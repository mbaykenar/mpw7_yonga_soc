magic
tech sky130B
magscale 12 1
timestamp 1598785131
<< metal5 >>
rect 0 100 20 105
rect 0 95 25 100
rect 0 85 30 95
rect 15 70 30 85
rect 15 60 35 70
rect 20 45 45 60
rect 15 35 35 45
rect 15 20 30 35
rect 0 10 30 20
rect 0 5 25 10
rect 0 0 20 5
<< properties >>
string FIXED_BBOX 0 -30 60 105
<< end >>
