VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO mba_core_region
  CLASS BLOCK ;
  FOREIGN mba_core_region ;
  ORIGIN 0.000 0.000 ;
  SIZE 1500.000 BY 1800.000 ;
  PIN boot_addr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1438.240 1500.000 1438.840 ;
    END
  END boot_addr_i[0]
  PIN boot_addr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 711.710 0.000 711.990 4.000 ;
    END
  END boot_addr_i[10]
  PIN boot_addr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 387.640 1500.000 388.240 ;
    END
  END boot_addr_i[11]
  PIN boot_addr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 190.070 1796.000 190.350 1800.000 ;
    END
  END boot_addr_i[12]
  PIN boot_addr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1251.240 1500.000 1251.840 ;
    END
  END boot_addr_i[13]
  PIN boot_addr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1298.840 1500.000 1299.440 ;
    END
  END boot_addr_i[14]
  PIN boot_addr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1098.240 4.000 1098.840 ;
    END
  END boot_addr_i[15]
  PIN boot_addr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 341.410 1796.000 341.690 1800.000 ;
    END
  END boot_addr_i[16]
  PIN boot_addr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1249.450 1796.000 1249.730 1800.000 ;
    END
  END boot_addr_i[17]
  PIN boot_addr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1017.610 1796.000 1017.890 1800.000 ;
    END
  END boot_addr_i[18]
  PIN boot_addr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 801.870 0.000 802.150 4.000 ;
    END
  END boot_addr_i[19]
  PIN boot_addr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1625.240 4.000 1625.840 ;
    END
  END boot_addr_i[1]
  PIN boot_addr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1278.440 4.000 1279.040 ;
    END
  END boot_addr_i[20]
  PIN boot_addr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 280.230 0.000 280.510 4.000 ;
    END
  END boot_addr_i[21]
  PIN boot_addr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 879.150 0.000 879.430 4.000 ;
    END
  END boot_addr_i[22]
  PIN boot_addr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 9.750 0.000 10.030 4.000 ;
    END
  END boot_addr_i[23]
  PIN boot_addr_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 408.040 4.000 408.640 ;
    END
  END boot_addr_i[24]
  PIN boot_addr_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1223.690 1796.000 1223.970 1800.000 ;
    END
  END boot_addr_i[25]
  PIN boot_addr_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 615.440 4.000 616.040 ;
    END
  END boot_addr_i[26]
  PIN boot_addr_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1046.590 1796.000 1046.870 1800.000 ;
    END
  END boot_addr_i[27]
  PIN boot_addr_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1329.440 1500.000 1330.040 ;
    END
  END boot_addr_i[28]
  PIN boot_addr_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 988.630 1796.000 988.910 1800.000 ;
    END
  END boot_addr_i[29]
  PIN boot_addr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1197.930 0.000 1198.210 4.000 ;
    END
  END boot_addr_i[2]
  PIN boot_addr_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 769.670 0.000 769.950 4.000 ;
    END
  END boot_addr_i[30]
  PIN boot_addr_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 927.450 0.000 927.730 4.000 ;
    END
  END boot_addr_i[31]
  PIN boot_addr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 377.440 1500.000 378.040 ;
    END
  END boot_addr_i[3]
  PIN boot_addr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1298.840 4.000 1299.440 ;
    END
  END boot_addr_i[4]
  PIN boot_addr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1485.840 4.000 1486.440 ;
    END
  END boot_addr_i[5]
  PIN boot_addr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 190.440 4.000 191.040 ;
    END
  END boot_addr_i[6]
  PIN boot_addr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 445.440 1500.000 446.040 ;
    END
  END boot_addr_i[7]
  PIN boot_addr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 629.040 1500.000 629.640 ;
    END
  END boot_addr_i[8]
  PIN boot_addr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 601.840 4.000 602.440 ;
    END
  END boot_addr_i[9]
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1011.170 1796.000 1011.450 1800.000 ;
    END
  END clk
  PIN clock_gating_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1132.240 1500.000 1132.840 ;
    END
  END clock_gating_i
  PIN core_busy_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1040.440 4.000 1041.040 ;
    END
  END core_busy_o
  PIN core_master_ar_addr[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.190 0.000 16.470 4.000 ;
    END
  END core_master_ar_addr[0]
  PIN core_master_ar_addr[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 591.640 1500.000 592.240 ;
    END
  END core_master_ar_addr[10]
  PIN core_master_ar_addr[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1492.640 1500.000 1493.240 ;
    END
  END core_master_ar_addr[11]
  PIN core_master_ar_addr[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1088.450 1796.000 1088.730 1800.000 ;
    END
  END core_master_ar_addr[12]
  PIN core_master_ar_addr[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 25.850 0.000 26.130 4.000 ;
    END
  END core_master_ar_addr[13]
  PIN core_master_ar_addr[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1315.840 1500.000 1316.440 ;
    END
  END core_master_ar_addr[14]
  PIN core_master_ar_addr[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 68.040 1500.000 68.640 ;
    END
  END core_master_ar_addr[15]
  PIN core_master_ar_addr[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 999.640 1500.000 1000.240 ;
    END
  END core_master_ar_addr[16]
  PIN core_master_ar_addr[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1285.240 1500.000 1285.840 ;
    END
  END core_master_ar_addr[17]
  PIN core_master_ar_addr[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 953.210 1796.000 953.490 1800.000 ;
    END
  END core_master_ar_addr[18]
  PIN core_master_ar_addr[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 953.210 0.000 953.490 4.000 ;
    END
  END core_master_ar_addr[19]
  PIN core_master_ar_addr[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1407.640 1500.000 1408.240 ;
    END
  END core_master_ar_addr[1]
  PIN core_master_ar_addr[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 553.930 0.000 554.210 4.000 ;
    END
  END core_master_ar_addr[20]
  PIN core_master_ar_addr[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1381.470 1796.000 1381.750 1800.000 ;
    END
  END core_master_ar_addr[21]
  PIN core_master_ar_addr[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 95.240 4.000 95.840 ;
    END
  END core_master_ar_addr[22]
  PIN core_master_ar_addr[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1499.440 4.000 1500.040 ;
    END
  END core_master_ar_addr[23]
  PIN core_master_ar_addr[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 737.470 1796.000 737.750 1800.000 ;
    END
  END core_master_ar_addr[24]
  PIN core_master_ar_addr[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 238.040 4.000 238.640 ;
    END
  END core_master_ar_addr[25]
  PIN core_master_ar_addr[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 386.490 1796.000 386.770 1800.000 ;
    END
  END core_master_ar_addr[26]
  PIN core_master_ar_addr[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 547.490 1796.000 547.770 1800.000 ;
    END
  END core_master_ar_addr[27]
  PIN core_master_ar_addr[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 112.240 4.000 112.840 ;
    END
  END core_master_ar_addr[28]
  PIN core_master_ar_addr[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 506.640 1500.000 507.240 ;
    END
  END core_master_ar_addr[29]
  PIN core_master_ar_addr[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1006.440 4.000 1007.040 ;
    END
  END core_master_ar_addr[2]
  PIN core_master_ar_addr[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 927.450 1796.000 927.730 1800.000 ;
    END
  END core_master_ar_addr[30]
  PIN core_master_ar_addr[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1744.240 4.000 1744.840 ;
    END
  END core_master_ar_addr[31]
  PIN core_master_ar_addr[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 799.040 4.000 799.640 ;
    END
  END core_master_ar_addr[3]
  PIN core_master_ar_addr[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 176.840 1500.000 177.440 ;
    END
  END core_master_ar_addr[4]
  PIN core_master_ar_addr[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1737.440 1500.000 1738.040 ;
    END
  END core_master_ar_addr[5]
  PIN core_master_ar_addr[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1434.840 4.000 1435.440 ;
    END
  END core_master_ar_addr[6]
  PIN core_master_ar_addr[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 669.850 1796.000 670.130 1800.000 ;
    END
  END core_master_ar_addr[7]
  PIN core_master_ar_addr[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 272.040 1500.000 272.640 ;
    END
  END core_master_ar_addr[8]
  PIN core_master_ar_addr[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1128.840 1500.000 1129.440 ;
    END
  END core_master_ar_addr[9]
  PIN core_master_ar_burst[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 180.410 1796.000 180.690 1800.000 ;
    END
  END core_master_ar_burst[0]
  PIN core_master_ar_burst[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 566.810 0.000 567.090 4.000 ;
    END
  END core_master_ar_burst[1]
  PIN core_master_ar_cache[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 870.440 4.000 871.040 ;
    END
  END core_master_ar_cache[0]
  PIN core_master_ar_cache[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 955.440 1500.000 956.040 ;
    END
  END core_master_ar_cache[1]
  PIN core_master_ar_cache[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 370.640 1500.000 371.240 ;
    END
  END core_master_ar_cache[2]
  PIN core_master_ar_cache[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1368.590 1796.000 1368.870 1800.000 ;
    END
  END core_master_ar_cache[3]
  PIN core_master_ar_id[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 769.670 1796.000 769.950 1800.000 ;
    END
  END core_master_ar_id[0]
  PIN core_master_ar_id[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1781.640 1500.000 1782.240 ;
    END
  END core_master_ar_id[1]
  PIN core_master_ar_id[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 743.910 1796.000 744.190 1800.000 ;
    END
  END core_master_ar_id[2]
  PIN core_master_ar_id[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1420.110 1796.000 1420.390 1800.000 ;
    END
  END core_master_ar_id[3]
  PIN core_master_ar_id[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 727.810 1796.000 728.090 1800.000 ;
    END
  END core_master_ar_id[4]
  PIN core_master_ar_id[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 409.030 1796.000 409.310 1800.000 ;
    END
  END core_master_ar_id[5]
  PIN core_master_ar_id[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1774.840 4.000 1775.440 ;
    END
  END core_master_ar_id[6]
  PIN core_master_ar_id[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1217.240 1500.000 1217.840 ;
    END
  END core_master_ar_id[7]
  PIN core_master_ar_id[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 877.240 1500.000 877.840 ;
    END
  END core_master_ar_id[8]
  PIN core_master_ar_id[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 363.840 4.000 364.440 ;
    END
  END core_master_ar_id[9]
  PIN core_master_ar_len[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 248.030 0.000 248.310 4.000 ;
    END
  END core_master_ar_len[0]
  PIN core_master_ar_len[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 20.440 4.000 21.040 ;
    END
  END core_master_ar_len[1]
  PIN core_master_ar_len[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 576.470 0.000 576.750 4.000 ;
    END
  END core_master_ar_len[2]
  PIN core_master_ar_len[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1785.040 4.000 1785.640 ;
    END
  END core_master_ar_len[3]
  PIN core_master_ar_len[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.970 0.000 13.250 4.000 ;
    END
  END core_master_ar_len[4]
  PIN core_master_ar_len[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 412.250 1796.000 412.530 1800.000 ;
    END
  END core_master_ar_len[5]
  PIN core_master_ar_len[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1133.530 1796.000 1133.810 1800.000 ;
    END
  END core_master_ar_len[6]
  PIN core_master_ar_len[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 202.950 0.000 203.230 4.000 ;
    END
  END core_master_ar_len[7]
  PIN core_master_ar_lock
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 901.040 4.000 901.640 ;
    END
  END core_master_ar_lock
  PIN core_master_ar_prot[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1145.840 4.000 1146.440 ;
    END
  END core_master_ar_prot[0]
  PIN core_master_ar_prot[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 557.640 1500.000 558.240 ;
    END
  END core_master_ar_prot[1]
  PIN core_master_ar_prot[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 251.640 1500.000 252.240 ;
    END
  END core_master_ar_prot[2]
  PIN core_master_ar_qos[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 605.450 0.000 605.730 4.000 ;
    END
  END core_master_ar_qos[0]
  PIN core_master_ar_qos[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 389.710 1796.000 389.990 1800.000 ;
    END
  END core_master_ar_qos[1]
  PIN core_master_ar_qos[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 839.840 4.000 840.440 ;
    END
  END core_master_ar_qos[2]
  PIN core_master_ar_qos[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 465.840 4.000 466.440 ;
    END
  END core_master_ar_qos[3]
  PIN core_master_ar_ready
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1094.840 1500.000 1095.440 ;
    END
  END core_master_ar_ready
  PIN core_master_ar_region[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 447.670 0.000 447.950 4.000 ;
    END
  END core_master_ar_region[0]
  PIN core_master_ar_region[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 315.650 0.000 315.930 4.000 ;
    END
  END core_master_ar_region[1]
  PIN core_master_ar_region[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 682.730 1796.000 683.010 1800.000 ;
    END
  END core_master_ar_region[2]
  PIN core_master_ar_region[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 148.210 1796.000 148.490 1800.000 ;
    END
  END core_master_ar_region[3]
  PIN core_master_ar_size[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1190.040 1500.000 1190.640 ;
    END
  END core_master_ar_size[0]
  PIN core_master_ar_size[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 931.640 4.000 932.240 ;
    END
  END core_master_ar_size[1]
  PIN core_master_ar_size[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1723.840 4.000 1724.440 ;
    END
  END core_master_ar_size[2]
  PIN core_master_ar_user[-1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 200.640 1500.000 201.240 ;
    END
  END core_master_ar_user[-1]
  PIN core_master_ar_user[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 710.640 4.000 711.240 ;
    END
  END core_master_ar_user[0]
  PIN core_master_ar_valid
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 731.030 1796.000 731.310 1800.000 ;
    END
  END core_master_ar_valid
  PIN core_master_aw_addr[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1497.390 1796.000 1497.670 1800.000 ;
    END
  END core_master_aw_addr[0]
  PIN core_master_aw_addr[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 272.040 4.000 272.640 ;
    END
  END core_master_aw_addr[10]
  PIN core_master_aw_addr[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 139.440 4.000 140.040 ;
    END
  END core_master_aw_addr[11]
  PIN core_master_aw_addr[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 834.070 0.000 834.350 4.000 ;
    END
  END core_master_aw_addr[12]
  PIN core_master_aw_addr[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 690.240 1500.000 690.840 ;
    END
  END core_master_aw_addr[13]
  PIN core_master_aw_addr[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 615.110 1796.000 615.390 1800.000 ;
    END
  END core_master_aw_addr[14]
  PIN core_master_aw_addr[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 153.040 1500.000 153.640 ;
    END
  END core_master_aw_addr[15]
  PIN core_master_aw_addr[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 979.240 1500.000 979.840 ;
    END
  END core_master_aw_addr[16]
  PIN core_master_aw_addr[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1285.240 4.000 1285.840 ;
    END
  END core_master_aw_addr[17]
  PIN core_master_aw_addr[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1655.840 4.000 1656.440 ;
    END
  END core_master_aw_addr[18]
  PIN core_master_aw_addr[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 721.370 1796.000 721.650 1800.000 ;
    END
  END core_master_aw_addr[19]
  PIN core_master_aw_addr[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 602.230 1796.000 602.510 1800.000 ;
    END
  END core_master_aw_addr[1]
  PIN core_master_aw_addr[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1026.840 1500.000 1027.440 ;
    END
  END core_master_aw_addr[20]
  PIN core_master_aw_addr[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 292.440 4.000 293.040 ;
    END
  END core_master_aw_addr[21]
  PIN core_master_aw_addr[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 336.640 1500.000 337.240 ;
    END
  END core_master_aw_addr[22]
  PIN core_master_aw_addr[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 937.110 1796.000 937.390 1800.000 ;
    END
  END core_master_aw_addr[23]
  PIN core_master_aw_addr[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 51.040 1500.000 51.640 ;
    END
  END core_master_aw_addr[24]
  PIN core_master_aw_addr[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1587.840 1500.000 1588.440 ;
    END
  END core_master_aw_addr[25]
  PIN core_master_aw_addr[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 901.040 1500.000 901.640 ;
    END
  END core_master_aw_addr[26]
  PIN core_master_aw_addr[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1377.040 1500.000 1377.640 ;
    END
  END core_master_aw_addr[27]
  PIN core_master_aw_addr[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 503.240 1500.000 503.840 ;
    END
  END core_master_aw_addr[28]
  PIN core_master_aw_addr[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1183.240 4.000 1183.840 ;
    END
  END core_master_aw_addr[29]
  PIN core_master_aw_addr[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 502.410 1796.000 502.690 1800.000 ;
    END
  END core_master_aw_addr[2]
  PIN core_master_aw_addr[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 27.240 1500.000 27.840 ;
    END
  END core_master_aw_addr[30]
  PIN core_master_aw_addr[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1077.840 4.000 1078.440 ;
    END
  END core_master_aw_addr[31]
  PIN core_master_aw_addr[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1540.240 1500.000 1540.840 ;
    END
  END core_master_aw_addr[3]
  PIN core_master_aw_addr[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1618.440 1500.000 1619.040 ;
    END
  END core_master_aw_addr[4]
  PIN core_master_aw_addr[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 78.240 4.000 78.840 ;
    END
  END core_master_aw_addr[5]
  PIN core_master_aw_addr[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 51.610 0.000 51.890 4.000 ;
    END
  END core_master_aw_addr[6]
  PIN core_master_aw_addr[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 697.040 4.000 697.640 ;
    END
  END core_master_aw_addr[7]
  PIN core_master_aw_addr[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1400.790 1796.000 1401.070 1800.000 ;
    END
  END core_master_aw_addr[8]
  PIN core_master_aw_addr[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 40.840 1500.000 41.440 ;
    END
  END core_master_aw_addr[9]
  PIN core_master_aw_burst[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 163.240 1500.000 163.840 ;
    END
  END core_master_aw_burst[0]
  PIN core_master_aw_burst[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 631.210 1796.000 631.490 1800.000 ;
    END
  END core_master_aw_burst[1]
  PIN core_master_aw_cache[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1127.090 0.000 1127.370 4.000 ;
    END
  END core_master_aw_cache[0]
  PIN core_master_aw_cache[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 814.750 0.000 815.030 4.000 ;
    END
  END core_master_aw_cache[1]
  PIN core_master_aw_cache[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 846.640 4.000 847.240 ;
    END
  END core_master_aw_cache[2]
  PIN core_master_aw_cache[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1247.840 4.000 1248.440 ;
    END
  END core_master_aw_cache[3]
  PIN core_master_aw_id[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1271.640 4.000 1272.240 ;
    END
  END core_master_aw_id[0]
  PIN core_master_aw_id[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 326.440 1500.000 327.040 ;
    END
  END core_master_aw_id[1]
  PIN core_master_aw_id[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1564.040 1500.000 1564.640 ;
    END
  END core_master_aw_id[2]
  PIN core_master_aw_id[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 61.240 1500.000 61.840 ;
    END
  END core_master_aw_id[3]
  PIN core_master_aw_id[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 394.440 4.000 395.040 ;
    END
  END core_master_aw_id[4]
  PIN core_master_aw_id[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 515.290 0.000 515.570 4.000 ;
    END
  END core_master_aw_id[5]
  PIN core_master_aw_id[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 567.840 1500.000 568.440 ;
    END
  END core_master_aw_id[6]
  PIN core_master_aw_id[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 132.110 1796.000 132.390 1800.000 ;
    END
  END core_master_aw_id[7]
  PIN core_master_aw_id[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 479.870 0.000 480.150 4.000 ;
    END
  END core_master_aw_id[8]
  PIN core_master_aw_id[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1696.640 4.000 1697.240 ;
    END
  END core_master_aw_id[9]
  PIN core_master_aw_len[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1230.130 0.000 1230.410 4.000 ;
    END
  END core_master_aw_len[0]
  PIN core_master_aw_len[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1734.040 4.000 1734.640 ;
    END
  END core_master_aw_len[1]
  PIN core_master_aw_len[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 860.240 4.000 860.840 ;
    END
  END core_master_aw_len[2]
  PIN core_master_aw_len[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 322.090 0.000 322.370 4.000 ;
    END
  END core_master_aw_len[3]
  PIN core_master_aw_len[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1751.040 4.000 1751.640 ;
    END
  END core_master_aw_len[4]
  PIN core_master_aw_len[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1123.870 1796.000 1124.150 1800.000 ;
    END
  END core_master_aw_len[5]
  PIN core_master_aw_len[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1451.840 4.000 1452.440 ;
    END
  END core_master_aw_len[6]
  PIN core_master_aw_len[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1040.150 0.000 1040.430 4.000 ;
    END
  END core_master_aw_len[7]
  PIN core_master_aw_lock
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 380.840 1500.000 381.440 ;
    END
  END core_master_aw_lock
  PIN core_master_aw_prot[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1003.040 4.000 1003.640 ;
    END
  END core_master_aw_prot[0]
  PIN core_master_aw_prot[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1332.840 4.000 1333.440 ;
    END
  END core_master_aw_prot[1]
  PIN core_master_aw_prot[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1036.930 1796.000 1037.210 1800.000 ;
    END
  END core_master_aw_prot[2]
  PIN core_master_aw_qos[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 718.150 1796.000 718.430 1800.000 ;
    END
  END core_master_aw_qos[0]
  PIN core_master_aw_qos[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 605.240 1500.000 605.840 ;
    END
  END core_master_aw_qos[1]
  PIN core_master_aw_qos[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 656.240 1500.000 656.840 ;
    END
  END core_master_aw_qos[2]
  PIN core_master_aw_qos[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 827.630 0.000 827.910 4.000 ;
    END
  END core_master_aw_qos[3]
  PIN core_master_aw_ready
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 187.040 4.000 187.640 ;
    END
  END core_master_aw_ready
  PIN core_master_aw_region[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 518.510 0.000 518.790 4.000 ;
    END
  END core_master_aw_region[0]
  PIN core_master_aw_region[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 469.240 1500.000 469.840 ;
    END
  END core_master_aw_region[1]
  PIN core_master_aw_region[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 564.440 1500.000 565.040 ;
    END
  END core_master_aw_region[2]
  PIN core_master_aw_region[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1098.240 1500.000 1098.840 ;
    END
  END core_master_aw_region[3]
  PIN core_master_aw_size[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1101.330 1796.000 1101.610 1800.000 ;
    END
  END core_master_aw_size[0]
  PIN core_master_aw_size[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 666.440 1500.000 667.040 ;
    END
  END core_master_aw_size[1]
  PIN core_master_aw_size[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 489.530 1796.000 489.810 1800.000 ;
    END
  END core_master_aw_size[2]
  PIN core_master_aw_user[-1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1078.790 1796.000 1079.070 1800.000 ;
    END
  END core_master_aw_user[-1]
  PIN core_master_aw_user[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 850.170 1796.000 850.450 1800.000 ;
    END
  END core_master_aw_user[0]
  PIN core_master_aw_valid
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1432.990 1796.000 1433.270 1800.000 ;
    END
  END core_master_aw_valid
  PIN core_master_b_id[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 621.550 1796.000 621.830 1800.000 ;
    END
  END core_master_b_id[0]
  PIN core_master_b_id[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 771.840 1500.000 772.440 ;
    END
  END core_master_b_id[1]
  PIN core_master_b_id[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1394.040 1500.000 1394.640 ;
    END
  END core_master_b_id[2]
  PIN core_master_b_id[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1494.170 0.000 1494.450 4.000 ;
    END
  END core_master_b_id[3]
  PIN core_master_b_id[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 455.640 4.000 456.240 ;
    END
  END core_master_b_id[4]
  PIN core_master_b_id[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1652.440 1500.000 1653.040 ;
    END
  END core_master_b_id[5]
  PIN core_master_b_id[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 632.440 1500.000 633.040 ;
    END
  END core_master_b_id[6]
  PIN core_master_b_id[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 508.850 0.000 509.130 4.000 ;
    END
  END core_master_b_id[7]
  PIN core_master_b_id[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1513.040 1500.000 1513.640 ;
    END
  END core_master_b_id[8]
  PIN core_master_b_id[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 136.040 1500.000 136.640 ;
    END
  END core_master_b_id[9]
  PIN core_master_b_ready
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1397.570 0.000 1397.850 4.000 ;
    END
  END core_master_b_ready
  PIN core_master_b_resp[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1162.840 4.000 1163.440 ;
    END
  END core_master_b_resp[0]
  PIN core_master_b_resp[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1669.440 4.000 1670.040 ;
    END
  END core_master_b_resp[1]
  PIN core_master_b_user[-1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 380.840 4.000 381.440 ;
    END
  END core_master_b_user[-1]
  PIN core_master_b_user[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 360.440 4.000 361.040 ;
    END
  END core_master_b_user[0]
  PIN core_master_b_valid
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1662.640 4.000 1663.240 ;
    END
  END core_master_b_valid
  PIN core_master_r_data[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1625.240 1500.000 1625.840 ;
    END
  END core_master_r_data[0]
  PIN core_master_r_data[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 282.240 4.000 282.840 ;
    END
  END core_master_r_data[10]
  PIN core_master_r_data[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 798.650 0.000 798.930 4.000 ;
    END
  END core_master_r_data[11]
  PIN core_master_r_data[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 615.440 1500.000 616.040 ;
    END
  END core_master_r_data[12]
  PIN core_master_r_data[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 383.270 1796.000 383.550 1800.000 ;
    END
  END core_master_r_data[13]
  PIN core_master_r_data[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1346.050 1796.000 1346.330 1800.000 ;
    END
  END core_master_r_data[14]
  PIN core_master_r_data[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 414.840 1500.000 415.440 ;
    END
  END core_master_r_data[15]
  PIN core_master_r_data[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1185.050 1796.000 1185.330 1800.000 ;
    END
  END core_master_r_data[16]
  PIN core_master_r_data[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1416.890 0.000 1417.170 4.000 ;
    END
  END core_master_r_data[17]
  PIN core_master_r_data[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 882.370 0.000 882.650 4.000 ;
    END
  END core_master_r_data[18]
  PIN core_master_r_data[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 486.310 0.000 486.590 4.000 ;
    END
  END core_master_r_data[19]
  PIN core_master_r_data[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1407.640 4.000 1408.240 ;
    END
  END core_master_r_data[1]
  PIN core_master_r_data[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 768.440 4.000 769.040 ;
    END
  END core_master_r_data[20]
  PIN core_master_r_data[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1065.910 0.000 1066.190 4.000 ;
    END
  END core_master_r_data[21]
  PIN core_master_r_data[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1074.440 4.000 1075.040 ;
    END
  END core_master_r_data[22]
  PIN core_master_r_data[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 557.150 0.000 557.430 4.000 ;
    END
  END core_master_r_data[23]
  PIN core_master_r_data[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 853.440 4.000 854.040 ;
    END
  END core_master_r_data[24]
  PIN core_master_r_data[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 589.350 0.000 589.630 4.000 ;
    END
  END core_master_r_data[25]
  PIN core_master_r_data[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 23.840 1500.000 24.440 ;
    END
  END core_master_r_data[26]
  PIN core_master_r_data[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1166.240 4.000 1166.840 ;
    END
  END core_master_r_data[27]
  PIN core_master_r_data[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1133.530 0.000 1133.810 4.000 ;
    END
  END core_master_r_data[28]
  PIN core_master_r_data[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1452.310 0.000 1452.590 4.000 ;
    END
  END core_master_r_data[29]
  PIN core_master_r_data[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1037.040 4.000 1037.640 ;
    END
  END core_master_r_data[2]
  PIN core_master_r_data[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 161.090 1796.000 161.370 1800.000 ;
    END
  END core_master_r_data[30]
  PIN core_master_r_data[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 595.790 1796.000 596.070 1800.000 ;
    END
  END core_master_r_data[31]
  PIN core_master_r_data[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1043.370 0.000 1043.650 4.000 ;
    END
  END core_master_r_data[32]
  PIN core_master_r_data[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 717.440 1500.000 718.040 ;
    END
  END core_master_r_data[33]
  PIN core_master_r_data[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 64.640 4.000 65.240 ;
    END
  END core_master_r_data[34]
  PIN core_master_r_data[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 260.910 1796.000 261.190 1800.000 ;
    END
  END core_master_r_data[35]
  PIN core_master_r_data[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 747.130 1796.000 747.410 1800.000 ;
    END
  END core_master_r_data[36]
  PIN core_master_r_data[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 834.070 1796.000 834.350 1800.000 ;
    END
  END core_master_r_data[37]
  PIN core_master_r_data[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 142.840 1500.000 143.440 ;
    END
  END core_master_r_data[38]
  PIN core_master_r_data[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 632.440 4.000 633.040 ;
    END
  END core_master_r_data[39]
  PIN core_master_r_data[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1024.050 1796.000 1024.330 1800.000 ;
    END
  END core_master_r_data[3]
  PIN core_master_r_data[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 457.330 1796.000 457.610 1800.000 ;
    END
  END core_master_r_data[40]
  PIN core_master_r_data[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 505.630 0.000 505.910 4.000 ;
    END
  END core_master_r_data[41]
  PIN core_master_r_data[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1747.640 4.000 1748.240 ;
    END
  END core_master_r_data[42]
  PIN core_master_r_data[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 472.640 4.000 473.240 ;
    END
  END core_master_r_data[43]
  PIN core_master_r_data[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 698.830 1796.000 699.110 1800.000 ;
    END
  END core_master_r_data[44]
  PIN core_master_r_data[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 483.090 0.000 483.370 4.000 ;
    END
  END core_master_r_data[45]
  PIN core_master_r_data[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1247.840 1500.000 1248.440 ;
    END
  END core_master_r_data[46]
  PIN core_master_r_data[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 193.840 4.000 194.440 ;
    END
  END core_master_r_data[47]
  PIN core_master_r_data[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 228.710 1796.000 228.990 1800.000 ;
    END
  END core_master_r_data[48]
  PIN core_master_r_data[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 106.350 1796.000 106.630 1800.000 ;
    END
  END core_master_r_data[49]
  PIN core_master_r_data[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 431.570 1796.000 431.850 1800.000 ;
    END
  END core_master_r_data[4]
  PIN core_master_r_data[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 695.610 1796.000 695.890 1800.000 ;
    END
  END core_master_r_data[50]
  PIN core_master_r_data[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 402.590 1796.000 402.870 1800.000 ;
    END
  END core_master_r_data[51]
  PIN core_master_r_data[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 863.050 1796.000 863.330 1800.000 ;
    END
  END core_master_r_data[52]
  PIN core_master_r_data[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 241.590 1796.000 241.870 1800.000 ;
    END
  END core_master_r_data[53]
  PIN core_master_r_data[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 44.240 4.000 44.840 ;
    END
  END core_master_r_data[54]
  PIN core_master_r_data[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 0.040 1500.000 0.640 ;
    END
  END core_master_r_data[55]
  PIN core_master_r_data[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1179.840 1500.000 1180.440 ;
    END
  END core_master_r_data[56]
  PIN core_master_r_data[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1237.640 1500.000 1238.240 ;
    END
  END core_master_r_data[57]
  PIN core_master_r_data[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1436.210 1796.000 1436.490 1800.000 ;
    END
  END core_master_r_data[58]
  PIN core_master_r_data[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1394.040 4.000 1394.640 ;
    END
  END core_master_r_data[59]
  PIN core_master_r_data[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 54.440 1500.000 55.040 ;
    END
  END core_master_r_data[5]
  PIN core_master_r_data[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 495.970 0.000 496.250 4.000 ;
    END
  END core_master_r_data[60]
  PIN core_master_r_data[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 778.640 4.000 779.240 ;
    END
  END core_master_r_data[61]
  PIN core_master_r_data[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1710.240 1500.000 1710.840 ;
    END
  END core_master_r_data[62]
  PIN core_master_r_data[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 659.640 4.000 660.240 ;
    END
  END core_master_r_data[63]
  PIN core_master_r_data[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 853.440 1500.000 854.040 ;
    END
  END core_master_r_data[6]
  PIN core_master_r_data[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 268.640 4.000 269.240 ;
    END
  END core_master_r_data[7]
  PIN core_master_r_data[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 985.410 0.000 985.690 4.000 ;
    END
  END core_master_r_data[8]
  PIN core_master_r_data[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 523.640 4.000 524.240 ;
    END
  END core_master_r_data[9]
  PIN core_master_r_id[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1343.040 1500.000 1343.640 ;
    END
  END core_master_r_id[0]
  PIN core_master_r_id[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 159.840 4.000 160.440 ;
    END
  END core_master_r_id[1]
  PIN core_master_r_id[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 833.040 1500.000 833.640 ;
    END
  END core_master_r_id[2]
  PIN core_master_r_id[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1781.640 4.000 1782.240 ;
    END
  END core_master_r_id[3]
  PIN core_master_r_id[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 795.430 0.000 795.710 4.000 ;
    END
  END core_master_r_id[4]
  PIN core_master_r_id[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 80.590 1796.000 80.870 1800.000 ;
    END
  END core_master_r_id[5]
  PIN core_master_r_id[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1246.230 0.000 1246.510 4.000 ;
    END
  END core_master_r_id[6]
  PIN core_master_r_id[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1587.840 4.000 1588.440 ;
    END
  END core_master_r_id[7]
  PIN core_master_r_id[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1703.440 4.000 1704.040 ;
    END
  END core_master_r_id[8]
  PIN core_master_r_id[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 418.240 1500.000 418.840 ;
    END
  END core_master_r_id[9]
  PIN core_master_r_last
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 586.130 0.000 586.410 4.000 ;
    END
  END core_master_r_last
  PIN core_master_r_ready
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 737.470 0.000 737.750 4.000 ;
    END
  END core_master_r_ready
  PIN core_master_r_resp[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1757.840 4.000 1758.440 ;
    END
  END core_master_r_resp[0]
  PIN core_master_r_resp[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 516.840 1500.000 517.440 ;
    END
  END core_master_r_resp[1]
  PIN core_master_r_user[-1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1465.440 1500.000 1466.040 ;
    END
  END core_master_r_user[-1]
  PIN core_master_r_user[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 392.930 0.000 393.210 4.000 ;
    END
  END core_master_r_user[0]
  PIN core_master_r_valid
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 186.850 0.000 187.130 4.000 ;
    END
  END core_master_r_valid
  PIN core_master_w_data[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1162.840 1500.000 1163.440 ;
    END
  END core_master_w_data[0]
  PIN core_master_w_data[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 988.630 0.000 988.910 4.000 ;
    END
  END core_master_w_data[10]
  PIN core_master_w_data[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1046.590 0.000 1046.870 4.000 ;
    END
  END core_master_w_data[11]
  PIN core_master_w_data[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1302.240 4.000 1302.840 ;
    END
  END core_master_w_data[12]
  PIN core_master_w_data[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 540.640 1500.000 541.240 ;
    END
  END core_master_w_data[13]
  PIN core_master_w_data[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 676.640 1500.000 677.240 ;
    END
  END core_master_w_data[14]
  PIN core_master_w_data[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 295.840 4.000 296.440 ;
    END
  END core_master_w_data[15]
  PIN core_master_w_data[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 642.640 1500.000 643.240 ;
    END
  END core_master_w_data[16]
  PIN core_master_w_data[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 805.090 0.000 805.370 4.000 ;
    END
  END core_master_w_data[17]
  PIN core_master_w_data[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1156.070 1796.000 1156.350 1800.000 ;
    END
  END core_master_w_data[18]
  PIN core_master_w_data[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 527.040 4.000 527.640 ;
    END
  END core_master_w_data[19]
  PIN core_master_w_data[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1014.390 0.000 1014.670 4.000 ;
    END
  END core_master_w_data[1]
  PIN core_master_w_data[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1145.840 1500.000 1146.440 ;
    END
  END core_master_w_data[20]
  PIN core_master_w_data[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1727.240 4.000 1727.840 ;
    END
  END core_master_w_data[21]
  PIN core_master_w_data[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 799.040 1500.000 799.640 ;
    END
  END core_master_w_data[22]
  PIN core_master_w_data[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 772.890 1796.000 773.170 1800.000 ;
    END
  END core_master_w_data[23]
  PIN core_master_w_data[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 938.440 4.000 939.040 ;
    END
  END core_master_w_data[24]
  PIN core_master_w_data[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 521.730 0.000 522.010 4.000 ;
    END
  END core_master_w_data[25]
  PIN core_master_w_data[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1482.440 1500.000 1483.040 ;
    END
  END core_master_w_data[26]
  PIN core_master_w_data[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 44.240 1500.000 44.840 ;
    END
  END core_master_w_data[27]
  PIN core_master_w_data[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 81.640 4.000 82.240 ;
    END
  END core_master_w_data[28]
  PIN core_master_w_data[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 3.440 1500.000 4.040 ;
    END
  END core_master_w_data[29]
  PIN core_master_w_data[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 989.440 4.000 990.040 ;
    END
  END core_master_w_data[2]
  PIN core_master_w_data[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 676.290 1796.000 676.570 1800.000 ;
    END
  END core_master_w_data[30]
  PIN core_master_w_data[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1067.640 4.000 1068.240 ;
    END
  END core_master_w_data[31]
  PIN core_master_w_data[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 170.040 4.000 170.640 ;
    END
  END core_master_w_data[32]
  PIN core_master_w_data[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 499.840 4.000 500.440 ;
    END
  END core_master_w_data[33]
  PIN core_master_w_data[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1710.240 4.000 1710.840 ;
    END
  END core_master_w_data[34]
  PIN core_master_w_data[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1368.590 0.000 1368.870 4.000 ;
    END
  END core_master_w_data[35]
  PIN core_master_w_data[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 941.840 4.000 942.440 ;
    END
  END core_master_w_data[36]
  PIN core_master_w_data[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 650.530 1796.000 650.810 1800.000 ;
    END
  END core_master_w_data[37]
  PIN core_master_w_data[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1795.240 1500.000 1795.840 ;
    END
  END core_master_w_data[38]
  PIN core_master_w_data[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1201.150 0.000 1201.430 4.000 ;
    END
  END core_master_w_data[39]
  PIN core_master_w_data[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 74.150 0.000 74.430 4.000 ;
    END
  END core_master_w_data[3]
  PIN core_master_w_data[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 640.870 0.000 641.150 4.000 ;
    END
  END core_master_w_data[40]
  PIN core_master_w_data[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1060.840 1500.000 1061.440 ;
    END
  END core_master_w_data[41]
  PIN core_master_w_data[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 483.090 1796.000 483.370 1800.000 ;
    END
  END core_master_w_data[42]
  PIN core_master_w_data[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 255.040 4.000 255.640 ;
    END
  END core_master_w_data[43]
  PIN core_master_w_data[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 537.240 4.000 537.840 ;
    END
  END core_master_w_data[44]
  PIN core_master_w_data[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 996.240 4.000 996.840 ;
    END
  END core_master_w_data[45]
  PIN core_master_w_data[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 647.310 1796.000 647.590 1800.000 ;
    END
  END core_master_w_data[46]
  PIN core_master_w_data[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 164.310 1796.000 164.590 1800.000 ;
    END
  END core_master_w_data[47]
  PIN core_master_w_data[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 386.490 0.000 386.770 4.000 ;
    END
  END core_master_w_data[48]
  PIN core_master_w_data[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 380.050 1796.000 380.330 1800.000 ;
    END
  END core_master_w_data[49]
  PIN core_master_w_data[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1481.290 1796.000 1481.570 1800.000 ;
    END
  END core_master_w_data[4]
  PIN core_master_w_data[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1397.440 4.000 1398.040 ;
    END
  END core_master_w_data[50]
  PIN core_master_w_data[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 615.110 0.000 615.390 4.000 ;
    END
  END core_master_w_data[51]
  PIN core_master_w_data[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1007.950 1796.000 1008.230 1800.000 ;
    END
  END core_master_w_data[52]
  PIN core_master_w_data[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 103.130 0.000 103.410 4.000 ;
    END
  END core_master_w_data[53]
  PIN core_master_w_data[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.710 1796.000 67.990 1800.000 ;
    END
  END core_master_w_data[54]
  PIN core_master_w_data[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1013.240 1500.000 1013.840 ;
    END
  END core_master_w_data[55]
  PIN core_master_w_data[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1516.440 4.000 1517.040 ;
    END
  END core_master_w_data[56]
  PIN core_master_w_data[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 824.410 1796.000 824.690 1800.000 ;
    END
  END core_master_w_data[57]
  PIN core_master_w_data[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 866.270 1796.000 866.550 1800.000 ;
    END
  END core_master_w_data[58]
  PIN core_master_w_data[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 428.350 1796.000 428.630 1800.000 ;
    END
  END core_master_w_data[59]
  PIN core_master_w_data[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 159.840 1500.000 160.440 ;
    END
  END core_master_w_data[5]
  PIN core_master_w_data[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1120.650 1796.000 1120.930 1800.000 ;
    END
  END core_master_w_data[60]
  PIN core_master_w_data[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1679.640 1500.000 1680.240 ;
    END
  END core_master_w_data[61]
  PIN core_master_w_data[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 724.590 1796.000 724.870 1800.000 ;
    END
  END core_master_w_data[62]
  PIN core_master_w_data[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1172.170 1796.000 1172.450 1800.000 ;
    END
  END core_master_w_data[63]
  PIN core_master_w_data[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 210.840 1500.000 211.440 ;
    END
  END core_master_w_data[6]
  PIN core_master_w_data[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 877.240 4.000 877.840 ;
    END
  END core_master_w_data[7]
  PIN core_master_w_data[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 207.440 4.000 208.040 ;
    END
  END core_master_w_data[8]
  PIN core_master_w_data[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 235.150 0.000 235.430 4.000 ;
    END
  END core_master_w_data[9]
  PIN core_master_w_last
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1252.670 1796.000 1252.950 1800.000 ;
    END
  END core_master_w_last
  PIN core_master_w_ready
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.530 1796.000 6.810 1800.000 ;
    END
  END core_master_w_ready
  PIN core_master_w_strb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 98.640 1500.000 99.240 ;
    END
  END core_master_w_strb[0]
  PIN core_master_w_strb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 829.640 1500.000 830.240 ;
    END
  END core_master_w_strb[1]
  PIN core_master_w_strb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 476.040 4.000 476.640 ;
    END
  END core_master_w_strb[2]
  PIN core_master_w_strb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1791.840 1500.000 1792.440 ;
    END
  END core_master_w_strb[3]
  PIN core_master_w_strb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 581.440 1500.000 582.040 ;
    END
  END core_master_w_strb[4]
  PIN core_master_w_strb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1689.840 1500.000 1690.440 ;
    END
  END core_master_w_strb[5]
  PIN core_master_w_strb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 405.810 1796.000 406.090 1800.000 ;
    END
  END core_master_w_strb[6]
  PIN core_master_w_strb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1204.370 1796.000 1204.650 1800.000 ;
    END
  END core_master_w_strb[7]
  PIN core_master_w_user[-1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 479.870 1796.000 480.150 1800.000 ;
    END
  END core_master_w_user[-1]
  PIN core_master_w_user[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 693.640 4.000 694.240 ;
    END
  END core_master_w_user[0]
  PIN core_master_w_valid
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 911.240 4.000 911.840 ;
    END
  END core_master_w_valid
  PIN data_slave_ar_addr[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1288.090 1796.000 1288.370 1800.000 ;
    END
  END data_slave_ar_addr[0]
  PIN data_slave_ar_addr[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 646.040 1500.000 646.640 ;
    END
  END data_slave_ar_addr[10]
  PIN data_slave_ar_addr[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 516.840 4.000 517.440 ;
    END
  END data_slave_ar_addr[11]
  PIN data_slave_ar_addr[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 257.690 1796.000 257.970 1800.000 ;
    END
  END data_slave_ar_addr[12]
  PIN data_slave_ar_addr[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 727.640 4.000 728.240 ;
    END
  END data_slave_ar_addr[13]
  PIN data_slave_ar_addr[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1261.440 1500.000 1262.040 ;
    END
  END data_slave_ar_addr[14]
  PIN data_slave_ar_addr[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1175.390 0.000 1175.670 4.000 ;
    END
  END data_slave_ar_addr[15]
  PIN data_slave_ar_addr[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 975.840 4.000 976.440 ;
    END
  END data_slave_ar_addr[16]
  PIN data_slave_ar_addr[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1105.040 4.000 1105.640 ;
    END
  END data_slave_ar_addr[17]
  PIN data_slave_ar_addr[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.270 1796.000 61.550 1800.000 ;
    END
  END data_slave_ar_addr[18]
  PIN data_slave_ar_addr[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 544.270 0.000 544.550 4.000 ;
    END
  END data_slave_ar_addr[19]
  PIN data_slave_ar_addr[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1233.350 0.000 1233.630 4.000 ;
    END
  END data_slave_ar_addr[1]
  PIN data_slave_ar_addr[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 938.440 1500.000 939.040 ;
    END
  END data_slave_ar_addr[20]
  PIN data_slave_ar_addr[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1638.840 4.000 1639.440 ;
    END
  END data_slave_ar_addr[21]
  PIN data_slave_ar_addr[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 17.040 1500.000 17.640 ;
    END
  END data_slave_ar_addr[22]
  PIN data_slave_ar_addr[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1391.130 1796.000 1391.410 1800.000 ;
    END
  END data_slave_ar_addr[23]
  PIN data_slave_ar_addr[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1356.640 4.000 1357.240 ;
    END
  END data_slave_ar_addr[24]
  PIN data_slave_ar_addr[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 431.840 4.000 432.440 ;
    END
  END data_slave_ar_addr[25]
  PIN data_slave_ar_addr[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 734.250 0.000 734.530 4.000 ;
    END
  END data_slave_ar_addr[26]
  PIN data_slave_ar_addr[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 285.640 4.000 286.240 ;
    END
  END data_slave_ar_addr[27]
  PIN data_slave_ar_addr[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 830.850 1796.000 831.130 1800.000 ;
    END
  END data_slave_ar_addr[28]
  PIN data_slave_ar_addr[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1271.640 1500.000 1272.240 ;
    END
  END data_slave_ar_addr[29]
  PIN data_slave_ar_addr[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1431.440 4.000 1432.040 ;
    END
  END data_slave_ar_addr[2]
  PIN data_slave_ar_addr[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 476.040 1500.000 476.640 ;
    END
  END data_slave_ar_addr[30]
  PIN data_slave_ar_addr[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 244.810 0.000 245.090 4.000 ;
    END
  END data_slave_ar_addr[31]
  PIN data_slave_ar_addr[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1672.840 4.000 1673.440 ;
    END
  END data_slave_ar_addr[3]
  PIN data_slave_ar_addr[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 409.030 0.000 409.310 4.000 ;
    END
  END data_slave_ar_addr[4]
  PIN data_slave_ar_addr[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1363.440 1500.000 1364.040 ;
    END
  END data_slave_ar_addr[5]
  PIN data_slave_ar_addr[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 459.040 4.000 459.640 ;
    END
  END data_slave_ar_addr[6]
  PIN data_slave_ar_addr[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 367.170 1796.000 367.450 1800.000 ;
    END
  END data_slave_ar_addr[7]
  PIN data_slave_ar_addr[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 318.870 1796.000 319.150 1800.000 ;
    END
  END data_slave_ar_addr[8]
  PIN data_slave_ar_addr[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 705.270 0.000 705.550 4.000 ;
    END
  END data_slave_ar_addr[9]
  PIN data_slave_ar_burst[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1577.640 4.000 1578.240 ;
    END
  END data_slave_ar_burst[0]
  PIN data_slave_ar_burst[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1497.390 0.000 1497.670 4.000 ;
    END
  END data_slave_ar_burst[1]
  PIN data_slave_ar_cache[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 222.270 0.000 222.550 4.000 ;
    END
  END data_slave_ar_cache[0]
  PIN data_slave_ar_cache[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1669.440 1500.000 1670.040 ;
    END
  END data_slave_ar_cache[1]
  PIN data_slave_ar_cache[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 367.240 1500.000 367.840 ;
    END
  END data_slave_ar_cache[2]
  PIN data_slave_ar_cache[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.530 0.000 6.810 4.000 ;
    END
  END data_slave_ar_cache[3]
  PIN data_slave_ar_id[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 550.710 1796.000 550.990 1800.000 ;
    END
  END data_slave_ar_id[0]
  PIN data_slave_ar_id[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1530.040 4.000 1530.640 ;
    END
  END data_slave_ar_id[1]
  PIN data_slave_ar_id[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 873.840 4.000 874.440 ;
    END
  END data_slave_ar_id[2]
  PIN data_slave_ar_id[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1645.640 1500.000 1646.240 ;
    END
  END data_slave_ar_id[3]
  PIN data_slave_ar_id[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 306.040 4.000 306.640 ;
    END
  END data_slave_ar_id[4]
  PIN data_slave_ar_id[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 316.240 4.000 316.840 ;
    END
  END data_slave_ar_id[5]
  PIN data_slave_ar_id[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 129.240 1500.000 129.840 ;
    END
  END data_slave_ar_id[6]
  PIN data_slave_ar_id[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1020.040 1500.000 1020.640 ;
    END
  END data_slave_ar_id[7]
  PIN data_slave_ar_id[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 802.440 4.000 803.040 ;
    END
  END data_slave_ar_id[8]
  PIN data_slave_ar_id[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 71.440 1500.000 72.040 ;
    END
  END data_slave_ar_id[9]
  PIN data_slave_ar_len[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 975.750 0.000 976.030 4.000 ;
    END
  END data_slave_ar_len[0]
  PIN data_slave_ar_len[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1365.370 0.000 1365.650 4.000 ;
    END
  END data_slave_ar_len[1]
  PIN data_slave_ar_len[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1455.240 1500.000 1455.840 ;
    END
  END data_slave_ar_len[2]
  PIN data_slave_ar_len[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1309.040 1500.000 1309.640 ;
    END
  END data_slave_ar_len[3]
  PIN data_slave_ar_len[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 598.440 1500.000 599.040 ;
    END
  END data_slave_ar_len[4]
  PIN data_slave_ar_len[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 959.650 1796.000 959.930 1800.000 ;
    END
  END data_slave_ar_len[5]
  PIN data_slave_ar_len[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 193.290 1796.000 193.570 1800.000 ;
    END
  END data_slave_ar_len[6]
  PIN data_slave_ar_len[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 493.040 4.000 493.640 ;
    END
  END data_slave_ar_len[7]
  PIN data_slave_ar_lock
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 846.950 1796.000 847.230 1800.000 ;
    END
  END data_slave_ar_lock
  PIN data_slave_ar_prot[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1057.440 4.000 1058.040 ;
    END
  END data_slave_ar_prot[0]
  PIN data_slave_ar_prot[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1333.170 1796.000 1333.450 1800.000 ;
    END
  END data_slave_ar_prot[1]
  PIN data_slave_ar_prot[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 125.840 1500.000 126.440 ;
    END
  END data_slave_ar_prot[2]
  PIN data_slave_ar_qos[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 914.570 0.000 914.850 4.000 ;
    END
  END data_slave_ar_qos[0]
  PIN data_slave_ar_qos[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 486.240 4.000 486.840 ;
    END
  END data_slave_ar_qos[1]
  PIN data_slave_ar_qos[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1519.840 1500.000 1520.440 ;
    END
  END data_slave_ar_qos[2]
  PIN data_slave_ar_qos[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 822.840 1500.000 823.440 ;
    END
  END data_slave_ar_qos[3]
  PIN data_slave_ar_ready
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 132.110 0.000 132.390 4.000 ;
    END
  END data_slave_ar_ready
  PIN data_slave_ar_region[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 193.840 1500.000 194.440 ;
    END
  END data_slave_ar_region[0]
  PIN data_slave_ar_region[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1128.840 4.000 1129.440 ;
    END
  END data_slave_ar_region[1]
  PIN data_slave_ar_region[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 10.240 4.000 10.840 ;
    END
  END data_slave_ar_region[2]
  PIN data_slave_ar_region[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1574.240 4.000 1574.840 ;
    END
  END data_slave_ar_region[3]
  PIN data_slave_ar_size[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 563.590 0.000 563.870 4.000 ;
    END
  END data_slave_ar_size[0]
  PIN data_slave_ar_size[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1397.570 1796.000 1397.850 1800.000 ;
    END
  END data_slave_ar_size[1]
  PIN data_slave_ar_size[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 999.640 4.000 1000.240 ;
    END
  END data_slave_ar_size[2]
  PIN data_slave_ar_user[-1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 802.440 1500.000 803.040 ;
    END
  END data_slave_ar_user[-1]
  PIN data_slave_ar_user[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 584.840 4.000 585.440 ;
    END
  END data_slave_ar_user[0]
  PIN data_slave_ar_valid
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1152.640 1500.000 1153.240 ;
    END
  END data_slave_ar_valid
  PIN data_slave_aw_addr[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1278.430 1796.000 1278.710 1800.000 ;
    END
  END data_slave_aw_addr[0]
  PIN data_slave_aw_addr[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1142.440 4.000 1143.040 ;
    END
  END data_slave_aw_addr[10]
  PIN data_slave_aw_addr[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 167.530 1796.000 167.810 1800.000 ;
    END
  END data_slave_aw_addr[11]
  PIN data_slave_aw_addr[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 531.390 0.000 531.670 4.000 ;
    END
  END data_slave_aw_addr[12]
  PIN data_slave_aw_addr[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 144.990 0.000 145.270 4.000 ;
    END
  END data_slave_aw_addr[13]
  PIN data_slave_aw_addr[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1091.440 4.000 1092.040 ;
    END
  END data_slave_aw_addr[14]
  PIN data_slave_aw_addr[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1349.840 4.000 1350.440 ;
    END
  END data_slave_aw_addr[15]
  PIN data_slave_aw_addr[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 442.040 4.000 442.640 ;
    END
  END data_slave_aw_addr[16]
  PIN data_slave_aw_addr[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 924.230 0.000 924.510 4.000 ;
    END
  END data_slave_aw_addr[17]
  PIN data_slave_aw_addr[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 962.870 1796.000 963.150 1800.000 ;
    END
  END data_slave_aw_addr[18]
  PIN data_slave_aw_addr[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 843.240 1500.000 843.840 ;
    END
  END data_slave_aw_addr[19]
  PIN data_slave_aw_addr[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1288.640 1500.000 1289.240 ;
    END
  END data_slave_aw_addr[1]
  PIN data_slave_aw_addr[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1223.690 0.000 1223.970 4.000 ;
    END
  END data_slave_aw_addr[20]
  PIN data_slave_aw_addr[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1207.590 1796.000 1207.870 1800.000 ;
    END
  END data_slave_aw_addr[21]
  PIN data_slave_aw_addr[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1169.640 4.000 1170.240 ;
    END
  END data_slave_aw_addr[22]
  PIN data_slave_aw_addr[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 402.590 0.000 402.870 4.000 ;
    END
  END data_slave_aw_addr[23]
  PIN data_slave_aw_addr[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 663.410 0.000 663.690 4.000 ;
    END
  END data_slave_aw_addr[24]
  PIN data_slave_aw_addr[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 892.030 0.000 892.310 4.000 ;
    END
  END data_slave_aw_addr[25]
  PIN data_slave_aw_addr[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 962.240 1500.000 962.840 ;
    END
  END data_slave_aw_addr[26]
  PIN data_slave_aw_addr[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1439.430 1796.000 1439.710 1800.000 ;
    END
  END data_slave_aw_addr[27]
  PIN data_slave_aw_addr[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1465.190 0.000 1465.470 4.000 ;
    END
  END data_slave_aw_addr[28]
  PIN data_slave_aw_addr[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1139.040 4.000 1139.640 ;
    END
  END data_slave_aw_addr[29]
  PIN data_slave_aw_addr[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 887.440 1500.000 888.040 ;
    END
  END data_slave_aw_addr[2]
  PIN data_slave_aw_addr[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 505.630 1796.000 505.910 1800.000 ;
    END
  END data_slave_aw_addr[30]
  PIN data_slave_aw_addr[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1278.430 0.000 1278.710 4.000 ;
    END
  END data_slave_aw_addr[31]
  PIN data_slave_aw_addr[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 872.710 0.000 872.990 4.000 ;
    END
  END data_slave_aw_addr[3]
  PIN data_slave_aw_addr[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1468.410 1796.000 1468.690 1800.000 ;
    END
  END data_slave_aw_addr[4]
  PIN data_slave_aw_addr[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 37.440 1500.000 38.040 ;
    END
  END data_slave_aw_addr[5]
  PIN data_slave_aw_addr[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 649.440 1500.000 650.040 ;
    END
  END data_slave_aw_addr[6]
  PIN data_slave_aw_addr[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 71.440 4.000 72.040 ;
    END
  END data_slave_aw_addr[7]
  PIN data_slave_aw_addr[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1757.840 1500.000 1758.440 ;
    END
  END data_slave_aw_addr[8]
  PIN data_slave_aw_addr[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 418.240 4.000 418.840 ;
    END
  END data_slave_aw_addr[9]
  PIN data_slave_aw_burst[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1655.840 1500.000 1656.440 ;
    END
  END data_slave_aw_burst[0]
  PIN data_slave_aw_burst[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 904.440 4.000 905.040 ;
    END
  END data_slave_aw_burst[1]
  PIN data_slave_aw_cache[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.970 1796.000 13.250 1800.000 ;
    END
  END data_slave_aw_cache[0]
  PIN data_slave_aw_cache[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 90.250 1796.000 90.530 1800.000 ;
    END
  END data_slave_aw_cache[1]
  PIN data_slave_aw_cache[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1332.840 1500.000 1333.440 ;
    END
  END data_slave_aw_cache[2]
  PIN data_slave_aw_cache[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1604.840 4.000 1605.440 ;
    END
  END data_slave_aw_cache[3]
  PIN data_slave_aw_id[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 227.840 4.000 228.440 ;
    END
  END data_slave_aw_id[0]
  PIN data_slave_aw_id[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 647.310 0.000 647.590 4.000 ;
    END
  END data_slave_aw_id[1]
  PIN data_slave_aw_id[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 666.440 4.000 667.040 ;
    END
  END data_slave_aw_id[2]
  PIN data_slave_aw_id[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1353.240 4.000 1353.840 ;
    END
  END data_slave_aw_id[3]
  PIN data_slave_aw_id[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 415.470 0.000 415.750 4.000 ;
    END
  END data_slave_aw_id[4]
  PIN data_slave_aw_id[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 856.610 0.000 856.890 4.000 ;
    END
  END data_slave_aw_id[5]
  PIN data_slave_aw_id[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1027.270 1796.000 1027.550 1800.000 ;
    END
  END data_slave_aw_id[6]
  PIN data_slave_aw_id[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 656.970 0.000 657.250 4.000 ;
    END
  END data_slave_aw_id[7]
  PIN data_slave_aw_id[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1077.840 1500.000 1078.440 ;
    END
  END data_slave_aw_id[8]
  PIN data_slave_aw_id[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 370.390 0.000 370.670 4.000 ;
    END
  END data_slave_aw_id[9]
  PIN data_slave_aw_len[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 795.640 1500.000 796.240 ;
    END
  END data_slave_aw_len[0]
  PIN data_slave_aw_len[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1130.310 1796.000 1130.590 1800.000 ;
    END
  END data_slave_aw_len[1]
  PIN data_slave_aw_len[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1072.350 0.000 1072.630 4.000 ;
    END
  END data_slave_aw_len[2]
  PIN data_slave_aw_len[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1108.440 4.000 1109.040 ;
    END
  END data_slave_aw_len[3]
  PIN data_slave_aw_len[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 578.040 1500.000 578.640 ;
    END
  END data_slave_aw_len[4]
  PIN data_slave_aw_len[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 907.840 1500.000 908.440 ;
    END
  END data_slave_aw_len[5]
  PIN data_slave_aw_len[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 78.240 1500.000 78.840 ;
    END
  END data_slave_aw_len[6]
  PIN data_slave_aw_len[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 499.190 0.000 499.470 4.000 ;
    END
  END data_slave_aw_len[7]
  PIN data_slave_aw_lock
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 108.840 4.000 109.440 ;
    END
  END data_slave_aw_lock
  PIN data_slave_aw_prot[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.050 1796.000 58.330 1800.000 ;
    END
  END data_slave_aw_prot[0]
  PIN data_slave_aw_prot[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 689.170 0.000 689.450 4.000 ;
    END
  END data_slave_aw_prot[1]
  PIN data_slave_aw_prot[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 197.240 1500.000 197.840 ;
    END
  END data_slave_aw_prot[2]
  PIN data_slave_aw_qos[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 231.240 4.000 231.840 ;
    END
  END data_slave_aw_qos[0]
  PIN data_slave_aw_qos[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1730.640 4.000 1731.240 ;
    END
  END data_slave_aw_qos[1]
  PIN data_slave_aw_qos[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 943.550 0.000 943.830 4.000 ;
    END
  END data_slave_aw_qos[2]
  PIN data_slave_aw_qos[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 148.210 0.000 148.490 4.000 ;
    END
  END data_slave_aw_qos[3]
  PIN data_slave_aw_ready
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1502.840 1500.000 1503.440 ;
    END
  END data_slave_aw_ready
  PIN data_slave_aw_region[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 880.640 1500.000 881.240 ;
    END
  END data_slave_aw_region[0]
  PIN data_slave_aw_region[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1013.240 4.000 1013.840 ;
    END
  END data_slave_aw_region[1]
  PIN data_slave_aw_region[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 573.250 1796.000 573.530 1800.000 ;
    END
  END data_slave_aw_region[2]
  PIN data_slave_aw_region[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 798.650 1796.000 798.930 1800.000 ;
    END
  END data_slave_aw_region[3]
  PIN data_slave_aw_size[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1584.440 4.000 1585.040 ;
    END
  END data_slave_aw_size[0]
  PIN data_slave_aw_size[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 982.190 1796.000 982.470 1800.000 ;
    END
  END data_slave_aw_size[1]
  PIN data_slave_aw_size[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1214.030 1796.000 1214.310 1800.000 ;
    END
  END data_slave_aw_size[2]
  PIN data_slave_aw_user[-1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 618.330 0.000 618.610 4.000 ;
    END
  END data_slave_aw_user[-1]
  PIN data_slave_aw_user[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 946.770 0.000 947.050 4.000 ;
    END
  END data_slave_aw_user[0]
  PIN data_slave_aw_valid
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1686.440 1500.000 1687.040 ;
    END
  END data_slave_aw_valid
  PIN data_slave_b_id[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1125.440 1500.000 1126.040 ;
    END
  END data_slave_b_id[0]
  PIN data_slave_b_id[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 659.640 1500.000 660.240 ;
    END
  END data_slave_b_id[1]
  PIN data_slave_b_id[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 389.710 0.000 389.990 4.000 ;
    END
  END data_slave_b_id[2]
  PIN data_slave_b_id[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 676.290 0.000 676.570 4.000 ;
    END
  END data_slave_b_id[3]
  PIN data_slave_b_id[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1458.640 4.000 1459.240 ;
    END
  END data_slave_b_id[4]
  PIN data_slave_b_id[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1423.330 1796.000 1423.610 1800.000 ;
    END
  END data_slave_b_id[5]
  PIN data_slave_b_id[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 228.710 0.000 228.990 4.000 ;
    END
  END data_slave_b_id[6]
  PIN data_slave_b_id[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 244.840 4.000 245.440 ;
    END
  END data_slave_b_id[7]
  PIN data_slave_b_id[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 144.990 1796.000 145.270 1800.000 ;
    END
  END data_slave_b_id[8]
  PIN data_slave_b_id[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.050 0.000 58.330 4.000 ;
    END
  END data_slave_b_id[9]
  PIN data_slave_b_ready
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1062.690 1796.000 1062.970 1800.000 ;
    END
  END data_slave_b_ready
  PIN data_slave_b_resp[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 948.640 4.000 949.240 ;
    END
  END data_slave_b_resp[0]
  PIN data_slave_b_resp[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 537.830 0.000 538.110 4.000 ;
    END
  END data_slave_b_resp[1]
  PIN data_slave_b_user[-1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 840.510 1796.000 840.790 1800.000 ;
    END
  END data_slave_b_user[-1]
  PIN data_slave_b_user[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 627.990 1796.000 628.270 1800.000 ;
    END
  END data_slave_b_user[0]
  PIN data_slave_b_valid
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 91.840 4.000 92.440 ;
    END
  END data_slave_b_valid
  PIN data_slave_r_data[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 77.370 0.000 77.650 4.000 ;
    END
  END data_slave_r_data[0]
  PIN data_slave_r_data[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 222.270 1796.000 222.550 1800.000 ;
    END
  END data_slave_r_data[10]
  PIN data_slave_r_data[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 513.440 4.000 514.040 ;
    END
  END data_slave_r_data[11]
  PIN data_slave_r_data[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1533.440 1500.000 1534.040 ;
    END
  END data_slave_r_data[12]
  PIN data_slave_r_data[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1313.850 1796.000 1314.130 1800.000 ;
    END
  END data_slave_r_data[13]
  PIN data_slave_r_data[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1258.040 4.000 1258.640 ;
    END
  END data_slave_r_data[14]
  PIN data_slave_r_data[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1050.640 4.000 1051.240 ;
    END
  END data_slave_r_data[15]
  PIN data_slave_r_data[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1017.610 0.000 1017.890 4.000 ;
    END
  END data_slave_r_data[16]
  PIN data_slave_r_data[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 940.330 0.000 940.610 4.000 ;
    END
  END data_slave_r_data[17]
  PIN data_slave_r_data[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 248.240 1500.000 248.840 ;
    END
  END data_slave_r_data[18]
  PIN data_slave_r_data[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1191.490 1796.000 1191.770 1800.000 ;
    END
  END data_slave_r_data[19]
  PIN data_slave_r_data[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 821.190 0.000 821.470 4.000 ;
    END
  END data_slave_r_data[1]
  PIN data_slave_r_data[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 685.950 0.000 686.230 4.000 ;
    END
  END data_slave_r_data[20]
  PIN data_slave_r_data[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1065.910 1796.000 1066.190 1800.000 ;
    END
  END data_slave_r_data[21]
  PIN data_slave_r_data[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 363.950 0.000 364.230 4.000 ;
    END
  END data_slave_r_data[22]
  PIN data_slave_r_data[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 624.770 1796.000 625.050 1800.000 ;
    END
  END data_slave_r_data[23]
  PIN data_slave_r_data[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 363.950 1796.000 364.230 1800.000 ;
    END
  END data_slave_r_data[24]
  PIN data_slave_r_data[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1234.240 4.000 1234.840 ;
    END
  END data_slave_r_data[25]
  PIN data_slave_r_data[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 277.010 0.000 277.290 4.000 ;
    END
  END data_slave_r_data[26]
  PIN data_slave_r_data[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 531.390 1796.000 531.670 1800.000 ;
    END
  END data_slave_r_data[27]
  PIN data_slave_r_data[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1484.510 1796.000 1484.790 1800.000 ;
    END
  END data_slave_r_data[28]
  PIN data_slave_r_data[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 720.840 4.000 721.440 ;
    END
  END data_slave_r_data[29]
  PIN data_slave_r_data[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3.310 1796.000 3.590 1800.000 ;
    END
  END data_slave_r_data[2]
  PIN data_slave_r_data[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1543.640 4.000 1544.240 ;
    END
  END data_slave_r_data[30]
  PIN data_slave_r_data[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 257.690 0.000 257.970 4.000 ;
    END
  END data_slave_r_data[31]
  PIN data_slave_r_data[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1101.330 0.000 1101.610 4.000 ;
    END
  END data_slave_r_data[32]
  PIN data_slave_r_data[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 415.470 1796.000 415.750 1800.000 ;
    END
  END data_slave_r_data[33]
  PIN data_slave_r_data[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 17.040 4.000 17.640 ;
    END
  END data_slave_r_data[34]
  PIN data_slave_r_data[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1621.840 4.000 1622.440 ;
    END
  END data_slave_r_data[35]
  PIN data_slave_r_data[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1342.830 1796.000 1343.110 1800.000 ;
    END
  END data_slave_r_data[36]
  PIN data_slave_r_data[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1307.410 0.000 1307.690 4.000 ;
    END
  END data_slave_r_data[37]
  PIN data_slave_r_data[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 570.030 1796.000 570.310 1800.000 ;
    END
  END data_slave_r_data[38]
  PIN data_slave_r_data[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1040.440 1500.000 1041.040 ;
    END
  END data_slave_r_data[39]
  PIN data_slave_r_data[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 700.440 4.000 701.040 ;
    END
  END data_slave_r_data[3]
  PIN data_slave_r_data[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1020.830 0.000 1021.110 4.000 ;
    END
  END data_slave_r_data[40]
  PIN data_slave_r_data[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1165.730 1796.000 1166.010 1800.000 ;
    END
  END data_slave_r_data[41]
  PIN data_slave_r_data[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 618.840 4.000 619.440 ;
    END
  END data_slave_r_data[42]
  PIN data_slave_r_data[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 90.250 0.000 90.530 4.000 ;
    END
  END data_slave_r_data[43]
  PIN data_slave_r_data[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 727.640 1500.000 728.240 ;
    END
  END data_slave_r_data[44]
  PIN data_slave_r_data[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 441.230 1796.000 441.510 1800.000 ;
    END
  END data_slave_r_data[45]
  PIN data_slave_r_data[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1082.010 1796.000 1082.290 1800.000 ;
    END
  END data_slave_r_data[46]
  PIN data_slave_r_data[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 392.930 1796.000 393.210 1800.000 ;
    END
  END data_slave_r_data[47]
  PIN data_slave_r_data[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1036.930 0.000 1037.210 4.000 ;
    END
  END data_slave_r_data[48]
  PIN data_slave_r_data[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1462.040 4.000 1462.640 ;
    END
  END data_slave_r_data[49]
  PIN data_slave_r_data[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 693.640 1500.000 694.240 ;
    END
  END data_slave_r_data[4]
  PIN data_slave_r_data[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 700.440 1500.000 701.040 ;
    END
  END data_slave_r_data[50]
  PIN data_slave_r_data[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1492.640 4.000 1493.240 ;
    END
  END data_slave_r_data[51]
  PIN data_slave_r_data[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 697.040 1500.000 697.640 ;
    END
  END data_slave_r_data[52]
  PIN data_slave_r_data[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1390.640 4.000 1391.240 ;
    END
  END data_slave_r_data[53]
  PIN data_slave_r_data[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1178.610 1796.000 1178.890 1800.000 ;
    END
  END data_slave_r_data[54]
  PIN data_slave_r_data[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 811.530 1796.000 811.810 1800.000 ;
    END
  END data_slave_r_data[55]
  PIN data_slave_r_data[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 315.650 1796.000 315.930 1800.000 ;
    END
  END data_slave_r_data[56]
  PIN data_slave_r_data[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1333.170 0.000 1333.450 4.000 ;
    END
  END data_slave_r_data[57]
  PIN data_slave_r_data[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 637.650 0.000 637.930 4.000 ;
    END
  END data_slave_r_data[58]
  PIN data_slave_r_data[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 850.170 0.000 850.450 4.000 ;
    END
  END data_slave_r_data[59]
  PIN data_slave_r_data[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 489.640 1500.000 490.240 ;
    END
  END data_slave_r_data[5]
  PIN data_slave_r_data[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 445.440 4.000 446.040 ;
    END
  END data_slave_r_data[60]
  PIN data_slave_r_data[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1004.730 1796.000 1005.010 1800.000 ;
    END
  END data_slave_r_data[61]
  PIN data_slave_r_data[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 387.640 4.000 388.240 ;
    END
  END data_slave_r_data[62]
  PIN data_slave_r_data[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1188.270 0.000 1188.550 4.000 ;
    END
  END data_slave_r_data[63]
  PIN data_slave_r_data[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 686.840 4.000 687.440 ;
    END
  END data_slave_r_data[6]
  PIN data_slave_r_data[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1434.840 1500.000 1435.440 ;
    END
  END data_slave_r_data[7]
  PIN data_slave_r_data[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1788.440 1500.000 1789.040 ;
    END
  END data_slave_r_data[8]
  PIN data_slave_r_data[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 196.510 0.000 196.790 4.000 ;
    END
  END data_slave_r_data[9]
  PIN data_slave_r_id[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1101.640 1500.000 1102.240 ;
    END
  END data_slave_r_id[0]
  PIN data_slave_r_id[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 792.210 1796.000 792.490 1800.000 ;
    END
  END data_slave_r_id[1]
  PIN data_slave_r_id[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 863.050 0.000 863.330 4.000 ;
    END
  END data_slave_r_id[2]
  PIN data_slave_r_id[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 826.240 4.000 826.840 ;
    END
  END data_slave_r_id[3]
  PIN data_slave_r_id[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1300.970 0.000 1301.250 4.000 ;
    END
  END data_slave_r_id[4]
  PIN data_slave_r_id[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1747.640 1500.000 1748.240 ;
    END
  END data_slave_r_id[5]
  PIN data_slave_r_id[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 772.890 0.000 773.170 4.000 ;
    END
  END data_slave_r_id[6]
  PIN data_slave_r_id[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1659.240 1500.000 1659.840 ;
    END
  END data_slave_r_id[7]
  PIN data_slave_r_id[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 567.840 4.000 568.440 ;
    END
  END data_slave_r_id[8]
  PIN data_slave_r_id[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1371.810 0.000 1372.090 4.000 ;
    END
  END data_slave_r_id[9]
  PIN data_slave_r_last
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1387.910 1796.000 1388.190 1800.000 ;
    END
  END data_slave_r_last
  PIN data_slave_r_ready
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 544.040 1500.000 544.640 ;
    END
  END data_slave_r_ready
  PIN data_slave_r_resp[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 985.410 1796.000 985.690 1800.000 ;
    END
  END data_slave_r_resp[0]
  PIN data_slave_r_resp[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 319.640 1500.000 320.240 ;
    END
  END data_slave_r_resp[1]
  PIN data_slave_r_user[-1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 690.240 4.000 690.840 ;
    END
  END data_slave_r_user[-1]
  PIN data_slave_r_user[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 177.190 1796.000 177.470 1800.000 ;
    END
  END data_slave_r_user[0]
  PIN data_slave_r_valid
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1394.350 0.000 1394.630 4.000 ;
    END
  END data_slave_r_valid
  PIN data_slave_w_data[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1713.640 4.000 1714.240 ;
    END
  END data_slave_w_data[0]
  PIN data_slave_w_data[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1339.640 1500.000 1340.240 ;
    END
  END data_slave_w_data[10]
  PIN data_slave_w_data[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 949.990 0.000 950.270 4.000 ;
    END
  END data_slave_w_data[11]
  PIN data_slave_w_data[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1056.250 1796.000 1056.530 1800.000 ;
    END
  END data_slave_w_data[12]
  PIN data_slave_w_data[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 642.640 4.000 643.240 ;
    END
  END data_slave_w_data[13]
  PIN data_slave_w_data[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.170 1796.000 45.450 1800.000 ;
    END
  END data_slave_w_data[14]
  PIN data_slave_w_data[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1342.830 0.000 1343.110 4.000 ;
    END
  END data_slave_w_data[15]
  PIN data_slave_w_data[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 917.790 0.000 918.070 4.000 ;
    END
  END data_slave_w_data[16]
  PIN data_slave_w_data[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 323.040 1500.000 323.640 ;
    END
  END data_slave_w_data[17]
  PIN data_slave_w_data[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 533.840 1500.000 534.440 ;
    END
  END data_slave_w_data[18]
  PIN data_slave_w_data[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1349.840 1500.000 1350.440 ;
    END
  END data_slave_w_data[19]
  PIN data_slave_w_data[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.470 1796.000 93.750 1800.000 ;
    END
  END data_slave_w_data[1]
  PIN data_slave_w_data[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 768.440 1500.000 769.040 ;
    END
  END data_slave_w_data[20]
  PIN data_slave_w_data[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1220.640 4.000 1221.240 ;
    END
  END data_slave_w_data[21]
  PIN data_slave_w_data[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 401.240 1500.000 401.840 ;
    END
  END data_slave_w_data[22]
  PIN data_slave_w_data[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 640.870 1796.000 641.150 1800.000 ;
    END
  END data_slave_w_data[23]
  PIN data_slave_w_data[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 708.490 0.000 708.770 4.000 ;
    END
  END data_slave_w_data[24]
  PIN data_slave_w_data[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1030.240 4.000 1030.840 ;
    END
  END data_slave_w_data[25]
  PIN data_slave_w_data[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 452.240 1500.000 452.840 ;
    END
  END data_slave_w_data[26]
  PIN data_slave_w_data[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 663.040 4.000 663.640 ;
    END
  END data_slave_w_data[27]
  PIN data_slave_w_data[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1107.770 0.000 1108.050 4.000 ;
    END
  END data_slave_w_data[28]
  PIN data_slave_w_data[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1210.810 0.000 1211.090 4.000 ;
    END
  END data_slave_w_data[29]
  PIN data_slave_w_data[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 581.440 4.000 582.040 ;
    END
  END data_slave_w_data[2]
  PIN data_slave_w_data[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 346.840 4.000 347.440 ;
    END
  END data_slave_w_data[30]
  PIN data_slave_w_data[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.390 0.000 48.670 4.000 ;
    END
  END data_slave_w_data[31]
  PIN data_slave_w_data[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1727.240 1500.000 1727.840 ;
    END
  END data_slave_w_data[32]
  PIN data_slave_w_data[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 714.040 4.000 714.640 ;
    END
  END data_slave_w_data[33]
  PIN data_slave_w_data[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 354.290 1796.000 354.570 1800.000 ;
    END
  END data_slave_w_data[34]
  PIN data_slave_w_data[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 106.350 0.000 106.630 4.000 ;
    END
  END data_slave_w_data[35]
  PIN data_slave_w_data[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1043.840 4.000 1044.440 ;
    END
  END data_slave_w_data[36]
  PIN data_slave_w_data[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 170.750 1796.000 171.030 1800.000 ;
    END
  END data_slave_w_data[37]
  PIN data_slave_w_data[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 95.240 1500.000 95.840 ;
    END
  END data_slave_w_data[38]
  PIN data_slave_w_data[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 618.840 1500.000 619.440 ;
    END
  END data_slave_w_data[39]
  PIN data_slave_w_data[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 541.050 0.000 541.330 4.000 ;
    END
  END data_slave_w_data[3]
  PIN data_slave_w_data[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 979.240 4.000 979.840 ;
    END
  END data_slave_w_data[40]
  PIN data_slave_w_data[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1115.240 4.000 1115.840 ;
    END
  END data_slave_w_data[41]
  PIN data_slave_w_data[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1506.240 1500.000 1506.840 ;
    END
  END data_slave_w_data[42]
  PIN data_slave_w_data[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 183.640 4.000 184.240 ;
    END
  END data_slave_w_data[43]
  PIN data_slave_w_data[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 238.370 1796.000 238.650 1800.000 ;
    END
  END data_slave_w_data[44]
  PIN data_slave_w_data[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 305.990 0.000 306.270 4.000 ;
    END
  END data_slave_w_data[45]
  PIN data_slave_w_data[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1373.640 4.000 1374.240 ;
    END
  END data_slave_w_data[46]
  PIN data_slave_w_data[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1676.240 4.000 1676.840 ;
    END
  END data_slave_w_data[47]
  PIN data_slave_w_data[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 579.690 0.000 579.970 4.000 ;
    END
  END data_slave_w_data[48]
  PIN data_slave_w_data[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 592.570 0.000 592.850 4.000 ;
    END
  END data_slave_w_data[49]
  PIN data_slave_w_data[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.510 1796.000 35.790 1800.000 ;
    END
  END data_slave_w_data[4]
  PIN data_slave_w_data[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 584.840 1500.000 585.440 ;
    END
  END data_slave_w_data[50]
  PIN data_slave_w_data[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 353.640 1500.000 354.240 ;
    END
  END data_slave_w_data[51]
  PIN data_slave_w_data[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 760.010 1796.000 760.290 1800.000 ;
    END
  END data_slave_w_data[52]
  PIN data_slave_w_data[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 54.440 4.000 55.040 ;
    END
  END data_slave_w_data[53]
  PIN data_slave_w_data[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 394.440 1500.000 395.040 ;
    END
  END data_slave_w_data[54]
  PIN data_slave_w_data[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 586.130 1796.000 586.410 1800.000 ;
    END
  END data_slave_w_data[55]
  PIN data_slave_w_data[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1355.710 0.000 1355.990 4.000 ;
    END
  END data_slave_w_data[56]
  PIN data_slave_w_data[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 334.970 1796.000 335.250 1800.000 ;
    END
  END data_slave_w_data[57]
  PIN data_slave_w_data[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 996.240 1500.000 996.840 ;
    END
  END data_slave_w_data[58]
  PIN data_slave_w_data[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 357.040 1500.000 357.640 ;
    END
  END data_slave_w_data[59]
  PIN data_slave_w_data[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1098.110 1796.000 1098.390 1800.000 ;
    END
  END data_slave_w_data[5]
  PIN data_slave_w_data[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1014.390 1796.000 1014.670 1800.000 ;
    END
  END data_slave_w_data[60]
  PIN data_slave_w_data[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 530.440 1500.000 531.040 ;
    END
  END data_slave_w_data[61]
  PIN data_slave_w_data[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1094.890 1796.000 1095.170 1800.000 ;
    END
  END data_slave_w_data[62]
  PIN data_slave_w_data[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1421.240 4.000 1421.840 ;
    END
  END data_slave_w_data[63]
  PIN data_slave_w_data[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 908.130 1796.000 908.410 1800.000 ;
    END
  END data_slave_w_data[6]
  PIN data_slave_w_data[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 270.570 1796.000 270.850 1800.000 ;
    END
  END data_slave_w_data[7]
  PIN data_slave_w_data[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1489.240 1500.000 1489.840 ;
    END
  END data_slave_w_data[8]
  PIN data_slave_w_data[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 808.310 1796.000 808.590 1800.000 ;
    END
  END data_slave_w_data[9]
  PIN data_slave_w_last
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 328.530 0.000 328.810 4.000 ;
    END
  END data_slave_w_last
  PIN data_slave_w_ready
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1033.710 0.000 1033.990 4.000 ;
    END
  END data_slave_w_ready
  PIN data_slave_w_strb[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 540.640 4.000 541.240 ;
    END
  END data_slave_w_strb[0]
  PIN data_slave_w_strb[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 448.840 4.000 449.440 ;
    END
  END data_slave_w_strb[1]
  PIN data_slave_w_strb[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 788.990 1796.000 789.270 1800.000 ;
    END
  END data_slave_w_strb[2]
  PIN data_slave_w_strb[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1375.030 1796.000 1375.310 1800.000 ;
    END
  END data_slave_w_strb[3]
  PIN data_slave_w_strb[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1455.530 1796.000 1455.810 1800.000 ;
    END
  END data_slave_w_strb[4]
  PIN data_slave_w_strb[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 496.440 4.000 497.040 ;
    END
  END data_slave_w_strb[5]
  PIN data_slave_w_strb[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 625.640 1500.000 626.240 ;
    END
  END data_slave_w_strb[6]
  PIN data_slave_w_strb[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1264.840 4.000 1265.440 ;
    END
  END data_slave_w_strb[7]
  PIN data_slave_w_user[-1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 40.840 4.000 41.440 ;
    END
  END data_slave_w_user[-1]
  PIN data_slave_w_user[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1292.040 1500.000 1292.640 ;
    END
  END data_slave_w_user[0]
  PIN data_slave_w_valid
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 421.640 1500.000 422.240 ;
    END
  END data_slave_w_valid
  PIN dbg_master_ar_addr[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 10.240 1500.000 10.840 ;
    END
  END dbg_master_ar_addr[0]
  PIN dbg_master_ar_addr[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 959.650 0.000 959.930 4.000 ;
    END
  END dbg_master_ar_addr[10]
  PIN dbg_master_ar_addr[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 383.270 0.000 383.550 4.000 ;
    END
  END dbg_master_ar_addr[11]
  PIN dbg_master_ar_addr[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1071.040 1500.000 1071.640 ;
    END
  END dbg_master_ar_addr[12]
  PIN dbg_master_ar_addr[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1200.240 4.000 1200.840 ;
    END
  END dbg_master_ar_addr[13]
  PIN dbg_master_ar_addr[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 411.440 4.000 412.040 ;
    END
  END dbg_master_ar_addr[14]
  PIN dbg_master_ar_addr[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 608.640 1500.000 609.240 ;
    END
  END dbg_master_ar_addr[15]
  PIN dbg_master_ar_addr[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 523.640 1500.000 524.240 ;
    END
  END dbg_master_ar_addr[16]
  PIN dbg_master_ar_addr[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 673.070 1796.000 673.350 1800.000 ;
    END
  END dbg_master_ar_addr[17]
  PIN dbg_master_ar_addr[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1428.040 4.000 1428.640 ;
    END
  END dbg_master_ar_addr[18]
  PIN dbg_master_ar_addr[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.490 0.000 64.770 4.000 ;
    END
  END dbg_master_ar_addr[19]
  PIN dbg_master_ar_addr[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1230.840 4.000 1231.440 ;
    END
  END dbg_master_ar_addr[1]
  PIN dbg_master_ar_addr[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 112.790 0.000 113.070 4.000 ;
    END
  END dbg_master_ar_addr[20]
  PIN dbg_master_ar_addr[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1426.550 0.000 1426.830 4.000 ;
    END
  END dbg_master_ar_addr[21]
  PIN dbg_master_ar_addr[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 785.440 1500.000 786.040 ;
    END
  END dbg_master_ar_addr[22]
  PIN dbg_master_ar_addr[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 819.440 1500.000 820.040 ;
    END
  END dbg_master_ar_addr[23]
  PIN dbg_master_ar_addr[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 975.840 1500.000 976.440 ;
    END
  END dbg_master_ar_addr[24]
  PIN dbg_master_ar_addr[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 312.840 4.000 313.440 ;
    END
  END dbg_master_ar_addr[25]
  PIN dbg_master_ar_addr[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1428.040 1500.000 1428.640 ;
    END
  END dbg_master_ar_addr[26]
  PIN dbg_master_ar_addr[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 952.040 1500.000 952.640 ;
    END
  END dbg_master_ar_addr[27]
  PIN dbg_master_ar_addr[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 108.840 1500.000 109.440 ;
    END
  END dbg_master_ar_addr[28]
  PIN dbg_master_ar_addr[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1458.640 1500.000 1459.240 ;
    END
  END dbg_master_ar_addr[29]
  PIN dbg_master_ar_addr[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 890.840 4.000 891.440 ;
    END
  END dbg_master_ar_addr[2]
  PIN dbg_master_ar_addr[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1091.670 0.000 1091.950 4.000 ;
    END
  END dbg_master_ar_addr[30]
  PIN dbg_master_ar_addr[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 163.240 4.000 163.840 ;
    END
  END dbg_master_ar_addr[31]
  PIN dbg_master_ar_addr[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1413.670 1796.000 1413.950 1800.000 ;
    END
  END dbg_master_ar_addr[3]
  PIN dbg_master_ar_addr[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1230.840 1500.000 1231.440 ;
    END
  END dbg_master_ar_addr[4]
  PIN dbg_master_ar_addr[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.930 1796.000 71.210 1800.000 ;
    END
  END dbg_master_ar_addr[5]
  PIN dbg_master_ar_addr[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 958.840 1500.000 959.440 ;
    END
  END dbg_master_ar_addr[6]
  PIN dbg_master_ar_addr[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1567.440 1500.000 1568.040 ;
    END
  END dbg_master_ar_addr[7]
  PIN dbg_master_ar_addr[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 608.640 4.000 609.240 ;
    END
  END dbg_master_ar_addr[8]
  PIN dbg_master_ar_addr[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1033.710 1796.000 1033.990 1800.000 ;
    END
  END dbg_master_ar_addr[9]
  PIN dbg_master_ar_burst[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 173.440 4.000 174.040 ;
    END
  END dbg_master_ar_burst[0]
  PIN dbg_master_ar_burst[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1125.440 4.000 1126.040 ;
    END
  END dbg_master_ar_burst[1]
  PIN dbg_master_ar_cache[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 595.040 4.000 595.640 ;
    END
  END dbg_master_ar_cache[0]
  PIN dbg_master_ar_cache[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1094.890 0.000 1095.170 4.000 ;
    END
  END dbg_master_ar_cache[1]
  PIN dbg_master_ar_cache[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1246.230 1796.000 1246.510 1800.000 ;
    END
  END dbg_master_ar_cache[2]
  PIN dbg_master_ar_cache[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 747.130 0.000 747.410 4.000 ;
    END
  END dbg_master_ar_cache[3]
  PIN dbg_master_ar_id[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1439.430 0.000 1439.710 4.000 ;
    END
  END dbg_master_ar_id[0]
  PIN dbg_master_ar_id[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1686.440 4.000 1687.040 ;
    END
  END dbg_master_ar_id[1]
  PIN dbg_master_ar_id[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 669.840 4.000 670.440 ;
    END
  END dbg_master_ar_id[2]
  PIN dbg_master_ar_id[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1230.130 1796.000 1230.410 1800.000 ;
    END
  END dbg_master_ar_id[3]
  PIN dbg_master_ar_id[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 54.830 1796.000 55.110 1800.000 ;
    END
  END dbg_master_ar_id[4]
  PIN dbg_master_ar_id[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1275.040 4.000 1275.640 ;
    END
  END dbg_master_ar_id[5]
  PIN dbg_master_ar_id[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1026.840 4.000 1027.440 ;
    END
  END dbg_master_ar_id[6]
  PIN dbg_master_ar_id[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 533.840 4.000 534.440 ;
    END
  END dbg_master_ar_id[7]
  PIN dbg_master_ar_id[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1441.640 1500.000 1442.240 ;
    END
  END dbg_master_ar_id[8]
  PIN dbg_master_ar_id[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 721.370 0.000 721.650 4.000 ;
    END
  END dbg_master_ar_id[9]
  PIN dbg_master_ar_len[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 289.890 1796.000 290.170 1800.000 ;
    END
  END dbg_master_ar_len[0]
  PIN dbg_master_ar_len[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1227.440 4.000 1228.040 ;
    END
  END dbg_master_ar_len[1]
  PIN dbg_master_ar_len[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1101.640 4.000 1102.240 ;
    END
  END dbg_master_ar_len[2]
  PIN dbg_master_ar_len[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1059.470 0.000 1059.750 4.000 ;
    END
  END dbg_master_ar_len[3]
  PIN dbg_master_ar_len[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1268.770 0.000 1269.050 4.000 ;
    END
  END dbg_master_ar_len[4]
  PIN dbg_master_ar_len[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 282.240 1500.000 282.840 ;
    END
  END dbg_master_ar_len[5]
  PIN dbg_master_ar_len[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 512.070 0.000 512.350 4.000 ;
    END
  END dbg_master_ar_len[6]
  PIN dbg_master_ar_len[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1496.040 4.000 1496.640 ;
    END
  END dbg_master_ar_len[7]
  PIN dbg_master_ar_lock
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1196.840 4.000 1197.440 ;
    END
  END dbg_master_ar_lock
  PIN dbg_master_ar_prot[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 921.010 0.000 921.290 4.000 ;
    END
  END dbg_master_ar_prot[0]
  PIN dbg_master_ar_prot[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 221.040 1500.000 221.640 ;
    END
  END dbg_master_ar_prot[1]
  PIN dbg_master_ar_prot[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 293.110 0.000 293.390 4.000 ;
    END
  END dbg_master_ar_prot[2]
  PIN dbg_master_ar_qos[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1259.110 0.000 1259.390 4.000 ;
    END
  END dbg_master_ar_qos[0]
  PIN dbg_master_ar_qos[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1300.970 1796.000 1301.250 1800.000 ;
    END
  END dbg_master_ar_qos[1]
  PIN dbg_master_ar_qos[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1023.440 1500.000 1024.040 ;
    END
  END dbg_master_ar_qos[2]
  PIN dbg_master_ar_qos[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 157.870 0.000 158.150 4.000 ;
    END
  END dbg_master_ar_qos[3]
  PIN dbg_master_ar_ready
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1536.840 4.000 1537.440 ;
    END
  END dbg_master_ar_ready
  PIN dbg_master_ar_region[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 863.640 4.000 864.240 ;
    END
  END dbg_master_ar_region[0]
  PIN dbg_master_ar_region[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1645.640 4.000 1646.240 ;
    END
  END dbg_master_ar_region[1]
  PIN dbg_master_ar_region[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 702.050 1796.000 702.330 1800.000 ;
    END
  END dbg_master_ar_region[2]
  PIN dbg_master_ar_region[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 454.110 1796.000 454.390 1800.000 ;
    END
  END dbg_master_ar_region[3]
  PIN dbg_master_ar_size[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 711.710 1796.000 711.990 1800.000 ;
    END
  END dbg_master_ar_size[0]
  PIN dbg_master_ar_size[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 283.450 1796.000 283.730 1800.000 ;
    END
  END dbg_master_ar_size[1]
  PIN dbg_master_ar_size[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1666.040 1500.000 1666.640 ;
    END
  END dbg_master_ar_size[2]
  PIN dbg_master_ar_user[-1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 592.570 1796.000 592.850 1800.000 ;
    END
  END dbg_master_ar_user[-1]
  PIN dbg_master_ar_user[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 125.670 1796.000 125.950 1800.000 ;
    END
  END dbg_master_ar_user[0]
  PIN dbg_master_ar_valid
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 278.840 1500.000 279.440 ;
    END
  END dbg_master_ar_valid
  PIN dbg_master_aw_addr[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1380.440 1500.000 1381.040 ;
    END
  END dbg_master_aw_addr[0]
  PIN dbg_master_aw_addr[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 57.840 4.000 58.440 ;
    END
  END dbg_master_aw_addr[10]
  PIN dbg_master_aw_addr[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 520.240 4.000 520.840 ;
    END
  END dbg_master_aw_addr[11]
  PIN dbg_master_aw_addr[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 496.440 1500.000 497.040 ;
    END
  END dbg_master_aw_addr[12]
  PIN dbg_master_aw_addr[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 921.010 1796.000 921.290 1800.000 ;
    END
  END dbg_master_aw_addr[13]
  PIN dbg_master_aw_addr[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1458.750 1796.000 1459.030 1800.000 ;
    END
  END dbg_master_aw_addr[14]
  PIN dbg_master_aw_addr[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 763.230 1796.000 763.510 1800.000 ;
    END
  END dbg_master_aw_addr[15]
  PIN dbg_master_aw_addr[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 19.410 1796.000 19.690 1800.000 ;
    END
  END dbg_master_aw_addr[16]
  PIN dbg_master_aw_addr[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 209.390 0.000 209.670 4.000 ;
    END
  END dbg_master_aw_addr[17]
  PIN dbg_master_aw_addr[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 214.240 4.000 214.840 ;
    END
  END dbg_master_aw_addr[18]
  PIN dbg_master_aw_addr[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 513.440 1500.000 514.040 ;
    END
  END dbg_master_aw_addr[19]
  PIN dbg_master_aw_addr[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 88.440 1500.000 89.040 ;
    END
  END dbg_master_aw_addr[1]
  PIN dbg_master_aw_addr[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 724.590 0.000 724.870 4.000 ;
    END
  END dbg_master_aw_addr[20]
  PIN dbg_master_aw_addr[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1322.640 4.000 1323.240 ;
    END
  END dbg_master_aw_addr[21]
  PIN dbg_master_aw_addr[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1203.640 1500.000 1204.240 ;
    END
  END dbg_master_aw_addr[22]
  PIN dbg_master_aw_addr[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1336.390 1796.000 1336.670 1800.000 ;
    END
  END dbg_master_aw_addr[23]
  PIN dbg_master_aw_addr[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1118.640 4.000 1119.240 ;
    END
  END dbg_master_aw_addr[24]
  PIN dbg_master_aw_addr[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 476.650 1796.000 476.930 1800.000 ;
    END
  END dbg_master_aw_addr[25]
  PIN dbg_master_aw_addr[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1475.640 1500.000 1476.240 ;
    END
  END dbg_master_aw_addr[26]
  PIN dbg_master_aw_addr[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 367.240 4.000 367.840 ;
    END
  END dbg_master_aw_addr[27]
  PIN dbg_master_aw_addr[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 965.640 4.000 966.240 ;
    END
  END dbg_master_aw_addr[28]
  PIN dbg_master_aw_addr[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 122.450 0.000 122.730 4.000 ;
    END
  END dbg_master_aw_addr[29]
  PIN dbg_master_aw_addr[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1442.650 1796.000 1442.930 1800.000 ;
    END
  END dbg_master_aw_addr[2]
  PIN dbg_master_aw_addr[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 683.440 4.000 684.040 ;
    END
  END dbg_master_aw_addr[30]
  PIN dbg_master_aw_addr[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1536.840 1500.000 1537.440 ;
    END
  END dbg_master_aw_addr[31]
  PIN dbg_master_aw_addr[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1601.440 1500.000 1602.040 ;
    END
  END dbg_master_aw_addr[3]
  PIN dbg_master_aw_addr[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 986.040 4.000 986.640 ;
    END
  END dbg_master_aw_addr[4]
  PIN dbg_master_aw_addr[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1744.240 1500.000 1744.840 ;
    END
  END dbg_master_aw_addr[5]
  PIN dbg_master_aw_addr[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1275.210 0.000 1275.490 4.000 ;
    END
  END dbg_master_aw_addr[6]
  PIN dbg_master_aw_addr[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 653.750 0.000 654.030 4.000 ;
    END
  END dbg_master_aw_addr[7]
  PIN dbg_master_aw_addr[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 47.640 1500.000 48.240 ;
    END
  END dbg_master_aw_addr[8]
  PIN dbg_master_aw_addr[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1108.440 1500.000 1109.040 ;
    END
  END dbg_master_aw_addr[9]
  PIN dbg_master_aw_burst[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 241.590 0.000 241.870 4.000 ;
    END
  END dbg_master_aw_burst[0]
  PIN dbg_master_aw_burst[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 840.510 0.000 840.790 4.000 ;
    END
  END dbg_master_aw_burst[1]
  PIN dbg_master_aw_cache[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 750.350 1796.000 750.630 1800.000 ;
    END
  END dbg_master_aw_cache[0]
  PIN dbg_master_aw_cache[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 180.240 4.000 180.840 ;
    END
  END dbg_master_aw_cache[1]
  PIN dbg_master_aw_cache[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1197.930 1796.000 1198.210 1800.000 ;
    END
  END dbg_master_aw_cache[2]
  PIN dbg_master_aw_cache[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1417.840 1500.000 1418.440 ;
    END
  END dbg_master_aw_cache[3]
  PIN dbg_master_aw_id[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1761.240 1500.000 1761.840 ;
    END
  END dbg_master_aw_id[0]
  PIN dbg_master_aw_id[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1533.440 4.000 1534.040 ;
    END
  END dbg_master_aw_id[1]
  PIN dbg_master_aw_id[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1445.040 4.000 1445.640 ;
    END
  END dbg_master_aw_id[2]
  PIN dbg_master_aw_id[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1243.010 1796.000 1243.290 1800.000 ;
    END
  END dbg_master_aw_id[3]
  PIN dbg_master_aw_id[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 534.610 1796.000 534.890 1800.000 ;
    END
  END dbg_master_aw_id[4]
  PIN dbg_master_aw_id[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1241.040 4.000 1241.640 ;
    END
  END dbg_master_aw_id[5]
  PIN dbg_master_aw_id[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1006.440 1500.000 1007.040 ;
    END
  END dbg_master_aw_id[6]
  PIN dbg_master_aw_id[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 347.850 0.000 348.130 4.000 ;
    END
  END dbg_master_aw_id[7]
  PIN dbg_master_aw_id[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1788.440 4.000 1789.040 ;
    END
  END dbg_master_aw_id[8]
  PIN dbg_master_aw_id[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 384.240 4.000 384.840 ;
    END
  END dbg_master_aw_id[9]
  PIN dbg_master_aw_len[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 819.440 4.000 820.040 ;
    END
  END dbg_master_aw_len[0]
  PIN dbg_master_aw_len[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 582.910 1796.000 583.190 1800.000 ;
    END
  END dbg_master_aw_len[1]
  PIN dbg_master_aw_len[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 227.840 1500.000 228.440 ;
    END
  END dbg_master_aw_len[2]
  PIN dbg_master_aw_len[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1407.230 0.000 1407.510 4.000 ;
    END
  END dbg_master_aw_len[3]
  PIN dbg_master_aw_len[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1075.570 1796.000 1075.850 1800.000 ;
    END
  END dbg_master_aw_len[4]
  PIN dbg_master_aw_len[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1323.510 1796.000 1323.790 1800.000 ;
    END
  END dbg_master_aw_len[5]
  PIN dbg_master_aw_len[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 186.850 1796.000 187.130 1800.000 ;
    END
  END dbg_master_aw_len[6]
  PIN dbg_master_aw_len[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1455.240 4.000 1455.840 ;
    END
  END dbg_master_aw_len[7]
  PIN dbg_master_aw_lock
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1317.070 1796.000 1317.350 1800.000 ;
    END
  END dbg_master_aw_lock
  PIN dbg_master_aw_prot[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 331.750 0.000 332.030 4.000 ;
    END
  END dbg_master_aw_prot[0]
  PIN dbg_master_aw_prot[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 998.290 0.000 998.570 4.000 ;
    END
  END dbg_master_aw_prot[1]
  PIN dbg_master_aw_prot[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1326.040 1500.000 1326.640 ;
    END
  END dbg_master_aw_prot[2]
  PIN dbg_master_aw_qos[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 753.570 0.000 753.850 4.000 ;
    END
  END dbg_master_aw_qos[0]
  PIN dbg_master_aw_qos[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1288.090 0.000 1288.370 4.000 ;
    END
  END dbg_master_aw_qos[1]
  PIN dbg_master_aw_qos[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 966.090 1796.000 966.370 1800.000 ;
    END
  END dbg_master_aw_qos[2]
  PIN dbg_master_aw_qos[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 217.640 1500.000 218.240 ;
    END
  END dbg_master_aw_qos[3]
  PIN dbg_master_aw_ready
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1662.640 1500.000 1663.240 ;
    END
  END dbg_master_aw_ready
  PIN dbg_master_aw_region[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 343.440 4.000 344.040 ;
    END
  END dbg_master_aw_region[0]
  PIN dbg_master_aw_region[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1173.040 4.000 1173.640 ;
    END
  END dbg_master_aw_region[1]
  PIN dbg_master_aw_region[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1734.040 1500.000 1734.640 ;
    END
  END dbg_master_aw_region[2]
  PIN dbg_master_aw_region[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1081.240 4.000 1081.840 ;
    END
  END dbg_master_aw_region[3]
  PIN dbg_master_aw_size[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1156.070 0.000 1156.350 4.000 ;
    END
  END dbg_master_aw_size[0]
  PIN dbg_master_aw_size[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1078.790 0.000 1079.070 4.000 ;
    END
  END dbg_master_aw_size[1]
  PIN dbg_master_aw_size[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.390 1796.000 48.670 1800.000 ;
    END
  END dbg_master_aw_size[2]
  PIN dbg_master_aw_user[-1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1176.440 4.000 1177.040 ;
    END
  END dbg_master_aw_user[-1]
  PIN dbg_master_aw_user[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 605.450 1796.000 605.730 1800.000 ;
    END
  END dbg_master_aw_user[0]
  PIN dbg_master_aw_valid
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1383.840 1500.000 1384.440 ;
    END
  END dbg_master_aw_valid
  PIN dbg_master_b_id[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1516.440 1500.000 1517.040 ;
    END
  END dbg_master_b_id[0]
  PIN dbg_master_b_id[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 689.170 1796.000 689.450 1800.000 ;
    END
  END dbg_master_b_id[1]
  PIN dbg_master_b_id[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1081.240 1500.000 1081.840 ;
    END
  END dbg_master_b_id[2]
  PIN dbg_master_b_id[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 344.630 1796.000 344.910 1800.000 ;
    END
  END dbg_master_b_id[3]
  PIN dbg_master_b_id[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 265.240 4.000 265.840 ;
    END
  END dbg_master_b_id[4]
  PIN dbg_master_b_id[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 309.440 4.000 310.040 ;
    END
  END dbg_master_b_id[5]
  PIN dbg_master_b_id[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 561.040 4.000 561.640 ;
    END
  END dbg_master_b_id[6]
  PIN dbg_master_b_id[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1618.440 4.000 1619.040 ;
    END
  END dbg_master_b_id[7]
  PIN dbg_master_b_id[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1441.640 4.000 1442.240 ;
    END
  END dbg_master_b_id[8]
  PIN dbg_master_b_id[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 727.810 0.000 728.090 4.000 ;
    END
  END dbg_master_b_id[9]
  PIN dbg_master_b_ready
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 795.430 1796.000 795.710 1800.000 ;
    END
  END dbg_master_b_ready
  PIN dbg_master_b_resp[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 933.890 1796.000 934.170 1800.000 ;
    END
  END dbg_master_b_resp[0]
  PIN dbg_master_b_resp[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 450.890 1796.000 451.170 1800.000 ;
    END
  END dbg_master_b_resp[1]
  PIN dbg_master_b_user[-1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 460.550 0.000 460.830 4.000 ;
    END
  END dbg_master_b_user[-1]
  PIN dbg_master_b_user[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1764.640 1500.000 1765.240 ;
    END
  END dbg_master_b_user[0]
  PIN dbg_master_b_valid
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 748.040 4.000 748.640 ;
    END
  END dbg_master_b_valid
  PIN dbg_master_r_data[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1265.550 1796.000 1265.830 1800.000 ;
    END
  END dbg_master_r_data[0]
  PIN dbg_master_r_data[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1252.670 0.000 1252.950 4.000 ;
    END
  END dbg_master_r_data[10]
  PIN dbg_master_r_data[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 751.440 4.000 752.040 ;
    END
  END dbg_master_r_data[11]
  PIN dbg_master_r_data[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 702.050 0.000 702.330 4.000 ;
    END
  END dbg_master_r_data[12]
  PIN dbg_master_r_data[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 761.640 1500.000 762.240 ;
    END
  END dbg_master_r_data[13]
  PIN dbg_master_r_data[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1352.490 0.000 1352.770 4.000 ;
    END
  END dbg_master_r_data[14]
  PIN dbg_master_r_data[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 930.670 1796.000 930.950 1800.000 ;
    END
  END dbg_master_r_data[15]
  PIN dbg_master_r_data[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1156.040 4.000 1156.640 ;
    END
  END dbg_master_r_data[16]
  PIN dbg_master_r_data[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 608.670 1796.000 608.950 1800.000 ;
    END
  END dbg_master_r_data[17]
  PIN dbg_master_r_data[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1336.240 1500.000 1336.840 ;
    END
  END dbg_master_r_data[18]
  PIN dbg_master_r_data[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 499.840 1500.000 500.440 ;
    END
  END dbg_master_r_data[19]
  PIN dbg_master_r_data[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1557.240 4.000 1557.840 ;
    END
  END dbg_master_r_data[1]
  PIN dbg_master_r_data[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 293.110 1796.000 293.390 1800.000 ;
    END
  END dbg_master_r_data[20]
  PIN dbg_master_r_data[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 744.640 1500.000 745.240 ;
    END
  END dbg_master_r_data[21]
  PIN dbg_master_r_data[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 457.330 0.000 457.610 4.000 ;
    END
  END dbg_master_r_data[22]
  PIN dbg_master_r_data[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1550.440 4.000 1551.040 ;
    END
  END dbg_master_r_data[23]
  PIN dbg_master_r_data[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 357.040 4.000 357.640 ;
    END
  END dbg_master_r_data[24]
  PIN dbg_master_r_data[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1023.440 4.000 1024.040 ;
    END
  END dbg_master_r_data[25]
  PIN dbg_master_r_data[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 945.240 4.000 945.840 ;
    END
  END dbg_master_r_data[26]
  PIN dbg_master_r_data[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 275.440 1500.000 276.040 ;
    END
  END dbg_master_r_data[27]
  PIN dbg_master_r_data[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 812.640 4.000 813.240 ;
    END
  END dbg_master_r_data[28]
  PIN dbg_master_r_data[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 931.640 1500.000 932.240 ;
    END
  END dbg_master_r_data[29]
  PIN dbg_master_r_data[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 116.010 1796.000 116.290 1800.000 ;
    END
  END dbg_master_r_data[2]
  PIN dbg_master_r_data[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1320.290 1796.000 1320.570 1800.000 ;
    END
  END dbg_master_r_data[30]
  PIN dbg_master_r_data[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.290 1796.000 32.570 1800.000 ;
    END
  END dbg_master_r_data[31]
  PIN dbg_master_r_data[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1326.730 1796.000 1327.010 1800.000 ;
    END
  END dbg_master_r_data[32]
  PIN dbg_master_r_data[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 740.690 1796.000 740.970 1800.000 ;
    END
  END dbg_master_r_data[33]
  PIN dbg_master_r_data[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1768.040 1500.000 1768.640 ;
    END
  END dbg_master_r_data[34]
  PIN dbg_master_r_data[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 482.840 4.000 483.440 ;
    END
  END dbg_master_r_data[35]
  PIN dbg_master_r_data[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1310.630 1796.000 1310.910 1800.000 ;
    END
  END dbg_master_r_data[36]
  PIN dbg_master_r_data[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 296.330 0.000 296.610 4.000 ;
    END
  END dbg_master_r_data[37]
  PIN dbg_master_r_data[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1049.810 1796.000 1050.090 1800.000 ;
    END
  END dbg_master_r_data[38]
  PIN dbg_master_r_data[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 370.390 1796.000 370.670 1800.000 ;
    END
  END dbg_master_r_data[39]
  PIN dbg_master_r_data[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1201.150 1796.000 1201.430 1800.000 ;
    END
  END dbg_master_r_data[3]
  PIN dbg_master_r_data[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1159.440 1500.000 1160.040 ;
    END
  END dbg_master_r_data[40]
  PIN dbg_master_r_data[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1224.040 4.000 1224.640 ;
    END
  END dbg_master_r_data[41]
  PIN dbg_master_r_data[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1030.240 1500.000 1030.840 ;
    END
  END dbg_master_r_data[42]
  PIN dbg_master_r_data[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1798.640 4.000 1799.240 ;
    END
  END dbg_master_r_data[43]
  PIN dbg_master_r_data[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 758.240 1500.000 758.840 ;
    END
  END dbg_master_r_data[44]
  PIN dbg_master_r_data[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1281.650 1796.000 1281.930 1800.000 ;
    END
  END dbg_master_r_data[45]
  PIN dbg_master_r_data[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1085.230 0.000 1085.510 4.000 ;
    END
  END dbg_master_r_data[46]
  PIN dbg_master_r_data[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 425.130 1796.000 425.410 1800.000 ;
    END
  END dbg_master_r_data[47]
  PIN dbg_master_r_data[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 969.310 0.000 969.590 4.000 ;
    END
  END dbg_master_r_data[48]
  PIN dbg_master_r_data[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 299.550 0.000 299.830 4.000 ;
    END
  END dbg_master_r_data[49]
  PIN dbg_master_r_data[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1487.730 0.000 1488.010 4.000 ;
    END
  END dbg_master_r_data[4]
  PIN dbg_master_r_data[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 273.790 0.000 274.070 4.000 ;
    END
  END dbg_master_r_data[50]
  PIN dbg_master_r_data[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 635.840 1500.000 636.440 ;
    END
  END dbg_master_r_data[51]
  PIN dbg_master_r_data[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 9.750 1796.000 10.030 1800.000 ;
    END
  END dbg_master_r_data[52]
  PIN dbg_master_r_data[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 129.240 4.000 129.840 ;
    END
  END dbg_master_r_data[53]
  PIN dbg_master_r_data[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 115.640 1500.000 116.240 ;
    END
  END dbg_master_r_data[54]
  PIN dbg_master_r_data[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 809.240 4.000 809.840 ;
    END
  END dbg_master_r_data[55]
  PIN dbg_master_r_data[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 805.840 1500.000 806.440 ;
    END
  END dbg_master_r_data[56]
  PIN dbg_master_r_data[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1778.240 1500.000 1778.840 ;
    END
  END dbg_master_r_data[57]
  PIN dbg_master_r_data[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 734.440 4.000 735.040 ;
    END
  END dbg_master_r_data[58]
  PIN dbg_master_r_data[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.950 1796.000 42.230 1800.000 ;
    END
  END dbg_master_r_data[59]
  PIN dbg_master_r_data[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1191.490 0.000 1191.770 4.000 ;
    END
  END dbg_master_r_data[5]
  PIN dbg_master_r_data[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 360.730 1796.000 361.010 1800.000 ;
    END
  END dbg_master_r_data[60]
  PIN dbg_master_r_data[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1431.440 1500.000 1432.040 ;
    END
  END dbg_master_r_data[61]
  PIN dbg_master_r_data[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1642.240 1500.000 1642.840 ;
    END
  END dbg_master_r_data[62]
  PIN dbg_master_r_data[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1795.240 4.000 1795.840 ;
    END
  END dbg_master_r_data[63]
  PIN dbg_master_r_data[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.290 0.000 32.570 4.000 ;
    END
  END dbg_master_r_data[6]
  PIN dbg_master_r_data[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 816.040 4.000 816.640 ;
    END
  END dbg_master_r_data[7]
  PIN dbg_master_r_data[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1317.070 0.000 1317.350 4.000 ;
    END
  END dbg_master_r_data[8]
  PIN dbg_master_r_data[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 338.190 0.000 338.470 4.000 ;
    END
  END dbg_master_r_data[9]
  PIN dbg_master_r_id[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 761.640 4.000 762.240 ;
    END
  END dbg_master_r_id[0]
  PIN dbg_master_r_id[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1114.210 1796.000 1114.490 1800.000 ;
    END
  END dbg_master_r_id[1]
  PIN dbg_master_r_id[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1088.450 0.000 1088.730 4.000 ;
    END
  END dbg_master_r_id[2]
  PIN dbg_master_r_id[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1326.730 0.000 1327.010 4.000 ;
    END
  END dbg_master_r_id[3]
  PIN dbg_master_r_id[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1390.640 1500.000 1391.240 ;
    END
  END dbg_master_r_id[4]
  PIN dbg_master_r_id[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 204.040 1500.000 204.640 ;
    END
  END dbg_master_r_id[5]
  PIN dbg_master_r_id[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 564.440 4.000 565.040 ;
    END
  END dbg_master_r_id[6]
  PIN dbg_master_r_id[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1047.240 4.000 1047.840 ;
    END
  END dbg_master_r_id[7]
  PIN dbg_master_r_id[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1683.040 1500.000 1683.640 ;
    END
  END dbg_master_r_id[8]
  PIN dbg_master_r_id[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 296.330 1796.000 296.610 1800.000 ;
    END
  END dbg_master_r_id[9]
  PIN dbg_master_r_last
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 351.070 0.000 351.350 4.000 ;
    END
  END dbg_master_r_last
  PIN dbg_master_r_ready
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 74.150 1796.000 74.430 1800.000 ;
    END
  END dbg_master_r_ready
  PIN dbg_master_r_resp[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1156.040 1500.000 1156.640 ;
    END
  END dbg_master_r_resp[0]
  PIN dbg_master_r_resp[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1105.040 1500.000 1105.640 ;
    END
  END dbg_master_r_resp[1]
  PIN dbg_master_r_user[-1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 917.790 1796.000 918.070 1800.000 ;
    END
  END dbg_master_r_user[-1]
  PIN dbg_master_r_user[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 894.240 1500.000 894.840 ;
    END
  END dbg_master_r_user[0]
  PIN dbg_master_r_valid
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1649.040 4.000 1649.640 ;
    END
  END dbg_master_r_valid
  PIN dbg_master_w_data[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 824.410 0.000 824.690 4.000 ;
    END
  END dbg_master_w_data[0]
  PIN dbg_master_w_data[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 758.240 4.000 758.840 ;
    END
  END dbg_master_w_data[10]
  PIN dbg_master_w_data[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 472.640 1500.000 473.240 ;
    END
  END dbg_master_w_data[11]
  PIN dbg_master_w_data[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1628.640 4.000 1629.240 ;
    END
  END dbg_master_w_data[12]
  PIN dbg_master_w_data[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 991.850 1796.000 992.130 1800.000 ;
    END
  END dbg_master_w_data[13]
  PIN dbg_master_w_data[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1181.830 0.000 1182.110 4.000 ;
    END
  END dbg_master_w_data[14]
  PIN dbg_master_w_data[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 547.440 1500.000 548.040 ;
    END
  END dbg_master_w_data[15]
  PIN dbg_master_w_data[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 397.840 4.000 398.440 ;
    END
  END dbg_master_w_data[16]
  PIN dbg_master_w_data[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 115.640 4.000 116.240 ;
    END
  END dbg_master_w_data[17]
  PIN dbg_master_w_data[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 469.240 4.000 469.840 ;
    END
  END dbg_master_w_data[18]
  PIN dbg_master_w_data[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 444.450 0.000 444.730 4.000 ;
    END
  END dbg_master_w_data[19]
  PIN dbg_master_w_data[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1442.650 0.000 1442.930 4.000 ;
    END
  END dbg_master_w_data[1]
  PIN dbg_master_w_data[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1122.040 1500.000 1122.640 ;
    END
  END dbg_master_w_data[20]
  PIN dbg_master_w_data[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 724.240 4.000 724.840 ;
    END
  END dbg_master_w_data[21]
  PIN dbg_master_w_data[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 998.290 1796.000 998.570 1800.000 ;
    END
  END dbg_master_w_data[22]
  PIN dbg_master_w_data[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 197.240 4.000 197.840 ;
    END
  END dbg_master_w_data[23]
  PIN dbg_master_w_data[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 527.040 1500.000 527.640 ;
    END
  END dbg_master_w_data[24]
  PIN dbg_master_w_data[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1207.040 1500.000 1207.640 ;
    END
  END dbg_master_w_data[25]
  PIN dbg_master_w_data[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 972.440 4.000 973.040 ;
    END
  END dbg_master_w_data[26]
  PIN dbg_master_w_data[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 753.570 1796.000 753.850 1800.000 ;
    END
  END dbg_master_w_data[27]
  PIN dbg_master_w_data[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 459.040 1500.000 459.640 ;
    END
  END dbg_master_w_data[28]
  PIN dbg_master_w_data[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 27.240 4.000 27.840 ;
    END
  END dbg_master_w_data[29]
  PIN dbg_master_w_data[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1683.040 4.000 1683.640 ;
    END
  END dbg_master_w_data[2]
  PIN dbg_master_w_data[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1424.640 1500.000 1425.240 ;
    END
  END dbg_master_w_data[30]
  PIN dbg_master_w_data[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1484.510 0.000 1484.790 4.000 ;
    END
  END dbg_master_w_data[31]
  PIN dbg_master_w_data[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 299.240 4.000 299.840 ;
    END
  END dbg_master_w_data[32]
  PIN dbg_master_w_data[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 135.330 0.000 135.610 4.000 ;
    END
  END dbg_master_w_data[33]
  PIN dbg_master_w_data[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1713.640 1500.000 1714.240 ;
    END
  END dbg_master_w_data[34]
  PIN dbg_master_w_data[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1365.370 1796.000 1365.650 1800.000 ;
    END
  END dbg_master_w_data[35]
  PIN dbg_master_w_data[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 782.040 1500.000 782.640 ;
    END
  END dbg_master_w_data[36]
  PIN dbg_master_w_data[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1244.440 4.000 1245.040 ;
    END
  END dbg_master_w_data[37]
  PIN dbg_master_w_data[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 396.150 1796.000 396.430 1800.000 ;
    END
  END dbg_master_w_data[38]
  PIN dbg_master_w_data[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1072.350 1796.000 1072.630 1800.000 ;
    END
  END dbg_master_w_data[39]
  PIN dbg_master_w_data[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 418.690 0.000 418.970 4.000 ;
    END
  END dbg_master_w_data[3]
  PIN dbg_master_w_data[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 598.440 4.000 599.040 ;
    END
  END dbg_master_w_data[40]
  PIN dbg_master_w_data[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1011.170 0.000 1011.450 4.000 ;
    END
  END dbg_master_w_data[41]
  PIN dbg_master_w_data[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1523.240 4.000 1523.840 ;
    END
  END dbg_master_w_data[42]
  PIN dbg_master_w_data[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1509.640 1500.000 1510.240 ;
    END
  END dbg_master_w_data[43]
  PIN dbg_master_w_data[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1226.910 0.000 1227.190 4.000 ;
    END
  END dbg_master_w_data[44]
  PIN dbg_master_w_data[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1346.440 4.000 1347.040 ;
    END
  END dbg_master_w_data[45]
  PIN dbg_master_w_data[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1009.840 1500.000 1010.440 ;
    END
  END dbg_master_w_data[46]
  PIN dbg_master_w_data[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1638.840 1500.000 1639.440 ;
    END
  END dbg_master_w_data[47]
  PIN dbg_master_w_data[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1391.130 0.000 1391.410 4.000 ;
    END
  END dbg_master_w_data[48]
  PIN dbg_master_w_data[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1771.440 4.000 1772.040 ;
    END
  END dbg_master_w_data[49]
  PIN dbg_master_w_data[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 414.840 4.000 415.440 ;
    END
  END dbg_master_w_data[4]
  PIN dbg_master_w_data[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 254.470 0.000 254.750 4.000 ;
    END
  END dbg_master_w_data[50]
  PIN dbg_master_w_data[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 261.840 4.000 262.440 ;
    END
  END dbg_master_w_data[51]
  PIN dbg_master_w_data[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1033.640 1500.000 1034.240 ;
    END
  END dbg_master_w_data[52]
  PIN dbg_master_w_data[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 544.270 1796.000 544.550 1800.000 ;
    END
  END dbg_master_w_data[53]
  PIN dbg_master_w_data[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 151.430 1796.000 151.710 1800.000 ;
    END
  END dbg_master_w_data[54]
  PIN dbg_master_w_data[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 771.840 4.000 772.440 ;
    END
  END dbg_master_w_data[55]
  PIN dbg_master_w_data[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 814.750 1796.000 815.030 1800.000 ;
    END
  END dbg_master_w_data[56]
  PIN dbg_master_w_data[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 199.730 1796.000 200.010 1800.000 ;
    END
  END dbg_master_w_data[57]
  PIN dbg_master_w_data[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 785.770 1796.000 786.050 1800.000 ;
    END
  END dbg_master_w_data[58]
  PIN dbg_master_w_data[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 822.840 4.000 823.440 ;
    END
  END dbg_master_w_data[59]
  PIN dbg_master_w_data[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 251.250 0.000 251.530 4.000 ;
    END
  END dbg_master_w_data[5]
  PIN dbg_master_w_data[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1001.510 0.000 1001.790 4.000 ;
    END
  END dbg_master_w_data[60]
  PIN dbg_master_w_data[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 718.150 0.000 718.430 4.000 ;
    END
  END dbg_master_w_data[61]
  PIN dbg_master_w_data[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 756.790 0.000 757.070 4.000 ;
    END
  END dbg_master_w_data[62]
  PIN dbg_master_w_data[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1371.810 1796.000 1372.090 1800.000 ;
    END
  END dbg_master_w_data[63]
  PIN dbg_master_w_data[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 3.440 4.000 4.040 ;
    END
  END dbg_master_w_data[6]
  PIN dbg_master_w_data[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1159.290 1796.000 1159.570 1800.000 ;
    END
  END dbg_master_w_data[7]
  PIN dbg_master_w_data[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1611.640 1500.000 1612.240 ;
    END
  END dbg_master_w_data[8]
  PIN dbg_master_w_data[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1423.330 0.000 1423.610 4.000 ;
    END
  END dbg_master_w_data[9]
  PIN dbg_master_w_last
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 856.840 1500.000 857.440 ;
    END
  END dbg_master_w_last
  PIN dbg_master_w_ready
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 676.640 4.000 677.240 ;
    END
  END dbg_master_w_ready
  PIN dbg_master_w_strb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1329.440 4.000 1330.040 ;
    END
  END dbg_master_w_strb[0]
  PIN dbg_master_w_strb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 550.840 1500.000 551.440 ;
    END
  END dbg_master_w_strb[1]
  PIN dbg_master_w_strb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 557.150 1796.000 557.430 1800.000 ;
    END
  END dbg_master_w_strb[2]
  PIN dbg_master_w_strb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1778.240 4.000 1778.840 ;
    END
  END dbg_master_w_strb[3]
  PIN dbg_master_w_strb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 473.430 0.000 473.710 4.000 ;
    END
  END dbg_master_w_strb[4]
  PIN dbg_master_w_strb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 945.240 1500.000 945.840 ;
    END
  END dbg_master_w_strb[5]
  PIN dbg_master_w_strb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 673.240 1500.000 673.840 ;
    END
  END dbg_master_w_strb[6]
  PIN dbg_master_w_strb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1445.870 0.000 1446.150 4.000 ;
    END
  END dbg_master_w_strb[7]
  PIN dbg_master_w_user[-1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 128.890 1796.000 129.170 1800.000 ;
    END
  END dbg_master_w_user[-1]
  PIN dbg_master_w_user[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 683.440 1500.000 684.040 ;
    END
  END dbg_master_w_user[0]
  PIN dbg_master_w_valid
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1581.040 1500.000 1581.640 ;
    END
  END dbg_master_w_valid
  PIN debug_addr[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 212.610 1796.000 212.890 1800.000 ;
    END
  END debug_addr[0]
  PIN debug_addr[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 892.030 1796.000 892.310 1800.000 ;
    END
  END debug_addr[10]
  PIN debug_addr[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 462.440 4.000 463.040 ;
    END
  END debug_addr[11]
  PIN debug_addr[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1445.870 1796.000 1446.150 1800.000 ;
    END
  END debug_addr[12]
  PIN debug_addr[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 88.440 4.000 89.040 ;
    END
  END debug_addr[13]
  PIN debug_addr[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1122.040 4.000 1122.640 ;
    END
  END debug_addr[14]
  PIN debug_addr[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 972.440 1500.000 973.040 ;
    END
  END debug_addr[1]
  PIN debug_addr[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 141.770 1796.000 142.050 1800.000 ;
    END
  END debug_addr[2]
  PIN debug_addr[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 264.130 0.000 264.410 4.000 ;
    END
  END debug_addr[3]
  PIN debug_addr[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 873.840 1500.000 874.440 ;
    END
  END debug_addr[4]
  PIN debug_addr[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 611.890 0.000 612.170 4.000 ;
    END
  END debug_addr[5]
  PIN debug_addr[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1475.640 4.000 1476.240 ;
    END
  END debug_addr[6]
  PIN debug_addr[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 547.440 4.000 548.040 ;
    END
  END debug_addr[7]
  PIN debug_addr[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 574.640 1500.000 575.240 ;
    END
  END debug_addr[8]
  PIN debug_addr[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1449.090 1796.000 1449.370 1800.000 ;
    END
  END debug_addr[9]
  PIN debug_gnt
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 425.040 1500.000 425.640 ;
    END
  END debug_gnt
  PIN debug_rdata[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1547.040 4.000 1547.640 ;
    END
  END debug_rdata[0]
  PIN debug_rdata[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1149.630 1796.000 1149.910 1800.000 ;
    END
  END debug_rdata[10]
  PIN debug_rdata[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 935.040 1500.000 935.640 ;
    END
  END debug_rdata[11]
  PIN debug_rdata[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 766.450 1796.000 766.730 1800.000 ;
    END
  END debug_rdata[12]
  PIN debug_rdata[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 264.130 1796.000 264.410 1800.000 ;
    END
  END debug_rdata[13]
  PIN debug_rdata[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 995.070 0.000 995.350 4.000 ;
    END
  END debug_rdata[14]
  PIN debug_rdata[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 170.750 0.000 171.030 4.000 ;
    END
  END debug_rdata[15]
  PIN debug_rdata[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 829.640 4.000 830.240 ;
    END
  END debug_rdata[16]
  PIN debug_rdata[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 986.040 1500.000 986.640 ;
    END
  END debug_rdata[17]
  PIN debug_rdata[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1059.470 1796.000 1059.750 1800.000 ;
    END
  END debug_rdata[18]
  PIN debug_rdata[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 911.240 1500.000 911.840 ;
    END
  END debug_rdata[19]
  PIN debug_rdata[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 180.410 0.000 180.690 4.000 ;
    END
  END debug_rdata[1]
  PIN debug_rdata[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 34.040 1500.000 34.640 ;
    END
  END debug_rdata[20]
  PIN debug_rdata[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1057.440 1500.000 1058.040 ;
    END
  END debug_rdata[21]
  PIN debug_rdata[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 180.240 1500.000 180.840 ;
    END
  END debug_rdata[22]
  PIN debug_rdata[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 306.040 1500.000 306.640 ;
    END
  END debug_rdata[23]
  PIN debug_rdata[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 666.630 0.000 666.910 4.000 ;
    END
  END debug_rdata[24]
  PIN debug_rdata[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 550.840 4.000 551.440 ;
    END
  END debug_rdata[25]
  PIN debug_rdata[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 350.240 1500.000 350.840 ;
    END
  END debug_rdata[26]
  PIN debug_rdata[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1717.040 1500.000 1717.640 ;
    END
  END debug_rdata[27]
  PIN debug_rdata[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 428.440 1500.000 429.040 ;
    END
  END debug_rdata[28]
  PIN debug_rdata[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1543.640 1500.000 1544.240 ;
    END
  END debug_rdata[29]
  PIN debug_rdata[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 376.830 0.000 377.110 4.000 ;
    END
  END debug_rdata[2]
  PIN debug_rdata[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.270 0.000 61.550 4.000 ;
    END
  END debug_rdata[30]
  PIN debug_rdata[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 309.210 1796.000 309.490 1800.000 ;
    END
  END debug_rdata[31]
  PIN debug_rdata[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 679.510 0.000 679.790 4.000 ;
    END
  END debug_rdata[3]
  PIN debug_rdata[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1312.440 1500.000 1313.040 ;
    END
  END debug_rdata[4]
  PIN debug_rdata[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 879.150 1796.000 879.430 1800.000 ;
    END
  END debug_rdata[5]
  PIN debug_rdata[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1362.150 1796.000 1362.430 1800.000 ;
    END
  END debug_rdata[6]
  PIN debug_rdata[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 173.970 1796.000 174.250 1800.000 ;
    END
  END debug_rdata[7]
  PIN debug_rdata[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 460.550 1796.000 460.830 1800.000 ;
    END
  END debug_rdata[8]
  PIN debug_rdata[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 652.840 4.000 653.440 ;
    END
  END debug_rdata[9]
  PIN debug_req
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 177.190 0.000 177.470 4.000 ;
    END
  END debug_req
  PIN debug_rvalid
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 360.730 0.000 361.010 4.000 ;
    END
  END debug_rvalid
  PIN debug_wdata[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 450.890 0.000 451.170 4.000 ;
    END
  END debug_wdata[0]
  PIN debug_wdata[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 737.840 4.000 738.440 ;
    END
  END debug_wdata[10]
  PIN debug_wdata[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 54.830 0.000 55.110 4.000 ;
    END
  END debug_wdata[11]
  PIN debug_wdata[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 470.210 0.000 470.490 4.000 ;
    END
  END debug_wdata[12]
  PIN debug_wdata[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1570.840 1500.000 1571.440 ;
    END
  END debug_wdata[13]
  PIN debug_wdata[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 914.640 4.000 915.240 ;
    END
  END debug_wdata[14]
  PIN debug_wdata[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 418.690 1796.000 418.970 1800.000 ;
    END
  END debug_wdata[15]
  PIN debug_wdata[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 778.640 1500.000 779.240 ;
    END
  END debug_wdata[16]
  PIN debug_wdata[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 982.190 0.000 982.470 4.000 ;
    END
  END debug_wdata[17]
  PIN debug_wdata[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 391.040 4.000 391.640 ;
    END
  END debug_wdata[18]
  PIN debug_wdata[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 506.640 4.000 507.240 ;
    END
  END debug_wdata[19]
  PIN debug_wdata[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1479.040 1500.000 1479.640 ;
    END
  END debug_wdata[1]
  PIN debug_wdata[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 765.040 4.000 765.640 ;
    END
  END debug_wdata[20]
  PIN debug_wdata[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 244.840 1500.000 245.440 ;
    END
  END debug_wdata[21]
  PIN debug_wdata[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 748.040 1500.000 748.640 ;
    END
  END debug_wdata[22]
  PIN debug_wdata[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1183.240 1500.000 1183.840 ;
    END
  END debug_wdata[23]
  PIN debug_wdata[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1526.640 1500.000 1527.240 ;
    END
  END debug_wdata[24]
  PIN debug_wdata[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 595.040 1500.000 595.640 ;
    END
  END debug_wdata[25]
  PIN debug_wdata[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 885.590 1796.000 885.870 1800.000 ;
    END
  END debug_wdata[26]
  PIN debug_wdata[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1111.840 1500.000 1112.440 ;
    END
  END debug_wdata[27]
  PIN debug_wdata[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1117.430 0.000 1117.710 4.000 ;
    END
  END debug_wdata[28]
  PIN debug_wdata[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 956.430 1796.000 956.710 1800.000 ;
    END
  END debug_wdata[29]
  PIN debug_wdata[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1479.040 4.000 1479.640 ;
    END
  END debug_wdata[2]
  PIN debug_wdata[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 731.030 0.000 731.310 4.000 ;
    END
  END debug_wdata[30]
  PIN debug_wdata[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1451.840 1500.000 1452.440 ;
    END
  END debug_wdata[31]
  PIN debug_wdata[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 373.610 0.000 373.890 4.000 ;
    END
  END debug_wdata[3]
  PIN debug_wdata[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 751.440 1500.000 752.040 ;
    END
  END debug_wdata[4]
  PIN debug_wdata[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 966.090 0.000 966.370 4.000 ;
    END
  END debug_wdata[5]
  PIN debug_wdata[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1007.950 0.000 1008.230 4.000 ;
    END
  END debug_wdata[6]
  PIN debug_wdata[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1366.840 4.000 1367.440 ;
    END
  END debug_wdata[7]
  PIN debug_wdata[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 631.210 0.000 631.490 4.000 ;
    END
  END debug_wdata[8]
  PIN debug_wdata[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1001.510 1796.000 1001.790 1800.000 ;
    END
  END debug_wdata[9]
  PIN debug_we
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 698.830 0.000 699.110 4.000 ;
    END
  END debug_we
  PIN fetch_enable_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 231.930 0.000 232.210 4.000 ;
    END
  END fetch_enable_i
  PIN instr_slave_ar_addr[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1305.640 4.000 1306.240 ;
    END
  END instr_slave_ar_addr[0]
  PIN instr_slave_ar_addr[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1366.840 1500.000 1367.440 ;
    END
  END instr_slave_ar_addr[10]
  PIN instr_slave_ar_addr[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1404.240 1500.000 1404.840 ;
    END
  END instr_slave_ar_addr[11]
  PIN instr_slave_ar_addr[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1754.440 4.000 1755.040 ;
    END
  END instr_slave_ar_addr[12]
  PIN instr_slave_ar_addr[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1297.750 1796.000 1298.030 1800.000 ;
    END
  END instr_slave_ar_addr[13]
  PIN instr_slave_ar_addr[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 325.310 0.000 325.590 4.000 ;
    END
  END instr_slave_ar_addr[14]
  PIN instr_slave_ar_addr[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 776.110 1796.000 776.390 1800.000 ;
    END
  END instr_slave_ar_addr[15]
  PIN instr_slave_ar_addr[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 750.350 0.000 750.630 4.000 ;
    END
  END instr_slave_ar_addr[16]
  PIN instr_slave_ar_addr[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 99.910 0.000 100.190 4.000 ;
    END
  END instr_slave_ar_addr[17]
  PIN instr_slave_ar_addr[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1024.050 0.000 1024.330 4.000 ;
    END
  END instr_slave_ar_addr[18]
  PIN instr_slave_ar_addr[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 318.870 0.000 319.150 4.000 ;
    END
  END instr_slave_ar_addr[19]
  PIN instr_slave_ar_addr[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1635.440 1500.000 1636.040 ;
    END
  END instr_slave_ar_addr[1]
  PIN instr_slave_ar_addr[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 316.240 1500.000 316.840 ;
    END
  END instr_slave_ar_addr[20]
  PIN instr_slave_ar_addr[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 295.840 1500.000 296.440 ;
    END
  END instr_slave_ar_addr[21]
  PIN instr_slave_ar_addr[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1110.990 0.000 1111.270 4.000 ;
    END
  END instr_slave_ar_addr[22]
  PIN instr_slave_ar_addr[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 146.240 1500.000 146.840 ;
    END
  END instr_slave_ar_addr[23]
  PIN instr_slave_ar_addr[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1601.440 4.000 1602.040 ;
    END
  END instr_slave_ar_addr[24]
  PIN instr_slave_ar_addr[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 164.310 0.000 164.590 4.000 ;
    END
  END instr_slave_ar_addr[25]
  PIN instr_slave_ar_addr[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1329.950 0.000 1330.230 4.000 ;
    END
  END instr_slave_ar_addr[26]
  PIN instr_slave_ar_addr[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1530.040 1500.000 1530.640 ;
    END
  END instr_slave_ar_addr[27]
  PIN instr_slave_ar_addr[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 669.840 1500.000 670.440 ;
    END
  END instr_slave_ar_addr[28]
  PIN instr_slave_ar_addr[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 692.390 1796.000 692.670 1800.000 ;
    END
  END instr_slave_ar_addr[29]
  PIN instr_slave_ar_addr[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 663.410 1796.000 663.690 1800.000 ;
    END
  END instr_slave_ar_addr[2]
  PIN instr_slave_ar_addr[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 649.440 4.000 650.040 ;
    END
  END instr_slave_ar_addr[30]
  PIN instr_slave_ar_addr[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1594.640 1500.000 1595.240 ;
    END
  END instr_slave_ar_addr[31]
  PIN instr_slave_ar_addr[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1424.640 4.000 1425.240 ;
    END
  END instr_slave_ar_addr[3]
  PIN instr_slave_ar_addr[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1210.440 1500.000 1211.040 ;
    END
  END instr_slave_ar_addr[4]
  PIN instr_slave_ar_addr[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1217.240 4.000 1217.840 ;
    END
  END instr_slave_ar_addr[5]
  PIN instr_slave_ar_addr[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 792.240 1500.000 792.840 ;
    END
  END instr_slave_ar_addr[6]
  PIN instr_slave_ar_addr[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 224.440 1500.000 225.040 ;
    END
  END instr_slave_ar_addr[7]
  PIN instr_slave_ar_addr[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 754.840 1500.000 755.440 ;
    END
  END instr_slave_ar_addr[8]
  PIN instr_slave_ar_addr[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 808.310 0.000 808.590 4.000 ;
    END
  END instr_slave_ar_addr[9]
  PIN instr_slave_ar_burst[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 215.830 0.000 216.110 4.000 ;
    END
  END instr_slave_ar_burst[0]
  PIN instr_slave_ar_burst[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1383.840 4.000 1384.440 ;
    END
  END instr_slave_ar_burst[1]
  PIN instr_slave_ar_cache[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1570.840 4.000 1571.440 ;
    END
  END instr_slave_ar_cache[0]
  PIN instr_slave_ar_cache[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 438.640 1500.000 439.240 ;
    END
  END instr_slave_ar_cache[1]
  PIN instr_slave_ar_cache[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1173.040 1500.000 1173.640 ;
    END
  END instr_slave_ar_cache[2]
  PIN instr_slave_ar_cache[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 653.750 1796.000 654.030 1800.000 ;
    END
  END instr_slave_ar_cache[3]
  PIN instr_slave_ar_id[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 68.040 4.000 68.640 ;
    END
  END instr_slave_ar_id[0]
  PIN instr_slave_ar_id[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1179.840 4.000 1180.440 ;
    END
  END instr_slave_ar_id[1]
  PIN instr_slave_ar_id[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1465.190 1796.000 1465.470 1800.000 ;
    END
  END instr_slave_ar_id[2]
  PIN instr_slave_ar_id[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 466.990 1796.000 467.270 1800.000 ;
    END
  END instr_slave_ar_id[3]
  PIN instr_slave_ar_id[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 741.240 1500.000 741.840 ;
    END
  END instr_slave_ar_id[4]
  PIN instr_slave_ar_id[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1375.030 0.000 1375.310 4.000 ;
    END
  END instr_slave_ar_id[5]
  PIN instr_slave_ar_id[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 534.610 0.000 534.890 4.000 ;
    END
  END instr_slave_ar_id[6]
  PIN instr_slave_ar_id[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 809.240 1500.000 809.840 ;
    END
  END instr_slave_ar_id[7]
  PIN instr_slave_ar_id[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1132.240 4.000 1132.840 ;
    END
  END instr_slave_ar_id[8]
  PIN instr_slave_ar_id[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 850.040 4.000 850.640 ;
    END
  END instr_slave_ar_id[9]
  PIN instr_slave_ar_len[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1339.640 4.000 1340.240 ;
    END
  END instr_slave_ar_len[0]
  PIN instr_slave_ar_len[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 161.090 0.000 161.370 4.000 ;
    END
  END instr_slave_ar_len[1]
  PIN instr_slave_ar_len[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 154.650 0.000 154.930 4.000 ;
    END
  END instr_slave_ar_len[2]
  PIN instr_slave_ar_len[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1062.690 0.000 1062.970 4.000 ;
    END
  END instr_slave_ar_len[3]
  PIN instr_slave_ar_len[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 125.670 0.000 125.950 4.000 ;
    END
  END instr_slave_ar_len[4]
  PIN instr_slave_ar_len[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1040.150 1796.000 1040.430 1800.000 ;
    END
  END instr_slave_ar_len[5]
  PIN instr_slave_ar_len[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1074.440 1500.000 1075.040 ;
    END
  END instr_slave_ar_len[6]
  PIN instr_slave_ar_len[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1706.840 4.000 1707.440 ;
    END
  END instr_slave_ar_len[7]
  PIN instr_slave_ar_lock
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1217.250 0.000 1217.530 4.000 ;
    END
  END instr_slave_ar_lock
  PIN instr_slave_ar_prot[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1254.640 4.000 1255.240 ;
    END
  END instr_slave_ar_prot[0]
  PIN instr_slave_ar_prot[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 867.040 1500.000 867.640 ;
    END
  END instr_slave_ar_prot[1]
  PIN instr_slave_ar_prot[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 660.190 0.000 660.470 4.000 ;
    END
  END instr_slave_ar_prot[2]
  PIN instr_slave_ar_qos[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1468.840 4.000 1469.440 ;
    END
  END instr_slave_ar_qos[0]
  PIN instr_slave_ar_qos[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1404.010 0.000 1404.290 4.000 ;
    END
  END instr_slave_ar_qos[1]
  PIN instr_slave_ar_qos[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 151.430 0.000 151.710 4.000 ;
    END
  END instr_slave_ar_qos[2]
  PIN instr_slave_ar_qos[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1462.040 1500.000 1462.640 ;
    END
  END instr_slave_ar_qos[3]
  PIN instr_slave_ar_ready
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1037.040 1500.000 1037.640 ;
    END
  END instr_slave_ar_ready
  PIN instr_slave_ar_region[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 404.640 1500.000 405.240 ;
    END
  END instr_slave_ar_region[0]
  PIN instr_slave_ar_region[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 399.370 0.000 399.650 4.000 ;
    END
  END instr_slave_ar_region[1]
  PIN instr_slave_ar_region[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 775.240 4.000 775.840 ;
    END
  END instr_slave_ar_region[2]
  PIN instr_slave_ar_region[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 867.040 4.000 867.640 ;
    END
  END instr_slave_ar_region[3]
  PIN instr_slave_ar_size[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 116.010 0.000 116.290 4.000 ;
    END
  END instr_slave_ar_size[0]
  PIN instr_slave_ar_size[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1455.530 0.000 1455.810 4.000 ;
    END
  END instr_slave_ar_size[1]
  PIN instr_slave_ar_size[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 869.490 1796.000 869.770 1800.000 ;
    END
  END instr_slave_ar_size[2]
  PIN instr_slave_ar_user[-1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1594.640 4.000 1595.240 ;
    END
  END instr_slave_ar_user[-1]
  PIN instr_slave_ar_user[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 219.050 0.000 219.330 4.000 ;
    END
  END instr_slave_ar_user[0]
  PIN instr_slave_ar_valid
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1255.890 1796.000 1256.170 1800.000 ;
    END
  END instr_slave_ar_valid
  PIN instr_slave_aw_addr[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 231.240 1500.000 231.840 ;
    END
  END instr_slave_aw_addr[0]
  PIN instr_slave_aw_addr[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1632.040 1500.000 1632.640 ;
    END
  END instr_slave_aw_addr[10]
  PIN instr_slave_aw_addr[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 302.770 0.000 303.050 4.000 ;
    END
  END instr_slave_aw_addr[11]
  PIN instr_slave_aw_addr[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1400.840 1500.000 1401.440 ;
    END
  END instr_slave_aw_addr[12]
  PIN instr_slave_aw_addr[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 843.730 0.000 844.010 4.000 ;
    END
  END instr_slave_aw_addr[13]
  PIN instr_slave_aw_addr[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 421.640 4.000 422.240 ;
    END
  END instr_slave_aw_addr[14]
  PIN instr_slave_aw_addr[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1305.640 1500.000 1306.240 ;
    END
  END instr_slave_aw_addr[15]
  PIN instr_slave_aw_addr[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 724.240 1500.000 724.840 ;
    END
  END instr_slave_aw_addr[16]
  PIN instr_slave_aw_addr[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1635.440 4.000 1636.040 ;
    END
  END instr_slave_aw_addr[17]
  PIN instr_slave_aw_addr[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 775.240 1500.000 775.840 ;
    END
  END instr_slave_aw_addr[18]
  PIN instr_slave_aw_addr[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 85.040 4.000 85.640 ;
    END
  END instr_slave_aw_addr[19]
  PIN instr_slave_aw_addr[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 705.270 1796.000 705.550 1800.000 ;
    END
  END instr_slave_aw_addr[1]
  PIN instr_slave_aw_addr[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1241.040 1500.000 1241.640 ;
    END
  END instr_slave_aw_addr[20]
  PIN instr_slave_aw_addr[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1094.840 4.000 1095.440 ;
    END
  END instr_slave_aw_addr[21]
  PIN instr_slave_aw_addr[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1120.650 0.000 1120.930 4.000 ;
    END
  END instr_slave_aw_addr[22]
  PIN instr_slave_aw_addr[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 574.640 4.000 575.240 ;
    END
  END instr_slave_aw_addr[23]
  PIN instr_slave_aw_addr[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 363.840 1500.000 364.440 ;
    END
  END instr_slave_aw_addr[24]
  PIN instr_slave_aw_addr[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1143.190 1796.000 1143.470 1800.000 ;
    END
  END instr_slave_aw_addr[25]
  PIN instr_slave_aw_addr[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 51.610 1796.000 51.890 1800.000 ;
    END
  END instr_slave_aw_addr[26]
  PIN instr_slave_aw_addr[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1294.530 0.000 1294.810 4.000 ;
    END
  END instr_slave_aw_addr[27]
  PIN instr_slave_aw_addr[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 989.440 1500.000 990.040 ;
    END
  END instr_slave_aw_addr[28]
  PIN instr_slave_aw_addr[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 91.840 1500.000 92.440 ;
    END
  END instr_slave_aw_addr[29]
  PIN instr_slave_aw_addr[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 209.390 1796.000 209.670 1800.000 ;
    END
  END instr_slave_aw_addr[2]
  PIN instr_slave_aw_addr[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1693.240 1500.000 1693.840 ;
    END
  END instr_slave_aw_addr[30]
  PIN instr_slave_aw_addr[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 969.040 4.000 969.640 ;
    END
  END instr_slave_aw_addr[31]
  PIN instr_slave_aw_addr[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1676.240 1500.000 1676.840 ;
    END
  END instr_slave_aw_addr[3]
  PIN instr_slave_aw_addr[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 940.330 1796.000 940.610 1800.000 ;
    END
  END instr_slave_aw_addr[4]
  PIN instr_slave_aw_addr[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 156.440 4.000 157.040 ;
    END
  END instr_slave_aw_addr[5]
  PIN instr_slave_aw_addr[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1429.770 0.000 1430.050 4.000 ;
    END
  END instr_slave_aw_addr[6]
  PIN instr_slave_aw_addr[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 801.870 1796.000 802.150 1800.000 ;
    END
  END instr_slave_aw_addr[7]
  PIN instr_slave_aw_addr[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1310.630 0.000 1310.910 4.000 ;
    END
  END instr_slave_aw_addr[8]
  PIN instr_slave_aw_addr[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 924.840 4.000 925.440 ;
    END
  END instr_slave_aw_addr[9]
  PIN instr_slave_aw_burst[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1343.040 4.000 1343.640 ;
    END
  END instr_slave_aw_burst[0]
  PIN instr_slave_aw_burst[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 624.770 0.000 625.050 4.000 ;
    END
  END instr_slave_aw_burst[1]
  PIN instr_slave_aw_cache[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 102.040 1500.000 102.640 ;
    END
  END instr_slave_aw_cache[0]
  PIN instr_slave_aw_cache[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1326.040 4.000 1326.640 ;
    END
  END instr_slave_aw_cache[1]
  PIN instr_slave_aw_cache[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1584.440 1500.000 1585.040 ;
    END
  END instr_slave_aw_cache[2]
  PIN instr_slave_aw_cache[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1322.640 1500.000 1323.240 ;
    END
  END instr_slave_aw_cache[3]
  PIN instr_slave_aw_id[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 933.890 0.000 934.170 4.000 ;
    END
  END instr_slave_aw_id[0]
  PIN instr_slave_aw_id[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 434.790 0.000 435.070 4.000 ;
    END
  END instr_slave_aw_id[1]
  PIN instr_slave_aw_id[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 312.430 0.000 312.710 4.000 ;
    END
  END instr_slave_aw_id[2]
  PIN instr_slave_aw_id[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1115.240 1500.000 1115.840 ;
    END
  END instr_slave_aw_id[3]
  PIN instr_slave_aw_id[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 524.950 1796.000 525.230 1800.000 ;
    END
  END instr_slave_aw_id[4]
  PIN instr_slave_aw_id[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 25.850 1796.000 26.130 1800.000 ;
    END
  END instr_slave_aw_id[5]
  PIN instr_slave_aw_id[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 904.910 1796.000 905.190 1800.000 ;
    END
  END instr_slave_aw_id[6]
  PIN instr_slave_aw_id[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 96.690 1796.000 96.970 1800.000 ;
    END
  END instr_slave_aw_id[7]
  PIN instr_slave_aw_id[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 292.440 1500.000 293.040 ;
    END
  END instr_slave_aw_id[8]
  PIN instr_slave_aw_id[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1064.240 1500.000 1064.840 ;
    END
  END instr_slave_aw_id[9]
  PIN instr_slave_aw_len[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1526.640 4.000 1527.240 ;
    END
  END instr_slave_aw_len[0]
  PIN instr_slave_aw_len[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 766.450 0.000 766.730 4.000 ;
    END
  END instr_slave_aw_len[1]
  PIN instr_slave_aw_len[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 731.040 1500.000 731.640 ;
    END
  END instr_slave_aw_len[2]
  PIN instr_slave_aw_len[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1436.210 0.000 1436.490 4.000 ;
    END
  END instr_slave_aw_len[3]
  PIN instr_slave_aw_len[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1214.030 0.000 1214.310 4.000 ;
    END
  END instr_slave_aw_len[4]
  PIN instr_slave_aw_len[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 843.730 1796.000 844.010 1800.000 ;
    END
  END instr_slave_aw_len[5]
  PIN instr_slave_aw_len[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 866.270 0.000 866.550 4.000 ;
    END
  END instr_slave_aw_len[6]
  PIN instr_slave_aw_len[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 962.240 4.000 962.840 ;
    END
  END instr_slave_aw_len[7]
  PIN instr_slave_aw_lock
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1384.690 0.000 1384.970 4.000 ;
    END
  END instr_slave_aw_lock
  PIN instr_slave_aw_prot[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 105.440 4.000 106.040 ;
    END
  END instr_slave_aw_prot[0]
  PIN instr_slave_aw_prot[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 341.410 0.000 341.690 4.000 ;
    END
  END instr_slave_aw_prot[1]
  PIN instr_slave_aw_prot[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 122.440 4.000 123.040 ;
    END
  END instr_slave_aw_prot[2]
  PIN instr_slave_aw_qos[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 235.150 1796.000 235.430 1800.000 ;
    END
  END instr_slave_aw_qos[0]
  PIN instr_slave_aw_qos[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 305.990 1796.000 306.270 1800.000 ;
    END
  END instr_slave_aw_qos[1]
  PIN instr_slave_aw_qos[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1176.440 1500.000 1177.040 ;
    END
  END instr_slave_aw_qos[2]
  PIN instr_slave_aw_qos[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 286.670 1796.000 286.950 1800.000 ;
    END
  END instr_slave_aw_qos[3]
  PIN instr_slave_aw_ready
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1084.640 1500.000 1085.240 ;
    END
  END instr_slave_aw_ready
  PIN instr_slave_aw_region[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 955.440 4.000 956.040 ;
    END
  END instr_slave_aw_region[0]
  PIN instr_slave_aw_region[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 13.640 1500.000 14.240 ;
    END
  END instr_slave_aw_region[1]
  PIN instr_slave_aw_region[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1404.240 4.000 1404.840 ;
    END
  END instr_slave_aw_region[2]
  PIN instr_slave_aw_region[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 328.530 1796.000 328.810 1800.000 ;
    END
  END instr_slave_aw_region[3]
  PIN instr_slave_aw_size[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.710 0.000 67.990 4.000 ;
    END
  END instr_slave_aw_size[0]
  PIN instr_slave_aw_size[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1268.770 1796.000 1269.050 1800.000 ;
    END
  END instr_slave_aw_size[1]
  PIN instr_slave_aw_size[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 214.240 1500.000 214.840 ;
    END
  END instr_slave_aw_size[2]
  PIN instr_slave_aw_user[-1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 634.430 1796.000 634.710 1800.000 ;
    END
  END instr_slave_aw_user[-1]
  PIN instr_slave_aw_user[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 486.310 1796.000 486.590 1800.000 ;
    END
  END instr_slave_aw_user[0]
  PIN instr_slave_aw_valid
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1284.870 0.000 1285.150 4.000 ;
    END
  END instr_slave_aw_valid
  PIN instr_slave_b_id[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1598.040 4.000 1598.640 ;
    END
  END instr_slave_b_id[0]
  PIN instr_slave_b_id[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 707.240 1500.000 707.840 ;
    END
  END instr_slave_b_id[1]
  PIN instr_slave_b_id[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 357.510 1796.000 357.790 1800.000 ;
    END
  END instr_slave_b_id[2]
  PIN instr_slave_b_id[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 99.910 1796.000 100.190 1800.000 ;
    END
  END instr_slave_b_id[3]
  PIN instr_slave_b_id[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 817.970 0.000 818.250 4.000 ;
    END
  END instr_slave_b_id[4]
  PIN instr_slave_b_id[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 199.730 0.000 200.010 4.000 ;
    END
  END instr_slave_b_id[5]
  PIN instr_slave_b_id[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1577.640 1500.000 1578.240 ;
    END
  END instr_slave_b_id[6]
  PIN instr_slave_b_id[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1136.750 1796.000 1137.030 1800.000 ;
    END
  END instr_slave_b_id[7]
  PIN instr_slave_b_id[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 109.570 0.000 109.850 4.000 ;
    END
  END instr_slave_b_id[8]
  PIN instr_slave_b_id[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1652.440 4.000 1653.040 ;
    END
  END instr_slave_b_id[9]
  PIN instr_slave_b_ready
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1482.440 4.000 1483.040 ;
    END
  END instr_slave_b_ready
  PIN instr_slave_b_resp[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 557.640 4.000 558.240 ;
    END
  END instr_slave_b_resp[0]
  PIN instr_slave_b_resp[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1339.610 1796.000 1339.890 1800.000 ;
    END
  END instr_slave_b_resp[1]
  PIN instr_slave_b_user[-1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1069.130 0.000 1069.410 4.000 ;
    END
  END instr_slave_b_user[-1]
  PIN instr_slave_b_user[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 911.350 0.000 911.630 4.000 ;
    END
  END instr_slave_b_user[0]
  PIN instr_slave_b_valid
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 666.630 1796.000 666.910 1800.000 ;
    END
  END instr_slave_b_valid
  PIN instr_slave_r_data[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 846.640 1500.000 847.240 ;
    END
  END instr_slave_r_data[0]
  PIN instr_slave_r_data[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1720.440 1500.000 1721.040 ;
    END
  END instr_slave_r_data[10]
  PIN instr_slave_r_data[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1264.840 1500.000 1265.440 ;
    END
  END instr_slave_r_data[11]
  PIN instr_slave_r_data[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 217.640 4.000 218.240 ;
    END
  END instr_slave_r_data[12]
  PIN instr_slave_r_data[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1207.040 4.000 1207.640 ;
    END
  END instr_slave_r_data[13]
  PIN instr_slave_r_data[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 894.240 4.000 894.840 ;
    END
  END instr_slave_r_data[14]
  PIN instr_slave_r_data[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 969.310 1796.000 969.590 1800.000 ;
    END
  END instr_slave_r_data[15]
  PIN instr_slave_r_data[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 571.240 1500.000 571.840 ;
    END
  END instr_slave_r_data[16]
  PIN instr_slave_r_data[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1553.840 1500.000 1554.440 ;
    END
  END instr_slave_r_data[17]
  PIN instr_slave_r_data[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 434.790 1796.000 435.070 1800.000 ;
    END
  END instr_slave_r_data[18]
  PIN instr_slave_r_data[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 241.440 4.000 242.040 ;
    END
  END instr_slave_r_data[19]
  PIN instr_slave_r_data[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 836.440 1500.000 837.040 ;
    END
  END instr_slave_r_data[1]
  PIN instr_slave_r_data[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 374.040 1500.000 374.640 ;
    END
  END instr_slave_r_data[20]
  PIN instr_slave_r_data[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 77.370 1796.000 77.650 1800.000 ;
    END
  END instr_slave_r_data[21]
  PIN instr_slave_r_data[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 103.130 1796.000 103.410 1800.000 ;
    END
  END instr_slave_r_data[22]
  PIN instr_slave_r_data[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1360.040 1500.000 1360.640 ;
    END
  END instr_slave_r_data[23]
  PIN instr_slave_r_data[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 119.040 4.000 119.640 ;
    END
  END instr_slave_r_data[24]
  PIN instr_slave_r_data[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1185.050 0.000 1185.330 4.000 ;
    END
  END instr_slave_r_data[25]
  PIN instr_slave_r_data[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 374.040 4.000 374.640 ;
    END
  END instr_slave_r_data[26]
  PIN instr_slave_r_data[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1604.840 1500.000 1605.440 ;
    END
  END instr_slave_r_data[27]
  PIN instr_slave_r_data[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 612.040 4.000 612.640 ;
    END
  END instr_slave_r_data[28]
  PIN instr_slave_r_data[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 969.040 1500.000 969.640 ;
    END
  END instr_slave_r_data[29]
  PIN instr_slave_r_data[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 441.230 0.000 441.510 4.000 ;
    END
  END instr_slave_r_data[2]
  PIN instr_slave_r_data[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1203.640 4.000 1204.240 ;
    END
  END instr_slave_r_data[30]
  PIN instr_slave_r_data[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1275.040 1500.000 1275.640 ;
    END
  END instr_slave_r_data[31]
  PIN instr_slave_r_data[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1468.410 0.000 1468.690 4.000 ;
    END
  END instr_slave_r_data[32]
  PIN instr_slave_r_data[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1730.640 1500.000 1731.240 ;
    END
  END instr_slave_r_data[33]
  PIN instr_slave_r_data[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1262.330 1796.000 1262.610 1800.000 ;
    END
  END instr_slave_r_data[34]
  PIN instr_slave_r_data[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 644.090 1796.000 644.370 1800.000 ;
    END
  END instr_slave_r_data[35]
  PIN instr_slave_r_data[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1146.410 1796.000 1146.690 1800.000 ;
    END
  END instr_slave_r_data[36]
  PIN instr_slave_r_data[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1696.640 1500.000 1697.240 ;
    END
  END instr_slave_r_data[37]
  PIN instr_slave_r_data[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 268.640 1500.000 269.240 ;
    END
  END instr_slave_r_data[38]
  PIN instr_slave_r_data[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1127.090 1796.000 1127.370 1800.000 ;
    END
  END instr_slave_r_data[39]
  PIN instr_slave_r_data[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 853.390 0.000 853.670 4.000 ;
    END
  END instr_slave_r_data[3]
  PIN instr_slave_r_data[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 64.640 1500.000 65.240 ;
    END
  END instr_slave_r_data[40]
  PIN instr_slave_r_data[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 921.440 1500.000 922.040 ;
    END
  END instr_slave_r_data[41]
  PIN instr_slave_r_data[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 785.440 4.000 786.040 ;
    END
  END instr_slave_r_data[42]
  PIN instr_slave_r_data[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 83.810 0.000 84.090 4.000 ;
    END
  END instr_slave_r_data[43]
  PIN instr_slave_r_data[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 792.240 4.000 792.840 ;
    END
  END instr_slave_r_data[44]
  PIN instr_slave_r_data[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 846.950 0.000 847.230 4.000 ;
    END
  END instr_slave_r_data[45]
  PIN instr_slave_r_data[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1082.010 0.000 1082.290 4.000 ;
    END
  END instr_slave_r_data[46]
  PIN instr_slave_r_data[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1054.040 4.000 1054.640 ;
    END
  END instr_slave_r_data[47]
  PIN instr_slave_r_data[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 278.840 4.000 279.440 ;
    END
  END instr_slave_r_data[48]
  PIN instr_slave_r_data[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 703.840 1500.000 704.440 ;
    END
  END instr_slave_r_data[49]
  PIN instr_slave_r_data[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1358.930 1796.000 1359.210 1800.000 ;
    END
  END instr_slave_r_data[4]
  PIN instr_slave_r_data[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 897.640 1500.000 898.240 ;
    END
  END instr_slave_r_data[50]
  PIN instr_slave_r_data[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1224.040 1500.000 1224.640 ;
    END
  END instr_slave_r_data[51]
  PIN instr_slave_r_data[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1478.070 0.000 1478.350 4.000 ;
    END
  END instr_slave_r_data[52]
  PIN instr_slave_r_data[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 779.330 0.000 779.610 4.000 ;
    END
  END instr_slave_r_data[53]
  PIN instr_slave_r_data[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1378.250 0.000 1378.530 4.000 ;
    END
  END instr_slave_r_data[54]
  PIN instr_slave_r_data[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 19.410 0.000 19.690 4.000 ;
    END
  END instr_slave_r_data[55]
  PIN instr_slave_r_data[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1764.640 4.000 1765.240 ;
    END
  END instr_slave_r_data[56]
  PIN instr_slave_r_data[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1471.630 1796.000 1471.910 1800.000 ;
    END
  END instr_slave_r_data[57]
  PIN instr_slave_r_data[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 122.450 1796.000 122.730 1800.000 ;
    END
  END instr_slave_r_data[58]
  PIN instr_slave_r_data[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 492.750 0.000 493.030 4.000 ;
    END
  END instr_slave_r_data[59]
  PIN instr_slave_r_data[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 329.840 1500.000 330.440 ;
    END
  END instr_slave_r_data[5]
  PIN instr_slave_r_data[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.950 0.000 42.230 4.000 ;
    END
  END instr_slave_r_data[60]
  PIN instr_slave_r_data[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1411.040 1500.000 1411.640 ;
    END
  END instr_slave_r_data[61]
  PIN instr_slave_r_data[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1550.440 1500.000 1551.040 ;
    END
  END instr_slave_r_data[62]
  PIN instr_slave_r_data[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1429.770 1796.000 1430.050 1800.000 ;
    END
  END instr_slave_r_data[63]
  PIN instr_slave_r_data[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 741.240 4.000 741.840 ;
    END
  END instr_slave_r_data[6]
  PIN instr_slave_r_data[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 856.610 1796.000 856.890 1800.000 ;
    END
  END instr_slave_r_data[7]
  PIN instr_slave_r_data[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 792.210 0.000 792.490 4.000 ;
    END
  END instr_slave_r_data[8]
  PIN instr_slave_r_data[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 112.790 1796.000 113.070 1800.000 ;
    END
  END instr_slave_r_data[9]
  PIN instr_slave_r_id[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 412.250 0.000 412.530 4.000 ;
    END
  END instr_slave_r_id[0]
  PIN instr_slave_r_id[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 521.730 1796.000 522.010 1800.000 ;
    END
  END instr_slave_r_id[1]
  PIN instr_slave_r_id[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1754.440 1500.000 1755.040 ;
    END
  END instr_slave_r_id[2]
  PIN instr_slave_r_id[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 331.750 1796.000 332.030 1800.000 ;
    END
  END instr_slave_r_id[3]
  PIN instr_slave_r_id[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 673.240 4.000 673.840 ;
    END
  END instr_slave_r_id[4]
  PIN instr_slave_r_id[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 520.240 1500.000 520.840 ;
    END
  END instr_slave_r_id[5]
  PIN instr_slave_r_id[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 322.090 1796.000 322.370 1800.000 ;
    END
  END instr_slave_r_id[6]
  PIN instr_slave_r_id[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 473.430 1796.000 473.710 1800.000 ;
    END
  END instr_slave_r_id[7]
  PIN instr_slave_r_id[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 267.350 1796.000 267.630 1800.000 ;
    END
  END instr_slave_r_id[8]
  PIN instr_slave_r_id[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 515.290 1796.000 515.570 1800.000 ;
    END
  END instr_slave_r_id[9]
  PIN instr_slave_r_last
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1319.240 4.000 1319.840 ;
    END
  END instr_slave_r_last
  PIN instr_slave_r_ready
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1233.350 1796.000 1233.630 1800.000 ;
    END
  END instr_slave_r_ready
  PIN instr_slave_r_resp[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1417.840 4.000 1418.440 ;
    END
  END instr_slave_r_resp[0]
  PIN instr_slave_r_resp[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1381.470 0.000 1381.750 4.000 ;
    END
  END instr_slave_r_resp[1]
  PIN instr_slave_r_user[-1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 190.440 1500.000 191.040 ;
    END
  END instr_slave_r_user[-1]
  PIN instr_slave_r_user[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 937.110 0.000 937.390 4.000 ;
    END
  END instr_slave_r_user[0]
  PIN instr_slave_r_valid
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 370.640 4.000 371.240 ;
    END
  END instr_slave_r_valid
  PIN instr_slave_w_data[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 312.430 1796.000 312.710 1800.000 ;
    END
  END instr_slave_w_data[0]
  PIN instr_slave_w_data[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 219.050 1796.000 219.330 1800.000 ;
    END
  END instr_slave_w_data[10]
  PIN instr_slave_w_data[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1016.640 4.000 1017.240 ;
    END
  END instr_slave_w_data[11]
  PIN instr_slave_w_data[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 992.840 4.000 993.440 ;
    END
  END instr_slave_w_data[12]
  PIN instr_slave_w_data[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1679.640 4.000 1680.240 ;
    END
  END instr_slave_w_data[13]
  PIN instr_slave_w_data[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 463.770 0.000 464.050 4.000 ;
    END
  END instr_slave_w_data[14]
  PIN instr_slave_w_data[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1509.640 4.000 1510.240 ;
    END
  END instr_slave_w_data[15]
  PIN instr_slave_w_data[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 918.040 4.000 918.640 ;
    END
  END instr_slave_w_data[16]
  PIN instr_slave_w_data[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1304.190 0.000 1304.470 4.000 ;
    END
  END instr_slave_w_data[17]
  PIN instr_slave_w_data[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1213.840 1500.000 1214.440 ;
    END
  END instr_slave_w_data[18]
  PIN instr_slave_w_data[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1149.240 1500.000 1149.840 ;
    END
  END instr_slave_w_data[19]
  PIN instr_slave_w_data[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1152.640 4.000 1153.240 ;
    END
  END instr_slave_w_data[1]
  PIN instr_slave_w_data[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1560.640 4.000 1561.240 ;
    END
  END instr_slave_w_data[20]
  PIN instr_slave_w_data[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 599.010 1796.000 599.290 1800.000 ;
    END
  END instr_slave_w_data[21]
  PIN instr_slave_w_data[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 875.930 0.000 876.210 4.000 ;
    END
  END instr_slave_w_data[22]
  PIN instr_slave_w_data[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1384.690 1796.000 1384.970 1800.000 ;
    END
  END instr_slave_w_data[23]
  PIN instr_slave_w_data[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1149.630 0.000 1149.910 4.000 ;
    END
  END instr_slave_w_data[24]
  PIN instr_slave_w_data[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1297.750 0.000 1298.030 4.000 ;
    END
  END instr_slave_w_data[25]
  PIN instr_slave_w_data[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1194.710 1796.000 1194.990 1800.000 ;
    END
  END instr_slave_w_data[26]
  PIN instr_slave_w_data[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 273.790 1796.000 274.070 1800.000 ;
    END
  END instr_slave_w_data[27]
  PIN instr_slave_w_data[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1302.240 1500.000 1302.840 ;
    END
  END instr_slave_w_data[28]
  PIN instr_slave_w_data[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 404.640 4.000 405.240 ;
    END
  END instr_slave_w_data[29]
  PIN instr_slave_w_data[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 336.640 4.000 337.240 ;
    END
  END instr_slave_w_data[2]
  PIN instr_slave_w_data[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 570.030 0.000 570.310 4.000 ;
    END
  END instr_slave_w_data[30]
  PIN instr_slave_w_data[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 319.640 4.000 320.240 ;
    END
  END instr_slave_w_data[31]
  PIN instr_slave_w_data[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 241.440 1500.000 242.040 ;
    END
  END instr_slave_w_data[32]
  PIN instr_slave_w_data[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1275.210 1796.000 1275.490 1800.000 ;
    END
  END instr_slave_w_data[33]
  PIN instr_slave_w_data[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 695.610 0.000 695.890 4.000 ;
    END
  END instr_slave_w_data[34]
  PIN instr_slave_w_data[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 447.670 1796.000 447.950 1800.000 ;
    END
  END instr_slave_w_data[35]
  PIN instr_slave_w_data[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1737.440 4.000 1738.040 ;
    END
  END instr_slave_w_data[36]
  PIN instr_slave_w_data[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1196.840 1500.000 1197.440 ;
    END
  END instr_slave_w_data[37]
  PIN instr_slave_w_data[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 493.040 1500.000 493.640 ;
    END
  END instr_slave_w_data[38]
  PIN instr_slave_w_data[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 554.240 1500.000 554.840 ;
    END
  END instr_slave_w_data[39]
  PIN instr_slave_w_data[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 897.640 4.000 898.240 ;
    END
  END instr_slave_w_data[3]
  PIN instr_slave_w_data[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1700.040 4.000 1700.640 ;
    END
  END instr_slave_w_data[40]
  PIN instr_slave_w_data[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 888.810 0.000 889.090 4.000 ;
    END
  END instr_slave_w_data[41]
  PIN instr_slave_w_data[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 489.530 0.000 489.810 4.000 ;
    END
  END instr_slave_w_data[42]
  PIN instr_slave_w_data[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1407.230 1796.000 1407.510 1800.000 ;
    END
  END instr_slave_w_data[43]
  PIN instr_slave_w_data[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 299.240 1500.000 299.840 ;
    END
  END instr_slave_w_data[44]
  PIN instr_slave_w_data[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1159.290 0.000 1159.570 4.000 ;
    END
  END instr_slave_w_data[45]
  PIN instr_slave_w_data[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 553.930 1796.000 554.210 1800.000 ;
    END
  END instr_slave_w_data[46]
  PIN instr_slave_w_data[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1309.040 4.000 1309.640 ;
    END
  END instr_slave_w_data[47]
  PIN instr_slave_w_data[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1053.030 1796.000 1053.310 1800.000 ;
    END
  END instr_slave_w_data[48]
  PIN instr_slave_w_data[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 571.240 4.000 571.840 ;
    END
  END instr_slave_w_data[49]
  PIN instr_slave_w_data[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1130.310 0.000 1130.590 4.000 ;
    END
  END instr_slave_w_data[4]
  PIN instr_slave_w_data[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1220.470 1796.000 1220.750 1800.000 ;
    END
  END instr_slave_w_data[50]
  PIN instr_slave_w_data[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 187.040 1500.000 187.640 ;
    END
  END instr_slave_w_data[51]
  PIN instr_slave_w_data[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1628.640 1500.000 1629.240 ;
    END
  END instr_slave_w_data[52]
  PIN instr_slave_w_data[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 280.230 1796.000 280.510 1800.000 ;
    END
  END instr_slave_w_data[53]
  PIN instr_slave_w_data[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 333.240 4.000 333.840 ;
    END
  END instr_slave_w_data[54]
  PIN instr_slave_w_data[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 425.040 4.000 425.640 ;
    END
  END instr_slave_w_data[55]
  PIN instr_slave_w_data[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 962.870 0.000 963.150 4.000 ;
    END
  END instr_slave_w_data[56]
  PIN instr_slave_w_data[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1186.640 1500.000 1187.240 ;
    END
  END instr_slave_w_data[57]
  PIN instr_slave_w_data[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 166.640 1500.000 167.240 ;
    END
  END instr_slave_w_data[58]
  PIN instr_slave_w_data[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 776.110 0.000 776.390 4.000 ;
    END
  END instr_slave_w_data[59]
  PIN instr_slave_w_data[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 376.830 1796.000 377.110 1800.000 ;
    END
  END instr_slave_w_data[5]
  PIN instr_slave_w_data[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 563.590 1796.000 563.870 1800.000 ;
    END
  END instr_slave_w_data[60]
  PIN instr_slave_w_data[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 466.990 0.000 467.270 4.000 ;
    END
  END instr_slave_w_data[61]
  PIN instr_slave_w_data[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 843.240 4.000 843.840 ;
    END
  END instr_slave_w_data[62]
  PIN instr_slave_w_data[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1356.640 1500.000 1357.240 ;
    END
  END instr_slave_w_data[63]
  PIN instr_slave_w_data[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 601.840 1500.000 602.440 ;
    END
  END instr_slave_w_data[6]
  PIN instr_slave_w_data[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1268.240 4.000 1268.840 ;
    END
  END instr_slave_w_data[7]
  PIN instr_slave_w_data[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1360.040 4.000 1360.640 ;
    END
  END instr_slave_w_data[8]
  PIN instr_slave_w_data[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 136.040 4.000 136.640 ;
    END
  END instr_slave_w_data[9]
  PIN instr_slave_w_last
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1003.040 1500.000 1003.640 ;
    END
  END instr_slave_w_last
  PIN instr_slave_w_ready
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 646.040 4.000 646.640 ;
    END
  END instr_slave_w_ready
  PIN instr_slave_w_strb[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 508.850 1796.000 509.130 1800.000 ;
    END
  END instr_slave_w_strb[0]
  PIN instr_slave_w_strb[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 898.470 1796.000 898.750 1800.000 ;
    END
  END instr_slave_w_strb[1]
  PIN instr_slave_w_strb[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1190.040 4.000 1190.640 ;
    END
  END instr_slave_w_strb[2]
  PIN instr_slave_w_strb[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1239.790 0.000 1240.070 4.000 ;
    END
  END instr_slave_w_strb[3]
  PIN instr_slave_w_strb[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 455.640 1500.000 456.240 ;
    END
  END instr_slave_w_strb[4]
  PIN instr_slave_w_strb[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 714.930 1796.000 715.210 1800.000 ;
    END
  END instr_slave_w_strb[5]
  PIN instr_slave_w_strb[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 421.910 0.000 422.190 4.000 ;
    END
  END instr_slave_w_strb[6]
  PIN instr_slave_w_strb[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1175.390 1796.000 1175.670 1800.000 ;
    END
  END instr_slave_w_strb[7]
  PIN instr_slave_w_user[-1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1703.440 1500.000 1704.040 ;
    END
  END instr_slave_w_user[-1]
  PIN instr_slave_w_user[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1271.990 0.000 1272.270 4.000 ;
    END
  END instr_slave_w_user[0]
  PIN instr_slave_w_valid
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1020.040 4.000 1020.640 ;
    END
  END instr_slave_w_valid
  PIN irq_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1292.040 4.000 1292.640 ;
    END
  END irq_i[0]
  PIN irq_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 904.440 1500.000 905.040 ;
    END
  END irq_i[10]
  PIN irq_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1139.040 1500.000 1139.640 ;
    END
  END irq_i[11]
  PIN irq_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1071.040 4.000 1071.640 ;
    END
  END irq_i[12]
  PIN irq_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 760.010 0.000 760.290 4.000 ;
    END
  END irq_i[13]
  PIN irq_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1107.770 1796.000 1108.050 1800.000 ;
    END
  END irq_i[14]
  PIN irq_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1262.330 0.000 1262.610 4.000 ;
    END
  END irq_i[15]
  PIN irq_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1349.270 1796.000 1349.550 1800.000 ;
    END
  END irq_i[16]
  PIN irq_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1689.840 4.000 1690.440 ;
    END
  END irq_i[17]
  PIN irq_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 153.040 4.000 153.640 ;
    END
  END irq_i[18]
  PIN irq_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1474.850 0.000 1475.130 4.000 ;
    END
  END irq_i[19]
  PIN irq_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 788.840 4.000 789.440 ;
    END
  END irq_i[1]
  PIN irq_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 270.570 0.000 270.850 4.000 ;
    END
  END irq_i[20]
  PIN irq_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 720.840 1500.000 721.440 ;
    END
  END irq_i[21]
  PIN irq_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1234.240 1500.000 1234.840 ;
    END
  END irq_i[22]
  PIN irq_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1281.840 4.000 1282.440 ;
    END
  END irq_i[23]
  PIN irq_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1461.970 1796.000 1462.250 1800.000 ;
    END
  END irq_i[24]
  PIN irq_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1420.110 0.000 1420.390 4.000 ;
    END
  END irq_i[25]
  PIN irq_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 193.290 0.000 193.570 4.000 ;
    END
  END irq_i[26]
  PIN irq_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 625.640 4.000 626.240 ;
    END
  END irq_i[27]
  PIN irq_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 20.440 1500.000 21.040 ;
    END
  END irq_i[28]
  PIN irq_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 785.770 0.000 786.050 4.000 ;
    END
  END irq_i[29]
  PIN irq_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 112.240 1500.000 112.840 ;
    END
  END irq_i[2]
  PIN irq_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 30.640 4.000 31.240 ;
    END
  END irq_i[30]
  PIN irq_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1227.440 1500.000 1228.040 ;
    END
  END irq_i[31]
  PIN irq_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 975.750 1796.000 976.030 1800.000 ;
    END
  END irq_i[3]
  PIN irq_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1349.270 0.000 1349.550 4.000 ;
    END
  END irq_i[4]
  PIN irq_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1323.510 0.000 1323.790 4.000 ;
    END
  END irq_i[5]
  PIN irq_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1315.840 4.000 1316.440 ;
    END
  END irq_i[6]
  PIN irq_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1358.930 0.000 1359.210 4.000 ;
    END
  END irq_i[7]
  PIN irq_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1251.240 4.000 1251.840 ;
    END
  END irq_i[8]
  PIN irq_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 344.630 0.000 344.910 4.000 ;
    END
  END irq_i[9]
  PIN mba_data_mem_addr0_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 438.640 4.000 439.240 ;
    END
  END mba_data_mem_addr0_o[0]
  PIN mba_data_mem_addr0_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 710.640 1500.000 711.240 ;
    END
  END mba_data_mem_addr0_o[10]
  PIN mba_data_mem_addr0_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 914.570 1796.000 914.850 1800.000 ;
    END
  END mba_data_mem_addr0_o[11]
  PIN mba_data_mem_addr0_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1591.240 1500.000 1591.840 ;
    END
  END mba_data_mem_addr0_o[12]
  PIN mba_data_mem_addr0_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1373.640 1500.000 1374.240 ;
    END
  END mba_data_mem_addr0_o[13]
  PIN mba_data_mem_addr0_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1178.610 0.000 1178.890 4.000 ;
    END
  END mba_data_mem_addr0_o[14]
  PIN mba_data_mem_addr0_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 255.040 1500.000 255.640 ;
    END
  END mba_data_mem_addr0_o[15]
  PIN mba_data_mem_addr0_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 904.910 0.000 905.190 4.000 ;
    END
  END mba_data_mem_addr0_o[16]
  PIN mba_data_mem_addr0_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 6.840 4.000 7.440 ;
    END
  END mba_data_mem_addr0_o[17]
  PIN mba_data_mem_addr0_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1320.290 0.000 1320.570 4.000 ;
    END
  END mba_data_mem_addr0_o[18]
  PIN mba_data_mem_addr0_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 346.840 1500.000 347.440 ;
    END
  END mba_data_mem_addr0_o[19]
  PIN mba_data_mem_addr0_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 744.640 4.000 745.240 ;
    END
  END mba_data_mem_addr0_o[1]
  PIN mba_data_mem_addr0_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 650.530 0.000 650.810 4.000 ;
    END
  END mba_data_mem_addr0_o[20]
  PIN mba_data_mem_addr0_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 943.550 1796.000 943.830 1800.000 ;
    END
  END mba_data_mem_addr0_o[21]
  PIN mba_data_mem_addr0_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1204.370 0.000 1204.650 4.000 ;
    END
  END mba_data_mem_addr0_o[22]
  PIN mba_data_mem_addr0_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1200.240 1500.000 1200.840 ;
    END
  END mba_data_mem_addr0_o[23]
  PIN mba_data_mem_addr0_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 812.640 1500.000 813.240 ;
    END
  END mba_data_mem_addr0_o[24]
  PIN mba_data_mem_addr0_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1485.840 1500.000 1486.440 ;
    END
  END mba_data_mem_addr0_o[25]
  PIN mba_data_mem_addr0_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 248.240 4.000 248.840 ;
    END
  END mba_data_mem_addr0_o[26]
  PIN mba_data_mem_addr0_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 895.250 0.000 895.530 4.000 ;
    END
  END mba_data_mem_addr0_o[27]
  PIN mba_data_mem_addr0_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.510 0.000 35.790 4.000 ;
    END
  END mba_data_mem_addr0_o[28]
  PIN mba_data_mem_addr0_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 170.040 1500.000 170.640 ;
    END
  END mba_data_mem_addr0_o[29]
  PIN mba_data_mem_addr0_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.090 1796.000 0.370 1800.000 ;
    END
  END mba_data_mem_addr0_o[2]
  PIN mba_data_mem_addr0_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 448.840 1500.000 449.440 ;
    END
  END mba_data_mem_addr0_o[30]
  PIN mba_data_mem_addr0_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 225.490 1796.000 225.770 1800.000 ;
    END
  END mba_data_mem_addr0_o[31]
  PIN mba_data_mem_addr0_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.090 0.000 0.370 4.000 ;
    END
  END mba_data_mem_addr0_o[3]
  PIN mba_data_mem_addr0_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 884.040 1500.000 884.640 ;
    END
  END mba_data_mem_addr0_o[4]
  PIN mba_data_mem_addr0_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1152.850 1796.000 1153.130 1800.000 ;
    END
  END mba_data_mem_addr0_o[5]
  PIN mba_data_mem_addr0_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1249.450 0.000 1249.730 4.000 ;
    END
  END mba_data_mem_addr0_o[6]
  PIN mba_data_mem_addr0_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1490.950 0.000 1491.230 4.000 ;
    END
  END mba_data_mem_addr0_o[7]
  PIN mba_data_mem_addr0_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 602.230 0.000 602.510 4.000 ;
    END
  END mba_data_mem_addr0_o[8]
  PIN mba_data_mem_addr0_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1502.840 4.000 1503.440 ;
    END
  END mba_data_mem_addr0_o[9]
  PIN mba_data_mem_addr1_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 261.840 1500.000 262.440 ;
    END
  END mba_data_mem_addr1_o[0]
  PIN mba_data_mem_addr1_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 482.840 1500.000 483.440 ;
    END
  END mba_data_mem_addr1_o[10]
  PIN mba_data_mem_addr1_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 435.240 4.000 435.840 ;
    END
  END mba_data_mem_addr1_o[11]
  PIN mba_data_mem_addr1_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 544.040 4.000 544.640 ;
    END
  END mba_data_mem_addr1_o[12]
  PIN mba_data_mem_addr1_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 248.030 1796.000 248.310 1800.000 ;
    END
  END mba_data_mem_addr1_o[13]
  PIN mba_data_mem_addr1_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 302.640 1500.000 303.240 ;
    END
  END mba_data_mem_addr1_o[14]
  PIN mba_data_mem_addr1_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1560.640 1500.000 1561.240 ;
    END
  END mba_data_mem_addr1_o[15]
  PIN mba_data_mem_addr1_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1611.640 4.000 1612.240 ;
    END
  END mba_data_mem_addr1_o[16]
  PIN mba_data_mem_addr1_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 635.840 4.000 636.440 ;
    END
  END mba_data_mem_addr1_o[17]
  PIN mba_data_mem_addr1_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 836.440 4.000 837.040 ;
    END
  END mba_data_mem_addr1_o[18]
  PIN mba_data_mem_addr1_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1030.490 0.000 1030.770 4.000 ;
    END
  END mba_data_mem_addr1_o[19]
  PIN mba_data_mem_addr1_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1207.590 0.000 1207.870 4.000 ;
    END
  END mba_data_mem_addr1_o[1]
  PIN mba_data_mem_addr1_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 244.810 1796.000 245.090 1800.000 ;
    END
  END mba_data_mem_addr1_o[20]
  PIN mba_data_mem_addr1_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1088.040 1500.000 1088.640 ;
    END
  END mba_data_mem_addr1_o[21]
  PIN mba_data_mem_addr1_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1659.240 4.000 1659.840 ;
    END
  END mba_data_mem_addr1_o[22]
  PIN mba_data_mem_addr1_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 582.910 0.000 583.190 4.000 ;
    END
  END mba_data_mem_addr1_o[23]
  PIN mba_data_mem_addr1_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1181.830 1796.000 1182.110 1800.000 ;
    END
  END mba_data_mem_addr1_o[24]
  PIN mba_data_mem_addr1_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 149.640 1500.000 150.240 ;
    END
  END mba_data_mem_addr1_o[25]
  PIN mba_data_mem_addr1_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 202.950 1796.000 203.230 1800.000 ;
    END
  END mba_data_mem_addr1_o[26]
  PIN mba_data_mem_addr1_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1226.910 1796.000 1227.190 1800.000 ;
    END
  END mba_data_mem_addr1_o[27]
  PIN mba_data_mem_addr1_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1295.440 4.000 1296.040 ;
    END
  END mba_data_mem_addr1_o[28]
  PIN mba_data_mem_addr1_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1581.040 4.000 1581.640 ;
    END
  END mba_data_mem_addr1_o[29]
  PIN mba_data_mem_addr1_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 898.470 0.000 898.750 4.000 ;
    END
  END mba_data_mem_addr1_o[2]
  PIN mba_data_mem_addr1_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 821.190 1796.000 821.470 1800.000 ;
    END
  END mba_data_mem_addr1_o[30]
  PIN mba_data_mem_addr1_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 122.440 1500.000 123.040 ;
    END
  END mba_data_mem_addr1_o[31]
  PIN mba_data_mem_addr1_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1352.490 1796.000 1352.770 1800.000 ;
    END
  END mba_data_mem_addr1_o[3]
  PIN mba_data_mem_addr1_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 425.130 0.000 425.410 4.000 ;
    END
  END mba_data_mem_addr1_o[4]
  PIN mba_data_mem_addr1_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1193.440 4.000 1194.040 ;
    END
  END mba_data_mem_addr1_o[5]
  PIN mba_data_mem_addr1_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1281.650 0.000 1281.930 4.000 ;
    END
  END mba_data_mem_addr1_o[6]
  PIN mba_data_mem_addr1_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1136.750 0.000 1137.030 4.000 ;
    END
  END mba_data_mem_addr1_o[7]
  PIN mba_data_mem_addr1_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 463.770 1796.000 464.050 1800.000 ;
    END
  END mba_data_mem_addr1_o[8]
  PIN mba_data_mem_addr1_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1615.040 1500.000 1615.640 ;
    END
  END mba_data_mem_addr1_o[9]
  PIN mba_data_mem_csb0_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 850.040 1500.000 850.640 ;
    END
  END mba_data_mem_csb0_o
  PIN mba_data_mem_csb1_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1304.190 1796.000 1304.470 1800.000 ;
    END
  END mba_data_mem_csb1_o
  PIN mba_data_mem_din0_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1400.790 0.000 1401.070 4.000 ;
    END
  END mba_data_mem_din0_o[0]
  PIN mba_data_mem_din0_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 782.550 0.000 782.830 4.000 ;
    END
  END mba_data_mem_din0_o[10]
  PIN mba_data_mem_din0_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1370.240 4.000 1370.840 ;
    END
  END mba_data_mem_din0_o[11]
  PIN mba_data_mem_din0_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 779.330 1796.000 779.610 1800.000 ;
    END
  END mba_data_mem_din0_o[12]
  PIN mba_data_mem_din0_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1448.440 1500.000 1449.040 ;
    END
  END mba_data_mem_din0_o[13]
  PIN mba_data_mem_din0_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1771.440 1500.000 1772.040 ;
    END
  END mba_data_mem_din0_o[14]
  PIN mba_data_mem_din0_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 289.040 1500.000 289.640 ;
    END
  END mba_data_mem_din0_o[15]
  PIN mba_data_mem_din0_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1254.640 1500.000 1255.240 ;
    END
  END mba_data_mem_din0_o[16]
  PIN mba_data_mem_din0_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 102.040 4.000 102.640 ;
    END
  END mba_data_mem_din0_o[17]
  PIN mba_data_mem_din0_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1411.040 4.000 1411.640 ;
    END
  END mba_data_mem_din0_o[18]
  PIN mba_data_mem_din0_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 173.970 0.000 174.250 4.000 ;
    END
  END mba_data_mem_din0_o[19]
  PIN mba_data_mem_din0_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1139.970 0.000 1140.250 4.000 ;
    END
  END mba_data_mem_din0_o[1]
  PIN mba_data_mem_din0_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 608.670 0.000 608.950 4.000 ;
    END
  END mba_data_mem_din0_o[20]
  PIN mba_data_mem_din0_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1047.240 1500.000 1047.840 ;
    END
  END mba_data_mem_din0_o[21]
  PIN mba_data_mem_din0_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 146.240 4.000 146.840 ;
    END
  END mba_data_mem_din0_o[22]
  PIN mba_data_mem_din0_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 627.990 0.000 628.270 4.000 ;
    END
  END mba_data_mem_din0_o[23]
  PIN mba_data_mem_din0_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 982.640 1500.000 983.240 ;
    END
  END mba_data_mem_din0_o[24]
  PIN mba_data_mem_din0_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 656.970 1796.000 657.250 1800.000 ;
    END
  END mba_data_mem_din0_o[25]
  PIN mba_data_mem_din0_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1557.240 1500.000 1557.840 ;
    END
  END mba_data_mem_din0_o[26]
  PIN mba_data_mem_din0_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 225.490 0.000 225.770 4.000 ;
    END
  END mba_data_mem_din0_o[27]
  PIN mba_data_mem_din0_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1387.240 1500.000 1387.840 ;
    END
  END mba_data_mem_din0_o[28]
  PIN mba_data_mem_din0_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1461.970 0.000 1462.250 4.000 ;
    END
  END mba_data_mem_din0_o[29]
  PIN mba_data_mem_din0_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 299.550 1796.000 299.830 1800.000 ;
    END
  END mba_data_mem_din0_o[2]
  PIN mba_data_mem_din0_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1346.050 0.000 1346.330 4.000 ;
    END
  END mba_data_mem_din0_o[30]
  PIN mba_data_mem_din0_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1494.170 1796.000 1494.450 1800.000 ;
    END
  END mba_data_mem_din0_o[31]
  PIN mba_data_mem_din0_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 576.470 1796.000 576.750 1800.000 ;
    END
  END mba_data_mem_din0_o[3]
  PIN mba_data_mem_din0_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 347.850 1796.000 348.130 1800.000 ;
    END
  END mba_data_mem_din0_o[4]
  PIN mba_data_mem_din0_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1632.040 4.000 1632.640 ;
    END
  END mba_data_mem_din0_o[5]
  PIN mba_data_mem_din0_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 618.330 1796.000 618.610 1800.000 ;
    END
  END mba_data_mem_din0_o[6]
  PIN mba_data_mem_din0_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 880.640 4.000 881.240 ;
    END
  END mba_data_mem_din0_o[7]
  PIN mba_data_mem_din0_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 682.730 0.000 683.010 4.000 ;
    END
  END mba_data_mem_din0_o[8]
  PIN mba_data_mem_din0_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 734.440 1500.000 735.040 ;
    END
  END mba_data_mem_din0_o[9]
  PIN mba_data_mem_dout0_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1281.840 1500.000 1282.440 ;
    END
  END mba_data_mem_dout0_i[0]
  PIN mba_data_mem_dout0_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1478.070 1796.000 1478.350 1800.000 ;
    END
  END mba_data_mem_dout0_i[10]
  PIN mba_data_mem_dout0_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1377.040 4.000 1377.640 ;
    END
  END mba_data_mem_dout0_i[11]
  PIN mba_data_mem_dout0_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 85.040 1500.000 85.640 ;
    END
  END mba_data_mem_dout0_i[12]
  PIN mba_data_mem_dout0_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 221.040 4.000 221.640 ;
    END
  END mba_data_mem_dout0_i[13]
  PIN mba_data_mem_dout0_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1294.530 1796.000 1294.810 1800.000 ;
    END
  END mba_data_mem_dout0_i[14]
  PIN mba_data_mem_dout0_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 495.970 1796.000 496.250 1800.000 ;
    END
  END mba_data_mem_dout0_i[15]
  PIN mba_data_mem_dout0_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 204.040 4.000 204.640 ;
    END
  END mba_data_mem_dout0_i[16]
  PIN mba_data_mem_dout0_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 397.840 1500.000 398.440 ;
    END
  END mba_data_mem_dout0_i[17]
  PIN mba_data_mem_dout0_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 837.290 1796.000 837.570 1800.000 ;
    END
  END mba_data_mem_dout0_i[18]
  PIN mba_data_mem_dout0_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 312.840 1500.000 313.440 ;
    END
  END mba_data_mem_dout0_i[19]
  PIN mba_data_mem_dout0_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 680.040 1500.000 680.640 ;
    END
  END mba_data_mem_dout0_i[1]
  PIN mba_data_mem_dout0_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 51.040 4.000 51.640 ;
    END
  END mba_data_mem_dout0_i[20]
  PIN mba_data_mem_dout0_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 550.710 0.000 550.990 4.000 ;
    END
  END mba_data_mem_dout0_i[21]
  PIN mba_data_mem_dout0_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 442.040 1500.000 442.640 ;
    END
  END mba_data_mem_dout0_i[22]
  PIN mba_data_mem_dout0_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1166.240 1500.000 1166.840 ;
    END
  END mba_data_mem_dout0_i[23]
  PIN mba_data_mem_dout0_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1085.230 1796.000 1085.510 1800.000 ;
    END
  END mba_data_mem_dout0_i[24]
  PIN mba_data_mem_dout0_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1553.840 4.000 1554.440 ;
    END
  END mba_data_mem_dout0_i[25]
  PIN mba_data_mem_dout0_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1472.240 4.000 1472.840 ;
    END
  END mba_data_mem_dout0_i[26]
  PIN mba_data_mem_dout0_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 234.640 4.000 235.240 ;
    END
  END mba_data_mem_dout0_i[27]
  PIN mba_data_mem_dout0_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 673.070 0.000 673.350 4.000 ;
    END
  END mba_data_mem_dout0_i[28]
  PIN mba_data_mem_dout0_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 911.350 1796.000 911.630 1800.000 ;
    END
  END mba_data_mem_dout0_i[29]
  PIN mba_data_mem_dout0_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 622.240 1500.000 622.840 ;
    END
  END mba_data_mem_dout0_i[2]
  PIN mba_data_mem_dout0_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1064.240 4.000 1064.840 ;
    END
  END mba_data_mem_dout0_i[30]
  PIN mba_data_mem_dout0_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 431.570 0.000 431.850 4.000 ;
    END
  END mba_data_mem_dout0_i[31]
  PIN mba_data_mem_dout0_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1168.950 1796.000 1169.230 1800.000 ;
    END
  END mba_data_mem_dout0_i[3]
  PIN mba_data_mem_dout0_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 196.510 1796.000 196.790 1800.000 ;
    END
  END mba_data_mem_dout0_i[4]
  PIN mba_data_mem_dout0_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 83.810 1796.000 84.090 1800.000 ;
    END
  END mba_data_mem_dout0_i[5]
  PIN mba_data_mem_dout0_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 438.010 1796.000 438.290 1800.000 ;
    END
  END mba_data_mem_dout0_i[6]
  PIN mba_data_mem_dout0_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 537.830 1796.000 538.110 1800.000 ;
    END
  END mba_data_mem_dout0_i[7]
  PIN mba_data_mem_dout0_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 560.370 1796.000 560.650 1800.000 ;
    END
  END mba_data_mem_dout0_i[8]
  PIN mba_data_mem_dout0_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1162.510 0.000 1162.790 4.000 ;
    END
  END mba_data_mem_dout0_i[9]
  PIN mba_data_mem_web0_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1720.440 4.000 1721.040 ;
    END
  END mba_data_mem_web0_o
  PIN mba_data_mem_wmask0_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 258.440 4.000 259.040 ;
    END
  END mba_data_mem_wmask0_o[0]
  PIN mba_data_mem_wmask0_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.070 0.000 29.350 4.000 ;
    END
  END mba_data_mem_wmask0_o[1]
  PIN mba_data_mem_wmask0_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 238.040 1500.000 238.640 ;
    END
  END mba_data_mem_wmask0_o[2]
  PIN mba_data_mem_wmask0_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1165.730 0.000 1166.010 4.000 ;
    END
  END mba_data_mem_wmask0_o[3]
  PIN mba_instr_mem_addr0_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 870.440 1500.000 871.040 ;
    END
  END mba_instr_mem_addr0_o[0]
  PIN mba_instr_mem_addr0_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 154.650 1796.000 154.930 1800.000 ;
    END
  END mba_instr_mem_addr0_o[10]
  PIN mba_instr_mem_addr0_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1050.640 1500.000 1051.240 ;
    END
  END mba_instr_mem_addr0_o[11]
  PIN mba_instr_mem_addr0_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 622.240 4.000 622.840 ;
    END
  END mba_instr_mem_addr0_o[12]
  PIN mba_instr_mem_addr0_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.030 0.000 87.310 4.000 ;
    END
  END mba_instr_mem_addr0_o[13]
  PIN mba_instr_mem_addr0_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 438.010 0.000 438.290 4.000 ;
    END
  END mba_instr_mem_addr0_o[14]
  PIN mba_instr_mem_addr0_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 972.530 0.000 972.810 4.000 ;
    END
  END mba_instr_mem_addr0_o[15]
  PIN mba_instr_mem_addr0_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1761.240 4.000 1761.840 ;
    END
  END mba_instr_mem_addr0_o[16]
  PIN mba_instr_mem_addr0_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 265.240 1500.000 265.840 ;
    END
  END mba_instr_mem_addr0_o[17]
  PIN mba_instr_mem_addr0_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 830.850 0.000 831.130 4.000 ;
    END
  END mba_instr_mem_addr0_o[18]
  PIN mba_instr_mem_addr0_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 139.440 1500.000 140.040 ;
    END
  END mba_instr_mem_addr0_o[19]
  PIN mba_instr_mem_addr0_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1487.730 1796.000 1488.010 1800.000 ;
    END
  END mba_instr_mem_addr0_o[1]
  PIN mba_instr_mem_addr0_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1104.550 1796.000 1104.830 1800.000 ;
    END
  END mba_instr_mem_addr0_o[20]
  PIN mba_instr_mem_addr0_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 173.440 1500.000 174.040 ;
    END
  END mba_instr_mem_addr0_o[21]
  PIN mba_instr_mem_addr0_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 717.440 4.000 718.040 ;
    END
  END mba_instr_mem_addr0_o[22]
  PIN mba_instr_mem_addr0_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 61.240 4.000 61.840 ;
    END
  END mba_instr_mem_addr0_o[23]
  PIN mba_instr_mem_addr0_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1217.250 1796.000 1217.530 1800.000 ;
    END
  END mba_instr_mem_addr0_o[24]
  PIN mba_instr_mem_addr0_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1567.440 4.000 1568.040 ;
    END
  END mba_instr_mem_addr0_o[25]
  PIN mba_instr_mem_addr0_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1490.950 1796.000 1491.230 1800.000 ;
    END
  END mba_instr_mem_addr0_o[26]
  PIN mba_instr_mem_addr0_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 119.040 1500.000 119.640 ;
    END
  END mba_instr_mem_addr0_o[27]
  PIN mba_instr_mem_addr0_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 251.250 1796.000 251.530 1800.000 ;
    END
  END mba_instr_mem_addr0_o[28]
  PIN mba_instr_mem_addr0_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 860.240 1500.000 860.840 ;
    END
  END mba_instr_mem_addr0_o[29]
  PIN mba_instr_mem_addr0_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1448.440 4.000 1449.040 ;
    END
  END mba_instr_mem_addr0_o[2]
  PIN mba_instr_mem_addr0_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 465.840 1500.000 466.440 ;
    END
  END mba_instr_mem_addr0_o[30]
  PIN mba_instr_mem_addr0_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 703.840 4.000 704.440 ;
    END
  END mba_instr_mem_addr0_o[31]
  PIN mba_instr_mem_addr0_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 267.350 0.000 267.630 4.000 ;
    END
  END mba_instr_mem_addr0_o[3]
  PIN mba_instr_mem_addr0_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1706.840 1500.000 1707.440 ;
    END
  END mba_instr_mem_addr0_o[4]
  PIN mba_instr_mem_addr0_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 13.640 4.000 14.240 ;
    END
  END mba_instr_mem_addr0_o[5]
  PIN mba_instr_mem_addr0_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1291.310 1796.000 1291.590 1800.000 ;
    END
  END mba_instr_mem_addr0_o[6]
  PIN mba_instr_mem_addr0_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 528.170 0.000 528.450 4.000 ;
    END
  END mba_instr_mem_addr0_o[7]
  PIN mba_instr_mem_addr0_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 479.440 1500.000 480.040 ;
    END
  END mba_instr_mem_addr0_o[8]
  PIN mba_instr_mem_addr0_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 928.240 4.000 928.840 ;
    END
  END mba_instr_mem_addr0_o[9]
  PIN mba_instr_mem_addr1_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 338.190 1796.000 338.470 1800.000 ;
    END
  END mba_instr_mem_addr1_o[0]
  PIN mba_instr_mem_addr1_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1110.990 1796.000 1111.270 1800.000 ;
    END
  END mba_instr_mem_addr1_o[10]
  PIN mba_instr_mem_addr1_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 887.440 4.000 888.040 ;
    END
  END mba_instr_mem_addr1_o[11]
  PIN mba_instr_mem_addr1_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1088.040 4.000 1088.640 ;
    END
  END mba_instr_mem_addr1_o[12]
  PIN mba_instr_mem_addr1_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 210.840 4.000 211.440 ;
    END
  END mba_instr_mem_addr1_o[13]
  PIN mba_instr_mem_addr1_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 795.640 4.000 796.240 ;
    END
  END mba_instr_mem_addr1_o[14]
  PIN mba_instr_mem_addr1_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 142.840 4.000 143.440 ;
    END
  END mba_instr_mem_addr1_o[15]
  PIN mba_instr_mem_addr1_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.070 1796.000 29.350 1800.000 ;
    END
  END mba_instr_mem_addr1_o[16]
  PIN mba_instr_mem_addr1_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 329.840 4.000 330.440 ;
    END
  END mba_instr_mem_addr1_o[17]
  PIN mba_instr_mem_addr1_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 588.240 4.000 588.840 ;
    END
  END mba_instr_mem_addr1_o[18]
  PIN mba_instr_mem_addr1_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 183.630 0.000 183.910 4.000 ;
    END
  END mba_instr_mem_addr1_o[19]
  PIN mba_instr_mem_addr1_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1114.210 0.000 1114.490 4.000 ;
    END
  END mba_instr_mem_addr1_o[1]
  PIN mba_instr_mem_addr1_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1271.990 1796.000 1272.270 1800.000 ;
    END
  END mba_instr_mem_addr1_o[20]
  PIN mba_instr_mem_addr1_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1394.350 1796.000 1394.630 1800.000 ;
    END
  END mba_instr_mem_addr1_o[21]
  PIN mba_instr_mem_addr1_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1255.890 0.000 1256.170 4.000 ;
    END
  END mba_instr_mem_addr1_o[22]
  PIN mba_instr_mem_addr1_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1740.840 1500.000 1741.440 ;
    END
  END mba_instr_mem_addr1_o[23]
  PIN mba_instr_mem_addr1_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1135.640 1500.000 1136.240 ;
    END
  END mba_instr_mem_addr1_o[24]
  PIN mba_instr_mem_addr1_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 408.040 1500.000 408.640 ;
    END
  END mba_instr_mem_addr1_o[25]
  PIN mba_instr_mem_addr1_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 119.230 1796.000 119.510 1800.000 ;
    END
  END mba_instr_mem_addr1_o[26]
  PIN mba_instr_mem_addr1_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 679.510 1796.000 679.790 1800.000 ;
    END
  END mba_instr_mem_addr1_o[27]
  PIN mba_instr_mem_addr1_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1104.550 0.000 1104.830 4.000 ;
    END
  END mba_instr_mem_addr1_o[28]
  PIN mba_instr_mem_addr1_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 74.840 1500.000 75.440 ;
    END
  END mba_instr_mem_addr1_o[29]
  PIN mba_instr_mem_addr1_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 928.240 1500.000 928.840 ;
    END
  END mba_instr_mem_addr1_o[2]
  PIN mba_instr_mem_addr1_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 921.440 4.000 922.040 ;
    END
  END mba_instr_mem_addr1_o[30]
  PIN mba_instr_mem_addr1_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1056.250 0.000 1056.530 4.000 ;
    END
  END mba_instr_mem_addr1_o[31]
  PIN mba_instr_mem_addr1_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 206.170 0.000 206.450 4.000 ;
    END
  END mba_instr_mem_addr1_o[3]
  PIN mba_instr_mem_addr1_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1400.840 4.000 1401.440 ;
    END
  END mba_instr_mem_addr1_o[4]
  PIN mba_instr_mem_addr1_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1608.240 1500.000 1608.840 ;
    END
  END mba_instr_mem_addr1_o[5]
  PIN mba_instr_mem_addr1_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 978.970 1796.000 979.250 1800.000 ;
    END
  END mba_instr_mem_addr1_o[6]
  PIN mba_instr_mem_addr1_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 743.910 0.000 744.190 4.000 ;
    END
  END mba_instr_mem_addr1_o[7]
  PIN mba_instr_mem_addr1_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 528.170 1796.000 528.450 1800.000 ;
    END
  END mba_instr_mem_addr1_o[8]
  PIN mba_instr_mem_addr1_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1258.040 1500.000 1258.640 ;
    END
  END mba_instr_mem_addr1_o[9]
  PIN mba_instr_mem_csb0_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1471.630 0.000 1471.910 4.000 ;
    END
  END mba_instr_mem_csb0_o
  PIN mba_instr_mem_csb1_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 512.070 1796.000 512.350 1800.000 ;
    END
  END mba_instr_mem_csb1_o
  PIN mba_instr_mem_din0_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1413.670 0.000 1413.950 4.000 ;
    END
  END mba_instr_mem_din0_o[0]
  PIN mba_instr_mem_din0_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 599.010 0.000 599.290 4.000 ;
    END
  END mba_instr_mem_din0_o[10]
  PIN mba_instr_mem_din0_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 96.690 0.000 96.970 4.000 ;
    END
  END mba_instr_mem_din0_o[11]
  PIN mba_instr_mem_din0_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 391.040 1500.000 391.640 ;
    END
  END mba_instr_mem_din0_o[12]
  PIN mba_instr_mem_din0_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 918.040 1500.000 918.640 ;
    END
  END mba_instr_mem_din0_o[13]
  PIN mba_instr_mem_din0_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1519.840 4.000 1520.440 ;
    END
  END mba_instr_mem_din0_o[14]
  PIN mba_instr_mem_din0_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1239.790 1796.000 1240.070 1800.000 ;
    END
  END mba_instr_mem_din0_o[15]
  PIN mba_instr_mem_din0_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 489.640 4.000 490.240 ;
    END
  END mba_instr_mem_din0_o[16]
  PIN mba_instr_mem_din0_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 639.240 4.000 639.840 ;
    END
  END mba_instr_mem_din0_o[17]
  PIN mba_instr_mem_din0_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 591.640 4.000 592.240 ;
    END
  END mba_instr_mem_din0_o[18]
  PIN mba_instr_mem_din0_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 80.590 0.000 80.870 4.000 ;
    END
  END mba_instr_mem_din0_o[19]
  PIN mba_instr_mem_din0_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 396.150 0.000 396.430 4.000 ;
    END
  END mba_instr_mem_din0_o[1]
  PIN mba_instr_mem_din0_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1353.240 1500.000 1353.840 ;
    END
  END mba_instr_mem_din0_o[20]
  PIN mba_instr_mem_din0_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1049.810 0.000 1050.090 4.000 ;
    END
  END mba_instr_mem_din0_o[21]
  PIN mba_instr_mem_din0_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 499.190 1796.000 499.470 1800.000 ;
    END
  END mba_instr_mem_din0_o[22]
  PIN mba_instr_mem_din0_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 946.770 1796.000 947.050 1800.000 ;
    END
  END mba_instr_mem_din0_o[23]
  PIN mba_instr_mem_din0_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1149.240 4.000 1149.840 ;
    END
  END mba_instr_mem_din0_o[24]
  PIN mba_instr_mem_din0_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 283.450 0.000 283.730 4.000 ;
    END
  END mba_instr_mem_din0_o[25]
  PIN mba_instr_mem_din0_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1468.840 1500.000 1469.440 ;
    END
  END mba_instr_mem_din0_o[26]
  PIN mba_instr_mem_din0_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1030.490 1796.000 1030.770 1800.000 ;
    END
  END mba_instr_mem_din0_o[27]
  PIN mba_instr_mem_din0_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 323.040 4.000 323.640 ;
    END
  END mba_instr_mem_din0_o[28]
  PIN mba_instr_mem_din0_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1785.040 1500.000 1785.640 ;
    END
  END mba_instr_mem_din0_o[29]
  PIN mba_instr_mem_din0_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 924.840 1500.000 925.440 ;
    END
  END mba_instr_mem_din0_o[2]
  PIN mba_instr_mem_din0_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1236.570 0.000 1236.850 4.000 ;
    END
  END mba_instr_mem_din0_o[30]
  PIN mba_instr_mem_din0_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 132.640 4.000 133.240 ;
    END
  END mba_instr_mem_din0_o[31]
  PIN mba_instr_mem_din0_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1608.240 4.000 1608.840 ;
    END
  END mba_instr_mem_din0_o[3]
  PIN mba_instr_mem_din0_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 560.370 0.000 560.650 4.000 ;
    END
  END mba_instr_mem_din0_o[4]
  PIN mba_instr_mem_din0_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 37.440 4.000 38.040 ;
    END
  END mba_instr_mem_din0_o[5]
  PIN mba_instr_mem_din0_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1449.090 0.000 1449.370 4.000 ;
    END
  END mba_instr_mem_din0_o[6]
  PIN mba_instr_mem_din0_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 826.240 1500.000 826.840 ;
    END
  END mba_instr_mem_din0_o[7]
  PIN mba_instr_mem_din0_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 350.240 4.000 350.840 ;
    END
  END mba_instr_mem_din0_o[8]
  PIN mba_instr_mem_din0_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 340.040 1500.000 340.640 ;
    END
  END mba_instr_mem_din0_o[9]
  PIN mba_instr_mem_dout0_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 289.890 0.000 290.170 4.000 ;
    END
  END mba_instr_mem_dout0_i[0]
  PIN mba_instr_mem_dout0_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 869.490 0.000 869.770 4.000 ;
    END
  END mba_instr_mem_dout0_i[10]
  PIN mba_instr_mem_dout0_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1054.040 1500.000 1054.640 ;
    END
  END mba_instr_mem_dout0_i[11]
  PIN mba_instr_mem_dout0_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 872.710 1796.000 872.990 1800.000 ;
    END
  END mba_instr_mem_dout0_i[12]
  PIN mba_instr_mem_dout0_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1416.890 1796.000 1417.170 1800.000 ;
    END
  END mba_instr_mem_dout0_i[13]
  PIN mba_instr_mem_dout0_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 343.440 1500.000 344.040 ;
    END
  END mba_instr_mem_dout0_i[14]
  PIN mba_instr_mem_dout0_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 138.550 0.000 138.830 4.000 ;
    END
  END mba_instr_mem_dout0_i[15]
  PIN mba_instr_mem_dout0_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1278.440 1500.000 1279.040 ;
    END
  END mba_instr_mem_dout0_i[16]
  PIN mba_instr_mem_dout0_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 38.730 0.000 39.010 4.000 ;
    END
  END mba_instr_mem_dout0_i[17]
  PIN mba_instr_mem_dout0_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1410.450 1796.000 1410.730 1800.000 ;
    END
  END mba_instr_mem_dout0_i[18]
  PIN mba_instr_mem_dout0_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 859.830 1796.000 860.110 1800.000 ;
    END
  END mba_instr_mem_dout0_i[19]
  PIN mba_instr_mem_dout0_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 431.840 1500.000 432.440 ;
    END
  END mba_instr_mem_dout0_i[1]
  PIN mba_instr_mem_dout0_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 817.970 1796.000 818.250 1800.000 ;
    END
  END mba_instr_mem_dout0_i[20]
  PIN mba_instr_mem_dout0_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1152.850 0.000 1153.130 4.000 ;
    END
  END mba_instr_mem_dout0_i[21]
  PIN mba_instr_mem_dout0_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 166.640 4.000 167.240 ;
    END
  END mba_instr_mem_dout0_i[22]
  PIN mba_instr_mem_dout0_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1143.190 0.000 1143.470 4.000 ;
    END
  END mba_instr_mem_dout0_i[23]
  PIN mba_instr_mem_dout0_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3.310 0.000 3.590 4.000 ;
    END
  END mba_instr_mem_dout0_i[24]
  PIN mba_instr_mem_dout0_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1336.390 0.000 1336.670 4.000 ;
    END
  END mba_instr_mem_dout0_i[25]
  PIN mba_instr_mem_dout0_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 510.040 4.000 510.640 ;
    END
  END mba_instr_mem_dout0_i[26]
  PIN mba_instr_mem_dout0_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1213.840 4.000 1214.440 ;
    END
  END mba_instr_mem_dout0_i[27]
  PIN mba_instr_mem_dout0_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 138.550 1796.000 138.830 1800.000 ;
    END
  END mba_instr_mem_dout0_i[28]
  PIN mba_instr_mem_dout0_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 289.040 4.000 289.640 ;
    END
  END mba_instr_mem_dout0_i[29]
  PIN mba_instr_mem_dout0_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 354.290 0.000 354.570 4.000 ;
    END
  END mba_instr_mem_dout0_i[2]
  PIN mba_instr_mem_dout0_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 128.890 0.000 129.170 4.000 ;
    END
  END mba_instr_mem_dout0_i[30]
  PIN mba_instr_mem_dout0_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 579.690 1796.000 579.970 1800.000 ;
    END
  END mba_instr_mem_dout0_i[31]
  PIN mba_instr_mem_dout0_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 215.830 1796.000 216.110 1800.000 ;
    END
  END mba_instr_mem_dout0_i[3]
  PIN mba_instr_mem_dout0_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 901.690 0.000 901.970 4.000 ;
    END
  END mba_instr_mem_dout0_i[4]
  PIN mba_instr_mem_dout0_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 888.810 1796.000 889.090 1800.000 ;
    END
  END mba_instr_mem_dout0_i[5]
  PIN mba_instr_mem_dout0_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 652.840 1500.000 653.440 ;
    END
  END mba_instr_mem_dout0_i[6]
  PIN mba_instr_mem_dout0_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 952.040 4.000 952.640 ;
    END
  END mba_instr_mem_dout0_i[7]
  PIN mba_instr_mem_dout0_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1499.440 1500.000 1500.040 ;
    END
  END mba_instr_mem_dout0_i[8]
  PIN mba_instr_mem_dout0_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 367.170 0.000 367.450 4.000 ;
    END
  END mba_instr_mem_dout0_i[9]
  PIN mba_instr_mem_web0_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 634.430 0.000 634.710 4.000 ;
    END
  END mba_instr_mem_web0_o
  PIN mba_instr_mem_wmask0_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 34.040 4.000 34.640 ;
    END
  END mba_instr_mem_wmask0_o[0]
  PIN mba_instr_mem_wmask0_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1414.440 1500.000 1415.040 ;
    END
  END mba_instr_mem_wmask0_o[1]
  PIN mba_instr_mem_wmask0_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 991.850 0.000 992.130 4.000 ;
    END
  END mba_instr_mem_wmask0_o[2]
  PIN mba_instr_mem_wmask0_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 895.250 1796.000 895.530 1800.000 ;
    END
  END mba_instr_mem_wmask0_o[3]
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 882.370 1796.000 882.650 1800.000 ;
    END
  END rst_n
  PIN tck_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1506.240 4.000 1506.840 ;
    END
  END tck_i
  PIN tdi_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.630 1796.000 22.910 1800.000 ;
    END
  END tdi_i
  PIN tdo_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1168.950 0.000 1169.230 4.000 ;
    END
  END tdo_o
  PIN testmode_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 340.040 4.000 340.640 ;
    END
  END testmode_i
  PIN tms_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1380.440 4.000 1381.040 ;
    END
  END tms_i
  PIN trstn_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 948.640 1500.000 949.240 ;
    END
  END trstn_i
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 1787.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 1787.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 1787.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 1787.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 635.440 10.640 637.040 1787.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 789.040 10.640 790.640 1787.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 942.640 10.640 944.240 1787.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 1096.240 10.640 1097.840 1787.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 1249.840 10.640 1251.440 1787.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 1403.440 10.640 1405.040 1787.280 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 1787.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 1787.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 1787.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 558.640 10.640 560.240 1787.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 712.240 10.640 713.840 1787.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 865.840 10.640 867.440 1787.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 1019.440 10.640 1021.040 1787.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 1173.040 10.640 1174.640 1787.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 1326.640 10.640 1328.240 1787.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 1480.240 10.640 1481.840 1787.280 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 1494.080 1787.125 ;
      LAYER met1 ;
        RECT 0.070 6.500 1498.150 1787.280 ;
      LAYER met2 ;
        RECT 0.650 1795.720 3.030 1799.125 ;
        RECT 3.870 1795.720 6.250 1799.125 ;
        RECT 7.090 1795.720 9.470 1799.125 ;
        RECT 10.310 1795.720 12.690 1799.125 ;
        RECT 13.530 1795.720 19.130 1799.125 ;
        RECT 19.970 1795.720 22.350 1799.125 ;
        RECT 23.190 1795.720 25.570 1799.125 ;
        RECT 26.410 1795.720 28.790 1799.125 ;
        RECT 29.630 1795.720 32.010 1799.125 ;
        RECT 32.850 1795.720 35.230 1799.125 ;
        RECT 36.070 1795.720 41.670 1799.125 ;
        RECT 42.510 1795.720 44.890 1799.125 ;
        RECT 45.730 1795.720 48.110 1799.125 ;
        RECT 48.950 1795.720 51.330 1799.125 ;
        RECT 52.170 1795.720 54.550 1799.125 ;
        RECT 55.390 1795.720 57.770 1799.125 ;
        RECT 58.610 1795.720 60.990 1799.125 ;
        RECT 61.830 1795.720 67.430 1799.125 ;
        RECT 68.270 1795.720 70.650 1799.125 ;
        RECT 71.490 1795.720 73.870 1799.125 ;
        RECT 74.710 1795.720 77.090 1799.125 ;
        RECT 77.930 1795.720 80.310 1799.125 ;
        RECT 81.150 1795.720 83.530 1799.125 ;
        RECT 84.370 1795.720 89.970 1799.125 ;
        RECT 90.810 1795.720 93.190 1799.125 ;
        RECT 94.030 1795.720 96.410 1799.125 ;
        RECT 97.250 1795.720 99.630 1799.125 ;
        RECT 100.470 1795.720 102.850 1799.125 ;
        RECT 103.690 1795.720 106.070 1799.125 ;
        RECT 106.910 1795.720 112.510 1799.125 ;
        RECT 113.350 1795.720 115.730 1799.125 ;
        RECT 116.570 1795.720 118.950 1799.125 ;
        RECT 119.790 1795.720 122.170 1799.125 ;
        RECT 123.010 1795.720 125.390 1799.125 ;
        RECT 126.230 1795.720 128.610 1799.125 ;
        RECT 129.450 1795.720 131.830 1799.125 ;
        RECT 132.670 1795.720 138.270 1799.125 ;
        RECT 139.110 1795.720 141.490 1799.125 ;
        RECT 142.330 1795.720 144.710 1799.125 ;
        RECT 145.550 1795.720 147.930 1799.125 ;
        RECT 148.770 1795.720 151.150 1799.125 ;
        RECT 151.990 1795.720 154.370 1799.125 ;
        RECT 155.210 1795.720 160.810 1799.125 ;
        RECT 161.650 1795.720 164.030 1799.125 ;
        RECT 164.870 1795.720 167.250 1799.125 ;
        RECT 168.090 1795.720 170.470 1799.125 ;
        RECT 171.310 1795.720 173.690 1799.125 ;
        RECT 174.530 1795.720 176.910 1799.125 ;
        RECT 177.750 1795.720 180.130 1799.125 ;
        RECT 180.970 1795.720 186.570 1799.125 ;
        RECT 187.410 1795.720 189.790 1799.125 ;
        RECT 190.630 1795.720 193.010 1799.125 ;
        RECT 193.850 1795.720 196.230 1799.125 ;
        RECT 197.070 1795.720 199.450 1799.125 ;
        RECT 200.290 1795.720 202.670 1799.125 ;
        RECT 203.510 1795.720 209.110 1799.125 ;
        RECT 209.950 1795.720 212.330 1799.125 ;
        RECT 213.170 1795.720 215.550 1799.125 ;
        RECT 216.390 1795.720 218.770 1799.125 ;
        RECT 219.610 1795.720 221.990 1799.125 ;
        RECT 222.830 1795.720 225.210 1799.125 ;
        RECT 226.050 1795.720 228.430 1799.125 ;
        RECT 229.270 1795.720 234.870 1799.125 ;
        RECT 235.710 1795.720 238.090 1799.125 ;
        RECT 238.930 1795.720 241.310 1799.125 ;
        RECT 242.150 1795.720 244.530 1799.125 ;
        RECT 245.370 1795.720 247.750 1799.125 ;
        RECT 248.590 1795.720 250.970 1799.125 ;
        RECT 251.810 1795.720 257.410 1799.125 ;
        RECT 258.250 1795.720 260.630 1799.125 ;
        RECT 261.470 1795.720 263.850 1799.125 ;
        RECT 264.690 1795.720 267.070 1799.125 ;
        RECT 267.910 1795.720 270.290 1799.125 ;
        RECT 271.130 1795.720 273.510 1799.125 ;
        RECT 274.350 1795.720 279.950 1799.125 ;
        RECT 280.790 1795.720 283.170 1799.125 ;
        RECT 284.010 1795.720 286.390 1799.125 ;
        RECT 287.230 1795.720 289.610 1799.125 ;
        RECT 290.450 1795.720 292.830 1799.125 ;
        RECT 293.670 1795.720 296.050 1799.125 ;
        RECT 296.890 1795.720 299.270 1799.125 ;
        RECT 300.110 1795.720 305.710 1799.125 ;
        RECT 306.550 1795.720 308.930 1799.125 ;
        RECT 309.770 1795.720 312.150 1799.125 ;
        RECT 312.990 1795.720 315.370 1799.125 ;
        RECT 316.210 1795.720 318.590 1799.125 ;
        RECT 319.430 1795.720 321.810 1799.125 ;
        RECT 322.650 1795.720 328.250 1799.125 ;
        RECT 329.090 1795.720 331.470 1799.125 ;
        RECT 332.310 1795.720 334.690 1799.125 ;
        RECT 335.530 1795.720 337.910 1799.125 ;
        RECT 338.750 1795.720 341.130 1799.125 ;
        RECT 341.970 1795.720 344.350 1799.125 ;
        RECT 345.190 1795.720 347.570 1799.125 ;
        RECT 348.410 1795.720 354.010 1799.125 ;
        RECT 354.850 1795.720 357.230 1799.125 ;
        RECT 358.070 1795.720 360.450 1799.125 ;
        RECT 361.290 1795.720 363.670 1799.125 ;
        RECT 364.510 1795.720 366.890 1799.125 ;
        RECT 367.730 1795.720 370.110 1799.125 ;
        RECT 370.950 1795.720 376.550 1799.125 ;
        RECT 377.390 1795.720 379.770 1799.125 ;
        RECT 380.610 1795.720 382.990 1799.125 ;
        RECT 383.830 1795.720 386.210 1799.125 ;
        RECT 387.050 1795.720 389.430 1799.125 ;
        RECT 390.270 1795.720 392.650 1799.125 ;
        RECT 393.490 1795.720 395.870 1799.125 ;
        RECT 396.710 1795.720 402.310 1799.125 ;
        RECT 403.150 1795.720 405.530 1799.125 ;
        RECT 406.370 1795.720 408.750 1799.125 ;
        RECT 409.590 1795.720 411.970 1799.125 ;
        RECT 412.810 1795.720 415.190 1799.125 ;
        RECT 416.030 1795.720 418.410 1799.125 ;
        RECT 419.250 1795.720 424.850 1799.125 ;
        RECT 425.690 1795.720 428.070 1799.125 ;
        RECT 428.910 1795.720 431.290 1799.125 ;
        RECT 432.130 1795.720 434.510 1799.125 ;
        RECT 435.350 1795.720 437.730 1799.125 ;
        RECT 438.570 1795.720 440.950 1799.125 ;
        RECT 441.790 1795.720 447.390 1799.125 ;
        RECT 448.230 1795.720 450.610 1799.125 ;
        RECT 451.450 1795.720 453.830 1799.125 ;
        RECT 454.670 1795.720 457.050 1799.125 ;
        RECT 457.890 1795.720 460.270 1799.125 ;
        RECT 461.110 1795.720 463.490 1799.125 ;
        RECT 464.330 1795.720 466.710 1799.125 ;
        RECT 467.550 1795.720 473.150 1799.125 ;
        RECT 473.990 1795.720 476.370 1799.125 ;
        RECT 477.210 1795.720 479.590 1799.125 ;
        RECT 480.430 1795.720 482.810 1799.125 ;
        RECT 483.650 1795.720 486.030 1799.125 ;
        RECT 486.870 1795.720 489.250 1799.125 ;
        RECT 490.090 1795.720 495.690 1799.125 ;
        RECT 496.530 1795.720 498.910 1799.125 ;
        RECT 499.750 1795.720 502.130 1799.125 ;
        RECT 502.970 1795.720 505.350 1799.125 ;
        RECT 506.190 1795.720 508.570 1799.125 ;
        RECT 509.410 1795.720 511.790 1799.125 ;
        RECT 512.630 1795.720 515.010 1799.125 ;
        RECT 515.850 1795.720 521.450 1799.125 ;
        RECT 522.290 1795.720 524.670 1799.125 ;
        RECT 525.510 1795.720 527.890 1799.125 ;
        RECT 528.730 1795.720 531.110 1799.125 ;
        RECT 531.950 1795.720 534.330 1799.125 ;
        RECT 535.170 1795.720 537.550 1799.125 ;
        RECT 538.390 1795.720 543.990 1799.125 ;
        RECT 544.830 1795.720 547.210 1799.125 ;
        RECT 548.050 1795.720 550.430 1799.125 ;
        RECT 551.270 1795.720 553.650 1799.125 ;
        RECT 554.490 1795.720 556.870 1799.125 ;
        RECT 557.710 1795.720 560.090 1799.125 ;
        RECT 560.930 1795.720 563.310 1799.125 ;
        RECT 564.150 1795.720 569.750 1799.125 ;
        RECT 570.590 1795.720 572.970 1799.125 ;
        RECT 573.810 1795.720 576.190 1799.125 ;
        RECT 577.030 1795.720 579.410 1799.125 ;
        RECT 580.250 1795.720 582.630 1799.125 ;
        RECT 583.470 1795.720 585.850 1799.125 ;
        RECT 586.690 1795.720 592.290 1799.125 ;
        RECT 593.130 1795.720 595.510 1799.125 ;
        RECT 596.350 1795.720 598.730 1799.125 ;
        RECT 599.570 1795.720 601.950 1799.125 ;
        RECT 602.790 1795.720 605.170 1799.125 ;
        RECT 606.010 1795.720 608.390 1799.125 ;
        RECT 609.230 1795.720 614.830 1799.125 ;
        RECT 615.670 1795.720 618.050 1799.125 ;
        RECT 618.890 1795.720 621.270 1799.125 ;
        RECT 622.110 1795.720 624.490 1799.125 ;
        RECT 625.330 1795.720 627.710 1799.125 ;
        RECT 628.550 1795.720 630.930 1799.125 ;
        RECT 631.770 1795.720 634.150 1799.125 ;
        RECT 634.990 1795.720 640.590 1799.125 ;
        RECT 641.430 1795.720 643.810 1799.125 ;
        RECT 644.650 1795.720 647.030 1799.125 ;
        RECT 647.870 1795.720 650.250 1799.125 ;
        RECT 651.090 1795.720 653.470 1799.125 ;
        RECT 654.310 1795.720 656.690 1799.125 ;
        RECT 657.530 1795.720 663.130 1799.125 ;
        RECT 663.970 1795.720 666.350 1799.125 ;
        RECT 667.190 1795.720 669.570 1799.125 ;
        RECT 670.410 1795.720 672.790 1799.125 ;
        RECT 673.630 1795.720 676.010 1799.125 ;
        RECT 676.850 1795.720 679.230 1799.125 ;
        RECT 680.070 1795.720 682.450 1799.125 ;
        RECT 683.290 1795.720 688.890 1799.125 ;
        RECT 689.730 1795.720 692.110 1799.125 ;
        RECT 692.950 1795.720 695.330 1799.125 ;
        RECT 696.170 1795.720 698.550 1799.125 ;
        RECT 699.390 1795.720 701.770 1799.125 ;
        RECT 702.610 1795.720 704.990 1799.125 ;
        RECT 705.830 1795.720 711.430 1799.125 ;
        RECT 712.270 1795.720 714.650 1799.125 ;
        RECT 715.490 1795.720 717.870 1799.125 ;
        RECT 718.710 1795.720 721.090 1799.125 ;
        RECT 721.930 1795.720 724.310 1799.125 ;
        RECT 725.150 1795.720 727.530 1799.125 ;
        RECT 728.370 1795.720 730.750 1799.125 ;
        RECT 731.590 1795.720 737.190 1799.125 ;
        RECT 738.030 1795.720 740.410 1799.125 ;
        RECT 741.250 1795.720 743.630 1799.125 ;
        RECT 744.470 1795.720 746.850 1799.125 ;
        RECT 747.690 1795.720 750.070 1799.125 ;
        RECT 750.910 1795.720 753.290 1799.125 ;
        RECT 754.130 1795.720 759.730 1799.125 ;
        RECT 760.570 1795.720 762.950 1799.125 ;
        RECT 763.790 1795.720 766.170 1799.125 ;
        RECT 767.010 1795.720 769.390 1799.125 ;
        RECT 770.230 1795.720 772.610 1799.125 ;
        RECT 773.450 1795.720 775.830 1799.125 ;
        RECT 776.670 1795.720 779.050 1799.125 ;
        RECT 779.890 1795.720 785.490 1799.125 ;
        RECT 786.330 1795.720 788.710 1799.125 ;
        RECT 789.550 1795.720 791.930 1799.125 ;
        RECT 792.770 1795.720 795.150 1799.125 ;
        RECT 795.990 1795.720 798.370 1799.125 ;
        RECT 799.210 1795.720 801.590 1799.125 ;
        RECT 802.430 1795.720 808.030 1799.125 ;
        RECT 808.870 1795.720 811.250 1799.125 ;
        RECT 812.090 1795.720 814.470 1799.125 ;
        RECT 815.310 1795.720 817.690 1799.125 ;
        RECT 818.530 1795.720 820.910 1799.125 ;
        RECT 821.750 1795.720 824.130 1799.125 ;
        RECT 824.970 1795.720 830.570 1799.125 ;
        RECT 831.410 1795.720 833.790 1799.125 ;
        RECT 834.630 1795.720 837.010 1799.125 ;
        RECT 837.850 1795.720 840.230 1799.125 ;
        RECT 841.070 1795.720 843.450 1799.125 ;
        RECT 844.290 1795.720 846.670 1799.125 ;
        RECT 847.510 1795.720 849.890 1799.125 ;
        RECT 850.730 1795.720 856.330 1799.125 ;
        RECT 857.170 1795.720 859.550 1799.125 ;
        RECT 860.390 1795.720 862.770 1799.125 ;
        RECT 863.610 1795.720 865.990 1799.125 ;
        RECT 866.830 1795.720 869.210 1799.125 ;
        RECT 870.050 1795.720 872.430 1799.125 ;
        RECT 873.270 1795.720 878.870 1799.125 ;
        RECT 879.710 1795.720 882.090 1799.125 ;
        RECT 882.930 1795.720 885.310 1799.125 ;
        RECT 886.150 1795.720 888.530 1799.125 ;
        RECT 889.370 1795.720 891.750 1799.125 ;
        RECT 892.590 1795.720 894.970 1799.125 ;
        RECT 895.810 1795.720 898.190 1799.125 ;
        RECT 899.030 1795.720 904.630 1799.125 ;
        RECT 905.470 1795.720 907.850 1799.125 ;
        RECT 908.690 1795.720 911.070 1799.125 ;
        RECT 911.910 1795.720 914.290 1799.125 ;
        RECT 915.130 1795.720 917.510 1799.125 ;
        RECT 918.350 1795.720 920.730 1799.125 ;
        RECT 921.570 1795.720 927.170 1799.125 ;
        RECT 928.010 1795.720 930.390 1799.125 ;
        RECT 931.230 1795.720 933.610 1799.125 ;
        RECT 934.450 1795.720 936.830 1799.125 ;
        RECT 937.670 1795.720 940.050 1799.125 ;
        RECT 940.890 1795.720 943.270 1799.125 ;
        RECT 944.110 1795.720 946.490 1799.125 ;
        RECT 947.330 1795.720 952.930 1799.125 ;
        RECT 953.770 1795.720 956.150 1799.125 ;
        RECT 956.990 1795.720 959.370 1799.125 ;
        RECT 960.210 1795.720 962.590 1799.125 ;
        RECT 963.430 1795.720 965.810 1799.125 ;
        RECT 966.650 1795.720 969.030 1799.125 ;
        RECT 969.870 1795.720 975.470 1799.125 ;
        RECT 976.310 1795.720 978.690 1799.125 ;
        RECT 979.530 1795.720 981.910 1799.125 ;
        RECT 982.750 1795.720 985.130 1799.125 ;
        RECT 985.970 1795.720 988.350 1799.125 ;
        RECT 989.190 1795.720 991.570 1799.125 ;
        RECT 992.410 1795.720 998.010 1799.125 ;
        RECT 998.850 1795.720 1001.230 1799.125 ;
        RECT 1002.070 1795.720 1004.450 1799.125 ;
        RECT 1005.290 1795.720 1007.670 1799.125 ;
        RECT 1008.510 1795.720 1010.890 1799.125 ;
        RECT 1011.730 1795.720 1014.110 1799.125 ;
        RECT 1014.950 1795.720 1017.330 1799.125 ;
        RECT 1018.170 1795.720 1023.770 1799.125 ;
        RECT 1024.610 1795.720 1026.990 1799.125 ;
        RECT 1027.830 1795.720 1030.210 1799.125 ;
        RECT 1031.050 1795.720 1033.430 1799.125 ;
        RECT 1034.270 1795.720 1036.650 1799.125 ;
        RECT 1037.490 1795.720 1039.870 1799.125 ;
        RECT 1040.710 1795.720 1046.310 1799.125 ;
        RECT 1047.150 1795.720 1049.530 1799.125 ;
        RECT 1050.370 1795.720 1052.750 1799.125 ;
        RECT 1053.590 1795.720 1055.970 1799.125 ;
        RECT 1056.810 1795.720 1059.190 1799.125 ;
        RECT 1060.030 1795.720 1062.410 1799.125 ;
        RECT 1063.250 1795.720 1065.630 1799.125 ;
        RECT 1066.470 1795.720 1072.070 1799.125 ;
        RECT 1072.910 1795.720 1075.290 1799.125 ;
        RECT 1076.130 1795.720 1078.510 1799.125 ;
        RECT 1079.350 1795.720 1081.730 1799.125 ;
        RECT 1082.570 1795.720 1084.950 1799.125 ;
        RECT 1085.790 1795.720 1088.170 1799.125 ;
        RECT 1089.010 1795.720 1094.610 1799.125 ;
        RECT 1095.450 1795.720 1097.830 1799.125 ;
        RECT 1098.670 1795.720 1101.050 1799.125 ;
        RECT 1101.890 1795.720 1104.270 1799.125 ;
        RECT 1105.110 1795.720 1107.490 1799.125 ;
        RECT 1108.330 1795.720 1110.710 1799.125 ;
        RECT 1111.550 1795.720 1113.930 1799.125 ;
        RECT 1114.770 1795.720 1120.370 1799.125 ;
        RECT 1121.210 1795.720 1123.590 1799.125 ;
        RECT 1124.430 1795.720 1126.810 1799.125 ;
        RECT 1127.650 1795.720 1130.030 1799.125 ;
        RECT 1130.870 1795.720 1133.250 1799.125 ;
        RECT 1134.090 1795.720 1136.470 1799.125 ;
        RECT 1137.310 1795.720 1142.910 1799.125 ;
        RECT 1143.750 1795.720 1146.130 1799.125 ;
        RECT 1146.970 1795.720 1149.350 1799.125 ;
        RECT 1150.190 1795.720 1152.570 1799.125 ;
        RECT 1153.410 1795.720 1155.790 1799.125 ;
        RECT 1156.630 1795.720 1159.010 1799.125 ;
        RECT 1159.850 1795.720 1165.450 1799.125 ;
        RECT 1166.290 1795.720 1168.670 1799.125 ;
        RECT 1169.510 1795.720 1171.890 1799.125 ;
        RECT 1172.730 1795.720 1175.110 1799.125 ;
        RECT 1175.950 1795.720 1178.330 1799.125 ;
        RECT 1179.170 1795.720 1181.550 1799.125 ;
        RECT 1182.390 1795.720 1184.770 1799.125 ;
        RECT 1185.610 1795.720 1191.210 1799.125 ;
        RECT 1192.050 1795.720 1194.430 1799.125 ;
        RECT 1195.270 1795.720 1197.650 1799.125 ;
        RECT 1198.490 1795.720 1200.870 1799.125 ;
        RECT 1201.710 1795.720 1204.090 1799.125 ;
        RECT 1204.930 1795.720 1207.310 1799.125 ;
        RECT 1208.150 1795.720 1213.750 1799.125 ;
        RECT 1214.590 1795.720 1216.970 1799.125 ;
        RECT 1217.810 1795.720 1220.190 1799.125 ;
        RECT 1221.030 1795.720 1223.410 1799.125 ;
        RECT 1224.250 1795.720 1226.630 1799.125 ;
        RECT 1227.470 1795.720 1229.850 1799.125 ;
        RECT 1230.690 1795.720 1233.070 1799.125 ;
        RECT 1233.910 1795.720 1239.510 1799.125 ;
        RECT 1240.350 1795.720 1242.730 1799.125 ;
        RECT 1243.570 1795.720 1245.950 1799.125 ;
        RECT 1246.790 1795.720 1249.170 1799.125 ;
        RECT 1250.010 1795.720 1252.390 1799.125 ;
        RECT 1253.230 1795.720 1255.610 1799.125 ;
        RECT 1256.450 1795.720 1262.050 1799.125 ;
        RECT 1262.890 1795.720 1265.270 1799.125 ;
        RECT 1266.110 1795.720 1268.490 1799.125 ;
        RECT 1269.330 1795.720 1271.710 1799.125 ;
        RECT 1272.550 1795.720 1274.930 1799.125 ;
        RECT 1275.770 1795.720 1278.150 1799.125 ;
        RECT 1278.990 1795.720 1281.370 1799.125 ;
        RECT 1282.210 1795.720 1287.810 1799.125 ;
        RECT 1288.650 1795.720 1291.030 1799.125 ;
        RECT 1291.870 1795.720 1294.250 1799.125 ;
        RECT 1295.090 1795.720 1297.470 1799.125 ;
        RECT 1298.310 1795.720 1300.690 1799.125 ;
        RECT 1301.530 1795.720 1303.910 1799.125 ;
        RECT 1304.750 1795.720 1310.350 1799.125 ;
        RECT 1311.190 1795.720 1313.570 1799.125 ;
        RECT 1314.410 1795.720 1316.790 1799.125 ;
        RECT 1317.630 1795.720 1320.010 1799.125 ;
        RECT 1320.850 1795.720 1323.230 1799.125 ;
        RECT 1324.070 1795.720 1326.450 1799.125 ;
        RECT 1327.290 1795.720 1332.890 1799.125 ;
        RECT 1333.730 1795.720 1336.110 1799.125 ;
        RECT 1336.950 1795.720 1339.330 1799.125 ;
        RECT 1340.170 1795.720 1342.550 1799.125 ;
        RECT 1343.390 1795.720 1345.770 1799.125 ;
        RECT 1346.610 1795.720 1348.990 1799.125 ;
        RECT 1349.830 1795.720 1352.210 1799.125 ;
        RECT 1353.050 1795.720 1358.650 1799.125 ;
        RECT 1359.490 1795.720 1361.870 1799.125 ;
        RECT 1362.710 1795.720 1365.090 1799.125 ;
        RECT 1365.930 1795.720 1368.310 1799.125 ;
        RECT 1369.150 1795.720 1371.530 1799.125 ;
        RECT 1372.370 1795.720 1374.750 1799.125 ;
        RECT 1375.590 1795.720 1381.190 1799.125 ;
        RECT 1382.030 1795.720 1384.410 1799.125 ;
        RECT 1385.250 1795.720 1387.630 1799.125 ;
        RECT 1388.470 1795.720 1390.850 1799.125 ;
        RECT 1391.690 1795.720 1394.070 1799.125 ;
        RECT 1394.910 1795.720 1397.290 1799.125 ;
        RECT 1398.130 1795.720 1400.510 1799.125 ;
        RECT 1401.350 1795.720 1406.950 1799.125 ;
        RECT 1407.790 1795.720 1410.170 1799.125 ;
        RECT 1411.010 1795.720 1413.390 1799.125 ;
        RECT 1414.230 1795.720 1416.610 1799.125 ;
        RECT 1417.450 1795.720 1419.830 1799.125 ;
        RECT 1420.670 1795.720 1423.050 1799.125 ;
        RECT 1423.890 1795.720 1429.490 1799.125 ;
        RECT 1430.330 1795.720 1432.710 1799.125 ;
        RECT 1433.550 1795.720 1435.930 1799.125 ;
        RECT 1436.770 1795.720 1439.150 1799.125 ;
        RECT 1439.990 1795.720 1442.370 1799.125 ;
        RECT 1443.210 1795.720 1445.590 1799.125 ;
        RECT 1446.430 1795.720 1448.810 1799.125 ;
        RECT 1449.650 1795.720 1455.250 1799.125 ;
        RECT 1456.090 1795.720 1458.470 1799.125 ;
        RECT 1459.310 1795.720 1461.690 1799.125 ;
        RECT 1462.530 1795.720 1464.910 1799.125 ;
        RECT 1465.750 1795.720 1468.130 1799.125 ;
        RECT 1468.970 1795.720 1471.350 1799.125 ;
        RECT 1472.190 1795.720 1477.790 1799.125 ;
        RECT 1478.630 1795.720 1481.010 1799.125 ;
        RECT 1481.850 1795.720 1484.230 1799.125 ;
        RECT 1485.070 1795.720 1487.450 1799.125 ;
        RECT 1488.290 1795.720 1490.670 1799.125 ;
        RECT 1491.510 1795.720 1493.890 1799.125 ;
        RECT 1494.730 1795.720 1497.110 1799.125 ;
        RECT 1497.950 1795.720 1498.120 1799.125 ;
        RECT 0.100 4.280 1498.120 1795.720 ;
        RECT 0.650 0.155 3.030 4.280 ;
        RECT 3.870 0.155 6.250 4.280 ;
        RECT 7.090 0.155 9.470 4.280 ;
        RECT 10.310 0.155 12.690 4.280 ;
        RECT 13.530 0.155 15.910 4.280 ;
        RECT 16.750 0.155 19.130 4.280 ;
        RECT 19.970 0.155 25.570 4.280 ;
        RECT 26.410 0.155 28.790 4.280 ;
        RECT 29.630 0.155 32.010 4.280 ;
        RECT 32.850 0.155 35.230 4.280 ;
        RECT 36.070 0.155 38.450 4.280 ;
        RECT 39.290 0.155 41.670 4.280 ;
        RECT 42.510 0.155 48.110 4.280 ;
        RECT 48.950 0.155 51.330 4.280 ;
        RECT 52.170 0.155 54.550 4.280 ;
        RECT 55.390 0.155 57.770 4.280 ;
        RECT 58.610 0.155 60.990 4.280 ;
        RECT 61.830 0.155 64.210 4.280 ;
        RECT 65.050 0.155 67.430 4.280 ;
        RECT 68.270 0.155 73.870 4.280 ;
        RECT 74.710 0.155 77.090 4.280 ;
        RECT 77.930 0.155 80.310 4.280 ;
        RECT 81.150 0.155 83.530 4.280 ;
        RECT 84.370 0.155 86.750 4.280 ;
        RECT 87.590 0.155 89.970 4.280 ;
        RECT 90.810 0.155 96.410 4.280 ;
        RECT 97.250 0.155 99.630 4.280 ;
        RECT 100.470 0.155 102.850 4.280 ;
        RECT 103.690 0.155 106.070 4.280 ;
        RECT 106.910 0.155 109.290 4.280 ;
        RECT 110.130 0.155 112.510 4.280 ;
        RECT 113.350 0.155 115.730 4.280 ;
        RECT 116.570 0.155 122.170 4.280 ;
        RECT 123.010 0.155 125.390 4.280 ;
        RECT 126.230 0.155 128.610 4.280 ;
        RECT 129.450 0.155 131.830 4.280 ;
        RECT 132.670 0.155 135.050 4.280 ;
        RECT 135.890 0.155 138.270 4.280 ;
        RECT 139.110 0.155 144.710 4.280 ;
        RECT 145.550 0.155 147.930 4.280 ;
        RECT 148.770 0.155 151.150 4.280 ;
        RECT 151.990 0.155 154.370 4.280 ;
        RECT 155.210 0.155 157.590 4.280 ;
        RECT 158.430 0.155 160.810 4.280 ;
        RECT 161.650 0.155 164.030 4.280 ;
        RECT 164.870 0.155 170.470 4.280 ;
        RECT 171.310 0.155 173.690 4.280 ;
        RECT 174.530 0.155 176.910 4.280 ;
        RECT 177.750 0.155 180.130 4.280 ;
        RECT 180.970 0.155 183.350 4.280 ;
        RECT 184.190 0.155 186.570 4.280 ;
        RECT 187.410 0.155 193.010 4.280 ;
        RECT 193.850 0.155 196.230 4.280 ;
        RECT 197.070 0.155 199.450 4.280 ;
        RECT 200.290 0.155 202.670 4.280 ;
        RECT 203.510 0.155 205.890 4.280 ;
        RECT 206.730 0.155 209.110 4.280 ;
        RECT 209.950 0.155 215.550 4.280 ;
        RECT 216.390 0.155 218.770 4.280 ;
        RECT 219.610 0.155 221.990 4.280 ;
        RECT 222.830 0.155 225.210 4.280 ;
        RECT 226.050 0.155 228.430 4.280 ;
        RECT 229.270 0.155 231.650 4.280 ;
        RECT 232.490 0.155 234.870 4.280 ;
        RECT 235.710 0.155 241.310 4.280 ;
        RECT 242.150 0.155 244.530 4.280 ;
        RECT 245.370 0.155 247.750 4.280 ;
        RECT 248.590 0.155 250.970 4.280 ;
        RECT 251.810 0.155 254.190 4.280 ;
        RECT 255.030 0.155 257.410 4.280 ;
        RECT 258.250 0.155 263.850 4.280 ;
        RECT 264.690 0.155 267.070 4.280 ;
        RECT 267.910 0.155 270.290 4.280 ;
        RECT 271.130 0.155 273.510 4.280 ;
        RECT 274.350 0.155 276.730 4.280 ;
        RECT 277.570 0.155 279.950 4.280 ;
        RECT 280.790 0.155 283.170 4.280 ;
        RECT 284.010 0.155 289.610 4.280 ;
        RECT 290.450 0.155 292.830 4.280 ;
        RECT 293.670 0.155 296.050 4.280 ;
        RECT 296.890 0.155 299.270 4.280 ;
        RECT 300.110 0.155 302.490 4.280 ;
        RECT 303.330 0.155 305.710 4.280 ;
        RECT 306.550 0.155 312.150 4.280 ;
        RECT 312.990 0.155 315.370 4.280 ;
        RECT 316.210 0.155 318.590 4.280 ;
        RECT 319.430 0.155 321.810 4.280 ;
        RECT 322.650 0.155 325.030 4.280 ;
        RECT 325.870 0.155 328.250 4.280 ;
        RECT 329.090 0.155 331.470 4.280 ;
        RECT 332.310 0.155 337.910 4.280 ;
        RECT 338.750 0.155 341.130 4.280 ;
        RECT 341.970 0.155 344.350 4.280 ;
        RECT 345.190 0.155 347.570 4.280 ;
        RECT 348.410 0.155 350.790 4.280 ;
        RECT 351.630 0.155 354.010 4.280 ;
        RECT 354.850 0.155 360.450 4.280 ;
        RECT 361.290 0.155 363.670 4.280 ;
        RECT 364.510 0.155 366.890 4.280 ;
        RECT 367.730 0.155 370.110 4.280 ;
        RECT 370.950 0.155 373.330 4.280 ;
        RECT 374.170 0.155 376.550 4.280 ;
        RECT 377.390 0.155 382.990 4.280 ;
        RECT 383.830 0.155 386.210 4.280 ;
        RECT 387.050 0.155 389.430 4.280 ;
        RECT 390.270 0.155 392.650 4.280 ;
        RECT 393.490 0.155 395.870 4.280 ;
        RECT 396.710 0.155 399.090 4.280 ;
        RECT 399.930 0.155 402.310 4.280 ;
        RECT 403.150 0.155 408.750 4.280 ;
        RECT 409.590 0.155 411.970 4.280 ;
        RECT 412.810 0.155 415.190 4.280 ;
        RECT 416.030 0.155 418.410 4.280 ;
        RECT 419.250 0.155 421.630 4.280 ;
        RECT 422.470 0.155 424.850 4.280 ;
        RECT 425.690 0.155 431.290 4.280 ;
        RECT 432.130 0.155 434.510 4.280 ;
        RECT 435.350 0.155 437.730 4.280 ;
        RECT 438.570 0.155 440.950 4.280 ;
        RECT 441.790 0.155 444.170 4.280 ;
        RECT 445.010 0.155 447.390 4.280 ;
        RECT 448.230 0.155 450.610 4.280 ;
        RECT 451.450 0.155 457.050 4.280 ;
        RECT 457.890 0.155 460.270 4.280 ;
        RECT 461.110 0.155 463.490 4.280 ;
        RECT 464.330 0.155 466.710 4.280 ;
        RECT 467.550 0.155 469.930 4.280 ;
        RECT 470.770 0.155 473.150 4.280 ;
        RECT 473.990 0.155 479.590 4.280 ;
        RECT 480.430 0.155 482.810 4.280 ;
        RECT 483.650 0.155 486.030 4.280 ;
        RECT 486.870 0.155 489.250 4.280 ;
        RECT 490.090 0.155 492.470 4.280 ;
        RECT 493.310 0.155 495.690 4.280 ;
        RECT 496.530 0.155 498.910 4.280 ;
        RECT 499.750 0.155 505.350 4.280 ;
        RECT 506.190 0.155 508.570 4.280 ;
        RECT 509.410 0.155 511.790 4.280 ;
        RECT 512.630 0.155 515.010 4.280 ;
        RECT 515.850 0.155 518.230 4.280 ;
        RECT 519.070 0.155 521.450 4.280 ;
        RECT 522.290 0.155 527.890 4.280 ;
        RECT 528.730 0.155 531.110 4.280 ;
        RECT 531.950 0.155 534.330 4.280 ;
        RECT 535.170 0.155 537.550 4.280 ;
        RECT 538.390 0.155 540.770 4.280 ;
        RECT 541.610 0.155 543.990 4.280 ;
        RECT 544.830 0.155 550.430 4.280 ;
        RECT 551.270 0.155 553.650 4.280 ;
        RECT 554.490 0.155 556.870 4.280 ;
        RECT 557.710 0.155 560.090 4.280 ;
        RECT 560.930 0.155 563.310 4.280 ;
        RECT 564.150 0.155 566.530 4.280 ;
        RECT 567.370 0.155 569.750 4.280 ;
        RECT 570.590 0.155 576.190 4.280 ;
        RECT 577.030 0.155 579.410 4.280 ;
        RECT 580.250 0.155 582.630 4.280 ;
        RECT 583.470 0.155 585.850 4.280 ;
        RECT 586.690 0.155 589.070 4.280 ;
        RECT 589.910 0.155 592.290 4.280 ;
        RECT 593.130 0.155 598.730 4.280 ;
        RECT 599.570 0.155 601.950 4.280 ;
        RECT 602.790 0.155 605.170 4.280 ;
        RECT 606.010 0.155 608.390 4.280 ;
        RECT 609.230 0.155 611.610 4.280 ;
        RECT 612.450 0.155 614.830 4.280 ;
        RECT 615.670 0.155 618.050 4.280 ;
        RECT 618.890 0.155 624.490 4.280 ;
        RECT 625.330 0.155 627.710 4.280 ;
        RECT 628.550 0.155 630.930 4.280 ;
        RECT 631.770 0.155 634.150 4.280 ;
        RECT 634.990 0.155 637.370 4.280 ;
        RECT 638.210 0.155 640.590 4.280 ;
        RECT 641.430 0.155 647.030 4.280 ;
        RECT 647.870 0.155 650.250 4.280 ;
        RECT 651.090 0.155 653.470 4.280 ;
        RECT 654.310 0.155 656.690 4.280 ;
        RECT 657.530 0.155 659.910 4.280 ;
        RECT 660.750 0.155 663.130 4.280 ;
        RECT 663.970 0.155 666.350 4.280 ;
        RECT 667.190 0.155 672.790 4.280 ;
        RECT 673.630 0.155 676.010 4.280 ;
        RECT 676.850 0.155 679.230 4.280 ;
        RECT 680.070 0.155 682.450 4.280 ;
        RECT 683.290 0.155 685.670 4.280 ;
        RECT 686.510 0.155 688.890 4.280 ;
        RECT 689.730 0.155 695.330 4.280 ;
        RECT 696.170 0.155 698.550 4.280 ;
        RECT 699.390 0.155 701.770 4.280 ;
        RECT 702.610 0.155 704.990 4.280 ;
        RECT 705.830 0.155 708.210 4.280 ;
        RECT 709.050 0.155 711.430 4.280 ;
        RECT 712.270 0.155 717.870 4.280 ;
        RECT 718.710 0.155 721.090 4.280 ;
        RECT 721.930 0.155 724.310 4.280 ;
        RECT 725.150 0.155 727.530 4.280 ;
        RECT 728.370 0.155 730.750 4.280 ;
        RECT 731.590 0.155 733.970 4.280 ;
        RECT 734.810 0.155 737.190 4.280 ;
        RECT 738.030 0.155 743.630 4.280 ;
        RECT 744.470 0.155 746.850 4.280 ;
        RECT 747.690 0.155 750.070 4.280 ;
        RECT 750.910 0.155 753.290 4.280 ;
        RECT 754.130 0.155 756.510 4.280 ;
        RECT 757.350 0.155 759.730 4.280 ;
        RECT 760.570 0.155 766.170 4.280 ;
        RECT 767.010 0.155 769.390 4.280 ;
        RECT 770.230 0.155 772.610 4.280 ;
        RECT 773.450 0.155 775.830 4.280 ;
        RECT 776.670 0.155 779.050 4.280 ;
        RECT 779.890 0.155 782.270 4.280 ;
        RECT 783.110 0.155 785.490 4.280 ;
        RECT 786.330 0.155 791.930 4.280 ;
        RECT 792.770 0.155 795.150 4.280 ;
        RECT 795.990 0.155 798.370 4.280 ;
        RECT 799.210 0.155 801.590 4.280 ;
        RECT 802.430 0.155 804.810 4.280 ;
        RECT 805.650 0.155 808.030 4.280 ;
        RECT 808.870 0.155 814.470 4.280 ;
        RECT 815.310 0.155 817.690 4.280 ;
        RECT 818.530 0.155 820.910 4.280 ;
        RECT 821.750 0.155 824.130 4.280 ;
        RECT 824.970 0.155 827.350 4.280 ;
        RECT 828.190 0.155 830.570 4.280 ;
        RECT 831.410 0.155 833.790 4.280 ;
        RECT 834.630 0.155 840.230 4.280 ;
        RECT 841.070 0.155 843.450 4.280 ;
        RECT 844.290 0.155 846.670 4.280 ;
        RECT 847.510 0.155 849.890 4.280 ;
        RECT 850.730 0.155 853.110 4.280 ;
        RECT 853.950 0.155 856.330 4.280 ;
        RECT 857.170 0.155 862.770 4.280 ;
        RECT 863.610 0.155 865.990 4.280 ;
        RECT 866.830 0.155 869.210 4.280 ;
        RECT 870.050 0.155 872.430 4.280 ;
        RECT 873.270 0.155 875.650 4.280 ;
        RECT 876.490 0.155 878.870 4.280 ;
        RECT 879.710 0.155 882.090 4.280 ;
        RECT 882.930 0.155 888.530 4.280 ;
        RECT 889.370 0.155 891.750 4.280 ;
        RECT 892.590 0.155 894.970 4.280 ;
        RECT 895.810 0.155 898.190 4.280 ;
        RECT 899.030 0.155 901.410 4.280 ;
        RECT 902.250 0.155 904.630 4.280 ;
        RECT 905.470 0.155 911.070 4.280 ;
        RECT 911.910 0.155 914.290 4.280 ;
        RECT 915.130 0.155 917.510 4.280 ;
        RECT 918.350 0.155 920.730 4.280 ;
        RECT 921.570 0.155 923.950 4.280 ;
        RECT 924.790 0.155 927.170 4.280 ;
        RECT 928.010 0.155 933.610 4.280 ;
        RECT 934.450 0.155 936.830 4.280 ;
        RECT 937.670 0.155 940.050 4.280 ;
        RECT 940.890 0.155 943.270 4.280 ;
        RECT 944.110 0.155 946.490 4.280 ;
        RECT 947.330 0.155 949.710 4.280 ;
        RECT 950.550 0.155 952.930 4.280 ;
        RECT 953.770 0.155 959.370 4.280 ;
        RECT 960.210 0.155 962.590 4.280 ;
        RECT 963.430 0.155 965.810 4.280 ;
        RECT 966.650 0.155 969.030 4.280 ;
        RECT 969.870 0.155 972.250 4.280 ;
        RECT 973.090 0.155 975.470 4.280 ;
        RECT 976.310 0.155 981.910 4.280 ;
        RECT 982.750 0.155 985.130 4.280 ;
        RECT 985.970 0.155 988.350 4.280 ;
        RECT 989.190 0.155 991.570 4.280 ;
        RECT 992.410 0.155 994.790 4.280 ;
        RECT 995.630 0.155 998.010 4.280 ;
        RECT 998.850 0.155 1001.230 4.280 ;
        RECT 1002.070 0.155 1007.670 4.280 ;
        RECT 1008.510 0.155 1010.890 4.280 ;
        RECT 1011.730 0.155 1014.110 4.280 ;
        RECT 1014.950 0.155 1017.330 4.280 ;
        RECT 1018.170 0.155 1020.550 4.280 ;
        RECT 1021.390 0.155 1023.770 4.280 ;
        RECT 1024.610 0.155 1030.210 4.280 ;
        RECT 1031.050 0.155 1033.430 4.280 ;
        RECT 1034.270 0.155 1036.650 4.280 ;
        RECT 1037.490 0.155 1039.870 4.280 ;
        RECT 1040.710 0.155 1043.090 4.280 ;
        RECT 1043.930 0.155 1046.310 4.280 ;
        RECT 1047.150 0.155 1049.530 4.280 ;
        RECT 1050.370 0.155 1055.970 4.280 ;
        RECT 1056.810 0.155 1059.190 4.280 ;
        RECT 1060.030 0.155 1062.410 4.280 ;
        RECT 1063.250 0.155 1065.630 4.280 ;
        RECT 1066.470 0.155 1068.850 4.280 ;
        RECT 1069.690 0.155 1072.070 4.280 ;
        RECT 1072.910 0.155 1078.510 4.280 ;
        RECT 1079.350 0.155 1081.730 4.280 ;
        RECT 1082.570 0.155 1084.950 4.280 ;
        RECT 1085.790 0.155 1088.170 4.280 ;
        RECT 1089.010 0.155 1091.390 4.280 ;
        RECT 1092.230 0.155 1094.610 4.280 ;
        RECT 1095.450 0.155 1101.050 4.280 ;
        RECT 1101.890 0.155 1104.270 4.280 ;
        RECT 1105.110 0.155 1107.490 4.280 ;
        RECT 1108.330 0.155 1110.710 4.280 ;
        RECT 1111.550 0.155 1113.930 4.280 ;
        RECT 1114.770 0.155 1117.150 4.280 ;
        RECT 1117.990 0.155 1120.370 4.280 ;
        RECT 1121.210 0.155 1126.810 4.280 ;
        RECT 1127.650 0.155 1130.030 4.280 ;
        RECT 1130.870 0.155 1133.250 4.280 ;
        RECT 1134.090 0.155 1136.470 4.280 ;
        RECT 1137.310 0.155 1139.690 4.280 ;
        RECT 1140.530 0.155 1142.910 4.280 ;
        RECT 1143.750 0.155 1149.350 4.280 ;
        RECT 1150.190 0.155 1152.570 4.280 ;
        RECT 1153.410 0.155 1155.790 4.280 ;
        RECT 1156.630 0.155 1159.010 4.280 ;
        RECT 1159.850 0.155 1162.230 4.280 ;
        RECT 1163.070 0.155 1165.450 4.280 ;
        RECT 1166.290 0.155 1168.670 4.280 ;
        RECT 1169.510 0.155 1175.110 4.280 ;
        RECT 1175.950 0.155 1178.330 4.280 ;
        RECT 1179.170 0.155 1181.550 4.280 ;
        RECT 1182.390 0.155 1184.770 4.280 ;
        RECT 1185.610 0.155 1187.990 4.280 ;
        RECT 1188.830 0.155 1191.210 4.280 ;
        RECT 1192.050 0.155 1197.650 4.280 ;
        RECT 1198.490 0.155 1200.870 4.280 ;
        RECT 1201.710 0.155 1204.090 4.280 ;
        RECT 1204.930 0.155 1207.310 4.280 ;
        RECT 1208.150 0.155 1210.530 4.280 ;
        RECT 1211.370 0.155 1213.750 4.280 ;
        RECT 1214.590 0.155 1216.970 4.280 ;
        RECT 1217.810 0.155 1223.410 4.280 ;
        RECT 1224.250 0.155 1226.630 4.280 ;
        RECT 1227.470 0.155 1229.850 4.280 ;
        RECT 1230.690 0.155 1233.070 4.280 ;
        RECT 1233.910 0.155 1236.290 4.280 ;
        RECT 1237.130 0.155 1239.510 4.280 ;
        RECT 1240.350 0.155 1245.950 4.280 ;
        RECT 1246.790 0.155 1249.170 4.280 ;
        RECT 1250.010 0.155 1252.390 4.280 ;
        RECT 1253.230 0.155 1255.610 4.280 ;
        RECT 1256.450 0.155 1258.830 4.280 ;
        RECT 1259.670 0.155 1262.050 4.280 ;
        RECT 1262.890 0.155 1268.490 4.280 ;
        RECT 1269.330 0.155 1271.710 4.280 ;
        RECT 1272.550 0.155 1274.930 4.280 ;
        RECT 1275.770 0.155 1278.150 4.280 ;
        RECT 1278.990 0.155 1281.370 4.280 ;
        RECT 1282.210 0.155 1284.590 4.280 ;
        RECT 1285.430 0.155 1287.810 4.280 ;
        RECT 1288.650 0.155 1294.250 4.280 ;
        RECT 1295.090 0.155 1297.470 4.280 ;
        RECT 1298.310 0.155 1300.690 4.280 ;
        RECT 1301.530 0.155 1303.910 4.280 ;
        RECT 1304.750 0.155 1307.130 4.280 ;
        RECT 1307.970 0.155 1310.350 4.280 ;
        RECT 1311.190 0.155 1316.790 4.280 ;
        RECT 1317.630 0.155 1320.010 4.280 ;
        RECT 1320.850 0.155 1323.230 4.280 ;
        RECT 1324.070 0.155 1326.450 4.280 ;
        RECT 1327.290 0.155 1329.670 4.280 ;
        RECT 1330.510 0.155 1332.890 4.280 ;
        RECT 1333.730 0.155 1336.110 4.280 ;
        RECT 1336.950 0.155 1342.550 4.280 ;
        RECT 1343.390 0.155 1345.770 4.280 ;
        RECT 1346.610 0.155 1348.990 4.280 ;
        RECT 1349.830 0.155 1352.210 4.280 ;
        RECT 1353.050 0.155 1355.430 4.280 ;
        RECT 1356.270 0.155 1358.650 4.280 ;
        RECT 1359.490 0.155 1365.090 4.280 ;
        RECT 1365.930 0.155 1368.310 4.280 ;
        RECT 1369.150 0.155 1371.530 4.280 ;
        RECT 1372.370 0.155 1374.750 4.280 ;
        RECT 1375.590 0.155 1377.970 4.280 ;
        RECT 1378.810 0.155 1381.190 4.280 ;
        RECT 1382.030 0.155 1384.410 4.280 ;
        RECT 1385.250 0.155 1390.850 4.280 ;
        RECT 1391.690 0.155 1394.070 4.280 ;
        RECT 1394.910 0.155 1397.290 4.280 ;
        RECT 1398.130 0.155 1400.510 4.280 ;
        RECT 1401.350 0.155 1403.730 4.280 ;
        RECT 1404.570 0.155 1406.950 4.280 ;
        RECT 1407.790 0.155 1413.390 4.280 ;
        RECT 1414.230 0.155 1416.610 4.280 ;
        RECT 1417.450 0.155 1419.830 4.280 ;
        RECT 1420.670 0.155 1423.050 4.280 ;
        RECT 1423.890 0.155 1426.270 4.280 ;
        RECT 1427.110 0.155 1429.490 4.280 ;
        RECT 1430.330 0.155 1435.930 4.280 ;
        RECT 1436.770 0.155 1439.150 4.280 ;
        RECT 1439.990 0.155 1442.370 4.280 ;
        RECT 1443.210 0.155 1445.590 4.280 ;
        RECT 1446.430 0.155 1448.810 4.280 ;
        RECT 1449.650 0.155 1452.030 4.280 ;
        RECT 1452.870 0.155 1455.250 4.280 ;
        RECT 1456.090 0.155 1461.690 4.280 ;
        RECT 1462.530 0.155 1464.910 4.280 ;
        RECT 1465.750 0.155 1468.130 4.280 ;
        RECT 1468.970 0.155 1471.350 4.280 ;
        RECT 1472.190 0.155 1474.570 4.280 ;
        RECT 1475.410 0.155 1477.790 4.280 ;
        RECT 1478.630 0.155 1484.230 4.280 ;
        RECT 1485.070 0.155 1487.450 4.280 ;
        RECT 1488.290 0.155 1490.670 4.280 ;
        RECT 1491.510 0.155 1493.890 4.280 ;
        RECT 1494.730 0.155 1497.110 4.280 ;
        RECT 1497.950 0.155 1498.120 4.280 ;
      LAYER met3 ;
        RECT 4.400 1798.240 1497.695 1799.105 ;
        RECT 2.365 1796.240 1497.695 1798.240 ;
        RECT 4.400 1794.840 1495.600 1796.240 ;
        RECT 2.365 1792.840 1497.695 1794.840 ;
        RECT 2.365 1791.440 1495.600 1792.840 ;
        RECT 2.365 1789.440 1497.695 1791.440 ;
        RECT 4.400 1788.040 1495.600 1789.440 ;
        RECT 2.365 1786.040 1497.695 1788.040 ;
        RECT 4.400 1784.640 1495.600 1786.040 ;
        RECT 2.365 1782.640 1497.695 1784.640 ;
        RECT 4.400 1781.240 1495.600 1782.640 ;
        RECT 2.365 1779.240 1497.695 1781.240 ;
        RECT 4.400 1777.840 1495.600 1779.240 ;
        RECT 2.365 1775.840 1497.695 1777.840 ;
        RECT 4.400 1774.440 1497.695 1775.840 ;
        RECT 2.365 1772.440 1497.695 1774.440 ;
        RECT 4.400 1771.040 1495.600 1772.440 ;
        RECT 2.365 1769.040 1497.695 1771.040 ;
        RECT 2.365 1767.640 1495.600 1769.040 ;
        RECT 2.365 1765.640 1497.695 1767.640 ;
        RECT 4.400 1764.240 1495.600 1765.640 ;
        RECT 2.365 1762.240 1497.695 1764.240 ;
        RECT 4.400 1760.840 1495.600 1762.240 ;
        RECT 2.365 1758.840 1497.695 1760.840 ;
        RECT 4.400 1757.440 1495.600 1758.840 ;
        RECT 2.365 1755.440 1497.695 1757.440 ;
        RECT 4.400 1754.040 1495.600 1755.440 ;
        RECT 2.365 1752.040 1497.695 1754.040 ;
        RECT 4.400 1750.640 1497.695 1752.040 ;
        RECT 2.365 1748.640 1497.695 1750.640 ;
        RECT 4.400 1747.240 1495.600 1748.640 ;
        RECT 2.365 1745.240 1497.695 1747.240 ;
        RECT 4.400 1743.840 1495.600 1745.240 ;
        RECT 2.365 1741.840 1497.695 1743.840 ;
        RECT 2.365 1740.440 1495.600 1741.840 ;
        RECT 2.365 1738.440 1497.695 1740.440 ;
        RECT 4.400 1737.040 1495.600 1738.440 ;
        RECT 2.365 1735.040 1497.695 1737.040 ;
        RECT 4.400 1733.640 1495.600 1735.040 ;
        RECT 2.365 1731.640 1497.695 1733.640 ;
        RECT 4.400 1730.240 1495.600 1731.640 ;
        RECT 2.365 1728.240 1497.695 1730.240 ;
        RECT 4.400 1726.840 1495.600 1728.240 ;
        RECT 2.365 1724.840 1497.695 1726.840 ;
        RECT 4.400 1723.440 1497.695 1724.840 ;
        RECT 2.365 1721.440 1497.695 1723.440 ;
        RECT 4.400 1720.040 1495.600 1721.440 ;
        RECT 2.365 1718.040 1497.695 1720.040 ;
        RECT 2.365 1716.640 1495.600 1718.040 ;
        RECT 2.365 1714.640 1497.695 1716.640 ;
        RECT 4.400 1713.240 1495.600 1714.640 ;
        RECT 2.365 1711.240 1497.695 1713.240 ;
        RECT 4.400 1709.840 1495.600 1711.240 ;
        RECT 2.365 1707.840 1497.695 1709.840 ;
        RECT 4.400 1706.440 1495.600 1707.840 ;
        RECT 2.365 1704.440 1497.695 1706.440 ;
        RECT 4.400 1703.040 1495.600 1704.440 ;
        RECT 2.365 1701.040 1497.695 1703.040 ;
        RECT 4.400 1699.640 1497.695 1701.040 ;
        RECT 2.365 1697.640 1497.695 1699.640 ;
        RECT 4.400 1696.240 1495.600 1697.640 ;
        RECT 2.365 1694.240 1497.695 1696.240 ;
        RECT 2.365 1692.840 1495.600 1694.240 ;
        RECT 2.365 1690.840 1497.695 1692.840 ;
        RECT 4.400 1689.440 1495.600 1690.840 ;
        RECT 2.365 1687.440 1497.695 1689.440 ;
        RECT 4.400 1686.040 1495.600 1687.440 ;
        RECT 2.365 1684.040 1497.695 1686.040 ;
        RECT 4.400 1682.640 1495.600 1684.040 ;
        RECT 2.365 1680.640 1497.695 1682.640 ;
        RECT 4.400 1679.240 1495.600 1680.640 ;
        RECT 2.365 1677.240 1497.695 1679.240 ;
        RECT 4.400 1675.840 1495.600 1677.240 ;
        RECT 2.365 1673.840 1497.695 1675.840 ;
        RECT 4.400 1672.440 1497.695 1673.840 ;
        RECT 2.365 1670.440 1497.695 1672.440 ;
        RECT 4.400 1669.040 1495.600 1670.440 ;
        RECT 2.365 1667.040 1497.695 1669.040 ;
        RECT 2.365 1665.640 1495.600 1667.040 ;
        RECT 2.365 1663.640 1497.695 1665.640 ;
        RECT 4.400 1662.240 1495.600 1663.640 ;
        RECT 2.365 1660.240 1497.695 1662.240 ;
        RECT 4.400 1658.840 1495.600 1660.240 ;
        RECT 2.365 1656.840 1497.695 1658.840 ;
        RECT 4.400 1655.440 1495.600 1656.840 ;
        RECT 2.365 1653.440 1497.695 1655.440 ;
        RECT 4.400 1652.040 1495.600 1653.440 ;
        RECT 2.365 1650.040 1497.695 1652.040 ;
        RECT 4.400 1648.640 1497.695 1650.040 ;
        RECT 2.365 1646.640 1497.695 1648.640 ;
        RECT 4.400 1645.240 1495.600 1646.640 ;
        RECT 2.365 1643.240 1497.695 1645.240 ;
        RECT 2.365 1641.840 1495.600 1643.240 ;
        RECT 2.365 1639.840 1497.695 1641.840 ;
        RECT 4.400 1638.440 1495.600 1639.840 ;
        RECT 2.365 1636.440 1497.695 1638.440 ;
        RECT 4.400 1635.040 1495.600 1636.440 ;
        RECT 2.365 1633.040 1497.695 1635.040 ;
        RECT 4.400 1631.640 1495.600 1633.040 ;
        RECT 2.365 1629.640 1497.695 1631.640 ;
        RECT 4.400 1628.240 1495.600 1629.640 ;
        RECT 2.365 1626.240 1497.695 1628.240 ;
        RECT 4.400 1624.840 1495.600 1626.240 ;
        RECT 2.365 1622.840 1497.695 1624.840 ;
        RECT 4.400 1621.440 1497.695 1622.840 ;
        RECT 2.365 1619.440 1497.695 1621.440 ;
        RECT 4.400 1618.040 1495.600 1619.440 ;
        RECT 2.365 1616.040 1497.695 1618.040 ;
        RECT 2.365 1614.640 1495.600 1616.040 ;
        RECT 2.365 1612.640 1497.695 1614.640 ;
        RECT 4.400 1611.240 1495.600 1612.640 ;
        RECT 2.365 1609.240 1497.695 1611.240 ;
        RECT 4.400 1607.840 1495.600 1609.240 ;
        RECT 2.365 1605.840 1497.695 1607.840 ;
        RECT 4.400 1604.440 1495.600 1605.840 ;
        RECT 2.365 1602.440 1497.695 1604.440 ;
        RECT 4.400 1601.040 1495.600 1602.440 ;
        RECT 2.365 1599.040 1497.695 1601.040 ;
        RECT 4.400 1597.640 1497.695 1599.040 ;
        RECT 2.365 1595.640 1497.695 1597.640 ;
        RECT 4.400 1594.240 1495.600 1595.640 ;
        RECT 2.365 1592.240 1497.695 1594.240 ;
        RECT 2.365 1590.840 1495.600 1592.240 ;
        RECT 2.365 1588.840 1497.695 1590.840 ;
        RECT 4.400 1587.440 1495.600 1588.840 ;
        RECT 2.365 1585.440 1497.695 1587.440 ;
        RECT 4.400 1584.040 1495.600 1585.440 ;
        RECT 2.365 1582.040 1497.695 1584.040 ;
        RECT 4.400 1580.640 1495.600 1582.040 ;
        RECT 2.365 1578.640 1497.695 1580.640 ;
        RECT 4.400 1577.240 1495.600 1578.640 ;
        RECT 2.365 1575.240 1497.695 1577.240 ;
        RECT 4.400 1573.840 1497.695 1575.240 ;
        RECT 2.365 1571.840 1497.695 1573.840 ;
        RECT 4.400 1570.440 1495.600 1571.840 ;
        RECT 2.365 1568.440 1497.695 1570.440 ;
        RECT 4.400 1567.040 1495.600 1568.440 ;
        RECT 2.365 1565.040 1497.695 1567.040 ;
        RECT 2.365 1563.640 1495.600 1565.040 ;
        RECT 2.365 1561.640 1497.695 1563.640 ;
        RECT 4.400 1560.240 1495.600 1561.640 ;
        RECT 2.365 1558.240 1497.695 1560.240 ;
        RECT 4.400 1556.840 1495.600 1558.240 ;
        RECT 2.365 1554.840 1497.695 1556.840 ;
        RECT 4.400 1553.440 1495.600 1554.840 ;
        RECT 2.365 1551.440 1497.695 1553.440 ;
        RECT 4.400 1550.040 1495.600 1551.440 ;
        RECT 2.365 1548.040 1497.695 1550.040 ;
        RECT 4.400 1546.640 1497.695 1548.040 ;
        RECT 2.365 1544.640 1497.695 1546.640 ;
        RECT 4.400 1543.240 1495.600 1544.640 ;
        RECT 2.365 1541.240 1497.695 1543.240 ;
        RECT 2.365 1539.840 1495.600 1541.240 ;
        RECT 2.365 1537.840 1497.695 1539.840 ;
        RECT 4.400 1536.440 1495.600 1537.840 ;
        RECT 2.365 1534.440 1497.695 1536.440 ;
        RECT 4.400 1533.040 1495.600 1534.440 ;
        RECT 2.365 1531.040 1497.695 1533.040 ;
        RECT 4.400 1529.640 1495.600 1531.040 ;
        RECT 2.365 1527.640 1497.695 1529.640 ;
        RECT 4.400 1526.240 1495.600 1527.640 ;
        RECT 2.365 1524.240 1497.695 1526.240 ;
        RECT 4.400 1522.840 1497.695 1524.240 ;
        RECT 2.365 1520.840 1497.695 1522.840 ;
        RECT 4.400 1519.440 1495.600 1520.840 ;
        RECT 2.365 1517.440 1497.695 1519.440 ;
        RECT 4.400 1516.040 1495.600 1517.440 ;
        RECT 2.365 1514.040 1497.695 1516.040 ;
        RECT 2.365 1512.640 1495.600 1514.040 ;
        RECT 2.365 1510.640 1497.695 1512.640 ;
        RECT 4.400 1509.240 1495.600 1510.640 ;
        RECT 2.365 1507.240 1497.695 1509.240 ;
        RECT 4.400 1505.840 1495.600 1507.240 ;
        RECT 2.365 1503.840 1497.695 1505.840 ;
        RECT 4.400 1502.440 1495.600 1503.840 ;
        RECT 2.365 1500.440 1497.695 1502.440 ;
        RECT 4.400 1499.040 1495.600 1500.440 ;
        RECT 2.365 1497.040 1497.695 1499.040 ;
        RECT 4.400 1495.640 1497.695 1497.040 ;
        RECT 2.365 1493.640 1497.695 1495.640 ;
        RECT 4.400 1492.240 1495.600 1493.640 ;
        RECT 2.365 1490.240 1497.695 1492.240 ;
        RECT 2.365 1488.840 1495.600 1490.240 ;
        RECT 2.365 1486.840 1497.695 1488.840 ;
        RECT 4.400 1485.440 1495.600 1486.840 ;
        RECT 2.365 1483.440 1497.695 1485.440 ;
        RECT 4.400 1482.040 1495.600 1483.440 ;
        RECT 2.365 1480.040 1497.695 1482.040 ;
        RECT 4.400 1478.640 1495.600 1480.040 ;
        RECT 2.365 1476.640 1497.695 1478.640 ;
        RECT 4.400 1475.240 1495.600 1476.640 ;
        RECT 2.365 1473.240 1497.695 1475.240 ;
        RECT 4.400 1471.840 1497.695 1473.240 ;
        RECT 2.365 1469.840 1497.695 1471.840 ;
        RECT 4.400 1468.440 1495.600 1469.840 ;
        RECT 2.365 1466.440 1497.695 1468.440 ;
        RECT 2.365 1465.040 1495.600 1466.440 ;
        RECT 2.365 1463.040 1497.695 1465.040 ;
        RECT 4.400 1461.640 1495.600 1463.040 ;
        RECT 2.365 1459.640 1497.695 1461.640 ;
        RECT 4.400 1458.240 1495.600 1459.640 ;
        RECT 2.365 1456.240 1497.695 1458.240 ;
        RECT 4.400 1454.840 1495.600 1456.240 ;
        RECT 2.365 1452.840 1497.695 1454.840 ;
        RECT 4.400 1451.440 1495.600 1452.840 ;
        RECT 2.365 1449.440 1497.695 1451.440 ;
        RECT 4.400 1448.040 1495.600 1449.440 ;
        RECT 2.365 1446.040 1497.695 1448.040 ;
        RECT 4.400 1444.640 1497.695 1446.040 ;
        RECT 2.365 1442.640 1497.695 1444.640 ;
        RECT 4.400 1441.240 1495.600 1442.640 ;
        RECT 2.365 1439.240 1497.695 1441.240 ;
        RECT 2.365 1437.840 1495.600 1439.240 ;
        RECT 2.365 1435.840 1497.695 1437.840 ;
        RECT 4.400 1434.440 1495.600 1435.840 ;
        RECT 2.365 1432.440 1497.695 1434.440 ;
        RECT 4.400 1431.040 1495.600 1432.440 ;
        RECT 2.365 1429.040 1497.695 1431.040 ;
        RECT 4.400 1427.640 1495.600 1429.040 ;
        RECT 2.365 1425.640 1497.695 1427.640 ;
        RECT 4.400 1424.240 1495.600 1425.640 ;
        RECT 2.365 1422.240 1497.695 1424.240 ;
        RECT 4.400 1420.840 1497.695 1422.240 ;
        RECT 2.365 1418.840 1497.695 1420.840 ;
        RECT 4.400 1417.440 1495.600 1418.840 ;
        RECT 2.365 1415.440 1497.695 1417.440 ;
        RECT 2.365 1414.040 1495.600 1415.440 ;
        RECT 2.365 1412.040 1497.695 1414.040 ;
        RECT 4.400 1410.640 1495.600 1412.040 ;
        RECT 2.365 1408.640 1497.695 1410.640 ;
        RECT 4.400 1407.240 1495.600 1408.640 ;
        RECT 2.365 1405.240 1497.695 1407.240 ;
        RECT 4.400 1403.840 1495.600 1405.240 ;
        RECT 2.365 1401.840 1497.695 1403.840 ;
        RECT 4.400 1400.440 1495.600 1401.840 ;
        RECT 2.365 1398.440 1497.695 1400.440 ;
        RECT 4.400 1397.040 1497.695 1398.440 ;
        RECT 2.365 1395.040 1497.695 1397.040 ;
        RECT 4.400 1393.640 1495.600 1395.040 ;
        RECT 2.365 1391.640 1497.695 1393.640 ;
        RECT 4.400 1390.240 1495.600 1391.640 ;
        RECT 2.365 1388.240 1497.695 1390.240 ;
        RECT 2.365 1386.840 1495.600 1388.240 ;
        RECT 2.365 1384.840 1497.695 1386.840 ;
        RECT 4.400 1383.440 1495.600 1384.840 ;
        RECT 2.365 1381.440 1497.695 1383.440 ;
        RECT 4.400 1380.040 1495.600 1381.440 ;
        RECT 2.365 1378.040 1497.695 1380.040 ;
        RECT 4.400 1376.640 1495.600 1378.040 ;
        RECT 2.365 1374.640 1497.695 1376.640 ;
        RECT 4.400 1373.240 1495.600 1374.640 ;
        RECT 2.365 1371.240 1497.695 1373.240 ;
        RECT 4.400 1369.840 1497.695 1371.240 ;
        RECT 2.365 1367.840 1497.695 1369.840 ;
        RECT 4.400 1366.440 1495.600 1367.840 ;
        RECT 2.365 1364.440 1497.695 1366.440 ;
        RECT 2.365 1363.040 1495.600 1364.440 ;
        RECT 2.365 1361.040 1497.695 1363.040 ;
        RECT 4.400 1359.640 1495.600 1361.040 ;
        RECT 2.365 1357.640 1497.695 1359.640 ;
        RECT 4.400 1356.240 1495.600 1357.640 ;
        RECT 2.365 1354.240 1497.695 1356.240 ;
        RECT 4.400 1352.840 1495.600 1354.240 ;
        RECT 2.365 1350.840 1497.695 1352.840 ;
        RECT 4.400 1349.440 1495.600 1350.840 ;
        RECT 2.365 1347.440 1497.695 1349.440 ;
        RECT 4.400 1346.040 1497.695 1347.440 ;
        RECT 2.365 1344.040 1497.695 1346.040 ;
        RECT 4.400 1342.640 1495.600 1344.040 ;
        RECT 2.365 1340.640 1497.695 1342.640 ;
        RECT 4.400 1339.240 1495.600 1340.640 ;
        RECT 2.365 1337.240 1497.695 1339.240 ;
        RECT 2.365 1335.840 1495.600 1337.240 ;
        RECT 2.365 1333.840 1497.695 1335.840 ;
        RECT 4.400 1332.440 1495.600 1333.840 ;
        RECT 2.365 1330.440 1497.695 1332.440 ;
        RECT 4.400 1329.040 1495.600 1330.440 ;
        RECT 2.365 1327.040 1497.695 1329.040 ;
        RECT 4.400 1325.640 1495.600 1327.040 ;
        RECT 2.365 1323.640 1497.695 1325.640 ;
        RECT 4.400 1322.240 1495.600 1323.640 ;
        RECT 2.365 1320.240 1497.695 1322.240 ;
        RECT 4.400 1318.840 1497.695 1320.240 ;
        RECT 2.365 1316.840 1497.695 1318.840 ;
        RECT 4.400 1315.440 1495.600 1316.840 ;
        RECT 2.365 1313.440 1497.695 1315.440 ;
        RECT 2.365 1312.040 1495.600 1313.440 ;
        RECT 2.365 1310.040 1497.695 1312.040 ;
        RECT 4.400 1308.640 1495.600 1310.040 ;
        RECT 2.365 1306.640 1497.695 1308.640 ;
        RECT 4.400 1305.240 1495.600 1306.640 ;
        RECT 2.365 1303.240 1497.695 1305.240 ;
        RECT 4.400 1301.840 1495.600 1303.240 ;
        RECT 2.365 1299.840 1497.695 1301.840 ;
        RECT 4.400 1298.440 1495.600 1299.840 ;
        RECT 2.365 1296.440 1497.695 1298.440 ;
        RECT 4.400 1295.040 1497.695 1296.440 ;
        RECT 2.365 1293.040 1497.695 1295.040 ;
        RECT 4.400 1291.640 1495.600 1293.040 ;
        RECT 2.365 1289.640 1497.695 1291.640 ;
        RECT 2.365 1288.240 1495.600 1289.640 ;
        RECT 2.365 1286.240 1497.695 1288.240 ;
        RECT 4.400 1284.840 1495.600 1286.240 ;
        RECT 2.365 1282.840 1497.695 1284.840 ;
        RECT 4.400 1281.440 1495.600 1282.840 ;
        RECT 2.365 1279.440 1497.695 1281.440 ;
        RECT 4.400 1278.040 1495.600 1279.440 ;
        RECT 2.365 1276.040 1497.695 1278.040 ;
        RECT 4.400 1274.640 1495.600 1276.040 ;
        RECT 2.365 1272.640 1497.695 1274.640 ;
        RECT 4.400 1271.240 1495.600 1272.640 ;
        RECT 2.365 1269.240 1497.695 1271.240 ;
        RECT 4.400 1267.840 1497.695 1269.240 ;
        RECT 2.365 1265.840 1497.695 1267.840 ;
        RECT 4.400 1264.440 1495.600 1265.840 ;
        RECT 2.365 1262.440 1497.695 1264.440 ;
        RECT 2.365 1261.040 1495.600 1262.440 ;
        RECT 2.365 1259.040 1497.695 1261.040 ;
        RECT 4.400 1257.640 1495.600 1259.040 ;
        RECT 2.365 1255.640 1497.695 1257.640 ;
        RECT 4.400 1254.240 1495.600 1255.640 ;
        RECT 2.365 1252.240 1497.695 1254.240 ;
        RECT 4.400 1250.840 1495.600 1252.240 ;
        RECT 2.365 1248.840 1497.695 1250.840 ;
        RECT 4.400 1247.440 1495.600 1248.840 ;
        RECT 2.365 1245.440 1497.695 1247.440 ;
        RECT 4.400 1244.040 1497.695 1245.440 ;
        RECT 2.365 1242.040 1497.695 1244.040 ;
        RECT 4.400 1240.640 1495.600 1242.040 ;
        RECT 2.365 1238.640 1497.695 1240.640 ;
        RECT 2.365 1237.240 1495.600 1238.640 ;
        RECT 2.365 1235.240 1497.695 1237.240 ;
        RECT 4.400 1233.840 1495.600 1235.240 ;
        RECT 2.365 1231.840 1497.695 1233.840 ;
        RECT 4.400 1230.440 1495.600 1231.840 ;
        RECT 2.365 1228.440 1497.695 1230.440 ;
        RECT 4.400 1227.040 1495.600 1228.440 ;
        RECT 2.365 1225.040 1497.695 1227.040 ;
        RECT 4.400 1223.640 1495.600 1225.040 ;
        RECT 2.365 1221.640 1497.695 1223.640 ;
        RECT 4.400 1220.240 1497.695 1221.640 ;
        RECT 2.365 1218.240 1497.695 1220.240 ;
        RECT 4.400 1216.840 1495.600 1218.240 ;
        RECT 2.365 1214.840 1497.695 1216.840 ;
        RECT 4.400 1213.440 1495.600 1214.840 ;
        RECT 2.365 1211.440 1497.695 1213.440 ;
        RECT 2.365 1210.040 1495.600 1211.440 ;
        RECT 2.365 1208.040 1497.695 1210.040 ;
        RECT 4.400 1206.640 1495.600 1208.040 ;
        RECT 2.365 1204.640 1497.695 1206.640 ;
        RECT 4.400 1203.240 1495.600 1204.640 ;
        RECT 2.365 1201.240 1497.695 1203.240 ;
        RECT 4.400 1199.840 1495.600 1201.240 ;
        RECT 2.365 1197.840 1497.695 1199.840 ;
        RECT 4.400 1196.440 1495.600 1197.840 ;
        RECT 2.365 1194.440 1497.695 1196.440 ;
        RECT 4.400 1193.040 1497.695 1194.440 ;
        RECT 2.365 1191.040 1497.695 1193.040 ;
        RECT 4.400 1189.640 1495.600 1191.040 ;
        RECT 2.365 1187.640 1497.695 1189.640 ;
        RECT 2.365 1186.240 1495.600 1187.640 ;
        RECT 2.365 1184.240 1497.695 1186.240 ;
        RECT 4.400 1182.840 1495.600 1184.240 ;
        RECT 2.365 1180.840 1497.695 1182.840 ;
        RECT 4.400 1179.440 1495.600 1180.840 ;
        RECT 2.365 1177.440 1497.695 1179.440 ;
        RECT 4.400 1176.040 1495.600 1177.440 ;
        RECT 2.365 1174.040 1497.695 1176.040 ;
        RECT 4.400 1172.640 1495.600 1174.040 ;
        RECT 2.365 1170.640 1497.695 1172.640 ;
        RECT 4.400 1169.240 1497.695 1170.640 ;
        RECT 2.365 1167.240 1497.695 1169.240 ;
        RECT 4.400 1165.840 1495.600 1167.240 ;
        RECT 2.365 1163.840 1497.695 1165.840 ;
        RECT 4.400 1162.440 1495.600 1163.840 ;
        RECT 2.365 1160.440 1497.695 1162.440 ;
        RECT 2.365 1159.040 1495.600 1160.440 ;
        RECT 2.365 1157.040 1497.695 1159.040 ;
        RECT 4.400 1155.640 1495.600 1157.040 ;
        RECT 2.365 1153.640 1497.695 1155.640 ;
        RECT 4.400 1152.240 1495.600 1153.640 ;
        RECT 2.365 1150.240 1497.695 1152.240 ;
        RECT 4.400 1148.840 1495.600 1150.240 ;
        RECT 2.365 1146.840 1497.695 1148.840 ;
        RECT 4.400 1145.440 1495.600 1146.840 ;
        RECT 2.365 1143.440 1497.695 1145.440 ;
        RECT 4.400 1142.040 1497.695 1143.440 ;
        RECT 2.365 1140.040 1497.695 1142.040 ;
        RECT 4.400 1138.640 1495.600 1140.040 ;
        RECT 2.365 1136.640 1497.695 1138.640 ;
        RECT 2.365 1135.240 1495.600 1136.640 ;
        RECT 2.365 1133.240 1497.695 1135.240 ;
        RECT 4.400 1131.840 1495.600 1133.240 ;
        RECT 2.365 1129.840 1497.695 1131.840 ;
        RECT 4.400 1128.440 1495.600 1129.840 ;
        RECT 2.365 1126.440 1497.695 1128.440 ;
        RECT 4.400 1125.040 1495.600 1126.440 ;
        RECT 2.365 1123.040 1497.695 1125.040 ;
        RECT 4.400 1121.640 1495.600 1123.040 ;
        RECT 2.365 1119.640 1497.695 1121.640 ;
        RECT 4.400 1118.240 1497.695 1119.640 ;
        RECT 2.365 1116.240 1497.695 1118.240 ;
        RECT 4.400 1114.840 1495.600 1116.240 ;
        RECT 2.365 1112.840 1497.695 1114.840 ;
        RECT 2.365 1111.440 1495.600 1112.840 ;
        RECT 2.365 1109.440 1497.695 1111.440 ;
        RECT 4.400 1108.040 1495.600 1109.440 ;
        RECT 2.365 1106.040 1497.695 1108.040 ;
        RECT 4.400 1104.640 1495.600 1106.040 ;
        RECT 2.365 1102.640 1497.695 1104.640 ;
        RECT 4.400 1101.240 1495.600 1102.640 ;
        RECT 2.365 1099.240 1497.695 1101.240 ;
        RECT 4.400 1097.840 1495.600 1099.240 ;
        RECT 2.365 1095.840 1497.695 1097.840 ;
        RECT 4.400 1094.440 1495.600 1095.840 ;
        RECT 2.365 1092.440 1497.695 1094.440 ;
        RECT 4.400 1091.040 1497.695 1092.440 ;
        RECT 2.365 1089.040 1497.695 1091.040 ;
        RECT 4.400 1087.640 1495.600 1089.040 ;
        RECT 2.365 1085.640 1497.695 1087.640 ;
        RECT 2.365 1084.240 1495.600 1085.640 ;
        RECT 2.365 1082.240 1497.695 1084.240 ;
        RECT 4.400 1080.840 1495.600 1082.240 ;
        RECT 2.365 1078.840 1497.695 1080.840 ;
        RECT 4.400 1077.440 1495.600 1078.840 ;
        RECT 2.365 1075.440 1497.695 1077.440 ;
        RECT 4.400 1074.040 1495.600 1075.440 ;
        RECT 2.365 1072.040 1497.695 1074.040 ;
        RECT 4.400 1070.640 1495.600 1072.040 ;
        RECT 2.365 1068.640 1497.695 1070.640 ;
        RECT 4.400 1067.240 1497.695 1068.640 ;
        RECT 2.365 1065.240 1497.695 1067.240 ;
        RECT 4.400 1063.840 1495.600 1065.240 ;
        RECT 2.365 1061.840 1497.695 1063.840 ;
        RECT 2.365 1060.440 1495.600 1061.840 ;
        RECT 2.365 1058.440 1497.695 1060.440 ;
        RECT 4.400 1057.040 1495.600 1058.440 ;
        RECT 2.365 1055.040 1497.695 1057.040 ;
        RECT 4.400 1053.640 1495.600 1055.040 ;
        RECT 2.365 1051.640 1497.695 1053.640 ;
        RECT 4.400 1050.240 1495.600 1051.640 ;
        RECT 2.365 1048.240 1497.695 1050.240 ;
        RECT 4.400 1046.840 1495.600 1048.240 ;
        RECT 2.365 1044.840 1497.695 1046.840 ;
        RECT 4.400 1043.440 1497.695 1044.840 ;
        RECT 2.365 1041.440 1497.695 1043.440 ;
        RECT 4.400 1040.040 1495.600 1041.440 ;
        RECT 2.365 1038.040 1497.695 1040.040 ;
        RECT 4.400 1036.640 1495.600 1038.040 ;
        RECT 2.365 1034.640 1497.695 1036.640 ;
        RECT 2.365 1033.240 1495.600 1034.640 ;
        RECT 2.365 1031.240 1497.695 1033.240 ;
        RECT 4.400 1029.840 1495.600 1031.240 ;
        RECT 2.365 1027.840 1497.695 1029.840 ;
        RECT 4.400 1026.440 1495.600 1027.840 ;
        RECT 2.365 1024.440 1497.695 1026.440 ;
        RECT 4.400 1023.040 1495.600 1024.440 ;
        RECT 2.365 1021.040 1497.695 1023.040 ;
        RECT 4.400 1019.640 1495.600 1021.040 ;
        RECT 2.365 1017.640 1497.695 1019.640 ;
        RECT 4.400 1016.240 1497.695 1017.640 ;
        RECT 2.365 1014.240 1497.695 1016.240 ;
        RECT 4.400 1012.840 1495.600 1014.240 ;
        RECT 2.365 1010.840 1497.695 1012.840 ;
        RECT 2.365 1009.440 1495.600 1010.840 ;
        RECT 2.365 1007.440 1497.695 1009.440 ;
        RECT 4.400 1006.040 1495.600 1007.440 ;
        RECT 2.365 1004.040 1497.695 1006.040 ;
        RECT 4.400 1002.640 1495.600 1004.040 ;
        RECT 2.365 1000.640 1497.695 1002.640 ;
        RECT 4.400 999.240 1495.600 1000.640 ;
        RECT 2.365 997.240 1497.695 999.240 ;
        RECT 4.400 995.840 1495.600 997.240 ;
        RECT 2.365 993.840 1497.695 995.840 ;
        RECT 4.400 992.440 1497.695 993.840 ;
        RECT 2.365 990.440 1497.695 992.440 ;
        RECT 4.400 989.040 1495.600 990.440 ;
        RECT 2.365 987.040 1497.695 989.040 ;
        RECT 4.400 985.640 1495.600 987.040 ;
        RECT 2.365 983.640 1497.695 985.640 ;
        RECT 2.365 982.240 1495.600 983.640 ;
        RECT 2.365 980.240 1497.695 982.240 ;
        RECT 4.400 978.840 1495.600 980.240 ;
        RECT 2.365 976.840 1497.695 978.840 ;
        RECT 4.400 975.440 1495.600 976.840 ;
        RECT 2.365 973.440 1497.695 975.440 ;
        RECT 4.400 972.040 1495.600 973.440 ;
        RECT 2.365 970.040 1497.695 972.040 ;
        RECT 4.400 968.640 1495.600 970.040 ;
        RECT 2.365 966.640 1497.695 968.640 ;
        RECT 4.400 965.240 1497.695 966.640 ;
        RECT 2.365 963.240 1497.695 965.240 ;
        RECT 4.400 961.840 1495.600 963.240 ;
        RECT 2.365 959.840 1497.695 961.840 ;
        RECT 2.365 958.440 1495.600 959.840 ;
        RECT 2.365 956.440 1497.695 958.440 ;
        RECT 4.400 955.040 1495.600 956.440 ;
        RECT 2.365 953.040 1497.695 955.040 ;
        RECT 4.400 951.640 1495.600 953.040 ;
        RECT 2.365 949.640 1497.695 951.640 ;
        RECT 4.400 948.240 1495.600 949.640 ;
        RECT 2.365 946.240 1497.695 948.240 ;
        RECT 4.400 944.840 1495.600 946.240 ;
        RECT 2.365 942.840 1497.695 944.840 ;
        RECT 4.400 941.440 1497.695 942.840 ;
        RECT 2.365 939.440 1497.695 941.440 ;
        RECT 4.400 938.040 1495.600 939.440 ;
        RECT 2.365 936.040 1497.695 938.040 ;
        RECT 2.365 934.640 1495.600 936.040 ;
        RECT 2.365 932.640 1497.695 934.640 ;
        RECT 4.400 931.240 1495.600 932.640 ;
        RECT 2.365 929.240 1497.695 931.240 ;
        RECT 4.400 927.840 1495.600 929.240 ;
        RECT 2.365 925.840 1497.695 927.840 ;
        RECT 4.400 924.440 1495.600 925.840 ;
        RECT 2.365 922.440 1497.695 924.440 ;
        RECT 4.400 921.040 1495.600 922.440 ;
        RECT 2.365 919.040 1497.695 921.040 ;
        RECT 4.400 917.640 1495.600 919.040 ;
        RECT 2.365 915.640 1497.695 917.640 ;
        RECT 4.400 914.240 1497.695 915.640 ;
        RECT 2.365 912.240 1497.695 914.240 ;
        RECT 4.400 910.840 1495.600 912.240 ;
        RECT 2.365 908.840 1497.695 910.840 ;
        RECT 2.365 907.440 1495.600 908.840 ;
        RECT 2.365 905.440 1497.695 907.440 ;
        RECT 4.400 904.040 1495.600 905.440 ;
        RECT 2.365 902.040 1497.695 904.040 ;
        RECT 4.400 900.640 1495.600 902.040 ;
        RECT 2.365 898.640 1497.695 900.640 ;
        RECT 4.400 897.240 1495.600 898.640 ;
        RECT 2.365 895.240 1497.695 897.240 ;
        RECT 4.400 893.840 1495.600 895.240 ;
        RECT 2.365 891.840 1497.695 893.840 ;
        RECT 4.400 890.440 1497.695 891.840 ;
        RECT 2.365 888.440 1497.695 890.440 ;
        RECT 4.400 887.040 1495.600 888.440 ;
        RECT 2.365 885.040 1497.695 887.040 ;
        RECT 2.365 883.640 1495.600 885.040 ;
        RECT 2.365 881.640 1497.695 883.640 ;
        RECT 4.400 880.240 1495.600 881.640 ;
        RECT 2.365 878.240 1497.695 880.240 ;
        RECT 4.400 876.840 1495.600 878.240 ;
        RECT 2.365 874.840 1497.695 876.840 ;
        RECT 4.400 873.440 1495.600 874.840 ;
        RECT 2.365 871.440 1497.695 873.440 ;
        RECT 4.400 870.040 1495.600 871.440 ;
        RECT 2.365 868.040 1497.695 870.040 ;
        RECT 4.400 866.640 1495.600 868.040 ;
        RECT 2.365 864.640 1497.695 866.640 ;
        RECT 4.400 863.240 1497.695 864.640 ;
        RECT 2.365 861.240 1497.695 863.240 ;
        RECT 4.400 859.840 1495.600 861.240 ;
        RECT 2.365 857.840 1497.695 859.840 ;
        RECT 2.365 856.440 1495.600 857.840 ;
        RECT 2.365 854.440 1497.695 856.440 ;
        RECT 4.400 853.040 1495.600 854.440 ;
        RECT 2.365 851.040 1497.695 853.040 ;
        RECT 4.400 849.640 1495.600 851.040 ;
        RECT 2.365 847.640 1497.695 849.640 ;
        RECT 4.400 846.240 1495.600 847.640 ;
        RECT 2.365 844.240 1497.695 846.240 ;
        RECT 4.400 842.840 1495.600 844.240 ;
        RECT 2.365 840.840 1497.695 842.840 ;
        RECT 4.400 839.440 1497.695 840.840 ;
        RECT 2.365 837.440 1497.695 839.440 ;
        RECT 4.400 836.040 1495.600 837.440 ;
        RECT 2.365 834.040 1497.695 836.040 ;
        RECT 2.365 832.640 1495.600 834.040 ;
        RECT 2.365 830.640 1497.695 832.640 ;
        RECT 4.400 829.240 1495.600 830.640 ;
        RECT 2.365 827.240 1497.695 829.240 ;
        RECT 4.400 825.840 1495.600 827.240 ;
        RECT 2.365 823.840 1497.695 825.840 ;
        RECT 4.400 822.440 1495.600 823.840 ;
        RECT 2.365 820.440 1497.695 822.440 ;
        RECT 4.400 819.040 1495.600 820.440 ;
        RECT 2.365 817.040 1497.695 819.040 ;
        RECT 4.400 815.640 1497.695 817.040 ;
        RECT 2.365 813.640 1497.695 815.640 ;
        RECT 4.400 812.240 1495.600 813.640 ;
        RECT 2.365 810.240 1497.695 812.240 ;
        RECT 4.400 808.840 1495.600 810.240 ;
        RECT 2.365 806.840 1497.695 808.840 ;
        RECT 2.365 805.440 1495.600 806.840 ;
        RECT 2.365 803.440 1497.695 805.440 ;
        RECT 4.400 802.040 1495.600 803.440 ;
        RECT 2.365 800.040 1497.695 802.040 ;
        RECT 4.400 798.640 1495.600 800.040 ;
        RECT 2.365 796.640 1497.695 798.640 ;
        RECT 4.400 795.240 1495.600 796.640 ;
        RECT 2.365 793.240 1497.695 795.240 ;
        RECT 4.400 791.840 1495.600 793.240 ;
        RECT 2.365 789.840 1497.695 791.840 ;
        RECT 4.400 788.440 1497.695 789.840 ;
        RECT 2.365 786.440 1497.695 788.440 ;
        RECT 4.400 785.040 1495.600 786.440 ;
        RECT 2.365 783.040 1497.695 785.040 ;
        RECT 2.365 781.640 1495.600 783.040 ;
        RECT 2.365 779.640 1497.695 781.640 ;
        RECT 4.400 778.240 1495.600 779.640 ;
        RECT 2.365 776.240 1497.695 778.240 ;
        RECT 4.400 774.840 1495.600 776.240 ;
        RECT 2.365 772.840 1497.695 774.840 ;
        RECT 4.400 771.440 1495.600 772.840 ;
        RECT 2.365 769.440 1497.695 771.440 ;
        RECT 4.400 768.040 1495.600 769.440 ;
        RECT 2.365 766.040 1497.695 768.040 ;
        RECT 4.400 764.640 1497.695 766.040 ;
        RECT 2.365 762.640 1497.695 764.640 ;
        RECT 4.400 761.240 1495.600 762.640 ;
        RECT 2.365 759.240 1497.695 761.240 ;
        RECT 4.400 757.840 1495.600 759.240 ;
        RECT 2.365 755.840 1497.695 757.840 ;
        RECT 2.365 754.440 1495.600 755.840 ;
        RECT 2.365 752.440 1497.695 754.440 ;
        RECT 4.400 751.040 1495.600 752.440 ;
        RECT 2.365 749.040 1497.695 751.040 ;
        RECT 4.400 747.640 1495.600 749.040 ;
        RECT 2.365 745.640 1497.695 747.640 ;
        RECT 4.400 744.240 1495.600 745.640 ;
        RECT 2.365 742.240 1497.695 744.240 ;
        RECT 4.400 740.840 1495.600 742.240 ;
        RECT 2.365 738.840 1497.695 740.840 ;
        RECT 4.400 737.440 1497.695 738.840 ;
        RECT 2.365 735.440 1497.695 737.440 ;
        RECT 4.400 734.040 1495.600 735.440 ;
        RECT 2.365 732.040 1497.695 734.040 ;
        RECT 2.365 730.640 1495.600 732.040 ;
        RECT 2.365 728.640 1497.695 730.640 ;
        RECT 4.400 727.240 1495.600 728.640 ;
        RECT 2.365 725.240 1497.695 727.240 ;
        RECT 4.400 723.840 1495.600 725.240 ;
        RECT 2.365 721.840 1497.695 723.840 ;
        RECT 4.400 720.440 1495.600 721.840 ;
        RECT 2.365 718.440 1497.695 720.440 ;
        RECT 4.400 717.040 1495.600 718.440 ;
        RECT 2.365 715.040 1497.695 717.040 ;
        RECT 4.400 713.640 1497.695 715.040 ;
        RECT 2.365 711.640 1497.695 713.640 ;
        RECT 4.400 710.240 1495.600 711.640 ;
        RECT 2.365 708.240 1497.695 710.240 ;
        RECT 2.365 706.840 1495.600 708.240 ;
        RECT 2.365 704.840 1497.695 706.840 ;
        RECT 4.400 703.440 1495.600 704.840 ;
        RECT 2.365 701.440 1497.695 703.440 ;
        RECT 4.400 700.040 1495.600 701.440 ;
        RECT 2.365 698.040 1497.695 700.040 ;
        RECT 4.400 696.640 1495.600 698.040 ;
        RECT 2.365 694.640 1497.695 696.640 ;
        RECT 4.400 693.240 1495.600 694.640 ;
        RECT 2.365 691.240 1497.695 693.240 ;
        RECT 4.400 689.840 1495.600 691.240 ;
        RECT 2.365 687.840 1497.695 689.840 ;
        RECT 4.400 686.440 1497.695 687.840 ;
        RECT 2.365 684.440 1497.695 686.440 ;
        RECT 4.400 683.040 1495.600 684.440 ;
        RECT 2.365 681.040 1497.695 683.040 ;
        RECT 2.365 679.640 1495.600 681.040 ;
        RECT 2.365 677.640 1497.695 679.640 ;
        RECT 4.400 676.240 1495.600 677.640 ;
        RECT 2.365 674.240 1497.695 676.240 ;
        RECT 4.400 672.840 1495.600 674.240 ;
        RECT 2.365 670.840 1497.695 672.840 ;
        RECT 4.400 669.440 1495.600 670.840 ;
        RECT 2.365 667.440 1497.695 669.440 ;
        RECT 4.400 666.040 1495.600 667.440 ;
        RECT 2.365 664.040 1497.695 666.040 ;
        RECT 4.400 662.640 1497.695 664.040 ;
        RECT 2.365 660.640 1497.695 662.640 ;
        RECT 4.400 659.240 1495.600 660.640 ;
        RECT 2.365 657.240 1497.695 659.240 ;
        RECT 2.365 655.840 1495.600 657.240 ;
        RECT 2.365 653.840 1497.695 655.840 ;
        RECT 4.400 652.440 1495.600 653.840 ;
        RECT 2.365 650.440 1497.695 652.440 ;
        RECT 4.400 649.040 1495.600 650.440 ;
        RECT 2.365 647.040 1497.695 649.040 ;
        RECT 4.400 645.640 1495.600 647.040 ;
        RECT 2.365 643.640 1497.695 645.640 ;
        RECT 4.400 642.240 1495.600 643.640 ;
        RECT 2.365 640.240 1497.695 642.240 ;
        RECT 4.400 638.840 1497.695 640.240 ;
        RECT 2.365 636.840 1497.695 638.840 ;
        RECT 4.400 635.440 1495.600 636.840 ;
        RECT 2.365 633.440 1497.695 635.440 ;
        RECT 4.400 632.040 1495.600 633.440 ;
        RECT 2.365 630.040 1497.695 632.040 ;
        RECT 2.365 628.640 1495.600 630.040 ;
        RECT 2.365 626.640 1497.695 628.640 ;
        RECT 4.400 625.240 1495.600 626.640 ;
        RECT 2.365 623.240 1497.695 625.240 ;
        RECT 4.400 621.840 1495.600 623.240 ;
        RECT 2.365 619.840 1497.695 621.840 ;
        RECT 4.400 618.440 1495.600 619.840 ;
        RECT 2.365 616.440 1497.695 618.440 ;
        RECT 4.400 615.040 1495.600 616.440 ;
        RECT 2.365 613.040 1497.695 615.040 ;
        RECT 4.400 611.640 1497.695 613.040 ;
        RECT 2.365 609.640 1497.695 611.640 ;
        RECT 4.400 608.240 1495.600 609.640 ;
        RECT 2.365 606.240 1497.695 608.240 ;
        RECT 2.365 604.840 1495.600 606.240 ;
        RECT 2.365 602.840 1497.695 604.840 ;
        RECT 4.400 601.440 1495.600 602.840 ;
        RECT 2.365 599.440 1497.695 601.440 ;
        RECT 4.400 598.040 1495.600 599.440 ;
        RECT 2.365 596.040 1497.695 598.040 ;
        RECT 4.400 594.640 1495.600 596.040 ;
        RECT 2.365 592.640 1497.695 594.640 ;
        RECT 4.400 591.240 1495.600 592.640 ;
        RECT 2.365 589.240 1497.695 591.240 ;
        RECT 4.400 587.840 1497.695 589.240 ;
        RECT 2.365 585.840 1497.695 587.840 ;
        RECT 4.400 584.440 1495.600 585.840 ;
        RECT 2.365 582.440 1497.695 584.440 ;
        RECT 4.400 581.040 1495.600 582.440 ;
        RECT 2.365 579.040 1497.695 581.040 ;
        RECT 2.365 577.640 1495.600 579.040 ;
        RECT 2.365 575.640 1497.695 577.640 ;
        RECT 4.400 574.240 1495.600 575.640 ;
        RECT 2.365 572.240 1497.695 574.240 ;
        RECT 4.400 570.840 1495.600 572.240 ;
        RECT 2.365 568.840 1497.695 570.840 ;
        RECT 4.400 567.440 1495.600 568.840 ;
        RECT 2.365 565.440 1497.695 567.440 ;
        RECT 4.400 564.040 1495.600 565.440 ;
        RECT 2.365 562.040 1497.695 564.040 ;
        RECT 4.400 560.640 1497.695 562.040 ;
        RECT 2.365 558.640 1497.695 560.640 ;
        RECT 4.400 557.240 1495.600 558.640 ;
        RECT 2.365 555.240 1497.695 557.240 ;
        RECT 2.365 553.840 1495.600 555.240 ;
        RECT 2.365 551.840 1497.695 553.840 ;
        RECT 4.400 550.440 1495.600 551.840 ;
        RECT 2.365 548.440 1497.695 550.440 ;
        RECT 4.400 547.040 1495.600 548.440 ;
        RECT 2.365 545.040 1497.695 547.040 ;
        RECT 4.400 543.640 1495.600 545.040 ;
        RECT 2.365 541.640 1497.695 543.640 ;
        RECT 4.400 540.240 1495.600 541.640 ;
        RECT 2.365 538.240 1497.695 540.240 ;
        RECT 4.400 536.840 1497.695 538.240 ;
        RECT 2.365 534.840 1497.695 536.840 ;
        RECT 4.400 533.440 1495.600 534.840 ;
        RECT 2.365 531.440 1497.695 533.440 ;
        RECT 2.365 530.040 1495.600 531.440 ;
        RECT 2.365 528.040 1497.695 530.040 ;
        RECT 4.400 526.640 1495.600 528.040 ;
        RECT 2.365 524.640 1497.695 526.640 ;
        RECT 4.400 523.240 1495.600 524.640 ;
        RECT 2.365 521.240 1497.695 523.240 ;
        RECT 4.400 519.840 1495.600 521.240 ;
        RECT 2.365 517.840 1497.695 519.840 ;
        RECT 4.400 516.440 1495.600 517.840 ;
        RECT 2.365 514.440 1497.695 516.440 ;
        RECT 4.400 513.040 1495.600 514.440 ;
        RECT 2.365 511.040 1497.695 513.040 ;
        RECT 4.400 509.640 1497.695 511.040 ;
        RECT 2.365 507.640 1497.695 509.640 ;
        RECT 4.400 506.240 1495.600 507.640 ;
        RECT 2.365 504.240 1497.695 506.240 ;
        RECT 2.365 502.840 1495.600 504.240 ;
        RECT 2.365 500.840 1497.695 502.840 ;
        RECT 4.400 499.440 1495.600 500.840 ;
        RECT 2.365 497.440 1497.695 499.440 ;
        RECT 4.400 496.040 1495.600 497.440 ;
        RECT 2.365 494.040 1497.695 496.040 ;
        RECT 4.400 492.640 1495.600 494.040 ;
        RECT 2.365 490.640 1497.695 492.640 ;
        RECT 4.400 489.240 1495.600 490.640 ;
        RECT 2.365 487.240 1497.695 489.240 ;
        RECT 4.400 485.840 1497.695 487.240 ;
        RECT 2.365 483.840 1497.695 485.840 ;
        RECT 4.400 482.440 1495.600 483.840 ;
        RECT 2.365 480.440 1497.695 482.440 ;
        RECT 2.365 479.040 1495.600 480.440 ;
        RECT 2.365 477.040 1497.695 479.040 ;
        RECT 4.400 475.640 1495.600 477.040 ;
        RECT 2.365 473.640 1497.695 475.640 ;
        RECT 4.400 472.240 1495.600 473.640 ;
        RECT 2.365 470.240 1497.695 472.240 ;
        RECT 4.400 468.840 1495.600 470.240 ;
        RECT 2.365 466.840 1497.695 468.840 ;
        RECT 4.400 465.440 1495.600 466.840 ;
        RECT 2.365 463.440 1497.695 465.440 ;
        RECT 4.400 462.040 1497.695 463.440 ;
        RECT 2.365 460.040 1497.695 462.040 ;
        RECT 4.400 458.640 1495.600 460.040 ;
        RECT 2.365 456.640 1497.695 458.640 ;
        RECT 4.400 455.240 1495.600 456.640 ;
        RECT 2.365 453.240 1497.695 455.240 ;
        RECT 2.365 451.840 1495.600 453.240 ;
        RECT 2.365 449.840 1497.695 451.840 ;
        RECT 4.400 448.440 1495.600 449.840 ;
        RECT 2.365 446.440 1497.695 448.440 ;
        RECT 4.400 445.040 1495.600 446.440 ;
        RECT 2.365 443.040 1497.695 445.040 ;
        RECT 4.400 441.640 1495.600 443.040 ;
        RECT 2.365 439.640 1497.695 441.640 ;
        RECT 4.400 438.240 1495.600 439.640 ;
        RECT 2.365 436.240 1497.695 438.240 ;
        RECT 4.400 434.840 1497.695 436.240 ;
        RECT 2.365 432.840 1497.695 434.840 ;
        RECT 4.400 431.440 1495.600 432.840 ;
        RECT 2.365 429.440 1497.695 431.440 ;
        RECT 2.365 428.040 1495.600 429.440 ;
        RECT 2.365 426.040 1497.695 428.040 ;
        RECT 4.400 424.640 1495.600 426.040 ;
        RECT 2.365 422.640 1497.695 424.640 ;
        RECT 4.400 421.240 1495.600 422.640 ;
        RECT 2.365 419.240 1497.695 421.240 ;
        RECT 4.400 417.840 1495.600 419.240 ;
        RECT 2.365 415.840 1497.695 417.840 ;
        RECT 4.400 414.440 1495.600 415.840 ;
        RECT 2.365 412.440 1497.695 414.440 ;
        RECT 4.400 411.040 1497.695 412.440 ;
        RECT 2.365 409.040 1497.695 411.040 ;
        RECT 4.400 407.640 1495.600 409.040 ;
        RECT 2.365 405.640 1497.695 407.640 ;
        RECT 4.400 404.240 1495.600 405.640 ;
        RECT 2.365 402.240 1497.695 404.240 ;
        RECT 2.365 400.840 1495.600 402.240 ;
        RECT 2.365 398.840 1497.695 400.840 ;
        RECT 4.400 397.440 1495.600 398.840 ;
        RECT 2.365 395.440 1497.695 397.440 ;
        RECT 4.400 394.040 1495.600 395.440 ;
        RECT 2.365 392.040 1497.695 394.040 ;
        RECT 4.400 390.640 1495.600 392.040 ;
        RECT 2.365 388.640 1497.695 390.640 ;
        RECT 4.400 387.240 1495.600 388.640 ;
        RECT 2.365 385.240 1497.695 387.240 ;
        RECT 4.400 383.840 1497.695 385.240 ;
        RECT 2.365 381.840 1497.695 383.840 ;
        RECT 4.400 380.440 1495.600 381.840 ;
        RECT 2.365 378.440 1497.695 380.440 ;
        RECT 2.365 377.040 1495.600 378.440 ;
        RECT 2.365 375.040 1497.695 377.040 ;
        RECT 4.400 373.640 1495.600 375.040 ;
        RECT 2.365 371.640 1497.695 373.640 ;
        RECT 4.400 370.240 1495.600 371.640 ;
        RECT 2.365 368.240 1497.695 370.240 ;
        RECT 4.400 366.840 1495.600 368.240 ;
        RECT 2.365 364.840 1497.695 366.840 ;
        RECT 4.400 363.440 1495.600 364.840 ;
        RECT 2.365 361.440 1497.695 363.440 ;
        RECT 4.400 360.040 1497.695 361.440 ;
        RECT 2.365 358.040 1497.695 360.040 ;
        RECT 4.400 356.640 1495.600 358.040 ;
        RECT 2.365 354.640 1497.695 356.640 ;
        RECT 2.365 353.240 1495.600 354.640 ;
        RECT 2.365 351.240 1497.695 353.240 ;
        RECT 4.400 349.840 1495.600 351.240 ;
        RECT 2.365 347.840 1497.695 349.840 ;
        RECT 4.400 346.440 1495.600 347.840 ;
        RECT 2.365 344.440 1497.695 346.440 ;
        RECT 4.400 343.040 1495.600 344.440 ;
        RECT 2.365 341.040 1497.695 343.040 ;
        RECT 4.400 339.640 1495.600 341.040 ;
        RECT 2.365 337.640 1497.695 339.640 ;
        RECT 4.400 336.240 1495.600 337.640 ;
        RECT 2.365 334.240 1497.695 336.240 ;
        RECT 4.400 332.840 1497.695 334.240 ;
        RECT 2.365 330.840 1497.695 332.840 ;
        RECT 4.400 329.440 1495.600 330.840 ;
        RECT 2.365 327.440 1497.695 329.440 ;
        RECT 2.365 326.040 1495.600 327.440 ;
        RECT 2.365 324.040 1497.695 326.040 ;
        RECT 4.400 322.640 1495.600 324.040 ;
        RECT 2.365 320.640 1497.695 322.640 ;
        RECT 4.400 319.240 1495.600 320.640 ;
        RECT 2.365 317.240 1497.695 319.240 ;
        RECT 4.400 315.840 1495.600 317.240 ;
        RECT 2.365 313.840 1497.695 315.840 ;
        RECT 4.400 312.440 1495.600 313.840 ;
        RECT 2.365 310.440 1497.695 312.440 ;
        RECT 4.400 309.040 1497.695 310.440 ;
        RECT 2.365 307.040 1497.695 309.040 ;
        RECT 4.400 305.640 1495.600 307.040 ;
        RECT 2.365 303.640 1497.695 305.640 ;
        RECT 2.365 302.240 1495.600 303.640 ;
        RECT 2.365 300.240 1497.695 302.240 ;
        RECT 4.400 298.840 1495.600 300.240 ;
        RECT 2.365 296.840 1497.695 298.840 ;
        RECT 4.400 295.440 1495.600 296.840 ;
        RECT 2.365 293.440 1497.695 295.440 ;
        RECT 4.400 292.040 1495.600 293.440 ;
        RECT 2.365 290.040 1497.695 292.040 ;
        RECT 4.400 288.640 1495.600 290.040 ;
        RECT 2.365 286.640 1497.695 288.640 ;
        RECT 4.400 285.240 1497.695 286.640 ;
        RECT 2.365 283.240 1497.695 285.240 ;
        RECT 4.400 281.840 1495.600 283.240 ;
        RECT 2.365 279.840 1497.695 281.840 ;
        RECT 4.400 278.440 1495.600 279.840 ;
        RECT 2.365 276.440 1497.695 278.440 ;
        RECT 2.365 275.040 1495.600 276.440 ;
        RECT 2.365 273.040 1497.695 275.040 ;
        RECT 4.400 271.640 1495.600 273.040 ;
        RECT 2.365 269.640 1497.695 271.640 ;
        RECT 4.400 268.240 1495.600 269.640 ;
        RECT 2.365 266.240 1497.695 268.240 ;
        RECT 4.400 264.840 1495.600 266.240 ;
        RECT 2.365 262.840 1497.695 264.840 ;
        RECT 4.400 261.440 1495.600 262.840 ;
        RECT 2.365 259.440 1497.695 261.440 ;
        RECT 4.400 258.040 1497.695 259.440 ;
        RECT 2.365 256.040 1497.695 258.040 ;
        RECT 4.400 254.640 1495.600 256.040 ;
        RECT 2.365 252.640 1497.695 254.640 ;
        RECT 2.365 251.240 1495.600 252.640 ;
        RECT 2.365 249.240 1497.695 251.240 ;
        RECT 4.400 247.840 1495.600 249.240 ;
        RECT 2.365 245.840 1497.695 247.840 ;
        RECT 4.400 244.440 1495.600 245.840 ;
        RECT 2.365 242.440 1497.695 244.440 ;
        RECT 4.400 241.040 1495.600 242.440 ;
        RECT 2.365 239.040 1497.695 241.040 ;
        RECT 4.400 237.640 1495.600 239.040 ;
        RECT 2.365 235.640 1497.695 237.640 ;
        RECT 4.400 234.240 1497.695 235.640 ;
        RECT 2.365 232.240 1497.695 234.240 ;
        RECT 4.400 230.840 1495.600 232.240 ;
        RECT 2.365 228.840 1497.695 230.840 ;
        RECT 4.400 227.440 1495.600 228.840 ;
        RECT 2.365 225.440 1497.695 227.440 ;
        RECT 2.365 224.040 1495.600 225.440 ;
        RECT 2.365 222.040 1497.695 224.040 ;
        RECT 4.400 220.640 1495.600 222.040 ;
        RECT 2.365 218.640 1497.695 220.640 ;
        RECT 4.400 217.240 1495.600 218.640 ;
        RECT 2.365 215.240 1497.695 217.240 ;
        RECT 4.400 213.840 1495.600 215.240 ;
        RECT 2.365 211.840 1497.695 213.840 ;
        RECT 4.400 210.440 1495.600 211.840 ;
        RECT 2.365 208.440 1497.695 210.440 ;
        RECT 4.400 207.040 1497.695 208.440 ;
        RECT 2.365 205.040 1497.695 207.040 ;
        RECT 4.400 203.640 1495.600 205.040 ;
        RECT 2.365 201.640 1497.695 203.640 ;
        RECT 2.365 200.240 1495.600 201.640 ;
        RECT 2.365 198.240 1497.695 200.240 ;
        RECT 4.400 196.840 1495.600 198.240 ;
        RECT 2.365 194.840 1497.695 196.840 ;
        RECT 4.400 193.440 1495.600 194.840 ;
        RECT 2.365 191.440 1497.695 193.440 ;
        RECT 4.400 190.040 1495.600 191.440 ;
        RECT 2.365 188.040 1497.695 190.040 ;
        RECT 4.400 186.640 1495.600 188.040 ;
        RECT 2.365 184.640 1497.695 186.640 ;
        RECT 4.400 183.240 1497.695 184.640 ;
        RECT 2.365 181.240 1497.695 183.240 ;
        RECT 4.400 179.840 1495.600 181.240 ;
        RECT 2.365 177.840 1497.695 179.840 ;
        RECT 2.365 176.440 1495.600 177.840 ;
        RECT 2.365 174.440 1497.695 176.440 ;
        RECT 4.400 173.040 1495.600 174.440 ;
        RECT 2.365 171.040 1497.695 173.040 ;
        RECT 4.400 169.640 1495.600 171.040 ;
        RECT 2.365 167.640 1497.695 169.640 ;
        RECT 4.400 166.240 1495.600 167.640 ;
        RECT 2.365 164.240 1497.695 166.240 ;
        RECT 4.400 162.840 1495.600 164.240 ;
        RECT 2.365 160.840 1497.695 162.840 ;
        RECT 4.400 159.440 1495.600 160.840 ;
        RECT 2.365 157.440 1497.695 159.440 ;
        RECT 4.400 156.040 1497.695 157.440 ;
        RECT 2.365 154.040 1497.695 156.040 ;
        RECT 4.400 152.640 1495.600 154.040 ;
        RECT 2.365 150.640 1497.695 152.640 ;
        RECT 2.365 149.240 1495.600 150.640 ;
        RECT 2.365 147.240 1497.695 149.240 ;
        RECT 4.400 145.840 1495.600 147.240 ;
        RECT 2.365 143.840 1497.695 145.840 ;
        RECT 4.400 142.440 1495.600 143.840 ;
        RECT 2.365 140.440 1497.695 142.440 ;
        RECT 4.400 139.040 1495.600 140.440 ;
        RECT 2.365 137.040 1497.695 139.040 ;
        RECT 4.400 135.640 1495.600 137.040 ;
        RECT 2.365 133.640 1497.695 135.640 ;
        RECT 4.400 132.240 1497.695 133.640 ;
        RECT 2.365 130.240 1497.695 132.240 ;
        RECT 4.400 128.840 1495.600 130.240 ;
        RECT 2.365 126.840 1497.695 128.840 ;
        RECT 2.365 125.440 1495.600 126.840 ;
        RECT 2.365 123.440 1497.695 125.440 ;
        RECT 4.400 122.040 1495.600 123.440 ;
        RECT 2.365 120.040 1497.695 122.040 ;
        RECT 4.400 118.640 1495.600 120.040 ;
        RECT 2.365 116.640 1497.695 118.640 ;
        RECT 4.400 115.240 1495.600 116.640 ;
        RECT 2.365 113.240 1497.695 115.240 ;
        RECT 4.400 111.840 1495.600 113.240 ;
        RECT 2.365 109.840 1497.695 111.840 ;
        RECT 4.400 108.440 1495.600 109.840 ;
        RECT 2.365 106.440 1497.695 108.440 ;
        RECT 4.400 105.040 1497.695 106.440 ;
        RECT 2.365 103.040 1497.695 105.040 ;
        RECT 4.400 101.640 1495.600 103.040 ;
        RECT 2.365 99.640 1497.695 101.640 ;
        RECT 2.365 98.240 1495.600 99.640 ;
        RECT 2.365 96.240 1497.695 98.240 ;
        RECT 4.400 94.840 1495.600 96.240 ;
        RECT 2.365 92.840 1497.695 94.840 ;
        RECT 4.400 91.440 1495.600 92.840 ;
        RECT 2.365 89.440 1497.695 91.440 ;
        RECT 4.400 88.040 1495.600 89.440 ;
        RECT 2.365 86.040 1497.695 88.040 ;
        RECT 4.400 84.640 1495.600 86.040 ;
        RECT 2.365 82.640 1497.695 84.640 ;
        RECT 4.400 81.240 1497.695 82.640 ;
        RECT 2.365 79.240 1497.695 81.240 ;
        RECT 4.400 77.840 1495.600 79.240 ;
        RECT 2.365 75.840 1497.695 77.840 ;
        RECT 2.365 74.440 1495.600 75.840 ;
        RECT 2.365 72.440 1497.695 74.440 ;
        RECT 4.400 71.040 1495.600 72.440 ;
        RECT 2.365 69.040 1497.695 71.040 ;
        RECT 4.400 67.640 1495.600 69.040 ;
        RECT 2.365 65.640 1497.695 67.640 ;
        RECT 4.400 64.240 1495.600 65.640 ;
        RECT 2.365 62.240 1497.695 64.240 ;
        RECT 4.400 60.840 1495.600 62.240 ;
        RECT 2.365 58.840 1497.695 60.840 ;
        RECT 4.400 57.440 1497.695 58.840 ;
        RECT 2.365 55.440 1497.695 57.440 ;
        RECT 4.400 54.040 1495.600 55.440 ;
        RECT 2.365 52.040 1497.695 54.040 ;
        RECT 4.400 50.640 1495.600 52.040 ;
        RECT 2.365 48.640 1497.695 50.640 ;
        RECT 2.365 47.240 1495.600 48.640 ;
        RECT 2.365 45.240 1497.695 47.240 ;
        RECT 4.400 43.840 1495.600 45.240 ;
        RECT 2.365 41.840 1497.695 43.840 ;
        RECT 4.400 40.440 1495.600 41.840 ;
        RECT 2.365 38.440 1497.695 40.440 ;
        RECT 4.400 37.040 1495.600 38.440 ;
        RECT 2.365 35.040 1497.695 37.040 ;
        RECT 4.400 33.640 1495.600 35.040 ;
        RECT 2.365 31.640 1497.695 33.640 ;
        RECT 4.400 30.240 1497.695 31.640 ;
        RECT 2.365 28.240 1497.695 30.240 ;
        RECT 4.400 26.840 1495.600 28.240 ;
        RECT 2.365 24.840 1497.695 26.840 ;
        RECT 2.365 23.440 1495.600 24.840 ;
        RECT 2.365 21.440 1497.695 23.440 ;
        RECT 4.400 20.040 1495.600 21.440 ;
        RECT 2.365 18.040 1497.695 20.040 ;
        RECT 4.400 16.640 1495.600 18.040 ;
        RECT 2.365 14.640 1497.695 16.640 ;
        RECT 4.400 13.240 1495.600 14.640 ;
        RECT 2.365 11.240 1497.695 13.240 ;
        RECT 4.400 9.840 1495.600 11.240 ;
        RECT 2.365 7.840 1497.695 9.840 ;
        RECT 4.400 6.440 1497.695 7.840 ;
        RECT 2.365 4.440 1497.695 6.440 ;
        RECT 4.400 3.040 1495.600 4.440 ;
        RECT 2.365 1.040 1497.695 3.040 ;
        RECT 2.365 0.175 1495.600 1.040 ;
      LAYER met4 ;
        RECT 3.055 10.240 20.640 1786.185 ;
        RECT 23.040 10.240 97.440 1786.185 ;
        RECT 99.840 10.240 174.240 1786.185 ;
        RECT 176.640 10.240 251.040 1786.185 ;
        RECT 253.440 10.240 327.840 1786.185 ;
        RECT 330.240 10.240 404.640 1786.185 ;
        RECT 407.040 10.240 481.440 1786.185 ;
        RECT 483.840 10.240 558.240 1786.185 ;
        RECT 560.640 10.240 635.040 1786.185 ;
        RECT 637.440 10.240 711.840 1786.185 ;
        RECT 714.240 10.240 788.640 1786.185 ;
        RECT 791.040 10.240 865.440 1786.185 ;
        RECT 867.840 10.240 942.240 1786.185 ;
        RECT 944.640 10.240 1019.040 1786.185 ;
        RECT 1021.440 10.240 1095.840 1786.185 ;
        RECT 1098.240 10.240 1172.640 1786.185 ;
        RECT 1175.040 10.240 1249.440 1786.185 ;
        RECT 1251.840 10.240 1326.240 1786.185 ;
        RECT 1328.640 10.240 1403.040 1786.185 ;
        RECT 1405.440 10.240 1479.840 1786.185 ;
        RECT 1482.240 10.240 1490.105 1786.185 ;
        RECT 3.055 6.975 1490.105 10.240 ;
  END
END mba_core_region
END LIBRARY

