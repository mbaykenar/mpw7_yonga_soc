magic
tech sky130B
magscale 1 2
timestamp 1649977179
<< nwell >>
rect -66 377 2562 897
<< pwell >>
rect 2032 225 2492 301
rect 1598 217 2492 225
rect 4 43 2492 217
rect -26 -43 2522 43
<< locali >>
rect 381 727 612 761
rect 113 500 179 583
rect 381 500 431 727
rect 113 466 431 500
rect 381 461 431 466
rect 217 305 303 430
rect 578 594 612 727
rect 537 560 612 594
rect 537 354 571 560
rect 697 460 769 583
rect 880 460 946 652
rect 1610 583 1858 611
rect 537 289 1084 354
rect 985 162 1084 289
rect 1354 310 1420 504
rect 1562 577 1858 583
rect 1562 384 1644 577
rect 1824 397 1858 577
rect 1824 263 1874 397
rect 2424 121 2474 747
<< obsli1 >>
rect 0 797 31 831
rect 65 797 127 831
rect 161 797 223 831
rect 257 797 319 831
rect 353 797 415 831
rect 449 797 511 831
rect 545 797 607 831
rect 641 797 703 831
rect 737 797 799 831
rect 833 797 895 831
rect 929 797 991 831
rect 1025 797 1087 831
rect 1121 797 1183 831
rect 1217 797 1279 831
rect 1313 797 1375 831
rect 1409 797 1471 831
rect 1505 797 1567 831
rect 1601 797 1663 831
rect 1697 797 1759 831
rect 1793 797 1855 831
rect 1889 797 1951 831
rect 1985 797 2047 831
rect 2081 797 2143 831
rect 2177 797 2239 831
rect 2273 797 2335 831
rect 2369 797 2431 831
rect 2465 797 2496 831
rect 124 735 314 741
rect 22 623 88 715
rect 124 701 130 735
rect 164 701 202 735
rect 236 701 274 735
rect 308 701 314 735
rect 22 269 56 623
rect 124 619 314 701
rect 467 635 542 691
rect 381 269 431 407
rect 22 235 431 269
rect 467 253 501 635
rect 654 735 844 741
rect 654 701 660 735
rect 694 701 732 735
rect 766 701 804 735
rect 838 701 844 735
rect 1266 735 1456 741
rect 654 619 844 701
rect 607 424 657 524
rect 1092 619 1158 719
rect 1266 701 1272 735
rect 1306 701 1344 735
rect 1378 701 1416 735
rect 1450 701 1456 735
rect 1664 727 2174 761
rect 1266 619 1456 701
rect 1492 623 1574 707
rect 1664 647 1730 727
rect 1894 623 1960 691
rect 1124 583 1158 619
rect 1492 583 1526 623
rect 1001 424 1067 583
rect 1124 549 1526 583
rect 607 390 1248 424
rect 22 103 88 235
rect 467 219 910 253
rect 124 113 314 199
rect 124 79 130 113
rect 164 79 202 113
rect 236 79 274 113
rect 308 79 314 113
rect 467 99 542 219
rect 650 113 840 183
rect 124 73 314 79
rect 650 79 656 113
rect 690 79 728 113
rect 762 79 800 113
rect 834 79 840 113
rect 650 73 840 79
rect 876 87 910 219
rect 1182 219 1248 390
rect 1284 183 1318 549
rect 1492 348 1526 549
rect 1492 314 1670 348
rect 1120 123 1318 183
rect 1354 235 1600 269
rect 1354 87 1388 235
rect 876 53 1388 87
rect 1424 113 1530 199
rect 1458 79 1496 113
rect 1424 73 1530 79
rect 1566 87 1600 235
rect 1636 123 1670 314
rect 1910 227 1944 623
rect 1980 531 2030 583
rect 1980 423 2104 531
rect 1706 207 1944 227
rect 1706 193 1998 207
rect 1706 87 1740 193
rect 1566 53 1740 87
rect 1776 87 1842 157
rect 1910 123 1998 193
rect 2054 183 2104 423
rect 2140 385 2174 727
rect 2210 735 2388 751
rect 2244 701 2282 735
rect 2316 701 2354 735
rect 2210 435 2388 701
rect 2140 319 2383 385
rect 2140 87 2174 319
rect 1776 53 2174 87
rect 2210 113 2388 283
rect 2244 79 2282 113
rect 2316 79 2354 113
rect 2210 73 2388 79
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2496 17
<< obsli1c >>
rect 31 797 65 831
rect 127 797 161 831
rect 223 797 257 831
rect 319 797 353 831
rect 415 797 449 831
rect 511 797 545 831
rect 607 797 641 831
rect 703 797 737 831
rect 799 797 833 831
rect 895 797 929 831
rect 991 797 1025 831
rect 1087 797 1121 831
rect 1183 797 1217 831
rect 1279 797 1313 831
rect 1375 797 1409 831
rect 1471 797 1505 831
rect 1567 797 1601 831
rect 1663 797 1697 831
rect 1759 797 1793 831
rect 1855 797 1889 831
rect 1951 797 1985 831
rect 2047 797 2081 831
rect 2143 797 2177 831
rect 2239 797 2273 831
rect 2335 797 2369 831
rect 2431 797 2465 831
rect 130 701 164 735
rect 202 701 236 735
rect 274 701 308 735
rect 660 701 694 735
rect 732 701 766 735
rect 804 701 838 735
rect 1272 701 1306 735
rect 1344 701 1378 735
rect 1416 701 1450 735
rect 130 79 164 113
rect 202 79 236 113
rect 274 79 308 113
rect 656 79 690 113
rect 728 79 762 113
rect 800 79 834 113
rect 1424 79 1458 113
rect 1496 79 1530 113
rect 2210 701 2244 735
rect 2282 701 2316 735
rect 2354 701 2388 735
rect 2210 79 2244 113
rect 2282 79 2316 113
rect 2354 79 2388 113
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
rect 2047 -17 2081 17
rect 2143 -17 2177 17
rect 2239 -17 2273 17
rect 2335 -17 2369 17
rect 2431 -17 2465 17
<< metal1 >>
rect 0 831 2496 837
rect 0 797 31 831
rect 65 797 127 831
rect 161 797 223 831
rect 257 797 319 831
rect 353 797 415 831
rect 449 797 511 831
rect 545 797 607 831
rect 641 797 703 831
rect 737 797 799 831
rect 833 797 895 831
rect 929 797 991 831
rect 1025 797 1087 831
rect 1121 797 1183 831
rect 1217 797 1279 831
rect 1313 797 1375 831
rect 1409 797 1471 831
rect 1505 797 1567 831
rect 1601 797 1663 831
rect 1697 797 1759 831
rect 1793 797 1855 831
rect 1889 797 1951 831
rect 1985 797 2047 831
rect 2081 797 2143 831
rect 2177 797 2239 831
rect 2273 797 2335 831
rect 2369 797 2431 831
rect 2465 797 2496 831
rect 0 791 2496 797
rect 0 735 2496 763
rect 0 701 130 735
rect 164 701 202 735
rect 236 701 274 735
rect 308 701 660 735
rect 694 701 732 735
rect 766 701 804 735
rect 838 701 1272 735
rect 1306 701 1344 735
rect 1378 701 1416 735
rect 1450 701 2210 735
rect 2244 701 2282 735
rect 2316 701 2354 735
rect 2388 701 2496 735
rect 0 689 2496 701
rect 0 113 2496 125
rect 0 79 130 113
rect 164 79 202 113
rect 236 79 274 113
rect 308 79 656 113
rect 690 79 728 113
rect 762 79 800 113
rect 834 79 1424 113
rect 1458 79 1496 113
rect 1530 79 2210 113
rect 2244 79 2282 113
rect 2316 79 2354 113
rect 2388 79 2496 113
rect 0 51 2496 79
rect 0 17 2496 23
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2496 17
rect 0 -23 2496 -17
<< labels >>
rlabel locali s 1354 310 1420 504 6 A0
port 1 nsew signal input
rlabel locali s 880 460 946 652 6 A1
port 2 nsew signal input
rlabel locali s 217 305 303 430 6 A2
port 3 nsew signal input
rlabel locali s 697 460 769 583 6 A3
port 4 nsew signal input
rlabel locali s 985 162 1084 289 6 S0
port 5 nsew signal input
rlabel locali s 537 289 1084 354 6 S0
port 5 nsew signal input
rlabel locali s 537 354 571 560 6 S0
port 5 nsew signal input
rlabel locali s 537 560 612 594 6 S0
port 5 nsew signal input
rlabel locali s 381 461 431 466 6 S0
port 5 nsew signal input
rlabel locali s 113 466 431 500 6 S0
port 5 nsew signal input
rlabel locali s 578 594 612 727 6 S0
port 5 nsew signal input
rlabel locali s 381 500 431 727 6 S0
port 5 nsew signal input
rlabel locali s 113 500 179 583 6 S0
port 5 nsew signal input
rlabel locali s 381 727 612 761 6 S0
port 5 nsew signal input
rlabel locali s 1824 263 1874 397 6 S1
port 6 nsew signal input
rlabel locali s 1824 397 1858 577 6 S1
port 6 nsew signal input
rlabel locali s 1562 384 1644 577 6 S1
port 6 nsew signal input
rlabel locali s 1562 577 1858 583 6 S1
port 6 nsew signal input
rlabel locali s 1610 583 1858 611 6 S1
port 6 nsew signal input
rlabel metal1 s 0 51 2496 125 6 VGND
port 7 nsew ground bidirectional
rlabel metal1 s 0 -23 2496 23 8 VNB
port 8 nsew ground bidirectional
rlabel pwell s -26 -43 2522 43 8 VNB
port 8 nsew ground bidirectional
rlabel pwell s 4 43 2492 217 6 VNB
port 8 nsew ground bidirectional
rlabel pwell s 1598 217 2492 225 6 VNB
port 8 nsew ground bidirectional
rlabel pwell s 2032 225 2492 301 6 VNB
port 8 nsew ground bidirectional
rlabel metal1 s 0 791 2496 837 6 VPB
port 9 nsew power bidirectional
rlabel nwell s -66 377 2562 897 6 VPB
port 9 nsew power bidirectional
rlabel metal1 s 0 689 2496 763 6 VPWR
port 10 nsew power bidirectional
rlabel locali s 2424 121 2474 747 6 X
port 11 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 2496 814
string LEFclass CORE
string LEFsite unithv
string LEFsymmetry X Y
string LEFview TRUE
string GDS_END 236664
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hvl/gds/sky130_fd_sc_hvl.gds
string GDS_START 211614
<< end >>
