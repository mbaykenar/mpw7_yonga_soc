magic
tech sky130B
magscale 12 1
timestamp 1598787603
<< metal5 >>
rect 0 60 60 75
rect 0 30 60 45
<< properties >>
string FIXED_BBOX 0 -30 75 105
<< end >>
