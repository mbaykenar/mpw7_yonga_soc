magic
tech sky130A
magscale 1 2
timestamp 1649977179
<< nwell >>
rect -38 261 682 582
<< pwell >>
rect 370 157 643 203
rect 1 21 643 157
rect 30 -17 64 21
<< scnmos >>
rect 79 47 109 131
rect 267 47 297 131
rect 351 47 381 131
rect 449 47 479 177
rect 533 47 563 177
<< scpmoshvt >>
rect 79 413 109 497
rect 182 413 212 497
rect 270 413 300 497
rect 449 297 479 497
rect 533 297 563 497
<< ndiff >>
rect 396 131 449 177
rect 27 106 79 131
rect 27 72 35 106
rect 69 72 79 106
rect 27 47 79 72
rect 109 106 161 131
rect 109 72 119 106
rect 153 72 161 106
rect 109 47 161 72
rect 215 106 267 131
rect 215 72 223 106
rect 257 72 267 106
rect 215 47 267 72
rect 297 47 351 131
rect 381 111 449 131
rect 381 77 405 111
rect 439 77 449 111
rect 381 47 449 77
rect 479 127 533 177
rect 479 93 489 127
rect 523 93 533 127
rect 479 47 533 93
rect 563 127 617 177
rect 563 93 573 127
rect 607 93 617 127
rect 563 47 617 93
<< pdiff >>
rect 27 462 79 497
rect 27 428 35 462
rect 69 428 79 462
rect 27 413 79 428
rect 109 471 182 497
rect 109 437 119 471
rect 153 437 182 471
rect 109 413 182 437
rect 212 462 270 497
rect 212 428 224 462
rect 258 428 270 462
rect 212 413 270 428
rect 300 483 449 497
rect 300 449 320 483
rect 354 449 388 483
rect 422 449 449 483
rect 300 413 449 449
rect 399 297 449 413
rect 479 457 533 497
rect 479 423 489 457
rect 523 423 533 457
rect 479 384 533 423
rect 479 350 489 384
rect 523 350 533 384
rect 479 297 533 350
rect 563 457 615 497
rect 563 423 573 457
rect 607 423 615 457
rect 563 389 615 423
rect 563 355 573 389
rect 607 355 615 389
rect 563 297 615 355
<< ndiffc >>
rect 35 72 69 106
rect 119 72 153 106
rect 223 72 257 106
rect 405 77 439 111
rect 489 93 523 127
rect 573 93 607 127
<< pdiffc >>
rect 35 428 69 462
rect 119 437 153 471
rect 224 428 258 462
rect 320 449 354 483
rect 388 449 422 483
rect 489 423 523 457
rect 489 350 523 384
rect 573 423 607 457
rect 573 355 607 389
<< poly >>
rect 79 497 109 523
rect 182 497 212 523
rect 270 497 300 523
rect 449 497 479 523
rect 533 497 563 523
rect 79 265 109 413
rect 40 249 109 265
rect 40 215 56 249
rect 90 215 109 249
rect 40 199 109 215
rect 79 131 109 199
rect 182 227 212 413
rect 270 379 300 413
rect 270 363 368 379
rect 270 329 317 363
rect 351 329 368 363
rect 270 305 368 329
rect 294 282 368 305
rect 294 233 381 282
rect 449 265 479 297
rect 533 265 563 297
rect 182 211 251 227
rect 182 177 201 211
rect 235 191 251 211
rect 235 177 297 191
rect 182 161 297 177
rect 267 131 297 161
rect 351 131 381 233
rect 423 249 563 265
rect 423 215 433 249
rect 467 215 563 249
rect 423 197 563 215
rect 449 177 479 197
rect 533 177 563 197
rect 79 21 109 47
rect 267 21 297 47
rect 351 21 381 47
rect 449 21 479 47
rect 533 21 563 47
<< polycont >>
rect 56 215 90 249
rect 317 329 351 363
rect 201 177 235 211
rect 433 215 467 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 644 561
rect 35 462 69 489
rect 103 471 169 527
rect 103 437 119 471
rect 153 437 169 471
rect 209 462 266 484
rect 35 403 69 428
rect 209 428 224 462
rect 258 428 266 462
rect 302 483 439 527
rect 302 449 320 483
rect 354 449 388 483
rect 422 449 439 483
rect 302 433 439 449
rect 475 457 536 473
rect 35 357 171 403
rect 30 249 90 323
rect 30 215 56 249
rect 30 153 90 215
rect 124 227 171 357
rect 209 295 266 428
rect 475 423 489 457
rect 523 423 536 457
rect 301 363 440 391
rect 301 329 317 363
rect 351 329 440 363
rect 475 384 536 423
rect 475 350 489 384
rect 523 350 536 384
rect 475 316 536 350
rect 573 457 627 527
rect 607 423 627 457
rect 573 389 627 423
rect 607 355 627 389
rect 573 336 627 355
rect 209 265 381 295
rect 209 261 467 265
rect 269 249 467 261
rect 124 211 235 227
rect 124 177 201 211
rect 124 161 235 177
rect 269 215 433 249
rect 269 189 467 215
rect 124 131 167 161
rect 19 106 85 118
rect 19 72 35 106
rect 69 72 85 106
rect 19 17 85 72
rect 119 106 167 131
rect 269 122 303 189
rect 501 155 536 316
rect 153 72 167 106
rect 119 56 167 72
rect 223 106 303 122
rect 489 127 536 155
rect 257 83 303 106
rect 375 111 455 116
rect 223 54 257 72
rect 375 77 405 111
rect 439 77 455 111
rect 375 17 455 77
rect 523 93 536 127
rect 489 51 536 93
rect 573 127 627 144
rect 607 93 627 127
rect 573 17 627 93
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 644 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
<< metal1 >>
rect 0 561 644 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 644 561
rect 0 496 644 527
rect 0 17 644 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 644 17
rect 0 -48 644 -17
<< labels >>
flabel pwell s 30 -17 64 17 0 FreeSans 200 0 0 0 VNB
port 4 nsew ground bidirectional
flabel nwell s 30 527 64 561 0 FreeSans 200 0 0 0 VPB
port 5 nsew power bidirectional
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 6 nsew power bidirectional abutment
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 3 nsew ground bidirectional abutment
flabel locali s 494 425 528 459 0 FreeSans 200 0 0 0 X
port 7 nsew signal output
flabel locali s 301 329 440 391 0 FreeSans 400 0 0 0 B
port 2 nsew signal input
flabel locali s 30 153 90 323 0 FreeSans 400 0 0 0 A_N
port 1 nsew signal input
flabel locali s 511 102 511 102 0 FreeSans 200 0 0 0 X
port 7 nsew
flabel locali s 310 357 344 391 0 FreeSans 400 0 0 0 B
port 2 nsew
flabel locali s 46 170 46 170 0 FreeSans 400 0 0 0 A_N
port 1 nsew
flabel locali s 30 289 64 323 0 FreeSans 400 0 0 0 A_N
port 1 nsew
flabel locali s 511 374 511 374 0 FreeSans 200 0 0 0 X
port 7 nsew
rlabel comment s 0 0 0 0 4 and2b_2
rlabel metal1 s 0 -48 644 48 1 VGND
port 3 nsew ground bidirectional abutment
rlabel metal1 s 0 496 644 592 1 VPWR
port 6 nsew power bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 644 544
string GDS_END 3839880
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 3834276
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string path 0.000 0.000 16.100 0.000 
<< end >>
