* NGSPICE file created from sky130_ef_sc_hd__fill_4.ext - technology: sky130A

.subckt sky130_ef_sc_hd__fill_4 VGND VPWR VPB VNB
.ends

