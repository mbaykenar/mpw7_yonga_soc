magic
tech sky130B
magscale 1 2
timestamp 1649977179
<< locali >>
rect 110 266 176 300
rect 0 176 66 210
rect 110 64 176 98
rect 1372 88 1406 170
rect 1477 103 2054 137
rect 767 54 1406 88
<< metal1 >>
rect 248 -44 294 418
rect 672 14 720 418
rect 1104 14 1152 418
rect 1496 0 1524 395
rect 1892 0 1920 395
use sky130_fd_bd_sram__openram_dp_nand3_dec_2  sky130_fd_bd_sram__openram_dp_nand3_dec_0
timestamp 1649977179
transform 1 0 0 0 1 0
box 0 -60 1322 474
use sky130_sram_1kbyte_1rw1r_8x1024_8_pinv_dec  sky130_sram_1kbyte_1rw1r_8x1024_8_pinv_dec_0
timestamp 1649977179
transform 1 0 1312 0 1 0
box 44 0 760 490
<< labels >>
rlabel metal1 s 1104 14 1152 418 4 vdd
port 1 nsew
rlabel metal1 s 672 14 720 418 4 vdd
port 1 nsew
rlabel metal1 s 1892 0 1920 395 4 vdd
port 1 nsew
rlabel metal1 s 1496 0 1524 395 4 gnd
port 2 nsew
rlabel metal1 s 248 -44 294 418 4 gnd
port 2 nsew
rlabel locali s 1765 120 1765 120 4 Z
port 3 nsew
rlabel locali s 143 81 143 81 4 A
port 4 nsew
rlabel locali s 33 193 33 193 4 B
port 5 nsew
rlabel locali s 143 283 143 283 4 C
port 6 nsew
<< properties >>
string FIXED_BBOX 0 0 2054 395
string GDS_END 51814
string GDS_FILE $PDKPATH/libs.ref/sky130_sram_macros/gds/sky130_sram_1kbyte_1rw1r_8x1024_8.gds
string GDS_START 50046
<< end >>
