magic
tech sky130B
magscale 1 2
timestamp 1662563211
<< obsli1 >>
rect 1104 2159 138828 437393
<< obsm1 >>
rect 14 1368 139992 437424
<< metal2 >>
rect 18 439200 74 440000
rect 662 439200 718 440000
rect 1950 439200 2006 440000
rect 2594 439200 2650 440000
rect 3238 439200 3294 440000
rect 3882 439200 3938 440000
rect 4526 439200 4582 440000
rect 5814 439200 5870 440000
rect 6458 439200 6514 440000
rect 7102 439200 7158 440000
rect 7746 439200 7802 440000
rect 8390 439200 8446 440000
rect 9034 439200 9090 440000
rect 10322 439200 10378 440000
rect 10966 439200 11022 440000
rect 11610 439200 11666 440000
rect 12254 439200 12310 440000
rect 12898 439200 12954 440000
rect 14186 439200 14242 440000
rect 14830 439200 14886 440000
rect 15474 439200 15530 440000
rect 16118 439200 16174 440000
rect 16762 439200 16818 440000
rect 18050 439200 18106 440000
rect 18694 439200 18750 440000
rect 19338 439200 19394 440000
rect 19982 439200 20038 440000
rect 20626 439200 20682 440000
rect 21914 439200 21970 440000
rect 22558 439200 22614 440000
rect 23202 439200 23258 440000
rect 23846 439200 23902 440000
rect 24490 439200 24546 440000
rect 25134 439200 25190 440000
rect 26422 439200 26478 440000
rect 27066 439200 27122 440000
rect 27710 439200 27766 440000
rect 28354 439200 28410 440000
rect 28998 439200 29054 440000
rect 30286 439200 30342 440000
rect 30930 439200 30986 440000
rect 31574 439200 31630 440000
rect 32218 439200 32274 440000
rect 32862 439200 32918 440000
rect 34150 439200 34206 440000
rect 34794 439200 34850 440000
rect 35438 439200 35494 440000
rect 36082 439200 36138 440000
rect 36726 439200 36782 440000
rect 38014 439200 38070 440000
rect 38658 439200 38714 440000
rect 39302 439200 39358 440000
rect 39946 439200 40002 440000
rect 40590 439200 40646 440000
rect 41878 439200 41934 440000
rect 42522 439200 42578 440000
rect 43166 439200 43222 440000
rect 43810 439200 43866 440000
rect 44454 439200 44510 440000
rect 45098 439200 45154 440000
rect 46386 439200 46442 440000
rect 47030 439200 47086 440000
rect 47674 439200 47730 440000
rect 48318 439200 48374 440000
rect 48962 439200 49018 440000
rect 50250 439200 50306 440000
rect 50894 439200 50950 440000
rect 51538 439200 51594 440000
rect 52182 439200 52238 440000
rect 52826 439200 52882 440000
rect 54114 439200 54170 440000
rect 54758 439200 54814 440000
rect 55402 439200 55458 440000
rect 56046 439200 56102 440000
rect 56690 439200 56746 440000
rect 57978 439200 58034 440000
rect 58622 439200 58678 440000
rect 59266 439200 59322 440000
rect 59910 439200 59966 440000
rect 60554 439200 60610 440000
rect 61198 439200 61254 440000
rect 62486 439200 62542 440000
rect 63130 439200 63186 440000
rect 63774 439200 63830 440000
rect 64418 439200 64474 440000
rect 65062 439200 65118 440000
rect 66350 439200 66406 440000
rect 66994 439200 67050 440000
rect 67638 439200 67694 440000
rect 68282 439200 68338 440000
rect 68926 439200 68982 440000
rect 70214 439200 70270 440000
rect 70858 439200 70914 440000
rect 71502 439200 71558 440000
rect 72146 439200 72202 440000
rect 72790 439200 72846 440000
rect 74078 439200 74134 440000
rect 74722 439200 74778 440000
rect 75366 439200 75422 440000
rect 76010 439200 76066 440000
rect 76654 439200 76710 440000
rect 77298 439200 77354 440000
rect 78586 439200 78642 440000
rect 79230 439200 79286 440000
rect 79874 439200 79930 440000
rect 80518 439200 80574 440000
rect 81162 439200 81218 440000
rect 82450 439200 82506 440000
rect 83094 439200 83150 440000
rect 83738 439200 83794 440000
rect 84382 439200 84438 440000
rect 85026 439200 85082 440000
rect 86314 439200 86370 440000
rect 86958 439200 87014 440000
rect 87602 439200 87658 440000
rect 88246 439200 88302 440000
rect 88890 439200 88946 440000
rect 90178 439200 90234 440000
rect 90822 439200 90878 440000
rect 91466 439200 91522 440000
rect 92110 439200 92166 440000
rect 92754 439200 92810 440000
rect 93398 439200 93454 440000
rect 94686 439200 94742 440000
rect 95330 439200 95386 440000
rect 95974 439200 96030 440000
rect 96618 439200 96674 440000
rect 97262 439200 97318 440000
rect 98550 439200 98606 440000
rect 99194 439200 99250 440000
rect 99838 439200 99894 440000
rect 100482 439200 100538 440000
rect 101126 439200 101182 440000
rect 102414 439200 102470 440000
rect 103058 439200 103114 440000
rect 103702 439200 103758 440000
rect 104346 439200 104402 440000
rect 104990 439200 105046 440000
rect 106278 439200 106334 440000
rect 106922 439200 106978 440000
rect 107566 439200 107622 440000
rect 108210 439200 108266 440000
rect 108854 439200 108910 440000
rect 109498 439200 109554 440000
rect 110786 439200 110842 440000
rect 111430 439200 111486 440000
rect 112074 439200 112130 440000
rect 112718 439200 112774 440000
rect 113362 439200 113418 440000
rect 114650 439200 114706 440000
rect 115294 439200 115350 440000
rect 115938 439200 115994 440000
rect 116582 439200 116638 440000
rect 117226 439200 117282 440000
rect 118514 439200 118570 440000
rect 119158 439200 119214 440000
rect 119802 439200 119858 440000
rect 120446 439200 120502 440000
rect 121090 439200 121146 440000
rect 122378 439200 122434 440000
rect 123022 439200 123078 440000
rect 123666 439200 123722 440000
rect 124310 439200 124366 440000
rect 124954 439200 125010 440000
rect 125598 439200 125654 440000
rect 126886 439200 126942 440000
rect 127530 439200 127586 440000
rect 128174 439200 128230 440000
rect 128818 439200 128874 440000
rect 129462 439200 129518 440000
rect 130750 439200 130806 440000
rect 131394 439200 131450 440000
rect 132038 439200 132094 440000
rect 132682 439200 132738 440000
rect 133326 439200 133382 440000
rect 134614 439200 134670 440000
rect 135258 439200 135314 440000
rect 135902 439200 135958 440000
rect 136546 439200 136602 440000
rect 137190 439200 137246 440000
rect 138478 439200 138534 440000
rect 139122 439200 139178 440000
rect 139766 439200 139822 440000
rect 18 0 74 800
rect 662 0 718 800
rect 1306 0 1362 800
rect 1950 0 2006 800
rect 2594 0 2650 800
rect 3238 0 3294 800
rect 4526 0 4582 800
rect 5170 0 5226 800
rect 5814 0 5870 800
rect 6458 0 6514 800
rect 7102 0 7158 800
rect 8390 0 8446 800
rect 9034 0 9090 800
rect 9678 0 9734 800
rect 10322 0 10378 800
rect 10966 0 11022 800
rect 12254 0 12310 800
rect 12898 0 12954 800
rect 13542 0 13598 800
rect 14186 0 14242 800
rect 14830 0 14886 800
rect 16118 0 16174 800
rect 16762 0 16818 800
rect 17406 0 17462 800
rect 18050 0 18106 800
rect 18694 0 18750 800
rect 19338 0 19394 800
rect 20626 0 20682 800
rect 21270 0 21326 800
rect 21914 0 21970 800
rect 22558 0 22614 800
rect 23202 0 23258 800
rect 24490 0 24546 800
rect 25134 0 25190 800
rect 25778 0 25834 800
rect 26422 0 26478 800
rect 27066 0 27122 800
rect 28354 0 28410 800
rect 28998 0 29054 800
rect 29642 0 29698 800
rect 30286 0 30342 800
rect 30930 0 30986 800
rect 32218 0 32274 800
rect 32862 0 32918 800
rect 33506 0 33562 800
rect 34150 0 34206 800
rect 34794 0 34850 800
rect 35438 0 35494 800
rect 36726 0 36782 800
rect 37370 0 37426 800
rect 38014 0 38070 800
rect 38658 0 38714 800
rect 39302 0 39358 800
rect 40590 0 40646 800
rect 41234 0 41290 800
rect 41878 0 41934 800
rect 42522 0 42578 800
rect 43166 0 43222 800
rect 44454 0 44510 800
rect 45098 0 45154 800
rect 45742 0 45798 800
rect 46386 0 46442 800
rect 47030 0 47086 800
rect 48318 0 48374 800
rect 48962 0 49018 800
rect 49606 0 49662 800
rect 50250 0 50306 800
rect 50894 0 50950 800
rect 51538 0 51594 800
rect 52826 0 52882 800
rect 53470 0 53526 800
rect 54114 0 54170 800
rect 54758 0 54814 800
rect 55402 0 55458 800
rect 56690 0 56746 800
rect 57334 0 57390 800
rect 57978 0 58034 800
rect 58622 0 58678 800
rect 59266 0 59322 800
rect 60554 0 60610 800
rect 61198 0 61254 800
rect 61842 0 61898 800
rect 62486 0 62542 800
rect 63130 0 63186 800
rect 64418 0 64474 800
rect 65062 0 65118 800
rect 65706 0 65762 800
rect 66350 0 66406 800
rect 66994 0 67050 800
rect 67638 0 67694 800
rect 68926 0 68982 800
rect 69570 0 69626 800
rect 70214 0 70270 800
rect 70858 0 70914 800
rect 71502 0 71558 800
rect 72790 0 72846 800
rect 73434 0 73490 800
rect 74078 0 74134 800
rect 74722 0 74778 800
rect 75366 0 75422 800
rect 76654 0 76710 800
rect 77298 0 77354 800
rect 77942 0 77998 800
rect 78586 0 78642 800
rect 79230 0 79286 800
rect 80518 0 80574 800
rect 81162 0 81218 800
rect 81806 0 81862 800
rect 82450 0 82506 800
rect 83094 0 83150 800
rect 83738 0 83794 800
rect 85026 0 85082 800
rect 85670 0 85726 800
rect 86314 0 86370 800
rect 86958 0 87014 800
rect 87602 0 87658 800
rect 88890 0 88946 800
rect 89534 0 89590 800
rect 90178 0 90234 800
rect 90822 0 90878 800
rect 91466 0 91522 800
rect 92754 0 92810 800
rect 93398 0 93454 800
rect 94042 0 94098 800
rect 94686 0 94742 800
rect 95330 0 95386 800
rect 96618 0 96674 800
rect 97262 0 97318 800
rect 97906 0 97962 800
rect 98550 0 98606 800
rect 99194 0 99250 800
rect 99838 0 99894 800
rect 101126 0 101182 800
rect 101770 0 101826 800
rect 102414 0 102470 800
rect 103058 0 103114 800
rect 103702 0 103758 800
rect 104990 0 105046 800
rect 105634 0 105690 800
rect 106278 0 106334 800
rect 106922 0 106978 800
rect 107566 0 107622 800
rect 108854 0 108910 800
rect 109498 0 109554 800
rect 110142 0 110198 800
rect 110786 0 110842 800
rect 111430 0 111486 800
rect 112718 0 112774 800
rect 113362 0 113418 800
rect 114006 0 114062 800
rect 114650 0 114706 800
rect 115294 0 115350 800
rect 115938 0 115994 800
rect 117226 0 117282 800
rect 117870 0 117926 800
rect 118514 0 118570 800
rect 119158 0 119214 800
rect 119802 0 119858 800
rect 121090 0 121146 800
rect 121734 0 121790 800
rect 122378 0 122434 800
rect 123022 0 123078 800
rect 123666 0 123722 800
rect 124954 0 125010 800
rect 125598 0 125654 800
rect 126242 0 126298 800
rect 126886 0 126942 800
rect 127530 0 127586 800
rect 128818 0 128874 800
rect 129462 0 129518 800
rect 130106 0 130162 800
rect 130750 0 130806 800
rect 131394 0 131450 800
rect 132038 0 132094 800
rect 133326 0 133382 800
rect 133970 0 134026 800
rect 134614 0 134670 800
rect 135258 0 135314 800
rect 135902 0 135958 800
rect 137190 0 137246 800
rect 137834 0 137890 800
rect 138478 0 138534 800
rect 139122 0 139178 800
rect 139766 0 139822 800
<< obsm2 >>
rect 130 439144 606 439385
rect 774 439144 1894 439385
rect 2062 439144 2538 439385
rect 2706 439144 3182 439385
rect 3350 439144 3826 439385
rect 3994 439144 4470 439385
rect 4638 439144 5758 439385
rect 5926 439144 6402 439385
rect 6570 439144 7046 439385
rect 7214 439144 7690 439385
rect 7858 439144 8334 439385
rect 8502 439144 8978 439385
rect 9146 439144 10266 439385
rect 10434 439144 10910 439385
rect 11078 439144 11554 439385
rect 11722 439144 12198 439385
rect 12366 439144 12842 439385
rect 13010 439144 14130 439385
rect 14298 439144 14774 439385
rect 14942 439144 15418 439385
rect 15586 439144 16062 439385
rect 16230 439144 16706 439385
rect 16874 439144 17994 439385
rect 18162 439144 18638 439385
rect 18806 439144 19282 439385
rect 19450 439144 19926 439385
rect 20094 439144 20570 439385
rect 20738 439144 21858 439385
rect 22026 439144 22502 439385
rect 22670 439144 23146 439385
rect 23314 439144 23790 439385
rect 23958 439144 24434 439385
rect 24602 439144 25078 439385
rect 25246 439144 26366 439385
rect 26534 439144 27010 439385
rect 27178 439144 27654 439385
rect 27822 439144 28298 439385
rect 28466 439144 28942 439385
rect 29110 439144 30230 439385
rect 30398 439144 30874 439385
rect 31042 439144 31518 439385
rect 31686 439144 32162 439385
rect 32330 439144 32806 439385
rect 32974 439144 34094 439385
rect 34262 439144 34738 439385
rect 34906 439144 35382 439385
rect 35550 439144 36026 439385
rect 36194 439144 36670 439385
rect 36838 439144 37958 439385
rect 38126 439144 38602 439385
rect 38770 439144 39246 439385
rect 39414 439144 39890 439385
rect 40058 439144 40534 439385
rect 40702 439144 41822 439385
rect 41990 439144 42466 439385
rect 42634 439144 43110 439385
rect 43278 439144 43754 439385
rect 43922 439144 44398 439385
rect 44566 439144 45042 439385
rect 45210 439144 46330 439385
rect 46498 439144 46974 439385
rect 47142 439144 47618 439385
rect 47786 439144 48262 439385
rect 48430 439144 48906 439385
rect 49074 439144 50194 439385
rect 50362 439144 50838 439385
rect 51006 439144 51482 439385
rect 51650 439144 52126 439385
rect 52294 439144 52770 439385
rect 52938 439144 54058 439385
rect 54226 439144 54702 439385
rect 54870 439144 55346 439385
rect 55514 439144 55990 439385
rect 56158 439144 56634 439385
rect 56802 439144 57922 439385
rect 58090 439144 58566 439385
rect 58734 439144 59210 439385
rect 59378 439144 59854 439385
rect 60022 439144 60498 439385
rect 60666 439144 61142 439385
rect 61310 439144 62430 439385
rect 62598 439144 63074 439385
rect 63242 439144 63718 439385
rect 63886 439144 64362 439385
rect 64530 439144 65006 439385
rect 65174 439144 66294 439385
rect 66462 439144 66938 439385
rect 67106 439144 67582 439385
rect 67750 439144 68226 439385
rect 68394 439144 68870 439385
rect 69038 439144 70158 439385
rect 70326 439144 70802 439385
rect 70970 439144 71446 439385
rect 71614 439144 72090 439385
rect 72258 439144 72734 439385
rect 72902 439144 74022 439385
rect 74190 439144 74666 439385
rect 74834 439144 75310 439385
rect 75478 439144 75954 439385
rect 76122 439144 76598 439385
rect 76766 439144 77242 439385
rect 77410 439144 78530 439385
rect 78698 439144 79174 439385
rect 79342 439144 79818 439385
rect 79986 439144 80462 439385
rect 80630 439144 81106 439385
rect 81274 439144 82394 439385
rect 82562 439144 83038 439385
rect 83206 439144 83682 439385
rect 83850 439144 84326 439385
rect 84494 439144 84970 439385
rect 85138 439144 86258 439385
rect 86426 439144 86902 439385
rect 87070 439144 87546 439385
rect 87714 439144 88190 439385
rect 88358 439144 88834 439385
rect 89002 439144 90122 439385
rect 90290 439144 90766 439385
rect 90934 439144 91410 439385
rect 91578 439144 92054 439385
rect 92222 439144 92698 439385
rect 92866 439144 93342 439385
rect 93510 439144 94630 439385
rect 94798 439144 95274 439385
rect 95442 439144 95918 439385
rect 96086 439144 96562 439385
rect 96730 439144 97206 439385
rect 97374 439144 98494 439385
rect 98662 439144 99138 439385
rect 99306 439144 99782 439385
rect 99950 439144 100426 439385
rect 100594 439144 101070 439385
rect 101238 439144 102358 439385
rect 102526 439144 103002 439385
rect 103170 439144 103646 439385
rect 103814 439144 104290 439385
rect 104458 439144 104934 439385
rect 105102 439144 106222 439385
rect 106390 439144 106866 439385
rect 107034 439144 107510 439385
rect 107678 439144 108154 439385
rect 108322 439144 108798 439385
rect 108966 439144 109442 439385
rect 109610 439144 110730 439385
rect 110898 439144 111374 439385
rect 111542 439144 112018 439385
rect 112186 439144 112662 439385
rect 112830 439144 113306 439385
rect 113474 439144 114594 439385
rect 114762 439144 115238 439385
rect 115406 439144 115882 439385
rect 116050 439144 116526 439385
rect 116694 439144 117170 439385
rect 117338 439144 118458 439385
rect 118626 439144 119102 439385
rect 119270 439144 119746 439385
rect 119914 439144 120390 439385
rect 120558 439144 121034 439385
rect 121202 439144 122322 439385
rect 122490 439144 122966 439385
rect 123134 439144 123610 439385
rect 123778 439144 124254 439385
rect 124422 439144 124898 439385
rect 125066 439144 125542 439385
rect 125710 439144 126830 439385
rect 126998 439144 127474 439385
rect 127642 439144 128118 439385
rect 128286 439144 128762 439385
rect 128930 439144 129406 439385
rect 129574 439144 130694 439385
rect 130862 439144 131338 439385
rect 131506 439144 131982 439385
rect 132150 439144 132626 439385
rect 132794 439144 133270 439385
rect 133438 439144 134558 439385
rect 134726 439144 135202 439385
rect 135370 439144 135846 439385
rect 136014 439144 136490 439385
rect 136658 439144 137134 439385
rect 137302 439144 138422 439385
rect 138590 439144 139066 439385
rect 139234 439144 139710 439385
rect 139878 439144 139992 439385
rect 20 856 139992 439144
rect 130 711 606 856
rect 774 711 1250 856
rect 1418 711 1894 856
rect 2062 711 2538 856
rect 2706 711 3182 856
rect 3350 711 4470 856
rect 4638 711 5114 856
rect 5282 711 5758 856
rect 5926 711 6402 856
rect 6570 711 7046 856
rect 7214 711 8334 856
rect 8502 711 8978 856
rect 9146 711 9622 856
rect 9790 711 10266 856
rect 10434 711 10910 856
rect 11078 711 12198 856
rect 12366 711 12842 856
rect 13010 711 13486 856
rect 13654 711 14130 856
rect 14298 711 14774 856
rect 14942 711 16062 856
rect 16230 711 16706 856
rect 16874 711 17350 856
rect 17518 711 17994 856
rect 18162 711 18638 856
rect 18806 711 19282 856
rect 19450 711 20570 856
rect 20738 711 21214 856
rect 21382 711 21858 856
rect 22026 711 22502 856
rect 22670 711 23146 856
rect 23314 711 24434 856
rect 24602 711 25078 856
rect 25246 711 25722 856
rect 25890 711 26366 856
rect 26534 711 27010 856
rect 27178 711 28298 856
rect 28466 711 28942 856
rect 29110 711 29586 856
rect 29754 711 30230 856
rect 30398 711 30874 856
rect 31042 711 32162 856
rect 32330 711 32806 856
rect 32974 711 33450 856
rect 33618 711 34094 856
rect 34262 711 34738 856
rect 34906 711 35382 856
rect 35550 711 36670 856
rect 36838 711 37314 856
rect 37482 711 37958 856
rect 38126 711 38602 856
rect 38770 711 39246 856
rect 39414 711 40534 856
rect 40702 711 41178 856
rect 41346 711 41822 856
rect 41990 711 42466 856
rect 42634 711 43110 856
rect 43278 711 44398 856
rect 44566 711 45042 856
rect 45210 711 45686 856
rect 45854 711 46330 856
rect 46498 711 46974 856
rect 47142 711 48262 856
rect 48430 711 48906 856
rect 49074 711 49550 856
rect 49718 711 50194 856
rect 50362 711 50838 856
rect 51006 711 51482 856
rect 51650 711 52770 856
rect 52938 711 53414 856
rect 53582 711 54058 856
rect 54226 711 54702 856
rect 54870 711 55346 856
rect 55514 711 56634 856
rect 56802 711 57278 856
rect 57446 711 57922 856
rect 58090 711 58566 856
rect 58734 711 59210 856
rect 59378 711 60498 856
rect 60666 711 61142 856
rect 61310 711 61786 856
rect 61954 711 62430 856
rect 62598 711 63074 856
rect 63242 711 64362 856
rect 64530 711 65006 856
rect 65174 711 65650 856
rect 65818 711 66294 856
rect 66462 711 66938 856
rect 67106 711 67582 856
rect 67750 711 68870 856
rect 69038 711 69514 856
rect 69682 711 70158 856
rect 70326 711 70802 856
rect 70970 711 71446 856
rect 71614 711 72734 856
rect 72902 711 73378 856
rect 73546 711 74022 856
rect 74190 711 74666 856
rect 74834 711 75310 856
rect 75478 711 76598 856
rect 76766 711 77242 856
rect 77410 711 77886 856
rect 78054 711 78530 856
rect 78698 711 79174 856
rect 79342 711 80462 856
rect 80630 711 81106 856
rect 81274 711 81750 856
rect 81918 711 82394 856
rect 82562 711 83038 856
rect 83206 711 83682 856
rect 83850 711 84970 856
rect 85138 711 85614 856
rect 85782 711 86258 856
rect 86426 711 86902 856
rect 87070 711 87546 856
rect 87714 711 88834 856
rect 89002 711 89478 856
rect 89646 711 90122 856
rect 90290 711 90766 856
rect 90934 711 91410 856
rect 91578 711 92698 856
rect 92866 711 93342 856
rect 93510 711 93986 856
rect 94154 711 94630 856
rect 94798 711 95274 856
rect 95442 711 96562 856
rect 96730 711 97206 856
rect 97374 711 97850 856
rect 98018 711 98494 856
rect 98662 711 99138 856
rect 99306 711 99782 856
rect 99950 711 101070 856
rect 101238 711 101714 856
rect 101882 711 102358 856
rect 102526 711 103002 856
rect 103170 711 103646 856
rect 103814 711 104934 856
rect 105102 711 105578 856
rect 105746 711 106222 856
rect 106390 711 106866 856
rect 107034 711 107510 856
rect 107678 711 108798 856
rect 108966 711 109442 856
rect 109610 711 110086 856
rect 110254 711 110730 856
rect 110898 711 111374 856
rect 111542 711 112662 856
rect 112830 711 113306 856
rect 113474 711 113950 856
rect 114118 711 114594 856
rect 114762 711 115238 856
rect 115406 711 115882 856
rect 116050 711 117170 856
rect 117338 711 117814 856
rect 117982 711 118458 856
rect 118626 711 119102 856
rect 119270 711 119746 856
rect 119914 711 121034 856
rect 121202 711 121678 856
rect 121846 711 122322 856
rect 122490 711 122966 856
rect 123134 711 123610 856
rect 123778 711 124898 856
rect 125066 711 125542 856
rect 125710 711 126186 856
rect 126354 711 126830 856
rect 126998 711 127474 856
rect 127642 711 128762 856
rect 128930 711 129406 856
rect 129574 711 130050 856
rect 130218 711 130694 856
rect 130862 711 131338 856
rect 131506 711 131982 856
rect 132150 711 133270 856
rect 133438 711 133914 856
rect 134082 711 134558 856
rect 134726 711 135202 856
rect 135370 711 135846 856
rect 136014 711 137134 856
rect 137302 711 137778 856
rect 137946 711 138422 856
rect 138590 711 139066 856
rect 139234 711 139710 856
rect 139878 711 139992 856
<< metal3 >>
rect 0 439288 800 439408
rect 139200 439288 140000 439408
rect 0 438608 800 438728
rect 139200 438608 140000 438728
rect 0 437928 800 438048
rect 139200 437928 140000 438048
rect 0 436568 800 436688
rect 139200 436568 140000 436688
rect 0 435888 800 436008
rect 139200 435888 140000 436008
rect 0 435208 800 435328
rect 139200 435208 140000 435328
rect 0 434528 800 434648
rect 139200 434528 140000 434648
rect 0 433848 800 433968
rect 139200 433848 140000 433968
rect 0 432488 800 432608
rect 139200 432488 140000 432608
rect 0 431808 800 431928
rect 139200 431808 140000 431928
rect 0 431128 800 431248
rect 139200 431128 140000 431248
rect 0 430448 800 430568
rect 139200 430448 140000 430568
rect 0 429768 800 429888
rect 139200 429768 140000 429888
rect 0 429088 800 429208
rect 139200 428408 140000 428528
rect 0 427728 800 427848
rect 139200 427728 140000 427848
rect 0 427048 800 427168
rect 139200 427048 140000 427168
rect 0 426368 800 426488
rect 139200 426368 140000 426488
rect 0 425688 800 425808
rect 139200 425688 140000 425808
rect 0 425008 800 425128
rect 139200 424328 140000 424448
rect 0 423648 800 423768
rect 139200 423648 140000 423768
rect 0 422968 800 423088
rect 139200 422968 140000 423088
rect 0 422288 800 422408
rect 139200 422288 140000 422408
rect 0 421608 800 421728
rect 139200 421608 140000 421728
rect 0 420928 800 421048
rect 139200 420928 140000 421048
rect 0 419568 800 419688
rect 139200 419568 140000 419688
rect 0 418888 800 419008
rect 139200 418888 140000 419008
rect 0 418208 800 418328
rect 139200 418208 140000 418328
rect 0 417528 800 417648
rect 139200 417528 140000 417648
rect 0 416848 800 416968
rect 139200 416848 140000 416968
rect 0 415488 800 415608
rect 139200 415488 140000 415608
rect 0 414808 800 414928
rect 139200 414808 140000 414928
rect 0 414128 800 414248
rect 139200 414128 140000 414248
rect 0 413448 800 413568
rect 139200 413448 140000 413568
rect 0 412768 800 412888
rect 139200 412768 140000 412888
rect 0 412088 800 412208
rect 139200 411408 140000 411528
rect 0 410728 800 410848
rect 139200 410728 140000 410848
rect 0 410048 800 410168
rect 139200 410048 140000 410168
rect 0 409368 800 409488
rect 139200 409368 140000 409488
rect 0 408688 800 408808
rect 139200 408688 140000 408808
rect 0 408008 800 408128
rect 139200 407328 140000 407448
rect 0 406648 800 406768
rect 139200 406648 140000 406768
rect 0 405968 800 406088
rect 139200 405968 140000 406088
rect 0 405288 800 405408
rect 139200 405288 140000 405408
rect 0 404608 800 404728
rect 139200 404608 140000 404728
rect 0 403928 800 404048
rect 139200 403928 140000 404048
rect 0 402568 800 402688
rect 139200 402568 140000 402688
rect 0 401888 800 402008
rect 139200 401888 140000 402008
rect 0 401208 800 401328
rect 139200 401208 140000 401328
rect 0 400528 800 400648
rect 139200 400528 140000 400648
rect 0 399848 800 399968
rect 139200 399848 140000 399968
rect 0 398488 800 398608
rect 139200 398488 140000 398608
rect 0 397808 800 397928
rect 139200 397808 140000 397928
rect 0 397128 800 397248
rect 139200 397128 140000 397248
rect 0 396448 800 396568
rect 139200 396448 140000 396568
rect 0 395768 800 395888
rect 139200 395768 140000 395888
rect 0 395088 800 395208
rect 139200 394408 140000 394528
rect 0 393728 800 393848
rect 139200 393728 140000 393848
rect 0 393048 800 393168
rect 139200 393048 140000 393168
rect 0 392368 800 392488
rect 139200 392368 140000 392488
rect 0 391688 800 391808
rect 139200 391688 140000 391808
rect 0 391008 800 391128
rect 139200 390328 140000 390448
rect 0 389648 800 389768
rect 139200 389648 140000 389768
rect 0 388968 800 389088
rect 139200 388968 140000 389088
rect 0 388288 800 388408
rect 139200 388288 140000 388408
rect 0 387608 800 387728
rect 139200 387608 140000 387728
rect 0 386928 800 387048
rect 139200 386928 140000 387048
rect 0 385568 800 385688
rect 139200 385568 140000 385688
rect 0 384888 800 385008
rect 139200 384888 140000 385008
rect 0 384208 800 384328
rect 139200 384208 140000 384328
rect 0 383528 800 383648
rect 139200 383528 140000 383648
rect 0 382848 800 382968
rect 139200 382848 140000 382968
rect 0 381488 800 381608
rect 139200 381488 140000 381608
rect 0 380808 800 380928
rect 139200 380808 140000 380928
rect 0 380128 800 380248
rect 139200 380128 140000 380248
rect 0 379448 800 379568
rect 139200 379448 140000 379568
rect 0 378768 800 378888
rect 139200 378768 140000 378888
rect 0 378088 800 378208
rect 139200 377408 140000 377528
rect 0 376728 800 376848
rect 139200 376728 140000 376848
rect 0 376048 800 376168
rect 139200 376048 140000 376168
rect 0 375368 800 375488
rect 139200 375368 140000 375488
rect 0 374688 800 374808
rect 139200 374688 140000 374808
rect 0 374008 800 374128
rect 139200 373328 140000 373448
rect 0 372648 800 372768
rect 139200 372648 140000 372768
rect 0 371968 800 372088
rect 139200 371968 140000 372088
rect 0 371288 800 371408
rect 139200 371288 140000 371408
rect 0 370608 800 370728
rect 139200 370608 140000 370728
rect 0 369928 800 370048
rect 139200 369928 140000 370048
rect 0 368568 800 368688
rect 139200 368568 140000 368688
rect 0 367888 800 368008
rect 139200 367888 140000 368008
rect 0 367208 800 367328
rect 139200 367208 140000 367328
rect 0 366528 800 366648
rect 139200 366528 140000 366648
rect 0 365848 800 365968
rect 139200 365848 140000 365968
rect 0 364488 800 364608
rect 139200 364488 140000 364608
rect 0 363808 800 363928
rect 139200 363808 140000 363928
rect 0 363128 800 363248
rect 139200 363128 140000 363248
rect 0 362448 800 362568
rect 139200 362448 140000 362568
rect 0 361768 800 361888
rect 139200 361768 140000 361888
rect 0 361088 800 361208
rect 139200 360408 140000 360528
rect 0 359728 800 359848
rect 139200 359728 140000 359848
rect 0 359048 800 359168
rect 139200 359048 140000 359168
rect 0 358368 800 358488
rect 139200 358368 140000 358488
rect 0 357688 800 357808
rect 139200 357688 140000 357808
rect 0 357008 800 357128
rect 139200 356328 140000 356448
rect 0 355648 800 355768
rect 139200 355648 140000 355768
rect 0 354968 800 355088
rect 139200 354968 140000 355088
rect 0 354288 800 354408
rect 139200 354288 140000 354408
rect 0 353608 800 353728
rect 139200 353608 140000 353728
rect 0 352928 800 353048
rect 139200 352928 140000 353048
rect 0 351568 800 351688
rect 139200 351568 140000 351688
rect 0 350888 800 351008
rect 139200 350888 140000 351008
rect 0 350208 800 350328
rect 139200 350208 140000 350328
rect 0 349528 800 349648
rect 139200 349528 140000 349648
rect 0 348848 800 348968
rect 139200 348848 140000 348968
rect 0 347488 800 347608
rect 139200 347488 140000 347608
rect 0 346808 800 346928
rect 139200 346808 140000 346928
rect 0 346128 800 346248
rect 139200 346128 140000 346248
rect 0 345448 800 345568
rect 139200 345448 140000 345568
rect 0 344768 800 344888
rect 139200 344768 140000 344888
rect 0 344088 800 344208
rect 139200 343408 140000 343528
rect 0 342728 800 342848
rect 139200 342728 140000 342848
rect 0 342048 800 342168
rect 139200 342048 140000 342168
rect 0 341368 800 341488
rect 139200 341368 140000 341488
rect 0 340688 800 340808
rect 139200 340688 140000 340808
rect 0 340008 800 340128
rect 139200 339328 140000 339448
rect 0 338648 800 338768
rect 139200 338648 140000 338768
rect 0 337968 800 338088
rect 139200 337968 140000 338088
rect 0 337288 800 337408
rect 139200 337288 140000 337408
rect 0 336608 800 336728
rect 139200 336608 140000 336728
rect 0 335928 800 336048
rect 139200 335928 140000 336048
rect 0 334568 800 334688
rect 139200 334568 140000 334688
rect 0 333888 800 334008
rect 139200 333888 140000 334008
rect 0 333208 800 333328
rect 139200 333208 140000 333328
rect 0 332528 800 332648
rect 139200 332528 140000 332648
rect 0 331848 800 331968
rect 139200 331848 140000 331968
rect 0 330488 800 330608
rect 139200 330488 140000 330608
rect 0 329808 800 329928
rect 139200 329808 140000 329928
rect 0 329128 800 329248
rect 139200 329128 140000 329248
rect 0 328448 800 328568
rect 139200 328448 140000 328568
rect 0 327768 800 327888
rect 139200 327768 140000 327888
rect 0 327088 800 327208
rect 139200 326408 140000 326528
rect 0 325728 800 325848
rect 139200 325728 140000 325848
rect 0 325048 800 325168
rect 139200 325048 140000 325168
rect 0 324368 800 324488
rect 139200 324368 140000 324488
rect 0 323688 800 323808
rect 139200 323688 140000 323808
rect 0 323008 800 323128
rect 139200 322328 140000 322448
rect 0 321648 800 321768
rect 139200 321648 140000 321768
rect 0 320968 800 321088
rect 139200 320968 140000 321088
rect 0 320288 800 320408
rect 139200 320288 140000 320408
rect 0 319608 800 319728
rect 139200 319608 140000 319728
rect 0 318928 800 319048
rect 139200 318248 140000 318368
rect 0 317568 800 317688
rect 139200 317568 140000 317688
rect 0 316888 800 317008
rect 139200 316888 140000 317008
rect 0 316208 800 316328
rect 139200 316208 140000 316328
rect 0 315528 800 315648
rect 139200 315528 140000 315648
rect 0 314848 800 314968
rect 139200 314848 140000 314968
rect 0 313488 800 313608
rect 139200 313488 140000 313608
rect 0 312808 800 312928
rect 139200 312808 140000 312928
rect 0 312128 800 312248
rect 139200 312128 140000 312248
rect 0 311448 800 311568
rect 139200 311448 140000 311568
rect 0 310768 800 310888
rect 139200 310768 140000 310888
rect 0 310088 800 310208
rect 139200 309408 140000 309528
rect 0 308728 800 308848
rect 139200 308728 140000 308848
rect 0 308048 800 308168
rect 139200 308048 140000 308168
rect 0 307368 800 307488
rect 139200 307368 140000 307488
rect 0 306688 800 306808
rect 139200 306688 140000 306808
rect 0 306008 800 306128
rect 139200 305328 140000 305448
rect 0 304648 800 304768
rect 139200 304648 140000 304768
rect 0 303968 800 304088
rect 139200 303968 140000 304088
rect 0 303288 800 303408
rect 139200 303288 140000 303408
rect 0 302608 800 302728
rect 139200 302608 140000 302728
rect 0 301928 800 302048
rect 139200 301248 140000 301368
rect 0 300568 800 300688
rect 139200 300568 140000 300688
rect 0 299888 800 300008
rect 139200 299888 140000 300008
rect 0 299208 800 299328
rect 139200 299208 140000 299328
rect 0 298528 800 298648
rect 139200 298528 140000 298648
rect 0 297848 800 297968
rect 139200 297848 140000 297968
rect 0 296488 800 296608
rect 139200 296488 140000 296608
rect 0 295808 800 295928
rect 139200 295808 140000 295928
rect 0 295128 800 295248
rect 139200 295128 140000 295248
rect 0 294448 800 294568
rect 139200 294448 140000 294568
rect 0 293768 800 293888
rect 139200 293768 140000 293888
rect 0 293088 800 293208
rect 139200 292408 140000 292528
rect 0 291728 800 291848
rect 139200 291728 140000 291848
rect 0 291048 800 291168
rect 139200 291048 140000 291168
rect 0 290368 800 290488
rect 139200 290368 140000 290488
rect 0 289688 800 289808
rect 139200 289688 140000 289808
rect 0 289008 800 289128
rect 139200 288328 140000 288448
rect 0 287648 800 287768
rect 139200 287648 140000 287768
rect 0 286968 800 287088
rect 139200 286968 140000 287088
rect 0 286288 800 286408
rect 139200 286288 140000 286408
rect 0 285608 800 285728
rect 139200 285608 140000 285728
rect 0 284928 800 285048
rect 139200 284248 140000 284368
rect 0 283568 800 283688
rect 139200 283568 140000 283688
rect 0 282888 800 283008
rect 139200 282888 140000 283008
rect 0 282208 800 282328
rect 139200 282208 140000 282328
rect 0 281528 800 281648
rect 139200 281528 140000 281648
rect 0 280848 800 280968
rect 139200 280848 140000 280968
rect 0 279488 800 279608
rect 139200 279488 140000 279608
rect 0 278808 800 278928
rect 139200 278808 140000 278928
rect 0 278128 800 278248
rect 139200 278128 140000 278248
rect 0 277448 800 277568
rect 139200 277448 140000 277568
rect 0 276768 800 276888
rect 139200 276768 140000 276888
rect 0 276088 800 276208
rect 139200 275408 140000 275528
rect 0 274728 800 274848
rect 139200 274728 140000 274848
rect 0 274048 800 274168
rect 139200 274048 140000 274168
rect 0 273368 800 273488
rect 139200 273368 140000 273488
rect 0 272688 800 272808
rect 139200 272688 140000 272808
rect 0 272008 800 272128
rect 139200 271328 140000 271448
rect 0 270648 800 270768
rect 139200 270648 140000 270768
rect 0 269968 800 270088
rect 139200 269968 140000 270088
rect 0 269288 800 269408
rect 139200 269288 140000 269408
rect 0 268608 800 268728
rect 139200 268608 140000 268728
rect 0 267928 800 268048
rect 139200 267248 140000 267368
rect 0 266568 800 266688
rect 139200 266568 140000 266688
rect 0 265888 800 266008
rect 139200 265888 140000 266008
rect 0 265208 800 265328
rect 139200 265208 140000 265328
rect 0 264528 800 264648
rect 139200 264528 140000 264648
rect 0 263848 800 263968
rect 139200 263848 140000 263968
rect 0 262488 800 262608
rect 139200 262488 140000 262608
rect 0 261808 800 261928
rect 139200 261808 140000 261928
rect 0 261128 800 261248
rect 139200 261128 140000 261248
rect 0 260448 800 260568
rect 139200 260448 140000 260568
rect 0 259768 800 259888
rect 139200 259768 140000 259888
rect 0 259088 800 259208
rect 139200 258408 140000 258528
rect 0 257728 800 257848
rect 139200 257728 140000 257848
rect 0 257048 800 257168
rect 139200 257048 140000 257168
rect 0 256368 800 256488
rect 139200 256368 140000 256488
rect 0 255688 800 255808
rect 139200 255688 140000 255808
rect 0 255008 800 255128
rect 139200 254328 140000 254448
rect 0 253648 800 253768
rect 139200 253648 140000 253768
rect 0 252968 800 253088
rect 139200 252968 140000 253088
rect 0 252288 800 252408
rect 139200 252288 140000 252408
rect 0 251608 800 251728
rect 139200 251608 140000 251728
rect 0 250928 800 251048
rect 139200 250248 140000 250368
rect 0 249568 800 249688
rect 139200 249568 140000 249688
rect 0 248888 800 249008
rect 139200 248888 140000 249008
rect 0 248208 800 248328
rect 139200 248208 140000 248328
rect 0 247528 800 247648
rect 139200 247528 140000 247648
rect 0 246848 800 246968
rect 139200 246848 140000 246968
rect 0 245488 800 245608
rect 139200 245488 140000 245608
rect 0 244808 800 244928
rect 139200 244808 140000 244928
rect 0 244128 800 244248
rect 139200 244128 140000 244248
rect 0 243448 800 243568
rect 139200 243448 140000 243568
rect 0 242768 800 242888
rect 139200 242768 140000 242888
rect 0 242088 800 242208
rect 139200 241408 140000 241528
rect 0 240728 800 240848
rect 139200 240728 140000 240848
rect 0 240048 800 240168
rect 139200 240048 140000 240168
rect 0 239368 800 239488
rect 139200 239368 140000 239488
rect 0 238688 800 238808
rect 139200 238688 140000 238808
rect 0 238008 800 238128
rect 139200 237328 140000 237448
rect 0 236648 800 236768
rect 139200 236648 140000 236768
rect 0 235968 800 236088
rect 139200 235968 140000 236088
rect 0 235288 800 235408
rect 139200 235288 140000 235408
rect 0 234608 800 234728
rect 139200 234608 140000 234728
rect 0 233928 800 234048
rect 139200 233248 140000 233368
rect 0 232568 800 232688
rect 139200 232568 140000 232688
rect 0 231888 800 232008
rect 139200 231888 140000 232008
rect 0 231208 800 231328
rect 139200 231208 140000 231328
rect 0 230528 800 230648
rect 139200 230528 140000 230648
rect 0 229848 800 229968
rect 139200 229848 140000 229968
rect 0 228488 800 228608
rect 139200 228488 140000 228608
rect 0 227808 800 227928
rect 139200 227808 140000 227928
rect 0 227128 800 227248
rect 139200 227128 140000 227248
rect 0 226448 800 226568
rect 139200 226448 140000 226568
rect 0 225768 800 225888
rect 139200 225768 140000 225888
rect 0 224408 800 224528
rect 139200 224408 140000 224528
rect 0 223728 800 223848
rect 139200 223728 140000 223848
rect 0 223048 800 223168
rect 139200 223048 140000 223168
rect 0 222368 800 222488
rect 139200 222368 140000 222488
rect 0 221688 800 221808
rect 139200 221688 140000 221808
rect 0 221008 800 221128
rect 139200 220328 140000 220448
rect 0 219648 800 219768
rect 139200 219648 140000 219768
rect 0 218968 800 219088
rect 139200 218968 140000 219088
rect 0 218288 800 218408
rect 139200 218288 140000 218408
rect 0 217608 800 217728
rect 139200 217608 140000 217728
rect 0 216928 800 217048
rect 139200 216248 140000 216368
rect 0 215568 800 215688
rect 139200 215568 140000 215688
rect 0 214888 800 215008
rect 139200 214888 140000 215008
rect 0 214208 800 214328
rect 139200 214208 140000 214328
rect 0 213528 800 213648
rect 139200 213528 140000 213648
rect 0 212848 800 212968
rect 139200 212848 140000 212968
rect 0 211488 800 211608
rect 139200 211488 140000 211608
rect 0 210808 800 210928
rect 139200 210808 140000 210928
rect 0 210128 800 210248
rect 139200 210128 140000 210248
rect 0 209448 800 209568
rect 139200 209448 140000 209568
rect 0 208768 800 208888
rect 139200 208768 140000 208888
rect 0 207408 800 207528
rect 139200 207408 140000 207528
rect 0 206728 800 206848
rect 139200 206728 140000 206848
rect 0 206048 800 206168
rect 139200 206048 140000 206168
rect 0 205368 800 205488
rect 139200 205368 140000 205488
rect 0 204688 800 204808
rect 139200 204688 140000 204808
rect 0 204008 800 204128
rect 139200 203328 140000 203448
rect 0 202648 800 202768
rect 139200 202648 140000 202768
rect 0 201968 800 202088
rect 139200 201968 140000 202088
rect 0 201288 800 201408
rect 139200 201288 140000 201408
rect 0 200608 800 200728
rect 139200 200608 140000 200728
rect 0 199928 800 200048
rect 139200 199248 140000 199368
rect 0 198568 800 198688
rect 139200 198568 140000 198688
rect 0 197888 800 198008
rect 139200 197888 140000 198008
rect 0 197208 800 197328
rect 139200 197208 140000 197328
rect 0 196528 800 196648
rect 139200 196528 140000 196648
rect 0 195848 800 195968
rect 139200 195848 140000 195968
rect 0 194488 800 194608
rect 139200 194488 140000 194608
rect 0 193808 800 193928
rect 139200 193808 140000 193928
rect 0 193128 800 193248
rect 139200 193128 140000 193248
rect 0 192448 800 192568
rect 139200 192448 140000 192568
rect 0 191768 800 191888
rect 139200 191768 140000 191888
rect 0 190408 800 190528
rect 139200 190408 140000 190528
rect 0 189728 800 189848
rect 139200 189728 140000 189848
rect 0 189048 800 189168
rect 139200 189048 140000 189168
rect 0 188368 800 188488
rect 139200 188368 140000 188488
rect 0 187688 800 187808
rect 139200 187688 140000 187808
rect 0 187008 800 187128
rect 139200 186328 140000 186448
rect 0 185648 800 185768
rect 139200 185648 140000 185768
rect 0 184968 800 185088
rect 139200 184968 140000 185088
rect 0 184288 800 184408
rect 139200 184288 140000 184408
rect 0 183608 800 183728
rect 139200 183608 140000 183728
rect 0 182928 800 183048
rect 139200 182248 140000 182368
rect 0 181568 800 181688
rect 139200 181568 140000 181688
rect 0 180888 800 181008
rect 139200 180888 140000 181008
rect 0 180208 800 180328
rect 139200 180208 140000 180328
rect 0 179528 800 179648
rect 139200 179528 140000 179648
rect 0 178848 800 178968
rect 139200 178848 140000 178968
rect 0 177488 800 177608
rect 139200 177488 140000 177608
rect 0 176808 800 176928
rect 139200 176808 140000 176928
rect 0 176128 800 176248
rect 139200 176128 140000 176248
rect 0 175448 800 175568
rect 139200 175448 140000 175568
rect 0 174768 800 174888
rect 139200 174768 140000 174888
rect 0 173408 800 173528
rect 139200 173408 140000 173528
rect 0 172728 800 172848
rect 139200 172728 140000 172848
rect 0 172048 800 172168
rect 139200 172048 140000 172168
rect 0 171368 800 171488
rect 139200 171368 140000 171488
rect 0 170688 800 170808
rect 139200 170688 140000 170808
rect 0 170008 800 170128
rect 139200 169328 140000 169448
rect 0 168648 800 168768
rect 139200 168648 140000 168768
rect 0 167968 800 168088
rect 139200 167968 140000 168088
rect 0 167288 800 167408
rect 139200 167288 140000 167408
rect 0 166608 800 166728
rect 139200 166608 140000 166728
rect 0 165928 800 166048
rect 139200 165248 140000 165368
rect 0 164568 800 164688
rect 139200 164568 140000 164688
rect 0 163888 800 164008
rect 139200 163888 140000 164008
rect 0 163208 800 163328
rect 139200 163208 140000 163328
rect 0 162528 800 162648
rect 139200 162528 140000 162648
rect 0 161848 800 161968
rect 139200 161848 140000 161968
rect 0 160488 800 160608
rect 139200 160488 140000 160608
rect 0 159808 800 159928
rect 139200 159808 140000 159928
rect 0 159128 800 159248
rect 139200 159128 140000 159248
rect 0 158448 800 158568
rect 139200 158448 140000 158568
rect 0 157768 800 157888
rect 139200 157768 140000 157888
rect 0 156408 800 156528
rect 139200 156408 140000 156528
rect 0 155728 800 155848
rect 139200 155728 140000 155848
rect 0 155048 800 155168
rect 139200 155048 140000 155168
rect 0 154368 800 154488
rect 139200 154368 140000 154488
rect 0 153688 800 153808
rect 139200 153688 140000 153808
rect 0 153008 800 153128
rect 139200 152328 140000 152448
rect 0 151648 800 151768
rect 139200 151648 140000 151768
rect 0 150968 800 151088
rect 139200 150968 140000 151088
rect 0 150288 800 150408
rect 139200 150288 140000 150408
rect 0 149608 800 149728
rect 139200 149608 140000 149728
rect 0 148928 800 149048
rect 139200 148248 140000 148368
rect 0 147568 800 147688
rect 139200 147568 140000 147688
rect 0 146888 800 147008
rect 139200 146888 140000 147008
rect 0 146208 800 146328
rect 139200 146208 140000 146328
rect 0 145528 800 145648
rect 139200 145528 140000 145648
rect 0 144848 800 144968
rect 139200 144848 140000 144968
rect 0 143488 800 143608
rect 139200 143488 140000 143608
rect 0 142808 800 142928
rect 139200 142808 140000 142928
rect 0 142128 800 142248
rect 139200 142128 140000 142248
rect 0 141448 800 141568
rect 139200 141448 140000 141568
rect 0 140768 800 140888
rect 139200 140768 140000 140888
rect 0 139408 800 139528
rect 139200 139408 140000 139528
rect 0 138728 800 138848
rect 139200 138728 140000 138848
rect 0 138048 800 138168
rect 139200 138048 140000 138168
rect 0 137368 800 137488
rect 139200 137368 140000 137488
rect 0 136688 800 136808
rect 139200 136688 140000 136808
rect 0 136008 800 136128
rect 139200 135328 140000 135448
rect 0 134648 800 134768
rect 139200 134648 140000 134768
rect 0 133968 800 134088
rect 139200 133968 140000 134088
rect 0 133288 800 133408
rect 139200 133288 140000 133408
rect 0 132608 800 132728
rect 139200 132608 140000 132728
rect 0 131928 800 132048
rect 139200 131248 140000 131368
rect 0 130568 800 130688
rect 139200 130568 140000 130688
rect 0 129888 800 130008
rect 139200 129888 140000 130008
rect 0 129208 800 129328
rect 139200 129208 140000 129328
rect 0 128528 800 128648
rect 139200 128528 140000 128648
rect 0 127848 800 127968
rect 139200 127848 140000 127968
rect 0 126488 800 126608
rect 139200 126488 140000 126608
rect 0 125808 800 125928
rect 139200 125808 140000 125928
rect 0 125128 800 125248
rect 139200 125128 140000 125248
rect 0 124448 800 124568
rect 139200 124448 140000 124568
rect 0 123768 800 123888
rect 139200 123768 140000 123888
rect 0 122408 800 122528
rect 139200 122408 140000 122528
rect 0 121728 800 121848
rect 139200 121728 140000 121848
rect 0 121048 800 121168
rect 139200 121048 140000 121168
rect 0 120368 800 120488
rect 139200 120368 140000 120488
rect 0 119688 800 119808
rect 139200 119688 140000 119808
rect 0 119008 800 119128
rect 139200 118328 140000 118448
rect 0 117648 800 117768
rect 139200 117648 140000 117768
rect 0 116968 800 117088
rect 139200 116968 140000 117088
rect 0 116288 800 116408
rect 139200 116288 140000 116408
rect 0 115608 800 115728
rect 139200 115608 140000 115728
rect 0 114928 800 115048
rect 139200 114248 140000 114368
rect 0 113568 800 113688
rect 139200 113568 140000 113688
rect 0 112888 800 113008
rect 139200 112888 140000 113008
rect 0 112208 800 112328
rect 139200 112208 140000 112328
rect 0 111528 800 111648
rect 139200 111528 140000 111648
rect 0 110848 800 110968
rect 139200 110848 140000 110968
rect 0 109488 800 109608
rect 139200 109488 140000 109608
rect 0 108808 800 108928
rect 139200 108808 140000 108928
rect 0 108128 800 108248
rect 139200 108128 140000 108248
rect 0 107448 800 107568
rect 139200 107448 140000 107568
rect 0 106768 800 106888
rect 139200 106768 140000 106888
rect 0 105408 800 105528
rect 139200 105408 140000 105528
rect 0 104728 800 104848
rect 139200 104728 140000 104848
rect 0 104048 800 104168
rect 139200 104048 140000 104168
rect 0 103368 800 103488
rect 139200 103368 140000 103488
rect 0 102688 800 102808
rect 139200 102688 140000 102808
rect 0 102008 800 102128
rect 139200 101328 140000 101448
rect 0 100648 800 100768
rect 139200 100648 140000 100768
rect 0 99968 800 100088
rect 139200 99968 140000 100088
rect 0 99288 800 99408
rect 139200 99288 140000 99408
rect 0 98608 800 98728
rect 139200 98608 140000 98728
rect 0 97928 800 98048
rect 139200 97248 140000 97368
rect 0 96568 800 96688
rect 139200 96568 140000 96688
rect 0 95888 800 96008
rect 139200 95888 140000 96008
rect 0 95208 800 95328
rect 139200 95208 140000 95328
rect 0 94528 800 94648
rect 139200 94528 140000 94648
rect 0 93848 800 93968
rect 139200 93848 140000 93968
rect 0 92488 800 92608
rect 139200 92488 140000 92608
rect 0 91808 800 91928
rect 139200 91808 140000 91928
rect 0 91128 800 91248
rect 139200 91128 140000 91248
rect 0 90448 800 90568
rect 139200 90448 140000 90568
rect 0 89768 800 89888
rect 139200 89768 140000 89888
rect 0 88408 800 88528
rect 139200 88408 140000 88528
rect 0 87728 800 87848
rect 139200 87728 140000 87848
rect 0 87048 800 87168
rect 139200 87048 140000 87168
rect 0 86368 800 86488
rect 139200 86368 140000 86488
rect 0 85688 800 85808
rect 139200 85688 140000 85808
rect 0 85008 800 85128
rect 139200 84328 140000 84448
rect 0 83648 800 83768
rect 139200 83648 140000 83768
rect 0 82968 800 83088
rect 139200 82968 140000 83088
rect 0 82288 800 82408
rect 139200 82288 140000 82408
rect 0 81608 800 81728
rect 139200 81608 140000 81728
rect 0 80928 800 81048
rect 139200 80248 140000 80368
rect 0 79568 800 79688
rect 139200 79568 140000 79688
rect 0 78888 800 79008
rect 139200 78888 140000 79008
rect 0 78208 800 78328
rect 139200 78208 140000 78328
rect 0 77528 800 77648
rect 139200 77528 140000 77648
rect 0 76848 800 76968
rect 139200 76168 140000 76288
rect 0 75488 800 75608
rect 139200 75488 140000 75608
rect 0 74808 800 74928
rect 139200 74808 140000 74928
rect 0 74128 800 74248
rect 139200 74128 140000 74248
rect 0 73448 800 73568
rect 139200 73448 140000 73568
rect 0 72768 800 72888
rect 139200 72768 140000 72888
rect 0 71408 800 71528
rect 139200 71408 140000 71528
rect 0 70728 800 70848
rect 139200 70728 140000 70848
rect 0 70048 800 70168
rect 139200 70048 140000 70168
rect 0 69368 800 69488
rect 139200 69368 140000 69488
rect 0 68688 800 68808
rect 139200 68688 140000 68808
rect 0 68008 800 68128
rect 139200 67328 140000 67448
rect 0 66648 800 66768
rect 139200 66648 140000 66768
rect 0 65968 800 66088
rect 139200 65968 140000 66088
rect 0 65288 800 65408
rect 139200 65288 140000 65408
rect 0 64608 800 64728
rect 139200 64608 140000 64728
rect 0 63928 800 64048
rect 139200 63248 140000 63368
rect 0 62568 800 62688
rect 139200 62568 140000 62688
rect 0 61888 800 62008
rect 139200 61888 140000 62008
rect 0 61208 800 61328
rect 139200 61208 140000 61328
rect 0 60528 800 60648
rect 139200 60528 140000 60648
rect 0 59848 800 59968
rect 139200 59168 140000 59288
rect 0 58488 800 58608
rect 139200 58488 140000 58608
rect 0 57808 800 57928
rect 139200 57808 140000 57928
rect 0 57128 800 57248
rect 139200 57128 140000 57248
rect 0 56448 800 56568
rect 139200 56448 140000 56568
rect 0 55768 800 55888
rect 139200 55768 140000 55888
rect 0 54408 800 54528
rect 139200 54408 140000 54528
rect 0 53728 800 53848
rect 139200 53728 140000 53848
rect 0 53048 800 53168
rect 139200 53048 140000 53168
rect 0 52368 800 52488
rect 139200 52368 140000 52488
rect 0 51688 800 51808
rect 139200 51688 140000 51808
rect 0 51008 800 51128
rect 139200 50328 140000 50448
rect 0 49648 800 49768
rect 139200 49648 140000 49768
rect 0 48968 800 49088
rect 139200 48968 140000 49088
rect 0 48288 800 48408
rect 139200 48288 140000 48408
rect 0 47608 800 47728
rect 139200 47608 140000 47728
rect 0 46928 800 47048
rect 139200 46248 140000 46368
rect 0 45568 800 45688
rect 139200 45568 140000 45688
rect 0 44888 800 45008
rect 139200 44888 140000 45008
rect 0 44208 800 44328
rect 139200 44208 140000 44328
rect 0 43528 800 43648
rect 139200 43528 140000 43648
rect 0 42848 800 42968
rect 139200 42168 140000 42288
rect 0 41488 800 41608
rect 139200 41488 140000 41608
rect 0 40808 800 40928
rect 139200 40808 140000 40928
rect 0 40128 800 40248
rect 139200 40128 140000 40248
rect 0 39448 800 39568
rect 139200 39448 140000 39568
rect 0 38768 800 38888
rect 139200 38768 140000 38888
rect 0 37408 800 37528
rect 139200 37408 140000 37528
rect 0 36728 800 36848
rect 139200 36728 140000 36848
rect 0 36048 800 36168
rect 139200 36048 140000 36168
rect 0 35368 800 35488
rect 139200 35368 140000 35488
rect 0 34688 800 34808
rect 139200 34688 140000 34808
rect 0 34008 800 34128
rect 139200 33328 140000 33448
rect 0 32648 800 32768
rect 139200 32648 140000 32768
rect 0 31968 800 32088
rect 139200 31968 140000 32088
rect 0 31288 800 31408
rect 139200 31288 140000 31408
rect 0 30608 800 30728
rect 139200 30608 140000 30728
rect 0 29928 800 30048
rect 139200 29248 140000 29368
rect 0 28568 800 28688
rect 139200 28568 140000 28688
rect 0 27888 800 28008
rect 139200 27888 140000 28008
rect 0 27208 800 27328
rect 139200 27208 140000 27328
rect 0 26528 800 26648
rect 139200 26528 140000 26648
rect 0 25848 800 25968
rect 139200 25168 140000 25288
rect 0 24488 800 24608
rect 139200 24488 140000 24608
rect 0 23808 800 23928
rect 139200 23808 140000 23928
rect 0 23128 800 23248
rect 139200 23128 140000 23248
rect 0 22448 800 22568
rect 139200 22448 140000 22568
rect 0 21768 800 21888
rect 139200 21768 140000 21888
rect 0 20408 800 20528
rect 139200 20408 140000 20528
rect 0 19728 800 19848
rect 139200 19728 140000 19848
rect 0 19048 800 19168
rect 139200 19048 140000 19168
rect 0 18368 800 18488
rect 139200 18368 140000 18488
rect 0 17688 800 17808
rect 139200 17688 140000 17808
rect 0 17008 800 17128
rect 139200 16328 140000 16448
rect 0 15648 800 15768
rect 139200 15648 140000 15768
rect 0 14968 800 15088
rect 139200 14968 140000 15088
rect 0 14288 800 14408
rect 139200 14288 140000 14408
rect 0 13608 800 13728
rect 139200 13608 140000 13728
rect 0 12928 800 13048
rect 139200 12248 140000 12368
rect 0 11568 800 11688
rect 139200 11568 140000 11688
rect 0 10888 800 11008
rect 139200 10888 140000 11008
rect 0 10208 800 10328
rect 139200 10208 140000 10328
rect 0 9528 800 9648
rect 139200 9528 140000 9648
rect 0 8848 800 8968
rect 139200 8168 140000 8288
rect 0 7488 800 7608
rect 139200 7488 140000 7608
rect 0 6808 800 6928
rect 139200 6808 140000 6928
rect 0 6128 800 6248
rect 139200 6128 140000 6248
rect 0 5448 800 5568
rect 139200 5448 140000 5568
rect 0 4768 800 4888
rect 139200 4768 140000 4888
rect 0 3408 800 3528
rect 139200 3408 140000 3528
rect 0 2728 800 2848
rect 139200 2728 140000 2848
rect 0 2048 800 2168
rect 139200 2048 140000 2168
rect 0 1368 800 1488
rect 139200 1368 140000 1488
rect 0 688 800 808
rect 139200 688 140000 808
<< obsm3 >>
rect 880 439208 139120 439381
rect 197 438808 139970 439208
rect 880 438528 139120 438808
rect 197 438128 139970 438528
rect 880 437848 139120 438128
rect 197 436768 139970 437848
rect 880 436488 139120 436768
rect 197 436088 139970 436488
rect 880 435808 139120 436088
rect 197 435408 139970 435808
rect 880 435128 139120 435408
rect 197 434728 139970 435128
rect 880 434448 139120 434728
rect 197 434048 139970 434448
rect 880 433768 139120 434048
rect 197 432688 139970 433768
rect 880 432408 139120 432688
rect 197 432008 139970 432408
rect 880 431728 139120 432008
rect 197 431328 139970 431728
rect 880 431048 139120 431328
rect 197 430648 139970 431048
rect 880 430368 139120 430648
rect 197 429968 139970 430368
rect 880 429688 139120 429968
rect 197 429288 139970 429688
rect 880 429008 139970 429288
rect 197 428608 139970 429008
rect 197 428328 139120 428608
rect 197 427928 139970 428328
rect 880 427648 139120 427928
rect 197 427248 139970 427648
rect 880 426968 139120 427248
rect 197 426568 139970 426968
rect 880 426288 139120 426568
rect 197 425888 139970 426288
rect 880 425608 139120 425888
rect 197 425208 139970 425608
rect 880 424928 139970 425208
rect 197 424528 139970 424928
rect 197 424248 139120 424528
rect 197 423848 139970 424248
rect 880 423568 139120 423848
rect 197 423168 139970 423568
rect 880 422888 139120 423168
rect 197 422488 139970 422888
rect 880 422208 139120 422488
rect 197 421808 139970 422208
rect 880 421528 139120 421808
rect 197 421128 139970 421528
rect 880 420848 139120 421128
rect 197 419768 139970 420848
rect 880 419488 139120 419768
rect 197 419088 139970 419488
rect 880 418808 139120 419088
rect 197 418408 139970 418808
rect 880 418128 139120 418408
rect 197 417728 139970 418128
rect 880 417448 139120 417728
rect 197 417048 139970 417448
rect 880 416768 139120 417048
rect 197 415688 139970 416768
rect 880 415408 139120 415688
rect 197 415008 139970 415408
rect 880 414728 139120 415008
rect 197 414328 139970 414728
rect 880 414048 139120 414328
rect 197 413648 139970 414048
rect 880 413368 139120 413648
rect 197 412968 139970 413368
rect 880 412688 139120 412968
rect 197 412288 139970 412688
rect 880 412008 139970 412288
rect 197 411608 139970 412008
rect 197 411328 139120 411608
rect 197 410928 139970 411328
rect 880 410648 139120 410928
rect 197 410248 139970 410648
rect 880 409968 139120 410248
rect 197 409568 139970 409968
rect 880 409288 139120 409568
rect 197 408888 139970 409288
rect 880 408608 139120 408888
rect 197 408208 139970 408608
rect 880 407928 139970 408208
rect 197 407528 139970 407928
rect 197 407248 139120 407528
rect 197 406848 139970 407248
rect 880 406568 139120 406848
rect 197 406168 139970 406568
rect 880 405888 139120 406168
rect 197 405488 139970 405888
rect 880 405208 139120 405488
rect 197 404808 139970 405208
rect 880 404528 139120 404808
rect 197 404128 139970 404528
rect 880 403848 139120 404128
rect 197 402768 139970 403848
rect 880 402488 139120 402768
rect 197 402088 139970 402488
rect 880 401808 139120 402088
rect 197 401408 139970 401808
rect 880 401128 139120 401408
rect 197 400728 139970 401128
rect 880 400448 139120 400728
rect 197 400048 139970 400448
rect 880 399768 139120 400048
rect 197 398688 139970 399768
rect 880 398408 139120 398688
rect 197 398008 139970 398408
rect 880 397728 139120 398008
rect 197 397328 139970 397728
rect 880 397048 139120 397328
rect 197 396648 139970 397048
rect 880 396368 139120 396648
rect 197 395968 139970 396368
rect 880 395688 139120 395968
rect 197 395288 139970 395688
rect 880 395008 139970 395288
rect 197 394608 139970 395008
rect 197 394328 139120 394608
rect 197 393928 139970 394328
rect 880 393648 139120 393928
rect 197 393248 139970 393648
rect 880 392968 139120 393248
rect 197 392568 139970 392968
rect 880 392288 139120 392568
rect 197 391888 139970 392288
rect 880 391608 139120 391888
rect 197 391208 139970 391608
rect 880 390928 139970 391208
rect 197 390528 139970 390928
rect 197 390248 139120 390528
rect 197 389848 139970 390248
rect 880 389568 139120 389848
rect 197 389168 139970 389568
rect 880 388888 139120 389168
rect 197 388488 139970 388888
rect 880 388208 139120 388488
rect 197 387808 139970 388208
rect 880 387528 139120 387808
rect 197 387128 139970 387528
rect 880 386848 139120 387128
rect 197 385768 139970 386848
rect 880 385488 139120 385768
rect 197 385088 139970 385488
rect 880 384808 139120 385088
rect 197 384408 139970 384808
rect 880 384128 139120 384408
rect 197 383728 139970 384128
rect 880 383448 139120 383728
rect 197 383048 139970 383448
rect 880 382768 139120 383048
rect 197 381688 139970 382768
rect 880 381408 139120 381688
rect 197 381008 139970 381408
rect 880 380728 139120 381008
rect 197 380328 139970 380728
rect 880 380048 139120 380328
rect 197 379648 139970 380048
rect 880 379368 139120 379648
rect 197 378968 139970 379368
rect 880 378688 139120 378968
rect 197 378288 139970 378688
rect 880 378008 139970 378288
rect 197 377608 139970 378008
rect 197 377328 139120 377608
rect 197 376928 139970 377328
rect 880 376648 139120 376928
rect 197 376248 139970 376648
rect 880 375968 139120 376248
rect 197 375568 139970 375968
rect 880 375288 139120 375568
rect 197 374888 139970 375288
rect 880 374608 139120 374888
rect 197 374208 139970 374608
rect 880 373928 139970 374208
rect 197 373528 139970 373928
rect 197 373248 139120 373528
rect 197 372848 139970 373248
rect 880 372568 139120 372848
rect 197 372168 139970 372568
rect 880 371888 139120 372168
rect 197 371488 139970 371888
rect 880 371208 139120 371488
rect 197 370808 139970 371208
rect 880 370528 139120 370808
rect 197 370128 139970 370528
rect 880 369848 139120 370128
rect 197 368768 139970 369848
rect 880 368488 139120 368768
rect 197 368088 139970 368488
rect 880 367808 139120 368088
rect 197 367408 139970 367808
rect 880 367128 139120 367408
rect 197 366728 139970 367128
rect 880 366448 139120 366728
rect 197 366048 139970 366448
rect 880 365768 139120 366048
rect 197 364688 139970 365768
rect 880 364408 139120 364688
rect 197 364008 139970 364408
rect 880 363728 139120 364008
rect 197 363328 139970 363728
rect 880 363048 139120 363328
rect 197 362648 139970 363048
rect 880 362368 139120 362648
rect 197 361968 139970 362368
rect 880 361688 139120 361968
rect 197 361288 139970 361688
rect 880 361008 139970 361288
rect 197 360608 139970 361008
rect 197 360328 139120 360608
rect 197 359928 139970 360328
rect 880 359648 139120 359928
rect 197 359248 139970 359648
rect 880 358968 139120 359248
rect 197 358568 139970 358968
rect 880 358288 139120 358568
rect 197 357888 139970 358288
rect 880 357608 139120 357888
rect 197 357208 139970 357608
rect 880 356928 139970 357208
rect 197 356528 139970 356928
rect 197 356248 139120 356528
rect 197 355848 139970 356248
rect 880 355568 139120 355848
rect 197 355168 139970 355568
rect 880 354888 139120 355168
rect 197 354488 139970 354888
rect 880 354208 139120 354488
rect 197 353808 139970 354208
rect 880 353528 139120 353808
rect 197 353128 139970 353528
rect 880 352848 139120 353128
rect 197 351768 139970 352848
rect 880 351488 139120 351768
rect 197 351088 139970 351488
rect 880 350808 139120 351088
rect 197 350408 139970 350808
rect 880 350128 139120 350408
rect 197 349728 139970 350128
rect 880 349448 139120 349728
rect 197 349048 139970 349448
rect 880 348768 139120 349048
rect 197 347688 139970 348768
rect 880 347408 139120 347688
rect 197 347008 139970 347408
rect 880 346728 139120 347008
rect 197 346328 139970 346728
rect 880 346048 139120 346328
rect 197 345648 139970 346048
rect 880 345368 139120 345648
rect 197 344968 139970 345368
rect 880 344688 139120 344968
rect 197 344288 139970 344688
rect 880 344008 139970 344288
rect 197 343608 139970 344008
rect 197 343328 139120 343608
rect 197 342928 139970 343328
rect 880 342648 139120 342928
rect 197 342248 139970 342648
rect 880 341968 139120 342248
rect 197 341568 139970 341968
rect 880 341288 139120 341568
rect 197 340888 139970 341288
rect 880 340608 139120 340888
rect 197 340208 139970 340608
rect 880 339928 139970 340208
rect 197 339528 139970 339928
rect 197 339248 139120 339528
rect 197 338848 139970 339248
rect 880 338568 139120 338848
rect 197 338168 139970 338568
rect 880 337888 139120 338168
rect 197 337488 139970 337888
rect 880 337208 139120 337488
rect 197 336808 139970 337208
rect 880 336528 139120 336808
rect 197 336128 139970 336528
rect 880 335848 139120 336128
rect 197 334768 139970 335848
rect 880 334488 139120 334768
rect 197 334088 139970 334488
rect 880 333808 139120 334088
rect 197 333408 139970 333808
rect 880 333128 139120 333408
rect 197 332728 139970 333128
rect 880 332448 139120 332728
rect 197 332048 139970 332448
rect 880 331768 139120 332048
rect 197 330688 139970 331768
rect 880 330408 139120 330688
rect 197 330008 139970 330408
rect 880 329728 139120 330008
rect 197 329328 139970 329728
rect 880 329048 139120 329328
rect 197 328648 139970 329048
rect 880 328368 139120 328648
rect 197 327968 139970 328368
rect 880 327688 139120 327968
rect 197 327288 139970 327688
rect 880 327008 139970 327288
rect 197 326608 139970 327008
rect 197 326328 139120 326608
rect 197 325928 139970 326328
rect 880 325648 139120 325928
rect 197 325248 139970 325648
rect 880 324968 139120 325248
rect 197 324568 139970 324968
rect 880 324288 139120 324568
rect 197 323888 139970 324288
rect 880 323608 139120 323888
rect 197 323208 139970 323608
rect 880 322928 139970 323208
rect 197 322528 139970 322928
rect 197 322248 139120 322528
rect 197 321848 139970 322248
rect 880 321568 139120 321848
rect 197 321168 139970 321568
rect 880 320888 139120 321168
rect 197 320488 139970 320888
rect 880 320208 139120 320488
rect 197 319808 139970 320208
rect 880 319528 139120 319808
rect 197 319128 139970 319528
rect 880 318848 139970 319128
rect 197 318448 139970 318848
rect 197 318168 139120 318448
rect 197 317768 139970 318168
rect 880 317488 139120 317768
rect 197 317088 139970 317488
rect 880 316808 139120 317088
rect 197 316408 139970 316808
rect 880 316128 139120 316408
rect 197 315728 139970 316128
rect 880 315448 139120 315728
rect 197 315048 139970 315448
rect 880 314768 139120 315048
rect 197 313688 139970 314768
rect 880 313408 139120 313688
rect 197 313008 139970 313408
rect 880 312728 139120 313008
rect 197 312328 139970 312728
rect 880 312048 139120 312328
rect 197 311648 139970 312048
rect 880 311368 139120 311648
rect 197 310968 139970 311368
rect 880 310688 139120 310968
rect 197 310288 139970 310688
rect 880 310008 139970 310288
rect 197 309608 139970 310008
rect 197 309328 139120 309608
rect 197 308928 139970 309328
rect 880 308648 139120 308928
rect 197 308248 139970 308648
rect 880 307968 139120 308248
rect 197 307568 139970 307968
rect 880 307288 139120 307568
rect 197 306888 139970 307288
rect 880 306608 139120 306888
rect 197 306208 139970 306608
rect 880 305928 139970 306208
rect 197 305528 139970 305928
rect 197 305248 139120 305528
rect 197 304848 139970 305248
rect 880 304568 139120 304848
rect 197 304168 139970 304568
rect 880 303888 139120 304168
rect 197 303488 139970 303888
rect 880 303208 139120 303488
rect 197 302808 139970 303208
rect 880 302528 139120 302808
rect 197 302128 139970 302528
rect 880 301848 139970 302128
rect 197 301448 139970 301848
rect 197 301168 139120 301448
rect 197 300768 139970 301168
rect 880 300488 139120 300768
rect 197 300088 139970 300488
rect 880 299808 139120 300088
rect 197 299408 139970 299808
rect 880 299128 139120 299408
rect 197 298728 139970 299128
rect 880 298448 139120 298728
rect 197 298048 139970 298448
rect 880 297768 139120 298048
rect 197 296688 139970 297768
rect 880 296408 139120 296688
rect 197 296008 139970 296408
rect 880 295728 139120 296008
rect 197 295328 139970 295728
rect 880 295048 139120 295328
rect 197 294648 139970 295048
rect 880 294368 139120 294648
rect 197 293968 139970 294368
rect 880 293688 139120 293968
rect 197 293288 139970 293688
rect 880 293008 139970 293288
rect 197 292608 139970 293008
rect 197 292328 139120 292608
rect 197 291928 139970 292328
rect 880 291648 139120 291928
rect 197 291248 139970 291648
rect 880 290968 139120 291248
rect 197 290568 139970 290968
rect 880 290288 139120 290568
rect 197 289888 139970 290288
rect 880 289608 139120 289888
rect 197 289208 139970 289608
rect 880 288928 139970 289208
rect 197 288528 139970 288928
rect 197 288248 139120 288528
rect 197 287848 139970 288248
rect 880 287568 139120 287848
rect 197 287168 139970 287568
rect 880 286888 139120 287168
rect 197 286488 139970 286888
rect 880 286208 139120 286488
rect 197 285808 139970 286208
rect 880 285528 139120 285808
rect 197 285128 139970 285528
rect 880 284848 139970 285128
rect 197 284448 139970 284848
rect 197 284168 139120 284448
rect 197 283768 139970 284168
rect 880 283488 139120 283768
rect 197 283088 139970 283488
rect 880 282808 139120 283088
rect 197 282408 139970 282808
rect 880 282128 139120 282408
rect 197 281728 139970 282128
rect 880 281448 139120 281728
rect 197 281048 139970 281448
rect 880 280768 139120 281048
rect 197 279688 139970 280768
rect 880 279408 139120 279688
rect 197 279008 139970 279408
rect 880 278728 139120 279008
rect 197 278328 139970 278728
rect 880 278048 139120 278328
rect 197 277648 139970 278048
rect 880 277368 139120 277648
rect 197 276968 139970 277368
rect 880 276688 139120 276968
rect 197 276288 139970 276688
rect 880 276008 139970 276288
rect 197 275608 139970 276008
rect 197 275328 139120 275608
rect 197 274928 139970 275328
rect 880 274648 139120 274928
rect 197 274248 139970 274648
rect 880 273968 139120 274248
rect 197 273568 139970 273968
rect 880 273288 139120 273568
rect 197 272888 139970 273288
rect 880 272608 139120 272888
rect 197 272208 139970 272608
rect 880 271928 139970 272208
rect 197 271528 139970 271928
rect 197 271248 139120 271528
rect 197 270848 139970 271248
rect 880 270568 139120 270848
rect 197 270168 139970 270568
rect 880 269888 139120 270168
rect 197 269488 139970 269888
rect 880 269208 139120 269488
rect 197 268808 139970 269208
rect 880 268528 139120 268808
rect 197 268128 139970 268528
rect 880 267848 139970 268128
rect 197 267448 139970 267848
rect 197 267168 139120 267448
rect 197 266768 139970 267168
rect 880 266488 139120 266768
rect 197 266088 139970 266488
rect 880 265808 139120 266088
rect 197 265408 139970 265808
rect 880 265128 139120 265408
rect 197 264728 139970 265128
rect 880 264448 139120 264728
rect 197 264048 139970 264448
rect 880 263768 139120 264048
rect 197 262688 139970 263768
rect 880 262408 139120 262688
rect 197 262008 139970 262408
rect 880 261728 139120 262008
rect 197 261328 139970 261728
rect 880 261048 139120 261328
rect 197 260648 139970 261048
rect 880 260368 139120 260648
rect 197 259968 139970 260368
rect 880 259688 139120 259968
rect 197 259288 139970 259688
rect 880 259008 139970 259288
rect 197 258608 139970 259008
rect 197 258328 139120 258608
rect 197 257928 139970 258328
rect 880 257648 139120 257928
rect 197 257248 139970 257648
rect 880 256968 139120 257248
rect 197 256568 139970 256968
rect 880 256288 139120 256568
rect 197 255888 139970 256288
rect 880 255608 139120 255888
rect 197 255208 139970 255608
rect 880 254928 139970 255208
rect 197 254528 139970 254928
rect 197 254248 139120 254528
rect 197 253848 139970 254248
rect 880 253568 139120 253848
rect 197 253168 139970 253568
rect 880 252888 139120 253168
rect 197 252488 139970 252888
rect 880 252208 139120 252488
rect 197 251808 139970 252208
rect 880 251528 139120 251808
rect 197 251128 139970 251528
rect 880 250848 139970 251128
rect 197 250448 139970 250848
rect 197 250168 139120 250448
rect 197 249768 139970 250168
rect 880 249488 139120 249768
rect 197 249088 139970 249488
rect 880 248808 139120 249088
rect 197 248408 139970 248808
rect 880 248128 139120 248408
rect 197 247728 139970 248128
rect 880 247448 139120 247728
rect 197 247048 139970 247448
rect 880 246768 139120 247048
rect 197 245688 139970 246768
rect 880 245408 139120 245688
rect 197 245008 139970 245408
rect 880 244728 139120 245008
rect 197 244328 139970 244728
rect 880 244048 139120 244328
rect 197 243648 139970 244048
rect 880 243368 139120 243648
rect 197 242968 139970 243368
rect 880 242688 139120 242968
rect 197 242288 139970 242688
rect 880 242008 139970 242288
rect 197 241608 139970 242008
rect 197 241328 139120 241608
rect 197 240928 139970 241328
rect 880 240648 139120 240928
rect 197 240248 139970 240648
rect 880 239968 139120 240248
rect 197 239568 139970 239968
rect 880 239288 139120 239568
rect 197 238888 139970 239288
rect 880 238608 139120 238888
rect 197 238208 139970 238608
rect 880 237928 139970 238208
rect 197 237528 139970 237928
rect 197 237248 139120 237528
rect 197 236848 139970 237248
rect 880 236568 139120 236848
rect 197 236168 139970 236568
rect 880 235888 139120 236168
rect 197 235488 139970 235888
rect 880 235208 139120 235488
rect 197 234808 139970 235208
rect 880 234528 139120 234808
rect 197 234128 139970 234528
rect 880 233848 139970 234128
rect 197 233448 139970 233848
rect 197 233168 139120 233448
rect 197 232768 139970 233168
rect 880 232488 139120 232768
rect 197 232088 139970 232488
rect 880 231808 139120 232088
rect 197 231408 139970 231808
rect 880 231128 139120 231408
rect 197 230728 139970 231128
rect 880 230448 139120 230728
rect 197 230048 139970 230448
rect 880 229768 139120 230048
rect 197 228688 139970 229768
rect 880 228408 139120 228688
rect 197 228008 139970 228408
rect 880 227728 139120 228008
rect 197 227328 139970 227728
rect 880 227048 139120 227328
rect 197 226648 139970 227048
rect 880 226368 139120 226648
rect 197 225968 139970 226368
rect 880 225688 139120 225968
rect 197 224608 139970 225688
rect 880 224328 139120 224608
rect 197 223928 139970 224328
rect 880 223648 139120 223928
rect 197 223248 139970 223648
rect 880 222968 139120 223248
rect 197 222568 139970 222968
rect 880 222288 139120 222568
rect 197 221888 139970 222288
rect 880 221608 139120 221888
rect 197 221208 139970 221608
rect 880 220928 139970 221208
rect 197 220528 139970 220928
rect 197 220248 139120 220528
rect 197 219848 139970 220248
rect 880 219568 139120 219848
rect 197 219168 139970 219568
rect 880 218888 139120 219168
rect 197 218488 139970 218888
rect 880 218208 139120 218488
rect 197 217808 139970 218208
rect 880 217528 139120 217808
rect 197 217128 139970 217528
rect 880 216848 139970 217128
rect 197 216448 139970 216848
rect 197 216168 139120 216448
rect 197 215768 139970 216168
rect 880 215488 139120 215768
rect 197 215088 139970 215488
rect 880 214808 139120 215088
rect 197 214408 139970 214808
rect 880 214128 139120 214408
rect 197 213728 139970 214128
rect 880 213448 139120 213728
rect 197 213048 139970 213448
rect 880 212768 139120 213048
rect 197 211688 139970 212768
rect 880 211408 139120 211688
rect 197 211008 139970 211408
rect 880 210728 139120 211008
rect 197 210328 139970 210728
rect 880 210048 139120 210328
rect 197 209648 139970 210048
rect 880 209368 139120 209648
rect 197 208968 139970 209368
rect 880 208688 139120 208968
rect 197 207608 139970 208688
rect 880 207328 139120 207608
rect 197 206928 139970 207328
rect 880 206648 139120 206928
rect 197 206248 139970 206648
rect 880 205968 139120 206248
rect 197 205568 139970 205968
rect 880 205288 139120 205568
rect 197 204888 139970 205288
rect 880 204608 139120 204888
rect 197 204208 139970 204608
rect 880 203928 139970 204208
rect 197 203528 139970 203928
rect 197 203248 139120 203528
rect 197 202848 139970 203248
rect 880 202568 139120 202848
rect 197 202168 139970 202568
rect 880 201888 139120 202168
rect 197 201488 139970 201888
rect 880 201208 139120 201488
rect 197 200808 139970 201208
rect 880 200528 139120 200808
rect 197 200128 139970 200528
rect 880 199848 139970 200128
rect 197 199448 139970 199848
rect 197 199168 139120 199448
rect 197 198768 139970 199168
rect 880 198488 139120 198768
rect 197 198088 139970 198488
rect 880 197808 139120 198088
rect 197 197408 139970 197808
rect 880 197128 139120 197408
rect 197 196728 139970 197128
rect 880 196448 139120 196728
rect 197 196048 139970 196448
rect 880 195768 139120 196048
rect 197 194688 139970 195768
rect 880 194408 139120 194688
rect 197 194008 139970 194408
rect 880 193728 139120 194008
rect 197 193328 139970 193728
rect 880 193048 139120 193328
rect 197 192648 139970 193048
rect 880 192368 139120 192648
rect 197 191968 139970 192368
rect 880 191688 139120 191968
rect 197 190608 139970 191688
rect 880 190328 139120 190608
rect 197 189928 139970 190328
rect 880 189648 139120 189928
rect 197 189248 139970 189648
rect 880 188968 139120 189248
rect 197 188568 139970 188968
rect 880 188288 139120 188568
rect 197 187888 139970 188288
rect 880 187608 139120 187888
rect 197 187208 139970 187608
rect 880 186928 139970 187208
rect 197 186528 139970 186928
rect 197 186248 139120 186528
rect 197 185848 139970 186248
rect 880 185568 139120 185848
rect 197 185168 139970 185568
rect 880 184888 139120 185168
rect 197 184488 139970 184888
rect 880 184208 139120 184488
rect 197 183808 139970 184208
rect 880 183528 139120 183808
rect 197 183128 139970 183528
rect 880 182848 139970 183128
rect 197 182448 139970 182848
rect 197 182168 139120 182448
rect 197 181768 139970 182168
rect 880 181488 139120 181768
rect 197 181088 139970 181488
rect 880 180808 139120 181088
rect 197 180408 139970 180808
rect 880 180128 139120 180408
rect 197 179728 139970 180128
rect 880 179448 139120 179728
rect 197 179048 139970 179448
rect 880 178768 139120 179048
rect 197 177688 139970 178768
rect 880 177408 139120 177688
rect 197 177008 139970 177408
rect 880 176728 139120 177008
rect 197 176328 139970 176728
rect 880 176048 139120 176328
rect 197 175648 139970 176048
rect 880 175368 139120 175648
rect 197 174968 139970 175368
rect 880 174688 139120 174968
rect 197 173608 139970 174688
rect 880 173328 139120 173608
rect 197 172928 139970 173328
rect 880 172648 139120 172928
rect 197 172248 139970 172648
rect 880 171968 139120 172248
rect 197 171568 139970 171968
rect 880 171288 139120 171568
rect 197 170888 139970 171288
rect 880 170608 139120 170888
rect 197 170208 139970 170608
rect 880 169928 139970 170208
rect 197 169528 139970 169928
rect 197 169248 139120 169528
rect 197 168848 139970 169248
rect 880 168568 139120 168848
rect 197 168168 139970 168568
rect 880 167888 139120 168168
rect 197 167488 139970 167888
rect 880 167208 139120 167488
rect 197 166808 139970 167208
rect 880 166528 139120 166808
rect 197 166128 139970 166528
rect 880 165848 139970 166128
rect 197 165448 139970 165848
rect 197 165168 139120 165448
rect 197 164768 139970 165168
rect 880 164488 139120 164768
rect 197 164088 139970 164488
rect 880 163808 139120 164088
rect 197 163408 139970 163808
rect 880 163128 139120 163408
rect 197 162728 139970 163128
rect 880 162448 139120 162728
rect 197 162048 139970 162448
rect 880 161768 139120 162048
rect 197 160688 139970 161768
rect 880 160408 139120 160688
rect 197 160008 139970 160408
rect 880 159728 139120 160008
rect 197 159328 139970 159728
rect 880 159048 139120 159328
rect 197 158648 139970 159048
rect 880 158368 139120 158648
rect 197 157968 139970 158368
rect 880 157688 139120 157968
rect 197 156608 139970 157688
rect 880 156328 139120 156608
rect 197 155928 139970 156328
rect 880 155648 139120 155928
rect 197 155248 139970 155648
rect 880 154968 139120 155248
rect 197 154568 139970 154968
rect 880 154288 139120 154568
rect 197 153888 139970 154288
rect 880 153608 139120 153888
rect 197 153208 139970 153608
rect 880 152928 139970 153208
rect 197 152528 139970 152928
rect 197 152248 139120 152528
rect 197 151848 139970 152248
rect 880 151568 139120 151848
rect 197 151168 139970 151568
rect 880 150888 139120 151168
rect 197 150488 139970 150888
rect 880 150208 139120 150488
rect 197 149808 139970 150208
rect 880 149528 139120 149808
rect 197 149128 139970 149528
rect 880 148848 139970 149128
rect 197 148448 139970 148848
rect 197 148168 139120 148448
rect 197 147768 139970 148168
rect 880 147488 139120 147768
rect 197 147088 139970 147488
rect 880 146808 139120 147088
rect 197 146408 139970 146808
rect 880 146128 139120 146408
rect 197 145728 139970 146128
rect 880 145448 139120 145728
rect 197 145048 139970 145448
rect 880 144768 139120 145048
rect 197 143688 139970 144768
rect 880 143408 139120 143688
rect 197 143008 139970 143408
rect 880 142728 139120 143008
rect 197 142328 139970 142728
rect 880 142048 139120 142328
rect 197 141648 139970 142048
rect 880 141368 139120 141648
rect 197 140968 139970 141368
rect 880 140688 139120 140968
rect 197 139608 139970 140688
rect 880 139328 139120 139608
rect 197 138928 139970 139328
rect 880 138648 139120 138928
rect 197 138248 139970 138648
rect 880 137968 139120 138248
rect 197 137568 139970 137968
rect 880 137288 139120 137568
rect 197 136888 139970 137288
rect 880 136608 139120 136888
rect 197 136208 139970 136608
rect 880 135928 139970 136208
rect 197 135528 139970 135928
rect 197 135248 139120 135528
rect 197 134848 139970 135248
rect 880 134568 139120 134848
rect 197 134168 139970 134568
rect 880 133888 139120 134168
rect 197 133488 139970 133888
rect 880 133208 139120 133488
rect 197 132808 139970 133208
rect 880 132528 139120 132808
rect 197 132128 139970 132528
rect 880 131848 139970 132128
rect 197 131448 139970 131848
rect 197 131168 139120 131448
rect 197 130768 139970 131168
rect 880 130488 139120 130768
rect 197 130088 139970 130488
rect 880 129808 139120 130088
rect 197 129408 139970 129808
rect 880 129128 139120 129408
rect 197 128728 139970 129128
rect 880 128448 139120 128728
rect 197 128048 139970 128448
rect 880 127768 139120 128048
rect 197 126688 139970 127768
rect 880 126408 139120 126688
rect 197 126008 139970 126408
rect 880 125728 139120 126008
rect 197 125328 139970 125728
rect 880 125048 139120 125328
rect 197 124648 139970 125048
rect 880 124368 139120 124648
rect 197 123968 139970 124368
rect 880 123688 139120 123968
rect 197 122608 139970 123688
rect 880 122328 139120 122608
rect 197 121928 139970 122328
rect 880 121648 139120 121928
rect 197 121248 139970 121648
rect 880 120968 139120 121248
rect 197 120568 139970 120968
rect 880 120288 139120 120568
rect 197 119888 139970 120288
rect 880 119608 139120 119888
rect 197 119208 139970 119608
rect 880 118928 139970 119208
rect 197 118528 139970 118928
rect 197 118248 139120 118528
rect 197 117848 139970 118248
rect 880 117568 139120 117848
rect 197 117168 139970 117568
rect 880 116888 139120 117168
rect 197 116488 139970 116888
rect 880 116208 139120 116488
rect 197 115808 139970 116208
rect 880 115528 139120 115808
rect 197 115128 139970 115528
rect 880 114848 139970 115128
rect 197 114448 139970 114848
rect 197 114168 139120 114448
rect 197 113768 139970 114168
rect 880 113488 139120 113768
rect 197 113088 139970 113488
rect 880 112808 139120 113088
rect 197 112408 139970 112808
rect 880 112128 139120 112408
rect 197 111728 139970 112128
rect 880 111448 139120 111728
rect 197 111048 139970 111448
rect 880 110768 139120 111048
rect 197 109688 139970 110768
rect 880 109408 139120 109688
rect 197 109008 139970 109408
rect 880 108728 139120 109008
rect 197 108328 139970 108728
rect 880 108048 139120 108328
rect 197 107648 139970 108048
rect 880 107368 139120 107648
rect 197 106968 139970 107368
rect 880 106688 139120 106968
rect 197 105608 139970 106688
rect 880 105328 139120 105608
rect 197 104928 139970 105328
rect 880 104648 139120 104928
rect 197 104248 139970 104648
rect 880 103968 139120 104248
rect 197 103568 139970 103968
rect 880 103288 139120 103568
rect 197 102888 139970 103288
rect 880 102608 139120 102888
rect 197 102208 139970 102608
rect 880 101928 139970 102208
rect 197 101528 139970 101928
rect 197 101248 139120 101528
rect 197 100848 139970 101248
rect 880 100568 139120 100848
rect 197 100168 139970 100568
rect 880 99888 139120 100168
rect 197 99488 139970 99888
rect 880 99208 139120 99488
rect 197 98808 139970 99208
rect 880 98528 139120 98808
rect 197 98128 139970 98528
rect 880 97848 139970 98128
rect 197 97448 139970 97848
rect 197 97168 139120 97448
rect 197 96768 139970 97168
rect 880 96488 139120 96768
rect 197 96088 139970 96488
rect 880 95808 139120 96088
rect 197 95408 139970 95808
rect 880 95128 139120 95408
rect 197 94728 139970 95128
rect 880 94448 139120 94728
rect 197 94048 139970 94448
rect 880 93768 139120 94048
rect 197 92688 139970 93768
rect 880 92408 139120 92688
rect 197 92008 139970 92408
rect 880 91728 139120 92008
rect 197 91328 139970 91728
rect 880 91048 139120 91328
rect 197 90648 139970 91048
rect 880 90368 139120 90648
rect 197 89968 139970 90368
rect 880 89688 139120 89968
rect 197 88608 139970 89688
rect 880 88328 139120 88608
rect 197 87928 139970 88328
rect 880 87648 139120 87928
rect 197 87248 139970 87648
rect 880 86968 139120 87248
rect 197 86568 139970 86968
rect 880 86288 139120 86568
rect 197 85888 139970 86288
rect 880 85608 139120 85888
rect 197 85208 139970 85608
rect 880 84928 139970 85208
rect 197 84528 139970 84928
rect 197 84248 139120 84528
rect 197 83848 139970 84248
rect 880 83568 139120 83848
rect 197 83168 139970 83568
rect 880 82888 139120 83168
rect 197 82488 139970 82888
rect 880 82208 139120 82488
rect 197 81808 139970 82208
rect 880 81528 139120 81808
rect 197 81128 139970 81528
rect 880 80848 139970 81128
rect 197 80448 139970 80848
rect 197 80168 139120 80448
rect 197 79768 139970 80168
rect 880 79488 139120 79768
rect 197 79088 139970 79488
rect 880 78808 139120 79088
rect 197 78408 139970 78808
rect 880 78128 139120 78408
rect 197 77728 139970 78128
rect 880 77448 139120 77728
rect 197 77048 139970 77448
rect 880 76768 139970 77048
rect 197 76368 139970 76768
rect 197 76088 139120 76368
rect 197 75688 139970 76088
rect 880 75408 139120 75688
rect 197 75008 139970 75408
rect 880 74728 139120 75008
rect 197 74328 139970 74728
rect 880 74048 139120 74328
rect 197 73648 139970 74048
rect 880 73368 139120 73648
rect 197 72968 139970 73368
rect 880 72688 139120 72968
rect 197 71608 139970 72688
rect 880 71328 139120 71608
rect 197 70928 139970 71328
rect 880 70648 139120 70928
rect 197 70248 139970 70648
rect 880 69968 139120 70248
rect 197 69568 139970 69968
rect 880 69288 139120 69568
rect 197 68888 139970 69288
rect 880 68608 139120 68888
rect 197 68208 139970 68608
rect 880 67928 139970 68208
rect 197 67528 139970 67928
rect 197 67248 139120 67528
rect 197 66848 139970 67248
rect 880 66568 139120 66848
rect 197 66168 139970 66568
rect 880 65888 139120 66168
rect 197 65488 139970 65888
rect 880 65208 139120 65488
rect 197 64808 139970 65208
rect 880 64528 139120 64808
rect 197 64128 139970 64528
rect 880 63848 139970 64128
rect 197 63448 139970 63848
rect 197 63168 139120 63448
rect 197 62768 139970 63168
rect 880 62488 139120 62768
rect 197 62088 139970 62488
rect 880 61808 139120 62088
rect 197 61408 139970 61808
rect 880 61128 139120 61408
rect 197 60728 139970 61128
rect 880 60448 139120 60728
rect 197 60048 139970 60448
rect 880 59768 139970 60048
rect 197 59368 139970 59768
rect 197 59088 139120 59368
rect 197 58688 139970 59088
rect 880 58408 139120 58688
rect 197 58008 139970 58408
rect 880 57728 139120 58008
rect 197 57328 139970 57728
rect 880 57048 139120 57328
rect 197 56648 139970 57048
rect 880 56368 139120 56648
rect 197 55968 139970 56368
rect 880 55688 139120 55968
rect 197 54608 139970 55688
rect 880 54328 139120 54608
rect 197 53928 139970 54328
rect 880 53648 139120 53928
rect 197 53248 139970 53648
rect 880 52968 139120 53248
rect 197 52568 139970 52968
rect 880 52288 139120 52568
rect 197 51888 139970 52288
rect 880 51608 139120 51888
rect 197 51208 139970 51608
rect 880 50928 139970 51208
rect 197 50528 139970 50928
rect 197 50248 139120 50528
rect 197 49848 139970 50248
rect 880 49568 139120 49848
rect 197 49168 139970 49568
rect 880 48888 139120 49168
rect 197 48488 139970 48888
rect 880 48208 139120 48488
rect 197 47808 139970 48208
rect 880 47528 139120 47808
rect 197 47128 139970 47528
rect 880 46848 139970 47128
rect 197 46448 139970 46848
rect 197 46168 139120 46448
rect 197 45768 139970 46168
rect 880 45488 139120 45768
rect 197 45088 139970 45488
rect 880 44808 139120 45088
rect 197 44408 139970 44808
rect 880 44128 139120 44408
rect 197 43728 139970 44128
rect 880 43448 139120 43728
rect 197 43048 139970 43448
rect 880 42768 139970 43048
rect 197 42368 139970 42768
rect 197 42088 139120 42368
rect 197 41688 139970 42088
rect 880 41408 139120 41688
rect 197 41008 139970 41408
rect 880 40728 139120 41008
rect 197 40328 139970 40728
rect 880 40048 139120 40328
rect 197 39648 139970 40048
rect 880 39368 139120 39648
rect 197 38968 139970 39368
rect 880 38688 139120 38968
rect 197 37608 139970 38688
rect 880 37328 139120 37608
rect 197 36928 139970 37328
rect 880 36648 139120 36928
rect 197 36248 139970 36648
rect 880 35968 139120 36248
rect 197 35568 139970 35968
rect 880 35288 139120 35568
rect 197 34888 139970 35288
rect 880 34608 139120 34888
rect 197 34208 139970 34608
rect 880 33928 139970 34208
rect 197 33528 139970 33928
rect 197 33248 139120 33528
rect 197 32848 139970 33248
rect 880 32568 139120 32848
rect 197 32168 139970 32568
rect 880 31888 139120 32168
rect 197 31488 139970 31888
rect 880 31208 139120 31488
rect 197 30808 139970 31208
rect 880 30528 139120 30808
rect 197 30128 139970 30528
rect 880 29848 139970 30128
rect 197 29448 139970 29848
rect 197 29168 139120 29448
rect 197 28768 139970 29168
rect 880 28488 139120 28768
rect 197 28088 139970 28488
rect 880 27808 139120 28088
rect 197 27408 139970 27808
rect 880 27128 139120 27408
rect 197 26728 139970 27128
rect 880 26448 139120 26728
rect 197 26048 139970 26448
rect 880 25768 139970 26048
rect 197 25368 139970 25768
rect 197 25088 139120 25368
rect 197 24688 139970 25088
rect 880 24408 139120 24688
rect 197 24008 139970 24408
rect 880 23728 139120 24008
rect 197 23328 139970 23728
rect 880 23048 139120 23328
rect 197 22648 139970 23048
rect 880 22368 139120 22648
rect 197 21968 139970 22368
rect 880 21688 139120 21968
rect 197 20608 139970 21688
rect 880 20328 139120 20608
rect 197 19928 139970 20328
rect 880 19648 139120 19928
rect 197 19248 139970 19648
rect 880 18968 139120 19248
rect 197 18568 139970 18968
rect 880 18288 139120 18568
rect 197 17888 139970 18288
rect 880 17608 139120 17888
rect 197 17208 139970 17608
rect 880 16928 139970 17208
rect 197 16528 139970 16928
rect 197 16248 139120 16528
rect 197 15848 139970 16248
rect 880 15568 139120 15848
rect 197 15168 139970 15568
rect 880 14888 139120 15168
rect 197 14488 139970 14888
rect 880 14208 139120 14488
rect 197 13808 139970 14208
rect 880 13528 139120 13808
rect 197 13128 139970 13528
rect 880 12848 139970 13128
rect 197 12448 139970 12848
rect 197 12168 139120 12448
rect 197 11768 139970 12168
rect 880 11488 139120 11768
rect 197 11088 139970 11488
rect 880 10808 139120 11088
rect 197 10408 139970 10808
rect 880 10128 139120 10408
rect 197 9728 139970 10128
rect 880 9448 139120 9728
rect 197 9048 139970 9448
rect 880 8768 139970 9048
rect 197 8368 139970 8768
rect 197 8088 139120 8368
rect 197 7688 139970 8088
rect 880 7408 139120 7688
rect 197 7008 139970 7408
rect 880 6728 139120 7008
rect 197 6328 139970 6728
rect 880 6048 139120 6328
rect 197 5648 139970 6048
rect 880 5368 139120 5648
rect 197 4968 139970 5368
rect 880 4688 139120 4968
rect 197 3608 139970 4688
rect 880 3328 139120 3608
rect 197 2928 139970 3328
rect 880 2648 139120 2928
rect 197 2248 139970 2648
rect 880 1968 139120 2248
rect 197 1568 139970 1968
rect 880 1288 139120 1568
rect 197 888 139970 1288
rect 880 715 139120 888
<< metal4 >>
rect 4208 2128 4528 437424
rect 19568 2128 19888 437424
rect 34928 2128 35248 437424
rect 50288 2128 50608 437424
rect 65648 2128 65968 437424
rect 81008 2128 81328 437424
rect 96368 2128 96688 437424
rect 111728 2128 112048 437424
rect 127088 2128 127408 437424
<< obsm4 >>
rect 427 2048 4128 437205
rect 4608 2048 19488 437205
rect 19968 2048 34848 437205
rect 35328 2048 50208 437205
rect 50688 2048 65568 437205
rect 66048 2048 80928 437205
rect 81408 2048 96288 437205
rect 96768 2048 111648 437205
rect 112128 2048 127008 437205
rect 127488 2048 139965 437205
rect 427 1667 139965 2048
<< labels >>
rlabel metal2 s 124310 439200 124366 440000 6 axi_spi_master_ar_addr[0]
port 1 nsew signal output
rlabel metal3 s 0 312808 800 312928 6 axi_spi_master_ar_addr[10]
port 2 nsew signal output
rlabel metal3 s 0 17688 800 17808 6 axi_spi_master_ar_addr[11]
port 3 nsew signal output
rlabel metal3 s 139200 36048 140000 36168 6 axi_spi_master_ar_addr[12]
port 4 nsew signal output
rlabel metal3 s 139200 197888 140000 198008 6 axi_spi_master_ar_addr[13]
port 5 nsew signal output
rlabel metal2 s 51538 0 51594 800 6 axi_spi_master_ar_addr[14]
port 6 nsew signal output
rlabel metal3 s 0 71408 800 71528 6 axi_spi_master_ar_addr[15]
port 7 nsew signal output
rlabel metal2 s 86958 0 87014 800 6 axi_spi_master_ar_addr[16]
port 8 nsew signal output
rlabel metal3 s 139200 410728 140000 410848 6 axi_spi_master_ar_addr[17]
port 9 nsew signal output
rlabel metal3 s 0 129208 800 129328 6 axi_spi_master_ar_addr[18]
port 10 nsew signal output
rlabel metal3 s 0 341368 800 341488 6 axi_spi_master_ar_addr[19]
port 11 nsew signal output
rlabel metal3 s 0 53728 800 53848 6 axi_spi_master_ar_addr[1]
port 12 nsew signal output
rlabel metal2 s 139122 439200 139178 440000 6 axi_spi_master_ar_addr[20]
port 13 nsew signal output
rlabel metal3 s 0 382848 800 382968 6 axi_spi_master_ar_addr[21]
port 14 nsew signal output
rlabel metal3 s 139200 327768 140000 327888 6 axi_spi_master_ar_addr[22]
port 15 nsew signal output
rlabel metal3 s 139200 22448 140000 22568 6 axi_spi_master_ar_addr[23]
port 16 nsew signal output
rlabel metal3 s 139200 141448 140000 141568 6 axi_spi_master_ar_addr[24]
port 17 nsew signal output
rlabel metal3 s 0 209448 800 209568 6 axi_spi_master_ar_addr[25]
port 18 nsew signal output
rlabel metal2 s 102414 439200 102470 440000 6 axi_spi_master_ar_addr[26]
port 19 nsew signal output
rlabel metal3 s 139200 57808 140000 57928 6 axi_spi_master_ar_addr[27]
port 20 nsew signal output
rlabel metal2 s 70214 439200 70270 440000 6 axi_spi_master_ar_addr[28]
port 21 nsew signal output
rlabel metal3 s 0 354968 800 355088 6 axi_spi_master_ar_addr[29]
port 22 nsew signal output
rlabel metal2 s 46386 0 46442 800 6 axi_spi_master_ar_addr[2]
port 23 nsew signal output
rlabel metal3 s 139200 113568 140000 113688 6 axi_spi_master_ar_addr[30]
port 24 nsew signal output
rlabel metal2 s 115294 439200 115350 440000 6 axi_spi_master_ar_addr[31]
port 25 nsew signal output
rlabel metal3 s 0 111528 800 111648 6 axi_spi_master_ar_addr[3]
port 26 nsew signal output
rlabel metal2 s 48962 439200 49018 440000 6 axi_spi_master_ar_addr[4]
port 27 nsew signal output
rlabel metal2 s 85026 439200 85082 440000 6 axi_spi_master_ar_addr[5]
port 28 nsew signal output
rlabel metal3 s 0 102688 800 102808 6 axi_spi_master_ar_addr[6]
port 29 nsew signal output
rlabel metal3 s 139200 376048 140000 376168 6 axi_spi_master_ar_addr[7]
port 30 nsew signal output
rlabel metal2 s 135258 439200 135314 440000 6 axi_spi_master_ar_addr[8]
port 31 nsew signal output
rlabel metal3 s 139200 129208 140000 129328 6 axi_spi_master_ar_addr[9]
port 32 nsew signal output
rlabel metal3 s 0 180208 800 180328 6 axi_spi_master_ar_burst[0]
port 33 nsew signal output
rlabel metal2 s 120446 439200 120502 440000 6 axi_spi_master_ar_burst[1]
port 34 nsew signal output
rlabel metal2 s 78586 0 78642 800 6 axi_spi_master_ar_cache[0]
port 35 nsew signal output
rlabel metal3 s 0 113568 800 113688 6 axi_spi_master_ar_cache[1]
port 36 nsew signal output
rlabel metal3 s 139200 437928 140000 438048 6 axi_spi_master_ar_cache[2]
port 37 nsew signal output
rlabel metal3 s 0 387608 800 387728 6 axi_spi_master_ar_cache[3]
port 38 nsew signal output
rlabel metal3 s 139200 418888 140000 419008 6 axi_spi_master_ar_id[0]
port 39 nsew signal output
rlabel metal3 s 139200 90448 140000 90568 6 axi_spi_master_ar_id[1]
port 40 nsew signal output
rlabel metal3 s 139200 91808 140000 91928 6 axi_spi_master_ar_id[2]
port 41 nsew signal output
rlabel metal3 s 139200 104728 140000 104848 6 axi_spi_master_ar_id[3]
port 42 nsew signal output
rlabel metal3 s 139200 249568 140000 249688 6 axi_spi_master_ar_id[4]
port 43 nsew signal output
rlabel metal3 s 0 369928 800 370048 6 axi_spi_master_ar_id[5]
port 44 nsew signal output
rlabel metal3 s 0 234608 800 234728 6 axi_spi_master_ar_len[0]
port 45 nsew signal output
rlabel metal3 s 139200 7488 140000 7608 6 axi_spi_master_ar_len[1]
port 46 nsew signal output
rlabel metal3 s 0 289008 800 289128 6 axi_spi_master_ar_len[2]
port 47 nsew signal output
rlabel metal2 s 88890 0 88946 800 6 axi_spi_master_ar_len[3]
port 48 nsew signal output
rlabel metal3 s 139200 26528 140000 26648 6 axi_spi_master_ar_len[4]
port 49 nsew signal output
rlabel metal3 s 0 238008 800 238128 6 axi_spi_master_ar_len[5]
port 50 nsew signal output
rlabel metal2 s 1306 0 1362 800 6 axi_spi_master_ar_len[6]
port 51 nsew signal output
rlabel metal3 s 0 252968 800 253088 6 axi_spi_master_ar_len[7]
port 52 nsew signal output
rlabel metal3 s 0 187688 800 187808 6 axi_spi_master_ar_lock
port 53 nsew signal output
rlabel metal3 s 139200 30608 140000 30728 6 axi_spi_master_ar_prot[0]
port 54 nsew signal output
rlabel metal3 s 139200 405968 140000 406088 6 axi_spi_master_ar_prot[1]
port 55 nsew signal output
rlabel metal3 s 0 27888 800 28008 6 axi_spi_master_ar_prot[2]
port 56 nsew signal output
rlabel metal3 s 0 412768 800 412888 6 axi_spi_master_ar_qos[0]
port 57 nsew signal output
rlabel metal3 s 139200 210128 140000 210248 6 axi_spi_master_ar_qos[1]
port 58 nsew signal output
rlabel metal3 s 0 248888 800 249008 6 axi_spi_master_ar_qos[2]
port 59 nsew signal output
rlabel metal3 s 139200 438608 140000 438728 6 axi_spi_master_ar_qos[3]
port 60 nsew signal output
rlabel metal2 s 74722 439200 74778 440000 6 axi_spi_master_ar_ready
port 61 nsew signal input
rlabel metal3 s 0 199928 800 200048 6 axi_spi_master_ar_region[0]
port 62 nsew signal output
rlabel metal3 s 139200 229848 140000 229968 6 axi_spi_master_ar_region[1]
port 63 nsew signal output
rlabel metal3 s 139200 126488 140000 126608 6 axi_spi_master_ar_region[2]
port 64 nsew signal output
rlabel metal3 s 0 295128 800 295248 6 axi_spi_master_ar_region[3]
port 65 nsew signal output
rlabel metal3 s 139200 362448 140000 362568 6 axi_spi_master_ar_size[0]
port 66 nsew signal output
rlabel metal3 s 139200 416848 140000 416968 6 axi_spi_master_ar_size[1]
port 67 nsew signal output
rlabel metal3 s 139200 180208 140000 180328 6 axi_spi_master_ar_size[2]
port 68 nsew signal output
rlabel metal2 s 128818 0 128874 800 6 axi_spi_master_ar_user[0]
port 69 nsew signal output
rlabel metal3 s 0 45568 800 45688 6 axi_spi_master_ar_user[1]
port 70 nsew signal output
rlabel metal3 s 139200 375368 140000 375488 6 axi_spi_master_ar_user[2]
port 71 nsew signal output
rlabel metal3 s 0 154368 800 154488 6 axi_spi_master_ar_user[3]
port 72 nsew signal output
rlabel metal3 s 0 139408 800 139528 6 axi_spi_master_ar_user[4]
port 73 nsew signal output
rlabel metal2 s 137190 0 137246 800 6 axi_spi_master_ar_user[5]
port 74 nsew signal output
rlabel metal3 s 139200 391688 140000 391808 6 axi_spi_master_ar_valid
port 75 nsew signal output
rlabel metal3 s 0 109488 800 109608 6 axi_spi_master_aw_addr[0]
port 76 nsew signal output
rlabel metal3 s 139200 86368 140000 86488 6 axi_spi_master_aw_addr[10]
port 77 nsew signal output
rlabel metal3 s 0 171368 800 171488 6 axi_spi_master_aw_addr[11]
port 78 nsew signal output
rlabel metal2 s 86314 439200 86370 440000 6 axi_spi_master_aw_addr[12]
port 79 nsew signal output
rlabel metal2 s 123022 439200 123078 440000 6 axi_spi_master_aw_addr[13]
port 80 nsew signal output
rlabel metal2 s 135902 439200 135958 440000 6 axi_spi_master_aw_addr[14]
port 81 nsew signal output
rlabel metal2 s 79230 0 79286 800 6 axi_spi_master_aw_addr[15]
port 82 nsew signal output
rlabel metal3 s 139200 299888 140000 300008 6 axi_spi_master_aw_addr[16]
port 83 nsew signal output
rlabel metal3 s 0 48968 800 49088 6 axi_spi_master_aw_addr[17]
port 84 nsew signal output
rlabel metal2 s 97906 0 97962 800 6 axi_spi_master_aw_addr[18]
port 85 nsew signal output
rlabel metal3 s 139200 118328 140000 118448 6 axi_spi_master_aw_addr[19]
port 86 nsew signal output
rlabel metal2 s 56690 439200 56746 440000 6 axi_spi_master_aw_addr[1]
port 87 nsew signal output
rlabel metal3 s 139200 374688 140000 374808 6 axi_spi_master_aw_addr[20]
port 88 nsew signal output
rlabel metal2 s 10966 0 11022 800 6 axi_spi_master_aw_addr[21]
port 89 nsew signal output
rlabel metal2 s 124954 439200 125010 440000 6 axi_spi_master_aw_addr[22]
port 90 nsew signal output
rlabel metal3 s 0 367208 800 367328 6 axi_spi_master_aw_addr[23]
port 91 nsew signal output
rlabel metal2 s 114006 0 114062 800 6 axi_spi_master_aw_addr[24]
port 92 nsew signal output
rlabel metal3 s 0 243448 800 243568 6 axi_spi_master_aw_addr[25]
port 93 nsew signal output
rlabel metal3 s 0 214888 800 215008 6 axi_spi_master_aw_addr[26]
port 94 nsew signal output
rlabel metal3 s 0 160488 800 160608 6 axi_spi_master_aw_addr[27]
port 95 nsew signal output
rlabel metal3 s 0 359048 800 359168 6 axi_spi_master_aw_addr[28]
port 96 nsew signal output
rlabel metal2 s 45098 439200 45154 440000 6 axi_spi_master_aw_addr[29]
port 97 nsew signal output
rlabel metal3 s 139200 325048 140000 325168 6 axi_spi_master_aw_addr[2]
port 98 nsew signal output
rlabel metal3 s 0 371288 800 371408 6 axi_spi_master_aw_addr[30]
port 99 nsew signal output
rlabel metal2 s 67638 0 67694 800 6 axi_spi_master_aw_addr[31]
port 100 nsew signal output
rlabel metal3 s 139200 235288 140000 235408 6 axi_spi_master_aw_addr[3]
port 101 nsew signal output
rlabel metal3 s 0 10888 800 11008 6 axi_spi_master_aw_addr[4]
port 102 nsew signal output
rlabel metal3 s 139200 351568 140000 351688 6 axi_spi_master_aw_addr[5]
port 103 nsew signal output
rlabel metal3 s 0 385568 800 385688 6 axi_spi_master_aw_addr[6]
port 104 nsew signal output
rlabel metal3 s 0 393728 800 393848 6 axi_spi_master_aw_addr[7]
port 105 nsew signal output
rlabel metal3 s 0 22448 800 22568 6 axi_spi_master_aw_addr[8]
port 106 nsew signal output
rlabel metal3 s 0 138728 800 138848 6 axi_spi_master_aw_addr[9]
port 107 nsew signal output
rlabel metal2 s 108854 439200 108910 440000 6 axi_spi_master_aw_burst[0]
port 108 nsew signal output
rlabel metal3 s 0 207408 800 207528 6 axi_spi_master_aw_burst[1]
port 109 nsew signal output
rlabel metal3 s 0 138048 800 138168 6 axi_spi_master_aw_cache[0]
port 110 nsew signal output
rlabel metal3 s 139200 303968 140000 304088 6 axi_spi_master_aw_cache[1]
port 111 nsew signal output
rlabel metal3 s 0 361088 800 361208 6 axi_spi_master_aw_cache[2]
port 112 nsew signal output
rlabel metal3 s 139200 219648 140000 219768 6 axi_spi_master_aw_cache[3]
port 113 nsew signal output
rlabel metal3 s 139200 277448 140000 277568 6 axi_spi_master_aw_id[0]
port 114 nsew signal output
rlabel metal3 s 0 376048 800 376168 6 axi_spi_master_aw_id[1]
port 115 nsew signal output
rlabel metal3 s 139200 376728 140000 376848 6 axi_spi_master_aw_id[2]
port 116 nsew signal output
rlabel metal3 s 139200 179528 140000 179648 6 axi_spi_master_aw_id[3]
port 117 nsew signal output
rlabel metal3 s 139200 407328 140000 407448 6 axi_spi_master_aw_id[4]
port 118 nsew signal output
rlabel metal3 s 139200 243448 140000 243568 6 axi_spi_master_aw_id[5]
port 119 nsew signal output
rlabel metal3 s 139200 208768 140000 208888 6 axi_spi_master_aw_len[0]
port 120 nsew signal output
rlabel metal3 s 0 364488 800 364608 6 axi_spi_master_aw_len[1]
port 121 nsew signal output
rlabel metal3 s 0 83648 800 83768 6 axi_spi_master_aw_len[2]
port 122 nsew signal output
rlabel metal3 s 139200 401208 140000 401328 6 axi_spi_master_aw_len[3]
port 123 nsew signal output
rlabel metal3 s 0 75488 800 75608 6 axi_spi_master_aw_len[4]
port 124 nsew signal output
rlabel metal3 s 139200 148248 140000 148368 6 axi_spi_master_aw_len[5]
port 125 nsew signal output
rlabel metal3 s 139200 28568 140000 28688 6 axi_spi_master_aw_len[6]
port 126 nsew signal output
rlabel metal3 s 0 212848 800 212968 6 axi_spi_master_aw_len[7]
port 127 nsew signal output
rlabel metal3 s 139200 291048 140000 291168 6 axi_spi_master_aw_lock
port 128 nsew signal output
rlabel metal2 s 59266 0 59322 800 6 axi_spi_master_aw_prot[0]
port 129 nsew signal output
rlabel metal3 s 139200 408688 140000 408808 6 axi_spi_master_aw_prot[1]
port 130 nsew signal output
rlabel metal2 s 133970 0 134026 800 6 axi_spi_master_aw_prot[2]
port 131 nsew signal output
rlabel metal2 s 60554 439200 60610 440000 6 axi_spi_master_aw_qos[0]
port 132 nsew signal output
rlabel metal3 s 0 397808 800 397928 6 axi_spi_master_aw_qos[1]
port 133 nsew signal output
rlabel metal2 s 30286 439200 30342 440000 6 axi_spi_master_aw_qos[2]
port 134 nsew signal output
rlabel metal2 s 117870 0 117926 800 6 axi_spi_master_aw_qos[3]
port 135 nsew signal output
rlabel metal3 s 0 195848 800 195968 6 axi_spi_master_aw_ready
port 136 nsew signal input
rlabel metal2 s 115294 0 115350 800 6 axi_spi_master_aw_region[0]
port 137 nsew signal output
rlabel metal3 s 0 92488 800 92608 6 axi_spi_master_aw_region[1]
port 138 nsew signal output
rlabel metal3 s 139200 232568 140000 232688 6 axi_spi_master_aw_region[2]
port 139 nsew signal output
rlabel metal2 s 134614 0 134670 800 6 axi_spi_master_aw_region[3]
port 140 nsew signal output
rlabel metal3 s 0 141448 800 141568 6 axi_spi_master_aw_size[0]
port 141 nsew signal output
rlabel metal3 s 0 95208 800 95328 6 axi_spi_master_aw_size[1]
port 142 nsew signal output
rlabel metal3 s 139200 114248 140000 114368 6 axi_spi_master_aw_size[2]
port 143 nsew signal output
rlabel metal2 s 106278 439200 106334 440000 6 axi_spi_master_aw_user[0]
port 144 nsew signal output
rlabel metal3 s 139200 350208 140000 350328 6 axi_spi_master_aw_user[1]
port 145 nsew signal output
rlabel metal3 s 0 172728 800 172848 6 axi_spi_master_aw_user[2]
port 146 nsew signal output
rlabel metal3 s 0 259088 800 259208 6 axi_spi_master_aw_user[3]
port 147 nsew signal output
rlabel metal2 s 133326 439200 133382 440000 6 axi_spi_master_aw_user[4]
port 148 nsew signal output
rlabel metal3 s 139200 44208 140000 44328 6 axi_spi_master_aw_user[5]
port 149 nsew signal output
rlabel metal2 s 52826 439200 52882 440000 6 axi_spi_master_aw_valid
port 150 nsew signal output
rlabel metal3 s 139200 353608 140000 353728 6 axi_spi_master_b_id[0]
port 151 nsew signal input
rlabel metal3 s 139200 221688 140000 221808 6 axi_spi_master_b_id[1]
port 152 nsew signal input
rlabel metal3 s 139200 29248 140000 29368 6 axi_spi_master_b_id[2]
port 153 nsew signal input
rlabel metal2 s 96618 439200 96674 440000 6 axi_spi_master_b_id[3]
port 154 nsew signal input
rlabel metal3 s 0 192448 800 192568 6 axi_spi_master_b_id[4]
port 155 nsew signal input
rlabel metal3 s 0 265888 800 266008 6 axi_spi_master_b_id[5]
port 156 nsew signal input
rlabel metal3 s 0 293768 800 293888 6 axi_spi_master_b_ready
port 157 nsew signal output
rlabel metal2 s 42522 0 42578 800 6 axi_spi_master_b_resp[0]
port 158 nsew signal input
rlabel metal3 s 139200 278808 140000 278928 6 axi_spi_master_b_resp[1]
port 159 nsew signal input
rlabel metal2 s 38658 439200 38714 440000 6 axi_spi_master_b_user[0]
port 160 nsew signal input
rlabel metal3 s 0 176808 800 176928 6 axi_spi_master_b_user[1]
port 161 nsew signal input
rlabel metal3 s 139200 99288 140000 99408 6 axi_spi_master_b_user[2]
port 162 nsew signal input
rlabel metal2 s 110786 0 110842 800 6 axi_spi_master_b_user[3]
port 163 nsew signal input
rlabel metal3 s 0 240728 800 240848 6 axi_spi_master_b_user[4]
port 164 nsew signal input
rlabel metal2 s 83738 439200 83794 440000 6 axi_spi_master_b_user[5]
port 165 nsew signal input
rlabel metal3 s 0 325728 800 325848 6 axi_spi_master_b_valid
port 166 nsew signal input
rlabel metal2 s 41234 0 41290 800 6 axi_spi_master_r_data[0]
port 167 nsew signal input
rlabel metal3 s 139200 207408 140000 207528 6 axi_spi_master_r_data[10]
port 168 nsew signal input
rlabel metal3 s 139200 31968 140000 32088 6 axi_spi_master_r_data[11]
port 169 nsew signal input
rlabel metal3 s 139200 84328 140000 84448 6 axi_spi_master_r_data[12]
port 170 nsew signal input
rlabel metal3 s 139200 343408 140000 343528 6 axi_spi_master_r_data[13]
port 171 nsew signal input
rlabel metal3 s 0 438608 800 438728 6 axi_spi_master_r_data[14]
port 172 nsew signal input
rlabel metal2 s 1950 0 2006 800 6 axi_spi_master_r_data[15]
port 173 nsew signal input
rlabel metal3 s 0 422968 800 423088 6 axi_spi_master_r_data[16]
port 174 nsew signal input
rlabel metal3 s 139200 424328 140000 424448 6 axi_spi_master_r_data[17]
port 175 nsew signal input
rlabel metal3 s 0 230528 800 230648 6 axi_spi_master_r_data[18]
port 176 nsew signal input
rlabel metal2 s 68926 439200 68982 440000 6 axi_spi_master_r_data[19]
port 177 nsew signal input
rlabel metal3 s 0 126488 800 126608 6 axi_spi_master_r_data[1]
port 178 nsew signal input
rlabel metal3 s 139200 271328 140000 271448 6 axi_spi_master_r_data[20]
port 179 nsew signal input
rlabel metal2 s 11610 439200 11666 440000 6 axi_spi_master_r_data[21]
port 180 nsew signal input
rlabel metal3 s 139200 176808 140000 176928 6 axi_spi_master_r_data[22]
port 181 nsew signal input
rlabel metal3 s 0 291048 800 291168 6 axi_spi_master_r_data[23]
port 182 nsew signal input
rlabel metal2 s 132682 439200 132738 440000 6 axi_spi_master_r_data[24]
port 183 nsew signal input
rlabel metal2 s 121734 0 121790 800 6 axi_spi_master_r_data[25]
port 184 nsew signal input
rlabel metal3 s 139200 88408 140000 88528 6 axi_spi_master_r_data[26]
port 185 nsew signal input
rlabel metal3 s 0 371968 800 372088 6 axi_spi_master_r_data[27]
port 186 nsew signal input
rlabel metal3 s 0 308048 800 308168 6 axi_spi_master_r_data[28]
port 187 nsew signal input
rlabel metal3 s 0 357688 800 357808 6 axi_spi_master_r_data[29]
port 188 nsew signal input
rlabel metal3 s 139200 78888 140000 79008 6 axi_spi_master_r_data[2]
port 189 nsew signal input
rlabel metal3 s 139200 44888 140000 45008 6 axi_spi_master_r_data[30]
port 190 nsew signal input
rlabel metal2 s 130106 0 130162 800 6 axi_spi_master_r_data[31]
port 191 nsew signal input
rlabel metal3 s 139200 349528 140000 349648 6 axi_spi_master_r_data[32]
port 192 nsew signal input
rlabel metal3 s 139200 134648 140000 134768 6 axi_spi_master_r_data[33]
port 193 nsew signal input
rlabel metal3 s 139200 177488 140000 177608 6 axi_spi_master_r_data[34]
port 194 nsew signal input
rlabel metal2 s 34150 439200 34206 440000 6 axi_spi_master_r_data[35]
port 195 nsew signal input
rlabel metal3 s 139200 108128 140000 108248 6 axi_spi_master_r_data[36]
port 196 nsew signal input
rlabel metal3 s 0 299208 800 299328 6 axi_spi_master_r_data[37]
port 197 nsew signal input
rlabel metal3 s 0 327088 800 327208 6 axi_spi_master_r_data[38]
port 198 nsew signal input
rlabel metal3 s 139200 272688 140000 272808 6 axi_spi_master_r_data[39]
port 199 nsew signal input
rlabel metal3 s 139200 247528 140000 247648 6 axi_spi_master_r_data[3]
port 200 nsew signal input
rlabel metal3 s 0 349528 800 349648 6 axi_spi_master_r_data[40]
port 201 nsew signal input
rlabel metal2 s 81806 0 81862 800 6 axi_spi_master_r_data[41]
port 202 nsew signal input
rlabel metal2 s 56690 0 56746 800 6 axi_spi_master_r_data[42]
port 203 nsew signal input
rlabel metal3 s 139200 59168 140000 59288 6 axi_spi_master_r_data[43]
port 204 nsew signal input
rlabel metal3 s 139200 257728 140000 257848 6 axi_spi_master_r_data[44]
port 205 nsew signal input
rlabel metal3 s 0 389648 800 389768 6 axi_spi_master_r_data[45]
port 206 nsew signal input
rlabel metal3 s 0 399848 800 399968 6 axi_spi_master_r_data[46]
port 207 nsew signal input
rlabel metal2 s 84382 439200 84438 440000 6 axi_spi_master_r_data[47]
port 208 nsew signal input
rlabel metal3 s 0 400528 800 400648 6 axi_spi_master_r_data[48]
port 209 nsew signal input
rlabel metal3 s 0 127848 800 127968 6 axi_spi_master_r_data[49]
port 210 nsew signal input
rlabel metal3 s 139200 323688 140000 323808 6 axi_spi_master_r_data[4]
port 211 nsew signal input
rlabel metal3 s 0 393048 800 393168 6 axi_spi_master_r_data[50]
port 212 nsew signal input
rlabel metal3 s 0 162528 800 162648 6 axi_spi_master_r_data[51]
port 213 nsew signal input
rlabel metal3 s 0 434528 800 434648 6 axi_spi_master_r_data[52]
port 214 nsew signal input
rlabel metal3 s 0 378088 800 378208 6 axi_spi_master_r_data[53]
port 215 nsew signal input
rlabel metal3 s 139200 388968 140000 389088 6 axi_spi_master_r_data[54]
port 216 nsew signal input
rlabel metal3 s 0 115608 800 115728 6 axi_spi_master_r_data[55]
port 217 nsew signal input
rlabel metal3 s 0 436568 800 436688 6 axi_spi_master_r_data[56]
port 218 nsew signal input
rlabel metal3 s 139200 397128 140000 397248 6 axi_spi_master_r_data[57]
port 219 nsew signal input
rlabel metal3 s 0 204008 800 204128 6 axi_spi_master_r_data[58]
port 220 nsew signal input
rlabel metal3 s 0 405968 800 406088 6 axi_spi_master_r_data[59]
port 221 nsew signal input
rlabel metal3 s 0 366528 800 366648 6 axi_spi_master_r_data[5]
port 222 nsew signal input
rlabel metal3 s 0 25848 800 25968 6 axi_spi_master_r_data[60]
port 223 nsew signal input
rlabel metal2 s 67638 439200 67694 440000 6 axi_spi_master_r_data[61]
port 224 nsew signal input
rlabel metal3 s 139200 274048 140000 274168 6 axi_spi_master_r_data[62]
port 225 nsew signal input
rlabel metal2 s 27066 439200 27122 440000 6 axi_spi_master_r_data[63]
port 226 nsew signal input
rlabel metal3 s 0 347488 800 347608 6 axi_spi_master_r_data[6]
port 227 nsew signal input
rlabel metal3 s 0 329128 800 329248 6 axi_spi_master_r_data[7]
port 228 nsew signal input
rlabel metal3 s 139200 158448 140000 158568 6 axi_spi_master_r_data[8]
port 229 nsew signal input
rlabel metal2 s 83738 0 83794 800 6 axi_spi_master_r_data[9]
port 230 nsew signal input
rlabel metal3 s 139200 383528 140000 383648 6 axi_spi_master_r_id[0]
port 231 nsew signal input
rlabel metal3 s 0 108808 800 108928 6 axi_spi_master_r_id[1]
port 232 nsew signal input
rlabel metal3 s 139200 366528 140000 366648 6 axi_spi_master_r_id[2]
port 233 nsew signal input
rlabel metal2 s 103702 439200 103758 440000 6 axi_spi_master_r_id[3]
port 234 nsew signal input
rlabel metal2 s 123666 0 123722 800 6 axi_spi_master_r_id[4]
port 235 nsew signal input
rlabel metal3 s 0 321648 800 321768 6 axi_spi_master_r_id[5]
port 236 nsew signal input
rlabel metal2 s 90822 0 90878 800 6 axi_spi_master_r_last
port 237 nsew signal input
rlabel metal3 s 139200 130568 140000 130688 6 axi_spi_master_r_ready
port 238 nsew signal output
rlabel metal3 s 139200 405288 140000 405408 6 axi_spi_master_r_resp[0]
port 239 nsew signal input
rlabel metal3 s 0 36728 800 36848 6 axi_spi_master_r_resp[1]
port 240 nsew signal input
rlabel metal3 s 139200 58488 140000 58608 6 axi_spi_master_r_user[0]
port 241 nsew signal input
rlabel metal3 s 139200 273368 140000 273488 6 axi_spi_master_r_user[1]
port 242 nsew signal input
rlabel metal2 s 85026 0 85082 800 6 axi_spi_master_r_user[2]
port 243 nsew signal input
rlabel metal3 s 0 184288 800 184408 6 axi_spi_master_r_user[3]
port 244 nsew signal input
rlabel metal3 s 139200 171368 140000 171488 6 axi_spi_master_r_user[4]
port 245 nsew signal input
rlabel metal3 s 139200 62568 140000 62688 6 axi_spi_master_r_user[5]
port 246 nsew signal input
rlabel metal3 s 0 405288 800 405408 6 axi_spi_master_r_valid
port 247 nsew signal input
rlabel metal2 s 83094 439200 83150 440000 6 axi_spi_master_w_data[0]
port 248 nsew signal output
rlabel metal3 s 139200 380808 140000 380928 6 axi_spi_master_w_data[10]
port 249 nsew signal output
rlabel metal3 s 0 396448 800 396568 6 axi_spi_master_w_data[11]
port 250 nsew signal output
rlabel metal3 s 0 205368 800 205488 6 axi_spi_master_w_data[12]
port 251 nsew signal output
rlabel metal2 s 65706 0 65762 800 6 axi_spi_master_w_data[13]
port 252 nsew signal output
rlabel metal2 s 50250 439200 50306 440000 6 axi_spi_master_w_data[14]
port 253 nsew signal output
rlabel metal3 s 0 159808 800 159928 6 axi_spi_master_w_data[15]
port 254 nsew signal output
rlabel metal3 s 0 28568 800 28688 6 axi_spi_master_w_data[16]
port 255 nsew signal output
rlabel metal3 s 139200 354288 140000 354408 6 axi_spi_master_w_data[17]
port 256 nsew signal output
rlabel metal2 s 8390 439200 8446 440000 6 axi_spi_master_w_data[18]
port 257 nsew signal output
rlabel metal3 s 139200 185648 140000 185768 6 axi_spi_master_w_data[19]
port 258 nsew signal output
rlabel metal3 s 0 331848 800 331968 6 axi_spi_master_w_data[1]
port 259 nsew signal output
rlabel metal3 s 139200 56448 140000 56568 6 axi_spi_master_w_data[20]
port 260 nsew signal output
rlabel metal2 s 7746 439200 7802 440000 6 axi_spi_master_w_data[21]
port 261 nsew signal output
rlabel metal3 s 139200 166608 140000 166728 6 axi_spi_master_w_data[22]
port 262 nsew signal output
rlabel metal3 s 0 312128 800 312248 6 axi_spi_master_w_data[23]
port 263 nsew signal output
rlabel metal2 s 76010 439200 76066 440000 6 axi_spi_master_w_data[24]
port 264 nsew signal output
rlabel metal3 s 139200 415488 140000 415608 6 axi_spi_master_w_data[25]
port 265 nsew signal output
rlabel metal3 s 139200 395768 140000 395888 6 axi_spi_master_w_data[26]
port 266 nsew signal output
rlabel metal3 s 0 253648 800 253768 6 axi_spi_master_w_data[27]
port 267 nsew signal output
rlabel metal3 s 0 107448 800 107568 6 axi_spi_master_w_data[28]
port 268 nsew signal output
rlabel metal3 s 139200 223728 140000 223848 6 axi_spi_master_w_data[29]
port 269 nsew signal output
rlabel metal3 s 139200 154368 140000 154488 6 axi_spi_master_w_data[2]
port 270 nsew signal output
rlabel metal3 s 139200 303288 140000 303408 6 axi_spi_master_w_data[30]
port 271 nsew signal output
rlabel metal3 s 0 300568 800 300688 6 axi_spi_master_w_data[31]
port 272 nsew signal output
rlabel metal3 s 0 248208 800 248328 6 axi_spi_master_w_data[32]
port 273 nsew signal output
rlabel metal3 s 139200 105408 140000 105528 6 axi_spi_master_w_data[33]
port 274 nsew signal output
rlabel metal2 s 30930 0 30986 800 6 axi_spi_master_w_data[34]
port 275 nsew signal output
rlabel metal3 s 139200 204688 140000 204808 6 axi_spi_master_w_data[35]
port 276 nsew signal output
rlabel metal3 s 139200 161848 140000 161968 6 axi_spi_master_w_data[36]
port 277 nsew signal output
rlabel metal2 s 52182 439200 52238 440000 6 axi_spi_master_w_data[37]
port 278 nsew signal output
rlabel metal3 s 139200 298528 140000 298648 6 axi_spi_master_w_data[38]
port 279 nsew signal output
rlabel metal3 s 0 290368 800 290488 6 axi_spi_master_w_data[39]
port 280 nsew signal output
rlabel metal3 s 0 391008 800 391128 6 axi_spi_master_w_data[3]
port 281 nsew signal output
rlabel metal3 s 0 125128 800 125248 6 axi_spi_master_w_data[40]
port 282 nsew signal output
rlabel metal3 s 139200 379448 140000 379568 6 axi_spi_master_w_data[41]
port 283 nsew signal output
rlabel metal2 s 125598 0 125654 800 6 axi_spi_master_w_data[42]
port 284 nsew signal output
rlabel metal3 s 139200 159808 140000 159928 6 axi_spi_master_w_data[43]
port 285 nsew signal output
rlabel metal3 s 139200 325728 140000 325848 6 axi_spi_master_w_data[44]
port 286 nsew signal output
rlabel metal3 s 0 231208 800 231328 6 axi_spi_master_w_data[45]
port 287 nsew signal output
rlabel metal2 s 76654 0 76710 800 6 axi_spi_master_w_data[46]
port 288 nsew signal output
rlabel metal3 s 139200 124448 140000 124568 6 axi_spi_master_w_data[47]
port 289 nsew signal output
rlabel metal3 s 139200 199248 140000 199368 6 axi_spi_master_w_data[48]
port 290 nsew signal output
rlabel metal2 s 46386 439200 46442 440000 6 axi_spi_master_w_data[49]
port 291 nsew signal output
rlabel metal3 s 0 184968 800 185088 6 axi_spi_master_w_data[4]
port 292 nsew signal output
rlabel metal3 s 0 210128 800 210248 6 axi_spi_master_w_data[50]
port 293 nsew signal output
rlabel metal3 s 0 74808 800 74928 6 axi_spi_master_w_data[51]
port 294 nsew signal output
rlabel metal3 s 0 279488 800 279608 6 axi_spi_master_w_data[52]
port 295 nsew signal output
rlabel metal3 s 0 294448 800 294568 6 axi_spi_master_w_data[53]
port 296 nsew signal output
rlabel metal2 s 111430 0 111486 800 6 axi_spi_master_w_data[54]
port 297 nsew signal output
rlabel metal3 s 0 280848 800 280968 6 axi_spi_master_w_data[55]
port 298 nsew signal output
rlabel metal3 s 0 302608 800 302728 6 axi_spi_master_w_data[56]
port 299 nsew signal output
rlabel metal3 s 139200 289688 140000 289808 6 axi_spi_master_w_data[57]
port 300 nsew signal output
rlabel metal3 s 0 86368 800 86488 6 axi_spi_master_w_data[58]
port 301 nsew signal output
rlabel metal2 s 65062 439200 65118 440000 6 axi_spi_master_w_data[59]
port 302 nsew signal output
rlabel metal3 s 139200 399848 140000 399968 6 axi_spi_master_w_data[5]
port 303 nsew signal output
rlabel metal3 s 0 287648 800 287768 6 axi_spi_master_w_data[60]
port 304 nsew signal output
rlabel metal2 s 68282 439200 68338 440000 6 axi_spi_master_w_data[61]
port 305 nsew signal output
rlabel metal3 s 0 167968 800 168088 6 axi_spi_master_w_data[62]
port 306 nsew signal output
rlabel metal3 s 139200 112208 140000 112328 6 axi_spi_master_w_data[63]
port 307 nsew signal output
rlabel metal3 s 139200 156408 140000 156528 6 axi_spi_master_w_data[6]
port 308 nsew signal output
rlabel metal3 s 0 34008 800 34128 6 axi_spi_master_w_data[7]
port 309 nsew signal output
rlabel metal3 s 0 274048 800 274168 6 axi_spi_master_w_data[8]
port 310 nsew signal output
rlabel metal2 s 98550 439200 98606 440000 6 axi_spi_master_w_data[9]
port 311 nsew signal output
rlabel metal3 s 0 143488 800 143608 6 axi_spi_master_w_last
port 312 nsew signal output
rlabel metal3 s 0 412088 800 412208 6 axi_spi_master_w_ready
port 313 nsew signal input
rlabel metal2 s 130750 0 130806 800 6 axi_spi_master_w_strb[0]
port 314 nsew signal output
rlabel metal3 s 0 242768 800 242888 6 axi_spi_master_w_strb[1]
port 315 nsew signal output
rlabel metal3 s 139200 36728 140000 36848 6 axi_spi_master_w_strb[2]
port 316 nsew signal output
rlabel metal3 s 139200 82968 140000 83088 6 axi_spi_master_w_strb[3]
port 317 nsew signal output
rlabel metal2 s 21270 0 21326 800 6 axi_spi_master_w_strb[4]
port 318 nsew signal output
rlabel metal3 s 0 158448 800 158568 6 axi_spi_master_w_strb[5]
port 319 nsew signal output
rlabel metal2 s 135258 0 135314 800 6 axi_spi_master_w_strb[6]
port 320 nsew signal output
rlabel metal3 s 0 415488 800 415608 6 axi_spi_master_w_strb[7]
port 321 nsew signal output
rlabel metal3 s 139200 16328 140000 16448 6 axi_spi_master_w_user[0]
port 322 nsew signal output
rlabel metal3 s 139200 5448 140000 5568 6 axi_spi_master_w_user[1]
port 323 nsew signal output
rlabel metal2 s 116582 439200 116638 440000 6 axi_spi_master_w_user[2]
port 324 nsew signal output
rlabel metal2 s 86314 0 86370 800 6 axi_spi_master_w_user[3]
port 325 nsew signal output
rlabel metal3 s 0 367888 800 368008 6 axi_spi_master_w_user[4]
port 326 nsew signal output
rlabel metal3 s 0 73448 800 73568 6 axi_spi_master_w_user[5]
port 327 nsew signal output
rlabel metal3 s 0 250928 800 251048 6 axi_spi_master_w_valid
port 328 nsew signal output
rlabel metal3 s 0 378768 800 378888 6 boot_addr_o[0]
port 329 nsew signal output
rlabel metal3 s 0 429088 800 429208 6 boot_addr_o[10]
port 330 nsew signal output
rlabel metal2 s 53470 0 53526 800 6 boot_addr_o[11]
port 331 nsew signal output
rlabel metal3 s 139200 290368 140000 290488 6 boot_addr_o[12]
port 332 nsew signal output
rlabel metal3 s 0 130568 800 130688 6 boot_addr_o[13]
port 333 nsew signal output
rlabel metal3 s 139200 23808 140000 23928 6 boot_addr_o[14]
port 334 nsew signal output
rlabel metal3 s 139200 19048 140000 19168 6 boot_addr_o[15]
port 335 nsew signal output
rlabel metal3 s 0 82288 800 82408 6 boot_addr_o[16]
port 336 nsew signal output
rlabel metal3 s 0 409368 800 409488 6 boot_addr_o[17]
port 337 nsew signal output
rlabel metal3 s 0 214208 800 214328 6 boot_addr_o[18]
port 338 nsew signal output
rlabel metal3 s 0 332528 800 332648 6 boot_addr_o[19]
port 339 nsew signal output
rlabel metal3 s 139200 348848 140000 348968 6 boot_addr_o[1]
port 340 nsew signal output
rlabel metal3 s 0 311448 800 311568 6 boot_addr_o[20]
port 341 nsew signal output
rlabel metal3 s 0 187008 800 187128 6 boot_addr_o[21]
port 342 nsew signal output
rlabel metal3 s 139200 218968 140000 219088 6 boot_addr_o[22]
port 343 nsew signal output
rlabel metal2 s 1950 439200 2006 440000 6 boot_addr_o[23]
port 344 nsew signal output
rlabel metal3 s 139200 95888 140000 96008 6 boot_addr_o[24]
port 345 nsew signal output
rlabel metal3 s 139200 285608 140000 285728 6 boot_addr_o[25]
port 346 nsew signal output
rlabel metal3 s 139200 8168 140000 8288 6 boot_addr_o[26]
port 347 nsew signal output
rlabel metal3 s 139200 123768 140000 123888 6 boot_addr_o[27]
port 348 nsew signal output
rlabel metal3 s 139200 401888 140000 402008 6 boot_addr_o[28]
port 349 nsew signal output
rlabel metal3 s 0 401888 800 402008 6 boot_addr_o[29]
port 350 nsew signal output
rlabel metal3 s 139200 93848 140000 93968 6 boot_addr_o[2]
port 351 nsew signal output
rlabel metal2 s 82450 0 82506 800 6 boot_addr_o[30]
port 352 nsew signal output
rlabel metal2 s 139766 0 139822 800 6 boot_addr_o[31]
port 353 nsew signal output
rlabel metal3 s 0 421608 800 421728 6 boot_addr_o[3]
port 354 nsew signal output
rlabel metal3 s 0 201288 800 201408 6 boot_addr_o[4]
port 355 nsew signal output
rlabel metal2 s 27710 439200 27766 440000 6 boot_addr_o[5]
port 356 nsew signal output
rlabel metal3 s 0 351568 800 351688 6 boot_addr_o[6]
port 357 nsew signal output
rlabel metal2 s 135902 0 135958 800 6 boot_addr_o[7]
port 358 nsew signal output
rlabel metal3 s 0 81608 800 81728 6 boot_addr_o[8]
port 359 nsew signal output
rlabel metal3 s 0 116968 800 117088 6 boot_addr_o[9]
port 360 nsew signal output
rlabel metal2 s 30286 0 30342 800 6 clk_gate_core_o
port 361 nsew signal output
rlabel metal2 s 74078 0 74134 800 6 clk_i
port 362 nsew signal input
rlabel metal3 s 139200 230528 140000 230648 6 clk_i_pll
port 363 nsew signal input
rlabel metal2 s 12898 0 12954 800 6 clk_o_pll
port 364 nsew signal output
rlabel metal3 s 0 281528 800 281648 6 clk_sel_i_pll
port 365 nsew signal input
rlabel metal3 s 139200 75488 140000 75608 6 clk_standalone_i_pll
port 366 nsew signal input
rlabel metal3 s 0 46928 800 47048 6 core_busy_i
port 367 nsew signal input
rlabel metal2 s 104990 439200 105046 440000 6 debug_addr[0]
port 368 nsew signal output
rlabel metal2 s 47674 439200 47730 440000 6 debug_addr[10]
port 369 nsew signal output
rlabel metal3 s 0 427728 800 427848 6 debug_addr[11]
port 370 nsew signal output
rlabel metal3 s 0 316888 800 317008 6 debug_addr[12]
port 371 nsew signal output
rlabel metal2 s 77942 0 77998 800 6 debug_addr[13]
port 372 nsew signal output
rlabel metal2 s 79874 439200 79930 440000 6 debug_addr[14]
port 373 nsew signal output
rlabel metal3 s 0 372648 800 372768 6 debug_addr[1]
port 374 nsew signal output
rlabel metal2 s 51538 439200 51594 440000 6 debug_addr[2]
port 375 nsew signal output
rlabel metal2 s 58622 0 58678 800 6 debug_addr[3]
port 376 nsew signal output
rlabel metal3 s 0 327768 800 327888 6 debug_addr[4]
port 377 nsew signal output
rlabel metal2 s 94686 439200 94742 440000 6 debug_addr[5]
port 378 nsew signal output
rlabel metal3 s 0 346808 800 346928 6 debug_addr[6]
port 379 nsew signal output
rlabel metal2 s 109498 0 109554 800 6 debug_addr[7]
port 380 nsew signal output
rlabel metal3 s 0 153688 800 153808 6 debug_addr[8]
port 381 nsew signal output
rlabel metal2 s 21914 439200 21970 440000 6 debug_addr[9]
port 382 nsew signal output
rlabel metal3 s 0 90448 800 90568 6 debug_gnt
port 383 nsew signal input
rlabel metal3 s 139200 76168 140000 76288 6 debug_rdata[0]
port 384 nsew signal input
rlabel metal3 s 0 315528 800 315648 6 debug_rdata[10]
port 385 nsew signal input
rlabel metal3 s 0 211488 800 211608 6 debug_rdata[11]
port 386 nsew signal input
rlabel metal3 s 139200 24488 140000 24608 6 debug_rdata[12]
port 387 nsew signal input
rlabel metal3 s 139200 138048 140000 138168 6 debug_rdata[13]
port 388 nsew signal input
rlabel metal3 s 139200 295808 140000 295928 6 debug_rdata[14]
port 389 nsew signal input
rlabel metal3 s 0 244128 800 244248 6 debug_rdata[15]
port 390 nsew signal input
rlabel metal3 s 139200 167288 140000 167408 6 debug_rdata[16]
port 391 nsew signal input
rlabel metal3 s 139200 274728 140000 274848 6 debug_rdata[17]
port 392 nsew signal input
rlabel metal3 s 139200 109488 140000 109608 6 debug_rdata[18]
port 393 nsew signal input
rlabel metal3 s 139200 71408 140000 71528 6 debug_rdata[19]
port 394 nsew signal input
rlabel metal3 s 0 376728 800 376848 6 debug_rdata[1]
port 395 nsew signal input
rlabel metal3 s 0 17008 800 17128 6 debug_rdata[20]
port 396 nsew signal input
rlabel metal3 s 0 2048 800 2168 6 debug_rdata[21]
port 397 nsew signal input
rlabel metal3 s 0 100648 800 100768 6 debug_rdata[22]
port 398 nsew signal input
rlabel metal3 s 0 23808 800 23928 6 debug_rdata[23]
port 399 nsew signal input
rlabel metal2 s 40590 0 40646 800 6 debug_rdata[24]
port 400 nsew signal input
rlabel metal3 s 0 308728 800 308848 6 debug_rdata[25]
port 401 nsew signal input
rlabel metal3 s 0 388968 800 389088 6 debug_rdata[26]
port 402 nsew signal input
rlabel metal3 s 139200 3408 140000 3528 6 debug_rdata[27]
port 403 nsew signal input
rlabel metal2 s 18694 0 18750 800 6 debug_rdata[28]
port 404 nsew signal input
rlabel metal3 s 139200 189728 140000 189848 6 debug_rdata[29]
port 405 nsew signal input
rlabel metal3 s 139200 38768 140000 38888 6 debug_rdata[2]
port 406 nsew signal input
rlabel metal2 s 38014 439200 38070 440000 6 debug_rdata[30]
port 407 nsew signal input
rlabel metal3 s 0 145528 800 145648 6 debug_rdata[31]
port 408 nsew signal input
rlabel metal3 s 139200 439288 140000 439408 6 debug_rdata[3]
port 409 nsew signal input
rlabel metal2 s 123022 0 123078 800 6 debug_rdata[4]
port 410 nsew signal input
rlabel metal2 s 119158 0 119214 800 6 debug_rdata[5]
port 411 nsew signal input
rlabel metal3 s 0 422288 800 422408 6 debug_rdata[6]
port 412 nsew signal input
rlabel metal3 s 139200 49648 140000 49768 6 debug_rdata[7]
port 413 nsew signal input
rlabel metal3 s 0 267928 800 268048 6 debug_rdata[8]
port 414 nsew signal input
rlabel metal3 s 0 260448 800 260568 6 debug_rdata[9]
port 415 nsew signal input
rlabel metal3 s 139200 306688 140000 306808 6 debug_req
port 416 nsew signal output
rlabel metal3 s 139200 335928 140000 336048 6 debug_rvalid
port 417 nsew signal input
rlabel metal3 s 139200 13608 140000 13728 6 debug_wdata[0]
port 418 nsew signal output
rlabel metal3 s 139200 125808 140000 125928 6 debug_wdata[10]
port 419 nsew signal output
rlabel metal3 s 139200 359728 140000 359848 6 debug_wdata[11]
port 420 nsew signal output
rlabel metal2 s 121090 0 121146 800 6 debug_wdata[12]
port 421 nsew signal output
rlabel metal3 s 0 70048 800 70168 6 debug_wdata[13]
port 422 nsew signal output
rlabel metal3 s 0 408688 800 408808 6 debug_wdata[14]
port 423 nsew signal output
rlabel metal3 s 0 301928 800 302048 6 debug_wdata[15]
port 424 nsew signal output
rlabel metal2 s 129462 439200 129518 440000 6 debug_wdata[16]
port 425 nsew signal output
rlabel metal3 s 139200 40808 140000 40928 6 debug_wdata[17]
port 426 nsew signal output
rlabel metal3 s 139200 150288 140000 150408 6 debug_wdata[18]
port 427 nsew signal output
rlabel metal3 s 139200 155048 140000 155168 6 debug_wdata[19]
port 428 nsew signal output
rlabel metal3 s 0 215568 800 215688 6 debug_wdata[1]
port 429 nsew signal output
rlabel metal3 s 0 329808 800 329928 6 debug_wdata[20]
port 430 nsew signal output
rlabel metal3 s 139200 226448 140000 226568 6 debug_wdata[21]
port 431 nsew signal output
rlabel metal3 s 0 43528 800 43648 6 debug_wdata[22]
port 432 nsew signal output
rlabel metal2 s 54114 439200 54170 440000 6 debug_wdata[23]
port 433 nsew signal output
rlabel metal3 s 139200 365848 140000 365968 6 debug_wdata[24]
port 434 nsew signal output
rlabel metal3 s 0 340008 800 340128 6 debug_wdata[25]
port 435 nsew signal output
rlabel metal3 s 139200 414128 140000 414248 6 debug_wdata[26]
port 436 nsew signal output
rlabel metal3 s 0 104728 800 104848 6 debug_wdata[27]
port 437 nsew signal output
rlabel metal3 s 0 310088 800 310208 6 debug_wdata[28]
port 438 nsew signal output
rlabel metal2 s 58622 439200 58678 440000 6 debug_wdata[29]
port 439 nsew signal output
rlabel metal3 s 0 96568 800 96688 6 debug_wdata[2]
port 440 nsew signal output
rlabel metal3 s 139200 176128 140000 176248 6 debug_wdata[30]
port 441 nsew signal output
rlabel metal2 s 44454 0 44510 800 6 debug_wdata[31]
port 442 nsew signal output
rlabel metal2 s 95330 439200 95386 440000 6 debug_wdata[3]
port 443 nsew signal output
rlabel metal3 s 0 66648 800 66768 6 debug_wdata[4]
port 444 nsew signal output
rlabel metal3 s 0 201968 800 202088 6 debug_wdata[5]
port 445 nsew signal output
rlabel metal3 s 0 150968 800 151088 6 debug_wdata[6]
port 446 nsew signal output
rlabel metal3 s 0 274728 800 274848 6 debug_wdata[7]
port 447 nsew signal output
rlabel metal3 s 139200 688 140000 808 6 debug_wdata[8]
port 448 nsew signal output
rlabel metal2 s 105634 0 105690 800 6 debug_wdata[9]
port 449 nsew signal output
rlabel metal2 s 90822 439200 90878 440000 6 debug_we
port 450 nsew signal output
rlabel metal3 s 139200 46248 140000 46368 6 fetch_enable_i
port 451 nsew signal input
rlabel metal3 s 0 395768 800 395888 6 fetch_enable_o
port 452 nsew signal output
rlabel metal3 s 139200 107448 140000 107568 6 fll1_ack_i
port 453 nsew signal input
rlabel metal3 s 0 14288 800 14408 6 fll1_add_o[0]
port 454 nsew signal output
rlabel metal3 s 139200 214208 140000 214328 6 fll1_add_o[1]
port 455 nsew signal output
rlabel metal3 s 0 20408 800 20528 6 fll1_lock_i
port 456 nsew signal input
rlabel metal3 s 139200 211488 140000 211608 6 fll1_rdata_i[0]
port 457 nsew signal input
rlabel metal2 s 44454 439200 44510 440000 6 fll1_rdata_i[10]
port 458 nsew signal input
rlabel metal2 s 26422 0 26478 800 6 fll1_rdata_i[11]
port 459 nsew signal input
rlabel metal3 s 0 133968 800 134088 6 fll1_rdata_i[12]
port 460 nsew signal input
rlabel metal3 s 0 124448 800 124568 6 fll1_rdata_i[13]
port 461 nsew signal input
rlabel metal3 s 0 333888 800 334008 6 fll1_rdata_i[14]
port 462 nsew signal input
rlabel metal3 s 0 190408 800 190528 6 fll1_rdata_i[15]
port 463 nsew signal input
rlabel metal3 s 139200 292408 140000 292528 6 fll1_rdata_i[16]
port 464 nsew signal input
rlabel metal3 s 0 276088 800 276208 6 fll1_rdata_i[17]
port 465 nsew signal input
rlabel metal2 s 14830 439200 14886 440000 6 fll1_rdata_i[18]
port 466 nsew signal input
rlabel metal2 s 66350 0 66406 800 6 fll1_rdata_i[19]
port 467 nsew signal input
rlabel metal2 s 60554 0 60610 800 6 fll1_rdata_i[1]
port 468 nsew signal input
rlabel metal3 s 0 425008 800 425128 6 fll1_rdata_i[20]
port 469 nsew signal input
rlabel metal3 s 139200 402568 140000 402688 6 fll1_rdata_i[21]
port 470 nsew signal input
rlabel metal3 s 139200 87728 140000 87848 6 fll1_rdata_i[22]
port 471 nsew signal input
rlabel metal3 s 139200 421608 140000 421728 6 fll1_rdata_i[23]
port 472 nsew signal input
rlabel metal3 s 139200 25168 140000 25288 6 fll1_rdata_i[24]
port 473 nsew signal input
rlabel metal3 s 139200 2728 140000 2848 6 fll1_rdata_i[25]
port 474 nsew signal input
rlabel metal2 s 26422 439200 26478 440000 6 fll1_rdata_i[26]
port 475 nsew signal input
rlabel metal3 s 139200 425688 140000 425808 6 fll1_rdata_i[27]
port 476 nsew signal input
rlabel metal2 s 113362 439200 113418 440000 6 fll1_rdata_i[28]
port 477 nsew signal input
rlabel metal2 s 47030 439200 47086 440000 6 fll1_rdata_i[29]
port 478 nsew signal input
rlabel metal3 s 0 60528 800 60648 6 fll1_rdata_i[2]
port 479 nsew signal input
rlabel metal3 s 139200 206728 140000 206848 6 fll1_rdata_i[30]
port 480 nsew signal input
rlabel metal3 s 139200 275408 140000 275528 6 fll1_rdata_i[31]
port 481 nsew signal input
rlabel metal3 s 0 325048 800 325168 6 fll1_rdata_i[3]
port 482 nsew signal input
rlabel metal3 s 139200 203328 140000 203448 6 fll1_rdata_i[4]
port 483 nsew signal input
rlabel metal3 s 0 137368 800 137488 6 fll1_rdata_i[5]
port 484 nsew signal input
rlabel metal3 s 139200 432488 140000 432608 6 fll1_rdata_i[6]
port 485 nsew signal input
rlabel metal3 s 139200 125128 140000 125248 6 fll1_rdata_i[7]
port 486 nsew signal input
rlabel metal3 s 139200 98608 140000 98728 6 fll1_rdata_i[8]
port 487 nsew signal input
rlabel metal3 s 0 221008 800 221128 6 fll1_rdata_i[9]
port 488 nsew signal input
rlabel metal3 s 139200 31288 140000 31408 6 fll1_req_o
port 489 nsew signal output
rlabel metal3 s 0 9528 800 9648 6 fll1_wdata_o[0]
port 490 nsew signal output
rlabel metal3 s 139200 127848 140000 127968 6 fll1_wdata_o[10]
port 491 nsew signal output
rlabel metal3 s 0 282888 800 283008 6 fll1_wdata_o[11]
port 492 nsew signal output
rlabel metal3 s 139200 102688 140000 102808 6 fll1_wdata_o[12]
port 493 nsew signal output
rlabel metal2 s 62486 0 62542 800 6 fll1_wdata_o[13]
port 494 nsew signal output
rlabel metal3 s 0 219648 800 219768 6 fll1_wdata_o[14]
port 495 nsew signal output
rlabel metal2 s 87602 439200 87658 440000 6 fll1_wdata_o[15]
port 496 nsew signal output
rlabel metal3 s 139200 410048 140000 410168 6 fll1_wdata_o[16]
port 497 nsew signal output
rlabel metal3 s 139200 131248 140000 131368 6 fll1_wdata_o[17]
port 498 nsew signal output
rlabel metal3 s 0 122408 800 122528 6 fll1_wdata_o[18]
port 499 nsew signal output
rlabel metal2 s 96618 0 96674 800 6 fll1_wdata_o[19]
port 500 nsew signal output
rlabel metal2 s 112074 439200 112130 440000 6 fll1_wdata_o[1]
port 501 nsew signal output
rlabel metal2 s 119802 439200 119858 440000 6 fll1_wdata_o[20]
port 502 nsew signal output
rlabel metal3 s 139200 255688 140000 255808 6 fll1_wdata_o[21]
port 503 nsew signal output
rlabel metal3 s 139200 228488 140000 228608 6 fll1_wdata_o[22]
port 504 nsew signal output
rlabel metal3 s 0 194488 800 194608 6 fll1_wdata_o[23]
port 505 nsew signal output
rlabel metal3 s 0 324368 800 324488 6 fll1_wdata_o[24]
port 506 nsew signal output
rlabel metal3 s 139200 216248 140000 216368 6 fll1_wdata_o[25]
port 507 nsew signal output
rlabel metal2 s 124954 0 125010 800 6 fll1_wdata_o[26]
port 508 nsew signal output
rlabel metal2 s 39946 439200 40002 440000 6 fll1_wdata_o[27]
port 509 nsew signal output
rlabel metal3 s 0 354288 800 354408 6 fll1_wdata_o[28]
port 510 nsew signal output
rlabel metal3 s 139200 293768 140000 293888 6 fll1_wdata_o[29]
port 511 nsew signal output
rlabel metal3 s 139200 256368 140000 256488 6 fll1_wdata_o[2]
port 512 nsew signal output
rlabel metal3 s 139200 288328 140000 288448 6 fll1_wdata_o[30]
port 513 nsew signal output
rlabel metal3 s 0 31288 800 31408 6 fll1_wdata_o[31]
port 514 nsew signal output
rlabel metal3 s 139200 252968 140000 253088 6 fll1_wdata_o[3]
port 515 nsew signal output
rlabel metal3 s 0 330488 800 330608 6 fll1_wdata_o[4]
port 516 nsew signal output
rlabel metal2 s 87602 0 87658 800 6 fll1_wdata_o[5]
port 517 nsew signal output
rlabel metal3 s 0 427048 800 427168 6 fll1_wdata_o[6]
port 518 nsew signal output
rlabel metal3 s 0 44888 800 45008 6 fll1_wdata_o[7]
port 519 nsew signal output
rlabel metal2 s 32862 0 32918 800 6 fll1_wdata_o[8]
port 520 nsew signal output
rlabel metal3 s 0 105408 800 105528 6 fll1_wdata_o[9]
port 521 nsew signal output
rlabel metal3 s 0 362448 800 362568 6 fll1_wrn_o
port 522 nsew signal output
rlabel metal3 s 0 249568 800 249688 6 fll_ack_o_pll
port 523 nsew signal output
rlabel metal3 s 0 303968 800 304088 6 fll_add_i_pll[0]
port 524 nsew signal input
rlabel metal3 s 139200 260448 140000 260568 6 fll_add_i_pll[1]
port 525 nsew signal input
rlabel metal2 s 94686 0 94742 800 6 fll_data_i_pll[0]
port 526 nsew signal input
rlabel metal3 s 139200 286288 140000 286408 6 fll_data_i_pll[10]
port 527 nsew signal input
rlabel metal3 s 0 51688 800 51808 6 fll_data_i_pll[11]
port 528 nsew signal input
rlabel metal3 s 139200 279488 140000 279608 6 fll_data_i_pll[12]
port 529 nsew signal input
rlabel metal3 s 139200 356328 140000 356448 6 fll_data_i_pll[13]
port 530 nsew signal input
rlabel metal3 s 139200 434528 140000 434648 6 fll_data_i_pll[14]
port 531 nsew signal input
rlabel metal3 s 0 236648 800 236768 6 fll_data_i_pll[15]
port 532 nsew signal input
rlabel metal2 s 47030 0 47086 800 6 fll_data_i_pll[16]
port 533 nsew signal input
rlabel metal3 s 139200 182248 140000 182368 6 fll_data_i_pll[17]
port 534 nsew signal input
rlabel metal3 s 0 318928 800 319048 6 fll_data_i_pll[18]
port 535 nsew signal input
rlabel metal3 s 139200 172728 140000 172848 6 fll_data_i_pll[19]
port 536 nsew signal input
rlabel metal2 s 22558 0 22614 800 6 fll_data_i_pll[1]
port 537 nsew signal input
rlabel metal3 s 139200 296488 140000 296608 6 fll_data_i_pll[20]
port 538 nsew signal input
rlabel metal3 s 0 161848 800 161968 6 fll_data_i_pll[21]
port 539 nsew signal input
rlabel metal2 s 28998 439200 29054 440000 6 fll_data_i_pll[22]
port 540 nsew signal input
rlabel metal3 s 0 375368 800 375488 6 fll_data_i_pll[23]
port 541 nsew signal input
rlabel metal2 s 104990 0 105046 800 6 fll_data_i_pll[24]
port 542 nsew signal input
rlabel metal3 s 139200 67328 140000 67448 6 fll_data_i_pll[25]
port 543 nsew signal input
rlabel metal3 s 139200 42168 140000 42288 6 fll_data_i_pll[26]
port 544 nsew signal input
rlabel metal3 s 0 94528 800 94648 6 fll_data_i_pll[27]
port 545 nsew signal input
rlabel metal3 s 0 346128 800 346248 6 fll_data_i_pll[28]
port 546 nsew signal input
rlabel metal3 s 139200 252288 140000 252408 6 fll_data_i_pll[29]
port 547 nsew signal input
rlabel metal3 s 0 217608 800 217728 6 fll_data_i_pll[2]
port 548 nsew signal input
rlabel metal3 s 139200 39448 140000 39568 6 fll_data_i_pll[30]
port 549 nsew signal input
rlabel metal3 s 0 333208 800 333328 6 fll_data_i_pll[31]
port 550 nsew signal input
rlabel metal3 s 139200 99968 140000 100088 6 fll_data_i_pll[3]
port 551 nsew signal input
rlabel metal2 s 61198 439200 61254 440000 6 fll_data_i_pll[4]
port 552 nsew signal input
rlabel metal3 s 139200 198568 140000 198688 6 fll_data_i_pll[5]
port 553 nsew signal input
rlabel metal3 s 0 78888 800 79008 6 fll_data_i_pll[6]
port 554 nsew signal input
rlabel metal3 s 0 336608 800 336728 6 fll_data_i_pll[7]
port 555 nsew signal input
rlabel metal3 s 0 193808 800 193928 6 fll_data_i_pll[8]
port 556 nsew signal input
rlabel metal3 s 139200 333888 140000 334008 6 fll_data_i_pll[9]
port 557 nsew signal input
rlabel metal3 s 139200 413448 140000 413568 6 fll_lock_o_pll
port 558 nsew signal output
rlabel metal3 s 139200 192448 140000 192568 6 fll_r_data_o_pll[0]
port 559 nsew signal output
rlabel metal3 s 0 269968 800 270088 6 fll_r_data_o_pll[10]
port 560 nsew signal output
rlabel metal3 s 139200 299208 140000 299328 6 fll_r_data_o_pll[11]
port 561 nsew signal output
rlabel metal3 s 139200 264528 140000 264648 6 fll_r_data_o_pll[12]
port 562 nsew signal output
rlabel metal2 s 40590 439200 40646 440000 6 fll_r_data_o_pll[13]
port 563 nsew signal output
rlabel metal3 s 139200 313488 140000 313608 6 fll_r_data_o_pll[14]
port 564 nsew signal output
rlabel metal2 s 125598 439200 125654 440000 6 fll_r_data_o_pll[15]
port 565 nsew signal output
rlabel metal3 s 0 374688 800 374808 6 fll_r_data_o_pll[16]
port 566 nsew signal output
rlabel metal3 s 139200 21768 140000 21888 6 fll_r_data_o_pll[17]
port 567 nsew signal output
rlabel metal3 s 0 188368 800 188488 6 fll_r_data_o_pll[18]
port 568 nsew signal output
rlabel metal3 s 139200 23128 140000 23248 6 fll_r_data_o_pll[19]
port 569 nsew signal output
rlabel metal3 s 139200 406648 140000 406768 6 fll_r_data_o_pll[1]
port 570 nsew signal output
rlabel metal3 s 139200 307368 140000 307488 6 fll_r_data_o_pll[20]
port 571 nsew signal output
rlabel metal3 s 0 131928 800 132048 6 fll_r_data_o_pll[21]
port 572 nsew signal output
rlabel metal2 s 36726 0 36782 800 6 fll_r_data_o_pll[22]
port 573 nsew signal output
rlabel metal3 s 0 337968 800 338088 6 fll_r_data_o_pll[23]
port 574 nsew signal output
rlabel metal2 s 34794 0 34850 800 6 fll_r_data_o_pll[24]
port 575 nsew signal output
rlabel metal3 s 0 78208 800 78328 6 fll_r_data_o_pll[25]
port 576 nsew signal output
rlabel metal3 s 0 365848 800 365968 6 fll_r_data_o_pll[26]
port 577 nsew signal output
rlabel metal3 s 0 37408 800 37528 6 fll_r_data_o_pll[27]
port 578 nsew signal output
rlabel metal3 s 0 239368 800 239488 6 fll_r_data_o_pll[28]
port 579 nsew signal output
rlabel metal3 s 0 345448 800 345568 6 fll_r_data_o_pll[29]
port 580 nsew signal output
rlabel metal3 s 0 153008 800 153128 6 fll_r_data_o_pll[2]
port 581 nsew signal output
rlabel metal3 s 0 185648 800 185768 6 fll_r_data_o_pll[30]
port 582 nsew signal output
rlabel metal3 s 139200 181568 140000 181688 6 fll_r_data_o_pll[31]
port 583 nsew signal output
rlabel metal2 s 99194 439200 99250 440000 6 fll_r_data_o_pll[3]
port 584 nsew signal output
rlabel metal3 s 0 27208 800 27328 6 fll_r_data_o_pll[4]
port 585 nsew signal output
rlabel metal3 s 139200 394408 140000 394528 6 fll_r_data_o_pll[5]
port 586 nsew signal output
rlabel metal3 s 0 1368 800 1488 6 fll_r_data_o_pll[6]
port 587 nsew signal output
rlabel metal3 s 0 172048 800 172168 6 fll_r_data_o_pll[7]
port 588 nsew signal output
rlabel metal3 s 0 106768 800 106888 6 fll_r_data_o_pll[8]
port 589 nsew signal output
rlabel metal3 s 139200 382848 140000 382968 6 fll_r_data_o_pll[9]
port 590 nsew signal output
rlabel metal2 s 24490 439200 24546 440000 6 fll_req_i_pll
port 591 nsew signal input
rlabel metal3 s 139200 180888 140000 181008 6 fll_wrn_i_pll
port 592 nsew signal input
rlabel metal2 s 64418 0 64474 800 6 gpio_dir[0]
port 593 nsew signal output
rlabel metal3 s 139200 371288 140000 371408 6 gpio_dir[10]
port 594 nsew signal output
rlabel metal3 s 0 247528 800 247648 6 gpio_dir[11]
port 595 nsew signal output
rlabel metal3 s 0 255688 800 255808 6 gpio_dir[12]
port 596 nsew signal output
rlabel metal3 s 139200 20408 140000 20528 6 gpio_dir[13]
port 597 nsew signal output
rlabel metal3 s 139200 115608 140000 115728 6 gpio_dir[14]
port 598 nsew signal output
rlabel metal3 s 139200 281528 140000 281648 6 gpio_dir[15]
port 599 nsew signal output
rlabel metal3 s 139200 209448 140000 209568 6 gpio_dir[16]
port 600 nsew signal output
rlabel metal3 s 0 2728 800 2848 6 gpio_dir[17]
port 601 nsew signal output
rlabel metal2 s 30930 439200 30986 440000 6 gpio_dir[18]
port 602 nsew signal output
rlabel metal3 s 0 233928 800 234048 6 gpio_dir[19]
port 603 nsew signal output
rlabel metal3 s 139200 337968 140000 338088 6 gpio_dir[1]
port 604 nsew signal output
rlabel metal3 s 139200 368568 140000 368688 6 gpio_dir[20]
port 605 nsew signal output
rlabel metal2 s 139766 439200 139822 440000 6 gpio_dir[21]
port 606 nsew signal output
rlabel metal3 s 0 49648 800 49768 6 gpio_dir[22]
port 607 nsew signal output
rlabel metal2 s 6458 439200 6514 440000 6 gpio_dir[23]
port 608 nsew signal output
rlabel metal2 s 41878 0 41934 800 6 gpio_dir[24]
port 609 nsew signal output
rlabel metal2 s 52826 0 52882 800 6 gpio_dir[25]
port 610 nsew signal output
rlabel metal3 s 0 76848 800 76968 6 gpio_dir[26]
port 611 nsew signal output
rlabel metal3 s 139200 238688 140000 238808 6 gpio_dir[27]
port 612 nsew signal output
rlabel metal3 s 0 193128 800 193248 6 gpio_dir[28]
port 613 nsew signal output
rlabel metal3 s 139200 320968 140000 321088 6 gpio_dir[29]
port 614 nsew signal output
rlabel metal2 s 3882 439200 3938 440000 6 gpio_dir[2]
port 615 nsew signal output
rlabel metal2 s 99838 0 99894 800 6 gpio_dir[30]
port 616 nsew signal output
rlabel metal3 s 139200 186328 140000 186448 6 gpio_dir[31]
port 617 nsew signal output
rlabel metal3 s 139200 128528 140000 128648 6 gpio_dir[3]
port 618 nsew signal output
rlabel metal3 s 0 403928 800 404048 6 gpio_dir[4]
port 619 nsew signal output
rlabel metal3 s 0 352928 800 353048 6 gpio_dir[5]
port 620 nsew signal output
rlabel metal3 s 0 350888 800 351008 6 gpio_dir[6]
port 621 nsew signal output
rlabel metal3 s 0 11568 800 11688 6 gpio_dir[7]
port 622 nsew signal output
rlabel metal3 s 0 149608 800 149728 6 gpio_dir[8]
port 623 nsew signal output
rlabel metal3 s 0 155048 800 155168 6 gpio_dir[9]
port 624 nsew signal output
rlabel metal3 s 139200 170688 140000 170808 6 gpio_in[0]
port 625 nsew signal input
rlabel metal3 s 139200 100648 140000 100768 6 gpio_in[10]
port 626 nsew signal input
rlabel metal3 s 0 269288 800 269408 6 gpio_in[11]
port 627 nsew signal input
rlabel metal3 s 0 21768 800 21888 6 gpio_in[12]
port 628 nsew signal input
rlabel metal3 s 0 307368 800 307488 6 gpio_in[13]
port 629 nsew signal input
rlabel metal3 s 0 133288 800 133408 6 gpio_in[14]
port 630 nsew signal input
rlabel metal2 s 14186 439200 14242 440000 6 gpio_in[15]
port 631 nsew signal input
rlabel metal3 s 139200 340688 140000 340808 6 gpio_in[16]
port 632 nsew signal input
rlabel metal3 s 139200 14968 140000 15088 6 gpio_in[17]
port 633 nsew signal input
rlabel metal2 s 79230 439200 79286 440000 6 gpio_in[18]
port 634 nsew signal input
rlabel metal2 s 43166 0 43222 800 6 gpio_in[19]
port 635 nsew signal input
rlabel metal3 s 0 157768 800 157888 6 gpio_in[1]
port 636 nsew signal input
rlabel metal3 s 139200 317568 140000 317688 6 gpio_in[20]
port 637 nsew signal input
rlabel metal3 s 139200 346128 140000 346248 6 gpio_in[21]
port 638 nsew signal input
rlabel metal2 s 4526 0 4582 800 6 gpio_in[22]
port 639 nsew signal input
rlabel metal2 s 115938 439200 115994 440000 6 gpio_in[23]
port 640 nsew signal input
rlabel metal3 s 139200 53048 140000 53168 6 gpio_in[24]
port 641 nsew signal input
rlabel metal3 s 0 47608 800 47728 6 gpio_in[25]
port 642 nsew signal input
rlabel metal3 s 139200 388288 140000 388408 6 gpio_in[26]
port 643 nsew signal input
rlabel metal3 s 139200 6128 140000 6248 6 gpio_in[27]
port 644 nsew signal input
rlabel metal3 s 139200 18368 140000 18488 6 gpio_in[28]
port 645 nsew signal input
rlabel metal2 s 25134 439200 25190 440000 6 gpio_in[29]
port 646 nsew signal input
rlabel metal2 s 77298 439200 77354 440000 6 gpio_in[2]
port 647 nsew signal input
rlabel metal3 s 0 242088 800 242208 6 gpio_in[30]
port 648 nsew signal input
rlabel metal3 s 0 38768 800 38888 6 gpio_in[31]
port 649 nsew signal input
rlabel metal3 s 0 183608 800 183728 6 gpio_in[3]
port 650 nsew signal input
rlabel metal3 s 139200 326408 140000 326528 6 gpio_in[4]
port 651 nsew signal input
rlabel metal3 s 139200 50328 140000 50448 6 gpio_in[5]
port 652 nsew signal input
rlabel metal2 s 50894 0 50950 800 6 gpio_in[6]
port 653 nsew signal input
rlabel metal2 s 118514 0 118570 800 6 gpio_in[7]
port 654 nsew signal input
rlabel metal3 s 139200 251608 140000 251728 6 gpio_in[8]
port 655 nsew signal input
rlabel metal3 s 0 368568 800 368688 6 gpio_in[9]
port 656 nsew signal input
rlabel metal2 s 70858 439200 70914 440000 6 gpio_out[0]
port 657 nsew signal output
rlabel metal3 s 139200 213528 140000 213648 6 gpio_out[10]
port 658 nsew signal output
rlabel metal2 s 90178 439200 90234 440000 6 gpio_out[11]
port 659 nsew signal output
rlabel metal2 s 119802 0 119858 800 6 gpio_out[12]
port 660 nsew signal output
rlabel metal3 s 0 55768 800 55888 6 gpio_out[13]
port 661 nsew signal output
rlabel metal3 s 0 414128 800 414248 6 gpio_out[14]
port 662 nsew signal output
rlabel metal3 s 139200 350888 140000 351008 6 gpio_out[15]
port 663 nsew signal output
rlabel metal3 s 139200 316888 140000 317008 6 gpio_out[16]
port 664 nsew signal output
rlabel metal2 s 57978 439200 58034 440000 6 gpio_out[17]
port 665 nsew signal output
rlabel metal3 s 139200 163888 140000 164008 6 gpio_out[18]
port 666 nsew signal output
rlabel metal3 s 139200 269968 140000 270088 6 gpio_out[19]
port 667 nsew signal output
rlabel metal3 s 0 65288 800 65408 6 gpio_out[1]
port 668 nsew signal output
rlabel metal3 s 0 72768 800 72888 6 gpio_out[20]
port 669 nsew signal output
rlabel metal2 s 65062 0 65118 800 6 gpio_out[21]
port 670 nsew signal output
rlabel metal3 s 0 181568 800 181688 6 gpio_out[22]
port 671 nsew signal output
rlabel metal3 s 139200 248888 140000 249008 6 gpio_out[23]
port 672 nsew signal output
rlabel metal3 s 0 357008 800 357128 6 gpio_out[24]
port 673 nsew signal output
rlabel metal2 s 18694 439200 18750 440000 6 gpio_out[25]
port 674 nsew signal output
rlabel metal3 s 0 688 800 808 6 gpio_out[26]
port 675 nsew signal output
rlabel metal3 s 0 197888 800 198008 6 gpio_out[27]
port 676 nsew signal output
rlabel metal3 s 139200 262488 140000 262608 6 gpio_out[28]
port 677 nsew signal output
rlabel metal3 s 139200 83648 140000 83768 6 gpio_out[29]
port 678 nsew signal output
rlabel metal2 s 91466 0 91522 800 6 gpio_out[2]
port 679 nsew signal output
rlabel metal3 s 0 291728 800 291848 6 gpio_out[30]
port 680 nsew signal output
rlabel metal3 s 0 379448 800 379568 6 gpio_out[31]
port 681 nsew signal output
rlabel metal3 s 0 155728 800 155848 6 gpio_out[3]
port 682 nsew signal output
rlabel metal2 s 100482 439200 100538 440000 6 gpio_out[4]
port 683 nsew signal output
rlabel metal3 s 139200 82288 140000 82408 6 gpio_out[5]
port 684 nsew signal output
rlabel metal3 s 139200 258408 140000 258528 6 gpio_out[6]
port 685 nsew signal output
rlabel metal3 s 0 402568 800 402688 6 gpio_out[7]
port 686 nsew signal output
rlabel metal3 s 0 144848 800 144968 6 gpio_out[8]
port 687 nsew signal output
rlabel metal3 s 139200 372648 140000 372768 6 gpio_out[9]
port 688 nsew signal output
rlabel metal3 s 139200 201968 140000 202088 6 gpio_padcfg[0]
port 689 nsew signal output
rlabel metal3 s 139200 45568 140000 45688 6 gpio_padcfg[100]
port 690 nsew signal output
rlabel metal3 s 139200 240728 140000 240848 6 gpio_padcfg[101]
port 691 nsew signal output
rlabel metal3 s 0 12928 800 13048 6 gpio_padcfg[102]
port 692 nsew signal output
rlabel metal3 s 0 134648 800 134768 6 gpio_padcfg[103]
port 693 nsew signal output
rlabel metal3 s 139200 129888 140000 130008 6 gpio_padcfg[104]
port 694 nsew signal output
rlabel metal2 s 74078 439200 74134 440000 6 gpio_padcfg[105]
port 695 nsew signal output
rlabel metal3 s 0 121728 800 121848 6 gpio_padcfg[106]
port 696 nsew signal output
rlabel metal3 s 0 278808 800 278928 6 gpio_padcfg[107]
port 697 nsew signal output
rlabel metal3 s 139200 422288 140000 422408 6 gpio_padcfg[108]
port 698 nsew signal output
rlabel metal2 s 12254 0 12310 800 6 gpio_padcfg[109]
port 699 nsew signal output
rlabel metal3 s 0 31968 800 32088 6 gpio_padcfg[10]
port 700 nsew signal output
rlabel metal3 s 139200 435208 140000 435328 6 gpio_padcfg[110]
port 701 nsew signal output
rlabel metal2 s 54758 439200 54814 440000 6 gpio_padcfg[111]
port 702 nsew signal output
rlabel metal3 s 139200 32648 140000 32768 6 gpio_padcfg[112]
port 703 nsew signal output
rlabel metal3 s 0 342728 800 342848 6 gpio_padcfg[113]
port 704 nsew signal output
rlabel metal2 s 38014 0 38070 800 6 gpio_padcfg[114]
port 705 nsew signal output
rlabel metal3 s 0 69368 800 69488 6 gpio_padcfg[115]
port 706 nsew signal output
rlabel metal3 s 139200 241408 140000 241528 6 gpio_padcfg[116]
port 707 nsew signal output
rlabel metal3 s 0 286288 800 286408 6 gpio_padcfg[117]
port 708 nsew signal output
rlabel metal2 s 64418 439200 64474 440000 6 gpio_padcfg[118]
port 709 nsew signal output
rlabel metal2 s 20626 0 20682 800 6 gpio_padcfg[119]
port 710 nsew signal output
rlabel metal2 s 9034 0 9090 800 6 gpio_padcfg[11]
port 711 nsew signal output
rlabel metal3 s 0 435888 800 436008 6 gpio_padcfg[120]
port 712 nsew signal output
rlabel metal3 s 0 191768 800 191888 6 gpio_padcfg[121]
port 713 nsew signal output
rlabel metal2 s 117226 0 117282 800 6 gpio_padcfg[122]
port 714 nsew signal output
rlabel metal2 s 37370 0 37426 800 6 gpio_padcfg[123]
port 715 nsew signal output
rlabel metal2 s 12898 439200 12954 440000 6 gpio_padcfg[124]
port 716 nsew signal output
rlabel metal2 s 106922 0 106978 800 6 gpio_padcfg[125]
port 717 nsew signal output
rlabel metal2 s 76654 439200 76710 440000 6 gpio_padcfg[126]
port 718 nsew signal output
rlabel metal3 s 0 433848 800 433968 6 gpio_padcfg[127]
port 719 nsew signal output
rlabel metal2 s 132038 439200 132094 440000 6 gpio_padcfg[128]
port 720 nsew signal output
rlabel metal3 s 139200 412768 140000 412888 6 gpio_padcfg[129]
port 721 nsew signal output
rlabel metal3 s 0 293088 800 293208 6 gpio_padcfg[12]
port 722 nsew signal output
rlabel metal3 s 0 298528 800 298648 6 gpio_padcfg[130]
port 723 nsew signal output
rlabel metal3 s 139200 218288 140000 218408 6 gpio_padcfg[131]
port 724 nsew signal output
rlabel metal3 s 139200 403928 140000 404048 6 gpio_padcfg[132]
port 725 nsew signal output
rlabel metal3 s 139200 333208 140000 333328 6 gpio_padcfg[133]
port 726 nsew signal output
rlabel metal3 s 139200 172048 140000 172168 6 gpio_padcfg[134]
port 727 nsew signal output
rlabel metal2 s 104346 439200 104402 440000 6 gpio_padcfg[135]
port 728 nsew signal output
rlabel metal3 s 0 257728 800 257848 6 gpio_padcfg[136]
port 729 nsew signal output
rlabel metal2 s 70858 0 70914 800 6 gpio_padcfg[137]
port 730 nsew signal output
rlabel metal3 s 139200 231888 140000 232008 6 gpio_padcfg[138]
port 731 nsew signal output
rlabel metal3 s 139200 190408 140000 190528 6 gpio_padcfg[139]
port 732 nsew signal output
rlabel metal3 s 139200 81608 140000 81728 6 gpio_padcfg[13]
port 733 nsew signal output
rlabel metal2 s 110786 439200 110842 440000 6 gpio_padcfg[140]
port 734 nsew signal output
rlabel metal3 s 139200 193128 140000 193248 6 gpio_padcfg[141]
port 735 nsew signal output
rlabel metal3 s 0 295808 800 295928 6 gpio_padcfg[142]
port 736 nsew signal output
rlabel metal3 s 139200 411408 140000 411528 6 gpio_padcfg[143]
port 737 nsew signal output
rlabel metal2 s 112718 439200 112774 440000 6 gpio_padcfg[144]
port 738 nsew signal output
rlabel metal3 s 0 26528 800 26648 6 gpio_padcfg[145]
port 739 nsew signal output
rlabel metal3 s 0 431128 800 431248 6 gpio_padcfg[146]
port 740 nsew signal output
rlabel metal2 s 14186 0 14242 800 6 gpio_padcfg[147]
port 741 nsew signal output
rlabel metal3 s 139200 418208 140000 418328 6 gpio_padcfg[148]
port 742 nsew signal output
rlabel metal3 s 139200 237328 140000 237448 6 gpio_padcfg[149]
port 743 nsew signal output
rlabel metal3 s 0 87048 800 87168 6 gpio_padcfg[14]
port 744 nsew signal output
rlabel metal2 s 39302 0 39358 800 6 gpio_padcfg[150]
port 745 nsew signal output
rlabel metal3 s 0 410728 800 410848 6 gpio_padcfg[151]
port 746 nsew signal output
rlabel metal2 s 92754 0 92810 800 6 gpio_padcfg[152]
port 747 nsew signal output
rlabel metal2 s 19338 439200 19394 440000 6 gpio_padcfg[153]
port 748 nsew signal output
rlabel metal3 s 139200 250248 140000 250368 6 gpio_padcfg[154]
port 749 nsew signal output
rlabel metal3 s 139200 178848 140000 178968 6 gpio_padcfg[155]
port 750 nsew signal output
rlabel metal3 s 0 7488 800 7608 6 gpio_padcfg[156]
port 751 nsew signal output
rlabel metal3 s 139200 155728 140000 155848 6 gpio_padcfg[157]
port 752 nsew signal output
rlabel metal3 s 139200 157768 140000 157888 6 gpio_padcfg[158]
port 753 nsew signal output
rlabel metal3 s 139200 420928 140000 421048 6 gpio_padcfg[159]
port 754 nsew signal output
rlabel metal3 s 139200 233248 140000 233368 6 gpio_padcfg[15]
port 755 nsew signal output
rlabel metal2 s 662 439200 718 440000 6 gpio_padcfg[160]
port 756 nsew signal output
rlabel metal3 s 0 146888 800 147008 6 gpio_padcfg[161]
port 757 nsew signal output
rlabel metal3 s 139200 10888 140000 11008 6 gpio_padcfg[162]
port 758 nsew signal output
rlabel metal2 s 55402 439200 55458 440000 6 gpio_padcfg[163]
port 759 nsew signal output
rlabel metal3 s 139200 396448 140000 396568 6 gpio_padcfg[164]
port 760 nsew signal output
rlabel metal3 s 139200 242768 140000 242888 6 gpio_padcfg[165]
port 761 nsew signal output
rlabel metal3 s 139200 436568 140000 436688 6 gpio_padcfg[166]
port 762 nsew signal output
rlabel metal3 s 139200 231208 140000 231328 6 gpio_padcfg[167]
port 763 nsew signal output
rlabel metal2 s 95974 439200 96030 440000 6 gpio_padcfg[168]
port 764 nsew signal output
rlabel metal3 s 139200 97248 140000 97368 6 gpio_padcfg[169]
port 765 nsew signal output
rlabel metal3 s 0 210808 800 210928 6 gpio_padcfg[16]
port 766 nsew signal output
rlabel metal3 s 0 350208 800 350328 6 gpio_padcfg[170]
port 767 nsew signal output
rlabel metal3 s 139200 139408 140000 139528 6 gpio_padcfg[171]
port 768 nsew signal output
rlabel metal2 s 101770 0 101826 800 6 gpio_padcfg[172]
port 769 nsew signal output
rlabel metal3 s 0 363128 800 363248 6 gpio_padcfg[173]
port 770 nsew signal output
rlabel metal2 s 59266 439200 59322 440000 6 gpio_padcfg[174]
port 771 nsew signal output
rlabel metal3 s 139200 354968 140000 355088 6 gpio_padcfg[175]
port 772 nsew signal output
rlabel metal3 s 139200 159128 140000 159248 6 gpio_padcfg[176]
port 773 nsew signal output
rlabel metal3 s 139200 329128 140000 329248 6 gpio_padcfg[177]
port 774 nsew signal output
rlabel metal2 s 57334 0 57390 800 6 gpio_padcfg[178]
port 775 nsew signal output
rlabel metal2 s 9678 0 9734 800 6 gpio_padcfg[179]
port 776 nsew signal output
rlabel metal3 s 139200 149608 140000 149728 6 gpio_padcfg[17]
port 777 nsew signal output
rlabel metal2 s 23202 439200 23258 440000 6 gpio_padcfg[180]
port 778 nsew signal output
rlabel metal3 s 0 129888 800 130008 6 gpio_padcfg[181]
port 779 nsew signal output
rlabel metal3 s 0 91808 800 91928 6 gpio_padcfg[182]
port 780 nsew signal output
rlabel metal3 s 139200 392368 140000 392488 6 gpio_padcfg[183]
port 781 nsew signal output
rlabel metal3 s 139200 48288 140000 48408 6 gpio_padcfg[184]
port 782 nsew signal output
rlabel metal2 s 20626 439200 20682 440000 6 gpio_padcfg[185]
port 783 nsew signal output
rlabel metal3 s 0 320288 800 320408 6 gpio_padcfg[186]
port 784 nsew signal output
rlabel metal2 s 27066 0 27122 800 6 gpio_padcfg[187]
port 785 nsew signal output
rlabel metal2 s 42522 439200 42578 440000 6 gpio_padcfg[188]
port 786 nsew signal output
rlabel metal2 s 69570 0 69626 800 6 gpio_padcfg[189]
port 787 nsew signal output
rlabel metal3 s 139200 69368 140000 69488 6 gpio_padcfg[18]
port 788 nsew signal output
rlabel metal2 s 8390 0 8446 800 6 gpio_padcfg[190]
port 789 nsew signal output
rlabel metal3 s 0 359728 800 359848 6 gpio_padcfg[191]
port 790 nsew signal output
rlabel metal3 s 0 148928 800 149048 6 gpio_padcfg[19]
port 791 nsew signal output
rlabel metal3 s 0 265208 800 265328 6 gpio_padcfg[1]
port 792 nsew signal output
rlabel metal3 s 0 13608 800 13728 6 gpio_padcfg[20]
port 793 nsew signal output
rlabel metal3 s 0 263848 800 263968 6 gpio_padcfg[21]
port 794 nsew signal output
rlabel metal3 s 0 208768 800 208888 6 gpio_padcfg[22]
port 795 nsew signal output
rlabel metal2 s 28354 0 28410 800 6 gpio_padcfg[23]
port 796 nsew signal output
rlabel metal3 s 139200 121728 140000 121848 6 gpio_padcfg[24]
port 797 nsew signal output
rlabel metal3 s 0 238688 800 238808 6 gpio_padcfg[25]
port 798 nsew signal output
rlabel metal3 s 139200 246848 140000 246968 6 gpio_padcfg[26]
port 799 nsew signal output
rlabel metal3 s 139200 133288 140000 133408 6 gpio_padcfg[27]
port 800 nsew signal output
rlabel metal3 s 139200 210808 140000 210928 6 gpio_padcfg[28]
port 801 nsew signal output
rlabel metal3 s 139200 278128 140000 278248 6 gpio_padcfg[29]
port 802 nsew signal output
rlabel metal3 s 139200 330488 140000 330608 6 gpio_padcfg[2]
port 803 nsew signal output
rlabel metal3 s 139200 187688 140000 187808 6 gpio_padcfg[30]
port 804 nsew signal output
rlabel metal2 s 108210 439200 108266 440000 6 gpio_padcfg[31]
port 805 nsew signal output
rlabel metal2 s 16762 439200 16818 440000 6 gpio_padcfg[32]
port 806 nsew signal output
rlabel metal3 s 0 8848 800 8968 6 gpio_padcfg[33]
port 807 nsew signal output
rlabel metal3 s 0 196528 800 196648 6 gpio_padcfg[34]
port 808 nsew signal output
rlabel metal3 s 0 89768 800 89888 6 gpio_padcfg[35]
port 809 nsew signal output
rlabel metal2 s 113362 0 113418 800 6 gpio_padcfg[36]
port 810 nsew signal output
rlabel metal3 s 0 132608 800 132728 6 gpio_padcfg[37]
port 811 nsew signal output
rlabel metal3 s 0 224408 800 224528 6 gpio_padcfg[38]
port 812 nsew signal output
rlabel metal3 s 139200 212848 140000 212968 6 gpio_padcfg[39]
port 813 nsew signal output
rlabel metal3 s 0 15648 800 15768 6 gpio_padcfg[3]
port 814 nsew signal output
rlabel metal3 s 139200 15648 140000 15768 6 gpio_padcfg[40]
port 815 nsew signal output
rlabel metal3 s 139200 142808 140000 142928 6 gpio_padcfg[41]
port 816 nsew signal output
rlabel metal3 s 0 40128 800 40248 6 gpio_padcfg[42]
port 817 nsew signal output
rlabel metal2 s 123666 439200 123722 440000 6 gpio_padcfg[43]
port 818 nsew signal output
rlabel metal2 s 107566 0 107622 800 6 gpio_padcfg[44]
port 819 nsew signal output
rlabel metal3 s 0 68688 800 68808 6 gpio_padcfg[45]
port 820 nsew signal output
rlabel metal3 s 139200 122408 140000 122528 6 gpio_padcfg[46]
port 821 nsew signal output
rlabel metal3 s 139200 308728 140000 308848 6 gpio_padcfg[47]
port 822 nsew signal output
rlabel metal3 s 139200 314848 140000 314968 6 gpio_padcfg[48]
port 823 nsew signal output
rlabel metal3 s 139200 136688 140000 136808 6 gpio_padcfg[49]
port 824 nsew signal output
rlabel metal3 s 0 335928 800 336048 6 gpio_padcfg[4]
port 825 nsew signal output
rlabel metal2 s 50250 0 50306 800 6 gpio_padcfg[50]
port 826 nsew signal output
rlabel metal3 s 0 163888 800 164008 6 gpio_padcfg[51]
port 827 nsew signal output
rlabel metal3 s 0 146208 800 146328 6 gpio_padcfg[52]
port 828 nsew signal output
rlabel metal2 s 16118 0 16174 800 6 gpio_padcfg[53]
port 829 nsew signal output
rlabel metal3 s 0 57128 800 57248 6 gpio_padcfg[54]
port 830 nsew signal output
rlabel metal3 s 0 323688 800 323808 6 gpio_padcfg[55]
port 831 nsew signal output
rlabel metal3 s 139200 352928 140000 353048 6 gpio_padcfg[56]
port 832 nsew signal output
rlabel metal3 s 0 206728 800 206848 6 gpio_padcfg[57]
port 833 nsew signal output
rlabel metal3 s 0 314848 800 314968 6 gpio_padcfg[58]
port 834 nsew signal output
rlabel metal3 s 0 380128 800 380248 6 gpio_padcfg[59]
port 835 nsew signal output
rlabel metal2 s 16118 439200 16174 440000 6 gpio_padcfg[5]
port 836 nsew signal output
rlabel metal3 s 139200 389648 140000 389768 6 gpio_padcfg[60]
port 837 nsew signal output
rlabel metal2 s 25778 0 25834 800 6 gpio_padcfg[61]
port 838 nsew signal output
rlabel metal3 s 0 256368 800 256488 6 gpio_padcfg[62]
port 839 nsew signal output
rlabel metal3 s 139200 337288 140000 337408 6 gpio_padcfg[63]
port 840 nsew signal output
rlabel metal3 s 0 95888 800 96008 6 gpio_padcfg[64]
port 841 nsew signal output
rlabel metal2 s 71502 439200 71558 440000 6 gpio_padcfg[65]
port 842 nsew signal output
rlabel metal3 s 0 323008 800 323128 6 gpio_padcfg[66]
port 843 nsew signal output
rlabel metal2 s 85670 0 85726 800 6 gpio_padcfg[67]
port 844 nsew signal output
rlabel metal3 s 139200 347488 140000 347608 6 gpio_padcfg[68]
port 845 nsew signal output
rlabel metal2 s 89534 0 89590 800 6 gpio_padcfg[69]
port 846 nsew signal output
rlabel metal3 s 139200 287648 140000 287768 6 gpio_padcfg[6]
port 847 nsew signal output
rlabel metal3 s 139200 331848 140000 331968 6 gpio_padcfg[70]
port 848 nsew signal output
rlabel metal3 s 139200 222368 140000 222488 6 gpio_padcfg[71]
port 849 nsew signal output
rlabel metal3 s 139200 133968 140000 134088 6 gpio_padcfg[72]
port 850 nsew signal output
rlabel metal3 s 0 98608 800 98728 6 gpio_padcfg[73]
port 851 nsew signal output
rlabel metal2 s 126242 0 126298 800 6 gpio_padcfg[74]
port 852 nsew signal output
rlabel metal2 s 33506 0 33562 800 6 gpio_padcfg[75]
port 853 nsew signal output
rlabel metal2 s 7102 439200 7158 440000 6 gpio_padcfg[76]
port 854 nsew signal output
rlabel metal2 s 54758 0 54814 800 6 gpio_padcfg[77]
port 855 nsew signal output
rlabel metal3 s 0 108128 800 108248 6 gpio_padcfg[78]
port 856 nsew signal output
rlabel metal3 s 139200 282888 140000 283008 6 gpio_padcfg[79]
port 857 nsew signal output
rlabel metal3 s 0 147568 800 147688 6 gpio_padcfg[7]
port 858 nsew signal output
rlabel metal3 s 139200 1368 140000 1488 6 gpio_padcfg[80]
port 859 nsew signal output
rlabel metal2 s 18 439200 74 440000 6 gpio_padcfg[81]
port 860 nsew signal output
rlabel metal3 s 139200 387608 140000 387728 6 gpio_padcfg[82]
port 861 nsew signal output
rlabel metal3 s 0 342048 800 342168 6 gpio_padcfg[83]
port 862 nsew signal output
rlabel metal3 s 139200 215568 140000 215688 6 gpio_padcfg[84]
port 863 nsew signal output
rlabel metal3 s 0 77528 800 77648 6 gpio_padcfg[85]
port 864 nsew signal output
rlabel metal2 s 83094 0 83150 800 6 gpio_padcfg[86]
port 865 nsew signal output
rlabel metal3 s 139200 227808 140000 227928 6 gpio_padcfg[87]
port 866 nsew signal output
rlabel metal3 s 139200 104048 140000 104168 6 gpio_padcfg[88]
port 867 nsew signal output
rlabel metal3 s 139200 64608 140000 64728 6 gpio_padcfg[89]
port 868 nsew signal output
rlabel metal3 s 0 180888 800 181008 6 gpio_padcfg[8]
port 869 nsew signal output
rlabel metal2 s 25134 0 25190 800 6 gpio_padcfg[90]
port 870 nsew signal output
rlabel metal3 s 0 30608 800 30728 6 gpio_padcfg[91]
port 871 nsew signal output
rlabel metal3 s 139200 27888 140000 28008 6 gpio_padcfg[92]
port 872 nsew signal output
rlabel metal2 s 19338 0 19394 800 6 gpio_padcfg[93]
port 873 nsew signal output
rlabel metal3 s 0 334568 800 334688 6 gpio_padcfg[94]
port 874 nsew signal output
rlabel metal3 s 139200 269288 140000 269408 6 gpio_padcfg[95]
port 875 nsew signal output
rlabel metal2 s 134614 439200 134670 440000 6 gpio_padcfg[96]
port 876 nsew signal output
rlabel metal3 s 0 123768 800 123888 6 gpio_padcfg[97]
port 877 nsew signal output
rlabel metal2 s 36082 439200 36138 440000 6 gpio_padcfg[98]
port 878 nsew signal output
rlabel metal3 s 0 136008 800 136128 6 gpio_padcfg[99]
port 879 nsew signal output
rlabel metal2 s 103702 0 103758 800 6 gpio_padcfg[9]
port 880 nsew signal output
rlabel metal3 s 139200 183608 140000 183728 6 io_oeb_pll[0]
port 881 nsew signal output
rlabel metal3 s 0 227808 800 227928 6 io_oeb_pll[10]
port 882 nsew signal output
rlabel metal3 s 0 159128 800 159248 6 io_oeb_pll[11]
port 883 nsew signal output
rlabel metal3 s 0 164568 800 164688 6 io_oeb_pll[12]
port 884 nsew signal output
rlabel metal3 s 139200 265208 140000 265328 6 io_oeb_pll[13]
port 885 nsew signal output
rlabel metal3 s 139200 165248 140000 165368 6 io_oeb_pll[14]
port 886 nsew signal output
rlabel metal3 s 0 10208 800 10328 6 io_oeb_pll[15]
port 887 nsew signal output
rlabel metal3 s 139200 267248 140000 267368 6 io_oeb_pll[16]
port 888 nsew signal output
rlabel metal3 s 0 423648 800 423768 6 io_oeb_pll[17]
port 889 nsew signal output
rlabel metal2 s 18050 0 18106 800 6 io_oeb_pll[18]
port 890 nsew signal output
rlabel metal3 s 139200 95208 140000 95328 6 io_oeb_pll[19]
port 891 nsew signal output
rlabel metal2 s 91466 439200 91522 440000 6 io_oeb_pll[1]
port 892 nsew signal output
rlabel metal2 s 88246 439200 88302 440000 6 io_oeb_pll[20]
port 893 nsew signal output
rlabel metal3 s 0 272688 800 272808 6 io_oeb_pll[21]
port 894 nsew signal output
rlabel metal3 s 0 282208 800 282328 6 io_oeb_pll[22]
port 895 nsew signal output
rlabel metal3 s 139200 138728 140000 138848 6 io_oeb_pll[23]
port 896 nsew signal output
rlabel metal3 s 139200 360408 140000 360528 6 io_oeb_pll[24]
port 897 nsew signal output
rlabel metal2 s 48318 0 48374 800 6 io_oeb_pll[25]
port 898 nsew signal output
rlabel metal3 s 139200 324368 140000 324488 6 io_oeb_pll[26]
port 899 nsew signal output
rlabel metal2 s 133326 0 133382 800 6 io_oeb_pll[27]
port 900 nsew signal output
rlabel metal3 s 0 44208 800 44328 6 io_oeb_pll[28]
port 901 nsew signal output
rlabel metal3 s 0 48288 800 48408 6 io_oeb_pll[29]
port 902 nsew signal output
rlabel metal3 s 139200 217608 140000 217728 6 io_oeb_pll[2]
port 903 nsew signal output
rlabel metal2 s 2594 0 2650 800 6 io_oeb_pll[30]
port 904 nsew signal output
rlabel metal3 s 139200 225768 140000 225888 6 io_oeb_pll[31]
port 905 nsew signal output
rlabel metal2 s 55402 0 55458 800 6 io_oeb_pll[32]
port 906 nsew signal output
rlabel metal3 s 0 222368 800 222488 6 io_oeb_pll[33]
port 907 nsew signal output
rlabel metal3 s 139200 300568 140000 300688 6 io_oeb_pll[34]
port 908 nsew signal output
rlabel metal2 s 92754 439200 92810 440000 6 io_oeb_pll[35]
port 909 nsew signal output
rlabel metal3 s 139200 40128 140000 40248 6 io_oeb_pll[36]
port 910 nsew signal output
rlabel metal3 s 0 437928 800 438048 6 io_oeb_pll[37]
port 911 nsew signal output
rlabel metal3 s 0 218968 800 219088 6 io_oeb_pll[3]
port 912 nsew signal output
rlabel metal2 s 131394 439200 131450 440000 6 io_oeb_pll[4]
port 913 nsew signal output
rlabel metal3 s 0 391688 800 391808 6 io_oeb_pll[5]
port 914 nsew signal output
rlabel metal3 s 139200 68688 140000 68808 6 io_oeb_pll[6]
port 915 nsew signal output
rlabel metal3 s 139200 261128 140000 261248 6 io_oeb_pll[7]
port 916 nsew signal output
rlabel metal3 s 139200 117648 140000 117768 6 io_oeb_pll[8]
port 917 nsew signal output
rlabel metal3 s 139200 377408 140000 377528 6 io_oeb_pll[9]
port 918 nsew signal output
rlabel metal3 s 139200 373328 140000 373448 6 io_out_pll[0]
port 919 nsew signal output
rlabel metal2 s 95330 0 95386 800 6 io_out_pll[10]
port 920 nsew signal output
rlabel metal3 s 139200 370608 140000 370728 6 io_out_pll[11]
port 921 nsew signal output
rlabel metal3 s 0 245488 800 245608 6 io_out_pll[12]
port 922 nsew signal output
rlabel metal3 s 139200 404608 140000 404728 6 io_out_pll[13]
port 923 nsew signal output
rlabel metal3 s 0 226448 800 226568 6 io_out_pll[14]
port 924 nsew signal output
rlabel metal2 s 75366 439200 75422 440000 6 io_out_pll[15]
port 925 nsew signal output
rlabel metal3 s 139200 72768 140000 72888 6 io_out_pll[16]
port 926 nsew signal output
rlabel metal3 s 139200 240048 140000 240168 6 io_out_pll[17]
port 927 nsew signal output
rlabel metal3 s 139200 41488 140000 41608 6 io_out_pll[18]
port 928 nsew signal output
rlabel metal2 s 99194 0 99250 800 6 io_out_pll[19]
port 929 nsew signal output
rlabel metal3 s 139200 121048 140000 121168 6 io_out_pll[1]
port 930 nsew signal output
rlabel metal3 s 0 430448 800 430568 6 io_out_pll[20]
port 931 nsew signal output
rlabel metal3 s 139200 357688 140000 357808 6 io_out_pll[21]
port 932 nsew signal output
rlabel metal3 s 139200 315528 140000 315648 6 io_out_pll[22]
port 933 nsew signal output
rlabel metal3 s 139200 9528 140000 9648 6 io_out_pll[23]
port 934 nsew signal output
rlabel metal3 s 0 52368 800 52488 6 io_out_pll[24]
port 935 nsew signal output
rlabel metal3 s 0 35368 800 35488 6 io_out_pll[25]
port 936 nsew signal output
rlabel metal3 s 0 70728 800 70848 6 io_out_pll[2]
port 937 nsew signal output
rlabel metal2 s 28354 439200 28410 440000 6 io_out_pll[3]
port 938 nsew signal output
rlabel metal3 s 139200 380128 140000 380248 6 io_out_pll[4]
port 939 nsew signal output
rlabel metal2 s 88890 439200 88946 440000 6 io_out_pll[5]
port 940 nsew signal output
rlabel metal2 s 22558 439200 22614 440000 6 io_out_pll[6]
port 941 nsew signal output
rlabel metal3 s 0 316208 800 316328 6 io_out_pll[7]
port 942 nsew signal output
rlabel metal3 s 139200 276768 140000 276888 6 io_out_pll[8]
port 943 nsew signal output
rlabel metal3 s 0 231888 800 232008 6 io_out_pll[9]
port 944 nsew signal output
rlabel metal2 s 122378 0 122434 800 6 irq_o[0]
port 945 nsew signal output
rlabel metal3 s 139200 223048 140000 223168 6 irq_o[10]
port 946 nsew signal output
rlabel metal3 s 139200 94528 140000 94648 6 irq_o[11]
port 947 nsew signal output
rlabel metal3 s 139200 57128 140000 57248 6 irq_o[12]
port 948 nsew signal output
rlabel metal2 s 78586 439200 78642 440000 6 irq_o[13]
port 949 nsew signal output
rlabel metal2 s 138478 0 138534 800 6 irq_o[14]
port 950 nsew signal output
rlabel metal3 s 139200 147568 140000 147688 6 irq_o[15]
port 951 nsew signal output
rlabel metal3 s 139200 87048 140000 87168 6 irq_o[16]
port 952 nsew signal output
rlabel metal3 s 0 306008 800 306128 6 irq_o[17]
port 953 nsew signal output
rlabel metal2 s 54114 0 54170 800 6 irq_o[18]
port 954 nsew signal output
rlabel metal3 s 0 229848 800 229968 6 irq_o[19]
port 955 nsew signal output
rlabel metal3 s 0 320968 800 321088 6 irq_o[1]
port 956 nsew signal output
rlabel metal3 s 0 120368 800 120488 6 irq_o[20]
port 957 nsew signal output
rlabel metal3 s 139200 295128 140000 295248 6 irq_o[21]
port 958 nsew signal output
rlabel metal3 s 0 121048 800 121168 6 irq_o[22]
port 959 nsew signal output
rlabel metal3 s 139200 280848 140000 280968 6 irq_o[23]
port 960 nsew signal output
rlabel metal3 s 0 36048 800 36168 6 irq_o[24]
port 961 nsew signal output
rlabel metal3 s 0 61208 800 61328 6 irq_o[25]
port 962 nsew signal output
rlabel metal2 s 12254 439200 12310 440000 6 irq_o[26]
port 963 nsew signal output
rlabel metal3 s 0 198568 800 198688 6 irq_o[27]
port 964 nsew signal output
rlabel metal2 s 10322 0 10378 800 6 irq_o[28]
port 965 nsew signal output
rlabel metal3 s 139200 435888 140000 436008 6 irq_o[29]
port 966 nsew signal output
rlabel metal3 s 0 178848 800 178968 6 irq_o[2]
port 967 nsew signal output
rlabel metal3 s 0 179528 800 179648 6 irq_o[30]
port 968 nsew signal output
rlabel metal2 s 18050 439200 18106 440000 6 irq_o[31]
port 969 nsew signal output
rlabel metal3 s 139200 70728 140000 70848 6 irq_o[3]
port 970 nsew signal output
rlabel metal3 s 0 426368 800 426488 6 irq_o[4]
port 971 nsew signal output
rlabel metal3 s 139200 220328 140000 220448 6 irq_o[5]
port 972 nsew signal output
rlabel metal3 s 0 85008 800 85128 6 irq_o[6]
port 973 nsew signal output
rlabel metal3 s 0 392368 800 392488 6 irq_o[7]
port 974 nsew signal output
rlabel metal3 s 0 176128 800 176248 6 irq_o[8]
port 975 nsew signal output
rlabel metal3 s 0 235288 800 235408 6 irq_o[9]
port 976 nsew signal output
rlabel metal3 s 139200 361768 140000 361888 6 la_data_out_pll[0]
port 977 nsew signal output
rlabel metal2 s 121090 439200 121146 440000 6 la_data_out_pll[10]
port 978 nsew signal output
rlabel metal2 s 17406 0 17462 800 6 la_data_out_pll[11]
port 979 nsew signal output
rlabel metal3 s 139200 304648 140000 304768 6 la_data_out_pll[12]
port 980 nsew signal output
rlabel metal3 s 0 257048 800 257168 6 la_data_out_pll[13]
port 981 nsew signal output
rlabel metal3 s 139200 248208 140000 248328 6 la_data_out_pll[14]
port 982 nsew signal output
rlabel metal3 s 139200 426368 140000 426488 6 la_data_out_pll[15]
port 983 nsew signal output
rlabel metal3 s 139200 34688 140000 34808 6 la_data_out_pll[16]
port 984 nsew signal output
rlabel metal3 s 0 283568 800 283688 6 la_data_out_pll[17]
port 985 nsew signal output
rlabel metal2 s 43810 439200 43866 440000 6 la_data_out_pll[18]
port 986 nsew signal output
rlabel metal3 s 139200 244808 140000 244928 6 la_data_out_pll[19]
port 987 nsew signal output
rlabel metal3 s 0 14968 800 15088 6 la_data_out_pll[1]
port 988 nsew signal output
rlabel metal3 s 0 304648 800 304768 6 la_data_out_pll[20]
port 989 nsew signal output
rlabel metal3 s 139200 367888 140000 368008 6 la_data_out_pll[21]
port 990 nsew signal output
rlabel metal3 s 139200 254328 140000 254448 6 la_data_out_pll[22]
port 991 nsew signal output
rlabel metal3 s 139200 132608 140000 132728 6 la_data_out_pll[23]
port 992 nsew signal output
rlabel metal3 s 0 278128 800 278248 6 la_data_out_pll[24]
port 993 nsew signal output
rlabel metal3 s 0 197208 800 197328 6 la_data_out_pll[25]
port 994 nsew signal output
rlabel metal3 s 139200 359048 140000 359168 6 la_data_out_pll[26]
port 995 nsew signal output
rlabel metal2 s 5814 439200 5870 440000 6 la_data_out_pll[27]
port 996 nsew signal output
rlabel metal2 s 15474 439200 15530 440000 6 la_data_out_pll[28]
port 997 nsew signal output
rlabel metal3 s 139200 244128 140000 244248 6 la_data_out_pll[29]
port 998 nsew signal output
rlabel metal3 s 0 165928 800 166048 6 la_data_out_pll[2]
port 999 nsew signal output
rlabel metal3 s 0 384208 800 384328 6 la_data_out_pll[30]
port 1000 nsew signal output
rlabel metal3 s 0 388288 800 388408 6 la_data_out_pll[31]
port 1001 nsew signal output
rlabel metal3 s 139200 329808 140000 329928 6 la_data_out_pll[32]
port 1002 nsew signal output
rlabel metal3 s 0 168648 800 168768 6 la_data_out_pll[33]
port 1003 nsew signal output
rlabel metal3 s 0 174768 800 174888 6 la_data_out_pll[34]
port 1004 nsew signal output
rlabel metal3 s 0 189048 800 189168 6 la_data_out_pll[35]
port 1005 nsew signal output
rlabel metal3 s 0 39448 800 39568 6 la_data_out_pll[36]
port 1006 nsew signal output
rlabel metal3 s 139200 150968 140000 151088 6 la_data_out_pll[37]
port 1007 nsew signal output
rlabel metal3 s 139200 265888 140000 266008 6 la_data_out_pll[38]
port 1008 nsew signal output
rlabel metal2 s 71502 0 71558 800 6 la_data_out_pll[39]
port 1009 nsew signal output
rlabel metal3 s 139200 294448 140000 294568 6 la_data_out_pll[3]
port 1010 nsew signal output
rlabel metal3 s 139200 316208 140000 316328 6 la_data_out_pll[40]
port 1011 nsew signal output
rlabel metal3 s 139200 103368 140000 103488 6 la_data_out_pll[41]
port 1012 nsew signal output
rlabel metal3 s 139200 390328 140000 390448 6 la_data_out_pll[42]
port 1013 nsew signal output
rlabel metal2 s 136546 439200 136602 440000 6 la_data_out_pll[43]
port 1014 nsew signal output
rlabel metal2 s 36726 439200 36782 440000 6 la_data_out_pll[44]
port 1015 nsew signal output
rlabel metal3 s 0 103368 800 103488 6 la_data_out_pll[45]
port 1016 nsew signal output
rlabel metal3 s 139200 385568 140000 385688 6 la_data_out_pll[46]
port 1017 nsew signal output
rlabel metal3 s 139200 153688 140000 153808 6 la_data_out_pll[47]
port 1018 nsew signal output
rlabel metal3 s 0 285608 800 285728 6 la_data_out_pll[48]
port 1019 nsew signal output
rlabel metal2 s 139122 0 139178 800 6 la_data_out_pll[49]
port 1020 nsew signal output
rlabel metal3 s 139200 120368 140000 120488 6 la_data_out_pll[4]
port 1021 nsew signal output
rlabel metal3 s 139200 259768 140000 259888 6 la_data_out_pll[50]
port 1022 nsew signal output
rlabel metal3 s 139200 47608 140000 47728 6 la_data_out_pll[51]
port 1023 nsew signal output
rlabel metal3 s 0 277448 800 277568 6 la_data_out_pll[52]
port 1024 nsew signal output
rlabel metal2 s 138478 439200 138534 440000 6 la_data_out_pll[53]
port 1025 nsew signal output
rlabel metal2 s 137834 0 137890 800 6 la_data_out_pll[54]
port 1026 nsew signal output
rlabel metal3 s 139200 37408 140000 37528 6 la_data_out_pll[55]
port 1027 nsew signal output
rlabel metal3 s 0 348848 800 348968 6 la_data_out_pll[56]
port 1028 nsew signal output
rlabel metal3 s 139200 393728 140000 393848 6 la_data_out_pll[57]
port 1029 nsew signal output
rlabel metal3 s 139200 224408 140000 224528 6 la_data_out_pll[58]
port 1030 nsew signal output
rlabel metal3 s 139200 428408 140000 428528 6 la_data_out_pll[59]
port 1031 nsew signal output
rlabel metal3 s 139200 257048 140000 257168 6 la_data_out_pll[5]
port 1032 nsew signal output
rlabel metal3 s 139200 309408 140000 309528 6 la_data_out_pll[60]
port 1033 nsew signal output
rlabel metal3 s 139200 106768 140000 106888 6 la_data_out_pll[61]
port 1034 nsew signal output
rlabel metal3 s 0 246848 800 246968 6 la_data_out_pll[62]
port 1035 nsew signal output
rlabel metal3 s 0 228488 800 228608 6 la_data_out_pll[63]
port 1036 nsew signal output
rlabel metal2 s 3238 0 3294 800 6 la_data_out_pll[6]
port 1037 nsew signal output
rlabel metal3 s 0 358368 800 358488 6 la_data_out_pll[7]
port 1038 nsew signal output
rlabel metal3 s 139200 409368 140000 409488 6 la_data_out_pll[8]
port 1039 nsew signal output
rlabel metal3 s 0 88408 800 88528 6 la_data_out_pll[9]
port 1040 nsew signal output
rlabel metal2 s 80518 0 80574 800 6 rst_n
port 1041 nsew signal input
rlabel metal3 s 139200 164568 140000 164688 6 rstn_i_pll
port 1042 nsew signal input
rlabel metal2 s 6458 0 6514 800 6 rstn_o_pll
port 1043 nsew signal output
rlabel metal3 s 139200 342048 140000 342168 6 scan_en_i_pll
port 1044 nsew signal input
rlabel metal3 s 139200 363808 140000 363928 6 scan_i_pll
port 1045 nsew signal input
rlabel metal3 s 139200 417528 140000 417648 6 scan_o_pll
port 1046 nsew signal output
rlabel metal3 s 0 414808 800 414928 6 scl_pad_i
port 1047 nsew signal input
rlabel metal3 s 0 19728 800 19848 6 scl_pad_o
port 1048 nsew signal output
rlabel metal3 s 0 163208 800 163328 6 scl_padoen_o
port 1049 nsew signal output
rlabel metal3 s 0 204688 800 204808 6 sda_pad_i
port 1050 nsew signal input
rlabel metal2 s 66994 0 67050 800 6 sda_pad_o
port 1051 nsew signal output
rlabel metal3 s 0 156408 800 156528 6 sda_padoen_o
port 1052 nsew signal output
rlabel metal3 s 0 225768 800 225888 6 slave_ar_addr[0]
port 1053 nsew signal input
rlabel metal3 s 0 418888 800 419008 6 slave_ar_addr[10]
port 1054 nsew signal input
rlabel metal2 s 66994 439200 67050 440000 6 slave_ar_addr[11]
port 1055 nsew signal input
rlabel metal3 s 0 223728 800 223848 6 slave_ar_addr[12]
port 1056 nsew signal input
rlabel metal3 s 0 417528 800 417648 6 slave_ar_addr[13]
port 1057 nsew signal input
rlabel metal2 s 3238 439200 3294 440000 6 slave_ar_addr[14]
port 1058 nsew signal input
rlabel metal3 s 0 406648 800 406768 6 slave_ar_addr[15]
port 1059 nsew signal input
rlabel metal3 s 0 266568 800 266688 6 slave_ar_addr[16]
port 1060 nsew signal input
rlabel metal2 s 106922 439200 106978 440000 6 slave_ar_addr[17]
port 1061 nsew signal input
rlabel metal2 s 127530 439200 127586 440000 6 slave_ar_addr[18]
port 1062 nsew signal input
rlabel metal3 s 139200 151648 140000 151768 6 slave_ar_addr[19]
port 1063 nsew signal input
rlabel metal3 s 139200 91128 140000 91248 6 slave_ar_addr[1]
port 1064 nsew signal input
rlabel metal3 s 0 99288 800 99408 6 slave_ar_addr[20]
port 1065 nsew signal input
rlabel metal3 s 139200 14288 140000 14408 6 slave_ar_addr[21]
port 1066 nsew signal input
rlabel metal3 s 139200 397808 140000 397928 6 slave_ar_addr[22]
port 1067 nsew signal input
rlabel metal3 s 0 61888 800 62008 6 slave_ar_addr[23]
port 1068 nsew signal input
rlabel metal3 s 0 397128 800 397248 6 slave_ar_addr[24]
port 1069 nsew signal input
rlabel metal3 s 139200 334568 140000 334688 6 slave_ar_addr[25]
port 1070 nsew signal input
rlabel metal3 s 0 398488 800 398608 6 slave_ar_addr[26]
port 1071 nsew signal input
rlabel metal3 s 0 338648 800 338768 6 slave_ar_addr[27]
port 1072 nsew signal input
rlabel metal2 s 75366 0 75422 800 6 slave_ar_addr[28]
port 1073 nsew signal input
rlabel metal3 s 0 310768 800 310888 6 slave_ar_addr[29]
port 1074 nsew signal input
rlabel metal3 s 0 54408 800 54528 6 slave_ar_addr[2]
port 1075 nsew signal input
rlabel metal3 s 139200 78208 140000 78328 6 slave_ar_addr[30]
port 1076 nsew signal input
rlabel metal3 s 139200 312808 140000 312928 6 slave_ar_addr[31]
port 1077 nsew signal input
rlabel metal3 s 0 112888 800 113008 6 slave_ar_addr[3]
port 1078 nsew signal input
rlabel metal3 s 139200 336608 140000 336728 6 slave_ar_addr[4]
port 1079 nsew signal input
rlabel metal3 s 0 3408 800 3528 6 slave_ar_addr[5]
port 1080 nsew signal input
rlabel metal2 s 19982 439200 20038 440000 6 slave_ar_addr[6]
port 1081 nsew signal input
rlabel metal3 s 139200 4768 140000 4888 6 slave_ar_addr[7]
port 1082 nsew signal input
rlabel metal3 s 139200 429768 140000 429888 6 slave_ar_addr[8]
port 1083 nsew signal input
rlabel metal3 s 139200 51688 140000 51808 6 slave_ar_addr[9]
port 1084 nsew signal input
rlabel metal3 s 0 42848 800 42968 6 slave_ar_burst[0]
port 1085 nsew signal input
rlabel metal2 s 118514 439200 118570 440000 6 slave_ar_burst[1]
port 1086 nsew signal input
rlabel metal3 s 0 404608 800 404728 6 slave_ar_cache[0]
port 1087 nsew signal input
rlabel metal3 s 139200 328448 140000 328568 6 slave_ar_cache[1]
port 1088 nsew signal input
rlabel metal3 s 0 361768 800 361888 6 slave_ar_cache[2]
port 1089 nsew signal input
rlabel metal3 s 0 189728 800 189848 6 slave_ar_cache[3]
port 1090 nsew signal input
rlabel metal2 s 94042 0 94098 800 6 slave_ar_id[0]
port 1091 nsew signal input
rlabel metal2 s 82450 439200 82506 440000 6 slave_ar_id[1]
port 1092 nsew signal input
rlabel metal3 s 0 104048 800 104168 6 slave_ar_id[2]
port 1093 nsew signal input
rlabel metal3 s 0 177488 800 177608 6 slave_ar_id[3]
port 1094 nsew signal input
rlabel metal3 s 0 128528 800 128648 6 slave_ar_id[4]
port 1095 nsew signal input
rlabel metal3 s 0 432488 800 432608 6 slave_ar_id[5]
port 1096 nsew signal input
rlabel metal3 s 0 344768 800 344888 6 slave_ar_len[0]
port 1097 nsew signal input
rlabel metal3 s 139200 311448 140000 311568 6 slave_ar_len[1]
port 1098 nsew signal input
rlabel metal3 s 139200 195848 140000 195968 6 slave_ar_len[2]
port 1099 nsew signal input
rlabel metal3 s 139200 205368 140000 205488 6 slave_ar_len[3]
port 1100 nsew signal input
rlabel metal2 s 114650 439200 114706 440000 6 slave_ar_len[4]
port 1101 nsew signal input
rlabel metal3 s 0 337288 800 337408 6 slave_ar_len[5]
port 1102 nsew signal input
rlabel metal3 s 139200 6808 140000 6928 6 slave_ar_len[6]
port 1103 nsew signal input
rlabel metal2 s 81162 0 81218 800 6 slave_ar_len[7]
port 1104 nsew signal input
rlabel metal3 s 139200 427728 140000 427848 6 slave_ar_lock
port 1105 nsew signal input
rlabel metal3 s 139200 163208 140000 163328 6 slave_ar_prot[0]
port 1106 nsew signal input
rlabel metal3 s 0 79568 800 79688 6 slave_ar_prot[1]
port 1107 nsew signal input
rlabel metal2 s 10322 439200 10378 440000 6 slave_ar_prot[2]
port 1108 nsew signal input
rlabel metal3 s 139200 310768 140000 310888 6 slave_ar_qos[0]
port 1109 nsew signal input
rlabel metal2 s 92110 439200 92166 440000 6 slave_ar_qos[1]
port 1110 nsew signal input
rlabel metal3 s 0 117648 800 117768 6 slave_ar_qos[2]
port 1111 nsew signal input
rlabel metal3 s 139200 48968 140000 49088 6 slave_ar_qos[3]
port 1112 nsew signal input
rlabel metal2 s 119158 439200 119214 440000 6 slave_ar_ready
port 1113 nsew signal output
rlabel metal3 s 139200 145528 140000 145648 6 slave_ar_region[0]
port 1114 nsew signal input
rlabel metal3 s 0 221688 800 221808 6 slave_ar_region[1]
port 1115 nsew signal input
rlabel metal3 s 0 401208 800 401328 6 slave_ar_region[2]
port 1116 nsew signal input
rlabel metal2 s 34150 0 34206 800 6 slave_ar_region[3]
port 1117 nsew signal input
rlabel metal2 s 101126 439200 101182 440000 6 slave_ar_size[0]
port 1118 nsew signal input
rlabel metal3 s 139200 19728 140000 19848 6 slave_ar_size[1]
port 1119 nsew signal input
rlabel metal3 s 139200 312128 140000 312248 6 slave_ar_size[2]
port 1120 nsew signal input
rlabel metal3 s 139200 142128 140000 142248 6 slave_ar_user[0]
port 1121 nsew signal input
rlabel metal2 s 129462 0 129518 800 6 slave_ar_user[1]
port 1122 nsew signal input
rlabel metal3 s 0 64608 800 64728 6 slave_ar_user[2]
port 1123 nsew signal input
rlabel metal2 s 9034 439200 9090 440000 6 slave_ar_user[3]
port 1124 nsew signal input
rlabel metal2 s 77298 0 77354 800 6 slave_ar_user[4]
port 1125 nsew signal input
rlabel metal3 s 0 431808 800 431928 6 slave_ar_user[5]
port 1126 nsew signal input
rlabel metal3 s 139200 339328 140000 339448 6 slave_ar_valid
port 1127 nsew signal input
rlabel metal3 s 139200 214888 140000 215008 6 slave_aw_addr[0]
port 1128 nsew signal input
rlabel metal3 s 0 261128 800 261248 6 slave_aw_addr[10]
port 1129 nsew signal input
rlabel metal3 s 0 276768 800 276888 6 slave_aw_addr[11]
port 1130 nsew signal input
rlabel metal3 s 139200 430448 140000 430568 6 slave_aw_addr[12]
port 1131 nsew signal input
rlabel metal3 s 0 85688 800 85808 6 slave_aw_addr[13]
port 1132 nsew signal input
rlabel metal3 s 139200 188368 140000 188488 6 slave_aw_addr[14]
port 1133 nsew signal input
rlabel metal3 s 0 439288 800 439408 6 slave_aw_addr[15]
port 1134 nsew signal input
rlabel metal2 s 63774 439200 63830 440000 6 slave_aw_addr[16]
port 1135 nsew signal input
rlabel metal3 s 0 244808 800 244928 6 slave_aw_addr[17]
port 1136 nsew signal input
rlabel metal3 s 139200 70048 140000 70168 6 slave_aw_addr[18]
port 1137 nsew signal input
rlabel metal3 s 0 58488 800 58608 6 slave_aw_addr[19]
port 1138 nsew signal input
rlabel metal2 s 32218 439200 32274 440000 6 slave_aw_addr[1]
port 1139 nsew signal input
rlabel metal2 s 70214 0 70270 800 6 slave_aw_addr[20]
port 1140 nsew signal input
rlabel metal3 s 0 182928 800 183048 6 slave_aw_addr[21]
port 1141 nsew signal input
rlabel metal3 s 139200 398488 140000 398608 6 slave_aw_addr[22]
port 1142 nsew signal input
rlabel metal3 s 139200 74808 140000 74928 6 slave_aw_addr[23]
port 1143 nsew signal input
rlabel metal3 s 139200 363128 140000 363248 6 slave_aw_addr[24]
port 1144 nsew signal input
rlabel metal3 s 0 227128 800 227248 6 slave_aw_addr[25]
port 1145 nsew signal input
rlabel metal3 s 0 112208 800 112328 6 slave_aw_addr[26]
port 1146 nsew signal input
rlabel metal3 s 139200 305328 140000 305448 6 slave_aw_addr[27]
port 1147 nsew signal input
rlabel metal3 s 139200 344768 140000 344888 6 slave_aw_addr[28]
port 1148 nsew signal input
rlabel metal2 s 126886 0 126942 800 6 slave_aw_addr[29]
port 1149 nsew signal input
rlabel metal2 s 97262 439200 97318 440000 6 slave_aw_addr[2]
port 1150 nsew signal input
rlabel metal3 s 139200 74128 140000 74248 6 slave_aw_addr[30]
port 1151 nsew signal input
rlabel metal2 s 137190 439200 137246 440000 6 slave_aw_addr[31]
port 1152 nsew signal input
rlabel metal3 s 0 82968 800 83088 6 slave_aw_addr[3]
port 1153 nsew signal input
rlabel metal3 s 139200 173408 140000 173528 6 slave_aw_addr[4]
port 1154 nsew signal input
rlabel metal3 s 139200 111528 140000 111648 6 slave_aw_addr[5]
port 1155 nsew signal input
rlabel metal2 s 28998 0 29054 800 6 slave_aw_addr[6]
port 1156 nsew signal input
rlabel metal2 s 45098 0 45154 800 6 slave_aw_addr[7]
port 1157 nsew signal input
rlabel metal3 s 0 223048 800 223168 6 slave_aw_addr[8]
port 1158 nsew signal input
rlabel metal3 s 139200 322328 140000 322448 6 slave_aw_addr[9]
port 1159 nsew signal input
rlabel metal3 s 0 142808 800 142928 6 slave_aw_burst[0]
port 1160 nsew signal input
rlabel metal3 s 139200 423648 140000 423768 6 slave_aw_burst[1]
port 1161 nsew signal input
rlabel metal3 s 0 170688 800 170808 6 slave_aw_cache[0]
port 1162 nsew signal input
rlabel metal3 s 0 80928 800 81048 6 slave_aw_cache[1]
port 1163 nsew signal input
rlabel metal3 s 0 235968 800 236088 6 slave_aw_cache[2]
port 1164 nsew signal input
rlabel metal3 s 0 62568 800 62688 6 slave_aw_cache[3]
port 1165 nsew signal input
rlabel metal2 s 131394 0 131450 800 6 slave_aw_id[0]
port 1166 nsew signal input
rlabel metal3 s 0 142128 800 142248 6 slave_aw_id[1]
port 1167 nsew signal input
rlabel metal2 s 59910 439200 59966 440000 6 slave_aw_id[2]
port 1168 nsew signal input
rlabel metal3 s 139200 321648 140000 321768 6 slave_aw_id[3]
port 1169 nsew signal input
rlabel metal2 s 72790 439200 72846 440000 6 slave_aw_id[4]
port 1170 nsew signal input
rlabel metal3 s 139200 89768 140000 89888 6 slave_aw_id[5]
port 1171 nsew signal input
rlabel metal3 s 0 216928 800 217048 6 slave_aw_len[0]
port 1172 nsew signal input
rlabel metal3 s 0 4768 800 4888 6 slave_aw_len[1]
port 1173 nsew signal input
rlabel metal3 s 0 151648 800 151768 6 slave_aw_len[2]
port 1174 nsew signal input
rlabel metal3 s 0 68008 800 68128 6 slave_aw_len[3]
port 1175 nsew signal input
rlabel metal2 s 57978 0 58034 800 6 slave_aw_len[4]
port 1176 nsew signal input
rlabel metal3 s 139200 197208 140000 197328 6 slave_aw_len[5]
port 1177 nsew signal input
rlabel metal3 s 139200 235968 140000 236088 6 slave_aw_len[6]
port 1178 nsew signal input
rlabel metal2 s 62486 439200 62542 440000 6 slave_aw_len[7]
port 1179 nsew signal input
rlabel metal3 s 139200 384208 140000 384328 6 slave_aw_lock
port 1180 nsew signal input
rlabel metal3 s 0 29928 800 30048 6 slave_aw_prot[0]
port 1181 nsew signal input
rlabel metal3 s 139200 60528 140000 60648 6 slave_aw_prot[1]
port 1182 nsew signal input
rlabel metal3 s 139200 160488 140000 160608 6 slave_aw_prot[2]
port 1183 nsew signal input
rlabel metal3 s 139200 12248 140000 12368 6 slave_aw_qos[0]
port 1184 nsew signal input
rlabel metal3 s 0 272008 800 272128 6 slave_aw_qos[1]
port 1185 nsew signal input
rlabel metal3 s 139200 85688 140000 85808 6 slave_aw_qos[2]
port 1186 nsew signal input
rlabel metal3 s 139200 175448 140000 175568 6 slave_aw_qos[3]
port 1187 nsew signal input
rlabel metal3 s 139200 110848 140000 110968 6 slave_aw_ready
port 1188 nsew signal output
rlabel metal2 s 108854 0 108910 800 6 slave_aw_region[0]
port 1189 nsew signal input
rlabel metal2 s 66350 439200 66406 440000 6 slave_aw_region[1]
port 1190 nsew signal input
rlabel metal3 s 139200 65288 140000 65408 6 slave_aw_region[2]
port 1191 nsew signal input
rlabel metal3 s 139200 318248 140000 318368 6 slave_aw_region[3]
port 1192 nsew signal input
rlabel metal3 s 139200 253648 140000 253768 6 slave_aw_size[0]
port 1193 nsew signal input
rlabel metal3 s 139200 367208 140000 367328 6 slave_aw_size[1]
port 1194 nsew signal input
rlabel metal3 s 139200 345448 140000 345568 6 slave_aw_size[2]
port 1195 nsew signal input
rlabel metal3 s 0 34688 800 34808 6 slave_aw_user[0]
port 1196 nsew signal input
rlabel metal2 s 5814 0 5870 800 6 slave_aw_user[1]
port 1197 nsew signal input
rlabel metal3 s 139200 146888 140000 147008 6 slave_aw_user[2]
port 1198 nsew signal input
rlabel metal3 s 0 19048 800 19168 6 slave_aw_user[3]
port 1199 nsew signal input
rlabel metal3 s 139200 193808 140000 193928 6 slave_aw_user[4]
port 1200 nsew signal input
rlabel metal3 s 0 380808 800 380928 6 slave_aw_user[5]
port 1201 nsew signal input
rlabel metal2 s 18 0 74 800 6 slave_aw_valid
port 1202 nsew signal input
rlabel metal3 s 139200 266568 140000 266688 6 slave_b_id[0]
port 1203 nsew signal output
rlabel metal3 s 0 102008 800 102128 6 slave_b_id[1]
port 1204 nsew signal output
rlabel metal3 s 139200 73448 140000 73568 6 slave_b_id[2]
port 1205 nsew signal output
rlabel metal3 s 139200 116968 140000 117088 6 slave_b_id[3]
port 1206 nsew signal output
rlabel metal2 s 101126 0 101182 800 6 slave_b_id[4]
port 1207 nsew signal output
rlabel metal3 s 0 289688 800 289808 6 slave_b_id[5]
port 1208 nsew signal output
rlabel metal3 s 0 116288 800 116408 6 slave_b_ready
port 1209 nsew signal input
rlabel metal3 s 139200 200608 140000 200728 6 slave_b_resp[0]
port 1210 nsew signal output
rlabel metal3 s 0 297848 800 297968 6 slave_b_resp[1]
port 1211 nsew signal output
rlabel metal2 s 112718 0 112774 800 6 slave_b_user[0]
port 1212 nsew signal output
rlabel metal3 s 0 383528 800 383648 6 slave_b_user[1]
port 1213 nsew signal output
rlabel metal3 s 139200 169328 140000 169448 6 slave_b_user[2]
port 1214 nsew signal output
rlabel metal3 s 139200 381488 140000 381608 6 slave_b_user[3]
port 1215 nsew signal output
rlabel metal3 s 0 306688 800 306808 6 slave_b_user[4]
port 1216 nsew signal output
rlabel metal3 s 0 296488 800 296608 6 slave_b_user[5]
port 1217 nsew signal output
rlabel metal3 s 139200 261808 140000 261928 6 slave_b_valid
port 1218 nsew signal output
rlabel metal3 s 139200 35368 140000 35488 6 slave_r_data[0]
port 1219 nsew signal output
rlabel metal3 s 139200 66648 140000 66768 6 slave_r_data[10]
port 1220 nsew signal output
rlabel metal3 s 0 381488 800 381608 6 slave_r_data[11]
port 1221 nsew signal output
rlabel metal3 s 139200 302608 140000 302728 6 slave_r_data[12]
port 1222 nsew signal output
rlabel metal3 s 0 119008 800 119128 6 slave_r_data[13]
port 1223 nsew signal output
rlabel metal2 s 98550 0 98606 800 6 slave_r_data[14]
port 1224 nsew signal output
rlabel metal2 s 103058 439200 103114 440000 6 slave_r_data[15]
port 1225 nsew signal output
rlabel metal3 s 139200 144848 140000 144968 6 slave_r_data[16]
port 1226 nsew signal output
rlabel metal3 s 0 374008 800 374128 6 slave_r_data[17]
port 1227 nsew signal output
rlabel metal2 s 109498 439200 109554 440000 6 slave_r_data[18]
port 1228 nsew signal output
rlabel metal3 s 0 251608 800 251728 6 slave_r_data[19]
port 1229 nsew signal output
rlabel metal3 s 0 299888 800 300008 6 slave_r_data[1]
port 1230 nsew signal output
rlabel metal3 s 139200 11568 140000 11688 6 slave_r_data[20]
port 1231 nsew signal output
rlabel metal2 s 41878 439200 41934 440000 6 slave_r_data[21]
port 1232 nsew signal output
rlabel metal3 s 139200 140768 140000 140888 6 slave_r_data[22]
port 1233 nsew signal output
rlabel metal2 s 130750 439200 130806 440000 6 slave_r_data[23]
port 1234 nsew signal output
rlabel metal2 s 72790 0 72846 800 6 slave_r_data[24]
port 1235 nsew signal output
rlabel metal3 s 0 232568 800 232688 6 slave_r_data[25]
port 1236 nsew signal output
rlabel metal3 s 139200 80248 140000 80368 6 slave_r_data[26]
port 1237 nsew signal output
rlabel metal3 s 139200 54408 140000 54528 6 slave_r_data[27]
port 1238 nsew signal output
rlabel metal3 s 0 418208 800 418328 6 slave_r_data[28]
port 1239 nsew signal output
rlabel metal3 s 139200 393048 140000 393168 6 slave_r_data[29]
port 1240 nsew signal output
rlabel metal3 s 139200 263848 140000 263968 6 slave_r_data[2]
port 1241 nsew signal output
rlabel metal2 s 122378 439200 122434 440000 6 slave_r_data[30]
port 1242 nsew signal output
rlabel metal3 s 139200 101328 140000 101448 6 slave_r_data[31]
port 1243 nsew signal output
rlabel metal2 s 132038 0 132094 800 6 slave_r_data[32]
port 1244 nsew signal output
rlabel metal3 s 0 261808 800 261928 6 slave_r_data[33]
port 1245 nsew signal output
rlabel metal3 s 0 41488 800 41608 6 slave_r_data[34]
port 1246 nsew signal output
rlabel metal3 s 139200 364488 140000 364608 6 slave_r_data[35]
port 1247 nsew signal output
rlabel metal3 s 139200 419568 140000 419688 6 slave_r_data[36]
port 1248 nsew signal output
rlabel metal3 s 139200 168648 140000 168768 6 slave_r_data[37]
port 1249 nsew signal output
rlabel metal3 s 139200 332528 140000 332648 6 slave_r_data[38]
port 1250 nsew signal output
rlabel metal2 s 86958 439200 87014 440000 6 slave_r_data[39]
port 1251 nsew signal output
rlabel metal3 s 0 268608 800 268728 6 slave_r_data[3]
port 1252 nsew signal output
rlabel metal2 s 29642 0 29698 800 6 slave_r_data[40]
port 1253 nsew signal output
rlabel metal3 s 139200 55768 140000 55888 6 slave_r_data[41]
port 1254 nsew signal output
rlabel metal2 s 103058 0 103114 800 6 slave_r_data[42]
port 1255 nsew signal output
rlabel metal3 s 139200 297848 140000 297968 6 slave_r_data[43]
port 1256 nsew signal output
rlabel metal2 s 23202 0 23258 800 6 slave_r_data[44]
port 1257 nsew signal output
rlabel metal2 s 106278 0 106334 800 6 slave_r_data[45]
port 1258 nsew signal output
rlabel metal3 s 139200 286968 140000 287088 6 slave_r_data[46]
port 1259 nsew signal output
rlabel metal2 s 10966 439200 11022 440000 6 slave_r_data[47]
port 1260 nsew signal output
rlabel metal3 s 139200 384888 140000 385008 6 slave_r_data[48]
port 1261 nsew signal output
rlabel metal2 s 38658 0 38714 800 6 slave_r_data[49]
port 1262 nsew signal output
rlabel metal3 s 139200 355648 140000 355768 6 slave_r_data[4]
port 1263 nsew signal output
rlabel metal3 s 139200 112888 140000 113008 6 slave_r_data[50]
port 1264 nsew signal output
rlabel metal3 s 0 386928 800 387048 6 slave_r_data[51]
port 1265 nsew signal output
rlabel metal3 s 139200 92488 140000 92608 6 slave_r_data[52]
port 1266 nsew signal output
rlabel metal3 s 139200 427048 140000 427168 6 slave_r_data[53]
port 1267 nsew signal output
rlabel metal3 s 0 435208 800 435328 6 slave_r_data[54]
port 1268 nsew signal output
rlabel metal3 s 0 395088 800 395208 6 slave_r_data[55]
port 1269 nsew signal output
rlabel metal3 s 0 303288 800 303408 6 slave_r_data[56]
port 1270 nsew signal output
rlabel metal2 s 2594 439200 2650 440000 6 slave_r_data[57]
port 1271 nsew signal output
rlabel metal3 s 0 175448 800 175568 6 slave_r_data[58]
port 1272 nsew signal output
rlabel metal2 s 115938 0 115994 800 6 slave_r_data[59]
port 1273 nsew signal output
rlabel metal3 s 139200 245488 140000 245608 6 slave_r_data[5]
port 1274 nsew signal output
rlabel metal3 s 139200 338648 140000 338768 6 slave_r_data[60]
port 1275 nsew signal output
rlabel metal3 s 139200 431128 140000 431248 6 slave_r_data[61]
port 1276 nsew signal output
rlabel metal3 s 0 259768 800 259888 6 slave_r_data[62]
port 1277 nsew signal output
rlabel metal3 s 139200 135328 140000 135448 6 slave_r_data[63]
port 1278 nsew signal output
rlabel metal2 s 72146 439200 72202 440000 6 slave_r_data[6]
port 1279 nsew signal output
rlabel metal2 s 117226 439200 117282 440000 6 slave_r_data[7]
port 1280 nsew signal output
rlabel metal3 s 0 419568 800 419688 6 slave_r_data[8]
port 1281 nsew signal output
rlabel metal2 s 43166 439200 43222 440000 6 slave_r_data[9]
port 1282 nsew signal output
rlabel metal3 s 139200 189048 140000 189168 6 slave_r_id[0]
port 1283 nsew signal output
rlabel metal2 s 39302 439200 39358 440000 6 slave_r_id[1]
port 1284 nsew signal output
rlabel metal3 s 139200 174768 140000 174888 6 slave_r_id[2]
port 1285 nsew signal output
rlabel metal3 s 139200 236648 140000 236768 6 slave_r_id[3]
port 1286 nsew signal output
rlabel metal2 s 61842 0 61898 800 6 slave_r_id[4]
port 1287 nsew signal output
rlabel metal2 s 93398 0 93454 800 6 slave_r_id[5]
port 1288 nsew signal output
rlabel metal3 s 139200 196528 140000 196648 6 slave_r_last
port 1289 nsew signal output
rlabel metal3 s 139200 320288 140000 320408 6 slave_r_ready
port 1290 nsew signal input
rlabel metal3 s 0 87728 800 87848 6 slave_r_resp[0]
port 1291 nsew signal output
rlabel metal3 s 0 286968 800 287088 6 slave_r_resp[1]
port 1292 nsew signal output
rlabel metal3 s 0 273368 800 273488 6 slave_r_user[0]
port 1293 nsew signal output
rlabel metal3 s 0 218288 800 218408 6 slave_r_user[1]
port 1294 nsew signal output
rlabel metal2 s 114650 0 114706 800 6 slave_r_user[2]
port 1295 nsew signal output
rlabel metal2 s 50894 439200 50950 440000 6 slave_r_user[3]
port 1296 nsew signal output
rlabel metal3 s 139200 227128 140000 227248 6 slave_r_user[4]
port 1297 nsew signal output
rlabel metal3 s 0 202648 800 202768 6 slave_r_user[5]
port 1298 nsew signal output
rlabel metal2 s 73434 0 73490 800 6 slave_r_valid
port 1299 nsew signal output
rlabel metal2 s 93398 439200 93454 440000 6 slave_w_data[0]
port 1300 nsew signal input
rlabel metal3 s 0 363808 800 363928 6 slave_w_data[10]
port 1301 nsew signal input
rlabel metal3 s 0 74128 800 74248 6 slave_w_data[11]
port 1302 nsew signal input
rlabel metal3 s 0 408008 800 408128 6 slave_w_data[12]
port 1303 nsew signal input
rlabel metal3 s 0 425688 800 425808 6 slave_w_data[13]
port 1304 nsew signal input
rlabel metal3 s 0 429768 800 429888 6 slave_w_data[14]
port 1305 nsew signal input
rlabel metal3 s 0 23128 800 23248 6 slave_w_data[15]
port 1306 nsew signal input
rlabel metal3 s 0 313488 800 313608 6 slave_w_data[16]
port 1307 nsew signal input
rlabel metal3 s 0 18368 800 18488 6 slave_w_data[17]
port 1308 nsew signal input
rlabel metal2 s 5170 0 5226 800 6 slave_w_data[18]
port 1309 nsew signal input
rlabel metal3 s 139200 162528 140000 162648 6 slave_w_data[19]
port 1310 nsew signal input
rlabel metal3 s 0 24488 800 24608 6 slave_w_data[1]
port 1311 nsew signal input
rlabel metal3 s 0 97928 800 98048 6 slave_w_data[20]
port 1312 nsew signal input
rlabel metal3 s 0 355648 800 355768 6 slave_w_data[21]
port 1313 nsew signal input
rlabel metal3 s 139200 301248 140000 301368 6 slave_w_data[22]
port 1314 nsew signal input
rlabel metal3 s 0 125808 800 125928 6 slave_w_data[23]
port 1315 nsew signal input
rlabel metal2 s 14830 0 14886 800 6 slave_w_data[24]
port 1316 nsew signal input
rlabel metal2 s 74722 0 74778 800 6 slave_w_data[25]
port 1317 nsew signal input
rlabel metal3 s 139200 27208 140000 27328 6 slave_w_data[26]
port 1318 nsew signal input
rlabel metal3 s 0 319608 800 319728 6 slave_w_data[27]
port 1319 nsew signal input
rlabel metal3 s 139200 167968 140000 168088 6 slave_w_data[28]
port 1320 nsew signal input
rlabel metal3 s 139200 2048 140000 2168 6 slave_w_data[29]
port 1321 nsew signal input
rlabel metal3 s 139200 146208 140000 146328 6 slave_w_data[2]
port 1322 nsew signal input
rlabel metal3 s 0 99968 800 100088 6 slave_w_data[30]
port 1323 nsew signal input
rlabel metal2 s 81162 439200 81218 440000 6 slave_w_data[31]
port 1324 nsew signal input
rlabel metal3 s 139200 152328 140000 152448 6 slave_w_data[32]
port 1325 nsew signal input
rlabel metal3 s 0 140768 800 140888 6 slave_w_data[33]
port 1326 nsew signal input
rlabel metal3 s 139200 234608 140000 234728 6 slave_w_data[34]
port 1327 nsew signal input
rlabel metal3 s 0 56448 800 56568 6 slave_w_data[35]
port 1328 nsew signal input
rlabel metal3 s 0 40808 800 40928 6 slave_w_data[36]
port 1329 nsew signal input
rlabel metal3 s 139200 431808 140000 431928 6 slave_w_data[37]
port 1330 nsew signal input
rlabel metal3 s 139200 143488 140000 143608 6 slave_w_data[38]
port 1331 nsew signal input
rlabel metal3 s 0 370608 800 370728 6 slave_w_data[39]
port 1332 nsew signal input
rlabel metal3 s 139200 270648 140000 270768 6 slave_w_data[3]
port 1333 nsew signal input
rlabel metal3 s 0 264528 800 264648 6 slave_w_data[40]
port 1334 nsew signal input
rlabel metal3 s 139200 202648 140000 202768 6 slave_w_data[41]
port 1335 nsew signal input
rlabel metal3 s 0 136688 800 136808 6 slave_w_data[42]
port 1336 nsew signal input
rlabel metal2 s 45742 0 45798 800 6 slave_w_data[43]
port 1337 nsew signal input
rlabel metal3 s 139200 414808 140000 414928 6 slave_w_data[44]
port 1338 nsew signal input
rlabel metal3 s 139200 63248 140000 63368 6 slave_w_data[45]
port 1339 nsew signal input
rlabel metal2 s 111430 439200 111486 440000 6 slave_w_data[46]
port 1340 nsew signal input
rlabel metal2 s 90178 0 90234 800 6 slave_w_data[47]
port 1341 nsew signal input
rlabel metal3 s 139200 206048 140000 206168 6 slave_w_data[48]
port 1342 nsew signal input
rlabel metal3 s 0 173408 800 173528 6 slave_w_data[49]
port 1343 nsew signal input
rlabel metal3 s 0 384888 800 385008 6 slave_w_data[4]
port 1344 nsew signal input
rlabel metal2 s 80518 439200 80574 440000 6 slave_w_data[50]
port 1345 nsew signal input
rlabel metal3 s 0 166608 800 166728 6 slave_w_data[51]
port 1346 nsew signal input
rlabel metal3 s 0 200608 800 200728 6 slave_w_data[52]
port 1347 nsew signal input
rlabel metal3 s 0 57808 800 57928 6 slave_w_data[53]
port 1348 nsew signal input
rlabel metal3 s 0 150288 800 150408 6 slave_w_data[54]
port 1349 nsew signal input
rlabel metal3 s 139200 342728 140000 342848 6 slave_w_data[55]
port 1350 nsew signal input
rlabel metal3 s 0 328448 800 328568 6 slave_w_data[56]
port 1351 nsew signal input
rlabel metal3 s 0 255008 800 255128 6 slave_w_data[57]
port 1352 nsew signal input
rlabel metal3 s 0 114928 800 115048 6 slave_w_data[58]
port 1353 nsew signal input
rlabel metal2 s 32218 0 32274 800 6 slave_w_data[59]
port 1354 nsew signal input
rlabel metal3 s 139200 53728 140000 53848 6 slave_w_data[5]
port 1355 nsew signal input
rlabel metal2 s 107566 439200 107622 440000 6 slave_w_data[60]
port 1356 nsew signal input
rlabel metal2 s 128818 439200 128874 440000 6 slave_w_data[61]
port 1357 nsew signal input
rlabel metal3 s 139200 79568 140000 79688 6 slave_w_data[62]
port 1358 nsew signal input
rlabel metal3 s 139200 422968 140000 423088 6 slave_w_data[63]
port 1359 nsew signal input
rlabel metal3 s 139200 319608 140000 319728 6 slave_w_data[6]
port 1360 nsew signal input
rlabel metal3 s 139200 194488 140000 194608 6 slave_w_data[7]
port 1361 nsew signal input
rlabel metal3 s 0 344088 800 344208 6 slave_w_data[8]
port 1362 nsew signal input
rlabel metal2 s 4526 439200 4582 440000 6 slave_w_data[9]
port 1363 nsew signal input
rlabel metal3 s 139200 52368 140000 52488 6 slave_w_last
port 1364 nsew signal input
rlabel metal3 s 139200 137368 140000 137488 6 slave_w_ready
port 1365 nsew signal output
rlabel metal3 s 139200 283568 140000 283688 6 slave_w_strb[0]
port 1366 nsew signal input
rlabel metal3 s 0 170008 800 170128 6 slave_w_strb[1]
port 1367 nsew signal input
rlabel metal3 s 0 51008 800 51128 6 slave_w_strb[2]
port 1368 nsew signal input
rlabel metal2 s 35438 0 35494 800 6 slave_w_strb[3]
port 1369 nsew signal input
rlabel metal3 s 0 252288 800 252408 6 slave_w_strb[4]
port 1370 nsew signal input
rlabel metal3 s 139200 400528 140000 400648 6 slave_w_strb[5]
port 1371 nsew signal input
rlabel metal2 s 56046 439200 56102 440000 6 slave_w_strb[6]
port 1372 nsew signal input
rlabel metal2 s 127530 0 127586 800 6 slave_w_strb[7]
port 1373 nsew signal input
rlabel metal3 s 0 416848 800 416968 6 slave_w_user[0]
port 1374 nsew signal input
rlabel metal3 s 139200 341368 140000 341488 6 slave_w_user[1]
port 1375 nsew signal input
rlabel metal3 s 139200 119688 140000 119808 6 slave_w_user[2]
port 1376 nsew signal input
rlabel metal3 s 0 413448 800 413568 6 slave_w_user[3]
port 1377 nsew signal input
rlabel metal3 s 139200 108808 140000 108928 6 slave_w_user[4]
port 1378 nsew signal input
rlabel metal2 s 102414 0 102470 800 6 slave_w_user[5]
port 1379 nsew signal input
rlabel metal2 s 16762 0 16818 800 6 slave_w_valid
port 1380 nsew signal input
rlabel metal3 s 139200 191768 140000 191888 6 spi_clk_i
port 1381 nsew signal input
rlabel metal3 s 139200 282208 140000 282328 6 spi_cs_i
port 1382 nsew signal input
rlabel metal3 s 0 270648 800 270768 6 spi_master_clk
port 1383 nsew signal output
rlabel metal2 s 99838 439200 99894 440000 6 spi_master_csn0
port 1384 nsew signal output
rlabel metal3 s 0 93848 800 93968 6 spi_master_csn1
port 1385 nsew signal output
rlabel metal3 s 0 119688 800 119808 6 spi_master_csn2
port 1386 nsew signal output
rlabel metal3 s 0 110848 800 110968 6 spi_master_csn3
port 1387 nsew signal output
rlabel metal2 s 13542 0 13598 800 6 spi_master_mode[0]
port 1388 nsew signal output
rlabel metal2 s 68926 0 68982 800 6 spi_master_mode[1]
port 1389 nsew signal output
rlabel metal3 s 139200 358368 140000 358488 6 spi_master_sdi0
port 1390 nsew signal input
rlabel metal3 s 139200 43528 140000 43648 6 spi_master_sdi1
port 1391 nsew signal input
rlabel metal3 s 0 410048 800 410168 6 spi_master_sdi2
port 1392 nsew signal input
rlabel metal2 s 48318 439200 48374 440000 6 spi_master_sdi3
port 1393 nsew signal input
rlabel metal3 s 0 206048 800 206168 6 spi_master_sdo0
port 1394 nsew signal output
rlabel metal2 s 48962 0 49018 800 6 spi_master_sdo1
port 1395 nsew signal output
rlabel metal3 s 139200 378768 140000 378888 6 spi_master_sdo2
port 1396 nsew signal output
rlabel metal2 s 63130 439200 63186 440000 6 spi_master_sdo3
port 1397 nsew signal output
rlabel metal3 s 0 63928 800 64048 6 spi_mode_o[0]
port 1398 nsew signal output
rlabel metal3 s 139200 433848 140000 433968 6 spi_mode_o[1]
port 1399 nsew signal output
rlabel metal3 s 139200 284248 140000 284368 6 spi_sdi0_i
port 1400 nsew signal input
rlabel metal3 s 139200 77528 140000 77648 6 spi_sdi1_i
port 1401 nsew signal input
rlabel metal3 s 0 5448 800 5568 6 spi_sdi2_i
port 1402 nsew signal input
rlabel metal3 s 0 284928 800 285048 6 spi_sdi3_i
port 1403 nsew signal input
rlabel metal2 s 97262 0 97318 800 6 spi_sdo0_o
port 1404 nsew signal output
rlabel metal3 s 139200 369928 140000 370048 6 spi_sdo1_o
port 1405 nsew signal output
rlabel metal3 s 139200 116288 140000 116408 6 spi_sdo2_o
port 1406 nsew signal output
rlabel metal3 s 139200 268608 140000 268728 6 spi_sdo3_o
port 1407 nsew signal output
rlabel metal3 s 0 65968 800 66088 6 testmode_i
port 1408 nsew signal input
rlabel metal3 s 139200 184288 140000 184408 6 testmode_i_pll
port 1409 nsew signal input
rlabel metal2 s 49606 0 49662 800 6 uart_cts
port 1410 nsew signal input
rlabel metal3 s 139200 10208 140000 10328 6 uart_dsr
port 1411 nsew signal input
rlabel metal3 s 139200 308048 140000 308168 6 uart_dtr
port 1412 nsew signal output
rlabel metal2 s 34794 439200 34850 440000 6 uart_rts
port 1413 nsew signal output
rlabel metal2 s 128174 439200 128230 440000 6 uart_rx
port 1414 nsew signal input
rlabel metal3 s 139200 184968 140000 185088 6 uart_tx
port 1415 nsew signal output
rlabel metal2 s 24490 0 24546 800 6 user_irq_pll[0]
port 1416 nsew signal output
rlabel metal3 s 139200 346808 140000 346928 6 user_irq_pll[1]
port 1417 nsew signal output
rlabel metal2 s 7102 0 7158 800 6 user_irq_pll[2]
port 1418 nsew signal output
rlabel metal2 s 126886 439200 126942 440000 6 vccd1
port 1419 nsew signal bidirectional
rlabel metal4 s 4208 2128 4528 437424 6 vccd1
port 1419 nsew signal bidirectional
rlabel metal4 s 34928 2128 35248 437424 6 vccd1
port 1419 nsew signal bidirectional
rlabel metal4 s 65648 2128 65968 437424 6 vccd1
port 1419 nsew signal bidirectional
rlabel metal4 s 96368 2128 96688 437424 6 vccd1
port 1419 nsew signal bidirectional
rlabel metal4 s 127088 2128 127408 437424 6 vccd1
port 1419 nsew signal bidirectional
rlabel metal2 s 31574 439200 31630 440000 6 vssd1
port 1420 nsew signal bidirectional
rlabel metal4 s 19568 2128 19888 437424 6 vssd1
port 1420 nsew signal bidirectional
rlabel metal4 s 50288 2128 50608 437424 6 vssd1
port 1420 nsew signal bidirectional
rlabel metal4 s 81008 2128 81328 437424 6 vssd1
port 1420 nsew signal bidirectional
rlabel metal4 s 111728 2128 112048 437424 6 vssd1
port 1420 nsew signal bidirectional
rlabel metal3 s 139200 201288 140000 201408 6 wbs_ack_o_pll
port 1421 nsew signal output
rlabel metal2 s 23846 439200 23902 440000 6 wbs_dat_o_pll[0]
port 1422 nsew signal output
rlabel metal3 s 139200 61888 140000 62008 6 wbs_dat_o_pll[10]
port 1423 nsew signal output
rlabel metal3 s 0 32648 800 32768 6 wbs_dat_o_pll[11]
port 1424 nsew signal output
rlabel metal3 s 139200 61208 140000 61328 6 wbs_dat_o_pll[12]
port 1425 nsew signal output
rlabel metal2 s 662 0 718 800 6 wbs_dat_o_pll[13]
port 1426 nsew signal output
rlabel metal3 s 139200 96568 140000 96688 6 wbs_dat_o_pll[14]
port 1427 nsew signal output
rlabel metal3 s 0 91128 800 91248 6 wbs_dat_o_pll[15]
port 1428 nsew signal output
rlabel metal3 s 0 213528 800 213648 6 wbs_dat_o_pll[16]
port 1429 nsew signal output
rlabel metal3 s 0 340688 800 340808 6 wbs_dat_o_pll[17]
port 1430 nsew signal output
rlabel metal3 s 0 53048 800 53168 6 wbs_dat_o_pll[18]
port 1431 nsew signal output
rlabel metal2 s 61198 0 61254 800 6 wbs_dat_o_pll[19]
port 1432 nsew signal output
rlabel metal2 s 21914 0 21970 800 6 wbs_dat_o_pll[1]
port 1433 nsew signal output
rlabel metal3 s 0 420928 800 421048 6 wbs_dat_o_pll[20]
port 1434 nsew signal output
rlabel metal3 s 0 353608 800 353728 6 wbs_dat_o_pll[21]
port 1435 nsew signal output
rlabel metal3 s 139200 17688 140000 17808 6 wbs_dat_o_pll[22]
port 1436 nsew signal output
rlabel metal3 s 0 6128 800 6248 6 wbs_dat_o_pll[23]
port 1437 nsew signal output
rlabel metal3 s 139200 239368 140000 239488 6 wbs_dat_o_pll[24]
port 1438 nsew signal output
rlabel metal3 s 0 167288 800 167408 6 wbs_dat_o_pll[25]
port 1439 nsew signal output
rlabel metal3 s 139200 386928 140000 387048 6 wbs_dat_o_pll[26]
port 1440 nsew signal output
rlabel metal2 s 63130 0 63186 800 6 wbs_dat_o_pll[27]
port 1441 nsew signal output
rlabel metal2 s 110142 0 110198 800 6 wbs_dat_o_pll[28]
port 1442 nsew signal output
rlabel metal3 s 0 6808 800 6928 6 wbs_dat_o_pll[29]
port 1443 nsew signal output
rlabel metal3 s 139200 371968 140000 372088 6 wbs_dat_o_pll[2]
port 1444 nsew signal output
rlabel metal3 s 139200 33328 140000 33448 6 wbs_dat_o_pll[30]
port 1445 nsew signal output
rlabel metal2 s 35438 439200 35494 440000 6 wbs_dat_o_pll[31]
port 1446 nsew signal output
rlabel metal2 s 32862 439200 32918 440000 6 wbs_dat_o_pll[3]
port 1447 nsew signal output
rlabel metal3 s 0 262488 800 262608 6 wbs_dat_o_pll[4]
port 1448 nsew signal output
rlabel metal3 s 0 317568 800 317688 6 wbs_dat_o_pll[5]
port 1449 nsew signal output
rlabel metal3 s 139200 65968 140000 66088 6 wbs_dat_o_pll[6]
port 1450 nsew signal output
rlabel metal3 s 0 59848 800 59968 6 wbs_dat_o_pll[7]
port 1451 nsew signal output
rlabel metal3 s 0 240048 800 240168 6 wbs_dat_o_pll[8]
port 1452 nsew signal output
rlabel metal3 s 139200 291728 140000 291848 6 wbs_dat_o_pll[9]
port 1453 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 140000 440000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 83802832
string GDS_FILE /home/mbaykenar/Desktop/workspace/mpw7_yonga_soc/openlane/peripherals_2/runs/22_09_07_17_47/results/signoff/peripherals.magic.gds
string GDS_START 1773840
<< end >>

