magic
tech sky130A
magscale 1 2
timestamp 1649977179
<< metal3 >>
rect 194 9244 4879 9246
rect 194 9180 200 9244
rect 264 9180 281 9244
rect 345 9180 362 9244
rect 426 9180 443 9244
rect 507 9180 524 9244
rect 588 9180 605 9244
rect 669 9180 686 9244
rect 750 9180 767 9244
rect 831 9180 848 9244
rect 912 9180 929 9244
rect 993 9180 1010 9244
rect 1074 9180 1091 9244
rect 1155 9180 1172 9244
rect 1236 9180 1253 9244
rect 1317 9180 1334 9244
rect 1398 9180 1415 9244
rect 1479 9180 1496 9244
rect 1560 9180 1577 9244
rect 1641 9180 1658 9244
rect 1722 9180 1739 9244
rect 1803 9180 1820 9244
rect 1884 9180 1901 9244
rect 1965 9180 1982 9244
rect 2046 9180 2063 9244
rect 2127 9180 2144 9244
rect 2208 9180 2225 9244
rect 2289 9180 2306 9244
rect 2370 9180 2387 9244
rect 2451 9180 2468 9244
rect 2532 9180 2549 9244
rect 2613 9180 2630 9244
rect 2694 9180 2711 9244
rect 2775 9180 2792 9244
rect 2856 9180 2873 9244
rect 2937 9180 2954 9244
rect 3018 9180 3035 9244
rect 3099 9180 3116 9244
rect 3180 9180 3197 9244
rect 3261 9180 3278 9244
rect 3342 9180 3359 9244
rect 3423 9180 3440 9244
rect 3504 9180 3521 9244
rect 3585 9180 3602 9244
rect 3666 9180 3683 9244
rect 3747 9180 3764 9244
rect 3828 9180 3845 9244
rect 3909 9180 3926 9244
rect 3990 9180 4007 9244
rect 4071 9180 4088 9244
rect 4152 9180 4169 9244
rect 4233 9180 4249 9244
rect 4313 9180 4329 9244
rect 4393 9180 4409 9244
rect 4473 9180 4489 9244
rect 4553 9180 4569 9244
rect 4633 9180 4649 9244
rect 4713 9180 4729 9244
rect 4793 9180 4809 9244
rect 4873 9180 4879 9244
rect 194 9158 4879 9180
rect 194 9094 200 9158
rect 264 9094 281 9158
rect 345 9094 362 9158
rect 426 9094 443 9158
rect 507 9094 524 9158
rect 588 9094 605 9158
rect 669 9094 686 9158
rect 750 9094 767 9158
rect 831 9094 848 9158
rect 912 9094 929 9158
rect 993 9094 1010 9158
rect 1074 9094 1091 9158
rect 1155 9094 1172 9158
rect 1236 9094 1253 9158
rect 1317 9094 1334 9158
rect 1398 9094 1415 9158
rect 1479 9094 1496 9158
rect 1560 9094 1577 9158
rect 1641 9094 1658 9158
rect 1722 9094 1739 9158
rect 1803 9094 1820 9158
rect 1884 9094 1901 9158
rect 1965 9094 1982 9158
rect 2046 9094 2063 9158
rect 2127 9094 2144 9158
rect 2208 9094 2225 9158
rect 2289 9094 2306 9158
rect 2370 9094 2387 9158
rect 2451 9094 2468 9158
rect 2532 9094 2549 9158
rect 2613 9094 2630 9158
rect 2694 9094 2711 9158
rect 2775 9094 2792 9158
rect 2856 9094 2873 9158
rect 2937 9094 2954 9158
rect 3018 9094 3035 9158
rect 3099 9094 3116 9158
rect 3180 9094 3197 9158
rect 3261 9094 3278 9158
rect 3342 9094 3359 9158
rect 3423 9094 3440 9158
rect 3504 9094 3521 9158
rect 3585 9094 3602 9158
rect 3666 9094 3683 9158
rect 3747 9094 3764 9158
rect 3828 9094 3845 9158
rect 3909 9094 3926 9158
rect 3990 9094 4007 9158
rect 4071 9094 4088 9158
rect 4152 9094 4169 9158
rect 4233 9094 4249 9158
rect 4313 9094 4329 9158
rect 4393 9094 4409 9158
rect 4473 9094 4489 9158
rect 4553 9094 4569 9158
rect 4633 9094 4649 9158
rect 4713 9094 4729 9158
rect 4793 9094 4809 9158
rect 4873 9094 4879 9158
rect 194 9072 4879 9094
rect 194 9008 200 9072
rect 264 9008 281 9072
rect 345 9008 362 9072
rect 426 9008 443 9072
rect 507 9008 524 9072
rect 588 9008 605 9072
rect 669 9008 686 9072
rect 750 9008 767 9072
rect 831 9008 848 9072
rect 912 9008 929 9072
rect 993 9008 1010 9072
rect 1074 9008 1091 9072
rect 1155 9008 1172 9072
rect 1236 9008 1253 9072
rect 1317 9008 1334 9072
rect 1398 9008 1415 9072
rect 1479 9008 1496 9072
rect 1560 9008 1577 9072
rect 1641 9008 1658 9072
rect 1722 9008 1739 9072
rect 1803 9008 1820 9072
rect 1884 9008 1901 9072
rect 1965 9008 1982 9072
rect 2046 9008 2063 9072
rect 2127 9008 2144 9072
rect 2208 9008 2225 9072
rect 2289 9008 2306 9072
rect 2370 9008 2387 9072
rect 2451 9008 2468 9072
rect 2532 9008 2549 9072
rect 2613 9008 2630 9072
rect 2694 9008 2711 9072
rect 2775 9008 2792 9072
rect 2856 9008 2873 9072
rect 2937 9008 2954 9072
rect 3018 9008 3035 9072
rect 3099 9008 3116 9072
rect 3180 9008 3197 9072
rect 3261 9008 3278 9072
rect 3342 9008 3359 9072
rect 3423 9008 3440 9072
rect 3504 9008 3521 9072
rect 3585 9008 3602 9072
rect 3666 9008 3683 9072
rect 3747 9008 3764 9072
rect 3828 9008 3845 9072
rect 3909 9008 3926 9072
rect 3990 9008 4007 9072
rect 4071 9008 4088 9072
rect 4152 9008 4169 9072
rect 4233 9008 4249 9072
rect 4313 9008 4329 9072
rect 4393 9008 4409 9072
rect 4473 9008 4489 9072
rect 4553 9008 4569 9072
rect 4633 9008 4649 9072
rect 4713 9008 4729 9072
rect 4793 9008 4809 9072
rect 4873 9008 4879 9072
rect 194 8986 4879 9008
rect 194 8922 200 8986
rect 264 8922 281 8986
rect 345 8922 362 8986
rect 426 8922 443 8986
rect 507 8922 524 8986
rect 588 8922 605 8986
rect 669 8922 686 8986
rect 750 8922 767 8986
rect 831 8922 848 8986
rect 912 8922 929 8986
rect 993 8922 1010 8986
rect 1074 8922 1091 8986
rect 1155 8922 1172 8986
rect 1236 8922 1253 8986
rect 1317 8922 1334 8986
rect 1398 8922 1415 8986
rect 1479 8922 1496 8986
rect 1560 8922 1577 8986
rect 1641 8922 1658 8986
rect 1722 8922 1739 8986
rect 1803 8922 1820 8986
rect 1884 8922 1901 8986
rect 1965 8922 1982 8986
rect 2046 8922 2063 8986
rect 2127 8922 2144 8986
rect 2208 8922 2225 8986
rect 2289 8922 2306 8986
rect 2370 8922 2387 8986
rect 2451 8922 2468 8986
rect 2532 8922 2549 8986
rect 2613 8922 2630 8986
rect 2694 8922 2711 8986
rect 2775 8922 2792 8986
rect 2856 8922 2873 8986
rect 2937 8922 2954 8986
rect 3018 8922 3035 8986
rect 3099 8922 3116 8986
rect 3180 8922 3197 8986
rect 3261 8922 3278 8986
rect 3342 8922 3359 8986
rect 3423 8922 3440 8986
rect 3504 8922 3521 8986
rect 3585 8922 3602 8986
rect 3666 8922 3683 8986
rect 3747 8922 3764 8986
rect 3828 8922 3845 8986
rect 3909 8922 3926 8986
rect 3990 8922 4007 8986
rect 4071 8922 4088 8986
rect 4152 8922 4169 8986
rect 4233 8922 4249 8986
rect 4313 8922 4329 8986
rect 4393 8922 4409 8986
rect 4473 8922 4489 8986
rect 4553 8922 4569 8986
rect 4633 8922 4649 8986
rect 4713 8922 4729 8986
rect 4793 8922 4809 8986
rect 4873 8922 4879 8986
rect 194 8900 4879 8922
rect 194 8836 200 8900
rect 264 8836 281 8900
rect 345 8836 362 8900
rect 426 8836 443 8900
rect 507 8836 524 8900
rect 588 8836 605 8900
rect 669 8836 686 8900
rect 750 8836 767 8900
rect 831 8836 848 8900
rect 912 8836 929 8900
rect 993 8836 1010 8900
rect 1074 8836 1091 8900
rect 1155 8836 1172 8900
rect 1236 8836 1253 8900
rect 1317 8836 1334 8900
rect 1398 8836 1415 8900
rect 1479 8836 1496 8900
rect 1560 8836 1577 8900
rect 1641 8836 1658 8900
rect 1722 8836 1739 8900
rect 1803 8836 1820 8900
rect 1884 8836 1901 8900
rect 1965 8836 1982 8900
rect 2046 8836 2063 8900
rect 2127 8836 2144 8900
rect 2208 8836 2225 8900
rect 2289 8836 2306 8900
rect 2370 8836 2387 8900
rect 2451 8836 2468 8900
rect 2532 8836 2549 8900
rect 2613 8836 2630 8900
rect 2694 8836 2711 8900
rect 2775 8836 2792 8900
rect 2856 8836 2873 8900
rect 2937 8836 2954 8900
rect 3018 8836 3035 8900
rect 3099 8836 3116 8900
rect 3180 8836 3197 8900
rect 3261 8836 3278 8900
rect 3342 8836 3359 8900
rect 3423 8836 3440 8900
rect 3504 8836 3521 8900
rect 3585 8836 3602 8900
rect 3666 8836 3683 8900
rect 3747 8836 3764 8900
rect 3828 8836 3845 8900
rect 3909 8836 3926 8900
rect 3990 8836 4007 8900
rect 4071 8836 4088 8900
rect 4152 8836 4169 8900
rect 4233 8836 4249 8900
rect 4313 8836 4329 8900
rect 4393 8836 4409 8900
rect 4473 8836 4489 8900
rect 4553 8836 4569 8900
rect 4633 8836 4649 8900
rect 4713 8836 4729 8900
rect 4793 8836 4809 8900
rect 4873 8836 4879 8900
rect 194 8814 4879 8836
rect 194 8750 200 8814
rect 264 8750 281 8814
rect 345 8750 362 8814
rect 426 8750 443 8814
rect 507 8750 524 8814
rect 588 8750 605 8814
rect 669 8750 686 8814
rect 750 8750 767 8814
rect 831 8750 848 8814
rect 912 8750 929 8814
rect 993 8750 1010 8814
rect 1074 8750 1091 8814
rect 1155 8750 1172 8814
rect 1236 8750 1253 8814
rect 1317 8750 1334 8814
rect 1398 8750 1415 8814
rect 1479 8750 1496 8814
rect 1560 8750 1577 8814
rect 1641 8750 1658 8814
rect 1722 8750 1739 8814
rect 1803 8750 1820 8814
rect 1884 8750 1901 8814
rect 1965 8750 1982 8814
rect 2046 8750 2063 8814
rect 2127 8750 2144 8814
rect 2208 8750 2225 8814
rect 2289 8750 2306 8814
rect 2370 8750 2387 8814
rect 2451 8750 2468 8814
rect 2532 8750 2549 8814
rect 2613 8750 2630 8814
rect 2694 8750 2711 8814
rect 2775 8750 2792 8814
rect 2856 8750 2873 8814
rect 2937 8750 2954 8814
rect 3018 8750 3035 8814
rect 3099 8750 3116 8814
rect 3180 8750 3197 8814
rect 3261 8750 3278 8814
rect 3342 8750 3359 8814
rect 3423 8750 3440 8814
rect 3504 8750 3521 8814
rect 3585 8750 3602 8814
rect 3666 8750 3683 8814
rect 3747 8750 3764 8814
rect 3828 8750 3845 8814
rect 3909 8750 3926 8814
rect 3990 8750 4007 8814
rect 4071 8750 4088 8814
rect 4152 8750 4169 8814
rect 4233 8750 4249 8814
rect 4313 8750 4329 8814
rect 4393 8750 4409 8814
rect 4473 8750 4489 8814
rect 4553 8750 4569 8814
rect 4633 8750 4649 8814
rect 4713 8750 4729 8814
rect 4793 8750 4809 8814
rect 4873 8750 4879 8814
rect 194 8728 4879 8750
rect 194 8664 200 8728
rect 264 8664 281 8728
rect 345 8664 362 8728
rect 426 8664 443 8728
rect 507 8664 524 8728
rect 588 8664 605 8728
rect 669 8664 686 8728
rect 750 8664 767 8728
rect 831 8664 848 8728
rect 912 8664 929 8728
rect 993 8664 1010 8728
rect 1074 8664 1091 8728
rect 1155 8664 1172 8728
rect 1236 8664 1253 8728
rect 1317 8664 1334 8728
rect 1398 8664 1415 8728
rect 1479 8664 1496 8728
rect 1560 8664 1577 8728
rect 1641 8664 1658 8728
rect 1722 8664 1739 8728
rect 1803 8664 1820 8728
rect 1884 8664 1901 8728
rect 1965 8664 1982 8728
rect 2046 8664 2063 8728
rect 2127 8664 2144 8728
rect 2208 8664 2225 8728
rect 2289 8664 2306 8728
rect 2370 8664 2387 8728
rect 2451 8664 2468 8728
rect 2532 8664 2549 8728
rect 2613 8664 2630 8728
rect 2694 8664 2711 8728
rect 2775 8664 2792 8728
rect 2856 8664 2873 8728
rect 2937 8664 2954 8728
rect 3018 8664 3035 8728
rect 3099 8664 3116 8728
rect 3180 8664 3197 8728
rect 3261 8664 3278 8728
rect 3342 8664 3359 8728
rect 3423 8664 3440 8728
rect 3504 8664 3521 8728
rect 3585 8664 3602 8728
rect 3666 8664 3683 8728
rect 3747 8664 3764 8728
rect 3828 8664 3845 8728
rect 3909 8664 3926 8728
rect 3990 8664 4007 8728
rect 4071 8664 4088 8728
rect 4152 8664 4169 8728
rect 4233 8664 4249 8728
rect 4313 8664 4329 8728
rect 4393 8664 4409 8728
rect 4473 8664 4489 8728
rect 4553 8664 4569 8728
rect 4633 8664 4649 8728
rect 4713 8664 4729 8728
rect 4793 8664 4809 8728
rect 4873 8664 4879 8728
rect 194 8642 4879 8664
rect 194 8578 200 8642
rect 264 8578 281 8642
rect 345 8578 362 8642
rect 426 8578 443 8642
rect 507 8578 524 8642
rect 588 8578 605 8642
rect 669 8578 686 8642
rect 750 8578 767 8642
rect 831 8578 848 8642
rect 912 8578 929 8642
rect 993 8578 1010 8642
rect 1074 8578 1091 8642
rect 1155 8578 1172 8642
rect 1236 8578 1253 8642
rect 1317 8578 1334 8642
rect 1398 8578 1415 8642
rect 1479 8578 1496 8642
rect 1560 8578 1577 8642
rect 1641 8578 1658 8642
rect 1722 8578 1739 8642
rect 1803 8578 1820 8642
rect 1884 8578 1901 8642
rect 1965 8578 1982 8642
rect 2046 8578 2063 8642
rect 2127 8578 2144 8642
rect 2208 8578 2225 8642
rect 2289 8578 2306 8642
rect 2370 8578 2387 8642
rect 2451 8578 2468 8642
rect 2532 8578 2549 8642
rect 2613 8578 2630 8642
rect 2694 8578 2711 8642
rect 2775 8578 2792 8642
rect 2856 8578 2873 8642
rect 2937 8578 2954 8642
rect 3018 8578 3035 8642
rect 3099 8578 3116 8642
rect 3180 8578 3197 8642
rect 3261 8578 3278 8642
rect 3342 8578 3359 8642
rect 3423 8578 3440 8642
rect 3504 8578 3521 8642
rect 3585 8578 3602 8642
rect 3666 8578 3683 8642
rect 3747 8578 3764 8642
rect 3828 8578 3845 8642
rect 3909 8578 3926 8642
rect 3990 8578 4007 8642
rect 4071 8578 4088 8642
rect 4152 8578 4169 8642
rect 4233 8578 4249 8642
rect 4313 8578 4329 8642
rect 4393 8578 4409 8642
rect 4473 8578 4489 8642
rect 4553 8578 4569 8642
rect 4633 8578 4649 8642
rect 4713 8578 4729 8642
rect 4793 8578 4809 8642
rect 4873 8578 4879 8642
rect 194 8556 4879 8578
rect 194 8492 200 8556
rect 264 8492 281 8556
rect 345 8492 362 8556
rect 426 8492 443 8556
rect 507 8492 524 8556
rect 588 8492 605 8556
rect 669 8492 686 8556
rect 750 8492 767 8556
rect 831 8492 848 8556
rect 912 8492 929 8556
rect 993 8492 1010 8556
rect 1074 8492 1091 8556
rect 1155 8492 1172 8556
rect 1236 8492 1253 8556
rect 1317 8492 1334 8556
rect 1398 8492 1415 8556
rect 1479 8492 1496 8556
rect 1560 8492 1577 8556
rect 1641 8492 1658 8556
rect 1722 8492 1739 8556
rect 1803 8492 1820 8556
rect 1884 8492 1901 8556
rect 1965 8492 1982 8556
rect 2046 8492 2063 8556
rect 2127 8492 2144 8556
rect 2208 8492 2225 8556
rect 2289 8492 2306 8556
rect 2370 8492 2387 8556
rect 2451 8492 2468 8556
rect 2532 8492 2549 8556
rect 2613 8492 2630 8556
rect 2694 8492 2711 8556
rect 2775 8492 2792 8556
rect 2856 8492 2873 8556
rect 2937 8492 2954 8556
rect 3018 8492 3035 8556
rect 3099 8492 3116 8556
rect 3180 8492 3197 8556
rect 3261 8492 3278 8556
rect 3342 8492 3359 8556
rect 3423 8492 3440 8556
rect 3504 8492 3521 8556
rect 3585 8492 3602 8556
rect 3666 8492 3683 8556
rect 3747 8492 3764 8556
rect 3828 8492 3845 8556
rect 3909 8492 3926 8556
rect 3990 8492 4007 8556
rect 4071 8492 4088 8556
rect 4152 8492 4169 8556
rect 4233 8492 4249 8556
rect 4313 8492 4329 8556
rect 4393 8492 4409 8556
rect 4473 8492 4489 8556
rect 4553 8492 4569 8556
rect 4633 8492 4649 8556
rect 4713 8492 4729 8556
rect 4793 8492 4809 8556
rect 4873 8492 4879 8556
rect 194 8470 4879 8492
rect 194 8406 200 8470
rect 264 8406 281 8470
rect 345 8406 362 8470
rect 426 8406 443 8470
rect 507 8406 524 8470
rect 588 8406 605 8470
rect 669 8406 686 8470
rect 750 8406 767 8470
rect 831 8406 848 8470
rect 912 8406 929 8470
rect 993 8406 1010 8470
rect 1074 8406 1091 8470
rect 1155 8406 1172 8470
rect 1236 8406 1253 8470
rect 1317 8406 1334 8470
rect 1398 8406 1415 8470
rect 1479 8406 1496 8470
rect 1560 8406 1577 8470
rect 1641 8406 1658 8470
rect 1722 8406 1739 8470
rect 1803 8406 1820 8470
rect 1884 8406 1901 8470
rect 1965 8406 1982 8470
rect 2046 8406 2063 8470
rect 2127 8406 2144 8470
rect 2208 8406 2225 8470
rect 2289 8406 2306 8470
rect 2370 8406 2387 8470
rect 2451 8406 2468 8470
rect 2532 8406 2549 8470
rect 2613 8406 2630 8470
rect 2694 8406 2711 8470
rect 2775 8406 2792 8470
rect 2856 8406 2873 8470
rect 2937 8406 2954 8470
rect 3018 8406 3035 8470
rect 3099 8406 3116 8470
rect 3180 8406 3197 8470
rect 3261 8406 3278 8470
rect 3342 8406 3359 8470
rect 3423 8406 3440 8470
rect 3504 8406 3521 8470
rect 3585 8406 3602 8470
rect 3666 8406 3683 8470
rect 3747 8406 3764 8470
rect 3828 8406 3845 8470
rect 3909 8406 3926 8470
rect 3990 8406 4007 8470
rect 4071 8406 4088 8470
rect 4152 8406 4169 8470
rect 4233 8406 4249 8470
rect 4313 8406 4329 8470
rect 4393 8406 4409 8470
rect 4473 8406 4489 8470
rect 4553 8406 4569 8470
rect 4633 8406 4649 8470
rect 4713 8406 4729 8470
rect 4793 8406 4809 8470
rect 4873 8406 4879 8470
rect 194 8384 4879 8406
rect 194 8320 200 8384
rect 264 8320 281 8384
rect 345 8320 362 8384
rect 426 8320 443 8384
rect 507 8320 524 8384
rect 588 8320 605 8384
rect 669 8320 686 8384
rect 750 8320 767 8384
rect 831 8320 848 8384
rect 912 8320 929 8384
rect 993 8320 1010 8384
rect 1074 8320 1091 8384
rect 1155 8320 1172 8384
rect 1236 8320 1253 8384
rect 1317 8320 1334 8384
rect 1398 8320 1415 8384
rect 1479 8320 1496 8384
rect 1560 8320 1577 8384
rect 1641 8320 1658 8384
rect 1722 8320 1739 8384
rect 1803 8320 1820 8384
rect 1884 8320 1901 8384
rect 1965 8320 1982 8384
rect 2046 8320 2063 8384
rect 2127 8320 2144 8384
rect 2208 8320 2225 8384
rect 2289 8320 2306 8384
rect 2370 8320 2387 8384
rect 2451 8320 2468 8384
rect 2532 8320 2549 8384
rect 2613 8320 2630 8384
rect 2694 8320 2711 8384
rect 2775 8320 2792 8384
rect 2856 8320 2873 8384
rect 2937 8320 2954 8384
rect 3018 8320 3035 8384
rect 3099 8320 3116 8384
rect 3180 8320 3197 8384
rect 3261 8320 3278 8384
rect 3342 8320 3359 8384
rect 3423 8320 3440 8384
rect 3504 8320 3521 8384
rect 3585 8320 3602 8384
rect 3666 8320 3683 8384
rect 3747 8320 3764 8384
rect 3828 8320 3845 8384
rect 3909 8320 3926 8384
rect 3990 8320 4007 8384
rect 4071 8320 4088 8384
rect 4152 8320 4169 8384
rect 4233 8320 4249 8384
rect 4313 8320 4329 8384
rect 4393 8320 4409 8384
rect 4473 8320 4489 8384
rect 4553 8320 4569 8384
rect 4633 8320 4649 8384
rect 4713 8320 4729 8384
rect 4793 8320 4809 8384
rect 4873 8320 4879 8384
rect 194 8318 4879 8320
rect 10078 9244 14858 9246
rect 10078 9180 10084 9244
rect 10148 9180 10166 9244
rect 10230 9180 10248 9244
rect 10312 9180 10330 9244
rect 10394 9180 10412 9244
rect 10476 9180 10494 9244
rect 10558 9180 10576 9244
rect 10640 9180 10657 9244
rect 10721 9180 10738 9244
rect 10802 9180 10819 9244
rect 10883 9180 10900 9244
rect 10964 9180 10981 9244
rect 11045 9180 11062 9244
rect 11126 9180 11143 9244
rect 11207 9180 11224 9244
rect 11288 9180 11305 9244
rect 11369 9180 11386 9244
rect 11450 9180 11467 9244
rect 11531 9180 11548 9244
rect 11612 9180 11629 9244
rect 11693 9180 11710 9244
rect 11774 9180 11791 9244
rect 11855 9180 11872 9244
rect 11936 9180 11953 9244
rect 12017 9180 12034 9244
rect 12098 9180 12115 9244
rect 12179 9180 12196 9244
rect 12260 9180 12277 9244
rect 12341 9180 12358 9244
rect 12422 9180 12439 9244
rect 12503 9180 12520 9244
rect 12584 9180 12601 9244
rect 12665 9180 12682 9244
rect 12746 9180 12763 9244
rect 12827 9180 12844 9244
rect 12908 9180 12925 9244
rect 12989 9180 13006 9244
rect 13070 9180 13087 9244
rect 13151 9180 13168 9244
rect 13232 9180 13249 9244
rect 13313 9180 13330 9244
rect 13394 9180 13411 9244
rect 13475 9180 13492 9244
rect 13556 9180 13573 9244
rect 13637 9180 13654 9244
rect 13718 9180 13735 9244
rect 13799 9180 13816 9244
rect 13880 9180 13897 9244
rect 13961 9180 13978 9244
rect 14042 9180 14059 9244
rect 14123 9180 14140 9244
rect 14204 9180 14221 9244
rect 14285 9180 14302 9244
rect 14366 9180 14383 9244
rect 14447 9180 14464 9244
rect 14528 9180 14545 9244
rect 14609 9180 14626 9244
rect 14690 9180 14707 9244
rect 14771 9180 14788 9244
rect 14852 9180 14858 9244
rect 10078 9158 14858 9180
rect 10078 9094 10084 9158
rect 10148 9094 10166 9158
rect 10230 9094 10248 9158
rect 10312 9094 10330 9158
rect 10394 9094 10412 9158
rect 10476 9094 10494 9158
rect 10558 9094 10576 9158
rect 10640 9094 10657 9158
rect 10721 9094 10738 9158
rect 10802 9094 10819 9158
rect 10883 9094 10900 9158
rect 10964 9094 10981 9158
rect 11045 9094 11062 9158
rect 11126 9094 11143 9158
rect 11207 9094 11224 9158
rect 11288 9094 11305 9158
rect 11369 9094 11386 9158
rect 11450 9094 11467 9158
rect 11531 9094 11548 9158
rect 11612 9094 11629 9158
rect 11693 9094 11710 9158
rect 11774 9094 11791 9158
rect 11855 9094 11872 9158
rect 11936 9094 11953 9158
rect 12017 9094 12034 9158
rect 12098 9094 12115 9158
rect 12179 9094 12196 9158
rect 12260 9094 12277 9158
rect 12341 9094 12358 9158
rect 12422 9094 12439 9158
rect 12503 9094 12520 9158
rect 12584 9094 12601 9158
rect 12665 9094 12682 9158
rect 12746 9094 12763 9158
rect 12827 9094 12844 9158
rect 12908 9094 12925 9158
rect 12989 9094 13006 9158
rect 13070 9094 13087 9158
rect 13151 9094 13168 9158
rect 13232 9094 13249 9158
rect 13313 9094 13330 9158
rect 13394 9094 13411 9158
rect 13475 9094 13492 9158
rect 13556 9094 13573 9158
rect 13637 9094 13654 9158
rect 13718 9094 13735 9158
rect 13799 9094 13816 9158
rect 13880 9094 13897 9158
rect 13961 9094 13978 9158
rect 14042 9094 14059 9158
rect 14123 9094 14140 9158
rect 14204 9094 14221 9158
rect 14285 9094 14302 9158
rect 14366 9094 14383 9158
rect 14447 9094 14464 9158
rect 14528 9094 14545 9158
rect 14609 9094 14626 9158
rect 14690 9094 14707 9158
rect 14771 9094 14788 9158
rect 14852 9094 14858 9158
rect 10078 9072 14858 9094
rect 10078 9008 10084 9072
rect 10148 9008 10166 9072
rect 10230 9008 10248 9072
rect 10312 9008 10330 9072
rect 10394 9008 10412 9072
rect 10476 9008 10494 9072
rect 10558 9008 10576 9072
rect 10640 9008 10657 9072
rect 10721 9008 10738 9072
rect 10802 9008 10819 9072
rect 10883 9008 10900 9072
rect 10964 9008 10981 9072
rect 11045 9008 11062 9072
rect 11126 9008 11143 9072
rect 11207 9008 11224 9072
rect 11288 9008 11305 9072
rect 11369 9008 11386 9072
rect 11450 9008 11467 9072
rect 11531 9008 11548 9072
rect 11612 9008 11629 9072
rect 11693 9008 11710 9072
rect 11774 9008 11791 9072
rect 11855 9008 11872 9072
rect 11936 9008 11953 9072
rect 12017 9008 12034 9072
rect 12098 9008 12115 9072
rect 12179 9008 12196 9072
rect 12260 9008 12277 9072
rect 12341 9008 12358 9072
rect 12422 9008 12439 9072
rect 12503 9008 12520 9072
rect 12584 9008 12601 9072
rect 12665 9008 12682 9072
rect 12746 9008 12763 9072
rect 12827 9008 12844 9072
rect 12908 9008 12925 9072
rect 12989 9008 13006 9072
rect 13070 9008 13087 9072
rect 13151 9008 13168 9072
rect 13232 9008 13249 9072
rect 13313 9008 13330 9072
rect 13394 9008 13411 9072
rect 13475 9008 13492 9072
rect 13556 9008 13573 9072
rect 13637 9008 13654 9072
rect 13718 9008 13735 9072
rect 13799 9008 13816 9072
rect 13880 9008 13897 9072
rect 13961 9008 13978 9072
rect 14042 9008 14059 9072
rect 14123 9008 14140 9072
rect 14204 9008 14221 9072
rect 14285 9008 14302 9072
rect 14366 9008 14383 9072
rect 14447 9008 14464 9072
rect 14528 9008 14545 9072
rect 14609 9008 14626 9072
rect 14690 9008 14707 9072
rect 14771 9008 14788 9072
rect 14852 9008 14858 9072
rect 10078 8986 14858 9008
rect 10078 8922 10084 8986
rect 10148 8922 10166 8986
rect 10230 8922 10248 8986
rect 10312 8922 10330 8986
rect 10394 8922 10412 8986
rect 10476 8922 10494 8986
rect 10558 8922 10576 8986
rect 10640 8922 10657 8986
rect 10721 8922 10738 8986
rect 10802 8922 10819 8986
rect 10883 8922 10900 8986
rect 10964 8922 10981 8986
rect 11045 8922 11062 8986
rect 11126 8922 11143 8986
rect 11207 8922 11224 8986
rect 11288 8922 11305 8986
rect 11369 8922 11386 8986
rect 11450 8922 11467 8986
rect 11531 8922 11548 8986
rect 11612 8922 11629 8986
rect 11693 8922 11710 8986
rect 11774 8922 11791 8986
rect 11855 8922 11872 8986
rect 11936 8922 11953 8986
rect 12017 8922 12034 8986
rect 12098 8922 12115 8986
rect 12179 8922 12196 8986
rect 12260 8922 12277 8986
rect 12341 8922 12358 8986
rect 12422 8922 12439 8986
rect 12503 8922 12520 8986
rect 12584 8922 12601 8986
rect 12665 8922 12682 8986
rect 12746 8922 12763 8986
rect 12827 8922 12844 8986
rect 12908 8922 12925 8986
rect 12989 8922 13006 8986
rect 13070 8922 13087 8986
rect 13151 8922 13168 8986
rect 13232 8922 13249 8986
rect 13313 8922 13330 8986
rect 13394 8922 13411 8986
rect 13475 8922 13492 8986
rect 13556 8922 13573 8986
rect 13637 8922 13654 8986
rect 13718 8922 13735 8986
rect 13799 8922 13816 8986
rect 13880 8922 13897 8986
rect 13961 8922 13978 8986
rect 14042 8922 14059 8986
rect 14123 8922 14140 8986
rect 14204 8922 14221 8986
rect 14285 8922 14302 8986
rect 14366 8922 14383 8986
rect 14447 8922 14464 8986
rect 14528 8922 14545 8986
rect 14609 8922 14626 8986
rect 14690 8922 14707 8986
rect 14771 8922 14788 8986
rect 14852 8922 14858 8986
rect 10078 8900 14858 8922
rect 10078 8836 10084 8900
rect 10148 8836 10166 8900
rect 10230 8836 10248 8900
rect 10312 8836 10330 8900
rect 10394 8836 10412 8900
rect 10476 8836 10494 8900
rect 10558 8836 10576 8900
rect 10640 8836 10657 8900
rect 10721 8836 10738 8900
rect 10802 8836 10819 8900
rect 10883 8836 10900 8900
rect 10964 8836 10981 8900
rect 11045 8836 11062 8900
rect 11126 8836 11143 8900
rect 11207 8836 11224 8900
rect 11288 8836 11305 8900
rect 11369 8836 11386 8900
rect 11450 8836 11467 8900
rect 11531 8836 11548 8900
rect 11612 8836 11629 8900
rect 11693 8836 11710 8900
rect 11774 8836 11791 8900
rect 11855 8836 11872 8900
rect 11936 8836 11953 8900
rect 12017 8836 12034 8900
rect 12098 8836 12115 8900
rect 12179 8836 12196 8900
rect 12260 8836 12277 8900
rect 12341 8836 12358 8900
rect 12422 8836 12439 8900
rect 12503 8836 12520 8900
rect 12584 8836 12601 8900
rect 12665 8836 12682 8900
rect 12746 8836 12763 8900
rect 12827 8836 12844 8900
rect 12908 8836 12925 8900
rect 12989 8836 13006 8900
rect 13070 8836 13087 8900
rect 13151 8836 13168 8900
rect 13232 8836 13249 8900
rect 13313 8836 13330 8900
rect 13394 8836 13411 8900
rect 13475 8836 13492 8900
rect 13556 8836 13573 8900
rect 13637 8836 13654 8900
rect 13718 8836 13735 8900
rect 13799 8836 13816 8900
rect 13880 8836 13897 8900
rect 13961 8836 13978 8900
rect 14042 8836 14059 8900
rect 14123 8836 14140 8900
rect 14204 8836 14221 8900
rect 14285 8836 14302 8900
rect 14366 8836 14383 8900
rect 14447 8836 14464 8900
rect 14528 8836 14545 8900
rect 14609 8836 14626 8900
rect 14690 8836 14707 8900
rect 14771 8836 14788 8900
rect 14852 8836 14858 8900
rect 10078 8814 14858 8836
rect 10078 8750 10084 8814
rect 10148 8750 10166 8814
rect 10230 8750 10248 8814
rect 10312 8750 10330 8814
rect 10394 8750 10412 8814
rect 10476 8750 10494 8814
rect 10558 8750 10576 8814
rect 10640 8750 10657 8814
rect 10721 8750 10738 8814
rect 10802 8750 10819 8814
rect 10883 8750 10900 8814
rect 10964 8750 10981 8814
rect 11045 8750 11062 8814
rect 11126 8750 11143 8814
rect 11207 8750 11224 8814
rect 11288 8750 11305 8814
rect 11369 8750 11386 8814
rect 11450 8750 11467 8814
rect 11531 8750 11548 8814
rect 11612 8750 11629 8814
rect 11693 8750 11710 8814
rect 11774 8750 11791 8814
rect 11855 8750 11872 8814
rect 11936 8750 11953 8814
rect 12017 8750 12034 8814
rect 12098 8750 12115 8814
rect 12179 8750 12196 8814
rect 12260 8750 12277 8814
rect 12341 8750 12358 8814
rect 12422 8750 12439 8814
rect 12503 8750 12520 8814
rect 12584 8750 12601 8814
rect 12665 8750 12682 8814
rect 12746 8750 12763 8814
rect 12827 8750 12844 8814
rect 12908 8750 12925 8814
rect 12989 8750 13006 8814
rect 13070 8750 13087 8814
rect 13151 8750 13168 8814
rect 13232 8750 13249 8814
rect 13313 8750 13330 8814
rect 13394 8750 13411 8814
rect 13475 8750 13492 8814
rect 13556 8750 13573 8814
rect 13637 8750 13654 8814
rect 13718 8750 13735 8814
rect 13799 8750 13816 8814
rect 13880 8750 13897 8814
rect 13961 8750 13978 8814
rect 14042 8750 14059 8814
rect 14123 8750 14140 8814
rect 14204 8750 14221 8814
rect 14285 8750 14302 8814
rect 14366 8750 14383 8814
rect 14447 8750 14464 8814
rect 14528 8750 14545 8814
rect 14609 8750 14626 8814
rect 14690 8750 14707 8814
rect 14771 8750 14788 8814
rect 14852 8750 14858 8814
rect 10078 8728 14858 8750
rect 10078 8664 10084 8728
rect 10148 8664 10166 8728
rect 10230 8664 10248 8728
rect 10312 8664 10330 8728
rect 10394 8664 10412 8728
rect 10476 8664 10494 8728
rect 10558 8664 10576 8728
rect 10640 8664 10657 8728
rect 10721 8664 10738 8728
rect 10802 8664 10819 8728
rect 10883 8664 10900 8728
rect 10964 8664 10981 8728
rect 11045 8664 11062 8728
rect 11126 8664 11143 8728
rect 11207 8664 11224 8728
rect 11288 8664 11305 8728
rect 11369 8664 11386 8728
rect 11450 8664 11467 8728
rect 11531 8664 11548 8728
rect 11612 8664 11629 8728
rect 11693 8664 11710 8728
rect 11774 8664 11791 8728
rect 11855 8664 11872 8728
rect 11936 8664 11953 8728
rect 12017 8664 12034 8728
rect 12098 8664 12115 8728
rect 12179 8664 12196 8728
rect 12260 8664 12277 8728
rect 12341 8664 12358 8728
rect 12422 8664 12439 8728
rect 12503 8664 12520 8728
rect 12584 8664 12601 8728
rect 12665 8664 12682 8728
rect 12746 8664 12763 8728
rect 12827 8664 12844 8728
rect 12908 8664 12925 8728
rect 12989 8664 13006 8728
rect 13070 8664 13087 8728
rect 13151 8664 13168 8728
rect 13232 8664 13249 8728
rect 13313 8664 13330 8728
rect 13394 8664 13411 8728
rect 13475 8664 13492 8728
rect 13556 8664 13573 8728
rect 13637 8664 13654 8728
rect 13718 8664 13735 8728
rect 13799 8664 13816 8728
rect 13880 8664 13897 8728
rect 13961 8664 13978 8728
rect 14042 8664 14059 8728
rect 14123 8664 14140 8728
rect 14204 8664 14221 8728
rect 14285 8664 14302 8728
rect 14366 8664 14383 8728
rect 14447 8664 14464 8728
rect 14528 8664 14545 8728
rect 14609 8664 14626 8728
rect 14690 8664 14707 8728
rect 14771 8664 14788 8728
rect 14852 8664 14858 8728
rect 10078 8642 14858 8664
rect 10078 8578 10084 8642
rect 10148 8578 10166 8642
rect 10230 8578 10248 8642
rect 10312 8578 10330 8642
rect 10394 8578 10412 8642
rect 10476 8578 10494 8642
rect 10558 8578 10576 8642
rect 10640 8578 10657 8642
rect 10721 8578 10738 8642
rect 10802 8578 10819 8642
rect 10883 8578 10900 8642
rect 10964 8578 10981 8642
rect 11045 8578 11062 8642
rect 11126 8578 11143 8642
rect 11207 8578 11224 8642
rect 11288 8578 11305 8642
rect 11369 8578 11386 8642
rect 11450 8578 11467 8642
rect 11531 8578 11548 8642
rect 11612 8578 11629 8642
rect 11693 8578 11710 8642
rect 11774 8578 11791 8642
rect 11855 8578 11872 8642
rect 11936 8578 11953 8642
rect 12017 8578 12034 8642
rect 12098 8578 12115 8642
rect 12179 8578 12196 8642
rect 12260 8578 12277 8642
rect 12341 8578 12358 8642
rect 12422 8578 12439 8642
rect 12503 8578 12520 8642
rect 12584 8578 12601 8642
rect 12665 8578 12682 8642
rect 12746 8578 12763 8642
rect 12827 8578 12844 8642
rect 12908 8578 12925 8642
rect 12989 8578 13006 8642
rect 13070 8578 13087 8642
rect 13151 8578 13168 8642
rect 13232 8578 13249 8642
rect 13313 8578 13330 8642
rect 13394 8578 13411 8642
rect 13475 8578 13492 8642
rect 13556 8578 13573 8642
rect 13637 8578 13654 8642
rect 13718 8578 13735 8642
rect 13799 8578 13816 8642
rect 13880 8578 13897 8642
rect 13961 8578 13978 8642
rect 14042 8578 14059 8642
rect 14123 8578 14140 8642
rect 14204 8578 14221 8642
rect 14285 8578 14302 8642
rect 14366 8578 14383 8642
rect 14447 8578 14464 8642
rect 14528 8578 14545 8642
rect 14609 8578 14626 8642
rect 14690 8578 14707 8642
rect 14771 8578 14788 8642
rect 14852 8578 14858 8642
rect 10078 8556 14858 8578
rect 10078 8492 10084 8556
rect 10148 8492 10166 8556
rect 10230 8492 10248 8556
rect 10312 8492 10330 8556
rect 10394 8492 10412 8556
rect 10476 8492 10494 8556
rect 10558 8492 10576 8556
rect 10640 8492 10657 8556
rect 10721 8492 10738 8556
rect 10802 8492 10819 8556
rect 10883 8492 10900 8556
rect 10964 8492 10981 8556
rect 11045 8492 11062 8556
rect 11126 8492 11143 8556
rect 11207 8492 11224 8556
rect 11288 8492 11305 8556
rect 11369 8492 11386 8556
rect 11450 8492 11467 8556
rect 11531 8492 11548 8556
rect 11612 8492 11629 8556
rect 11693 8492 11710 8556
rect 11774 8492 11791 8556
rect 11855 8492 11872 8556
rect 11936 8492 11953 8556
rect 12017 8492 12034 8556
rect 12098 8492 12115 8556
rect 12179 8492 12196 8556
rect 12260 8492 12277 8556
rect 12341 8492 12358 8556
rect 12422 8492 12439 8556
rect 12503 8492 12520 8556
rect 12584 8492 12601 8556
rect 12665 8492 12682 8556
rect 12746 8492 12763 8556
rect 12827 8492 12844 8556
rect 12908 8492 12925 8556
rect 12989 8492 13006 8556
rect 13070 8492 13087 8556
rect 13151 8492 13168 8556
rect 13232 8492 13249 8556
rect 13313 8492 13330 8556
rect 13394 8492 13411 8556
rect 13475 8492 13492 8556
rect 13556 8492 13573 8556
rect 13637 8492 13654 8556
rect 13718 8492 13735 8556
rect 13799 8492 13816 8556
rect 13880 8492 13897 8556
rect 13961 8492 13978 8556
rect 14042 8492 14059 8556
rect 14123 8492 14140 8556
rect 14204 8492 14221 8556
rect 14285 8492 14302 8556
rect 14366 8492 14383 8556
rect 14447 8492 14464 8556
rect 14528 8492 14545 8556
rect 14609 8492 14626 8556
rect 14690 8492 14707 8556
rect 14771 8492 14788 8556
rect 14852 8492 14858 8556
rect 10078 8470 14858 8492
rect 10078 8406 10084 8470
rect 10148 8406 10166 8470
rect 10230 8406 10248 8470
rect 10312 8406 10330 8470
rect 10394 8406 10412 8470
rect 10476 8406 10494 8470
rect 10558 8406 10576 8470
rect 10640 8406 10657 8470
rect 10721 8406 10738 8470
rect 10802 8406 10819 8470
rect 10883 8406 10900 8470
rect 10964 8406 10981 8470
rect 11045 8406 11062 8470
rect 11126 8406 11143 8470
rect 11207 8406 11224 8470
rect 11288 8406 11305 8470
rect 11369 8406 11386 8470
rect 11450 8406 11467 8470
rect 11531 8406 11548 8470
rect 11612 8406 11629 8470
rect 11693 8406 11710 8470
rect 11774 8406 11791 8470
rect 11855 8406 11872 8470
rect 11936 8406 11953 8470
rect 12017 8406 12034 8470
rect 12098 8406 12115 8470
rect 12179 8406 12196 8470
rect 12260 8406 12277 8470
rect 12341 8406 12358 8470
rect 12422 8406 12439 8470
rect 12503 8406 12520 8470
rect 12584 8406 12601 8470
rect 12665 8406 12682 8470
rect 12746 8406 12763 8470
rect 12827 8406 12844 8470
rect 12908 8406 12925 8470
rect 12989 8406 13006 8470
rect 13070 8406 13087 8470
rect 13151 8406 13168 8470
rect 13232 8406 13249 8470
rect 13313 8406 13330 8470
rect 13394 8406 13411 8470
rect 13475 8406 13492 8470
rect 13556 8406 13573 8470
rect 13637 8406 13654 8470
rect 13718 8406 13735 8470
rect 13799 8406 13816 8470
rect 13880 8406 13897 8470
rect 13961 8406 13978 8470
rect 14042 8406 14059 8470
rect 14123 8406 14140 8470
rect 14204 8406 14221 8470
rect 14285 8406 14302 8470
rect 14366 8406 14383 8470
rect 14447 8406 14464 8470
rect 14528 8406 14545 8470
rect 14609 8406 14626 8470
rect 14690 8406 14707 8470
rect 14771 8406 14788 8470
rect 14852 8406 14858 8470
rect 10078 8384 14858 8406
rect 10078 8320 10084 8384
rect 10148 8320 10166 8384
rect 10230 8320 10248 8384
rect 10312 8320 10330 8384
rect 10394 8320 10412 8384
rect 10476 8320 10494 8384
rect 10558 8320 10576 8384
rect 10640 8320 10657 8384
rect 10721 8320 10738 8384
rect 10802 8320 10819 8384
rect 10883 8320 10900 8384
rect 10964 8320 10981 8384
rect 11045 8320 11062 8384
rect 11126 8320 11143 8384
rect 11207 8320 11224 8384
rect 11288 8320 11305 8384
rect 11369 8320 11386 8384
rect 11450 8320 11467 8384
rect 11531 8320 11548 8384
rect 11612 8320 11629 8384
rect 11693 8320 11710 8384
rect 11774 8320 11791 8384
rect 11855 8320 11872 8384
rect 11936 8320 11953 8384
rect 12017 8320 12034 8384
rect 12098 8320 12115 8384
rect 12179 8320 12196 8384
rect 12260 8320 12277 8384
rect 12341 8320 12358 8384
rect 12422 8320 12439 8384
rect 12503 8320 12520 8384
rect 12584 8320 12601 8384
rect 12665 8320 12682 8384
rect 12746 8320 12763 8384
rect 12827 8320 12844 8384
rect 12908 8320 12925 8384
rect 12989 8320 13006 8384
rect 13070 8320 13087 8384
rect 13151 8320 13168 8384
rect 13232 8320 13249 8384
rect 13313 8320 13330 8384
rect 13394 8320 13411 8384
rect 13475 8320 13492 8384
rect 13556 8320 13573 8384
rect 13637 8320 13654 8384
rect 13718 8320 13735 8384
rect 13799 8320 13816 8384
rect 13880 8320 13897 8384
rect 13961 8320 13978 8384
rect 14042 8320 14059 8384
rect 14123 8320 14140 8384
rect 14204 8320 14221 8384
rect 14285 8320 14302 8384
rect 14366 8320 14383 8384
rect 14447 8320 14464 8384
rect 14528 8320 14545 8384
rect 14609 8320 14626 8384
rect 14690 8320 14707 8384
rect 14771 8320 14788 8384
rect 14852 8320 14858 8384
rect 10078 8318 14858 8320
<< via3 >>
rect 200 9180 264 9244
rect 281 9180 345 9244
rect 362 9180 426 9244
rect 443 9180 507 9244
rect 524 9180 588 9244
rect 605 9180 669 9244
rect 686 9180 750 9244
rect 767 9180 831 9244
rect 848 9180 912 9244
rect 929 9180 993 9244
rect 1010 9180 1074 9244
rect 1091 9180 1155 9244
rect 1172 9180 1236 9244
rect 1253 9180 1317 9244
rect 1334 9180 1398 9244
rect 1415 9180 1479 9244
rect 1496 9180 1560 9244
rect 1577 9180 1641 9244
rect 1658 9180 1722 9244
rect 1739 9180 1803 9244
rect 1820 9180 1884 9244
rect 1901 9180 1965 9244
rect 1982 9180 2046 9244
rect 2063 9180 2127 9244
rect 2144 9180 2208 9244
rect 2225 9180 2289 9244
rect 2306 9180 2370 9244
rect 2387 9180 2451 9244
rect 2468 9180 2532 9244
rect 2549 9180 2613 9244
rect 2630 9180 2694 9244
rect 2711 9180 2775 9244
rect 2792 9180 2856 9244
rect 2873 9180 2937 9244
rect 2954 9180 3018 9244
rect 3035 9180 3099 9244
rect 3116 9180 3180 9244
rect 3197 9180 3261 9244
rect 3278 9180 3342 9244
rect 3359 9180 3423 9244
rect 3440 9180 3504 9244
rect 3521 9180 3585 9244
rect 3602 9180 3666 9244
rect 3683 9180 3747 9244
rect 3764 9180 3828 9244
rect 3845 9180 3909 9244
rect 3926 9180 3990 9244
rect 4007 9180 4071 9244
rect 4088 9180 4152 9244
rect 4169 9180 4233 9244
rect 4249 9180 4313 9244
rect 4329 9180 4393 9244
rect 4409 9180 4473 9244
rect 4489 9180 4553 9244
rect 4569 9180 4633 9244
rect 4649 9180 4713 9244
rect 4729 9180 4793 9244
rect 4809 9180 4873 9244
rect 200 9094 264 9158
rect 281 9094 345 9158
rect 362 9094 426 9158
rect 443 9094 507 9158
rect 524 9094 588 9158
rect 605 9094 669 9158
rect 686 9094 750 9158
rect 767 9094 831 9158
rect 848 9094 912 9158
rect 929 9094 993 9158
rect 1010 9094 1074 9158
rect 1091 9094 1155 9158
rect 1172 9094 1236 9158
rect 1253 9094 1317 9158
rect 1334 9094 1398 9158
rect 1415 9094 1479 9158
rect 1496 9094 1560 9158
rect 1577 9094 1641 9158
rect 1658 9094 1722 9158
rect 1739 9094 1803 9158
rect 1820 9094 1884 9158
rect 1901 9094 1965 9158
rect 1982 9094 2046 9158
rect 2063 9094 2127 9158
rect 2144 9094 2208 9158
rect 2225 9094 2289 9158
rect 2306 9094 2370 9158
rect 2387 9094 2451 9158
rect 2468 9094 2532 9158
rect 2549 9094 2613 9158
rect 2630 9094 2694 9158
rect 2711 9094 2775 9158
rect 2792 9094 2856 9158
rect 2873 9094 2937 9158
rect 2954 9094 3018 9158
rect 3035 9094 3099 9158
rect 3116 9094 3180 9158
rect 3197 9094 3261 9158
rect 3278 9094 3342 9158
rect 3359 9094 3423 9158
rect 3440 9094 3504 9158
rect 3521 9094 3585 9158
rect 3602 9094 3666 9158
rect 3683 9094 3747 9158
rect 3764 9094 3828 9158
rect 3845 9094 3909 9158
rect 3926 9094 3990 9158
rect 4007 9094 4071 9158
rect 4088 9094 4152 9158
rect 4169 9094 4233 9158
rect 4249 9094 4313 9158
rect 4329 9094 4393 9158
rect 4409 9094 4473 9158
rect 4489 9094 4553 9158
rect 4569 9094 4633 9158
rect 4649 9094 4713 9158
rect 4729 9094 4793 9158
rect 4809 9094 4873 9158
rect 200 9008 264 9072
rect 281 9008 345 9072
rect 362 9008 426 9072
rect 443 9008 507 9072
rect 524 9008 588 9072
rect 605 9008 669 9072
rect 686 9008 750 9072
rect 767 9008 831 9072
rect 848 9008 912 9072
rect 929 9008 993 9072
rect 1010 9008 1074 9072
rect 1091 9008 1155 9072
rect 1172 9008 1236 9072
rect 1253 9008 1317 9072
rect 1334 9008 1398 9072
rect 1415 9008 1479 9072
rect 1496 9008 1560 9072
rect 1577 9008 1641 9072
rect 1658 9008 1722 9072
rect 1739 9008 1803 9072
rect 1820 9008 1884 9072
rect 1901 9008 1965 9072
rect 1982 9008 2046 9072
rect 2063 9008 2127 9072
rect 2144 9008 2208 9072
rect 2225 9008 2289 9072
rect 2306 9008 2370 9072
rect 2387 9008 2451 9072
rect 2468 9008 2532 9072
rect 2549 9008 2613 9072
rect 2630 9008 2694 9072
rect 2711 9008 2775 9072
rect 2792 9008 2856 9072
rect 2873 9008 2937 9072
rect 2954 9008 3018 9072
rect 3035 9008 3099 9072
rect 3116 9008 3180 9072
rect 3197 9008 3261 9072
rect 3278 9008 3342 9072
rect 3359 9008 3423 9072
rect 3440 9008 3504 9072
rect 3521 9008 3585 9072
rect 3602 9008 3666 9072
rect 3683 9008 3747 9072
rect 3764 9008 3828 9072
rect 3845 9008 3909 9072
rect 3926 9008 3990 9072
rect 4007 9008 4071 9072
rect 4088 9008 4152 9072
rect 4169 9008 4233 9072
rect 4249 9008 4313 9072
rect 4329 9008 4393 9072
rect 4409 9008 4473 9072
rect 4489 9008 4553 9072
rect 4569 9008 4633 9072
rect 4649 9008 4713 9072
rect 4729 9008 4793 9072
rect 4809 9008 4873 9072
rect 200 8922 264 8986
rect 281 8922 345 8986
rect 362 8922 426 8986
rect 443 8922 507 8986
rect 524 8922 588 8986
rect 605 8922 669 8986
rect 686 8922 750 8986
rect 767 8922 831 8986
rect 848 8922 912 8986
rect 929 8922 993 8986
rect 1010 8922 1074 8986
rect 1091 8922 1155 8986
rect 1172 8922 1236 8986
rect 1253 8922 1317 8986
rect 1334 8922 1398 8986
rect 1415 8922 1479 8986
rect 1496 8922 1560 8986
rect 1577 8922 1641 8986
rect 1658 8922 1722 8986
rect 1739 8922 1803 8986
rect 1820 8922 1884 8986
rect 1901 8922 1965 8986
rect 1982 8922 2046 8986
rect 2063 8922 2127 8986
rect 2144 8922 2208 8986
rect 2225 8922 2289 8986
rect 2306 8922 2370 8986
rect 2387 8922 2451 8986
rect 2468 8922 2532 8986
rect 2549 8922 2613 8986
rect 2630 8922 2694 8986
rect 2711 8922 2775 8986
rect 2792 8922 2856 8986
rect 2873 8922 2937 8986
rect 2954 8922 3018 8986
rect 3035 8922 3099 8986
rect 3116 8922 3180 8986
rect 3197 8922 3261 8986
rect 3278 8922 3342 8986
rect 3359 8922 3423 8986
rect 3440 8922 3504 8986
rect 3521 8922 3585 8986
rect 3602 8922 3666 8986
rect 3683 8922 3747 8986
rect 3764 8922 3828 8986
rect 3845 8922 3909 8986
rect 3926 8922 3990 8986
rect 4007 8922 4071 8986
rect 4088 8922 4152 8986
rect 4169 8922 4233 8986
rect 4249 8922 4313 8986
rect 4329 8922 4393 8986
rect 4409 8922 4473 8986
rect 4489 8922 4553 8986
rect 4569 8922 4633 8986
rect 4649 8922 4713 8986
rect 4729 8922 4793 8986
rect 4809 8922 4873 8986
rect 200 8836 264 8900
rect 281 8836 345 8900
rect 362 8836 426 8900
rect 443 8836 507 8900
rect 524 8836 588 8900
rect 605 8836 669 8900
rect 686 8836 750 8900
rect 767 8836 831 8900
rect 848 8836 912 8900
rect 929 8836 993 8900
rect 1010 8836 1074 8900
rect 1091 8836 1155 8900
rect 1172 8836 1236 8900
rect 1253 8836 1317 8900
rect 1334 8836 1398 8900
rect 1415 8836 1479 8900
rect 1496 8836 1560 8900
rect 1577 8836 1641 8900
rect 1658 8836 1722 8900
rect 1739 8836 1803 8900
rect 1820 8836 1884 8900
rect 1901 8836 1965 8900
rect 1982 8836 2046 8900
rect 2063 8836 2127 8900
rect 2144 8836 2208 8900
rect 2225 8836 2289 8900
rect 2306 8836 2370 8900
rect 2387 8836 2451 8900
rect 2468 8836 2532 8900
rect 2549 8836 2613 8900
rect 2630 8836 2694 8900
rect 2711 8836 2775 8900
rect 2792 8836 2856 8900
rect 2873 8836 2937 8900
rect 2954 8836 3018 8900
rect 3035 8836 3099 8900
rect 3116 8836 3180 8900
rect 3197 8836 3261 8900
rect 3278 8836 3342 8900
rect 3359 8836 3423 8900
rect 3440 8836 3504 8900
rect 3521 8836 3585 8900
rect 3602 8836 3666 8900
rect 3683 8836 3747 8900
rect 3764 8836 3828 8900
rect 3845 8836 3909 8900
rect 3926 8836 3990 8900
rect 4007 8836 4071 8900
rect 4088 8836 4152 8900
rect 4169 8836 4233 8900
rect 4249 8836 4313 8900
rect 4329 8836 4393 8900
rect 4409 8836 4473 8900
rect 4489 8836 4553 8900
rect 4569 8836 4633 8900
rect 4649 8836 4713 8900
rect 4729 8836 4793 8900
rect 4809 8836 4873 8900
rect 200 8750 264 8814
rect 281 8750 345 8814
rect 362 8750 426 8814
rect 443 8750 507 8814
rect 524 8750 588 8814
rect 605 8750 669 8814
rect 686 8750 750 8814
rect 767 8750 831 8814
rect 848 8750 912 8814
rect 929 8750 993 8814
rect 1010 8750 1074 8814
rect 1091 8750 1155 8814
rect 1172 8750 1236 8814
rect 1253 8750 1317 8814
rect 1334 8750 1398 8814
rect 1415 8750 1479 8814
rect 1496 8750 1560 8814
rect 1577 8750 1641 8814
rect 1658 8750 1722 8814
rect 1739 8750 1803 8814
rect 1820 8750 1884 8814
rect 1901 8750 1965 8814
rect 1982 8750 2046 8814
rect 2063 8750 2127 8814
rect 2144 8750 2208 8814
rect 2225 8750 2289 8814
rect 2306 8750 2370 8814
rect 2387 8750 2451 8814
rect 2468 8750 2532 8814
rect 2549 8750 2613 8814
rect 2630 8750 2694 8814
rect 2711 8750 2775 8814
rect 2792 8750 2856 8814
rect 2873 8750 2937 8814
rect 2954 8750 3018 8814
rect 3035 8750 3099 8814
rect 3116 8750 3180 8814
rect 3197 8750 3261 8814
rect 3278 8750 3342 8814
rect 3359 8750 3423 8814
rect 3440 8750 3504 8814
rect 3521 8750 3585 8814
rect 3602 8750 3666 8814
rect 3683 8750 3747 8814
rect 3764 8750 3828 8814
rect 3845 8750 3909 8814
rect 3926 8750 3990 8814
rect 4007 8750 4071 8814
rect 4088 8750 4152 8814
rect 4169 8750 4233 8814
rect 4249 8750 4313 8814
rect 4329 8750 4393 8814
rect 4409 8750 4473 8814
rect 4489 8750 4553 8814
rect 4569 8750 4633 8814
rect 4649 8750 4713 8814
rect 4729 8750 4793 8814
rect 4809 8750 4873 8814
rect 200 8664 264 8728
rect 281 8664 345 8728
rect 362 8664 426 8728
rect 443 8664 507 8728
rect 524 8664 588 8728
rect 605 8664 669 8728
rect 686 8664 750 8728
rect 767 8664 831 8728
rect 848 8664 912 8728
rect 929 8664 993 8728
rect 1010 8664 1074 8728
rect 1091 8664 1155 8728
rect 1172 8664 1236 8728
rect 1253 8664 1317 8728
rect 1334 8664 1398 8728
rect 1415 8664 1479 8728
rect 1496 8664 1560 8728
rect 1577 8664 1641 8728
rect 1658 8664 1722 8728
rect 1739 8664 1803 8728
rect 1820 8664 1884 8728
rect 1901 8664 1965 8728
rect 1982 8664 2046 8728
rect 2063 8664 2127 8728
rect 2144 8664 2208 8728
rect 2225 8664 2289 8728
rect 2306 8664 2370 8728
rect 2387 8664 2451 8728
rect 2468 8664 2532 8728
rect 2549 8664 2613 8728
rect 2630 8664 2694 8728
rect 2711 8664 2775 8728
rect 2792 8664 2856 8728
rect 2873 8664 2937 8728
rect 2954 8664 3018 8728
rect 3035 8664 3099 8728
rect 3116 8664 3180 8728
rect 3197 8664 3261 8728
rect 3278 8664 3342 8728
rect 3359 8664 3423 8728
rect 3440 8664 3504 8728
rect 3521 8664 3585 8728
rect 3602 8664 3666 8728
rect 3683 8664 3747 8728
rect 3764 8664 3828 8728
rect 3845 8664 3909 8728
rect 3926 8664 3990 8728
rect 4007 8664 4071 8728
rect 4088 8664 4152 8728
rect 4169 8664 4233 8728
rect 4249 8664 4313 8728
rect 4329 8664 4393 8728
rect 4409 8664 4473 8728
rect 4489 8664 4553 8728
rect 4569 8664 4633 8728
rect 4649 8664 4713 8728
rect 4729 8664 4793 8728
rect 4809 8664 4873 8728
rect 200 8578 264 8642
rect 281 8578 345 8642
rect 362 8578 426 8642
rect 443 8578 507 8642
rect 524 8578 588 8642
rect 605 8578 669 8642
rect 686 8578 750 8642
rect 767 8578 831 8642
rect 848 8578 912 8642
rect 929 8578 993 8642
rect 1010 8578 1074 8642
rect 1091 8578 1155 8642
rect 1172 8578 1236 8642
rect 1253 8578 1317 8642
rect 1334 8578 1398 8642
rect 1415 8578 1479 8642
rect 1496 8578 1560 8642
rect 1577 8578 1641 8642
rect 1658 8578 1722 8642
rect 1739 8578 1803 8642
rect 1820 8578 1884 8642
rect 1901 8578 1965 8642
rect 1982 8578 2046 8642
rect 2063 8578 2127 8642
rect 2144 8578 2208 8642
rect 2225 8578 2289 8642
rect 2306 8578 2370 8642
rect 2387 8578 2451 8642
rect 2468 8578 2532 8642
rect 2549 8578 2613 8642
rect 2630 8578 2694 8642
rect 2711 8578 2775 8642
rect 2792 8578 2856 8642
rect 2873 8578 2937 8642
rect 2954 8578 3018 8642
rect 3035 8578 3099 8642
rect 3116 8578 3180 8642
rect 3197 8578 3261 8642
rect 3278 8578 3342 8642
rect 3359 8578 3423 8642
rect 3440 8578 3504 8642
rect 3521 8578 3585 8642
rect 3602 8578 3666 8642
rect 3683 8578 3747 8642
rect 3764 8578 3828 8642
rect 3845 8578 3909 8642
rect 3926 8578 3990 8642
rect 4007 8578 4071 8642
rect 4088 8578 4152 8642
rect 4169 8578 4233 8642
rect 4249 8578 4313 8642
rect 4329 8578 4393 8642
rect 4409 8578 4473 8642
rect 4489 8578 4553 8642
rect 4569 8578 4633 8642
rect 4649 8578 4713 8642
rect 4729 8578 4793 8642
rect 4809 8578 4873 8642
rect 200 8492 264 8556
rect 281 8492 345 8556
rect 362 8492 426 8556
rect 443 8492 507 8556
rect 524 8492 588 8556
rect 605 8492 669 8556
rect 686 8492 750 8556
rect 767 8492 831 8556
rect 848 8492 912 8556
rect 929 8492 993 8556
rect 1010 8492 1074 8556
rect 1091 8492 1155 8556
rect 1172 8492 1236 8556
rect 1253 8492 1317 8556
rect 1334 8492 1398 8556
rect 1415 8492 1479 8556
rect 1496 8492 1560 8556
rect 1577 8492 1641 8556
rect 1658 8492 1722 8556
rect 1739 8492 1803 8556
rect 1820 8492 1884 8556
rect 1901 8492 1965 8556
rect 1982 8492 2046 8556
rect 2063 8492 2127 8556
rect 2144 8492 2208 8556
rect 2225 8492 2289 8556
rect 2306 8492 2370 8556
rect 2387 8492 2451 8556
rect 2468 8492 2532 8556
rect 2549 8492 2613 8556
rect 2630 8492 2694 8556
rect 2711 8492 2775 8556
rect 2792 8492 2856 8556
rect 2873 8492 2937 8556
rect 2954 8492 3018 8556
rect 3035 8492 3099 8556
rect 3116 8492 3180 8556
rect 3197 8492 3261 8556
rect 3278 8492 3342 8556
rect 3359 8492 3423 8556
rect 3440 8492 3504 8556
rect 3521 8492 3585 8556
rect 3602 8492 3666 8556
rect 3683 8492 3747 8556
rect 3764 8492 3828 8556
rect 3845 8492 3909 8556
rect 3926 8492 3990 8556
rect 4007 8492 4071 8556
rect 4088 8492 4152 8556
rect 4169 8492 4233 8556
rect 4249 8492 4313 8556
rect 4329 8492 4393 8556
rect 4409 8492 4473 8556
rect 4489 8492 4553 8556
rect 4569 8492 4633 8556
rect 4649 8492 4713 8556
rect 4729 8492 4793 8556
rect 4809 8492 4873 8556
rect 200 8406 264 8470
rect 281 8406 345 8470
rect 362 8406 426 8470
rect 443 8406 507 8470
rect 524 8406 588 8470
rect 605 8406 669 8470
rect 686 8406 750 8470
rect 767 8406 831 8470
rect 848 8406 912 8470
rect 929 8406 993 8470
rect 1010 8406 1074 8470
rect 1091 8406 1155 8470
rect 1172 8406 1236 8470
rect 1253 8406 1317 8470
rect 1334 8406 1398 8470
rect 1415 8406 1479 8470
rect 1496 8406 1560 8470
rect 1577 8406 1641 8470
rect 1658 8406 1722 8470
rect 1739 8406 1803 8470
rect 1820 8406 1884 8470
rect 1901 8406 1965 8470
rect 1982 8406 2046 8470
rect 2063 8406 2127 8470
rect 2144 8406 2208 8470
rect 2225 8406 2289 8470
rect 2306 8406 2370 8470
rect 2387 8406 2451 8470
rect 2468 8406 2532 8470
rect 2549 8406 2613 8470
rect 2630 8406 2694 8470
rect 2711 8406 2775 8470
rect 2792 8406 2856 8470
rect 2873 8406 2937 8470
rect 2954 8406 3018 8470
rect 3035 8406 3099 8470
rect 3116 8406 3180 8470
rect 3197 8406 3261 8470
rect 3278 8406 3342 8470
rect 3359 8406 3423 8470
rect 3440 8406 3504 8470
rect 3521 8406 3585 8470
rect 3602 8406 3666 8470
rect 3683 8406 3747 8470
rect 3764 8406 3828 8470
rect 3845 8406 3909 8470
rect 3926 8406 3990 8470
rect 4007 8406 4071 8470
rect 4088 8406 4152 8470
rect 4169 8406 4233 8470
rect 4249 8406 4313 8470
rect 4329 8406 4393 8470
rect 4409 8406 4473 8470
rect 4489 8406 4553 8470
rect 4569 8406 4633 8470
rect 4649 8406 4713 8470
rect 4729 8406 4793 8470
rect 4809 8406 4873 8470
rect 200 8320 264 8384
rect 281 8320 345 8384
rect 362 8320 426 8384
rect 443 8320 507 8384
rect 524 8320 588 8384
rect 605 8320 669 8384
rect 686 8320 750 8384
rect 767 8320 831 8384
rect 848 8320 912 8384
rect 929 8320 993 8384
rect 1010 8320 1074 8384
rect 1091 8320 1155 8384
rect 1172 8320 1236 8384
rect 1253 8320 1317 8384
rect 1334 8320 1398 8384
rect 1415 8320 1479 8384
rect 1496 8320 1560 8384
rect 1577 8320 1641 8384
rect 1658 8320 1722 8384
rect 1739 8320 1803 8384
rect 1820 8320 1884 8384
rect 1901 8320 1965 8384
rect 1982 8320 2046 8384
rect 2063 8320 2127 8384
rect 2144 8320 2208 8384
rect 2225 8320 2289 8384
rect 2306 8320 2370 8384
rect 2387 8320 2451 8384
rect 2468 8320 2532 8384
rect 2549 8320 2613 8384
rect 2630 8320 2694 8384
rect 2711 8320 2775 8384
rect 2792 8320 2856 8384
rect 2873 8320 2937 8384
rect 2954 8320 3018 8384
rect 3035 8320 3099 8384
rect 3116 8320 3180 8384
rect 3197 8320 3261 8384
rect 3278 8320 3342 8384
rect 3359 8320 3423 8384
rect 3440 8320 3504 8384
rect 3521 8320 3585 8384
rect 3602 8320 3666 8384
rect 3683 8320 3747 8384
rect 3764 8320 3828 8384
rect 3845 8320 3909 8384
rect 3926 8320 3990 8384
rect 4007 8320 4071 8384
rect 4088 8320 4152 8384
rect 4169 8320 4233 8384
rect 4249 8320 4313 8384
rect 4329 8320 4393 8384
rect 4409 8320 4473 8384
rect 4489 8320 4553 8384
rect 4569 8320 4633 8384
rect 4649 8320 4713 8384
rect 4729 8320 4793 8384
rect 4809 8320 4873 8384
rect 10084 9180 10148 9244
rect 10166 9180 10230 9244
rect 10248 9180 10312 9244
rect 10330 9180 10394 9244
rect 10412 9180 10476 9244
rect 10494 9180 10558 9244
rect 10576 9180 10640 9244
rect 10657 9180 10721 9244
rect 10738 9180 10802 9244
rect 10819 9180 10883 9244
rect 10900 9180 10964 9244
rect 10981 9180 11045 9244
rect 11062 9180 11126 9244
rect 11143 9180 11207 9244
rect 11224 9180 11288 9244
rect 11305 9180 11369 9244
rect 11386 9180 11450 9244
rect 11467 9180 11531 9244
rect 11548 9180 11612 9244
rect 11629 9180 11693 9244
rect 11710 9180 11774 9244
rect 11791 9180 11855 9244
rect 11872 9180 11936 9244
rect 11953 9180 12017 9244
rect 12034 9180 12098 9244
rect 12115 9180 12179 9244
rect 12196 9180 12260 9244
rect 12277 9180 12341 9244
rect 12358 9180 12422 9244
rect 12439 9180 12503 9244
rect 12520 9180 12584 9244
rect 12601 9180 12665 9244
rect 12682 9180 12746 9244
rect 12763 9180 12827 9244
rect 12844 9180 12908 9244
rect 12925 9180 12989 9244
rect 13006 9180 13070 9244
rect 13087 9180 13151 9244
rect 13168 9180 13232 9244
rect 13249 9180 13313 9244
rect 13330 9180 13394 9244
rect 13411 9180 13475 9244
rect 13492 9180 13556 9244
rect 13573 9180 13637 9244
rect 13654 9180 13718 9244
rect 13735 9180 13799 9244
rect 13816 9180 13880 9244
rect 13897 9180 13961 9244
rect 13978 9180 14042 9244
rect 14059 9180 14123 9244
rect 14140 9180 14204 9244
rect 14221 9180 14285 9244
rect 14302 9180 14366 9244
rect 14383 9180 14447 9244
rect 14464 9180 14528 9244
rect 14545 9180 14609 9244
rect 14626 9180 14690 9244
rect 14707 9180 14771 9244
rect 14788 9180 14852 9244
rect 10084 9094 10148 9158
rect 10166 9094 10230 9158
rect 10248 9094 10312 9158
rect 10330 9094 10394 9158
rect 10412 9094 10476 9158
rect 10494 9094 10558 9158
rect 10576 9094 10640 9158
rect 10657 9094 10721 9158
rect 10738 9094 10802 9158
rect 10819 9094 10883 9158
rect 10900 9094 10964 9158
rect 10981 9094 11045 9158
rect 11062 9094 11126 9158
rect 11143 9094 11207 9158
rect 11224 9094 11288 9158
rect 11305 9094 11369 9158
rect 11386 9094 11450 9158
rect 11467 9094 11531 9158
rect 11548 9094 11612 9158
rect 11629 9094 11693 9158
rect 11710 9094 11774 9158
rect 11791 9094 11855 9158
rect 11872 9094 11936 9158
rect 11953 9094 12017 9158
rect 12034 9094 12098 9158
rect 12115 9094 12179 9158
rect 12196 9094 12260 9158
rect 12277 9094 12341 9158
rect 12358 9094 12422 9158
rect 12439 9094 12503 9158
rect 12520 9094 12584 9158
rect 12601 9094 12665 9158
rect 12682 9094 12746 9158
rect 12763 9094 12827 9158
rect 12844 9094 12908 9158
rect 12925 9094 12989 9158
rect 13006 9094 13070 9158
rect 13087 9094 13151 9158
rect 13168 9094 13232 9158
rect 13249 9094 13313 9158
rect 13330 9094 13394 9158
rect 13411 9094 13475 9158
rect 13492 9094 13556 9158
rect 13573 9094 13637 9158
rect 13654 9094 13718 9158
rect 13735 9094 13799 9158
rect 13816 9094 13880 9158
rect 13897 9094 13961 9158
rect 13978 9094 14042 9158
rect 14059 9094 14123 9158
rect 14140 9094 14204 9158
rect 14221 9094 14285 9158
rect 14302 9094 14366 9158
rect 14383 9094 14447 9158
rect 14464 9094 14528 9158
rect 14545 9094 14609 9158
rect 14626 9094 14690 9158
rect 14707 9094 14771 9158
rect 14788 9094 14852 9158
rect 10084 9008 10148 9072
rect 10166 9008 10230 9072
rect 10248 9008 10312 9072
rect 10330 9008 10394 9072
rect 10412 9008 10476 9072
rect 10494 9008 10558 9072
rect 10576 9008 10640 9072
rect 10657 9008 10721 9072
rect 10738 9008 10802 9072
rect 10819 9008 10883 9072
rect 10900 9008 10964 9072
rect 10981 9008 11045 9072
rect 11062 9008 11126 9072
rect 11143 9008 11207 9072
rect 11224 9008 11288 9072
rect 11305 9008 11369 9072
rect 11386 9008 11450 9072
rect 11467 9008 11531 9072
rect 11548 9008 11612 9072
rect 11629 9008 11693 9072
rect 11710 9008 11774 9072
rect 11791 9008 11855 9072
rect 11872 9008 11936 9072
rect 11953 9008 12017 9072
rect 12034 9008 12098 9072
rect 12115 9008 12179 9072
rect 12196 9008 12260 9072
rect 12277 9008 12341 9072
rect 12358 9008 12422 9072
rect 12439 9008 12503 9072
rect 12520 9008 12584 9072
rect 12601 9008 12665 9072
rect 12682 9008 12746 9072
rect 12763 9008 12827 9072
rect 12844 9008 12908 9072
rect 12925 9008 12989 9072
rect 13006 9008 13070 9072
rect 13087 9008 13151 9072
rect 13168 9008 13232 9072
rect 13249 9008 13313 9072
rect 13330 9008 13394 9072
rect 13411 9008 13475 9072
rect 13492 9008 13556 9072
rect 13573 9008 13637 9072
rect 13654 9008 13718 9072
rect 13735 9008 13799 9072
rect 13816 9008 13880 9072
rect 13897 9008 13961 9072
rect 13978 9008 14042 9072
rect 14059 9008 14123 9072
rect 14140 9008 14204 9072
rect 14221 9008 14285 9072
rect 14302 9008 14366 9072
rect 14383 9008 14447 9072
rect 14464 9008 14528 9072
rect 14545 9008 14609 9072
rect 14626 9008 14690 9072
rect 14707 9008 14771 9072
rect 14788 9008 14852 9072
rect 10084 8922 10148 8986
rect 10166 8922 10230 8986
rect 10248 8922 10312 8986
rect 10330 8922 10394 8986
rect 10412 8922 10476 8986
rect 10494 8922 10558 8986
rect 10576 8922 10640 8986
rect 10657 8922 10721 8986
rect 10738 8922 10802 8986
rect 10819 8922 10883 8986
rect 10900 8922 10964 8986
rect 10981 8922 11045 8986
rect 11062 8922 11126 8986
rect 11143 8922 11207 8986
rect 11224 8922 11288 8986
rect 11305 8922 11369 8986
rect 11386 8922 11450 8986
rect 11467 8922 11531 8986
rect 11548 8922 11612 8986
rect 11629 8922 11693 8986
rect 11710 8922 11774 8986
rect 11791 8922 11855 8986
rect 11872 8922 11936 8986
rect 11953 8922 12017 8986
rect 12034 8922 12098 8986
rect 12115 8922 12179 8986
rect 12196 8922 12260 8986
rect 12277 8922 12341 8986
rect 12358 8922 12422 8986
rect 12439 8922 12503 8986
rect 12520 8922 12584 8986
rect 12601 8922 12665 8986
rect 12682 8922 12746 8986
rect 12763 8922 12827 8986
rect 12844 8922 12908 8986
rect 12925 8922 12989 8986
rect 13006 8922 13070 8986
rect 13087 8922 13151 8986
rect 13168 8922 13232 8986
rect 13249 8922 13313 8986
rect 13330 8922 13394 8986
rect 13411 8922 13475 8986
rect 13492 8922 13556 8986
rect 13573 8922 13637 8986
rect 13654 8922 13718 8986
rect 13735 8922 13799 8986
rect 13816 8922 13880 8986
rect 13897 8922 13961 8986
rect 13978 8922 14042 8986
rect 14059 8922 14123 8986
rect 14140 8922 14204 8986
rect 14221 8922 14285 8986
rect 14302 8922 14366 8986
rect 14383 8922 14447 8986
rect 14464 8922 14528 8986
rect 14545 8922 14609 8986
rect 14626 8922 14690 8986
rect 14707 8922 14771 8986
rect 14788 8922 14852 8986
rect 10084 8836 10148 8900
rect 10166 8836 10230 8900
rect 10248 8836 10312 8900
rect 10330 8836 10394 8900
rect 10412 8836 10476 8900
rect 10494 8836 10558 8900
rect 10576 8836 10640 8900
rect 10657 8836 10721 8900
rect 10738 8836 10802 8900
rect 10819 8836 10883 8900
rect 10900 8836 10964 8900
rect 10981 8836 11045 8900
rect 11062 8836 11126 8900
rect 11143 8836 11207 8900
rect 11224 8836 11288 8900
rect 11305 8836 11369 8900
rect 11386 8836 11450 8900
rect 11467 8836 11531 8900
rect 11548 8836 11612 8900
rect 11629 8836 11693 8900
rect 11710 8836 11774 8900
rect 11791 8836 11855 8900
rect 11872 8836 11936 8900
rect 11953 8836 12017 8900
rect 12034 8836 12098 8900
rect 12115 8836 12179 8900
rect 12196 8836 12260 8900
rect 12277 8836 12341 8900
rect 12358 8836 12422 8900
rect 12439 8836 12503 8900
rect 12520 8836 12584 8900
rect 12601 8836 12665 8900
rect 12682 8836 12746 8900
rect 12763 8836 12827 8900
rect 12844 8836 12908 8900
rect 12925 8836 12989 8900
rect 13006 8836 13070 8900
rect 13087 8836 13151 8900
rect 13168 8836 13232 8900
rect 13249 8836 13313 8900
rect 13330 8836 13394 8900
rect 13411 8836 13475 8900
rect 13492 8836 13556 8900
rect 13573 8836 13637 8900
rect 13654 8836 13718 8900
rect 13735 8836 13799 8900
rect 13816 8836 13880 8900
rect 13897 8836 13961 8900
rect 13978 8836 14042 8900
rect 14059 8836 14123 8900
rect 14140 8836 14204 8900
rect 14221 8836 14285 8900
rect 14302 8836 14366 8900
rect 14383 8836 14447 8900
rect 14464 8836 14528 8900
rect 14545 8836 14609 8900
rect 14626 8836 14690 8900
rect 14707 8836 14771 8900
rect 14788 8836 14852 8900
rect 10084 8750 10148 8814
rect 10166 8750 10230 8814
rect 10248 8750 10312 8814
rect 10330 8750 10394 8814
rect 10412 8750 10476 8814
rect 10494 8750 10558 8814
rect 10576 8750 10640 8814
rect 10657 8750 10721 8814
rect 10738 8750 10802 8814
rect 10819 8750 10883 8814
rect 10900 8750 10964 8814
rect 10981 8750 11045 8814
rect 11062 8750 11126 8814
rect 11143 8750 11207 8814
rect 11224 8750 11288 8814
rect 11305 8750 11369 8814
rect 11386 8750 11450 8814
rect 11467 8750 11531 8814
rect 11548 8750 11612 8814
rect 11629 8750 11693 8814
rect 11710 8750 11774 8814
rect 11791 8750 11855 8814
rect 11872 8750 11936 8814
rect 11953 8750 12017 8814
rect 12034 8750 12098 8814
rect 12115 8750 12179 8814
rect 12196 8750 12260 8814
rect 12277 8750 12341 8814
rect 12358 8750 12422 8814
rect 12439 8750 12503 8814
rect 12520 8750 12584 8814
rect 12601 8750 12665 8814
rect 12682 8750 12746 8814
rect 12763 8750 12827 8814
rect 12844 8750 12908 8814
rect 12925 8750 12989 8814
rect 13006 8750 13070 8814
rect 13087 8750 13151 8814
rect 13168 8750 13232 8814
rect 13249 8750 13313 8814
rect 13330 8750 13394 8814
rect 13411 8750 13475 8814
rect 13492 8750 13556 8814
rect 13573 8750 13637 8814
rect 13654 8750 13718 8814
rect 13735 8750 13799 8814
rect 13816 8750 13880 8814
rect 13897 8750 13961 8814
rect 13978 8750 14042 8814
rect 14059 8750 14123 8814
rect 14140 8750 14204 8814
rect 14221 8750 14285 8814
rect 14302 8750 14366 8814
rect 14383 8750 14447 8814
rect 14464 8750 14528 8814
rect 14545 8750 14609 8814
rect 14626 8750 14690 8814
rect 14707 8750 14771 8814
rect 14788 8750 14852 8814
rect 10084 8664 10148 8728
rect 10166 8664 10230 8728
rect 10248 8664 10312 8728
rect 10330 8664 10394 8728
rect 10412 8664 10476 8728
rect 10494 8664 10558 8728
rect 10576 8664 10640 8728
rect 10657 8664 10721 8728
rect 10738 8664 10802 8728
rect 10819 8664 10883 8728
rect 10900 8664 10964 8728
rect 10981 8664 11045 8728
rect 11062 8664 11126 8728
rect 11143 8664 11207 8728
rect 11224 8664 11288 8728
rect 11305 8664 11369 8728
rect 11386 8664 11450 8728
rect 11467 8664 11531 8728
rect 11548 8664 11612 8728
rect 11629 8664 11693 8728
rect 11710 8664 11774 8728
rect 11791 8664 11855 8728
rect 11872 8664 11936 8728
rect 11953 8664 12017 8728
rect 12034 8664 12098 8728
rect 12115 8664 12179 8728
rect 12196 8664 12260 8728
rect 12277 8664 12341 8728
rect 12358 8664 12422 8728
rect 12439 8664 12503 8728
rect 12520 8664 12584 8728
rect 12601 8664 12665 8728
rect 12682 8664 12746 8728
rect 12763 8664 12827 8728
rect 12844 8664 12908 8728
rect 12925 8664 12989 8728
rect 13006 8664 13070 8728
rect 13087 8664 13151 8728
rect 13168 8664 13232 8728
rect 13249 8664 13313 8728
rect 13330 8664 13394 8728
rect 13411 8664 13475 8728
rect 13492 8664 13556 8728
rect 13573 8664 13637 8728
rect 13654 8664 13718 8728
rect 13735 8664 13799 8728
rect 13816 8664 13880 8728
rect 13897 8664 13961 8728
rect 13978 8664 14042 8728
rect 14059 8664 14123 8728
rect 14140 8664 14204 8728
rect 14221 8664 14285 8728
rect 14302 8664 14366 8728
rect 14383 8664 14447 8728
rect 14464 8664 14528 8728
rect 14545 8664 14609 8728
rect 14626 8664 14690 8728
rect 14707 8664 14771 8728
rect 14788 8664 14852 8728
rect 10084 8578 10148 8642
rect 10166 8578 10230 8642
rect 10248 8578 10312 8642
rect 10330 8578 10394 8642
rect 10412 8578 10476 8642
rect 10494 8578 10558 8642
rect 10576 8578 10640 8642
rect 10657 8578 10721 8642
rect 10738 8578 10802 8642
rect 10819 8578 10883 8642
rect 10900 8578 10964 8642
rect 10981 8578 11045 8642
rect 11062 8578 11126 8642
rect 11143 8578 11207 8642
rect 11224 8578 11288 8642
rect 11305 8578 11369 8642
rect 11386 8578 11450 8642
rect 11467 8578 11531 8642
rect 11548 8578 11612 8642
rect 11629 8578 11693 8642
rect 11710 8578 11774 8642
rect 11791 8578 11855 8642
rect 11872 8578 11936 8642
rect 11953 8578 12017 8642
rect 12034 8578 12098 8642
rect 12115 8578 12179 8642
rect 12196 8578 12260 8642
rect 12277 8578 12341 8642
rect 12358 8578 12422 8642
rect 12439 8578 12503 8642
rect 12520 8578 12584 8642
rect 12601 8578 12665 8642
rect 12682 8578 12746 8642
rect 12763 8578 12827 8642
rect 12844 8578 12908 8642
rect 12925 8578 12989 8642
rect 13006 8578 13070 8642
rect 13087 8578 13151 8642
rect 13168 8578 13232 8642
rect 13249 8578 13313 8642
rect 13330 8578 13394 8642
rect 13411 8578 13475 8642
rect 13492 8578 13556 8642
rect 13573 8578 13637 8642
rect 13654 8578 13718 8642
rect 13735 8578 13799 8642
rect 13816 8578 13880 8642
rect 13897 8578 13961 8642
rect 13978 8578 14042 8642
rect 14059 8578 14123 8642
rect 14140 8578 14204 8642
rect 14221 8578 14285 8642
rect 14302 8578 14366 8642
rect 14383 8578 14447 8642
rect 14464 8578 14528 8642
rect 14545 8578 14609 8642
rect 14626 8578 14690 8642
rect 14707 8578 14771 8642
rect 14788 8578 14852 8642
rect 10084 8492 10148 8556
rect 10166 8492 10230 8556
rect 10248 8492 10312 8556
rect 10330 8492 10394 8556
rect 10412 8492 10476 8556
rect 10494 8492 10558 8556
rect 10576 8492 10640 8556
rect 10657 8492 10721 8556
rect 10738 8492 10802 8556
rect 10819 8492 10883 8556
rect 10900 8492 10964 8556
rect 10981 8492 11045 8556
rect 11062 8492 11126 8556
rect 11143 8492 11207 8556
rect 11224 8492 11288 8556
rect 11305 8492 11369 8556
rect 11386 8492 11450 8556
rect 11467 8492 11531 8556
rect 11548 8492 11612 8556
rect 11629 8492 11693 8556
rect 11710 8492 11774 8556
rect 11791 8492 11855 8556
rect 11872 8492 11936 8556
rect 11953 8492 12017 8556
rect 12034 8492 12098 8556
rect 12115 8492 12179 8556
rect 12196 8492 12260 8556
rect 12277 8492 12341 8556
rect 12358 8492 12422 8556
rect 12439 8492 12503 8556
rect 12520 8492 12584 8556
rect 12601 8492 12665 8556
rect 12682 8492 12746 8556
rect 12763 8492 12827 8556
rect 12844 8492 12908 8556
rect 12925 8492 12989 8556
rect 13006 8492 13070 8556
rect 13087 8492 13151 8556
rect 13168 8492 13232 8556
rect 13249 8492 13313 8556
rect 13330 8492 13394 8556
rect 13411 8492 13475 8556
rect 13492 8492 13556 8556
rect 13573 8492 13637 8556
rect 13654 8492 13718 8556
rect 13735 8492 13799 8556
rect 13816 8492 13880 8556
rect 13897 8492 13961 8556
rect 13978 8492 14042 8556
rect 14059 8492 14123 8556
rect 14140 8492 14204 8556
rect 14221 8492 14285 8556
rect 14302 8492 14366 8556
rect 14383 8492 14447 8556
rect 14464 8492 14528 8556
rect 14545 8492 14609 8556
rect 14626 8492 14690 8556
rect 14707 8492 14771 8556
rect 14788 8492 14852 8556
rect 10084 8406 10148 8470
rect 10166 8406 10230 8470
rect 10248 8406 10312 8470
rect 10330 8406 10394 8470
rect 10412 8406 10476 8470
rect 10494 8406 10558 8470
rect 10576 8406 10640 8470
rect 10657 8406 10721 8470
rect 10738 8406 10802 8470
rect 10819 8406 10883 8470
rect 10900 8406 10964 8470
rect 10981 8406 11045 8470
rect 11062 8406 11126 8470
rect 11143 8406 11207 8470
rect 11224 8406 11288 8470
rect 11305 8406 11369 8470
rect 11386 8406 11450 8470
rect 11467 8406 11531 8470
rect 11548 8406 11612 8470
rect 11629 8406 11693 8470
rect 11710 8406 11774 8470
rect 11791 8406 11855 8470
rect 11872 8406 11936 8470
rect 11953 8406 12017 8470
rect 12034 8406 12098 8470
rect 12115 8406 12179 8470
rect 12196 8406 12260 8470
rect 12277 8406 12341 8470
rect 12358 8406 12422 8470
rect 12439 8406 12503 8470
rect 12520 8406 12584 8470
rect 12601 8406 12665 8470
rect 12682 8406 12746 8470
rect 12763 8406 12827 8470
rect 12844 8406 12908 8470
rect 12925 8406 12989 8470
rect 13006 8406 13070 8470
rect 13087 8406 13151 8470
rect 13168 8406 13232 8470
rect 13249 8406 13313 8470
rect 13330 8406 13394 8470
rect 13411 8406 13475 8470
rect 13492 8406 13556 8470
rect 13573 8406 13637 8470
rect 13654 8406 13718 8470
rect 13735 8406 13799 8470
rect 13816 8406 13880 8470
rect 13897 8406 13961 8470
rect 13978 8406 14042 8470
rect 14059 8406 14123 8470
rect 14140 8406 14204 8470
rect 14221 8406 14285 8470
rect 14302 8406 14366 8470
rect 14383 8406 14447 8470
rect 14464 8406 14528 8470
rect 14545 8406 14609 8470
rect 14626 8406 14690 8470
rect 14707 8406 14771 8470
rect 14788 8406 14852 8470
rect 10084 8320 10148 8384
rect 10166 8320 10230 8384
rect 10248 8320 10312 8384
rect 10330 8320 10394 8384
rect 10412 8320 10476 8384
rect 10494 8320 10558 8384
rect 10576 8320 10640 8384
rect 10657 8320 10721 8384
rect 10738 8320 10802 8384
rect 10819 8320 10883 8384
rect 10900 8320 10964 8384
rect 10981 8320 11045 8384
rect 11062 8320 11126 8384
rect 11143 8320 11207 8384
rect 11224 8320 11288 8384
rect 11305 8320 11369 8384
rect 11386 8320 11450 8384
rect 11467 8320 11531 8384
rect 11548 8320 11612 8384
rect 11629 8320 11693 8384
rect 11710 8320 11774 8384
rect 11791 8320 11855 8384
rect 11872 8320 11936 8384
rect 11953 8320 12017 8384
rect 12034 8320 12098 8384
rect 12115 8320 12179 8384
rect 12196 8320 12260 8384
rect 12277 8320 12341 8384
rect 12358 8320 12422 8384
rect 12439 8320 12503 8384
rect 12520 8320 12584 8384
rect 12601 8320 12665 8384
rect 12682 8320 12746 8384
rect 12763 8320 12827 8384
rect 12844 8320 12908 8384
rect 12925 8320 12989 8384
rect 13006 8320 13070 8384
rect 13087 8320 13151 8384
rect 13168 8320 13232 8384
rect 13249 8320 13313 8384
rect 13330 8320 13394 8384
rect 13411 8320 13475 8384
rect 13492 8320 13556 8384
rect 13573 8320 13637 8384
rect 13654 8320 13718 8384
rect 13735 8320 13799 8384
rect 13816 8320 13880 8384
rect 13897 8320 13961 8384
rect 13978 8320 14042 8384
rect 14059 8320 14123 8384
rect 14140 8320 14204 8384
rect 14221 8320 14285 8384
rect 14302 8320 14366 8384
rect 14383 8320 14447 8384
rect 14464 8320 14528 8384
rect 14545 8320 14609 8384
rect 14626 8320 14690 8384
rect 14707 8320 14771 8384
rect 14788 8320 14852 8384
<< metal4 >>
rect 0 35157 254 40000
rect 14746 35157 15000 40000
rect 0 14007 254 19000
rect 14746 14007 15000 19000
rect 0 12817 254 13707
rect 14746 12817 15000 13707
rect 0 11647 254 12537
rect 14746 11647 15000 12537
rect 0 11281 254 11347
rect 14746 11281 15000 11347
rect 0 10625 254 11221
rect 14746 10625 15000 11221
rect 0 10329 254 10565
rect 14746 10329 15000 10565
rect 0 9673 254 10269
rect 14746 9673 15000 10269
rect 0 9547 254 9613
rect 14746 9547 15000 9613
rect 0 9244 4874 9247
rect 0 9180 200 9244
rect 264 9180 281 9244
rect 345 9180 362 9244
rect 426 9180 443 9244
rect 507 9180 524 9244
rect 588 9180 605 9244
rect 669 9180 686 9244
rect 750 9180 767 9244
rect 831 9180 848 9244
rect 912 9180 929 9244
rect 993 9180 1010 9244
rect 1074 9180 1091 9244
rect 1155 9180 1172 9244
rect 1236 9180 1253 9244
rect 1317 9180 1334 9244
rect 1398 9180 1415 9244
rect 1479 9180 1496 9244
rect 1560 9180 1577 9244
rect 1641 9180 1658 9244
rect 1722 9180 1739 9244
rect 1803 9180 1820 9244
rect 1884 9180 1901 9244
rect 1965 9180 1982 9244
rect 2046 9180 2063 9244
rect 2127 9180 2144 9244
rect 2208 9180 2225 9244
rect 2289 9180 2306 9244
rect 2370 9180 2387 9244
rect 2451 9180 2468 9244
rect 2532 9180 2549 9244
rect 2613 9180 2630 9244
rect 2694 9180 2711 9244
rect 2775 9180 2792 9244
rect 2856 9180 2873 9244
rect 2937 9180 2954 9244
rect 3018 9180 3035 9244
rect 3099 9180 3116 9244
rect 3180 9180 3197 9244
rect 3261 9180 3278 9244
rect 3342 9180 3359 9244
rect 3423 9180 3440 9244
rect 3504 9180 3521 9244
rect 3585 9180 3602 9244
rect 3666 9180 3683 9244
rect 3747 9180 3764 9244
rect 3828 9180 3845 9244
rect 3909 9180 3926 9244
rect 3990 9180 4007 9244
rect 4071 9180 4088 9244
rect 4152 9180 4169 9244
rect 4233 9180 4249 9244
rect 4313 9180 4329 9244
rect 4393 9180 4409 9244
rect 4473 9180 4489 9244
rect 4553 9180 4569 9244
rect 4633 9180 4649 9244
rect 4713 9180 4729 9244
rect 4793 9180 4809 9244
rect 4873 9180 4874 9244
rect 0 9158 4874 9180
rect 0 9094 200 9158
rect 264 9094 281 9158
rect 345 9094 362 9158
rect 426 9094 443 9158
rect 507 9094 524 9158
rect 588 9094 605 9158
rect 669 9094 686 9158
rect 750 9094 767 9158
rect 831 9094 848 9158
rect 912 9094 929 9158
rect 993 9094 1010 9158
rect 1074 9094 1091 9158
rect 1155 9094 1172 9158
rect 1236 9094 1253 9158
rect 1317 9094 1334 9158
rect 1398 9094 1415 9158
rect 1479 9094 1496 9158
rect 1560 9094 1577 9158
rect 1641 9094 1658 9158
rect 1722 9094 1739 9158
rect 1803 9094 1820 9158
rect 1884 9094 1901 9158
rect 1965 9094 1982 9158
rect 2046 9094 2063 9158
rect 2127 9094 2144 9158
rect 2208 9094 2225 9158
rect 2289 9094 2306 9158
rect 2370 9094 2387 9158
rect 2451 9094 2468 9158
rect 2532 9094 2549 9158
rect 2613 9094 2630 9158
rect 2694 9094 2711 9158
rect 2775 9094 2792 9158
rect 2856 9094 2873 9158
rect 2937 9094 2954 9158
rect 3018 9094 3035 9158
rect 3099 9094 3116 9158
rect 3180 9094 3197 9158
rect 3261 9094 3278 9158
rect 3342 9094 3359 9158
rect 3423 9094 3440 9158
rect 3504 9094 3521 9158
rect 3585 9094 3602 9158
rect 3666 9094 3683 9158
rect 3747 9094 3764 9158
rect 3828 9094 3845 9158
rect 3909 9094 3926 9158
rect 3990 9094 4007 9158
rect 4071 9094 4088 9158
rect 4152 9094 4169 9158
rect 4233 9094 4249 9158
rect 4313 9094 4329 9158
rect 4393 9094 4409 9158
rect 4473 9094 4489 9158
rect 4553 9094 4569 9158
rect 4633 9094 4649 9158
rect 4713 9094 4729 9158
rect 4793 9094 4809 9158
rect 4873 9094 4874 9158
rect 0 9072 4874 9094
rect 0 9008 200 9072
rect 264 9008 281 9072
rect 345 9008 362 9072
rect 426 9008 443 9072
rect 507 9008 524 9072
rect 588 9008 605 9072
rect 669 9008 686 9072
rect 750 9008 767 9072
rect 831 9008 848 9072
rect 912 9008 929 9072
rect 993 9008 1010 9072
rect 1074 9008 1091 9072
rect 1155 9008 1172 9072
rect 1236 9008 1253 9072
rect 1317 9008 1334 9072
rect 1398 9008 1415 9072
rect 1479 9008 1496 9072
rect 1560 9008 1577 9072
rect 1641 9008 1658 9072
rect 1722 9008 1739 9072
rect 1803 9008 1820 9072
rect 1884 9008 1901 9072
rect 1965 9008 1982 9072
rect 2046 9008 2063 9072
rect 2127 9008 2144 9072
rect 2208 9008 2225 9072
rect 2289 9008 2306 9072
rect 2370 9008 2387 9072
rect 2451 9008 2468 9072
rect 2532 9008 2549 9072
rect 2613 9008 2630 9072
rect 2694 9008 2711 9072
rect 2775 9008 2792 9072
rect 2856 9008 2873 9072
rect 2937 9008 2954 9072
rect 3018 9008 3035 9072
rect 3099 9008 3116 9072
rect 3180 9008 3197 9072
rect 3261 9008 3278 9072
rect 3342 9008 3359 9072
rect 3423 9008 3440 9072
rect 3504 9008 3521 9072
rect 3585 9008 3602 9072
rect 3666 9008 3683 9072
rect 3747 9008 3764 9072
rect 3828 9008 3845 9072
rect 3909 9008 3926 9072
rect 3990 9008 4007 9072
rect 4071 9008 4088 9072
rect 4152 9008 4169 9072
rect 4233 9008 4249 9072
rect 4313 9008 4329 9072
rect 4393 9008 4409 9072
rect 4473 9008 4489 9072
rect 4553 9008 4569 9072
rect 4633 9008 4649 9072
rect 4713 9008 4729 9072
rect 4793 9008 4809 9072
rect 4873 9008 4874 9072
rect 0 8986 4874 9008
rect 0 8922 200 8986
rect 264 8922 281 8986
rect 345 8922 362 8986
rect 426 8922 443 8986
rect 507 8922 524 8986
rect 588 8922 605 8986
rect 669 8922 686 8986
rect 750 8922 767 8986
rect 831 8922 848 8986
rect 912 8922 929 8986
rect 993 8922 1010 8986
rect 1074 8922 1091 8986
rect 1155 8922 1172 8986
rect 1236 8922 1253 8986
rect 1317 8922 1334 8986
rect 1398 8922 1415 8986
rect 1479 8922 1496 8986
rect 1560 8922 1577 8986
rect 1641 8922 1658 8986
rect 1722 8922 1739 8986
rect 1803 8922 1820 8986
rect 1884 8922 1901 8986
rect 1965 8922 1982 8986
rect 2046 8922 2063 8986
rect 2127 8922 2144 8986
rect 2208 8922 2225 8986
rect 2289 8922 2306 8986
rect 2370 8922 2387 8986
rect 2451 8922 2468 8986
rect 2532 8922 2549 8986
rect 2613 8922 2630 8986
rect 2694 8922 2711 8986
rect 2775 8922 2792 8986
rect 2856 8922 2873 8986
rect 2937 8922 2954 8986
rect 3018 8922 3035 8986
rect 3099 8922 3116 8986
rect 3180 8922 3197 8986
rect 3261 8922 3278 8986
rect 3342 8922 3359 8986
rect 3423 8922 3440 8986
rect 3504 8922 3521 8986
rect 3585 8922 3602 8986
rect 3666 8922 3683 8986
rect 3747 8922 3764 8986
rect 3828 8922 3845 8986
rect 3909 8922 3926 8986
rect 3990 8922 4007 8986
rect 4071 8922 4088 8986
rect 4152 8922 4169 8986
rect 4233 8922 4249 8986
rect 4313 8922 4329 8986
rect 4393 8922 4409 8986
rect 4473 8922 4489 8986
rect 4553 8922 4569 8986
rect 4633 8922 4649 8986
rect 4713 8922 4729 8986
rect 4793 8922 4809 8986
rect 4873 8922 4874 8986
rect 0 8900 4874 8922
rect 0 8836 200 8900
rect 264 8836 281 8900
rect 345 8836 362 8900
rect 426 8836 443 8900
rect 507 8836 524 8900
rect 588 8836 605 8900
rect 669 8836 686 8900
rect 750 8836 767 8900
rect 831 8836 848 8900
rect 912 8836 929 8900
rect 993 8836 1010 8900
rect 1074 8836 1091 8900
rect 1155 8836 1172 8900
rect 1236 8836 1253 8900
rect 1317 8836 1334 8900
rect 1398 8836 1415 8900
rect 1479 8836 1496 8900
rect 1560 8836 1577 8900
rect 1641 8836 1658 8900
rect 1722 8836 1739 8900
rect 1803 8836 1820 8900
rect 1884 8836 1901 8900
rect 1965 8836 1982 8900
rect 2046 8836 2063 8900
rect 2127 8836 2144 8900
rect 2208 8836 2225 8900
rect 2289 8836 2306 8900
rect 2370 8836 2387 8900
rect 2451 8836 2468 8900
rect 2532 8836 2549 8900
rect 2613 8836 2630 8900
rect 2694 8836 2711 8900
rect 2775 8836 2792 8900
rect 2856 8836 2873 8900
rect 2937 8836 2954 8900
rect 3018 8836 3035 8900
rect 3099 8836 3116 8900
rect 3180 8836 3197 8900
rect 3261 8836 3278 8900
rect 3342 8836 3359 8900
rect 3423 8836 3440 8900
rect 3504 8836 3521 8900
rect 3585 8836 3602 8900
rect 3666 8836 3683 8900
rect 3747 8836 3764 8900
rect 3828 8836 3845 8900
rect 3909 8836 3926 8900
rect 3990 8836 4007 8900
rect 4071 8836 4088 8900
rect 4152 8836 4169 8900
rect 4233 8836 4249 8900
rect 4313 8836 4329 8900
rect 4393 8836 4409 8900
rect 4473 8836 4489 8900
rect 4553 8836 4569 8900
rect 4633 8836 4649 8900
rect 4713 8836 4729 8900
rect 4793 8836 4809 8900
rect 4873 8836 4874 8900
rect 0 8814 4874 8836
rect 0 8750 200 8814
rect 264 8750 281 8814
rect 345 8750 362 8814
rect 426 8750 443 8814
rect 507 8750 524 8814
rect 588 8750 605 8814
rect 669 8750 686 8814
rect 750 8750 767 8814
rect 831 8750 848 8814
rect 912 8750 929 8814
rect 993 8750 1010 8814
rect 1074 8750 1091 8814
rect 1155 8750 1172 8814
rect 1236 8750 1253 8814
rect 1317 8750 1334 8814
rect 1398 8750 1415 8814
rect 1479 8750 1496 8814
rect 1560 8750 1577 8814
rect 1641 8750 1658 8814
rect 1722 8750 1739 8814
rect 1803 8750 1820 8814
rect 1884 8750 1901 8814
rect 1965 8750 1982 8814
rect 2046 8750 2063 8814
rect 2127 8750 2144 8814
rect 2208 8750 2225 8814
rect 2289 8750 2306 8814
rect 2370 8750 2387 8814
rect 2451 8750 2468 8814
rect 2532 8750 2549 8814
rect 2613 8750 2630 8814
rect 2694 8750 2711 8814
rect 2775 8750 2792 8814
rect 2856 8750 2873 8814
rect 2937 8750 2954 8814
rect 3018 8750 3035 8814
rect 3099 8750 3116 8814
rect 3180 8750 3197 8814
rect 3261 8750 3278 8814
rect 3342 8750 3359 8814
rect 3423 8750 3440 8814
rect 3504 8750 3521 8814
rect 3585 8750 3602 8814
rect 3666 8750 3683 8814
rect 3747 8750 3764 8814
rect 3828 8750 3845 8814
rect 3909 8750 3926 8814
rect 3990 8750 4007 8814
rect 4071 8750 4088 8814
rect 4152 8750 4169 8814
rect 4233 8750 4249 8814
rect 4313 8750 4329 8814
rect 4393 8750 4409 8814
rect 4473 8750 4489 8814
rect 4553 8750 4569 8814
rect 4633 8750 4649 8814
rect 4713 8750 4729 8814
rect 4793 8750 4809 8814
rect 4873 8750 4874 8814
rect 0 8728 4874 8750
rect 0 8664 200 8728
rect 264 8664 281 8728
rect 345 8664 362 8728
rect 426 8664 443 8728
rect 507 8664 524 8728
rect 588 8664 605 8728
rect 669 8664 686 8728
rect 750 8664 767 8728
rect 831 8664 848 8728
rect 912 8664 929 8728
rect 993 8664 1010 8728
rect 1074 8664 1091 8728
rect 1155 8664 1172 8728
rect 1236 8664 1253 8728
rect 1317 8664 1334 8728
rect 1398 8664 1415 8728
rect 1479 8664 1496 8728
rect 1560 8664 1577 8728
rect 1641 8664 1658 8728
rect 1722 8664 1739 8728
rect 1803 8664 1820 8728
rect 1884 8664 1901 8728
rect 1965 8664 1982 8728
rect 2046 8664 2063 8728
rect 2127 8664 2144 8728
rect 2208 8664 2225 8728
rect 2289 8664 2306 8728
rect 2370 8664 2387 8728
rect 2451 8664 2468 8728
rect 2532 8664 2549 8728
rect 2613 8664 2630 8728
rect 2694 8664 2711 8728
rect 2775 8664 2792 8728
rect 2856 8664 2873 8728
rect 2937 8664 2954 8728
rect 3018 8664 3035 8728
rect 3099 8664 3116 8728
rect 3180 8664 3197 8728
rect 3261 8664 3278 8728
rect 3342 8664 3359 8728
rect 3423 8664 3440 8728
rect 3504 8664 3521 8728
rect 3585 8664 3602 8728
rect 3666 8664 3683 8728
rect 3747 8664 3764 8728
rect 3828 8664 3845 8728
rect 3909 8664 3926 8728
rect 3990 8664 4007 8728
rect 4071 8664 4088 8728
rect 4152 8664 4169 8728
rect 4233 8664 4249 8728
rect 4313 8664 4329 8728
rect 4393 8664 4409 8728
rect 4473 8664 4489 8728
rect 4553 8664 4569 8728
rect 4633 8664 4649 8728
rect 4713 8664 4729 8728
rect 4793 8664 4809 8728
rect 4873 8664 4874 8728
rect 0 8642 4874 8664
rect 0 8578 200 8642
rect 264 8578 281 8642
rect 345 8578 362 8642
rect 426 8578 443 8642
rect 507 8578 524 8642
rect 588 8578 605 8642
rect 669 8578 686 8642
rect 750 8578 767 8642
rect 831 8578 848 8642
rect 912 8578 929 8642
rect 993 8578 1010 8642
rect 1074 8578 1091 8642
rect 1155 8578 1172 8642
rect 1236 8578 1253 8642
rect 1317 8578 1334 8642
rect 1398 8578 1415 8642
rect 1479 8578 1496 8642
rect 1560 8578 1577 8642
rect 1641 8578 1658 8642
rect 1722 8578 1739 8642
rect 1803 8578 1820 8642
rect 1884 8578 1901 8642
rect 1965 8578 1982 8642
rect 2046 8578 2063 8642
rect 2127 8578 2144 8642
rect 2208 8578 2225 8642
rect 2289 8578 2306 8642
rect 2370 8578 2387 8642
rect 2451 8578 2468 8642
rect 2532 8578 2549 8642
rect 2613 8578 2630 8642
rect 2694 8578 2711 8642
rect 2775 8578 2792 8642
rect 2856 8578 2873 8642
rect 2937 8578 2954 8642
rect 3018 8578 3035 8642
rect 3099 8578 3116 8642
rect 3180 8578 3197 8642
rect 3261 8578 3278 8642
rect 3342 8578 3359 8642
rect 3423 8578 3440 8642
rect 3504 8578 3521 8642
rect 3585 8578 3602 8642
rect 3666 8578 3683 8642
rect 3747 8578 3764 8642
rect 3828 8578 3845 8642
rect 3909 8578 3926 8642
rect 3990 8578 4007 8642
rect 4071 8578 4088 8642
rect 4152 8578 4169 8642
rect 4233 8578 4249 8642
rect 4313 8578 4329 8642
rect 4393 8578 4409 8642
rect 4473 8578 4489 8642
rect 4553 8578 4569 8642
rect 4633 8578 4649 8642
rect 4713 8578 4729 8642
rect 4793 8578 4809 8642
rect 4873 8578 4874 8642
rect 0 8556 4874 8578
rect 0 8492 200 8556
rect 264 8492 281 8556
rect 345 8492 362 8556
rect 426 8492 443 8556
rect 507 8492 524 8556
rect 588 8492 605 8556
rect 669 8492 686 8556
rect 750 8492 767 8556
rect 831 8492 848 8556
rect 912 8492 929 8556
rect 993 8492 1010 8556
rect 1074 8492 1091 8556
rect 1155 8492 1172 8556
rect 1236 8492 1253 8556
rect 1317 8492 1334 8556
rect 1398 8492 1415 8556
rect 1479 8492 1496 8556
rect 1560 8492 1577 8556
rect 1641 8492 1658 8556
rect 1722 8492 1739 8556
rect 1803 8492 1820 8556
rect 1884 8492 1901 8556
rect 1965 8492 1982 8556
rect 2046 8492 2063 8556
rect 2127 8492 2144 8556
rect 2208 8492 2225 8556
rect 2289 8492 2306 8556
rect 2370 8492 2387 8556
rect 2451 8492 2468 8556
rect 2532 8492 2549 8556
rect 2613 8492 2630 8556
rect 2694 8492 2711 8556
rect 2775 8492 2792 8556
rect 2856 8492 2873 8556
rect 2937 8492 2954 8556
rect 3018 8492 3035 8556
rect 3099 8492 3116 8556
rect 3180 8492 3197 8556
rect 3261 8492 3278 8556
rect 3342 8492 3359 8556
rect 3423 8492 3440 8556
rect 3504 8492 3521 8556
rect 3585 8492 3602 8556
rect 3666 8492 3683 8556
rect 3747 8492 3764 8556
rect 3828 8492 3845 8556
rect 3909 8492 3926 8556
rect 3990 8492 4007 8556
rect 4071 8492 4088 8556
rect 4152 8492 4169 8556
rect 4233 8492 4249 8556
rect 4313 8492 4329 8556
rect 4393 8492 4409 8556
rect 4473 8492 4489 8556
rect 4553 8492 4569 8556
rect 4633 8492 4649 8556
rect 4713 8492 4729 8556
rect 4793 8492 4809 8556
rect 4873 8492 4874 8556
rect 0 8470 4874 8492
rect 0 8406 200 8470
rect 264 8406 281 8470
rect 345 8406 362 8470
rect 426 8406 443 8470
rect 507 8406 524 8470
rect 588 8406 605 8470
rect 669 8406 686 8470
rect 750 8406 767 8470
rect 831 8406 848 8470
rect 912 8406 929 8470
rect 993 8406 1010 8470
rect 1074 8406 1091 8470
rect 1155 8406 1172 8470
rect 1236 8406 1253 8470
rect 1317 8406 1334 8470
rect 1398 8406 1415 8470
rect 1479 8406 1496 8470
rect 1560 8406 1577 8470
rect 1641 8406 1658 8470
rect 1722 8406 1739 8470
rect 1803 8406 1820 8470
rect 1884 8406 1901 8470
rect 1965 8406 1982 8470
rect 2046 8406 2063 8470
rect 2127 8406 2144 8470
rect 2208 8406 2225 8470
rect 2289 8406 2306 8470
rect 2370 8406 2387 8470
rect 2451 8406 2468 8470
rect 2532 8406 2549 8470
rect 2613 8406 2630 8470
rect 2694 8406 2711 8470
rect 2775 8406 2792 8470
rect 2856 8406 2873 8470
rect 2937 8406 2954 8470
rect 3018 8406 3035 8470
rect 3099 8406 3116 8470
rect 3180 8406 3197 8470
rect 3261 8406 3278 8470
rect 3342 8406 3359 8470
rect 3423 8406 3440 8470
rect 3504 8406 3521 8470
rect 3585 8406 3602 8470
rect 3666 8406 3683 8470
rect 3747 8406 3764 8470
rect 3828 8406 3845 8470
rect 3909 8406 3926 8470
rect 3990 8406 4007 8470
rect 4071 8406 4088 8470
rect 4152 8406 4169 8470
rect 4233 8406 4249 8470
rect 4313 8406 4329 8470
rect 4393 8406 4409 8470
rect 4473 8406 4489 8470
rect 4553 8406 4569 8470
rect 4633 8406 4649 8470
rect 4713 8406 4729 8470
rect 4793 8406 4809 8470
rect 4873 8406 4874 8470
rect 0 8384 4874 8406
rect 0 8320 200 8384
rect 264 8320 281 8384
rect 345 8320 362 8384
rect 426 8320 443 8384
rect 507 8320 524 8384
rect 588 8320 605 8384
rect 669 8320 686 8384
rect 750 8320 767 8384
rect 831 8320 848 8384
rect 912 8320 929 8384
rect 993 8320 1010 8384
rect 1074 8320 1091 8384
rect 1155 8320 1172 8384
rect 1236 8320 1253 8384
rect 1317 8320 1334 8384
rect 1398 8320 1415 8384
rect 1479 8320 1496 8384
rect 1560 8320 1577 8384
rect 1641 8320 1658 8384
rect 1722 8320 1739 8384
rect 1803 8320 1820 8384
rect 1884 8320 1901 8384
rect 1965 8320 1982 8384
rect 2046 8320 2063 8384
rect 2127 8320 2144 8384
rect 2208 8320 2225 8384
rect 2289 8320 2306 8384
rect 2370 8320 2387 8384
rect 2451 8320 2468 8384
rect 2532 8320 2549 8384
rect 2613 8320 2630 8384
rect 2694 8320 2711 8384
rect 2775 8320 2792 8384
rect 2856 8320 2873 8384
rect 2937 8320 2954 8384
rect 3018 8320 3035 8384
rect 3099 8320 3116 8384
rect 3180 8320 3197 8384
rect 3261 8320 3278 8384
rect 3342 8320 3359 8384
rect 3423 8320 3440 8384
rect 3504 8320 3521 8384
rect 3585 8320 3602 8384
rect 3666 8320 3683 8384
rect 3747 8320 3764 8384
rect 3828 8320 3845 8384
rect 3909 8320 3926 8384
rect 3990 8320 4007 8384
rect 4071 8320 4088 8384
rect 4152 8320 4169 8384
rect 4233 8320 4249 8384
rect 4313 8320 4329 8384
rect 4393 8320 4409 8384
rect 4473 8320 4489 8384
rect 4553 8320 4569 8384
rect 4633 8320 4649 8384
rect 4713 8320 4729 8384
rect 4793 8320 4809 8384
rect 4873 8320 4874 8384
rect 0 8317 4874 8320
rect 10083 9244 15000 9247
rect 10083 9180 10084 9244
rect 10148 9180 10166 9244
rect 10230 9180 10248 9244
rect 10312 9180 10330 9244
rect 10394 9180 10412 9244
rect 10476 9180 10494 9244
rect 10558 9180 10576 9244
rect 10640 9180 10657 9244
rect 10721 9180 10738 9244
rect 10802 9180 10819 9244
rect 10883 9180 10900 9244
rect 10964 9180 10981 9244
rect 11045 9180 11062 9244
rect 11126 9180 11143 9244
rect 11207 9180 11224 9244
rect 11288 9180 11305 9244
rect 11369 9180 11386 9244
rect 11450 9180 11467 9244
rect 11531 9180 11548 9244
rect 11612 9180 11629 9244
rect 11693 9180 11710 9244
rect 11774 9180 11791 9244
rect 11855 9180 11872 9244
rect 11936 9180 11953 9244
rect 12017 9180 12034 9244
rect 12098 9180 12115 9244
rect 12179 9180 12196 9244
rect 12260 9180 12277 9244
rect 12341 9180 12358 9244
rect 12422 9180 12439 9244
rect 12503 9180 12520 9244
rect 12584 9180 12601 9244
rect 12665 9180 12682 9244
rect 12746 9180 12763 9244
rect 12827 9180 12844 9244
rect 12908 9180 12925 9244
rect 12989 9180 13006 9244
rect 13070 9180 13087 9244
rect 13151 9180 13168 9244
rect 13232 9180 13249 9244
rect 13313 9180 13330 9244
rect 13394 9180 13411 9244
rect 13475 9180 13492 9244
rect 13556 9180 13573 9244
rect 13637 9180 13654 9244
rect 13718 9180 13735 9244
rect 13799 9180 13816 9244
rect 13880 9180 13897 9244
rect 13961 9180 13978 9244
rect 14042 9180 14059 9244
rect 14123 9180 14140 9244
rect 14204 9180 14221 9244
rect 14285 9180 14302 9244
rect 14366 9180 14383 9244
rect 14447 9180 14464 9244
rect 14528 9180 14545 9244
rect 14609 9180 14626 9244
rect 14690 9180 14707 9244
rect 14771 9180 14788 9244
rect 14852 9180 15000 9244
rect 10083 9158 15000 9180
rect 10083 9094 10084 9158
rect 10148 9094 10166 9158
rect 10230 9094 10248 9158
rect 10312 9094 10330 9158
rect 10394 9094 10412 9158
rect 10476 9094 10494 9158
rect 10558 9094 10576 9158
rect 10640 9094 10657 9158
rect 10721 9094 10738 9158
rect 10802 9094 10819 9158
rect 10883 9094 10900 9158
rect 10964 9094 10981 9158
rect 11045 9094 11062 9158
rect 11126 9094 11143 9158
rect 11207 9094 11224 9158
rect 11288 9094 11305 9158
rect 11369 9094 11386 9158
rect 11450 9094 11467 9158
rect 11531 9094 11548 9158
rect 11612 9094 11629 9158
rect 11693 9094 11710 9158
rect 11774 9094 11791 9158
rect 11855 9094 11872 9158
rect 11936 9094 11953 9158
rect 12017 9094 12034 9158
rect 12098 9094 12115 9158
rect 12179 9094 12196 9158
rect 12260 9094 12277 9158
rect 12341 9094 12358 9158
rect 12422 9094 12439 9158
rect 12503 9094 12520 9158
rect 12584 9094 12601 9158
rect 12665 9094 12682 9158
rect 12746 9094 12763 9158
rect 12827 9094 12844 9158
rect 12908 9094 12925 9158
rect 12989 9094 13006 9158
rect 13070 9094 13087 9158
rect 13151 9094 13168 9158
rect 13232 9094 13249 9158
rect 13313 9094 13330 9158
rect 13394 9094 13411 9158
rect 13475 9094 13492 9158
rect 13556 9094 13573 9158
rect 13637 9094 13654 9158
rect 13718 9094 13735 9158
rect 13799 9094 13816 9158
rect 13880 9094 13897 9158
rect 13961 9094 13978 9158
rect 14042 9094 14059 9158
rect 14123 9094 14140 9158
rect 14204 9094 14221 9158
rect 14285 9094 14302 9158
rect 14366 9094 14383 9158
rect 14447 9094 14464 9158
rect 14528 9094 14545 9158
rect 14609 9094 14626 9158
rect 14690 9094 14707 9158
rect 14771 9094 14788 9158
rect 14852 9094 15000 9158
rect 10083 9072 15000 9094
rect 10083 9008 10084 9072
rect 10148 9008 10166 9072
rect 10230 9008 10248 9072
rect 10312 9008 10330 9072
rect 10394 9008 10412 9072
rect 10476 9008 10494 9072
rect 10558 9008 10576 9072
rect 10640 9008 10657 9072
rect 10721 9008 10738 9072
rect 10802 9008 10819 9072
rect 10883 9008 10900 9072
rect 10964 9008 10981 9072
rect 11045 9008 11062 9072
rect 11126 9008 11143 9072
rect 11207 9008 11224 9072
rect 11288 9008 11305 9072
rect 11369 9008 11386 9072
rect 11450 9008 11467 9072
rect 11531 9008 11548 9072
rect 11612 9008 11629 9072
rect 11693 9008 11710 9072
rect 11774 9008 11791 9072
rect 11855 9008 11872 9072
rect 11936 9008 11953 9072
rect 12017 9008 12034 9072
rect 12098 9008 12115 9072
rect 12179 9008 12196 9072
rect 12260 9008 12277 9072
rect 12341 9008 12358 9072
rect 12422 9008 12439 9072
rect 12503 9008 12520 9072
rect 12584 9008 12601 9072
rect 12665 9008 12682 9072
rect 12746 9008 12763 9072
rect 12827 9008 12844 9072
rect 12908 9008 12925 9072
rect 12989 9008 13006 9072
rect 13070 9008 13087 9072
rect 13151 9008 13168 9072
rect 13232 9008 13249 9072
rect 13313 9008 13330 9072
rect 13394 9008 13411 9072
rect 13475 9008 13492 9072
rect 13556 9008 13573 9072
rect 13637 9008 13654 9072
rect 13718 9008 13735 9072
rect 13799 9008 13816 9072
rect 13880 9008 13897 9072
rect 13961 9008 13978 9072
rect 14042 9008 14059 9072
rect 14123 9008 14140 9072
rect 14204 9008 14221 9072
rect 14285 9008 14302 9072
rect 14366 9008 14383 9072
rect 14447 9008 14464 9072
rect 14528 9008 14545 9072
rect 14609 9008 14626 9072
rect 14690 9008 14707 9072
rect 14771 9008 14788 9072
rect 14852 9008 15000 9072
rect 10083 8986 15000 9008
rect 10083 8922 10084 8986
rect 10148 8922 10166 8986
rect 10230 8922 10248 8986
rect 10312 8922 10330 8986
rect 10394 8922 10412 8986
rect 10476 8922 10494 8986
rect 10558 8922 10576 8986
rect 10640 8922 10657 8986
rect 10721 8922 10738 8986
rect 10802 8922 10819 8986
rect 10883 8922 10900 8986
rect 10964 8922 10981 8986
rect 11045 8922 11062 8986
rect 11126 8922 11143 8986
rect 11207 8922 11224 8986
rect 11288 8922 11305 8986
rect 11369 8922 11386 8986
rect 11450 8922 11467 8986
rect 11531 8922 11548 8986
rect 11612 8922 11629 8986
rect 11693 8922 11710 8986
rect 11774 8922 11791 8986
rect 11855 8922 11872 8986
rect 11936 8922 11953 8986
rect 12017 8922 12034 8986
rect 12098 8922 12115 8986
rect 12179 8922 12196 8986
rect 12260 8922 12277 8986
rect 12341 8922 12358 8986
rect 12422 8922 12439 8986
rect 12503 8922 12520 8986
rect 12584 8922 12601 8986
rect 12665 8922 12682 8986
rect 12746 8922 12763 8986
rect 12827 8922 12844 8986
rect 12908 8922 12925 8986
rect 12989 8922 13006 8986
rect 13070 8922 13087 8986
rect 13151 8922 13168 8986
rect 13232 8922 13249 8986
rect 13313 8922 13330 8986
rect 13394 8922 13411 8986
rect 13475 8922 13492 8986
rect 13556 8922 13573 8986
rect 13637 8922 13654 8986
rect 13718 8922 13735 8986
rect 13799 8922 13816 8986
rect 13880 8922 13897 8986
rect 13961 8922 13978 8986
rect 14042 8922 14059 8986
rect 14123 8922 14140 8986
rect 14204 8922 14221 8986
rect 14285 8922 14302 8986
rect 14366 8922 14383 8986
rect 14447 8922 14464 8986
rect 14528 8922 14545 8986
rect 14609 8922 14626 8986
rect 14690 8922 14707 8986
rect 14771 8922 14788 8986
rect 14852 8922 15000 8986
rect 10083 8900 15000 8922
rect 10083 8836 10084 8900
rect 10148 8836 10166 8900
rect 10230 8836 10248 8900
rect 10312 8836 10330 8900
rect 10394 8836 10412 8900
rect 10476 8836 10494 8900
rect 10558 8836 10576 8900
rect 10640 8836 10657 8900
rect 10721 8836 10738 8900
rect 10802 8836 10819 8900
rect 10883 8836 10900 8900
rect 10964 8836 10981 8900
rect 11045 8836 11062 8900
rect 11126 8836 11143 8900
rect 11207 8836 11224 8900
rect 11288 8836 11305 8900
rect 11369 8836 11386 8900
rect 11450 8836 11467 8900
rect 11531 8836 11548 8900
rect 11612 8836 11629 8900
rect 11693 8836 11710 8900
rect 11774 8836 11791 8900
rect 11855 8836 11872 8900
rect 11936 8836 11953 8900
rect 12017 8836 12034 8900
rect 12098 8836 12115 8900
rect 12179 8836 12196 8900
rect 12260 8836 12277 8900
rect 12341 8836 12358 8900
rect 12422 8836 12439 8900
rect 12503 8836 12520 8900
rect 12584 8836 12601 8900
rect 12665 8836 12682 8900
rect 12746 8836 12763 8900
rect 12827 8836 12844 8900
rect 12908 8836 12925 8900
rect 12989 8836 13006 8900
rect 13070 8836 13087 8900
rect 13151 8836 13168 8900
rect 13232 8836 13249 8900
rect 13313 8836 13330 8900
rect 13394 8836 13411 8900
rect 13475 8836 13492 8900
rect 13556 8836 13573 8900
rect 13637 8836 13654 8900
rect 13718 8836 13735 8900
rect 13799 8836 13816 8900
rect 13880 8836 13897 8900
rect 13961 8836 13978 8900
rect 14042 8836 14059 8900
rect 14123 8836 14140 8900
rect 14204 8836 14221 8900
rect 14285 8836 14302 8900
rect 14366 8836 14383 8900
rect 14447 8836 14464 8900
rect 14528 8836 14545 8900
rect 14609 8836 14626 8900
rect 14690 8836 14707 8900
rect 14771 8836 14788 8900
rect 14852 8836 15000 8900
rect 10083 8814 15000 8836
rect 10083 8750 10084 8814
rect 10148 8750 10166 8814
rect 10230 8750 10248 8814
rect 10312 8750 10330 8814
rect 10394 8750 10412 8814
rect 10476 8750 10494 8814
rect 10558 8750 10576 8814
rect 10640 8750 10657 8814
rect 10721 8750 10738 8814
rect 10802 8750 10819 8814
rect 10883 8750 10900 8814
rect 10964 8750 10981 8814
rect 11045 8750 11062 8814
rect 11126 8750 11143 8814
rect 11207 8750 11224 8814
rect 11288 8750 11305 8814
rect 11369 8750 11386 8814
rect 11450 8750 11467 8814
rect 11531 8750 11548 8814
rect 11612 8750 11629 8814
rect 11693 8750 11710 8814
rect 11774 8750 11791 8814
rect 11855 8750 11872 8814
rect 11936 8750 11953 8814
rect 12017 8750 12034 8814
rect 12098 8750 12115 8814
rect 12179 8750 12196 8814
rect 12260 8750 12277 8814
rect 12341 8750 12358 8814
rect 12422 8750 12439 8814
rect 12503 8750 12520 8814
rect 12584 8750 12601 8814
rect 12665 8750 12682 8814
rect 12746 8750 12763 8814
rect 12827 8750 12844 8814
rect 12908 8750 12925 8814
rect 12989 8750 13006 8814
rect 13070 8750 13087 8814
rect 13151 8750 13168 8814
rect 13232 8750 13249 8814
rect 13313 8750 13330 8814
rect 13394 8750 13411 8814
rect 13475 8750 13492 8814
rect 13556 8750 13573 8814
rect 13637 8750 13654 8814
rect 13718 8750 13735 8814
rect 13799 8750 13816 8814
rect 13880 8750 13897 8814
rect 13961 8750 13978 8814
rect 14042 8750 14059 8814
rect 14123 8750 14140 8814
rect 14204 8750 14221 8814
rect 14285 8750 14302 8814
rect 14366 8750 14383 8814
rect 14447 8750 14464 8814
rect 14528 8750 14545 8814
rect 14609 8750 14626 8814
rect 14690 8750 14707 8814
rect 14771 8750 14788 8814
rect 14852 8750 15000 8814
rect 10083 8728 15000 8750
rect 10083 8664 10084 8728
rect 10148 8664 10166 8728
rect 10230 8664 10248 8728
rect 10312 8664 10330 8728
rect 10394 8664 10412 8728
rect 10476 8664 10494 8728
rect 10558 8664 10576 8728
rect 10640 8664 10657 8728
rect 10721 8664 10738 8728
rect 10802 8664 10819 8728
rect 10883 8664 10900 8728
rect 10964 8664 10981 8728
rect 11045 8664 11062 8728
rect 11126 8664 11143 8728
rect 11207 8664 11224 8728
rect 11288 8664 11305 8728
rect 11369 8664 11386 8728
rect 11450 8664 11467 8728
rect 11531 8664 11548 8728
rect 11612 8664 11629 8728
rect 11693 8664 11710 8728
rect 11774 8664 11791 8728
rect 11855 8664 11872 8728
rect 11936 8664 11953 8728
rect 12017 8664 12034 8728
rect 12098 8664 12115 8728
rect 12179 8664 12196 8728
rect 12260 8664 12277 8728
rect 12341 8664 12358 8728
rect 12422 8664 12439 8728
rect 12503 8664 12520 8728
rect 12584 8664 12601 8728
rect 12665 8664 12682 8728
rect 12746 8664 12763 8728
rect 12827 8664 12844 8728
rect 12908 8664 12925 8728
rect 12989 8664 13006 8728
rect 13070 8664 13087 8728
rect 13151 8664 13168 8728
rect 13232 8664 13249 8728
rect 13313 8664 13330 8728
rect 13394 8664 13411 8728
rect 13475 8664 13492 8728
rect 13556 8664 13573 8728
rect 13637 8664 13654 8728
rect 13718 8664 13735 8728
rect 13799 8664 13816 8728
rect 13880 8664 13897 8728
rect 13961 8664 13978 8728
rect 14042 8664 14059 8728
rect 14123 8664 14140 8728
rect 14204 8664 14221 8728
rect 14285 8664 14302 8728
rect 14366 8664 14383 8728
rect 14447 8664 14464 8728
rect 14528 8664 14545 8728
rect 14609 8664 14626 8728
rect 14690 8664 14707 8728
rect 14771 8664 14788 8728
rect 14852 8664 15000 8728
rect 10083 8642 15000 8664
rect 10083 8578 10084 8642
rect 10148 8578 10166 8642
rect 10230 8578 10248 8642
rect 10312 8578 10330 8642
rect 10394 8578 10412 8642
rect 10476 8578 10494 8642
rect 10558 8578 10576 8642
rect 10640 8578 10657 8642
rect 10721 8578 10738 8642
rect 10802 8578 10819 8642
rect 10883 8578 10900 8642
rect 10964 8578 10981 8642
rect 11045 8578 11062 8642
rect 11126 8578 11143 8642
rect 11207 8578 11224 8642
rect 11288 8578 11305 8642
rect 11369 8578 11386 8642
rect 11450 8578 11467 8642
rect 11531 8578 11548 8642
rect 11612 8578 11629 8642
rect 11693 8578 11710 8642
rect 11774 8578 11791 8642
rect 11855 8578 11872 8642
rect 11936 8578 11953 8642
rect 12017 8578 12034 8642
rect 12098 8578 12115 8642
rect 12179 8578 12196 8642
rect 12260 8578 12277 8642
rect 12341 8578 12358 8642
rect 12422 8578 12439 8642
rect 12503 8578 12520 8642
rect 12584 8578 12601 8642
rect 12665 8578 12682 8642
rect 12746 8578 12763 8642
rect 12827 8578 12844 8642
rect 12908 8578 12925 8642
rect 12989 8578 13006 8642
rect 13070 8578 13087 8642
rect 13151 8578 13168 8642
rect 13232 8578 13249 8642
rect 13313 8578 13330 8642
rect 13394 8578 13411 8642
rect 13475 8578 13492 8642
rect 13556 8578 13573 8642
rect 13637 8578 13654 8642
rect 13718 8578 13735 8642
rect 13799 8578 13816 8642
rect 13880 8578 13897 8642
rect 13961 8578 13978 8642
rect 14042 8578 14059 8642
rect 14123 8578 14140 8642
rect 14204 8578 14221 8642
rect 14285 8578 14302 8642
rect 14366 8578 14383 8642
rect 14447 8578 14464 8642
rect 14528 8578 14545 8642
rect 14609 8578 14626 8642
rect 14690 8578 14707 8642
rect 14771 8578 14788 8642
rect 14852 8578 15000 8642
rect 10083 8556 15000 8578
rect 10083 8492 10084 8556
rect 10148 8492 10166 8556
rect 10230 8492 10248 8556
rect 10312 8492 10330 8556
rect 10394 8492 10412 8556
rect 10476 8492 10494 8556
rect 10558 8492 10576 8556
rect 10640 8492 10657 8556
rect 10721 8492 10738 8556
rect 10802 8492 10819 8556
rect 10883 8492 10900 8556
rect 10964 8492 10981 8556
rect 11045 8492 11062 8556
rect 11126 8492 11143 8556
rect 11207 8492 11224 8556
rect 11288 8492 11305 8556
rect 11369 8492 11386 8556
rect 11450 8492 11467 8556
rect 11531 8492 11548 8556
rect 11612 8492 11629 8556
rect 11693 8492 11710 8556
rect 11774 8492 11791 8556
rect 11855 8492 11872 8556
rect 11936 8492 11953 8556
rect 12017 8492 12034 8556
rect 12098 8492 12115 8556
rect 12179 8492 12196 8556
rect 12260 8492 12277 8556
rect 12341 8492 12358 8556
rect 12422 8492 12439 8556
rect 12503 8492 12520 8556
rect 12584 8492 12601 8556
rect 12665 8492 12682 8556
rect 12746 8492 12763 8556
rect 12827 8492 12844 8556
rect 12908 8492 12925 8556
rect 12989 8492 13006 8556
rect 13070 8492 13087 8556
rect 13151 8492 13168 8556
rect 13232 8492 13249 8556
rect 13313 8492 13330 8556
rect 13394 8492 13411 8556
rect 13475 8492 13492 8556
rect 13556 8492 13573 8556
rect 13637 8492 13654 8556
rect 13718 8492 13735 8556
rect 13799 8492 13816 8556
rect 13880 8492 13897 8556
rect 13961 8492 13978 8556
rect 14042 8492 14059 8556
rect 14123 8492 14140 8556
rect 14204 8492 14221 8556
rect 14285 8492 14302 8556
rect 14366 8492 14383 8556
rect 14447 8492 14464 8556
rect 14528 8492 14545 8556
rect 14609 8492 14626 8556
rect 14690 8492 14707 8556
rect 14771 8492 14788 8556
rect 14852 8492 15000 8556
rect 10083 8470 15000 8492
rect 10083 8406 10084 8470
rect 10148 8406 10166 8470
rect 10230 8406 10248 8470
rect 10312 8406 10330 8470
rect 10394 8406 10412 8470
rect 10476 8406 10494 8470
rect 10558 8406 10576 8470
rect 10640 8406 10657 8470
rect 10721 8406 10738 8470
rect 10802 8406 10819 8470
rect 10883 8406 10900 8470
rect 10964 8406 10981 8470
rect 11045 8406 11062 8470
rect 11126 8406 11143 8470
rect 11207 8406 11224 8470
rect 11288 8406 11305 8470
rect 11369 8406 11386 8470
rect 11450 8406 11467 8470
rect 11531 8406 11548 8470
rect 11612 8406 11629 8470
rect 11693 8406 11710 8470
rect 11774 8406 11791 8470
rect 11855 8406 11872 8470
rect 11936 8406 11953 8470
rect 12017 8406 12034 8470
rect 12098 8406 12115 8470
rect 12179 8406 12196 8470
rect 12260 8406 12277 8470
rect 12341 8406 12358 8470
rect 12422 8406 12439 8470
rect 12503 8406 12520 8470
rect 12584 8406 12601 8470
rect 12665 8406 12682 8470
rect 12746 8406 12763 8470
rect 12827 8406 12844 8470
rect 12908 8406 12925 8470
rect 12989 8406 13006 8470
rect 13070 8406 13087 8470
rect 13151 8406 13168 8470
rect 13232 8406 13249 8470
rect 13313 8406 13330 8470
rect 13394 8406 13411 8470
rect 13475 8406 13492 8470
rect 13556 8406 13573 8470
rect 13637 8406 13654 8470
rect 13718 8406 13735 8470
rect 13799 8406 13816 8470
rect 13880 8406 13897 8470
rect 13961 8406 13978 8470
rect 14042 8406 14059 8470
rect 14123 8406 14140 8470
rect 14204 8406 14221 8470
rect 14285 8406 14302 8470
rect 14366 8406 14383 8470
rect 14447 8406 14464 8470
rect 14528 8406 14545 8470
rect 14609 8406 14626 8470
rect 14690 8406 14707 8470
rect 14771 8406 14788 8470
rect 14852 8406 15000 8470
rect 10083 8384 15000 8406
rect 10083 8320 10084 8384
rect 10148 8320 10166 8384
rect 10230 8320 10248 8384
rect 10312 8320 10330 8384
rect 10394 8320 10412 8384
rect 10476 8320 10494 8384
rect 10558 8320 10576 8384
rect 10640 8320 10657 8384
rect 10721 8320 10738 8384
rect 10802 8320 10819 8384
rect 10883 8320 10900 8384
rect 10964 8320 10981 8384
rect 11045 8320 11062 8384
rect 11126 8320 11143 8384
rect 11207 8320 11224 8384
rect 11288 8320 11305 8384
rect 11369 8320 11386 8384
rect 11450 8320 11467 8384
rect 11531 8320 11548 8384
rect 11612 8320 11629 8384
rect 11693 8320 11710 8384
rect 11774 8320 11791 8384
rect 11855 8320 11872 8384
rect 11936 8320 11953 8384
rect 12017 8320 12034 8384
rect 12098 8320 12115 8384
rect 12179 8320 12196 8384
rect 12260 8320 12277 8384
rect 12341 8320 12358 8384
rect 12422 8320 12439 8384
rect 12503 8320 12520 8384
rect 12584 8320 12601 8384
rect 12665 8320 12682 8384
rect 12746 8320 12763 8384
rect 12827 8320 12844 8384
rect 12908 8320 12925 8384
rect 12989 8320 13006 8384
rect 13070 8320 13087 8384
rect 13151 8320 13168 8384
rect 13232 8320 13249 8384
rect 13313 8320 13330 8384
rect 13394 8320 13411 8384
rect 13475 8320 13492 8384
rect 13556 8320 13573 8384
rect 13637 8320 13654 8384
rect 13718 8320 13735 8384
rect 13799 8320 13816 8384
rect 13880 8320 13897 8384
rect 13961 8320 13978 8384
rect 14042 8320 14059 8384
rect 14123 8320 14140 8384
rect 14204 8320 14221 8384
rect 14285 8320 14302 8384
rect 14366 8320 14383 8384
rect 14447 8320 14464 8384
rect 14528 8320 14545 8384
rect 14609 8320 14626 8384
rect 14690 8320 14707 8384
rect 14771 8320 14788 8384
rect 14852 8320 15000 8384
rect 10083 8317 15000 8320
rect 0 7347 254 8037
rect 14746 7347 15000 8037
rect 0 6377 254 7067
rect 14746 6377 15000 7067
rect 0 5167 254 6097
rect 14746 5167 15000 6097
rect 0 3957 254 4887
rect 14746 3957 15000 4887
rect 0 2987 193 3677
rect 14807 2987 15000 3677
rect 0 1777 254 2707
rect 14746 1777 15000 2707
rect 0 407 254 1497
rect 14746 407 15000 1497
<< metal5 >>
rect 0 35157 254 40000
rect 14746 35157 15000 40000
rect 0 14007 254 18997
rect 14746 14007 15000 18997
rect 0 12837 254 13687
rect 14746 12837 15000 13687
rect 0 11667 254 12517
rect 14746 11667 15000 12517
rect 0 9547 254 11347
rect 14746 9547 15000 11347
rect 0 8337 254 9227
rect 14746 8337 15000 9227
rect 0 7368 254 8017
rect 14746 7368 15000 8017
rect 0 6397 254 7047
rect 14746 6397 15000 7047
rect 0 5187 254 6077
rect 14746 5187 15000 6077
rect 0 3977 254 4867
rect 14746 3977 15000 4867
rect 0 3007 193 3657
rect 14807 3007 15000 3657
rect 0 1797 254 2687
rect 14746 1797 15000 2687
rect 0 427 254 1477
rect 14746 427 15000 1477
use sky130_fd_io__com_bus_hookup  sky130_fd_io__com_bus_hookup_0
timestamp 1649977179
transform 1 0 0 0 1 549
box 0 -142 15000 39451
<< labels >>
flabel metal5 s 0 12837 254 13687 3 FreeSans 520 0 0 0 VDDIO_Q
port 1 nsew power bidirectional
flabel metal5 s 14746 1797 15000 2687 3 FreeSans 520 180 0 0 VCCD
port 2 nsew power bidirectional
flabel metal5 s 14746 9547 15000 11347 3 FreeSans 520 180 0 0 VSSA
port 3 nsew ground bidirectional
flabel metal5 s 14746 7368 15000 8017 3 FreeSans 520 180 0 0 VSSA
port 3 nsew ground bidirectional
flabel metal5 s 0 9547 254 11347 3 FreeSans 520 0 0 0 VSSA
port 3 nsew ground bidirectional
flabel metal5 s 0 7368 254 8017 3 FreeSans 520 0 0 0 VSSA
port 3 nsew ground bidirectional
flabel metal5 s 14746 8337 15000 9227 3 FreeSans 520 180 0 0 VSSD
port 4 nsew ground bidirectional
flabel metal5 s 0 8337 254 9227 3 FreeSans 520 0 0 0 VSSD
port 4 nsew ground bidirectional
flabel metal5 s 14746 35157 15000 40000 3 FreeSans 520 180 0 0 VSSIO
port 5 nsew ground bidirectional
flabel metal5 s 14746 5187 15000 6077 3 FreeSans 520 180 0 0 VSSIO
port 5 nsew ground bidirectional
flabel metal5 s 0 35157 254 40000 3 FreeSans 520 0 0 0 VSSIO
port 5 nsew ground bidirectional
flabel metal5 s 0 5187 254 6077 3 FreeSans 520 0 0 0 VSSIO
port 5 nsew ground bidirectional
flabel metal5 s 14746 11667 15000 12517 3 FreeSans 520 180 0 0 VSSIO_Q
port 6 nsew ground bidirectional
flabel metal5 s 0 11667 254 12517 3 FreeSans 520 0 0 0 VSSIO_Q
port 6 nsew ground bidirectional
flabel metal5 s 14746 6397 15000 7047 3 FreeSans 520 180 0 0 VSWITCH
port 7 nsew power bidirectional
flabel metal5 s 0 1797 254 2687 3 FreeSans 520 0 0 0 VCCD
port 2 nsew power bidirectional
flabel metal5 s 14746 427 15000 1477 3 FreeSans 520 180 0 0 VCCHIB
port 8 nsew power bidirectional
flabel metal5 s 0 427 254 1477 3 FreeSans 520 0 0 0 VCCHIB
port 8 nsew power bidirectional
flabel metal5 s 14807 3007 15000 3657 3 FreeSans 520 180 0 0 VDDA
port 9 nsew power bidirectional
flabel metal5 s 0 3007 193 3657 3 FreeSans 520 0 0 0 VDDA
port 9 nsew power bidirectional
flabel metal5 s 14746 14007 15000 18997 3 FreeSans 520 180 0 0 VDDIO
port 10 nsew power bidirectional
flabel metal5 s 14746 3977 15000 4867 3 FreeSans 520 180 0 0 VDDIO
port 10 nsew power bidirectional
flabel metal5 s 0 14007 254 18997 3 FreeSans 520 0 0 0 VDDIO
port 10 nsew power bidirectional
flabel metal5 s 0 3977 254 4867 3 FreeSans 520 0 0 0 VDDIO
port 10 nsew power bidirectional
flabel metal5 s 0 6397 254 7047 3 FreeSans 520 0 0 0 VSWITCH
port 7 nsew power bidirectional
flabel metal5 s 14746 12837 15000 13687 3 FreeSans 520 180 0 0 VDDIO_Q
port 1 nsew power bidirectional
flabel metal4 s 14746 7347 15000 8037 3 FreeSans 520 180 0 0 VSSA
port 3 nsew ground bidirectional
flabel metal4 s 14746 9547 15000 9613 3 FreeSans 520 180 0 0 VSSA
port 3 nsew ground bidirectional
flabel metal4 s 14746 11281 15000 11347 3 FreeSans 520 180 0 0 VSSA
port 3 nsew ground bidirectional
flabel metal4 s 14746 10329 15000 10565 3 FreeSans 520 180 0 0 VSSA
port 3 nsew ground bidirectional
flabel metal4 s 0 9547 254 9613 3 FreeSans 520 0 0 0 VSSA
port 3 nsew ground bidirectional
flabel metal4 s 0 407 254 1497 3 FreeSans 520 0 0 0 VCCHIB
port 8 nsew power bidirectional
flabel metal4 s 0 10329 254 10565 3 FreeSans 520 0 0 0 VSSA
port 3 nsew ground bidirectional
flabel metal4 s 0 11281 254 11347 3 FreeSans 520 0 0 0 VSSA
port 3 nsew ground bidirectional
flabel metal4 s 0 7347 254 8037 3 FreeSans 520 0 0 0 VSSA
port 3 nsew ground bidirectional
flabel metal4 s 14746 8317 15000 9247 3 FreeSans 520 180 0 0 VSSD
port 4 nsew ground bidirectional
flabel metal4 s 0 8317 254 9247 3 FreeSans 520 0 0 0 VSSD
port 4 nsew ground bidirectional
flabel metal4 s 14746 35157 15000 40000 3 FreeSans 520 180 0 0 VSSIO
port 5 nsew ground bidirectional
flabel metal4 s 14746 5167 15000 6097 3 FreeSans 520 180 0 0 VSSIO
port 5 nsew ground bidirectional
flabel metal4 s 0 35157 254 40000 3 FreeSans 520 0 0 0 VSSIO
port 5 nsew ground bidirectional
flabel metal4 s 0 5167 254 6097 3 FreeSans 520 0 0 0 VSSIO
port 5 nsew ground bidirectional
flabel metal4 s 14746 11647 15000 12537 3 FreeSans 520 180 0 0 VSSIO_Q
port 6 nsew ground bidirectional
flabel metal4 s 0 11647 254 12537 3 FreeSans 520 0 0 0 VSSIO_Q
port 6 nsew ground bidirectional
flabel metal4 s 14746 6377 15000 7067 3 FreeSans 520 180 0 0 VSWITCH
port 7 nsew power bidirectional
flabel metal4 s 14746 10625 15000 11221 3 FreeSans 520 180 0 0 AMUXBUS_A
port 11 nsew signal bidirectional
flabel metal4 s 0 10625 254 11221 3 FreeSans 520 0 0 0 AMUXBUS_A
port 11 nsew signal bidirectional
flabel metal4 s 14746 9673 15000 10269 3 FreeSans 520 180 0 0 AMUXBUS_B
port 12 nsew signal bidirectional
flabel metal4 s 0 9673 254 10269 3 FreeSans 520 0 0 0 AMUXBUS_B
port 12 nsew signal bidirectional
flabel metal4 s 14746 1777 15000 2707 3 FreeSans 520 180 0 0 VCCD
port 2 nsew power bidirectional
flabel metal4 s 0 1777 254 2707 3 FreeSans 520 0 0 0 VCCD
port 2 nsew power bidirectional
flabel metal4 s 14746 407 15000 1497 3 FreeSans 520 180 0 0 VCCHIB
port 8 nsew power bidirectional
flabel metal4 s 14807 2987 15000 3677 3 FreeSans 520 180 0 0 VDDA
port 9 nsew power bidirectional
flabel metal4 s 0 2987 193 3677 3 FreeSans 520 0 0 0 VDDA
port 9 nsew power bidirectional
flabel metal4 s 14746 3957 15000 4887 3 FreeSans 520 180 0 0 VDDIO
port 10 nsew power bidirectional
flabel metal4 s 14746 14007 15000 19000 3 FreeSans 520 180 0 0 VDDIO
port 10 nsew power bidirectional
flabel metal4 s 0 3957 254 4887 3 FreeSans 520 0 0 0 VDDIO
port 10 nsew power bidirectional
flabel metal4 s 0 14007 254 19000 3 FreeSans 520 0 0 0 VDDIO
port 10 nsew power bidirectional
flabel metal4 s 14746 12817 15000 13707 3 FreeSans 520 180 0 0 VDDIO_Q
port 1 nsew power bidirectional
flabel metal4 s 0 6377 254 7067 3 FreeSans 520 0 0 0 VSWITCH
port 7 nsew power bidirectional
flabel metal4 s 0 12817 254 13707 3 FreeSans 520 0 0 0 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 14746 10625 15000 11221 1 AMUXBUS_A
port 11 nsew signal bidirectional
rlabel metal4 s 14746 9673 15000 10269 1 AMUXBUS_B
port 12 nsew signal bidirectional
rlabel metal4 s 14746 1777 15000 2707 1 VCCD
port 2 nsew power bidirectional
rlabel metal5 s 0 1797 254 2687 1 VCCD
port 2 nsew power bidirectional
rlabel metal5 s 14746 1797 15000 2687 1 VCCD
port 2 nsew power bidirectional
rlabel metal4 s 14746 407 15000 1497 1 VCCHIB
port 8 nsew power bidirectional
rlabel metal5 s 0 427 254 1477 1 VCCHIB
port 8 nsew power bidirectional
rlabel metal5 s 14746 427 15000 1477 1 VCCHIB
port 8 nsew power bidirectional
rlabel metal4 s 14807 2987 15000 3677 1 VDDA
port 9 nsew power bidirectional
rlabel metal5 s 0 3007 193 3657 1 VDDA
port 9 nsew power bidirectional
rlabel metal5 s 14807 3007 15000 3657 1 VDDA
port 9 nsew power bidirectional
rlabel metal4 s 0 14007 254 19000 1 VDDIO
port 10 nsew power bidirectional
rlabel metal4 s 14746 3957 15000 4887 1 VDDIO
port 10 nsew power bidirectional
rlabel metal4 s 14746 14007 15000 19000 1 VDDIO
port 10 nsew power bidirectional
rlabel metal5 s 0 3977 254 4867 1 VDDIO
port 10 nsew power bidirectional
rlabel metal5 s 0 14007 254 18997 1 VDDIO
port 10 nsew power bidirectional
rlabel metal5 s 14746 3977 15000 4867 1 VDDIO
port 10 nsew power bidirectional
rlabel metal5 s 14746 14007 15000 18997 1 VDDIO
port 10 nsew power bidirectional
rlabel metal4 s 14746 12817 15000 13707 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal5 s 0 12837 254 13687 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal5 s 14746 12837 15000 13687 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 0 9547 254 9613 1 VSSA
port 3 nsew ground bidirectional
rlabel metal4 s 0 10329 254 10565 1 VSSA
port 3 nsew ground bidirectional
rlabel metal4 s 0 11281 254 11347 1 VSSA
port 3 nsew ground bidirectional
rlabel metal4 s 14746 7347 15000 8037 1 VSSA
port 3 nsew ground bidirectional
rlabel metal4 s 14746 9547 15000 9613 1 VSSA
port 3 nsew ground bidirectional
rlabel metal4 s 14746 10329 15000 10565 1 VSSA
port 3 nsew ground bidirectional
rlabel metal4 s 14746 11281 15000 11347 1 VSSA
port 3 nsew ground bidirectional
rlabel metal5 s 0 7368 254 8017 1 VSSA
port 3 nsew ground bidirectional
rlabel metal5 s 0 9547 254 11347 1 VSSA
port 3 nsew ground bidirectional
rlabel metal5 s 14746 7368 15000 8017 1 VSSA
port 3 nsew ground bidirectional
rlabel metal5 s 14746 9547 15000 11347 1 VSSA
port 3 nsew ground bidirectional
rlabel metal3 s 10078 8318 14858 9246 1 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 0 8317 4874 9247 1 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 10083 8317 15000 9247 1 VSSD
port 4 nsew ground bidirectional
rlabel metal5 s 0 8337 254 9227 1 VSSD
port 4 nsew ground bidirectional
rlabel metal5 s 14746 8337 15000 9227 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 14800 9192 14840 9232 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 14800 9106 14840 9146 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 14800 9020 14840 9060 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 14800 8934 14840 8974 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 14800 8848 14840 8888 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 14800 8762 14840 8802 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 14800 8676 14840 8716 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 14800 8590 14840 8630 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 14800 8504 14840 8544 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 14800 8418 14840 8458 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 14800 8332 14840 8372 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 14719 9192 14759 9232 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 14719 9106 14759 9146 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 14719 9020 14759 9060 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 14719 8934 14759 8974 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 14719 8848 14759 8888 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 14719 8762 14759 8802 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 14719 8676 14759 8716 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 14719 8590 14759 8630 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 14719 8504 14759 8544 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 14719 8418 14759 8458 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 14719 8332 14759 8372 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 14638 9192 14678 9232 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 14638 9106 14678 9146 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 14638 9020 14678 9060 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 14638 8934 14678 8974 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 14638 8848 14678 8888 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 14638 8762 14678 8802 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 14638 8676 14678 8716 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 14638 8590 14678 8630 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 14638 8504 14678 8544 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 14638 8418 14678 8458 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 14638 8332 14678 8372 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 14557 9192 14597 9232 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 14557 9106 14597 9146 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 14557 9020 14597 9060 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 14557 8934 14597 8974 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 14557 8848 14597 8888 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 14557 8762 14597 8802 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 14557 8676 14597 8716 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 14557 8590 14597 8630 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 14557 8504 14597 8544 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 14557 8418 14597 8458 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 14557 8332 14597 8372 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 14476 9192 14516 9232 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 14476 9106 14516 9146 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 14476 9020 14516 9060 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 14476 8934 14516 8974 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 14476 8848 14516 8888 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 14476 8762 14516 8802 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 14476 8676 14516 8716 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 14476 8590 14516 8630 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 14476 8504 14516 8544 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 14476 8418 14516 8458 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 14476 8332 14516 8372 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 14395 9192 14435 9232 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 14395 9106 14435 9146 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 14395 9020 14435 9060 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 14395 8934 14435 8974 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 14395 8848 14435 8888 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 14395 8762 14435 8802 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 14395 8676 14435 8716 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 14395 8590 14435 8630 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 14395 8504 14435 8544 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 14395 8418 14435 8458 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 14395 8332 14435 8372 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 14314 9192 14354 9232 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 14314 9106 14354 9146 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 14314 9020 14354 9060 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 14314 8934 14354 8974 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 14314 8848 14354 8888 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 14314 8762 14354 8802 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 14314 8676 14354 8716 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 14314 8590 14354 8630 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 14314 8504 14354 8544 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 14314 8418 14354 8458 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 14314 8332 14354 8372 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 14233 9192 14273 9232 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 14233 9106 14273 9146 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 14233 9020 14273 9060 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 14233 8934 14273 8974 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 14233 8848 14273 8888 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 14233 8762 14273 8802 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 14233 8676 14273 8716 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 14233 8590 14273 8630 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 14233 8504 14273 8544 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 14233 8418 14273 8458 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 14233 8332 14273 8372 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 14152 9192 14192 9232 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 14152 9106 14192 9146 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 14152 9020 14192 9060 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 14152 8934 14192 8974 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 14152 8848 14192 8888 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 14152 8762 14192 8802 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 14152 8676 14192 8716 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 14152 8590 14192 8630 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 14152 8504 14192 8544 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 14152 8418 14192 8458 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 14152 8332 14192 8372 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 14071 9192 14111 9232 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 14071 9106 14111 9146 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 14071 9020 14111 9060 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 14071 8934 14111 8974 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 14071 8848 14111 8888 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 14071 8762 14111 8802 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 14071 8676 14111 8716 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 14071 8590 14111 8630 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 14071 8504 14111 8544 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 14071 8418 14111 8458 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 14071 8332 14111 8372 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13990 9192 14030 9232 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13990 9106 14030 9146 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13990 9020 14030 9060 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13990 8934 14030 8974 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13990 8848 14030 8888 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13990 8762 14030 8802 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13990 8676 14030 8716 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13990 8590 14030 8630 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13990 8504 14030 8544 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13990 8418 14030 8458 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13990 8332 14030 8372 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13909 9192 13949 9232 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13909 9106 13949 9146 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13909 9020 13949 9060 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13909 8934 13949 8974 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13909 8848 13949 8888 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13909 8762 13949 8802 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13909 8676 13949 8716 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13909 8590 13949 8630 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13909 8504 13949 8544 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13909 8418 13949 8458 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13909 8332 13949 8372 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13828 9192 13868 9232 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13828 9106 13868 9146 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13828 9020 13868 9060 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13828 8934 13868 8974 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13828 8848 13868 8888 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13828 8762 13868 8802 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13828 8676 13868 8716 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13828 8590 13868 8630 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13828 8504 13868 8544 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13828 8418 13868 8458 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13828 8332 13868 8372 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13747 9192 13787 9232 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13747 9106 13787 9146 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13747 9020 13787 9060 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13747 8934 13787 8974 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13747 8848 13787 8888 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13747 8762 13787 8802 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13747 8676 13787 8716 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13747 8590 13787 8630 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13747 8504 13787 8544 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13747 8418 13787 8458 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13747 8332 13787 8372 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13666 9192 13706 9232 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13666 9106 13706 9146 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13666 9020 13706 9060 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13666 8934 13706 8974 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13666 8848 13706 8888 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13666 8762 13706 8802 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13666 8676 13706 8716 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13666 8590 13706 8630 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13666 8504 13706 8544 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13666 8418 13706 8458 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13666 8332 13706 8372 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13585 9192 13625 9232 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13585 9106 13625 9146 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13585 9020 13625 9060 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13585 8934 13625 8974 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13585 8848 13625 8888 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13585 8762 13625 8802 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13585 8676 13625 8716 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13585 8590 13625 8630 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13585 8504 13625 8544 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13585 8418 13625 8458 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13585 8332 13625 8372 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13504 9192 13544 9232 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13504 9106 13544 9146 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13504 9020 13544 9060 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13504 8934 13544 8974 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13504 8848 13544 8888 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13504 8762 13544 8802 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13504 8676 13544 8716 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13504 8590 13544 8630 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13504 8504 13544 8544 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13504 8418 13544 8458 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13504 8332 13544 8372 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13423 9192 13463 9232 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13423 9106 13463 9146 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13423 9020 13463 9060 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13423 8934 13463 8974 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13423 8848 13463 8888 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13423 8762 13463 8802 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13423 8676 13463 8716 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13423 8590 13463 8630 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13423 8504 13463 8544 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13423 8418 13463 8458 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13423 8332 13463 8372 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13342 9192 13382 9232 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13342 9106 13382 9146 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13342 9020 13382 9060 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13342 8934 13382 8974 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13342 8848 13382 8888 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13342 8762 13382 8802 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13342 8676 13382 8716 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13342 8590 13382 8630 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13342 8504 13382 8544 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13342 8418 13382 8458 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13342 8332 13382 8372 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13261 9192 13301 9232 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13261 9106 13301 9146 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13261 9020 13301 9060 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13261 8934 13301 8974 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13261 8848 13301 8888 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13261 8762 13301 8802 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13261 8676 13301 8716 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13261 8590 13301 8630 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13261 8504 13301 8544 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13261 8418 13301 8458 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13261 8332 13301 8372 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13180 9192 13220 9232 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13180 9106 13220 9146 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13180 9020 13220 9060 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13180 8934 13220 8974 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13180 8848 13220 8888 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13180 8762 13220 8802 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13180 8676 13220 8716 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13180 8590 13220 8630 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13180 8504 13220 8544 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13180 8418 13220 8458 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13180 8332 13220 8372 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13099 9192 13139 9232 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13099 9106 13139 9146 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13099 9020 13139 9060 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13099 8934 13139 8974 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13099 8848 13139 8888 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13099 8762 13139 8802 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13099 8676 13139 8716 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13099 8590 13139 8630 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13099 8504 13139 8544 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13099 8418 13139 8458 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13099 8332 13139 8372 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13018 9192 13058 9232 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13018 9106 13058 9146 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13018 9020 13058 9060 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13018 8934 13058 8974 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13018 8848 13058 8888 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13018 8762 13058 8802 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13018 8676 13058 8716 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13018 8590 13058 8630 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13018 8504 13058 8544 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13018 8418 13058 8458 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13018 8332 13058 8372 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 12937 9192 12977 9232 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 12937 9106 12977 9146 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 12937 9020 12977 9060 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 12937 8934 12977 8974 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 12937 8848 12977 8888 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 12937 8762 12977 8802 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 12937 8676 12977 8716 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 12937 8590 12977 8630 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 12937 8504 12977 8544 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 12937 8418 12977 8458 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 12937 8332 12977 8372 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 12856 9192 12896 9232 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 12856 9106 12896 9146 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 12856 9020 12896 9060 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 12856 8934 12896 8974 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 12856 8848 12896 8888 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 12856 8762 12896 8802 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 12856 8676 12896 8716 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 12856 8590 12896 8630 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 12856 8504 12896 8544 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 12856 8418 12896 8458 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 12856 8332 12896 8372 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 12775 9192 12815 9232 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 12775 9106 12815 9146 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 12775 9020 12815 9060 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 12775 8934 12815 8974 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 12775 8848 12815 8888 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 12775 8762 12815 8802 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 12775 8676 12815 8716 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 12775 8590 12815 8630 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 12775 8504 12815 8544 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 12775 8418 12815 8458 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 12775 8332 12815 8372 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 12694 9192 12734 9232 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 12694 9106 12734 9146 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 12694 9020 12734 9060 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 12694 8934 12734 8974 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 12694 8848 12734 8888 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 12694 8762 12734 8802 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 12694 8676 12734 8716 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 12694 8590 12734 8630 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 12694 8504 12734 8544 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 12694 8418 12734 8458 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 12694 8332 12734 8372 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 12613 9192 12653 9232 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 12613 9106 12653 9146 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 12613 9020 12653 9060 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 12613 8934 12653 8974 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 12613 8848 12653 8888 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 12613 8762 12653 8802 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 12613 8676 12653 8716 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 12613 8590 12653 8630 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 12613 8504 12653 8544 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 12613 8418 12653 8458 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 12613 8332 12653 8372 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 12532 9192 12572 9232 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 12532 9106 12572 9146 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 12532 9020 12572 9060 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 12532 8934 12572 8974 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 12532 8848 12572 8888 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 12532 8762 12572 8802 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 12532 8676 12572 8716 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 12532 8590 12572 8630 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 12532 8504 12572 8544 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 12532 8418 12572 8458 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 12532 8332 12572 8372 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 12451 9192 12491 9232 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 12451 9106 12491 9146 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 12451 9020 12491 9060 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 12451 8934 12491 8974 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 12451 8848 12491 8888 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 12451 8762 12491 8802 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 12451 8676 12491 8716 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 12451 8590 12491 8630 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 12451 8504 12491 8544 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 12451 8418 12491 8458 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 12451 8332 12491 8372 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 12370 9192 12410 9232 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 12370 9106 12410 9146 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 12370 9020 12410 9060 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 12370 8934 12410 8974 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 12370 8848 12410 8888 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 12370 8762 12410 8802 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 12370 8676 12410 8716 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 12370 8590 12410 8630 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 12370 8504 12410 8544 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 12370 8418 12410 8458 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 12370 8332 12410 8372 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 12289 9192 12329 9232 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 12289 9106 12329 9146 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 12289 9020 12329 9060 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 12289 8934 12329 8974 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 12289 8848 12329 8888 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 12289 8762 12329 8802 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 12289 8676 12329 8716 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 12289 8590 12329 8630 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 12289 8504 12329 8544 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 12289 8418 12329 8458 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 12289 8332 12329 8372 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 12208 9192 12248 9232 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 12208 9106 12248 9146 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 12208 9020 12248 9060 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 12208 8934 12248 8974 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 12208 8848 12248 8888 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 12208 8762 12248 8802 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 12208 8676 12248 8716 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 12208 8590 12248 8630 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 12208 8504 12248 8544 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 12208 8418 12248 8458 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 12208 8332 12248 8372 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 12127 9192 12167 9232 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 12127 9106 12167 9146 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 12127 9020 12167 9060 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 12127 8934 12167 8974 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 12127 8848 12167 8888 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 12127 8762 12167 8802 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 12127 8676 12167 8716 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 12127 8590 12167 8630 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 12127 8504 12167 8544 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 12127 8418 12167 8458 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 12127 8332 12167 8372 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 12046 9192 12086 9232 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 12046 9106 12086 9146 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 12046 9020 12086 9060 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 12046 8934 12086 8974 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 12046 8848 12086 8888 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 12046 8762 12086 8802 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 12046 8676 12086 8716 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 12046 8590 12086 8630 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 12046 8504 12086 8544 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 12046 8418 12086 8458 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 12046 8332 12086 8372 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 11965 9192 12005 9232 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 11965 9106 12005 9146 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 11965 9020 12005 9060 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 11965 8934 12005 8974 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 11965 8848 12005 8888 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 11965 8762 12005 8802 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 11965 8676 12005 8716 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 11965 8590 12005 8630 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 11965 8504 12005 8544 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 11965 8418 12005 8458 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 11965 8332 12005 8372 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 11884 9192 11924 9232 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 11884 9106 11924 9146 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 11884 9020 11924 9060 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 11884 8934 11924 8974 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 11884 8848 11924 8888 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 11884 8762 11924 8802 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 11884 8676 11924 8716 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 11884 8590 11924 8630 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 11884 8504 11924 8544 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 11884 8418 11924 8458 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 11884 8332 11924 8372 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 11803 9192 11843 9232 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 11803 9106 11843 9146 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 11803 9020 11843 9060 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 11803 8934 11843 8974 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 11803 8848 11843 8888 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 11803 8762 11843 8802 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 11803 8676 11843 8716 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 11803 8590 11843 8630 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 11803 8504 11843 8544 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 11803 8418 11843 8458 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 11803 8332 11843 8372 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 11722 9192 11762 9232 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 11722 9106 11762 9146 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 11722 9020 11762 9060 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 11722 8934 11762 8974 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 11722 8848 11762 8888 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 11722 8762 11762 8802 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 11722 8676 11762 8716 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 11722 8590 11762 8630 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 11722 8504 11762 8544 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 11722 8418 11762 8458 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 11722 8332 11762 8372 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 11641 9192 11681 9232 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 11641 9106 11681 9146 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 11641 9020 11681 9060 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 11641 8934 11681 8974 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 11641 8848 11681 8888 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 11641 8762 11681 8802 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 11641 8676 11681 8716 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 11641 8590 11681 8630 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 11641 8504 11681 8544 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 11641 8418 11681 8458 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 11641 8332 11681 8372 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 11560 9192 11600 9232 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 11560 9106 11600 9146 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 11560 9020 11600 9060 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 11560 8934 11600 8974 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 11560 8848 11600 8888 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 11560 8762 11600 8802 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 11560 8676 11600 8716 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 11560 8590 11600 8630 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 11560 8504 11600 8544 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 11560 8418 11600 8458 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 11560 8332 11600 8372 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 11479 9192 11519 9232 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 11479 9106 11519 9146 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 11479 9020 11519 9060 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 11479 8934 11519 8974 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 11479 8848 11519 8888 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 11479 8762 11519 8802 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 11479 8676 11519 8716 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 11479 8590 11519 8630 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 11479 8504 11519 8544 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 11479 8418 11519 8458 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 11479 8332 11519 8372 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 11398 9192 11438 9232 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 11398 9106 11438 9146 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 11398 9020 11438 9060 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 11398 8934 11438 8974 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 11398 8848 11438 8888 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 11398 8762 11438 8802 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 11398 8676 11438 8716 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 11398 8590 11438 8630 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 11398 8504 11438 8544 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 11398 8418 11438 8458 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 11398 8332 11438 8372 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 11317 9192 11357 9232 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 11317 9106 11357 9146 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 11317 9020 11357 9060 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 11317 8934 11357 8974 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 11317 8848 11357 8888 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 11317 8762 11357 8802 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 11317 8676 11357 8716 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 11317 8590 11357 8630 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 11317 8504 11357 8544 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 11317 8418 11357 8458 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 11317 8332 11357 8372 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 11236 9192 11276 9232 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 11236 9106 11276 9146 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 11236 9020 11276 9060 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 11236 8934 11276 8974 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 11236 8848 11276 8888 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 11236 8762 11276 8802 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 11236 8676 11276 8716 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 11236 8590 11276 8630 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 11236 8504 11276 8544 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 11236 8418 11276 8458 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 11236 8332 11276 8372 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 11155 9192 11195 9232 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 11155 9106 11195 9146 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 11155 9020 11195 9060 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 11155 8934 11195 8974 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 11155 8848 11195 8888 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 11155 8762 11195 8802 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 11155 8676 11195 8716 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 11155 8590 11195 8630 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 11155 8504 11195 8544 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 11155 8418 11195 8458 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 11155 8332 11195 8372 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 11074 9192 11114 9232 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 11074 9106 11114 9146 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 11074 9020 11114 9060 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 11074 8934 11114 8974 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 11074 8848 11114 8888 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 11074 8762 11114 8802 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 11074 8676 11114 8716 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 11074 8590 11114 8630 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 11074 8504 11114 8544 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 11074 8418 11114 8458 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 11074 8332 11114 8372 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 10993 9192 11033 9232 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 10993 9106 11033 9146 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 10993 9020 11033 9060 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 10993 8934 11033 8974 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 10993 8848 11033 8888 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 10993 8762 11033 8802 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 10993 8676 11033 8716 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 10993 8590 11033 8630 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 10993 8504 11033 8544 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 10993 8418 11033 8458 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 10993 8332 11033 8372 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 10912 9192 10952 9232 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 10912 9106 10952 9146 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 10912 9020 10952 9060 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 10912 8934 10952 8974 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 10912 8848 10952 8888 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 10912 8762 10952 8802 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 10912 8676 10952 8716 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 10912 8590 10952 8630 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 10912 8504 10952 8544 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 10912 8418 10952 8458 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 10912 8332 10952 8372 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 10831 9192 10871 9232 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 10831 9106 10871 9146 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 10831 9020 10871 9060 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 10831 8934 10871 8974 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 10831 8848 10871 8888 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 10831 8762 10871 8802 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 10831 8676 10871 8716 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 10831 8590 10871 8630 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 10831 8504 10871 8544 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 10831 8418 10871 8458 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 10831 8332 10871 8372 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 10750 9192 10790 9232 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 10750 9106 10790 9146 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 10750 9020 10790 9060 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 10750 8934 10790 8974 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 10750 8848 10790 8888 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 10750 8762 10790 8802 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 10750 8676 10790 8716 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 10750 8590 10790 8630 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 10750 8504 10790 8544 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 10750 8418 10790 8458 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 10750 8332 10790 8372 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 10669 9192 10709 9232 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 10669 9106 10709 9146 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 10669 9020 10709 9060 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 10669 8934 10709 8974 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 10669 8848 10709 8888 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 10669 8762 10709 8802 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 10669 8676 10709 8716 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 10669 8590 10709 8630 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 10669 8504 10709 8544 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 10669 8418 10709 8458 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 10669 8332 10709 8372 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 10588 9192 10628 9232 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 10588 9106 10628 9146 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 10588 9020 10628 9060 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 10588 8934 10628 8974 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 10588 8848 10628 8888 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 10588 8762 10628 8802 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 10588 8676 10628 8716 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 10588 8590 10628 8630 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 10588 8504 10628 8544 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 10588 8418 10628 8458 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 10588 8332 10628 8372 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 10506 9192 10546 9232 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 10506 9106 10546 9146 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 10506 9020 10546 9060 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 10506 8934 10546 8974 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 10506 8848 10546 8888 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 10506 8762 10546 8802 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 10506 8676 10546 8716 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 10506 8590 10546 8630 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 10506 8504 10546 8544 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 10506 8418 10546 8458 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 10506 8332 10546 8372 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 10424 9192 10464 9232 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 10424 9106 10464 9146 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 10424 9020 10464 9060 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 10424 8934 10464 8974 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 10424 8848 10464 8888 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 10424 8762 10464 8802 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 10424 8676 10464 8716 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 10424 8590 10464 8630 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 10424 8504 10464 8544 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 10424 8418 10464 8458 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 10424 8332 10464 8372 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 10342 9192 10382 9232 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 10342 9106 10382 9146 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 10342 9020 10382 9060 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 10342 8934 10382 8974 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 10342 8848 10382 8888 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 10342 8762 10382 8802 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 10342 8676 10382 8716 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 10342 8590 10382 8630 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 10342 8504 10382 8544 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 10342 8418 10382 8458 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 10342 8332 10382 8372 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 10260 9192 10300 9232 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 10260 9106 10300 9146 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 10260 9020 10300 9060 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 10260 8934 10300 8974 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 10260 8848 10300 8888 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 10260 8762 10300 8802 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 10260 8676 10300 8716 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 10260 8590 10300 8630 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 10260 8504 10300 8544 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 10260 8418 10300 8458 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 10260 8332 10300 8372 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 10178 9192 10218 9232 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 10178 9106 10218 9146 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 10178 9020 10218 9060 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 10178 8934 10218 8974 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 10178 8848 10218 8888 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 10178 8762 10218 8802 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 10178 8676 10218 8716 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 10178 8590 10218 8630 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 10178 8504 10218 8544 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 10178 8418 10218 8458 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 10178 8332 10218 8372 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 10096 9192 10136 9232 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 10096 9106 10136 9146 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 10096 9020 10136 9060 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 10096 8934 10136 8974 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 10096 8848 10136 8888 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 10096 8762 10136 8802 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 10096 8676 10136 8716 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 10096 8590 10136 8630 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 10096 8504 10136 8544 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 10096 8418 10136 8458 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 10096 8332 10136 8372 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 4821 9192 4861 9232 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 4821 9106 4861 9146 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 4821 9020 4861 9060 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 4821 8934 4861 8974 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 4821 8848 4861 8888 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 4821 8762 4861 8802 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 4821 8676 4861 8716 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 4821 8590 4861 8630 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 4821 8504 4861 8544 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 4821 8418 4861 8458 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 4821 8332 4861 8372 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 4741 9192 4781 9232 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 4741 9106 4781 9146 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 4741 9020 4781 9060 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 4741 8934 4781 8974 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 4741 8848 4781 8888 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 4741 8762 4781 8802 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 4741 8676 4781 8716 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 4741 8590 4781 8630 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 4741 8504 4781 8544 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 4741 8418 4781 8458 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 4741 8332 4781 8372 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 4661 9192 4701 9232 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 4661 9106 4701 9146 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 4661 9020 4701 9060 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 4661 8934 4701 8974 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 4661 8848 4701 8888 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 4661 8762 4701 8802 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 4661 8676 4701 8716 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 4661 8590 4701 8630 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 4661 8504 4701 8544 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 4661 8418 4701 8458 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 4661 8332 4701 8372 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 4581 9192 4621 9232 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 4581 9106 4621 9146 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 4581 9020 4621 9060 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 4581 8934 4621 8974 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 4581 8848 4621 8888 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 4581 8762 4621 8802 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 4581 8676 4621 8716 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 4581 8590 4621 8630 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 4581 8504 4621 8544 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 4581 8418 4621 8458 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 4581 8332 4621 8372 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 4501 9192 4541 9232 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 4501 9106 4541 9146 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 4501 9020 4541 9060 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 4501 8934 4541 8974 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 4501 8848 4541 8888 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 4501 8762 4541 8802 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 4501 8676 4541 8716 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 4501 8590 4541 8630 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 4501 8504 4541 8544 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 4501 8418 4541 8458 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 4501 8332 4541 8372 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 4421 9192 4461 9232 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 4421 9106 4461 9146 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 4421 9020 4461 9060 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 4421 8934 4461 8974 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 4421 8848 4461 8888 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 4421 8762 4461 8802 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 4421 8676 4461 8716 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 4421 8590 4461 8630 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 4421 8504 4461 8544 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 4421 8418 4461 8458 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 4421 8332 4461 8372 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 4341 9192 4381 9232 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 4341 9106 4381 9146 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 4341 9020 4381 9060 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 4341 8934 4381 8974 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 4341 8848 4381 8888 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 4341 8762 4381 8802 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 4341 8676 4381 8716 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 4341 8590 4381 8630 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 4341 8504 4381 8544 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 4341 8418 4381 8458 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 4341 8332 4381 8372 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 4261 9192 4301 9232 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 4261 9106 4301 9146 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 4261 9020 4301 9060 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 4261 8934 4301 8974 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 4261 8848 4301 8888 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 4261 8762 4301 8802 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 4261 8676 4301 8716 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 4261 8590 4301 8630 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 4261 8504 4301 8544 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 4261 8418 4301 8458 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 4261 8332 4301 8372 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 4181 9192 4221 9232 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 4181 9106 4221 9146 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 4181 9020 4221 9060 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 4181 8934 4221 8974 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 4181 8848 4221 8888 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 4181 8762 4221 8802 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 4181 8676 4221 8716 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 4181 8590 4221 8630 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 4181 8504 4221 8544 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 4181 8418 4221 8458 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 4181 8332 4221 8372 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 4100 9192 4140 9232 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 4100 9106 4140 9146 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 4100 9020 4140 9060 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 4100 8934 4140 8974 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 4100 8848 4140 8888 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 4100 8762 4140 8802 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 4100 8676 4140 8716 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 4100 8590 4140 8630 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 4100 8504 4140 8544 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 4100 8418 4140 8458 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 4100 8332 4140 8372 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 4019 9192 4059 9232 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 4019 9106 4059 9146 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 4019 9020 4059 9060 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 4019 8934 4059 8974 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 4019 8848 4059 8888 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 4019 8762 4059 8802 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 4019 8676 4059 8716 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 4019 8590 4059 8630 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 4019 8504 4059 8544 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 4019 8418 4059 8458 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 4019 8332 4059 8372 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3938 9192 3978 9232 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3938 9106 3978 9146 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3938 9020 3978 9060 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3938 8934 3978 8974 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3938 8848 3978 8888 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3938 8762 3978 8802 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3938 8676 3978 8716 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3938 8590 3978 8630 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3938 8504 3978 8544 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3938 8418 3978 8458 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3938 8332 3978 8372 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3857 9192 3897 9232 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3857 9106 3897 9146 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3857 9020 3897 9060 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3857 8934 3897 8974 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3857 8848 3897 8888 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3857 8762 3897 8802 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3857 8676 3897 8716 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3857 8590 3897 8630 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3857 8504 3897 8544 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3857 8418 3897 8458 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3857 8332 3897 8372 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3776 9192 3816 9232 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3776 9106 3816 9146 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3776 9020 3816 9060 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3776 8934 3816 8974 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3776 8848 3816 8888 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3776 8762 3816 8802 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3776 8676 3816 8716 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3776 8590 3816 8630 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3776 8504 3816 8544 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3776 8418 3816 8458 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3776 8332 3816 8372 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3695 9192 3735 9232 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3695 9106 3735 9146 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3695 9020 3735 9060 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3695 8934 3735 8974 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3695 8848 3735 8888 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3695 8762 3735 8802 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3695 8676 3735 8716 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3695 8590 3735 8630 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3695 8504 3735 8544 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3695 8418 3735 8458 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3695 8332 3735 8372 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3614 9192 3654 9232 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3614 9106 3654 9146 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3614 9020 3654 9060 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3614 8934 3654 8974 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3614 8848 3654 8888 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3614 8762 3654 8802 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3614 8676 3654 8716 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3614 8590 3654 8630 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3614 8504 3654 8544 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3614 8418 3654 8458 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3614 8332 3654 8372 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3533 9192 3573 9232 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3533 9106 3573 9146 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3533 9020 3573 9060 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3533 8934 3573 8974 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3533 8848 3573 8888 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3533 8762 3573 8802 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3533 8676 3573 8716 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3533 8590 3573 8630 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3533 8504 3573 8544 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3533 8418 3573 8458 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3533 8332 3573 8372 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3452 9192 3492 9232 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3452 9106 3492 9146 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3452 9020 3492 9060 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3452 8934 3492 8974 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3452 8848 3492 8888 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3452 8762 3492 8802 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3452 8676 3492 8716 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3452 8590 3492 8630 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3452 8504 3492 8544 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3452 8418 3492 8458 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3452 8332 3492 8372 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3371 9192 3411 9232 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3371 9106 3411 9146 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3371 9020 3411 9060 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3371 8934 3411 8974 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3371 8848 3411 8888 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3371 8762 3411 8802 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3371 8676 3411 8716 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3371 8590 3411 8630 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3371 8504 3411 8544 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3371 8418 3411 8458 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3371 8332 3411 8372 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3290 9192 3330 9232 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3290 9106 3330 9146 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3290 9020 3330 9060 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3290 8934 3330 8974 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3290 8848 3330 8888 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3290 8762 3330 8802 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3290 8676 3330 8716 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3290 8590 3330 8630 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3290 8504 3330 8544 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3290 8418 3330 8458 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3290 8332 3330 8372 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3209 9192 3249 9232 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3209 9106 3249 9146 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3209 9020 3249 9060 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3209 8934 3249 8974 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3209 8848 3249 8888 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3209 8762 3249 8802 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3209 8676 3249 8716 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3209 8590 3249 8630 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3209 8504 3249 8544 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3209 8418 3249 8458 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3209 8332 3249 8372 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3128 9192 3168 9232 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3128 9106 3168 9146 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3128 9020 3168 9060 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3128 8934 3168 8974 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3128 8848 3168 8888 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3128 8762 3168 8802 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3128 8676 3168 8716 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3128 8590 3168 8630 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3128 8504 3168 8544 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3128 8418 3168 8458 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3128 8332 3168 8372 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3047 9192 3087 9232 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3047 9106 3087 9146 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3047 9020 3087 9060 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3047 8934 3087 8974 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3047 8848 3087 8888 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3047 8762 3087 8802 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3047 8676 3087 8716 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3047 8590 3087 8630 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3047 8504 3087 8544 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3047 8418 3087 8458 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3047 8332 3087 8372 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 2966 9192 3006 9232 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 2966 9106 3006 9146 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 2966 9020 3006 9060 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 2966 8934 3006 8974 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 2966 8848 3006 8888 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 2966 8762 3006 8802 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 2966 8676 3006 8716 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 2966 8590 3006 8630 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 2966 8504 3006 8544 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 2966 8418 3006 8458 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 2966 8332 3006 8372 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 2885 9192 2925 9232 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 2885 9106 2925 9146 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 2885 9020 2925 9060 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 2885 8934 2925 8974 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 2885 8848 2925 8888 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 2885 8762 2925 8802 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 2885 8676 2925 8716 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 2885 8590 2925 8630 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 2885 8504 2925 8544 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 2885 8418 2925 8458 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 2885 8332 2925 8372 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 2804 9192 2844 9232 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 2804 9106 2844 9146 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 2804 9020 2844 9060 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 2804 8934 2844 8974 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 2804 8848 2844 8888 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 2804 8762 2844 8802 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 2804 8676 2844 8716 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 2804 8590 2844 8630 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 2804 8504 2844 8544 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 2804 8418 2844 8458 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 2804 8332 2844 8372 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 2723 9192 2763 9232 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 2723 9106 2763 9146 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 2723 9020 2763 9060 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 2723 8934 2763 8974 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 2723 8848 2763 8888 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 2723 8762 2763 8802 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 2723 8676 2763 8716 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 2723 8590 2763 8630 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 2723 8504 2763 8544 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 2723 8418 2763 8458 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 2723 8332 2763 8372 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 2642 9192 2682 9232 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 2642 9106 2682 9146 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 2642 9020 2682 9060 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 2642 8934 2682 8974 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 2642 8848 2682 8888 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 2642 8762 2682 8802 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 2642 8676 2682 8716 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 2642 8590 2682 8630 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 2642 8504 2682 8544 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 2642 8418 2682 8458 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 2642 8332 2682 8372 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 2561 9192 2601 9232 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 2561 9106 2601 9146 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 2561 9020 2601 9060 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 2561 8934 2601 8974 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 2561 8848 2601 8888 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 2561 8762 2601 8802 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 2561 8676 2601 8716 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 2561 8590 2601 8630 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 2561 8504 2601 8544 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 2561 8418 2601 8458 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 2561 8332 2601 8372 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 2480 9192 2520 9232 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 2480 9106 2520 9146 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 2480 9020 2520 9060 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 2480 8934 2520 8974 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 2480 8848 2520 8888 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 2480 8762 2520 8802 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 2480 8676 2520 8716 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 2480 8590 2520 8630 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 2480 8504 2520 8544 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 2480 8418 2520 8458 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 2480 8332 2520 8372 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 2399 9192 2439 9232 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 2399 9106 2439 9146 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 2399 9020 2439 9060 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 2399 8934 2439 8974 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 2399 8848 2439 8888 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 2399 8762 2439 8802 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 2399 8676 2439 8716 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 2399 8590 2439 8630 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 2399 8504 2439 8544 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 2399 8418 2439 8458 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 2399 8332 2439 8372 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 2318 9192 2358 9232 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 2318 9106 2358 9146 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 2318 9020 2358 9060 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 2318 8934 2358 8974 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 2318 8848 2358 8888 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 2318 8762 2358 8802 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 2318 8676 2358 8716 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 2318 8590 2358 8630 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 2318 8504 2358 8544 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 2318 8418 2358 8458 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 2318 8332 2358 8372 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 2237 9192 2277 9232 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 2237 9106 2277 9146 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 2237 9020 2277 9060 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 2237 8934 2277 8974 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 2237 8848 2277 8888 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 2237 8762 2277 8802 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 2237 8676 2277 8716 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 2237 8590 2277 8630 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 2237 8504 2277 8544 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 2237 8418 2277 8458 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 2237 8332 2277 8372 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 2156 9192 2196 9232 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 2156 9106 2196 9146 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 2156 9020 2196 9060 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 2156 8934 2196 8974 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 2156 8848 2196 8888 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 2156 8762 2196 8802 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 2156 8676 2196 8716 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 2156 8590 2196 8630 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 2156 8504 2196 8544 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 2156 8418 2196 8458 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 2156 8332 2196 8372 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 2075 9192 2115 9232 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 2075 9106 2115 9146 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 2075 9020 2115 9060 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 2075 8934 2115 8974 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 2075 8848 2115 8888 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 2075 8762 2115 8802 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 2075 8676 2115 8716 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 2075 8590 2115 8630 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 2075 8504 2115 8544 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 2075 8418 2115 8458 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 2075 8332 2115 8372 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1994 9192 2034 9232 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1994 9106 2034 9146 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1994 9020 2034 9060 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1994 8934 2034 8974 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1994 8848 2034 8888 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1994 8762 2034 8802 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1994 8676 2034 8716 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1994 8590 2034 8630 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1994 8504 2034 8544 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1994 8418 2034 8458 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1994 8332 2034 8372 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1913 9192 1953 9232 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1913 9106 1953 9146 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1913 9020 1953 9060 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1913 8934 1953 8974 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1913 8848 1953 8888 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1913 8762 1953 8802 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1913 8676 1953 8716 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1913 8590 1953 8630 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1913 8504 1953 8544 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1913 8418 1953 8458 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1913 8332 1953 8372 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1832 9192 1872 9232 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1832 9106 1872 9146 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1832 9020 1872 9060 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1832 8934 1872 8974 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1832 8848 1872 8888 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1832 8762 1872 8802 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1832 8676 1872 8716 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1832 8590 1872 8630 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1832 8504 1872 8544 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1832 8418 1872 8458 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1832 8332 1872 8372 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1751 9192 1791 9232 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1751 9106 1791 9146 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1751 9020 1791 9060 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1751 8934 1791 8974 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1751 8848 1791 8888 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1751 8762 1791 8802 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1751 8676 1791 8716 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1751 8590 1791 8630 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1751 8504 1791 8544 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1751 8418 1791 8458 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1751 8332 1791 8372 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1670 9192 1710 9232 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1670 9106 1710 9146 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1670 9020 1710 9060 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1670 8934 1710 8974 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1670 8848 1710 8888 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1670 8762 1710 8802 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1670 8676 1710 8716 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1670 8590 1710 8630 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1670 8504 1710 8544 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1670 8418 1710 8458 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1670 8332 1710 8372 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1589 9192 1629 9232 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1589 9106 1629 9146 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1589 9020 1629 9060 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1589 8934 1629 8974 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1589 8848 1629 8888 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1589 8762 1629 8802 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1589 8676 1629 8716 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1589 8590 1629 8630 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1589 8504 1629 8544 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1589 8418 1629 8458 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1589 8332 1629 8372 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1508 9192 1548 9232 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1508 9106 1548 9146 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1508 9020 1548 9060 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1508 8934 1548 8974 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1508 8848 1548 8888 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1508 8762 1548 8802 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1508 8676 1548 8716 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1508 8590 1548 8630 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1508 8504 1548 8544 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1508 8418 1548 8458 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1508 8332 1548 8372 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1427 9192 1467 9232 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1427 9106 1467 9146 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1427 9020 1467 9060 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1427 8934 1467 8974 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1427 8848 1467 8888 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1427 8762 1467 8802 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1427 8676 1467 8716 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1427 8590 1467 8630 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1427 8504 1467 8544 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1427 8418 1467 8458 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1427 8332 1467 8372 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1346 9192 1386 9232 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1346 9106 1386 9146 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1346 9020 1386 9060 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1346 8934 1386 8974 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1346 8848 1386 8888 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1346 8762 1386 8802 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1346 8676 1386 8716 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1346 8590 1386 8630 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1346 8504 1386 8544 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1346 8418 1386 8458 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1346 8332 1386 8372 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1265 9192 1305 9232 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1265 9106 1305 9146 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1265 9020 1305 9060 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1265 8934 1305 8974 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1265 8848 1305 8888 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1265 8762 1305 8802 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1265 8676 1305 8716 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1265 8590 1305 8630 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1265 8504 1305 8544 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1265 8418 1305 8458 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1265 8332 1305 8372 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1184 9192 1224 9232 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1184 9106 1224 9146 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1184 9020 1224 9060 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1184 8934 1224 8974 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1184 8848 1224 8888 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1184 8762 1224 8802 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1184 8676 1224 8716 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1184 8590 1224 8630 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1184 8504 1224 8544 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1184 8418 1224 8458 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1184 8332 1224 8372 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1103 9192 1143 9232 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1103 9106 1143 9146 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1103 9020 1143 9060 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1103 8934 1143 8974 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1103 8848 1143 8888 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1103 8762 1143 8802 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1103 8676 1143 8716 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1103 8590 1143 8630 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1103 8504 1143 8544 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1103 8418 1143 8458 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1103 8332 1143 8372 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1022 9192 1062 9232 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1022 9106 1062 9146 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1022 9020 1062 9060 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1022 8934 1062 8974 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1022 8848 1062 8888 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1022 8762 1062 8802 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1022 8676 1062 8716 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1022 8590 1062 8630 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1022 8504 1062 8544 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1022 8418 1062 8458 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1022 8332 1062 8372 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 941 9192 981 9232 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 941 9106 981 9146 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 941 9020 981 9060 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 941 8934 981 8974 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 941 8848 981 8888 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 941 8762 981 8802 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 941 8676 981 8716 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 941 8590 981 8630 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 941 8504 981 8544 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 941 8418 981 8458 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 941 8332 981 8372 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 860 9192 900 9232 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 860 9106 900 9146 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 860 9020 900 9060 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 860 8934 900 8974 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 860 8848 900 8888 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 860 8762 900 8802 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 860 8676 900 8716 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 860 8590 900 8630 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 860 8504 900 8544 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 860 8418 900 8458 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 860 8332 900 8372 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 779 9192 819 9232 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 779 9106 819 9146 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 779 9020 819 9060 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 779 8934 819 8974 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 779 8848 819 8888 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 779 8762 819 8802 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 779 8676 819 8716 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 779 8590 819 8630 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 779 8504 819 8544 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 779 8418 819 8458 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 779 8332 819 8372 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 698 9192 738 9232 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 698 9106 738 9146 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 698 9020 738 9060 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 698 8934 738 8974 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 698 8848 738 8888 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 698 8762 738 8802 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 698 8676 738 8716 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 698 8590 738 8630 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 698 8504 738 8544 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 698 8418 738 8458 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 698 8332 738 8372 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 617 9192 657 9232 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 617 9106 657 9146 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 617 9020 657 9060 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 617 8934 657 8974 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 617 8848 657 8888 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 617 8762 657 8802 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 617 8676 657 8716 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 617 8590 657 8630 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 617 8504 657 8544 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 617 8418 657 8458 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 617 8332 657 8372 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 536 9192 576 9232 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 536 9106 576 9146 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 536 9020 576 9060 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 536 8934 576 8974 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 536 8848 576 8888 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 536 8762 576 8802 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 536 8676 576 8716 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 536 8590 576 8630 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 536 8504 576 8544 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 536 8418 576 8458 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 536 8332 576 8372 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 455 9192 495 9232 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 455 9106 495 9146 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 455 9020 495 9060 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 455 8934 495 8974 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 455 8848 495 8888 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 455 8762 495 8802 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 455 8676 495 8716 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 455 8590 495 8630 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 455 8504 495 8544 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 455 8418 495 8458 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 455 8332 495 8372 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 374 9192 414 9232 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 374 9106 414 9146 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 374 9020 414 9060 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 374 8934 414 8974 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 374 8848 414 8888 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 374 8762 414 8802 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 374 8676 414 8716 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 374 8590 414 8630 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 374 8504 414 8544 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 374 8418 414 8458 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 374 8332 414 8372 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 293 9192 333 9232 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 293 9106 333 9146 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 293 9020 333 9060 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 293 8934 333 8974 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 293 8848 333 8888 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 293 8762 333 8802 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 293 8676 333 8716 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 293 8590 333 8630 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 293 8504 333 8544 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 293 8418 333 8458 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 293 8332 333 8372 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 212 9192 252 9232 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 212 9106 252 9146 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 212 9020 252 9060 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 212 8934 252 8974 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 212 8848 252 8888 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 212 8762 252 8802 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 212 8676 252 8716 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 212 8590 252 8630 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 212 8504 252 8544 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 212 8418 252 8458 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 212 8332 252 8372 1 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 0 5167 254 6097 1 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 14746 35157 15000 40000 1 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 14746 5167 15000 6097 1 VSSIO
port 5 nsew ground bidirectional
rlabel metal5 s 0 35157 254 40000 1 VSSIO
port 5 nsew ground bidirectional
rlabel metal5 s 0 5187 254 6077 1 VSSIO
port 5 nsew ground bidirectional
rlabel metal5 s 14746 35157 15000 40000 1 VSSIO
port 5 nsew ground bidirectional
rlabel metal5 s 14746 5187 15000 6077 1 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 14746 11647 15000 12537 1 VSSIO_Q
port 6 nsew ground bidirectional
rlabel metal5 s 0 11667 254 12517 1 VSSIO_Q
port 6 nsew ground bidirectional
rlabel metal5 s 14746 11667 15000 12517 1 VSSIO_Q
port 6 nsew ground bidirectional
rlabel metal4 s 14746 6377 15000 7067 1 VSWITCH
port 7 nsew power bidirectional
rlabel metal5 s 0 6397 254 7047 1 VSWITCH
port 7 nsew power bidirectional
rlabel metal5 s 14746 6397 15000 7047 1 VSWITCH
port 7 nsew power bidirectional
<< properties >>
string FIXED_BBOX 0 0 15000 40000
string GDS_END 2174082
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 2083250
string LEFclass PAD
string LEFsymmetry X Y R90
<< end >>
