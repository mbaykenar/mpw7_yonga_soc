magic
tech sky130B
magscale 1 2
timestamp 1649977179
<< metal3 >>
rect 10078 8318 14858 9246
<< obsm3 >>
rect 194 8318 4879 9246
<< metal4 >>
rect 0 35157 254 40000
rect 14746 35157 15000 40000
rect 0 14007 254 19000
rect 14746 14007 15000 19000
rect 0 12817 254 13707
rect 14746 12817 15000 13707
rect 0 11647 254 12537
rect 14746 11647 15000 12537
rect 0 11281 15000 11347
rect 0 10625 15000 11221
rect 0 10329 254 10565
rect 14746 10329 15000 10565
rect 0 9673 15000 10269
rect 0 9547 15000 9613
rect 0 9244 254 9247
rect 0 9180 264 9244
rect 281 9180 345 9244
rect 362 9180 426 9244
rect 443 9180 507 9244
rect 524 9180 588 9244
rect 605 9180 669 9244
rect 686 9180 750 9244
rect 767 9180 831 9244
rect 848 9180 912 9244
rect 929 9180 993 9244
rect 1010 9180 1074 9244
rect 1091 9180 1155 9244
rect 1172 9180 1236 9244
rect 1253 9180 1317 9244
rect 1334 9180 1398 9244
rect 1415 9180 1479 9244
rect 1496 9180 1560 9244
rect 1577 9180 1641 9244
rect 1658 9180 1722 9244
rect 1739 9180 1803 9244
rect 1820 9180 1884 9244
rect 1901 9180 1965 9244
rect 1982 9180 2046 9244
rect 2063 9180 2127 9244
rect 2144 9180 2208 9244
rect 2225 9180 2289 9244
rect 2306 9180 2370 9244
rect 2387 9180 2451 9244
rect 2468 9180 2532 9244
rect 2549 9180 2613 9244
rect 2630 9180 2694 9244
rect 2711 9180 2775 9244
rect 2792 9180 2856 9244
rect 2873 9180 2937 9244
rect 2954 9180 3018 9244
rect 3035 9180 3099 9244
rect 3116 9180 3180 9244
rect 3197 9180 3261 9244
rect 3278 9180 3342 9244
rect 3359 9180 3423 9244
rect 3440 9180 3504 9244
rect 3521 9180 3585 9244
rect 3602 9180 3666 9244
rect 3683 9180 3747 9244
rect 3764 9180 3828 9244
rect 3845 9180 3909 9244
rect 3926 9180 3990 9244
rect 4007 9180 4071 9244
rect 4088 9180 4152 9244
rect 4169 9180 4233 9244
rect 4249 9180 4313 9244
rect 4329 9180 4393 9244
rect 4409 9180 4473 9244
rect 4489 9180 4553 9244
rect 4569 9180 4633 9244
rect 4649 9180 4713 9244
rect 4729 9180 4793 9244
rect 4809 9180 4873 9244
rect 0 9158 254 9180
rect 0 9094 264 9158
rect 281 9094 345 9158
rect 362 9094 426 9158
rect 443 9094 507 9158
rect 524 9094 588 9158
rect 605 9094 669 9158
rect 686 9094 750 9158
rect 767 9094 831 9158
rect 848 9094 912 9158
rect 929 9094 993 9158
rect 1010 9094 1074 9158
rect 1091 9094 1155 9158
rect 1172 9094 1236 9158
rect 1253 9094 1317 9158
rect 1334 9094 1398 9158
rect 1415 9094 1479 9158
rect 1496 9094 1560 9158
rect 1577 9094 1641 9158
rect 1658 9094 1722 9158
rect 1739 9094 1803 9158
rect 1820 9094 1884 9158
rect 1901 9094 1965 9158
rect 1982 9094 2046 9158
rect 2063 9094 2127 9158
rect 2144 9094 2208 9158
rect 2225 9094 2289 9158
rect 2306 9094 2370 9158
rect 2387 9094 2451 9158
rect 2468 9094 2532 9158
rect 2549 9094 2613 9158
rect 2630 9094 2694 9158
rect 2711 9094 2775 9158
rect 2792 9094 2856 9158
rect 2873 9094 2937 9158
rect 2954 9094 3018 9158
rect 3035 9094 3099 9158
rect 3116 9094 3180 9158
rect 3197 9094 3261 9158
rect 3278 9094 3342 9158
rect 3359 9094 3423 9158
rect 3440 9094 3504 9158
rect 3521 9094 3585 9158
rect 3602 9094 3666 9158
rect 3683 9094 3747 9158
rect 3764 9094 3828 9158
rect 3845 9094 3909 9158
rect 3926 9094 3990 9158
rect 4007 9094 4071 9158
rect 4088 9094 4152 9158
rect 4169 9094 4233 9158
rect 4249 9094 4313 9158
rect 4329 9094 4393 9158
rect 4409 9094 4473 9158
rect 4489 9094 4553 9158
rect 4569 9094 4633 9158
rect 4649 9094 4713 9158
rect 4729 9094 4793 9158
rect 4809 9094 4873 9158
rect 0 9072 254 9094
rect 0 9008 264 9072
rect 281 9008 345 9072
rect 362 9008 426 9072
rect 443 9008 507 9072
rect 524 9008 588 9072
rect 605 9008 669 9072
rect 686 9008 750 9072
rect 767 9008 831 9072
rect 848 9008 912 9072
rect 929 9008 993 9072
rect 1010 9008 1074 9072
rect 1091 9008 1155 9072
rect 1172 9008 1236 9072
rect 1253 9008 1317 9072
rect 1334 9008 1398 9072
rect 1415 9008 1479 9072
rect 1496 9008 1560 9072
rect 1577 9008 1641 9072
rect 1658 9008 1722 9072
rect 1739 9008 1803 9072
rect 1820 9008 1884 9072
rect 1901 9008 1965 9072
rect 1982 9008 2046 9072
rect 2063 9008 2127 9072
rect 2144 9008 2208 9072
rect 2225 9008 2289 9072
rect 2306 9008 2370 9072
rect 2387 9008 2451 9072
rect 2468 9008 2532 9072
rect 2549 9008 2613 9072
rect 2630 9008 2694 9072
rect 2711 9008 2775 9072
rect 2792 9008 2856 9072
rect 2873 9008 2937 9072
rect 2954 9008 3018 9072
rect 3035 9008 3099 9072
rect 3116 9008 3180 9072
rect 3197 9008 3261 9072
rect 3278 9008 3342 9072
rect 3359 9008 3423 9072
rect 3440 9008 3504 9072
rect 3521 9008 3585 9072
rect 3602 9008 3666 9072
rect 3683 9008 3747 9072
rect 3764 9008 3828 9072
rect 3845 9008 3909 9072
rect 3926 9008 3990 9072
rect 4007 9008 4071 9072
rect 4088 9008 4152 9072
rect 4169 9008 4233 9072
rect 4249 9008 4313 9072
rect 4329 9008 4393 9072
rect 4409 9008 4473 9072
rect 4489 9008 4553 9072
rect 4569 9008 4633 9072
rect 4649 9008 4713 9072
rect 4729 9008 4793 9072
rect 4809 9008 4873 9072
rect 0 8986 254 9008
rect 0 8922 264 8986
rect 281 8922 345 8986
rect 362 8922 426 8986
rect 443 8922 507 8986
rect 524 8922 588 8986
rect 605 8922 669 8986
rect 686 8922 750 8986
rect 767 8922 831 8986
rect 848 8922 912 8986
rect 929 8922 993 8986
rect 1010 8922 1074 8986
rect 1091 8922 1155 8986
rect 1172 8922 1236 8986
rect 1253 8922 1317 8986
rect 1334 8922 1398 8986
rect 1415 8922 1479 8986
rect 1496 8922 1560 8986
rect 1577 8922 1641 8986
rect 1658 8922 1722 8986
rect 1739 8922 1803 8986
rect 1820 8922 1884 8986
rect 1901 8922 1965 8986
rect 1982 8922 2046 8986
rect 2063 8922 2127 8986
rect 2144 8922 2208 8986
rect 2225 8922 2289 8986
rect 2306 8922 2370 8986
rect 2387 8922 2451 8986
rect 2468 8922 2532 8986
rect 2549 8922 2613 8986
rect 2630 8922 2694 8986
rect 2711 8922 2775 8986
rect 2792 8922 2856 8986
rect 2873 8922 2937 8986
rect 2954 8922 3018 8986
rect 3035 8922 3099 8986
rect 3116 8922 3180 8986
rect 3197 8922 3261 8986
rect 3278 8922 3342 8986
rect 3359 8922 3423 8986
rect 3440 8922 3504 8986
rect 3521 8922 3585 8986
rect 3602 8922 3666 8986
rect 3683 8922 3747 8986
rect 3764 8922 3828 8986
rect 3845 8922 3909 8986
rect 3926 8922 3990 8986
rect 4007 8922 4071 8986
rect 4088 8922 4152 8986
rect 4169 8922 4233 8986
rect 4249 8922 4313 8986
rect 4329 8922 4393 8986
rect 4409 8922 4473 8986
rect 4489 8922 4553 8986
rect 4569 8922 4633 8986
rect 4649 8922 4713 8986
rect 4729 8922 4793 8986
rect 4809 8922 4873 8986
rect 0 8900 254 8922
rect 0 8836 264 8900
rect 281 8836 345 8900
rect 362 8836 426 8900
rect 443 8836 507 8900
rect 524 8836 588 8900
rect 605 8836 669 8900
rect 686 8836 750 8900
rect 767 8836 831 8900
rect 848 8836 912 8900
rect 929 8836 993 8900
rect 1010 8836 1074 8900
rect 1091 8836 1155 8900
rect 1172 8836 1236 8900
rect 1253 8836 1317 8900
rect 1334 8836 1398 8900
rect 1415 8836 1479 8900
rect 1496 8836 1560 8900
rect 1577 8836 1641 8900
rect 1658 8836 1722 8900
rect 1739 8836 1803 8900
rect 1820 8836 1884 8900
rect 1901 8836 1965 8900
rect 1982 8836 2046 8900
rect 2063 8836 2127 8900
rect 2144 8836 2208 8900
rect 2225 8836 2289 8900
rect 2306 8836 2370 8900
rect 2387 8836 2451 8900
rect 2468 8836 2532 8900
rect 2549 8836 2613 8900
rect 2630 8836 2694 8900
rect 2711 8836 2775 8900
rect 2792 8836 2856 8900
rect 2873 8836 2937 8900
rect 2954 8836 3018 8900
rect 3035 8836 3099 8900
rect 3116 8836 3180 8900
rect 3197 8836 3261 8900
rect 3278 8836 3342 8900
rect 3359 8836 3423 8900
rect 3440 8836 3504 8900
rect 3521 8836 3585 8900
rect 3602 8836 3666 8900
rect 3683 8836 3747 8900
rect 3764 8836 3828 8900
rect 3845 8836 3909 8900
rect 3926 8836 3990 8900
rect 4007 8836 4071 8900
rect 4088 8836 4152 8900
rect 4169 8836 4233 8900
rect 4249 8836 4313 8900
rect 4329 8836 4393 8900
rect 4409 8836 4473 8900
rect 4489 8836 4553 8900
rect 4569 8836 4633 8900
rect 4649 8836 4713 8900
rect 4729 8836 4793 8900
rect 4809 8836 4873 8900
rect 0 8814 254 8836
rect 0 8750 264 8814
rect 281 8750 345 8814
rect 362 8750 426 8814
rect 443 8750 507 8814
rect 524 8750 588 8814
rect 605 8750 669 8814
rect 686 8750 750 8814
rect 767 8750 831 8814
rect 848 8750 912 8814
rect 929 8750 993 8814
rect 1010 8750 1074 8814
rect 1091 8750 1155 8814
rect 1172 8750 1236 8814
rect 1253 8750 1317 8814
rect 1334 8750 1398 8814
rect 1415 8750 1479 8814
rect 1496 8750 1560 8814
rect 1577 8750 1641 8814
rect 1658 8750 1722 8814
rect 1739 8750 1803 8814
rect 1820 8750 1884 8814
rect 1901 8750 1965 8814
rect 1982 8750 2046 8814
rect 2063 8750 2127 8814
rect 2144 8750 2208 8814
rect 2225 8750 2289 8814
rect 2306 8750 2370 8814
rect 2387 8750 2451 8814
rect 2468 8750 2532 8814
rect 2549 8750 2613 8814
rect 2630 8750 2694 8814
rect 2711 8750 2775 8814
rect 2792 8750 2856 8814
rect 2873 8750 2937 8814
rect 2954 8750 3018 8814
rect 3035 8750 3099 8814
rect 3116 8750 3180 8814
rect 3197 8750 3261 8814
rect 3278 8750 3342 8814
rect 3359 8750 3423 8814
rect 3440 8750 3504 8814
rect 3521 8750 3585 8814
rect 3602 8750 3666 8814
rect 3683 8750 3747 8814
rect 3764 8750 3828 8814
rect 3845 8750 3909 8814
rect 3926 8750 3990 8814
rect 4007 8750 4071 8814
rect 4088 8750 4152 8814
rect 4169 8750 4233 8814
rect 4249 8750 4313 8814
rect 4329 8750 4393 8814
rect 4409 8750 4473 8814
rect 4489 8750 4553 8814
rect 4569 8750 4633 8814
rect 4649 8750 4713 8814
rect 4729 8750 4793 8814
rect 4809 8750 4873 8814
rect 0 8728 254 8750
rect 0 8664 264 8728
rect 281 8664 345 8728
rect 362 8664 426 8728
rect 443 8664 507 8728
rect 524 8664 588 8728
rect 605 8664 669 8728
rect 686 8664 750 8728
rect 767 8664 831 8728
rect 848 8664 912 8728
rect 929 8664 993 8728
rect 1010 8664 1074 8728
rect 1091 8664 1155 8728
rect 1172 8664 1236 8728
rect 1253 8664 1317 8728
rect 1334 8664 1398 8728
rect 1415 8664 1479 8728
rect 1496 8664 1560 8728
rect 1577 8664 1641 8728
rect 1658 8664 1722 8728
rect 1739 8664 1803 8728
rect 1820 8664 1884 8728
rect 1901 8664 1965 8728
rect 1982 8664 2046 8728
rect 2063 8664 2127 8728
rect 2144 8664 2208 8728
rect 2225 8664 2289 8728
rect 2306 8664 2370 8728
rect 2387 8664 2451 8728
rect 2468 8664 2532 8728
rect 2549 8664 2613 8728
rect 2630 8664 2694 8728
rect 2711 8664 2775 8728
rect 2792 8664 2856 8728
rect 2873 8664 2937 8728
rect 2954 8664 3018 8728
rect 3035 8664 3099 8728
rect 3116 8664 3180 8728
rect 3197 8664 3261 8728
rect 3278 8664 3342 8728
rect 3359 8664 3423 8728
rect 3440 8664 3504 8728
rect 3521 8664 3585 8728
rect 3602 8664 3666 8728
rect 3683 8664 3747 8728
rect 3764 8664 3828 8728
rect 3845 8664 3909 8728
rect 3926 8664 3990 8728
rect 4007 8664 4071 8728
rect 4088 8664 4152 8728
rect 4169 8664 4233 8728
rect 4249 8664 4313 8728
rect 4329 8664 4393 8728
rect 4409 8664 4473 8728
rect 4489 8664 4553 8728
rect 4569 8664 4633 8728
rect 4649 8664 4713 8728
rect 4729 8664 4793 8728
rect 4809 8664 4873 8728
rect 0 8642 254 8664
rect 0 8578 264 8642
rect 281 8578 345 8642
rect 362 8578 426 8642
rect 443 8578 507 8642
rect 524 8578 588 8642
rect 605 8578 669 8642
rect 686 8578 750 8642
rect 767 8578 831 8642
rect 848 8578 912 8642
rect 929 8578 993 8642
rect 1010 8578 1074 8642
rect 1091 8578 1155 8642
rect 1172 8578 1236 8642
rect 1253 8578 1317 8642
rect 1334 8578 1398 8642
rect 1415 8578 1479 8642
rect 1496 8578 1560 8642
rect 1577 8578 1641 8642
rect 1658 8578 1722 8642
rect 1739 8578 1803 8642
rect 1820 8578 1884 8642
rect 1901 8578 1965 8642
rect 1982 8578 2046 8642
rect 2063 8578 2127 8642
rect 2144 8578 2208 8642
rect 2225 8578 2289 8642
rect 2306 8578 2370 8642
rect 2387 8578 2451 8642
rect 2468 8578 2532 8642
rect 2549 8578 2613 8642
rect 2630 8578 2694 8642
rect 2711 8578 2775 8642
rect 2792 8578 2856 8642
rect 2873 8578 2937 8642
rect 2954 8578 3018 8642
rect 3035 8578 3099 8642
rect 3116 8578 3180 8642
rect 3197 8578 3261 8642
rect 3278 8578 3342 8642
rect 3359 8578 3423 8642
rect 3440 8578 3504 8642
rect 3521 8578 3585 8642
rect 3602 8578 3666 8642
rect 3683 8578 3747 8642
rect 3764 8578 3828 8642
rect 3845 8578 3909 8642
rect 3926 8578 3990 8642
rect 4007 8578 4071 8642
rect 4088 8578 4152 8642
rect 4169 8578 4233 8642
rect 4249 8578 4313 8642
rect 4329 8578 4393 8642
rect 4409 8578 4473 8642
rect 4489 8578 4553 8642
rect 4569 8578 4633 8642
rect 4649 8578 4713 8642
rect 4729 8578 4793 8642
rect 4809 8578 4873 8642
rect 0 8556 254 8578
rect 0 8492 264 8556
rect 281 8492 345 8556
rect 362 8492 426 8556
rect 443 8492 507 8556
rect 524 8492 588 8556
rect 605 8492 669 8556
rect 686 8492 750 8556
rect 767 8492 831 8556
rect 848 8492 912 8556
rect 929 8492 993 8556
rect 1010 8492 1074 8556
rect 1091 8492 1155 8556
rect 1172 8492 1236 8556
rect 1253 8492 1317 8556
rect 1334 8492 1398 8556
rect 1415 8492 1479 8556
rect 1496 8492 1560 8556
rect 1577 8492 1641 8556
rect 1658 8492 1722 8556
rect 1739 8492 1803 8556
rect 1820 8492 1884 8556
rect 1901 8492 1965 8556
rect 1982 8492 2046 8556
rect 2063 8492 2127 8556
rect 2144 8492 2208 8556
rect 2225 8492 2289 8556
rect 2306 8492 2370 8556
rect 2387 8492 2451 8556
rect 2468 8492 2532 8556
rect 2549 8492 2613 8556
rect 2630 8492 2694 8556
rect 2711 8492 2775 8556
rect 2792 8492 2856 8556
rect 2873 8492 2937 8556
rect 2954 8492 3018 8556
rect 3035 8492 3099 8556
rect 3116 8492 3180 8556
rect 3197 8492 3261 8556
rect 3278 8492 3342 8556
rect 3359 8492 3423 8556
rect 3440 8492 3504 8556
rect 3521 8492 3585 8556
rect 3602 8492 3666 8556
rect 3683 8492 3747 8556
rect 3764 8492 3828 8556
rect 3845 8492 3909 8556
rect 3926 8492 3990 8556
rect 4007 8492 4071 8556
rect 4088 8492 4152 8556
rect 4169 8492 4233 8556
rect 4249 8492 4313 8556
rect 4329 8492 4393 8556
rect 4409 8492 4473 8556
rect 4489 8492 4553 8556
rect 4569 8492 4633 8556
rect 4649 8492 4713 8556
rect 4729 8492 4793 8556
rect 4809 8492 4873 8556
rect 0 8470 254 8492
rect 0 8406 264 8470
rect 281 8406 345 8470
rect 362 8406 426 8470
rect 443 8406 507 8470
rect 524 8406 588 8470
rect 605 8406 669 8470
rect 686 8406 750 8470
rect 767 8406 831 8470
rect 848 8406 912 8470
rect 929 8406 993 8470
rect 1010 8406 1074 8470
rect 1091 8406 1155 8470
rect 1172 8406 1236 8470
rect 1253 8406 1317 8470
rect 1334 8406 1398 8470
rect 1415 8406 1479 8470
rect 1496 8406 1560 8470
rect 1577 8406 1641 8470
rect 1658 8406 1722 8470
rect 1739 8406 1803 8470
rect 1820 8406 1884 8470
rect 1901 8406 1965 8470
rect 1982 8406 2046 8470
rect 2063 8406 2127 8470
rect 2144 8406 2208 8470
rect 2225 8406 2289 8470
rect 2306 8406 2370 8470
rect 2387 8406 2451 8470
rect 2468 8406 2532 8470
rect 2549 8406 2613 8470
rect 2630 8406 2694 8470
rect 2711 8406 2775 8470
rect 2792 8406 2856 8470
rect 2873 8406 2937 8470
rect 2954 8406 3018 8470
rect 3035 8406 3099 8470
rect 3116 8406 3180 8470
rect 3197 8406 3261 8470
rect 3278 8406 3342 8470
rect 3359 8406 3423 8470
rect 3440 8406 3504 8470
rect 3521 8406 3585 8470
rect 3602 8406 3666 8470
rect 3683 8406 3747 8470
rect 3764 8406 3828 8470
rect 3845 8406 3909 8470
rect 3926 8406 3990 8470
rect 4007 8406 4071 8470
rect 4088 8406 4152 8470
rect 4169 8406 4233 8470
rect 4249 8406 4313 8470
rect 4329 8406 4393 8470
rect 4409 8406 4473 8470
rect 4489 8406 4553 8470
rect 4569 8406 4633 8470
rect 4649 8406 4713 8470
rect 4729 8406 4793 8470
rect 4809 8406 4873 8470
rect 0 8384 254 8406
rect 0 8320 264 8384
rect 281 8320 345 8384
rect 362 8320 426 8384
rect 443 8320 507 8384
rect 524 8320 588 8384
rect 605 8320 669 8384
rect 686 8320 750 8384
rect 767 8320 831 8384
rect 848 8320 912 8384
rect 929 8320 993 8384
rect 1010 8320 1074 8384
rect 1091 8320 1155 8384
rect 1172 8320 1236 8384
rect 1253 8320 1317 8384
rect 1334 8320 1398 8384
rect 1415 8320 1479 8384
rect 1496 8320 1560 8384
rect 1577 8320 1641 8384
rect 1658 8320 1722 8384
rect 1739 8320 1803 8384
rect 1820 8320 1884 8384
rect 1901 8320 1965 8384
rect 1982 8320 2046 8384
rect 2063 8320 2127 8384
rect 2144 8320 2208 8384
rect 2225 8320 2289 8384
rect 2306 8320 2370 8384
rect 2387 8320 2451 8384
rect 2468 8320 2532 8384
rect 2549 8320 2613 8384
rect 2630 8320 2694 8384
rect 2711 8320 2775 8384
rect 2792 8320 2856 8384
rect 2873 8320 2937 8384
rect 2954 8320 3018 8384
rect 3035 8320 3099 8384
rect 3116 8320 3180 8384
rect 3197 8320 3261 8384
rect 3278 8320 3342 8384
rect 3359 8320 3423 8384
rect 3440 8320 3504 8384
rect 3521 8320 3585 8384
rect 3602 8320 3666 8384
rect 3683 8320 3747 8384
rect 3764 8320 3828 8384
rect 3845 8320 3909 8384
rect 3926 8320 3990 8384
rect 4007 8320 4071 8384
rect 4088 8320 4152 8384
rect 4169 8320 4233 8384
rect 4249 8320 4313 8384
rect 4329 8320 4393 8384
rect 4409 8320 4473 8384
rect 4489 8320 4553 8384
rect 4569 8320 4633 8384
rect 4649 8320 4713 8384
rect 4729 8320 4793 8384
rect 4809 8320 4873 8384
rect 0 8317 254 8320
rect 14746 8317 15000 9247
rect 0 7347 254 8037
rect 14746 7347 15000 8037
rect 0 6377 254 7067
rect 14746 6377 15000 7067
rect 0 5167 254 6097
rect 14746 5167 15000 6097
rect 0 3957 254 4887
rect 14746 3957 15000 4887
rect 0 2987 193 3677
rect 14807 2987 15000 3677
rect 0 1777 254 2707
rect 14746 1777 15000 2707
rect 0 407 254 1497
rect 14746 407 15000 1497
<< obsm4 >>
rect 334 35077 14666 40000
rect 193 19080 14807 35077
rect 334 13927 14666 19080
rect 193 13787 14807 13927
rect 334 12737 14666 13787
rect 193 12617 14807 12737
rect 334 11567 14666 12617
rect 193 11427 14807 11567
rect 334 10349 14666 10545
rect 193 9327 14807 9467
rect 334 9244 14666 9327
rect 345 9180 362 9244
rect 426 9180 443 9244
rect 507 9180 524 9244
rect 588 9180 605 9244
rect 669 9180 686 9244
rect 750 9180 767 9244
rect 831 9180 848 9244
rect 912 9180 929 9244
rect 993 9180 1010 9244
rect 1074 9180 1091 9244
rect 1155 9180 1172 9244
rect 1236 9180 1253 9244
rect 1317 9180 1334 9244
rect 1398 9180 1415 9244
rect 1479 9180 1496 9244
rect 1560 9180 1577 9244
rect 1641 9180 1658 9244
rect 1722 9180 1739 9244
rect 1803 9180 1820 9244
rect 1884 9180 1901 9244
rect 1965 9180 1982 9244
rect 2046 9180 2063 9244
rect 2127 9180 2144 9244
rect 2208 9180 2225 9244
rect 2289 9180 2306 9244
rect 2370 9180 2387 9244
rect 2451 9180 2468 9244
rect 2532 9180 2549 9244
rect 2613 9180 2630 9244
rect 2694 9180 2711 9244
rect 2775 9180 2792 9244
rect 2856 9180 2873 9244
rect 2937 9180 2954 9244
rect 3018 9180 3035 9244
rect 3099 9180 3116 9244
rect 3180 9180 3197 9244
rect 3261 9180 3278 9244
rect 3342 9180 3359 9244
rect 3423 9180 3440 9244
rect 3504 9180 3521 9244
rect 3585 9180 3602 9244
rect 3666 9180 3683 9244
rect 3747 9180 3764 9244
rect 3828 9180 3845 9244
rect 3909 9180 3926 9244
rect 3990 9180 4007 9244
rect 4071 9180 4088 9244
rect 4152 9180 4169 9244
rect 4233 9180 4249 9244
rect 4313 9180 4329 9244
rect 4393 9180 4409 9244
rect 4473 9180 4489 9244
rect 4553 9180 4569 9244
rect 4633 9180 4649 9244
rect 4713 9180 4729 9244
rect 4793 9180 4809 9244
rect 4873 9180 14666 9244
rect 334 9158 14666 9180
rect 345 9094 362 9158
rect 426 9094 443 9158
rect 507 9094 524 9158
rect 588 9094 605 9158
rect 669 9094 686 9158
rect 750 9094 767 9158
rect 831 9094 848 9158
rect 912 9094 929 9158
rect 993 9094 1010 9158
rect 1074 9094 1091 9158
rect 1155 9094 1172 9158
rect 1236 9094 1253 9158
rect 1317 9094 1334 9158
rect 1398 9094 1415 9158
rect 1479 9094 1496 9158
rect 1560 9094 1577 9158
rect 1641 9094 1658 9158
rect 1722 9094 1739 9158
rect 1803 9094 1820 9158
rect 1884 9094 1901 9158
rect 1965 9094 1982 9158
rect 2046 9094 2063 9158
rect 2127 9094 2144 9158
rect 2208 9094 2225 9158
rect 2289 9094 2306 9158
rect 2370 9094 2387 9158
rect 2451 9094 2468 9158
rect 2532 9094 2549 9158
rect 2613 9094 2630 9158
rect 2694 9094 2711 9158
rect 2775 9094 2792 9158
rect 2856 9094 2873 9158
rect 2937 9094 2954 9158
rect 3018 9094 3035 9158
rect 3099 9094 3116 9158
rect 3180 9094 3197 9158
rect 3261 9094 3278 9158
rect 3342 9094 3359 9158
rect 3423 9094 3440 9158
rect 3504 9094 3521 9158
rect 3585 9094 3602 9158
rect 3666 9094 3683 9158
rect 3747 9094 3764 9158
rect 3828 9094 3845 9158
rect 3909 9094 3926 9158
rect 3990 9094 4007 9158
rect 4071 9094 4088 9158
rect 4152 9094 4169 9158
rect 4233 9094 4249 9158
rect 4313 9094 4329 9158
rect 4393 9094 4409 9158
rect 4473 9094 4489 9158
rect 4553 9094 4569 9158
rect 4633 9094 4649 9158
rect 4713 9094 4729 9158
rect 4793 9094 4809 9158
rect 4873 9094 14666 9158
rect 334 9072 14666 9094
rect 345 9008 362 9072
rect 426 9008 443 9072
rect 507 9008 524 9072
rect 588 9008 605 9072
rect 669 9008 686 9072
rect 750 9008 767 9072
rect 831 9008 848 9072
rect 912 9008 929 9072
rect 993 9008 1010 9072
rect 1074 9008 1091 9072
rect 1155 9008 1172 9072
rect 1236 9008 1253 9072
rect 1317 9008 1334 9072
rect 1398 9008 1415 9072
rect 1479 9008 1496 9072
rect 1560 9008 1577 9072
rect 1641 9008 1658 9072
rect 1722 9008 1739 9072
rect 1803 9008 1820 9072
rect 1884 9008 1901 9072
rect 1965 9008 1982 9072
rect 2046 9008 2063 9072
rect 2127 9008 2144 9072
rect 2208 9008 2225 9072
rect 2289 9008 2306 9072
rect 2370 9008 2387 9072
rect 2451 9008 2468 9072
rect 2532 9008 2549 9072
rect 2613 9008 2630 9072
rect 2694 9008 2711 9072
rect 2775 9008 2792 9072
rect 2856 9008 2873 9072
rect 2937 9008 2954 9072
rect 3018 9008 3035 9072
rect 3099 9008 3116 9072
rect 3180 9008 3197 9072
rect 3261 9008 3278 9072
rect 3342 9008 3359 9072
rect 3423 9008 3440 9072
rect 3504 9008 3521 9072
rect 3585 9008 3602 9072
rect 3666 9008 3683 9072
rect 3747 9008 3764 9072
rect 3828 9008 3845 9072
rect 3909 9008 3926 9072
rect 3990 9008 4007 9072
rect 4071 9008 4088 9072
rect 4152 9008 4169 9072
rect 4233 9008 4249 9072
rect 4313 9008 4329 9072
rect 4393 9008 4409 9072
rect 4473 9008 4489 9072
rect 4553 9008 4569 9072
rect 4633 9008 4649 9072
rect 4713 9008 4729 9072
rect 4793 9008 4809 9072
rect 4873 9008 14666 9072
rect 334 8986 14666 9008
rect 345 8922 362 8986
rect 426 8922 443 8986
rect 507 8922 524 8986
rect 588 8922 605 8986
rect 669 8922 686 8986
rect 750 8922 767 8986
rect 831 8922 848 8986
rect 912 8922 929 8986
rect 993 8922 1010 8986
rect 1074 8922 1091 8986
rect 1155 8922 1172 8986
rect 1236 8922 1253 8986
rect 1317 8922 1334 8986
rect 1398 8922 1415 8986
rect 1479 8922 1496 8986
rect 1560 8922 1577 8986
rect 1641 8922 1658 8986
rect 1722 8922 1739 8986
rect 1803 8922 1820 8986
rect 1884 8922 1901 8986
rect 1965 8922 1982 8986
rect 2046 8922 2063 8986
rect 2127 8922 2144 8986
rect 2208 8922 2225 8986
rect 2289 8922 2306 8986
rect 2370 8922 2387 8986
rect 2451 8922 2468 8986
rect 2532 8922 2549 8986
rect 2613 8922 2630 8986
rect 2694 8922 2711 8986
rect 2775 8922 2792 8986
rect 2856 8922 2873 8986
rect 2937 8922 2954 8986
rect 3018 8922 3035 8986
rect 3099 8922 3116 8986
rect 3180 8922 3197 8986
rect 3261 8922 3278 8986
rect 3342 8922 3359 8986
rect 3423 8922 3440 8986
rect 3504 8922 3521 8986
rect 3585 8922 3602 8986
rect 3666 8922 3683 8986
rect 3747 8922 3764 8986
rect 3828 8922 3845 8986
rect 3909 8922 3926 8986
rect 3990 8922 4007 8986
rect 4071 8922 4088 8986
rect 4152 8922 4169 8986
rect 4233 8922 4249 8986
rect 4313 8922 4329 8986
rect 4393 8922 4409 8986
rect 4473 8922 4489 8986
rect 4553 8922 4569 8986
rect 4633 8922 4649 8986
rect 4713 8922 4729 8986
rect 4793 8922 4809 8986
rect 4873 8922 14666 8986
rect 334 8900 14666 8922
rect 345 8836 362 8900
rect 426 8836 443 8900
rect 507 8836 524 8900
rect 588 8836 605 8900
rect 669 8836 686 8900
rect 750 8836 767 8900
rect 831 8836 848 8900
rect 912 8836 929 8900
rect 993 8836 1010 8900
rect 1074 8836 1091 8900
rect 1155 8836 1172 8900
rect 1236 8836 1253 8900
rect 1317 8836 1334 8900
rect 1398 8836 1415 8900
rect 1479 8836 1496 8900
rect 1560 8836 1577 8900
rect 1641 8836 1658 8900
rect 1722 8836 1739 8900
rect 1803 8836 1820 8900
rect 1884 8836 1901 8900
rect 1965 8836 1982 8900
rect 2046 8836 2063 8900
rect 2127 8836 2144 8900
rect 2208 8836 2225 8900
rect 2289 8836 2306 8900
rect 2370 8836 2387 8900
rect 2451 8836 2468 8900
rect 2532 8836 2549 8900
rect 2613 8836 2630 8900
rect 2694 8836 2711 8900
rect 2775 8836 2792 8900
rect 2856 8836 2873 8900
rect 2937 8836 2954 8900
rect 3018 8836 3035 8900
rect 3099 8836 3116 8900
rect 3180 8836 3197 8900
rect 3261 8836 3278 8900
rect 3342 8836 3359 8900
rect 3423 8836 3440 8900
rect 3504 8836 3521 8900
rect 3585 8836 3602 8900
rect 3666 8836 3683 8900
rect 3747 8836 3764 8900
rect 3828 8836 3845 8900
rect 3909 8836 3926 8900
rect 3990 8836 4007 8900
rect 4071 8836 4088 8900
rect 4152 8836 4169 8900
rect 4233 8836 4249 8900
rect 4313 8836 4329 8900
rect 4393 8836 4409 8900
rect 4473 8836 4489 8900
rect 4553 8836 4569 8900
rect 4633 8836 4649 8900
rect 4713 8836 4729 8900
rect 4793 8836 4809 8900
rect 4873 8836 14666 8900
rect 334 8814 14666 8836
rect 345 8750 362 8814
rect 426 8750 443 8814
rect 507 8750 524 8814
rect 588 8750 605 8814
rect 669 8750 686 8814
rect 750 8750 767 8814
rect 831 8750 848 8814
rect 912 8750 929 8814
rect 993 8750 1010 8814
rect 1074 8750 1091 8814
rect 1155 8750 1172 8814
rect 1236 8750 1253 8814
rect 1317 8750 1334 8814
rect 1398 8750 1415 8814
rect 1479 8750 1496 8814
rect 1560 8750 1577 8814
rect 1641 8750 1658 8814
rect 1722 8750 1739 8814
rect 1803 8750 1820 8814
rect 1884 8750 1901 8814
rect 1965 8750 1982 8814
rect 2046 8750 2063 8814
rect 2127 8750 2144 8814
rect 2208 8750 2225 8814
rect 2289 8750 2306 8814
rect 2370 8750 2387 8814
rect 2451 8750 2468 8814
rect 2532 8750 2549 8814
rect 2613 8750 2630 8814
rect 2694 8750 2711 8814
rect 2775 8750 2792 8814
rect 2856 8750 2873 8814
rect 2937 8750 2954 8814
rect 3018 8750 3035 8814
rect 3099 8750 3116 8814
rect 3180 8750 3197 8814
rect 3261 8750 3278 8814
rect 3342 8750 3359 8814
rect 3423 8750 3440 8814
rect 3504 8750 3521 8814
rect 3585 8750 3602 8814
rect 3666 8750 3683 8814
rect 3747 8750 3764 8814
rect 3828 8750 3845 8814
rect 3909 8750 3926 8814
rect 3990 8750 4007 8814
rect 4071 8750 4088 8814
rect 4152 8750 4169 8814
rect 4233 8750 4249 8814
rect 4313 8750 4329 8814
rect 4393 8750 4409 8814
rect 4473 8750 4489 8814
rect 4553 8750 4569 8814
rect 4633 8750 4649 8814
rect 4713 8750 4729 8814
rect 4793 8750 4809 8814
rect 4873 8750 14666 8814
rect 334 8728 14666 8750
rect 345 8664 362 8728
rect 426 8664 443 8728
rect 507 8664 524 8728
rect 588 8664 605 8728
rect 669 8664 686 8728
rect 750 8664 767 8728
rect 831 8664 848 8728
rect 912 8664 929 8728
rect 993 8664 1010 8728
rect 1074 8664 1091 8728
rect 1155 8664 1172 8728
rect 1236 8664 1253 8728
rect 1317 8664 1334 8728
rect 1398 8664 1415 8728
rect 1479 8664 1496 8728
rect 1560 8664 1577 8728
rect 1641 8664 1658 8728
rect 1722 8664 1739 8728
rect 1803 8664 1820 8728
rect 1884 8664 1901 8728
rect 1965 8664 1982 8728
rect 2046 8664 2063 8728
rect 2127 8664 2144 8728
rect 2208 8664 2225 8728
rect 2289 8664 2306 8728
rect 2370 8664 2387 8728
rect 2451 8664 2468 8728
rect 2532 8664 2549 8728
rect 2613 8664 2630 8728
rect 2694 8664 2711 8728
rect 2775 8664 2792 8728
rect 2856 8664 2873 8728
rect 2937 8664 2954 8728
rect 3018 8664 3035 8728
rect 3099 8664 3116 8728
rect 3180 8664 3197 8728
rect 3261 8664 3278 8728
rect 3342 8664 3359 8728
rect 3423 8664 3440 8728
rect 3504 8664 3521 8728
rect 3585 8664 3602 8728
rect 3666 8664 3683 8728
rect 3747 8664 3764 8728
rect 3828 8664 3845 8728
rect 3909 8664 3926 8728
rect 3990 8664 4007 8728
rect 4071 8664 4088 8728
rect 4152 8664 4169 8728
rect 4233 8664 4249 8728
rect 4313 8664 4329 8728
rect 4393 8664 4409 8728
rect 4473 8664 4489 8728
rect 4553 8664 4569 8728
rect 4633 8664 4649 8728
rect 4713 8664 4729 8728
rect 4793 8664 4809 8728
rect 4873 8664 14666 8728
rect 334 8642 14666 8664
rect 345 8578 362 8642
rect 426 8578 443 8642
rect 507 8578 524 8642
rect 588 8578 605 8642
rect 669 8578 686 8642
rect 750 8578 767 8642
rect 831 8578 848 8642
rect 912 8578 929 8642
rect 993 8578 1010 8642
rect 1074 8578 1091 8642
rect 1155 8578 1172 8642
rect 1236 8578 1253 8642
rect 1317 8578 1334 8642
rect 1398 8578 1415 8642
rect 1479 8578 1496 8642
rect 1560 8578 1577 8642
rect 1641 8578 1658 8642
rect 1722 8578 1739 8642
rect 1803 8578 1820 8642
rect 1884 8578 1901 8642
rect 1965 8578 1982 8642
rect 2046 8578 2063 8642
rect 2127 8578 2144 8642
rect 2208 8578 2225 8642
rect 2289 8578 2306 8642
rect 2370 8578 2387 8642
rect 2451 8578 2468 8642
rect 2532 8578 2549 8642
rect 2613 8578 2630 8642
rect 2694 8578 2711 8642
rect 2775 8578 2792 8642
rect 2856 8578 2873 8642
rect 2937 8578 2954 8642
rect 3018 8578 3035 8642
rect 3099 8578 3116 8642
rect 3180 8578 3197 8642
rect 3261 8578 3278 8642
rect 3342 8578 3359 8642
rect 3423 8578 3440 8642
rect 3504 8578 3521 8642
rect 3585 8578 3602 8642
rect 3666 8578 3683 8642
rect 3747 8578 3764 8642
rect 3828 8578 3845 8642
rect 3909 8578 3926 8642
rect 3990 8578 4007 8642
rect 4071 8578 4088 8642
rect 4152 8578 4169 8642
rect 4233 8578 4249 8642
rect 4313 8578 4329 8642
rect 4393 8578 4409 8642
rect 4473 8578 4489 8642
rect 4553 8578 4569 8642
rect 4633 8578 4649 8642
rect 4713 8578 4729 8642
rect 4793 8578 4809 8642
rect 4873 8578 14666 8642
rect 334 8556 14666 8578
rect 345 8492 362 8556
rect 426 8492 443 8556
rect 507 8492 524 8556
rect 588 8492 605 8556
rect 669 8492 686 8556
rect 750 8492 767 8556
rect 831 8492 848 8556
rect 912 8492 929 8556
rect 993 8492 1010 8556
rect 1074 8492 1091 8556
rect 1155 8492 1172 8556
rect 1236 8492 1253 8556
rect 1317 8492 1334 8556
rect 1398 8492 1415 8556
rect 1479 8492 1496 8556
rect 1560 8492 1577 8556
rect 1641 8492 1658 8556
rect 1722 8492 1739 8556
rect 1803 8492 1820 8556
rect 1884 8492 1901 8556
rect 1965 8492 1982 8556
rect 2046 8492 2063 8556
rect 2127 8492 2144 8556
rect 2208 8492 2225 8556
rect 2289 8492 2306 8556
rect 2370 8492 2387 8556
rect 2451 8492 2468 8556
rect 2532 8492 2549 8556
rect 2613 8492 2630 8556
rect 2694 8492 2711 8556
rect 2775 8492 2792 8556
rect 2856 8492 2873 8556
rect 2937 8492 2954 8556
rect 3018 8492 3035 8556
rect 3099 8492 3116 8556
rect 3180 8492 3197 8556
rect 3261 8492 3278 8556
rect 3342 8492 3359 8556
rect 3423 8492 3440 8556
rect 3504 8492 3521 8556
rect 3585 8492 3602 8556
rect 3666 8492 3683 8556
rect 3747 8492 3764 8556
rect 3828 8492 3845 8556
rect 3909 8492 3926 8556
rect 3990 8492 4007 8556
rect 4071 8492 4088 8556
rect 4152 8492 4169 8556
rect 4233 8492 4249 8556
rect 4313 8492 4329 8556
rect 4393 8492 4409 8556
rect 4473 8492 4489 8556
rect 4553 8492 4569 8556
rect 4633 8492 4649 8556
rect 4713 8492 4729 8556
rect 4793 8492 4809 8556
rect 4873 8492 14666 8556
rect 334 8470 14666 8492
rect 345 8406 362 8470
rect 426 8406 443 8470
rect 507 8406 524 8470
rect 588 8406 605 8470
rect 669 8406 686 8470
rect 750 8406 767 8470
rect 831 8406 848 8470
rect 912 8406 929 8470
rect 993 8406 1010 8470
rect 1074 8406 1091 8470
rect 1155 8406 1172 8470
rect 1236 8406 1253 8470
rect 1317 8406 1334 8470
rect 1398 8406 1415 8470
rect 1479 8406 1496 8470
rect 1560 8406 1577 8470
rect 1641 8406 1658 8470
rect 1722 8406 1739 8470
rect 1803 8406 1820 8470
rect 1884 8406 1901 8470
rect 1965 8406 1982 8470
rect 2046 8406 2063 8470
rect 2127 8406 2144 8470
rect 2208 8406 2225 8470
rect 2289 8406 2306 8470
rect 2370 8406 2387 8470
rect 2451 8406 2468 8470
rect 2532 8406 2549 8470
rect 2613 8406 2630 8470
rect 2694 8406 2711 8470
rect 2775 8406 2792 8470
rect 2856 8406 2873 8470
rect 2937 8406 2954 8470
rect 3018 8406 3035 8470
rect 3099 8406 3116 8470
rect 3180 8406 3197 8470
rect 3261 8406 3278 8470
rect 3342 8406 3359 8470
rect 3423 8406 3440 8470
rect 3504 8406 3521 8470
rect 3585 8406 3602 8470
rect 3666 8406 3683 8470
rect 3747 8406 3764 8470
rect 3828 8406 3845 8470
rect 3909 8406 3926 8470
rect 3990 8406 4007 8470
rect 4071 8406 4088 8470
rect 4152 8406 4169 8470
rect 4233 8406 4249 8470
rect 4313 8406 4329 8470
rect 4393 8406 4409 8470
rect 4473 8406 4489 8470
rect 4553 8406 4569 8470
rect 4633 8406 4649 8470
rect 4713 8406 4729 8470
rect 4793 8406 4809 8470
rect 4873 8406 14666 8470
rect 334 8384 14666 8406
rect 345 8320 362 8384
rect 426 8320 443 8384
rect 507 8320 524 8384
rect 588 8320 605 8384
rect 669 8320 686 8384
rect 750 8320 767 8384
rect 831 8320 848 8384
rect 912 8320 929 8384
rect 993 8320 1010 8384
rect 1074 8320 1091 8384
rect 1155 8320 1172 8384
rect 1236 8320 1253 8384
rect 1317 8320 1334 8384
rect 1398 8320 1415 8384
rect 1479 8320 1496 8384
rect 1560 8320 1577 8384
rect 1641 8320 1658 8384
rect 1722 8320 1739 8384
rect 1803 8320 1820 8384
rect 1884 8320 1901 8384
rect 1965 8320 1982 8384
rect 2046 8320 2063 8384
rect 2127 8320 2144 8384
rect 2208 8320 2225 8384
rect 2289 8320 2306 8384
rect 2370 8320 2387 8384
rect 2451 8320 2468 8384
rect 2532 8320 2549 8384
rect 2613 8320 2630 8384
rect 2694 8320 2711 8384
rect 2775 8320 2792 8384
rect 2856 8320 2873 8384
rect 2937 8320 2954 8384
rect 3018 8320 3035 8384
rect 3099 8320 3116 8384
rect 3180 8320 3197 8384
rect 3261 8320 3278 8384
rect 3342 8320 3359 8384
rect 3423 8320 3440 8384
rect 3504 8320 3521 8384
rect 3585 8320 3602 8384
rect 3666 8320 3683 8384
rect 3747 8320 3764 8384
rect 3828 8320 3845 8384
rect 3909 8320 3926 8384
rect 3990 8320 4007 8384
rect 4071 8320 4088 8384
rect 4152 8320 4169 8384
rect 4233 8320 4249 8384
rect 4313 8320 4329 8384
rect 4393 8320 4409 8384
rect 4473 8320 4489 8384
rect 4553 8320 4569 8384
rect 4633 8320 4649 8384
rect 4713 8320 4729 8384
rect 4793 8320 4809 8384
rect 4873 8320 14666 8384
rect 334 8237 14666 8320
rect 193 8117 14807 8237
rect 334 7267 14666 8117
rect 193 7147 14807 7267
rect 334 6297 14666 7147
rect 193 6177 14807 6297
rect 334 5087 14666 6177
rect 193 4967 14807 5087
rect 334 3877 14666 4967
rect 193 3757 14807 3877
rect 273 2907 14727 3757
rect 193 2787 14807 2907
rect 334 1697 14666 2787
rect 193 1577 14807 1697
rect 334 407 14666 1577
<< metal5 >>
rect 0 35157 254 40000
rect 14746 35157 15000 40000
rect 0 14007 254 18997
rect 0 12837 254 13687
rect 0 11667 254 12517
rect 0 9547 254 11347
rect 0 8337 254 9227
rect 0 7368 254 8017
rect 14746 14007 15000 18997
rect 14746 12837 15000 13687
rect 14746 11667 15000 12517
rect 14746 9547 15000 11347
rect 14746 8337 15000 9227
rect 14746 7368 15000 8017
rect 0 6397 254 7047
rect 0 5187 254 6077
rect 0 3977 254 4867
rect 14746 6397 15000 7047
rect 14746 5187 15000 6077
rect 14746 3977 15000 4867
rect 0 3007 193 3657
rect 14807 3007 15000 3657
rect 0 1797 254 2687
rect 0 427 254 1477
rect 14746 1797 15000 2687
rect 14746 427 15000 1477
<< obsm5 >>
rect 574 34837 14426 40000
rect 0 19317 15000 34837
rect 574 7368 14426 19317
rect 0 7367 15000 7368
rect 574 3657 14426 7367
rect 513 3007 14487 3657
rect 574 427 14426 3007
<< labels >>
rlabel metal5 s 0 12837 254 13687 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal5 s 14746 12837 15000 13687 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 14746 12817 15000 13707 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 0 12817 254 13707 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal5 s 14746 1797 15000 2687 6 VCCD
port 2 nsew power bidirectional
rlabel metal5 s 0 1797 254 2687 6 VCCD
port 2 nsew power bidirectional
rlabel metal4 s 14746 1777 15000 2707 6 VCCD
port 2 nsew power bidirectional
rlabel metal4 s 0 1777 254 2707 6 VCCD
port 2 nsew power bidirectional
rlabel metal5 s 14746 9547 15000 11347 6 VSSA
port 3 nsew ground bidirectional
rlabel metal5 s 14746 7368 15000 8017 6 VSSA
port 3 nsew ground bidirectional
rlabel metal5 s 0 9547 254 11347 6 VSSA
port 3 nsew ground bidirectional
rlabel metal5 s 0 7368 254 8017 6 VSSA
port 3 nsew ground bidirectional
rlabel metal4 s 14746 7347 15000 8037 6 VSSA
port 3 nsew ground bidirectional
rlabel metal4 s 0 9547 15000 9613 6 VSSA
port 3 nsew ground bidirectional
rlabel metal4 s 0 11281 15000 11347 6 VSSA
port 3 nsew ground bidirectional
rlabel metal4 s 14746 10329 15000 10565 6 VSSA
port 3 nsew ground bidirectional
rlabel metal4 s 0 10329 254 10565 6 VSSA
port 3 nsew ground bidirectional
rlabel metal4 s 0 7347 254 8037 6 VSSA
port 3 nsew ground bidirectional
rlabel metal5 s 14746 8337 15000 9227 6 VSSD
port 4 nsew ground bidirectional
rlabel metal5 s 0 8337 254 9227 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 14746 8317 15000 9247 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 0 8317 254 9247 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 10078 8318 14858 9246 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 14800 9192 14840 9232 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 14800 9106 14840 9146 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 14800 9020 14840 9060 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 14800 8934 14840 8974 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 14800 8848 14840 8888 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 14800 8762 14840 8802 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 14800 8676 14840 8716 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 14800 8590 14840 8630 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 14800 8504 14840 8544 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 14800 8418 14840 8458 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 14800 8332 14840 8372 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 14719 9192 14759 9232 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 14719 9106 14759 9146 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 14719 9020 14759 9060 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 14719 8934 14759 8974 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 14719 8848 14759 8888 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 14719 8762 14759 8802 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 14719 8676 14759 8716 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 14719 8590 14759 8630 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 14719 8504 14759 8544 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 14719 8418 14759 8458 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 14719 8332 14759 8372 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 14638 9192 14678 9232 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 14638 9106 14678 9146 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 14638 9020 14678 9060 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 14638 8934 14678 8974 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 14638 8848 14678 8888 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 14638 8762 14678 8802 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 14638 8676 14678 8716 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 14638 8590 14678 8630 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 14638 8504 14678 8544 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 14638 8418 14678 8458 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 14638 8332 14678 8372 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 14557 9192 14597 9232 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 14557 9106 14597 9146 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 14557 9020 14597 9060 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 14557 8934 14597 8974 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 14557 8848 14597 8888 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 14557 8762 14597 8802 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 14557 8676 14597 8716 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 14557 8590 14597 8630 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 14557 8504 14597 8544 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 14557 8418 14597 8458 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 14557 8332 14597 8372 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 14476 9192 14516 9232 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 14476 9106 14516 9146 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 14476 9020 14516 9060 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 14476 8934 14516 8974 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 14476 8848 14516 8888 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 14476 8762 14516 8802 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 14476 8676 14516 8716 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 14476 8590 14516 8630 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 14476 8504 14516 8544 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 14476 8418 14516 8458 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 14476 8332 14516 8372 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 14395 9192 14435 9232 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 14395 9106 14435 9146 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 14395 9020 14435 9060 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 14395 8934 14435 8974 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 14395 8848 14435 8888 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 14395 8762 14435 8802 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 14395 8676 14435 8716 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 14395 8590 14435 8630 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 14395 8504 14435 8544 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 14395 8418 14435 8458 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 14395 8332 14435 8372 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 14314 9192 14354 9232 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 14314 9106 14354 9146 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 14314 9020 14354 9060 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 14314 8934 14354 8974 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 14314 8848 14354 8888 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 14314 8762 14354 8802 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 14314 8676 14354 8716 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 14314 8590 14354 8630 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 14314 8504 14354 8544 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 14314 8418 14354 8458 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 14314 8332 14354 8372 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 14233 9192 14273 9232 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 14233 9106 14273 9146 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 14233 9020 14273 9060 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 14233 8934 14273 8974 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 14233 8848 14273 8888 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 14233 8762 14273 8802 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 14233 8676 14273 8716 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 14233 8590 14273 8630 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 14233 8504 14273 8544 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 14233 8418 14273 8458 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 14233 8332 14273 8372 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 14152 9192 14192 9232 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 14152 9106 14192 9146 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 14152 9020 14192 9060 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 14152 8934 14192 8974 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 14152 8848 14192 8888 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 14152 8762 14192 8802 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 14152 8676 14192 8716 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 14152 8590 14192 8630 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 14152 8504 14192 8544 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 14152 8418 14192 8458 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 14152 8332 14192 8372 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 14071 9192 14111 9232 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 14071 9106 14111 9146 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 14071 9020 14111 9060 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 14071 8934 14111 8974 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 14071 8848 14111 8888 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 14071 8762 14111 8802 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 14071 8676 14111 8716 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 14071 8590 14111 8630 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 14071 8504 14111 8544 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 14071 8418 14111 8458 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 14071 8332 14111 8372 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13990 9192 14030 9232 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13990 9106 14030 9146 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13990 9020 14030 9060 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13990 8934 14030 8974 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13990 8848 14030 8888 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13990 8762 14030 8802 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13990 8676 14030 8716 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13990 8590 14030 8630 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13990 8504 14030 8544 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13990 8418 14030 8458 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13990 8332 14030 8372 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13909 9192 13949 9232 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13909 9106 13949 9146 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13909 9020 13949 9060 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13909 8934 13949 8974 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13909 8848 13949 8888 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13909 8762 13949 8802 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13909 8676 13949 8716 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13909 8590 13949 8630 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13909 8504 13949 8544 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13909 8418 13949 8458 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13909 8332 13949 8372 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13828 9192 13868 9232 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13828 9106 13868 9146 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13828 9020 13868 9060 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13828 8934 13868 8974 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13828 8848 13868 8888 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13828 8762 13868 8802 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13828 8676 13868 8716 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13828 8590 13868 8630 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13828 8504 13868 8544 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13828 8418 13868 8458 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13828 8332 13868 8372 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13747 9192 13787 9232 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13747 9106 13787 9146 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13747 9020 13787 9060 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13747 8934 13787 8974 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13747 8848 13787 8888 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13747 8762 13787 8802 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13747 8676 13787 8716 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13747 8590 13787 8630 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13747 8504 13787 8544 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13747 8418 13787 8458 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13747 8332 13787 8372 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13666 9192 13706 9232 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13666 9106 13706 9146 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13666 9020 13706 9060 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13666 8934 13706 8974 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13666 8848 13706 8888 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13666 8762 13706 8802 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13666 8676 13706 8716 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13666 8590 13706 8630 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13666 8504 13706 8544 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13666 8418 13706 8458 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13666 8332 13706 8372 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13585 9192 13625 9232 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13585 9106 13625 9146 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13585 9020 13625 9060 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13585 8934 13625 8974 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13585 8848 13625 8888 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13585 8762 13625 8802 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13585 8676 13625 8716 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13585 8590 13625 8630 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13585 8504 13625 8544 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13585 8418 13625 8458 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13585 8332 13625 8372 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13504 9192 13544 9232 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13504 9106 13544 9146 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13504 9020 13544 9060 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13504 8934 13544 8974 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13504 8848 13544 8888 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13504 8762 13544 8802 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13504 8676 13544 8716 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13504 8590 13544 8630 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13504 8504 13544 8544 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13504 8418 13544 8458 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13504 8332 13544 8372 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13423 9192 13463 9232 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13423 9106 13463 9146 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13423 9020 13463 9060 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13423 8934 13463 8974 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13423 8848 13463 8888 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13423 8762 13463 8802 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13423 8676 13463 8716 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13423 8590 13463 8630 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13423 8504 13463 8544 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13423 8418 13463 8458 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13423 8332 13463 8372 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13342 9192 13382 9232 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13342 9106 13382 9146 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13342 9020 13382 9060 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13342 8934 13382 8974 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13342 8848 13382 8888 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13342 8762 13382 8802 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13342 8676 13382 8716 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13342 8590 13382 8630 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13342 8504 13382 8544 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13342 8418 13382 8458 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13342 8332 13382 8372 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13261 9192 13301 9232 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13261 9106 13301 9146 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13261 9020 13301 9060 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13261 8934 13301 8974 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13261 8848 13301 8888 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13261 8762 13301 8802 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13261 8676 13301 8716 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13261 8590 13301 8630 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13261 8504 13301 8544 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13261 8418 13301 8458 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13261 8332 13301 8372 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13180 9192 13220 9232 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13180 9106 13220 9146 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13180 9020 13220 9060 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13180 8934 13220 8974 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13180 8848 13220 8888 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13180 8762 13220 8802 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13180 8676 13220 8716 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13180 8590 13220 8630 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13180 8504 13220 8544 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13180 8418 13220 8458 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13180 8332 13220 8372 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13099 9192 13139 9232 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13099 9106 13139 9146 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13099 9020 13139 9060 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13099 8934 13139 8974 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13099 8848 13139 8888 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13099 8762 13139 8802 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13099 8676 13139 8716 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13099 8590 13139 8630 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13099 8504 13139 8544 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13099 8418 13139 8458 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13099 8332 13139 8372 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13018 9192 13058 9232 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13018 9106 13058 9146 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13018 9020 13058 9060 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13018 8934 13058 8974 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13018 8848 13058 8888 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13018 8762 13058 8802 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13018 8676 13058 8716 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13018 8590 13058 8630 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13018 8504 13058 8544 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13018 8418 13058 8458 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13018 8332 13058 8372 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 12937 9192 12977 9232 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 12937 9106 12977 9146 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 12937 9020 12977 9060 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 12937 8934 12977 8974 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 12937 8848 12977 8888 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 12937 8762 12977 8802 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 12937 8676 12977 8716 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 12937 8590 12977 8630 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 12937 8504 12977 8544 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 12937 8418 12977 8458 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 12937 8332 12977 8372 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 12856 9192 12896 9232 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 12856 9106 12896 9146 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 12856 9020 12896 9060 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 12856 8934 12896 8974 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 12856 8848 12896 8888 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 12856 8762 12896 8802 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 12856 8676 12896 8716 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 12856 8590 12896 8630 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 12856 8504 12896 8544 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 12856 8418 12896 8458 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 12856 8332 12896 8372 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 12775 9192 12815 9232 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 12775 9106 12815 9146 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 12775 9020 12815 9060 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 12775 8934 12815 8974 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 12775 8848 12815 8888 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 12775 8762 12815 8802 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 12775 8676 12815 8716 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 12775 8590 12815 8630 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 12775 8504 12815 8544 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 12775 8418 12815 8458 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 12775 8332 12815 8372 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 12694 9192 12734 9232 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 12694 9106 12734 9146 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 12694 9020 12734 9060 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 12694 8934 12734 8974 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 12694 8848 12734 8888 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 12694 8762 12734 8802 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 12694 8676 12734 8716 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 12694 8590 12734 8630 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 12694 8504 12734 8544 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 12694 8418 12734 8458 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 12694 8332 12734 8372 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 12613 9192 12653 9232 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 12613 9106 12653 9146 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 12613 9020 12653 9060 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 12613 8934 12653 8974 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 12613 8848 12653 8888 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 12613 8762 12653 8802 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 12613 8676 12653 8716 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 12613 8590 12653 8630 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 12613 8504 12653 8544 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 12613 8418 12653 8458 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 12613 8332 12653 8372 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 12532 9192 12572 9232 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 12532 9106 12572 9146 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 12532 9020 12572 9060 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 12532 8934 12572 8974 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 12532 8848 12572 8888 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 12532 8762 12572 8802 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 12532 8676 12572 8716 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 12532 8590 12572 8630 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 12532 8504 12572 8544 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 12532 8418 12572 8458 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 12532 8332 12572 8372 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 12451 9192 12491 9232 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 12451 9106 12491 9146 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 12451 9020 12491 9060 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 12451 8934 12491 8974 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 12451 8848 12491 8888 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 12451 8762 12491 8802 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 12451 8676 12491 8716 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 12451 8590 12491 8630 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 12451 8504 12491 8544 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 12451 8418 12491 8458 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 12451 8332 12491 8372 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 12370 9192 12410 9232 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 12370 9106 12410 9146 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 12370 9020 12410 9060 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 12370 8934 12410 8974 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 12370 8848 12410 8888 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 12370 8762 12410 8802 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 12370 8676 12410 8716 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 12370 8590 12410 8630 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 12370 8504 12410 8544 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 12370 8418 12410 8458 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 12370 8332 12410 8372 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 12289 9192 12329 9232 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 12289 9106 12329 9146 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 12289 9020 12329 9060 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 12289 8934 12329 8974 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 12289 8848 12329 8888 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 12289 8762 12329 8802 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 12289 8676 12329 8716 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 12289 8590 12329 8630 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 12289 8504 12329 8544 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 12289 8418 12329 8458 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 12289 8332 12329 8372 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 12208 9192 12248 9232 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 12208 9106 12248 9146 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 12208 9020 12248 9060 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 12208 8934 12248 8974 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 12208 8848 12248 8888 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 12208 8762 12248 8802 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 12208 8676 12248 8716 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 12208 8590 12248 8630 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 12208 8504 12248 8544 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 12208 8418 12248 8458 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 12208 8332 12248 8372 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 12127 9192 12167 9232 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 12127 9106 12167 9146 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 12127 9020 12167 9060 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 12127 8934 12167 8974 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 12127 8848 12167 8888 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 12127 8762 12167 8802 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 12127 8676 12167 8716 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 12127 8590 12167 8630 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 12127 8504 12167 8544 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 12127 8418 12167 8458 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 12127 8332 12167 8372 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 12046 9192 12086 9232 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 12046 9106 12086 9146 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 12046 9020 12086 9060 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 12046 8934 12086 8974 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 12046 8848 12086 8888 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 12046 8762 12086 8802 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 12046 8676 12086 8716 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 12046 8590 12086 8630 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 12046 8504 12086 8544 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 12046 8418 12086 8458 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 12046 8332 12086 8372 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 11965 9192 12005 9232 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 11965 9106 12005 9146 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 11965 9020 12005 9060 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 11965 8934 12005 8974 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 11965 8848 12005 8888 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 11965 8762 12005 8802 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 11965 8676 12005 8716 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 11965 8590 12005 8630 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 11965 8504 12005 8544 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 11965 8418 12005 8458 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 11965 8332 12005 8372 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 11884 9192 11924 9232 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 11884 9106 11924 9146 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 11884 9020 11924 9060 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 11884 8934 11924 8974 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 11884 8848 11924 8888 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 11884 8762 11924 8802 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 11884 8676 11924 8716 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 11884 8590 11924 8630 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 11884 8504 11924 8544 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 11884 8418 11924 8458 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 11884 8332 11924 8372 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 11803 9192 11843 9232 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 11803 9106 11843 9146 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 11803 9020 11843 9060 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 11803 8934 11843 8974 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 11803 8848 11843 8888 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 11803 8762 11843 8802 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 11803 8676 11843 8716 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 11803 8590 11843 8630 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 11803 8504 11843 8544 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 11803 8418 11843 8458 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 11803 8332 11843 8372 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 11722 9192 11762 9232 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 11722 9106 11762 9146 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 11722 9020 11762 9060 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 11722 8934 11762 8974 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 11722 8848 11762 8888 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 11722 8762 11762 8802 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 11722 8676 11762 8716 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 11722 8590 11762 8630 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 11722 8504 11762 8544 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 11722 8418 11762 8458 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 11722 8332 11762 8372 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 11641 9192 11681 9232 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 11641 9106 11681 9146 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 11641 9020 11681 9060 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 11641 8934 11681 8974 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 11641 8848 11681 8888 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 11641 8762 11681 8802 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 11641 8676 11681 8716 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 11641 8590 11681 8630 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 11641 8504 11681 8544 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 11641 8418 11681 8458 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 11641 8332 11681 8372 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 11560 9192 11600 9232 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 11560 9106 11600 9146 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 11560 9020 11600 9060 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 11560 8934 11600 8974 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 11560 8848 11600 8888 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 11560 8762 11600 8802 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 11560 8676 11600 8716 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 11560 8590 11600 8630 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 11560 8504 11600 8544 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 11560 8418 11600 8458 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 11560 8332 11600 8372 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 11479 9192 11519 9232 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 11479 9106 11519 9146 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 11479 9020 11519 9060 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 11479 8934 11519 8974 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 11479 8848 11519 8888 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 11479 8762 11519 8802 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 11479 8676 11519 8716 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 11479 8590 11519 8630 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 11479 8504 11519 8544 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 11479 8418 11519 8458 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 11479 8332 11519 8372 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 11398 9192 11438 9232 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 11398 9106 11438 9146 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 11398 9020 11438 9060 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 11398 8934 11438 8974 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 11398 8848 11438 8888 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 11398 8762 11438 8802 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 11398 8676 11438 8716 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 11398 8590 11438 8630 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 11398 8504 11438 8544 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 11398 8418 11438 8458 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 11398 8332 11438 8372 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 11317 9192 11357 9232 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 11317 9106 11357 9146 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 11317 9020 11357 9060 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 11317 8934 11357 8974 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 11317 8848 11357 8888 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 11317 8762 11357 8802 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 11317 8676 11357 8716 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 11317 8590 11357 8630 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 11317 8504 11357 8544 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 11317 8418 11357 8458 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 11317 8332 11357 8372 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 11236 9192 11276 9232 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 11236 9106 11276 9146 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 11236 9020 11276 9060 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 11236 8934 11276 8974 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 11236 8848 11276 8888 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 11236 8762 11276 8802 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 11236 8676 11276 8716 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 11236 8590 11276 8630 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 11236 8504 11276 8544 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 11236 8418 11276 8458 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 11236 8332 11276 8372 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 11155 9192 11195 9232 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 11155 9106 11195 9146 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 11155 9020 11195 9060 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 11155 8934 11195 8974 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 11155 8848 11195 8888 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 11155 8762 11195 8802 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 11155 8676 11195 8716 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 11155 8590 11195 8630 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 11155 8504 11195 8544 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 11155 8418 11195 8458 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 11155 8332 11195 8372 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 11074 9192 11114 9232 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 11074 9106 11114 9146 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 11074 9020 11114 9060 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 11074 8934 11114 8974 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 11074 8848 11114 8888 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 11074 8762 11114 8802 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 11074 8676 11114 8716 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 11074 8590 11114 8630 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 11074 8504 11114 8544 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 11074 8418 11114 8458 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 11074 8332 11114 8372 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 10993 9192 11033 9232 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 10993 9106 11033 9146 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 10993 9020 11033 9060 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 10993 8934 11033 8974 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 10993 8848 11033 8888 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 10993 8762 11033 8802 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 10993 8676 11033 8716 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 10993 8590 11033 8630 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 10993 8504 11033 8544 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 10993 8418 11033 8458 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 10993 8332 11033 8372 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 10912 9192 10952 9232 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 10912 9106 10952 9146 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 10912 9020 10952 9060 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 10912 8934 10952 8974 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 10912 8848 10952 8888 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 10912 8762 10952 8802 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 10912 8676 10952 8716 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 10912 8590 10952 8630 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 10912 8504 10952 8544 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 10912 8418 10952 8458 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 10912 8332 10952 8372 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 10831 9192 10871 9232 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 10831 9106 10871 9146 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 10831 9020 10871 9060 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 10831 8934 10871 8974 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 10831 8848 10871 8888 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 10831 8762 10871 8802 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 10831 8676 10871 8716 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 10831 8590 10871 8630 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 10831 8504 10871 8544 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 10831 8418 10871 8458 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 10831 8332 10871 8372 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 10750 9192 10790 9232 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 10750 9106 10790 9146 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 10750 9020 10790 9060 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 10750 8934 10790 8974 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 10750 8848 10790 8888 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 10750 8762 10790 8802 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 10750 8676 10790 8716 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 10750 8590 10790 8630 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 10750 8504 10790 8544 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 10750 8418 10790 8458 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 10750 8332 10790 8372 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 10669 9192 10709 9232 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 10669 9106 10709 9146 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 10669 9020 10709 9060 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 10669 8934 10709 8974 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 10669 8848 10709 8888 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 10669 8762 10709 8802 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 10669 8676 10709 8716 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 10669 8590 10709 8630 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 10669 8504 10709 8544 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 10669 8418 10709 8458 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 10669 8332 10709 8372 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 10588 9192 10628 9232 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 10588 9106 10628 9146 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 10588 9020 10628 9060 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 10588 8934 10628 8974 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 10588 8848 10628 8888 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 10588 8762 10628 8802 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 10588 8676 10628 8716 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 10588 8590 10628 8630 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 10588 8504 10628 8544 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 10588 8418 10628 8458 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 10588 8332 10628 8372 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 10506 9192 10546 9232 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 10506 9106 10546 9146 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 10506 9020 10546 9060 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 10506 8934 10546 8974 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 10506 8848 10546 8888 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 10506 8762 10546 8802 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 10506 8676 10546 8716 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 10506 8590 10546 8630 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 10506 8504 10546 8544 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 10506 8418 10546 8458 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 10506 8332 10546 8372 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 10424 9192 10464 9232 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 10424 9106 10464 9146 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 10424 9020 10464 9060 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 10424 8934 10464 8974 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 10424 8848 10464 8888 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 10424 8762 10464 8802 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 10424 8676 10464 8716 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 10424 8590 10464 8630 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 10424 8504 10464 8544 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 10424 8418 10464 8458 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 10424 8332 10464 8372 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 10342 9192 10382 9232 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 10342 9106 10382 9146 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 10342 9020 10382 9060 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 10342 8934 10382 8974 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 10342 8848 10382 8888 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 10342 8762 10382 8802 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 10342 8676 10382 8716 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 10342 8590 10382 8630 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 10342 8504 10382 8544 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 10342 8418 10382 8458 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 10342 8332 10382 8372 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 10260 9192 10300 9232 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 10260 9106 10300 9146 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 10260 9020 10300 9060 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 10260 8934 10300 8974 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 10260 8848 10300 8888 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 10260 8762 10300 8802 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 10260 8676 10300 8716 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 10260 8590 10300 8630 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 10260 8504 10300 8544 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 10260 8418 10300 8458 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 10260 8332 10300 8372 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 10178 9192 10218 9232 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 10178 9106 10218 9146 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 10178 9020 10218 9060 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 10178 8934 10218 8974 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 10178 8848 10218 8888 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 10178 8762 10218 8802 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 10178 8676 10218 8716 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 10178 8590 10218 8630 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 10178 8504 10218 8544 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 10178 8418 10218 8458 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 10178 8332 10218 8372 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 10096 9192 10136 9232 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 10096 9106 10136 9146 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 10096 9020 10136 9060 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 10096 8934 10136 8974 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 10096 8848 10136 8888 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 10096 8762 10136 8802 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 10096 8676 10136 8716 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 10096 8590 10136 8630 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 10096 8504 10136 8544 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 10096 8418 10136 8458 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 10096 8332 10136 8372 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 4809 9180 4873 9244 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 4809 9180 4873 9244 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 4809 9094 4873 9158 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 4809 9094 4873 9158 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 4809 9008 4873 9072 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 4809 9008 4873 9072 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 4809 8922 4873 8986 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 4809 8922 4873 8986 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 4809 8836 4873 8900 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 4809 8836 4873 8900 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 4809 8750 4873 8814 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 4809 8750 4873 8814 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 4809 8664 4873 8728 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 4809 8664 4873 8728 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 4809 8578 4873 8642 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 4809 8578 4873 8642 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 4809 8492 4873 8556 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 4809 8492 4873 8556 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 4809 8406 4873 8470 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 4809 8406 4873 8470 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 4809 8320 4873 8384 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 4809 8320 4873 8384 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 4729 9180 4793 9244 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 4729 9180 4793 9244 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 4729 9094 4793 9158 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 4729 9094 4793 9158 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 4729 9008 4793 9072 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 4729 9008 4793 9072 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 4729 8922 4793 8986 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 4729 8922 4793 8986 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 4729 8836 4793 8900 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 4729 8836 4793 8900 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 4729 8750 4793 8814 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 4729 8750 4793 8814 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 4729 8664 4793 8728 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 4729 8664 4793 8728 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 4729 8578 4793 8642 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 4729 8578 4793 8642 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 4729 8492 4793 8556 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 4729 8492 4793 8556 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 4729 8406 4793 8470 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 4729 8406 4793 8470 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 4729 8320 4793 8384 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 4729 8320 4793 8384 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 4649 9180 4713 9244 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 4649 9180 4713 9244 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 4649 9094 4713 9158 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 4649 9094 4713 9158 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 4649 9008 4713 9072 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 4649 9008 4713 9072 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 4649 8922 4713 8986 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 4649 8922 4713 8986 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 4649 8836 4713 8900 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 4649 8836 4713 8900 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 4649 8750 4713 8814 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 4649 8750 4713 8814 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 4649 8664 4713 8728 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 4649 8664 4713 8728 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 4649 8578 4713 8642 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 4649 8578 4713 8642 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 4649 8492 4713 8556 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 4649 8492 4713 8556 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 4649 8406 4713 8470 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 4649 8406 4713 8470 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 4649 8320 4713 8384 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 4649 8320 4713 8384 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 4569 9180 4633 9244 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 4569 9180 4633 9244 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 4569 9094 4633 9158 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 4569 9094 4633 9158 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 4569 9008 4633 9072 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 4569 9008 4633 9072 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 4569 8922 4633 8986 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 4569 8922 4633 8986 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 4569 8836 4633 8900 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 4569 8836 4633 8900 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 4569 8750 4633 8814 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 4569 8750 4633 8814 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 4569 8664 4633 8728 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 4569 8664 4633 8728 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 4569 8578 4633 8642 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 4569 8578 4633 8642 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 4569 8492 4633 8556 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 4569 8492 4633 8556 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 4569 8406 4633 8470 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 4569 8406 4633 8470 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 4569 8320 4633 8384 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 4569 8320 4633 8384 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 4489 9180 4553 9244 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 4489 9180 4553 9244 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 4489 9094 4553 9158 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 4489 9094 4553 9158 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 4489 9008 4553 9072 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 4489 9008 4553 9072 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 4489 8922 4553 8986 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 4489 8922 4553 8986 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 4489 8836 4553 8900 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 4489 8836 4553 8900 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 4489 8750 4553 8814 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 4489 8750 4553 8814 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 4489 8664 4553 8728 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 4489 8664 4553 8728 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 4489 8578 4553 8642 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 4489 8578 4553 8642 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 4489 8492 4553 8556 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 4489 8492 4553 8556 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 4489 8406 4553 8470 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 4489 8406 4553 8470 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 4489 8320 4553 8384 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 4489 8320 4553 8384 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 4409 9180 4473 9244 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 4409 9180 4473 9244 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 4409 9094 4473 9158 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 4409 9094 4473 9158 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 4409 9008 4473 9072 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 4409 9008 4473 9072 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 4409 8922 4473 8986 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 4409 8922 4473 8986 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 4409 8836 4473 8900 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 4409 8836 4473 8900 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 4409 8750 4473 8814 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 4409 8750 4473 8814 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 4409 8664 4473 8728 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 4409 8664 4473 8728 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 4409 8578 4473 8642 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 4409 8578 4473 8642 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 4409 8492 4473 8556 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 4409 8492 4473 8556 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 4409 8406 4473 8470 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 4409 8406 4473 8470 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 4409 8320 4473 8384 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 4409 8320 4473 8384 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 4329 9180 4393 9244 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 4329 9180 4393 9244 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 4329 9094 4393 9158 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 4329 9094 4393 9158 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 4329 9008 4393 9072 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 4329 9008 4393 9072 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 4329 8922 4393 8986 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 4329 8922 4393 8986 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 4329 8836 4393 8900 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 4329 8836 4393 8900 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 4329 8750 4393 8814 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 4329 8750 4393 8814 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 4329 8664 4393 8728 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 4329 8664 4393 8728 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 4329 8578 4393 8642 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 4329 8578 4393 8642 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 4329 8492 4393 8556 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 4329 8492 4393 8556 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 4329 8406 4393 8470 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 4329 8406 4393 8470 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 4329 8320 4393 8384 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 4329 8320 4393 8384 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 4249 9180 4313 9244 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 4249 9180 4313 9244 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 4249 9094 4313 9158 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 4249 9094 4313 9158 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 4249 9008 4313 9072 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 4249 9008 4313 9072 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 4249 8922 4313 8986 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 4249 8922 4313 8986 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 4249 8836 4313 8900 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 4249 8836 4313 8900 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 4249 8750 4313 8814 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 4249 8750 4313 8814 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 4249 8664 4313 8728 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 4249 8664 4313 8728 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 4249 8578 4313 8642 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 4249 8578 4313 8642 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 4249 8492 4313 8556 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 4249 8492 4313 8556 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 4249 8406 4313 8470 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 4249 8406 4313 8470 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 4249 8320 4313 8384 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 4249 8320 4313 8384 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 4169 9180 4233 9244 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 4169 9180 4233 9244 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 4169 9094 4233 9158 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 4169 9094 4233 9158 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 4169 9008 4233 9072 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 4169 9008 4233 9072 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 4169 8922 4233 8986 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 4169 8922 4233 8986 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 4169 8836 4233 8900 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 4169 8836 4233 8900 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 4169 8750 4233 8814 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 4169 8750 4233 8814 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 4169 8664 4233 8728 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 4169 8664 4233 8728 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 4169 8578 4233 8642 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 4169 8578 4233 8642 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 4169 8492 4233 8556 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 4169 8492 4233 8556 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 4169 8406 4233 8470 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 4169 8406 4233 8470 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 4169 8320 4233 8384 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 4169 8320 4233 8384 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 4088 9180 4152 9244 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 4088 9180 4152 9244 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 4088 9094 4152 9158 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 4088 9094 4152 9158 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 4088 9008 4152 9072 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 4088 9008 4152 9072 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 4088 8922 4152 8986 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 4088 8922 4152 8986 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 4088 8836 4152 8900 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 4088 8836 4152 8900 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 4088 8750 4152 8814 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 4088 8750 4152 8814 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 4088 8664 4152 8728 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 4088 8664 4152 8728 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 4088 8578 4152 8642 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 4088 8578 4152 8642 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 4088 8492 4152 8556 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 4088 8492 4152 8556 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 4088 8406 4152 8470 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 4088 8406 4152 8470 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 4088 8320 4152 8384 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 4088 8320 4152 8384 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 4007 9180 4071 9244 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 4007 9180 4071 9244 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 4007 9094 4071 9158 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 4007 9094 4071 9158 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 4007 9008 4071 9072 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 4007 9008 4071 9072 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 4007 8922 4071 8986 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 4007 8922 4071 8986 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 4007 8836 4071 8900 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 4007 8836 4071 8900 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 4007 8750 4071 8814 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 4007 8750 4071 8814 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 4007 8664 4071 8728 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 4007 8664 4071 8728 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 4007 8578 4071 8642 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 4007 8578 4071 8642 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 4007 8492 4071 8556 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 4007 8492 4071 8556 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 4007 8406 4071 8470 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 4007 8406 4071 8470 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 4007 8320 4071 8384 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 4007 8320 4071 8384 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 3926 9180 3990 9244 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 3926 9180 3990 9244 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 3926 9094 3990 9158 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 3926 9094 3990 9158 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 3926 9008 3990 9072 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 3926 9008 3990 9072 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 3926 8922 3990 8986 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 3926 8922 3990 8986 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 3926 8836 3990 8900 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 3926 8836 3990 8900 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 3926 8750 3990 8814 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 3926 8750 3990 8814 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 3926 8664 3990 8728 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 3926 8664 3990 8728 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 3926 8578 3990 8642 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 3926 8578 3990 8642 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 3926 8492 3990 8556 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 3926 8492 3990 8556 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 3926 8406 3990 8470 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 3926 8406 3990 8470 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 3926 8320 3990 8384 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 3926 8320 3990 8384 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 3845 9180 3909 9244 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 3845 9180 3909 9244 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 3845 9094 3909 9158 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 3845 9094 3909 9158 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 3845 9008 3909 9072 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 3845 9008 3909 9072 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 3845 8922 3909 8986 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 3845 8922 3909 8986 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 3845 8836 3909 8900 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 3845 8836 3909 8900 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 3845 8750 3909 8814 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 3845 8750 3909 8814 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 3845 8664 3909 8728 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 3845 8664 3909 8728 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 3845 8578 3909 8642 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 3845 8578 3909 8642 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 3845 8492 3909 8556 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 3845 8492 3909 8556 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 3845 8406 3909 8470 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 3845 8406 3909 8470 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 3845 8320 3909 8384 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 3845 8320 3909 8384 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 3764 9180 3828 9244 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 3764 9180 3828 9244 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 3764 9094 3828 9158 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 3764 9094 3828 9158 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 3764 9008 3828 9072 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 3764 9008 3828 9072 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 3764 8922 3828 8986 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 3764 8922 3828 8986 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 3764 8836 3828 8900 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 3764 8836 3828 8900 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 3764 8750 3828 8814 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 3764 8750 3828 8814 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 3764 8664 3828 8728 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 3764 8664 3828 8728 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 3764 8578 3828 8642 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 3764 8578 3828 8642 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 3764 8492 3828 8556 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 3764 8492 3828 8556 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 3764 8406 3828 8470 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 3764 8406 3828 8470 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 3764 8320 3828 8384 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 3764 8320 3828 8384 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 3683 9180 3747 9244 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 3683 9180 3747 9244 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 3683 9094 3747 9158 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 3683 9094 3747 9158 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 3683 9008 3747 9072 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 3683 9008 3747 9072 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 3683 8922 3747 8986 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 3683 8922 3747 8986 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 3683 8836 3747 8900 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 3683 8836 3747 8900 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 3683 8750 3747 8814 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 3683 8750 3747 8814 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 3683 8664 3747 8728 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 3683 8664 3747 8728 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 3683 8578 3747 8642 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 3683 8578 3747 8642 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 3683 8492 3747 8556 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 3683 8492 3747 8556 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 3683 8406 3747 8470 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 3683 8406 3747 8470 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 3683 8320 3747 8384 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 3683 8320 3747 8384 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 3602 9180 3666 9244 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 3602 9180 3666 9244 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 3602 9094 3666 9158 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 3602 9094 3666 9158 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 3602 9008 3666 9072 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 3602 9008 3666 9072 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 3602 8922 3666 8986 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 3602 8922 3666 8986 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 3602 8836 3666 8900 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 3602 8836 3666 8900 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 3602 8750 3666 8814 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 3602 8750 3666 8814 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 3602 8664 3666 8728 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 3602 8664 3666 8728 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 3602 8578 3666 8642 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 3602 8578 3666 8642 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 3602 8492 3666 8556 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 3602 8492 3666 8556 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 3602 8406 3666 8470 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 3602 8406 3666 8470 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 3602 8320 3666 8384 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 3602 8320 3666 8384 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 3521 9180 3585 9244 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 3521 9180 3585 9244 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 3521 9094 3585 9158 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 3521 9094 3585 9158 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 3521 9008 3585 9072 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 3521 9008 3585 9072 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 3521 8922 3585 8986 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 3521 8922 3585 8986 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 3521 8836 3585 8900 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 3521 8836 3585 8900 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 3521 8750 3585 8814 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 3521 8750 3585 8814 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 3521 8664 3585 8728 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 3521 8664 3585 8728 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 3521 8578 3585 8642 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 3521 8578 3585 8642 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 3521 8492 3585 8556 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 3521 8492 3585 8556 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 3521 8406 3585 8470 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 3521 8406 3585 8470 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 3521 8320 3585 8384 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 3521 8320 3585 8384 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 3440 9180 3504 9244 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 3440 9180 3504 9244 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 3440 9094 3504 9158 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 3440 9094 3504 9158 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 3440 9008 3504 9072 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 3440 9008 3504 9072 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 3440 8922 3504 8986 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 3440 8922 3504 8986 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 3440 8836 3504 8900 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 3440 8836 3504 8900 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 3440 8750 3504 8814 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 3440 8750 3504 8814 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 3440 8664 3504 8728 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 3440 8664 3504 8728 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 3440 8578 3504 8642 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 3440 8578 3504 8642 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 3440 8492 3504 8556 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 3440 8492 3504 8556 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 3440 8406 3504 8470 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 3440 8406 3504 8470 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 3440 8320 3504 8384 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 3440 8320 3504 8384 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 3359 9180 3423 9244 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 3359 9180 3423 9244 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 3359 9094 3423 9158 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 3359 9094 3423 9158 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 3359 9008 3423 9072 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 3359 9008 3423 9072 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 3359 8922 3423 8986 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 3359 8922 3423 8986 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 3359 8836 3423 8900 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 3359 8836 3423 8900 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 3359 8750 3423 8814 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 3359 8750 3423 8814 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 3359 8664 3423 8728 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 3359 8664 3423 8728 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 3359 8578 3423 8642 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 3359 8578 3423 8642 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 3359 8492 3423 8556 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 3359 8492 3423 8556 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 3359 8406 3423 8470 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 3359 8406 3423 8470 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 3359 8320 3423 8384 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 3359 8320 3423 8384 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 3278 9180 3342 9244 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 3278 9180 3342 9244 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 3278 9094 3342 9158 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 3278 9094 3342 9158 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 3278 9008 3342 9072 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 3278 9008 3342 9072 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 3278 8922 3342 8986 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 3278 8922 3342 8986 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 3278 8836 3342 8900 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 3278 8836 3342 8900 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 3278 8750 3342 8814 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 3278 8750 3342 8814 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 3278 8664 3342 8728 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 3278 8664 3342 8728 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 3278 8578 3342 8642 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 3278 8578 3342 8642 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 3278 8492 3342 8556 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 3278 8492 3342 8556 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 3278 8406 3342 8470 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 3278 8406 3342 8470 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 3278 8320 3342 8384 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 3278 8320 3342 8384 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 3197 9180 3261 9244 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 3197 9180 3261 9244 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 3197 9094 3261 9158 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 3197 9094 3261 9158 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 3197 9008 3261 9072 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 3197 9008 3261 9072 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 3197 8922 3261 8986 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 3197 8922 3261 8986 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 3197 8836 3261 8900 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 3197 8836 3261 8900 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 3197 8750 3261 8814 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 3197 8750 3261 8814 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 3197 8664 3261 8728 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 3197 8664 3261 8728 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 3197 8578 3261 8642 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 3197 8578 3261 8642 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 3197 8492 3261 8556 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 3197 8492 3261 8556 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 3197 8406 3261 8470 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 3197 8406 3261 8470 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 3197 8320 3261 8384 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 3197 8320 3261 8384 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 3116 9180 3180 9244 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 3116 9180 3180 9244 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 3116 9094 3180 9158 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 3116 9094 3180 9158 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 3116 9008 3180 9072 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 3116 9008 3180 9072 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 3116 8922 3180 8986 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 3116 8922 3180 8986 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 3116 8836 3180 8900 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 3116 8836 3180 8900 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 3116 8750 3180 8814 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 3116 8750 3180 8814 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 3116 8664 3180 8728 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 3116 8664 3180 8728 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 3116 8578 3180 8642 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 3116 8578 3180 8642 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 3116 8492 3180 8556 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 3116 8492 3180 8556 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 3116 8406 3180 8470 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 3116 8406 3180 8470 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 3116 8320 3180 8384 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 3116 8320 3180 8384 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 3035 9180 3099 9244 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 3035 9180 3099 9244 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 3035 9094 3099 9158 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 3035 9094 3099 9158 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 3035 9008 3099 9072 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 3035 9008 3099 9072 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 3035 8922 3099 8986 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 3035 8922 3099 8986 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 3035 8836 3099 8900 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 3035 8836 3099 8900 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 3035 8750 3099 8814 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 3035 8750 3099 8814 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 3035 8664 3099 8728 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 3035 8664 3099 8728 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 3035 8578 3099 8642 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 3035 8578 3099 8642 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 3035 8492 3099 8556 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 3035 8492 3099 8556 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 3035 8406 3099 8470 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 3035 8406 3099 8470 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 3035 8320 3099 8384 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 3035 8320 3099 8384 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2954 9180 3018 9244 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2954 9180 3018 9244 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2954 9094 3018 9158 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2954 9094 3018 9158 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2954 9008 3018 9072 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2954 9008 3018 9072 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2954 8922 3018 8986 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2954 8922 3018 8986 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2954 8836 3018 8900 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2954 8836 3018 8900 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2954 8750 3018 8814 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2954 8750 3018 8814 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2954 8664 3018 8728 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2954 8664 3018 8728 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2954 8578 3018 8642 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2954 8578 3018 8642 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2954 8492 3018 8556 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2954 8492 3018 8556 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2954 8406 3018 8470 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2954 8406 3018 8470 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2954 8320 3018 8384 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2954 8320 3018 8384 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2873 9180 2937 9244 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2873 9180 2937 9244 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2873 9094 2937 9158 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2873 9094 2937 9158 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2873 9008 2937 9072 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2873 9008 2937 9072 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2873 8922 2937 8986 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2873 8922 2937 8986 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2873 8836 2937 8900 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2873 8836 2937 8900 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2873 8750 2937 8814 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2873 8750 2937 8814 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2873 8664 2937 8728 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2873 8664 2937 8728 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2873 8578 2937 8642 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2873 8578 2937 8642 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2873 8492 2937 8556 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2873 8492 2937 8556 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2873 8406 2937 8470 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2873 8406 2937 8470 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2873 8320 2937 8384 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2873 8320 2937 8384 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2792 9180 2856 9244 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2792 9180 2856 9244 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2792 9094 2856 9158 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2792 9094 2856 9158 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2792 9008 2856 9072 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2792 9008 2856 9072 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2792 8922 2856 8986 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2792 8922 2856 8986 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2792 8836 2856 8900 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2792 8836 2856 8900 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2792 8750 2856 8814 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2792 8750 2856 8814 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2792 8664 2856 8728 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2792 8664 2856 8728 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2792 8578 2856 8642 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2792 8578 2856 8642 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2792 8492 2856 8556 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2792 8492 2856 8556 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2792 8406 2856 8470 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2792 8406 2856 8470 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2792 8320 2856 8384 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2792 8320 2856 8384 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2711 9180 2775 9244 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2711 9180 2775 9244 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2711 9094 2775 9158 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2711 9094 2775 9158 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2711 9008 2775 9072 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2711 9008 2775 9072 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2711 8922 2775 8986 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2711 8922 2775 8986 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2711 8836 2775 8900 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2711 8836 2775 8900 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2711 8750 2775 8814 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2711 8750 2775 8814 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2711 8664 2775 8728 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2711 8664 2775 8728 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2711 8578 2775 8642 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2711 8578 2775 8642 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2711 8492 2775 8556 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2711 8492 2775 8556 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2711 8406 2775 8470 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2711 8406 2775 8470 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2711 8320 2775 8384 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2711 8320 2775 8384 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2630 9180 2694 9244 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2630 9180 2694 9244 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2630 9094 2694 9158 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2630 9094 2694 9158 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2630 9008 2694 9072 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2630 9008 2694 9072 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2630 8922 2694 8986 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2630 8922 2694 8986 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2630 8836 2694 8900 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2630 8836 2694 8900 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2630 8750 2694 8814 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2630 8750 2694 8814 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2630 8664 2694 8728 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2630 8664 2694 8728 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2630 8578 2694 8642 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2630 8578 2694 8642 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2630 8492 2694 8556 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2630 8492 2694 8556 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2630 8406 2694 8470 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2630 8406 2694 8470 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2630 8320 2694 8384 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2630 8320 2694 8384 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2549 9180 2613 9244 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2549 9180 2613 9244 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2549 9094 2613 9158 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2549 9094 2613 9158 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2549 9008 2613 9072 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2549 9008 2613 9072 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2549 8922 2613 8986 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2549 8922 2613 8986 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2549 8836 2613 8900 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2549 8836 2613 8900 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2549 8750 2613 8814 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2549 8750 2613 8814 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2549 8664 2613 8728 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2549 8664 2613 8728 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2549 8578 2613 8642 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2549 8578 2613 8642 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2549 8492 2613 8556 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2549 8492 2613 8556 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2549 8406 2613 8470 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2549 8406 2613 8470 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2549 8320 2613 8384 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2549 8320 2613 8384 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2468 9180 2532 9244 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2468 9180 2532 9244 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2468 9094 2532 9158 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2468 9094 2532 9158 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2468 9008 2532 9072 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2468 9008 2532 9072 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2468 8922 2532 8986 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2468 8922 2532 8986 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2468 8836 2532 8900 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2468 8836 2532 8900 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2468 8750 2532 8814 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2468 8750 2532 8814 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2468 8664 2532 8728 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2468 8664 2532 8728 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2468 8578 2532 8642 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2468 8578 2532 8642 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2468 8492 2532 8556 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2468 8492 2532 8556 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2468 8406 2532 8470 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2468 8406 2532 8470 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2468 8320 2532 8384 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2468 8320 2532 8384 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2387 9180 2451 9244 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2387 9180 2451 9244 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2387 9094 2451 9158 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2387 9094 2451 9158 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2387 9008 2451 9072 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2387 9008 2451 9072 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2387 8922 2451 8986 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2387 8922 2451 8986 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2387 8836 2451 8900 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2387 8836 2451 8900 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2387 8750 2451 8814 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2387 8750 2451 8814 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2387 8664 2451 8728 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2387 8664 2451 8728 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2387 8578 2451 8642 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2387 8578 2451 8642 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2387 8492 2451 8556 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2387 8492 2451 8556 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2387 8406 2451 8470 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2387 8406 2451 8470 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2387 8320 2451 8384 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2387 8320 2451 8384 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2306 9180 2370 9244 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2306 9180 2370 9244 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2306 9094 2370 9158 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2306 9094 2370 9158 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2306 9008 2370 9072 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2306 9008 2370 9072 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2306 8922 2370 8986 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2306 8922 2370 8986 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2306 8836 2370 8900 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2306 8836 2370 8900 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2306 8750 2370 8814 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2306 8750 2370 8814 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2306 8664 2370 8728 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2306 8664 2370 8728 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2306 8578 2370 8642 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2306 8578 2370 8642 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2306 8492 2370 8556 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2306 8492 2370 8556 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2306 8406 2370 8470 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2306 8406 2370 8470 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2306 8320 2370 8384 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2306 8320 2370 8384 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2225 9180 2289 9244 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2225 9180 2289 9244 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2225 9094 2289 9158 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2225 9094 2289 9158 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2225 9008 2289 9072 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2225 9008 2289 9072 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2225 8922 2289 8986 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2225 8922 2289 8986 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2225 8836 2289 8900 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2225 8836 2289 8900 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2225 8750 2289 8814 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2225 8750 2289 8814 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2225 8664 2289 8728 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2225 8664 2289 8728 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2225 8578 2289 8642 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2225 8578 2289 8642 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2225 8492 2289 8556 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2225 8492 2289 8556 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2225 8406 2289 8470 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2225 8406 2289 8470 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2225 8320 2289 8384 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2225 8320 2289 8384 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2144 9180 2208 9244 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2144 9180 2208 9244 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2144 9094 2208 9158 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2144 9094 2208 9158 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2144 9008 2208 9072 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2144 9008 2208 9072 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2144 8922 2208 8986 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2144 8922 2208 8986 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2144 8836 2208 8900 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2144 8836 2208 8900 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2144 8750 2208 8814 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2144 8750 2208 8814 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2144 8664 2208 8728 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2144 8664 2208 8728 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2144 8578 2208 8642 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2144 8578 2208 8642 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2144 8492 2208 8556 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2144 8492 2208 8556 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2144 8406 2208 8470 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2144 8406 2208 8470 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2144 8320 2208 8384 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2144 8320 2208 8384 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2063 9180 2127 9244 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2063 9180 2127 9244 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2063 9094 2127 9158 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2063 9094 2127 9158 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2063 9008 2127 9072 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2063 9008 2127 9072 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2063 8922 2127 8986 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2063 8922 2127 8986 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2063 8836 2127 8900 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2063 8836 2127 8900 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2063 8750 2127 8814 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2063 8750 2127 8814 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2063 8664 2127 8728 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2063 8664 2127 8728 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2063 8578 2127 8642 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2063 8578 2127 8642 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2063 8492 2127 8556 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2063 8492 2127 8556 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2063 8406 2127 8470 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2063 8406 2127 8470 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2063 8320 2127 8384 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2063 8320 2127 8384 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1982 9180 2046 9244 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1982 9180 2046 9244 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1982 9094 2046 9158 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1982 9094 2046 9158 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1982 9008 2046 9072 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1982 9008 2046 9072 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1982 8922 2046 8986 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1982 8922 2046 8986 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1982 8836 2046 8900 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1982 8836 2046 8900 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1982 8750 2046 8814 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1982 8750 2046 8814 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1982 8664 2046 8728 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1982 8664 2046 8728 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1982 8578 2046 8642 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1982 8578 2046 8642 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1982 8492 2046 8556 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1982 8492 2046 8556 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1982 8406 2046 8470 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1982 8406 2046 8470 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1982 8320 2046 8384 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1982 8320 2046 8384 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1901 9180 1965 9244 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1901 9180 1965 9244 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1901 9094 1965 9158 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1901 9094 1965 9158 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1901 9008 1965 9072 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1901 9008 1965 9072 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1901 8922 1965 8986 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1901 8922 1965 8986 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1901 8836 1965 8900 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1901 8836 1965 8900 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1901 8750 1965 8814 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1901 8750 1965 8814 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1901 8664 1965 8728 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1901 8664 1965 8728 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1901 8578 1965 8642 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1901 8578 1965 8642 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1901 8492 1965 8556 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1901 8492 1965 8556 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1901 8406 1965 8470 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1901 8406 1965 8470 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1901 8320 1965 8384 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1901 8320 1965 8384 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1820 9180 1884 9244 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1820 9180 1884 9244 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1820 9094 1884 9158 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1820 9094 1884 9158 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1820 9008 1884 9072 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1820 9008 1884 9072 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1820 8922 1884 8986 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1820 8922 1884 8986 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1820 8836 1884 8900 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1820 8836 1884 8900 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1820 8750 1884 8814 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1820 8750 1884 8814 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1820 8664 1884 8728 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1820 8664 1884 8728 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1820 8578 1884 8642 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1820 8578 1884 8642 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1820 8492 1884 8556 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1820 8492 1884 8556 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1820 8406 1884 8470 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1820 8406 1884 8470 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1820 8320 1884 8384 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1820 8320 1884 8384 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1739 9180 1803 9244 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1739 9180 1803 9244 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1739 9094 1803 9158 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1739 9094 1803 9158 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1739 9008 1803 9072 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1739 9008 1803 9072 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1739 8922 1803 8986 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1739 8922 1803 8986 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1739 8836 1803 8900 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1739 8836 1803 8900 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1739 8750 1803 8814 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1739 8750 1803 8814 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1739 8664 1803 8728 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1739 8664 1803 8728 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1739 8578 1803 8642 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1739 8578 1803 8642 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1739 8492 1803 8556 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1739 8492 1803 8556 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1739 8406 1803 8470 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1739 8406 1803 8470 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1739 8320 1803 8384 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1739 8320 1803 8384 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1658 9180 1722 9244 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1658 9180 1722 9244 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1658 9094 1722 9158 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1658 9094 1722 9158 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1658 9008 1722 9072 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1658 9008 1722 9072 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1658 8922 1722 8986 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1658 8922 1722 8986 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1658 8836 1722 8900 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1658 8836 1722 8900 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1658 8750 1722 8814 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1658 8750 1722 8814 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1658 8664 1722 8728 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1658 8664 1722 8728 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1658 8578 1722 8642 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1658 8578 1722 8642 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1658 8492 1722 8556 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1658 8492 1722 8556 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1658 8406 1722 8470 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1658 8406 1722 8470 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1658 8320 1722 8384 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1658 8320 1722 8384 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1577 9180 1641 9244 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1577 9180 1641 9244 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1577 9094 1641 9158 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1577 9094 1641 9158 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1577 9008 1641 9072 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1577 9008 1641 9072 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1577 8922 1641 8986 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1577 8922 1641 8986 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1577 8836 1641 8900 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1577 8836 1641 8900 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1577 8750 1641 8814 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1577 8750 1641 8814 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1577 8664 1641 8728 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1577 8664 1641 8728 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1577 8578 1641 8642 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1577 8578 1641 8642 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1577 8492 1641 8556 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1577 8492 1641 8556 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1577 8406 1641 8470 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1577 8406 1641 8470 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1577 8320 1641 8384 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1577 8320 1641 8384 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1496 9180 1560 9244 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1496 9180 1560 9244 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1496 9094 1560 9158 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1496 9094 1560 9158 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1496 9008 1560 9072 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1496 9008 1560 9072 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1496 8922 1560 8986 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1496 8922 1560 8986 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1496 8836 1560 8900 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1496 8836 1560 8900 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1496 8750 1560 8814 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1496 8750 1560 8814 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1496 8664 1560 8728 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1496 8664 1560 8728 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1496 8578 1560 8642 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1496 8578 1560 8642 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1496 8492 1560 8556 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1496 8492 1560 8556 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1496 8406 1560 8470 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1496 8406 1560 8470 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1496 8320 1560 8384 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1496 8320 1560 8384 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1415 9180 1479 9244 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1415 9180 1479 9244 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1415 9094 1479 9158 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1415 9094 1479 9158 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1415 9008 1479 9072 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1415 9008 1479 9072 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1415 8922 1479 8986 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1415 8922 1479 8986 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1415 8836 1479 8900 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1415 8836 1479 8900 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1415 8750 1479 8814 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1415 8750 1479 8814 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1415 8664 1479 8728 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1415 8664 1479 8728 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1415 8578 1479 8642 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1415 8578 1479 8642 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1415 8492 1479 8556 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1415 8492 1479 8556 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1415 8406 1479 8470 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1415 8406 1479 8470 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1415 8320 1479 8384 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1415 8320 1479 8384 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1334 9180 1398 9244 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1334 9180 1398 9244 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1334 9094 1398 9158 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1334 9094 1398 9158 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1334 9008 1398 9072 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1334 9008 1398 9072 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1334 8922 1398 8986 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1334 8922 1398 8986 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1334 8836 1398 8900 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1334 8836 1398 8900 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1334 8750 1398 8814 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1334 8750 1398 8814 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1334 8664 1398 8728 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1334 8664 1398 8728 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1334 8578 1398 8642 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1334 8578 1398 8642 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1334 8492 1398 8556 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1334 8492 1398 8556 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1334 8406 1398 8470 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1334 8406 1398 8470 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1334 8320 1398 8384 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1334 8320 1398 8384 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1253 9180 1317 9244 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1253 9180 1317 9244 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1253 9094 1317 9158 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1253 9094 1317 9158 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1253 9008 1317 9072 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1253 9008 1317 9072 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1253 8922 1317 8986 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1253 8922 1317 8986 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1253 8836 1317 8900 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1253 8836 1317 8900 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1253 8750 1317 8814 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1253 8750 1317 8814 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1253 8664 1317 8728 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1253 8664 1317 8728 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1253 8578 1317 8642 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1253 8578 1317 8642 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1253 8492 1317 8556 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1253 8492 1317 8556 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1253 8406 1317 8470 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1253 8406 1317 8470 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1253 8320 1317 8384 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1253 8320 1317 8384 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1172 9180 1236 9244 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1172 9180 1236 9244 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1172 9094 1236 9158 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1172 9094 1236 9158 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1172 9008 1236 9072 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1172 9008 1236 9072 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1172 8922 1236 8986 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1172 8922 1236 8986 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1172 8836 1236 8900 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1172 8836 1236 8900 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1172 8750 1236 8814 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1172 8750 1236 8814 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1172 8664 1236 8728 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1172 8664 1236 8728 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1172 8578 1236 8642 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1172 8578 1236 8642 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1172 8492 1236 8556 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1172 8492 1236 8556 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1172 8406 1236 8470 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1172 8406 1236 8470 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1172 8320 1236 8384 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1172 8320 1236 8384 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1091 9180 1155 9244 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1091 9180 1155 9244 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1091 9094 1155 9158 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1091 9094 1155 9158 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1091 9008 1155 9072 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1091 9008 1155 9072 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1091 8922 1155 8986 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1091 8922 1155 8986 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1091 8836 1155 8900 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1091 8836 1155 8900 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1091 8750 1155 8814 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1091 8750 1155 8814 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1091 8664 1155 8728 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1091 8664 1155 8728 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1091 8578 1155 8642 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1091 8578 1155 8642 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1091 8492 1155 8556 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1091 8492 1155 8556 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1091 8406 1155 8470 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1091 8406 1155 8470 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1091 8320 1155 8384 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1091 8320 1155 8384 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1010 9180 1074 9244 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1010 9180 1074 9244 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1010 9094 1074 9158 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1010 9094 1074 9158 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1010 9008 1074 9072 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1010 9008 1074 9072 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1010 8922 1074 8986 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1010 8922 1074 8986 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1010 8836 1074 8900 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1010 8836 1074 8900 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1010 8750 1074 8814 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1010 8750 1074 8814 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1010 8664 1074 8728 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1010 8664 1074 8728 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1010 8578 1074 8642 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1010 8578 1074 8642 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1010 8492 1074 8556 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1010 8492 1074 8556 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1010 8406 1074 8470 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1010 8406 1074 8470 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1010 8320 1074 8384 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1010 8320 1074 8384 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 929 9180 993 9244 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 929 9180 993 9244 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 929 9094 993 9158 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 929 9094 993 9158 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 929 9008 993 9072 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 929 9008 993 9072 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 929 8922 993 8986 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 929 8922 993 8986 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 929 8836 993 8900 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 929 8836 993 8900 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 929 8750 993 8814 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 929 8750 993 8814 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 929 8664 993 8728 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 929 8664 993 8728 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 929 8578 993 8642 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 929 8578 993 8642 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 929 8492 993 8556 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 929 8492 993 8556 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 929 8406 993 8470 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 929 8406 993 8470 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 929 8320 993 8384 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 929 8320 993 8384 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 848 9180 912 9244 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 848 9180 912 9244 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 848 9094 912 9158 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 848 9094 912 9158 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 848 9008 912 9072 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 848 9008 912 9072 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 848 8922 912 8986 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 848 8922 912 8986 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 848 8836 912 8900 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 848 8836 912 8900 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 848 8750 912 8814 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 848 8750 912 8814 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 848 8664 912 8728 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 848 8664 912 8728 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 848 8578 912 8642 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 848 8578 912 8642 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 848 8492 912 8556 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 848 8492 912 8556 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 848 8406 912 8470 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 848 8406 912 8470 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 848 8320 912 8384 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 848 8320 912 8384 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 767 9180 831 9244 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 767 9180 831 9244 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 767 9094 831 9158 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 767 9094 831 9158 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 767 9008 831 9072 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 767 9008 831 9072 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 767 8922 831 8986 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 767 8922 831 8986 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 767 8836 831 8900 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 767 8836 831 8900 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 767 8750 831 8814 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 767 8750 831 8814 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 767 8664 831 8728 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 767 8664 831 8728 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 767 8578 831 8642 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 767 8578 831 8642 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 767 8492 831 8556 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 767 8492 831 8556 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 767 8406 831 8470 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 767 8406 831 8470 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 767 8320 831 8384 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 767 8320 831 8384 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 686 9180 750 9244 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 686 9180 750 9244 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 686 9094 750 9158 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 686 9094 750 9158 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 686 9008 750 9072 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 686 9008 750 9072 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 686 8922 750 8986 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 686 8922 750 8986 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 686 8836 750 8900 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 686 8836 750 8900 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 686 8750 750 8814 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 686 8750 750 8814 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 686 8664 750 8728 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 686 8664 750 8728 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 686 8578 750 8642 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 686 8578 750 8642 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 686 8492 750 8556 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 686 8492 750 8556 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 686 8406 750 8470 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 686 8406 750 8470 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 686 8320 750 8384 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 686 8320 750 8384 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 605 9180 669 9244 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 605 9180 669 9244 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 605 9094 669 9158 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 605 9094 669 9158 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 605 9008 669 9072 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 605 9008 669 9072 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 605 8922 669 8986 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 605 8922 669 8986 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 605 8836 669 8900 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 605 8836 669 8900 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 605 8750 669 8814 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 605 8750 669 8814 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 605 8664 669 8728 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 605 8664 669 8728 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 605 8578 669 8642 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 605 8578 669 8642 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 605 8492 669 8556 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 605 8492 669 8556 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 605 8406 669 8470 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 605 8406 669 8470 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 605 8320 669 8384 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 605 8320 669 8384 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 524 9180 588 9244 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 524 9180 588 9244 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 524 9094 588 9158 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 524 9094 588 9158 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 524 9008 588 9072 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 524 9008 588 9072 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 524 8922 588 8986 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 524 8922 588 8986 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 524 8836 588 8900 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 524 8836 588 8900 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 524 8750 588 8814 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 524 8750 588 8814 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 524 8664 588 8728 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 524 8664 588 8728 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 524 8578 588 8642 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 524 8578 588 8642 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 524 8492 588 8556 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 524 8492 588 8556 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 524 8406 588 8470 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 524 8406 588 8470 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 524 8320 588 8384 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 524 8320 588 8384 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 443 9180 507 9244 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 443 9180 507 9244 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 443 9094 507 9158 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 443 9094 507 9158 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 443 9008 507 9072 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 443 9008 507 9072 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 443 8922 507 8986 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 443 8922 507 8986 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 443 8836 507 8900 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 443 8836 507 8900 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 443 8750 507 8814 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 443 8750 507 8814 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 443 8664 507 8728 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 443 8664 507 8728 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 443 8578 507 8642 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 443 8578 507 8642 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 443 8492 507 8556 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 443 8492 507 8556 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 443 8406 507 8470 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 443 8406 507 8470 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 443 8320 507 8384 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 443 8320 507 8384 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 362 9180 426 9244 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 362 9180 426 9244 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 362 9094 426 9158 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 362 9094 426 9158 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 362 9008 426 9072 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 362 9008 426 9072 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 362 8922 426 8986 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 362 8922 426 8986 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 362 8836 426 8900 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 362 8836 426 8900 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 362 8750 426 8814 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 362 8750 426 8814 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 362 8664 426 8728 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 362 8664 426 8728 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 362 8578 426 8642 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 362 8578 426 8642 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 362 8492 426 8556 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 362 8492 426 8556 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 362 8406 426 8470 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 362 8406 426 8470 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 362 8320 426 8384 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 362 8320 426 8384 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 281 9180 345 9244 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 281 9180 345 9244 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 281 9094 345 9158 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 281 9094 345 9158 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 281 9008 345 9072 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 281 9008 345 9072 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 281 8922 345 8986 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 281 8922 345 8986 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 281 8836 345 8900 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 281 8836 345 8900 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 281 8750 345 8814 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 281 8750 345 8814 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 281 8664 345 8728 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 281 8664 345 8728 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 281 8578 345 8642 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 281 8578 345 8642 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 281 8492 345 8556 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 281 8492 345 8556 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 281 8406 345 8470 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 281 8406 345 8470 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 281 8320 345 8384 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 281 8320 345 8384 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 254 9180 264 9244 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 200 9180 264 9244 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 254 9094 264 9158 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 200 9094 264 9158 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 254 9008 264 9072 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 200 9008 264 9072 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 254 8922 264 8986 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 200 8922 264 8986 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 254 8836 264 8900 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 200 8836 264 8900 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 254 8750 264 8814 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 200 8750 264 8814 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 254 8664 264 8728 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 200 8664 264 8728 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 254 8578 264 8642 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 200 8578 264 8642 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 254 8492 264 8556 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 200 8492 264 8556 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 254 8406 264 8470 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 200 8406 264 8470 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 254 8320 264 8384 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 200 8320 264 8384 6 VSSD
port 4 nsew ground bidirectional
rlabel metal5 s 14746 35157 15000 40000 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal5 s 14746 5187 15000 6077 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal5 s 0 35157 254 40000 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal5 s 0 5187 254 6077 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 14746 35157 15000 40000 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 14746 5167 15000 6097 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 0 35157 254 40000 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 0 5167 254 6097 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal5 s 14746 11667 15000 12517 6 VSSIO_Q
port 6 nsew ground bidirectional
rlabel metal5 s 0 11667 254 12517 6 VSSIO_Q
port 6 nsew ground bidirectional
rlabel metal4 s 14746 11647 15000 12537 6 VSSIO_Q
port 6 nsew ground bidirectional
rlabel metal4 s 0 11647 254 12537 6 VSSIO_Q
port 6 nsew ground bidirectional
rlabel metal5 s 14746 6397 15000 7047 6 VSWITCH
port 7 nsew power bidirectional
rlabel metal5 s 0 6397 254 7047 6 VSWITCH
port 7 nsew power bidirectional
rlabel metal4 s 14746 6377 15000 7067 6 VSWITCH
port 7 nsew power bidirectional
rlabel metal4 s 0 6377 254 7067 6 VSWITCH
port 7 nsew power bidirectional
rlabel metal5 s 14746 427 15000 1477 6 VCCHIB
port 8 nsew power bidirectional
rlabel metal5 s 0 427 254 1477 6 VCCHIB
port 8 nsew power bidirectional
rlabel metal4 s 0 407 254 1497 6 VCCHIB
port 8 nsew power bidirectional
rlabel metal4 s 14746 407 15000 1497 6 VCCHIB
port 8 nsew power bidirectional
rlabel metal5 s 14807 3007 15000 3657 6 VDDA
port 9 nsew power bidirectional
rlabel metal5 s 0 3007 193 3657 6 VDDA
port 9 nsew power bidirectional
rlabel metal4 s 14807 2987 15000 3677 6 VDDA
port 9 nsew power bidirectional
rlabel metal4 s 0 2987 193 3677 6 VDDA
port 9 nsew power bidirectional
rlabel metal5 s 14746 14007 15000 18997 6 VDDIO
port 10 nsew power bidirectional
rlabel metal5 s 14746 3977 15000 4867 6 VDDIO
port 10 nsew power bidirectional
rlabel metal5 s 0 14007 254 18997 6 VDDIO
port 10 nsew power bidirectional
rlabel metal5 s 0 3977 254 4867 6 VDDIO
port 10 nsew power bidirectional
rlabel metal4 s 14746 3957 15000 4887 6 VDDIO
port 10 nsew power bidirectional
rlabel metal4 s 14746 14007 15000 19000 6 VDDIO
port 10 nsew power bidirectional
rlabel metal4 s 0 3957 254 4887 6 VDDIO
port 10 nsew power bidirectional
rlabel metal4 s 0 14007 254 19000 6 VDDIO
port 10 nsew power bidirectional
rlabel metal4 s 0 10625 15000 11221 6 AMUXBUS_A
port 11 nsew signal bidirectional
rlabel metal4 s 0 9673 15000 10269 6 AMUXBUS_B
port 12 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 15000 40000
string LEFclass PAD
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_END 2174082
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 2083250
<< end >>
