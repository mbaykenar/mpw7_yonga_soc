magic
tech sky130A
magscale 1 2
timestamp 1649977179
<< labels >>
flabel comment s 62 25 62 25 2 FreeSans 50 0 0 0 EM1O
flabel comment s 118 27 118 27 0 FreeSans 50 0 0 0 B
flabel comment s 50 27 50 27 0 FreeSans 50 0 0 0 A
<< properties >>
string GDS_END 43806398
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 43805630
<< end >>
