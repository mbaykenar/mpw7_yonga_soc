magic
tech sky130B
magscale 1 2
timestamp 1649977179
<< nwell >>
rect -42 416 1632 1116
<< pwell >>
rect 40 118 1550 310
<< mvnmos >>
rect 119 144 239 284
rect 295 144 415 284
rect 471 144 591 284
rect 647 144 767 284
rect 823 144 943 284
rect 999 144 1119 284
rect 1175 144 1295 284
rect 1351 144 1471 284
<< mvpmos >>
rect 119 750 239 950
rect 295 750 415 950
rect 471 750 591 950
rect 647 750 767 950
rect 823 750 943 950
rect 999 750 1119 950
rect 1175 750 1295 950
rect 1351 750 1471 950
rect 119 482 239 682
rect 295 482 415 682
rect 471 482 591 682
rect 647 482 767 682
rect 823 482 943 682
rect 999 482 1119 682
rect 1175 482 1295 682
rect 1351 482 1471 682
<< mvndiff >>
rect 66 272 119 284
rect 66 238 74 272
rect 108 238 119 272
rect 66 204 119 238
rect 66 170 74 204
rect 108 170 119 204
rect 66 144 119 170
rect 239 272 295 284
rect 239 238 250 272
rect 284 238 295 272
rect 239 204 295 238
rect 239 170 250 204
rect 284 170 295 204
rect 239 144 295 170
rect 415 272 471 284
rect 415 238 426 272
rect 460 238 471 272
rect 415 204 471 238
rect 415 170 426 204
rect 460 170 471 204
rect 415 144 471 170
rect 591 272 647 284
rect 591 238 602 272
rect 636 238 647 272
rect 591 204 647 238
rect 591 170 602 204
rect 636 170 647 204
rect 591 144 647 170
rect 767 272 823 284
rect 767 238 778 272
rect 812 238 823 272
rect 767 204 823 238
rect 767 170 778 204
rect 812 170 823 204
rect 767 144 823 170
rect 943 272 999 284
rect 943 238 954 272
rect 988 238 999 272
rect 943 204 999 238
rect 943 170 954 204
rect 988 170 999 204
rect 943 144 999 170
rect 1119 272 1175 284
rect 1119 238 1130 272
rect 1164 238 1175 272
rect 1119 204 1175 238
rect 1119 170 1130 204
rect 1164 170 1175 204
rect 1119 144 1175 170
rect 1295 272 1351 284
rect 1295 238 1306 272
rect 1340 238 1351 272
rect 1295 204 1351 238
rect 1295 170 1306 204
rect 1340 170 1351 204
rect 1295 144 1351 170
rect 1471 272 1524 284
rect 1471 238 1482 272
rect 1516 238 1524 272
rect 1471 204 1524 238
rect 1471 170 1482 204
rect 1516 170 1524 204
rect 1471 144 1524 170
<< mvpdiff >>
rect 66 932 119 950
rect 66 898 74 932
rect 108 898 119 932
rect 66 864 119 898
rect 66 830 74 864
rect 108 830 119 864
rect 66 796 119 830
rect 66 762 74 796
rect 108 762 119 796
rect 66 750 119 762
rect 239 932 295 950
rect 239 898 250 932
rect 284 898 295 932
rect 239 864 295 898
rect 239 830 250 864
rect 284 830 295 864
rect 239 796 295 830
rect 239 762 250 796
rect 284 762 295 796
rect 239 750 295 762
rect 415 932 471 950
rect 415 898 426 932
rect 460 898 471 932
rect 415 864 471 898
rect 415 830 426 864
rect 460 830 471 864
rect 415 796 471 830
rect 415 762 426 796
rect 460 762 471 796
rect 415 750 471 762
rect 591 932 647 950
rect 591 898 602 932
rect 636 898 647 932
rect 591 864 647 898
rect 591 830 602 864
rect 636 830 647 864
rect 591 796 647 830
rect 591 762 602 796
rect 636 762 647 796
rect 591 750 647 762
rect 767 932 823 950
rect 767 898 778 932
rect 812 898 823 932
rect 767 864 823 898
rect 767 830 778 864
rect 812 830 823 864
rect 767 796 823 830
rect 767 762 778 796
rect 812 762 823 796
rect 767 750 823 762
rect 943 932 999 950
rect 943 898 954 932
rect 988 898 999 932
rect 943 864 999 898
rect 943 830 954 864
rect 988 830 999 864
rect 943 796 999 830
rect 943 762 954 796
rect 988 762 999 796
rect 943 750 999 762
rect 1119 932 1175 950
rect 1119 898 1130 932
rect 1164 898 1175 932
rect 1119 864 1175 898
rect 1119 830 1130 864
rect 1164 830 1175 864
rect 1119 796 1175 830
rect 1119 762 1130 796
rect 1164 762 1175 796
rect 1119 750 1175 762
rect 1295 932 1351 950
rect 1295 898 1306 932
rect 1340 898 1351 932
rect 1295 864 1351 898
rect 1295 830 1306 864
rect 1340 830 1351 864
rect 1295 796 1351 830
rect 1295 762 1306 796
rect 1340 762 1351 796
rect 1295 750 1351 762
rect 1471 932 1524 950
rect 1471 898 1482 932
rect 1516 898 1524 932
rect 1471 864 1524 898
rect 1471 830 1482 864
rect 1516 830 1524 864
rect 1471 796 1524 830
rect 1471 762 1482 796
rect 1516 762 1524 796
rect 1471 750 1524 762
rect 66 670 119 682
rect 66 636 74 670
rect 108 636 119 670
rect 66 602 119 636
rect 66 568 74 602
rect 108 568 119 602
rect 66 534 119 568
rect 66 500 74 534
rect 108 500 119 534
rect 66 482 119 500
rect 239 670 295 682
rect 239 636 250 670
rect 284 636 295 670
rect 239 602 295 636
rect 239 568 250 602
rect 284 568 295 602
rect 239 534 295 568
rect 239 500 250 534
rect 284 500 295 534
rect 239 482 295 500
rect 415 670 471 682
rect 415 636 426 670
rect 460 636 471 670
rect 415 602 471 636
rect 415 568 426 602
rect 460 568 471 602
rect 415 534 471 568
rect 415 500 426 534
rect 460 500 471 534
rect 415 482 471 500
rect 591 670 647 682
rect 591 636 602 670
rect 636 636 647 670
rect 591 602 647 636
rect 591 568 602 602
rect 636 568 647 602
rect 591 534 647 568
rect 591 500 602 534
rect 636 500 647 534
rect 591 482 647 500
rect 767 670 823 682
rect 767 636 778 670
rect 812 636 823 670
rect 767 602 823 636
rect 767 568 778 602
rect 812 568 823 602
rect 767 534 823 568
rect 767 500 778 534
rect 812 500 823 534
rect 767 482 823 500
rect 943 670 999 682
rect 943 636 954 670
rect 988 636 999 670
rect 943 602 999 636
rect 943 568 954 602
rect 988 568 999 602
rect 943 534 999 568
rect 943 500 954 534
rect 988 500 999 534
rect 943 482 999 500
rect 1119 670 1175 682
rect 1119 636 1130 670
rect 1164 636 1175 670
rect 1119 602 1175 636
rect 1119 568 1130 602
rect 1164 568 1175 602
rect 1119 534 1175 568
rect 1119 500 1130 534
rect 1164 500 1175 534
rect 1119 482 1175 500
rect 1295 670 1351 682
rect 1295 636 1306 670
rect 1340 636 1351 670
rect 1295 602 1351 636
rect 1295 568 1306 602
rect 1340 568 1351 602
rect 1295 534 1351 568
rect 1295 500 1306 534
rect 1340 500 1351 534
rect 1295 482 1351 500
rect 1471 670 1524 682
rect 1471 636 1482 670
rect 1516 636 1524 670
rect 1471 602 1524 636
rect 1471 568 1482 602
rect 1516 568 1524 602
rect 1471 534 1524 568
rect 1471 500 1482 534
rect 1516 500 1524 534
rect 1471 482 1524 500
<< mvndiffc >>
rect 74 238 108 272
rect 74 170 108 204
rect 250 238 284 272
rect 250 170 284 204
rect 426 238 460 272
rect 426 170 460 204
rect 602 238 636 272
rect 602 170 636 204
rect 778 238 812 272
rect 778 170 812 204
rect 954 238 988 272
rect 954 170 988 204
rect 1130 238 1164 272
rect 1130 170 1164 204
rect 1306 238 1340 272
rect 1306 170 1340 204
rect 1482 238 1516 272
rect 1482 170 1516 204
<< mvpdiffc >>
rect 74 898 108 932
rect 74 830 108 864
rect 74 762 108 796
rect 250 898 284 932
rect 250 830 284 864
rect 250 762 284 796
rect 426 898 460 932
rect 426 830 460 864
rect 426 762 460 796
rect 602 898 636 932
rect 602 830 636 864
rect 602 762 636 796
rect 778 898 812 932
rect 778 830 812 864
rect 778 762 812 796
rect 954 898 988 932
rect 954 830 988 864
rect 954 762 988 796
rect 1130 898 1164 932
rect 1130 830 1164 864
rect 1130 762 1164 796
rect 1306 898 1340 932
rect 1306 830 1340 864
rect 1306 762 1340 796
rect 1482 898 1516 932
rect 1482 830 1516 864
rect 1482 762 1516 796
rect 74 636 108 670
rect 74 568 108 602
rect 74 500 108 534
rect 250 636 284 670
rect 250 568 284 602
rect 250 500 284 534
rect 426 636 460 670
rect 426 568 460 602
rect 426 500 460 534
rect 602 636 636 670
rect 602 568 636 602
rect 602 500 636 534
rect 778 636 812 670
rect 778 568 812 602
rect 778 500 812 534
rect 954 636 988 670
rect 954 568 988 602
rect 954 500 988 534
rect 1130 636 1164 670
rect 1130 568 1164 602
rect 1130 500 1164 534
rect 1306 636 1340 670
rect 1306 568 1340 602
rect 1306 500 1340 534
rect 1482 636 1516 670
rect 1482 568 1516 602
rect 1482 500 1516 534
<< poly >>
rect 119 950 239 976
rect 295 950 415 976
rect 471 950 591 976
rect 647 950 767 976
rect 823 950 943 976
rect 999 950 1119 976
rect 1175 950 1295 976
rect 1351 950 1471 976
rect 119 682 239 750
rect 295 682 415 750
rect 471 682 591 750
rect 647 682 767 750
rect 823 682 943 750
rect 999 682 1119 750
rect 1175 682 1295 750
rect 1351 682 1471 750
rect 119 434 239 482
rect 119 400 166 434
rect 200 400 239 434
rect 119 366 239 400
rect 119 332 166 366
rect 200 332 239 366
rect 119 284 239 332
rect 295 450 415 482
rect 471 450 591 482
rect 295 434 591 450
rect 295 400 318 434
rect 352 400 386 434
rect 420 400 454 434
rect 488 400 522 434
rect 556 400 591 434
rect 295 384 591 400
rect 295 284 415 384
rect 471 284 591 384
rect 647 450 767 482
rect 823 450 943 482
rect 647 434 943 450
rect 647 400 673 434
rect 707 400 741 434
rect 775 400 809 434
rect 843 400 877 434
rect 911 400 943 434
rect 647 384 943 400
rect 647 284 767 384
rect 823 284 943 384
rect 999 450 1119 482
rect 1175 450 1295 482
rect 999 434 1295 450
rect 999 400 1022 434
rect 1056 400 1090 434
rect 1124 400 1158 434
rect 1192 400 1226 434
rect 1260 400 1295 434
rect 999 384 1295 400
rect 999 284 1119 384
rect 1175 284 1295 384
rect 1351 434 1471 482
rect 1351 400 1397 434
rect 1431 400 1471 434
rect 1351 366 1471 400
rect 1351 332 1397 366
rect 1431 332 1471 366
rect 1351 284 1471 332
rect 119 118 239 144
rect 295 118 415 144
rect 471 118 591 144
rect 647 118 767 144
rect 823 118 943 144
rect 999 118 1119 144
rect 1175 118 1295 144
rect 1351 118 1471 144
<< polycont >>
rect 166 400 200 434
rect 166 332 200 366
rect 318 400 352 434
rect 386 400 420 434
rect 454 400 488 434
rect 522 400 556 434
rect 673 400 707 434
rect 741 400 775 434
rect 809 400 843 434
rect 877 400 911 434
rect 1022 400 1056 434
rect 1090 400 1124 434
rect 1158 400 1192 434
rect 1226 400 1260 434
rect 1397 400 1431 434
rect 1397 332 1431 366
<< locali >>
rect 74 932 108 944
rect 74 864 108 872
rect 74 796 108 830
rect 74 670 108 762
rect 74 602 108 636
rect 74 534 108 568
rect 250 932 284 950
rect 250 864 284 898
rect 250 796 284 830
rect 250 670 284 762
rect 250 602 284 636
rect 250 534 284 568
rect 74 484 108 500
rect 249 500 250 519
rect 426 932 460 944
rect 426 864 460 872
rect 426 796 460 830
rect 426 670 460 762
rect 426 602 460 636
rect 426 534 460 568
rect 284 500 287 519
rect 249 485 287 500
rect 602 932 636 950
rect 602 864 636 898
rect 602 796 636 830
rect 602 670 636 762
rect 602 602 636 636
rect 602 534 636 568
rect 150 433 166 434
rect 200 433 216 434
rect 144 400 166 433
rect 144 399 182 400
rect 150 366 216 399
rect 150 332 166 366
rect 200 332 216 366
rect 74 272 108 288
rect 74 227 108 238
rect 74 155 108 170
rect 250 272 284 485
rect 426 484 460 500
rect 600 500 602 519
rect 778 932 812 944
rect 778 864 812 872
rect 778 796 812 830
rect 778 670 812 762
rect 778 602 812 636
rect 778 534 812 568
rect 636 500 638 519
rect 600 485 638 500
rect 954 932 988 950
rect 954 864 988 898
rect 954 796 988 830
rect 954 670 988 762
rect 954 602 988 636
rect 954 534 988 568
rect 318 434 556 450
rect 352 433 386 434
rect 353 400 386 433
rect 420 433 454 434
rect 420 400 421 433
rect 488 400 522 434
rect 318 399 319 400
rect 353 399 421 400
rect 455 399 522 400
rect 318 384 556 399
rect 250 204 284 238
rect 250 154 284 170
rect 426 272 460 288
rect 426 227 460 238
rect 426 155 460 170
rect 602 272 636 485
rect 778 484 812 500
rect 952 500 954 519
rect 1130 932 1164 944
rect 1130 864 1164 872
rect 1130 796 1164 830
rect 1130 670 1164 762
rect 1130 602 1164 636
rect 1130 534 1164 568
rect 988 500 990 519
rect 952 485 990 500
rect 1306 932 1340 950
rect 1306 864 1340 898
rect 1306 796 1340 830
rect 1306 670 1340 762
rect 1306 602 1340 636
rect 1306 534 1340 568
rect 673 434 911 450
rect 707 433 741 434
rect 712 400 741 433
rect 775 433 809 434
rect 673 399 678 400
rect 712 399 775 400
rect 843 433 877 434
rect 843 400 872 433
rect 809 399 872 400
rect 906 399 911 400
rect 673 384 911 399
rect 602 204 636 238
rect 602 154 636 170
rect 778 272 812 288
rect 778 227 812 238
rect 778 155 812 170
rect 954 272 988 485
rect 1130 484 1164 500
rect 1305 500 1306 519
rect 1482 932 1516 944
rect 1482 864 1516 872
rect 1482 796 1516 830
rect 1482 670 1516 762
rect 1482 602 1516 636
rect 1482 534 1516 568
rect 1340 500 1343 519
rect 1305 485 1343 500
rect 1022 434 1260 450
rect 1056 433 1090 434
rect 1057 400 1090 433
rect 1124 433 1158 434
rect 1124 400 1125 433
rect 1192 400 1226 434
rect 1022 399 1023 400
rect 1057 399 1125 400
rect 1159 399 1226 400
rect 1022 384 1260 399
rect 954 204 988 238
rect 954 154 988 170
rect 1130 272 1164 288
rect 1130 227 1164 238
rect 1130 155 1164 170
rect 1306 272 1340 485
rect 1482 484 1516 500
rect 1381 433 1397 434
rect 1431 433 1447 434
rect 1431 400 1446 433
rect 1408 399 1446 400
rect 1381 366 1447 399
rect 1381 332 1397 366
rect 1431 332 1447 366
rect 1306 204 1340 238
rect 1306 154 1340 170
rect 1482 272 1516 288
rect 1482 227 1516 238
rect 1482 155 1516 170
<< viali >>
rect 74 944 108 978
rect 74 898 108 906
rect 74 872 108 898
rect 215 485 249 519
rect 426 944 460 978
rect 426 898 460 906
rect 426 872 460 898
rect 287 485 321 519
rect 110 399 144 433
rect 182 400 200 433
rect 200 400 216 433
rect 182 399 216 400
rect 74 204 108 227
rect 74 193 108 204
rect 74 121 108 155
rect 566 485 600 519
rect 778 944 812 978
rect 778 898 812 906
rect 778 872 812 898
rect 638 485 672 519
rect 319 400 352 433
rect 352 400 353 433
rect 421 400 454 433
rect 454 400 455 433
rect 522 400 556 433
rect 319 399 353 400
rect 421 399 455 400
rect 522 399 556 400
rect 426 204 460 227
rect 426 193 460 204
rect 426 121 460 155
rect 918 485 952 519
rect 1130 944 1164 978
rect 1130 898 1164 906
rect 1130 872 1164 898
rect 990 485 1024 519
rect 678 400 707 433
rect 707 400 712 433
rect 678 399 712 400
rect 775 399 809 433
rect 872 400 877 433
rect 877 400 906 433
rect 872 399 906 400
rect 778 204 812 227
rect 778 193 812 204
rect 778 121 812 155
rect 1271 485 1305 519
rect 1482 944 1516 978
rect 1482 898 1516 906
rect 1482 872 1516 898
rect 1343 485 1377 519
rect 1023 400 1056 433
rect 1056 400 1057 433
rect 1125 400 1158 433
rect 1158 400 1159 433
rect 1226 400 1260 433
rect 1023 399 1057 400
rect 1125 399 1159 400
rect 1226 399 1260 400
rect 1130 204 1164 227
rect 1130 193 1164 204
rect 1130 121 1164 155
rect 1374 400 1397 433
rect 1397 400 1408 433
rect 1374 399 1408 400
rect 1446 399 1480 433
rect 1482 204 1516 227
rect 1482 193 1516 204
rect 1482 121 1516 155
<< metal1 >>
rect 24 978 1566 1062
rect 24 944 74 978
rect 108 944 426 978
rect 460 944 778 978
rect 812 944 1130 978
rect 1164 944 1482 978
rect 1516 944 1566 978
rect 24 906 1566 944
rect 24 872 74 906
rect 108 872 426 906
rect 460 872 778 906
rect 812 872 1130 906
rect 1164 872 1482 906
rect 1516 872 1566 906
rect 24 859 1566 872
rect 203 519 1389 525
rect 203 485 215 519
rect 249 485 287 519
rect 321 485 566 519
rect 600 485 638 519
rect 672 485 918 519
rect 952 485 990 519
rect 1024 485 1271 519
rect 1305 485 1343 519
rect 1377 485 1389 519
rect 203 479 1389 485
rect 98 433 1492 439
rect 98 399 110 433
rect 144 399 182 433
rect 216 399 319 433
rect 353 399 421 433
rect 455 399 522 433
rect 556 399 678 433
rect 712 399 775 433
rect 809 399 872 433
rect 906 399 1023 433
rect 1057 399 1125 433
rect 1159 399 1226 433
rect 1260 399 1374 433
rect 1408 399 1446 433
rect 1480 399 1492 433
rect 98 393 1492 399
rect 24 227 1566 239
rect 24 193 74 227
rect 108 193 426 227
rect 460 193 778 227
rect 812 193 1130 227
rect 1164 193 1482 227
rect 1516 193 1566 227
rect 24 155 1566 193
rect 24 121 74 155
rect 108 121 426 155
rect 460 121 778 155
rect 812 121 1130 155
rect 1164 121 1482 155
rect 1516 121 1566 155
rect 24 24 1566 121
use sky130_fd_pr__model__nfet_highvoltage__example_55959141808613  sky130_fd_pr__model__nfet_highvoltage__example_55959141808613_0
timestamp 1649977179
transform 1 0 119 0 -1 284
box -28 0 1380 63
use sky130_fd_pr__model__pfet_highvoltage__example_55959141808614  sky130_fd_pr__model__pfet_highvoltage__example_55959141808614_0
timestamp 1649977179
transform 1 0 119 0 -1 682
box -28 0 1380 97
use sky130_fd_pr__model__pfet_highvoltage__example_55959141808614  sky130_fd_pr__model__pfet_highvoltage__example_55959141808614_1
timestamp 1649977179
transform 1 0 119 0 1 750
box -28 0 1380 97
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_0
timestamp 1649977179
transform 0 -1 108 1 0 872
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_1
timestamp 1649977179
transform 0 -1 812 1 0 872
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_2
timestamp 1649977179
transform 0 -1 812 -1 0 227
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_3
timestamp 1649977179
transform 0 -1 460 1 0 872
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_4
timestamp 1649977179
transform 0 -1 460 -1 0 227
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_5
timestamp 1649977179
transform 0 -1 108 -1 0 227
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_6
timestamp 1649977179
transform 0 -1 1516 -1 0 227
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_7
timestamp 1649977179
transform 0 -1 1164 -1 0 227
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_8
timestamp 1649977179
transform 0 -1 1516 1 0 872
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_9
timestamp 1649977179
transform 0 -1 1164 1 0 872
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_559591418083  sky130_fd_pr__via_pol1__example_559591418083_0
timestamp 1649977179
transform 0 -1 1447 -1 0 450
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_559591418083  sky130_fd_pr__via_pol1__example_559591418083_1
timestamp 1649977179
transform 0 -1 216 -1 0 450
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_55959141808612  sky130_fd_pr__via_pol1__example_55959141808612_0
timestamp 1649977179
transform 1 0 657 0 1 384
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_55959141808612  sky130_fd_pr__via_pol1__example_55959141808612_1
timestamp 1649977179
transform 1 0 1006 0 1 384
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_55959141808612  sky130_fd_pr__via_pol1__example_55959141808612_2
timestamp 1649977179
transform 1 0 302 0 1 384
box 0 0 1 1
<< labels >>
flabel metal1 s 149 396 200 437 0 FreeSans 400 0 0 0 IN
port 1 nsew
flabel metal1 s 24 1004 1566 1062 3 FreeSans 520 0 0 0 VPWR
port 2 nsew
flabel metal1 s 24 24 1566 82 3 FreeSans 520 0 0 0 VGND
port 3 nsew
flabel metal1 s 352 488 401 522 0 FreeSans 200 0 0 0 OUT
port 4 nsew
<< properties >>
string GDS_END 7978984
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 7972158
<< end >>
