magic
tech sky130A
magscale 1 2
timestamp 1649977179
<< nwell >>
rect -38 261 2062 582
<< pwell >>
rect 1 21 2013 203
rect 30 -17 64 21
<< scnmos >>
rect 79 47 109 177
rect 163 47 193 177
rect 247 47 277 177
rect 331 47 361 177
rect 418 47 448 177
rect 502 47 532 177
rect 586 47 616 177
rect 670 47 700 177
rect 754 47 784 177
rect 838 47 868 177
rect 922 47 952 177
rect 1038 47 1068 177
rect 1194 47 1224 177
rect 1278 47 1308 177
rect 1362 47 1392 177
rect 1446 47 1476 177
rect 1634 47 1664 177
rect 1718 47 1748 177
rect 1802 47 1832 177
rect 1905 47 1935 177
<< scpmoshvt >>
rect 79 297 109 497
rect 163 297 193 497
rect 247 297 277 497
rect 331 297 361 497
rect 418 297 448 497
rect 502 297 532 497
rect 586 297 616 497
rect 670 297 700 497
rect 858 297 888 497
rect 942 297 972 497
rect 1026 297 1056 497
rect 1110 297 1140 497
rect 1194 297 1224 497
rect 1278 297 1308 497
rect 1362 297 1392 497
rect 1446 297 1476 497
rect 1634 297 1664 497
rect 1718 297 1748 497
rect 1802 297 1832 497
rect 1905 297 1935 497
<< ndiff >>
rect 27 161 79 177
rect 27 127 35 161
rect 69 127 79 161
rect 27 93 79 127
rect 27 59 35 93
rect 69 59 79 93
rect 27 47 79 59
rect 109 165 163 177
rect 109 131 119 165
rect 153 131 163 165
rect 109 47 163 131
rect 193 93 247 177
rect 193 59 203 93
rect 237 59 247 93
rect 193 47 247 59
rect 277 165 331 177
rect 277 131 287 165
rect 321 131 331 165
rect 277 47 331 131
rect 361 93 418 177
rect 361 59 371 93
rect 405 59 418 93
rect 361 47 418 59
rect 448 165 502 177
rect 448 131 458 165
rect 492 131 502 165
rect 448 47 502 131
rect 532 93 586 177
rect 532 59 542 93
rect 576 59 586 93
rect 532 47 586 59
rect 616 165 670 177
rect 616 131 626 165
rect 660 131 670 165
rect 616 47 670 131
rect 700 165 754 177
rect 700 131 710 165
rect 744 131 754 165
rect 700 93 754 131
rect 700 59 710 93
rect 744 59 754 93
rect 700 47 754 59
rect 784 93 838 177
rect 784 59 794 93
rect 828 59 838 93
rect 784 47 838 59
rect 868 165 922 177
rect 868 131 878 165
rect 912 131 922 165
rect 868 93 922 131
rect 868 59 878 93
rect 912 59 922 93
rect 868 47 922 59
rect 952 93 1038 177
rect 952 59 978 93
rect 1012 59 1038 93
rect 952 47 1038 59
rect 1068 165 1194 177
rect 1068 131 1078 165
rect 1112 131 1146 165
rect 1180 131 1194 165
rect 1068 93 1194 131
rect 1068 59 1078 93
rect 1112 59 1146 93
rect 1180 59 1194 93
rect 1068 47 1194 59
rect 1224 93 1278 177
rect 1224 59 1234 93
rect 1268 59 1278 93
rect 1224 47 1278 59
rect 1308 165 1362 177
rect 1308 131 1318 165
rect 1352 131 1362 165
rect 1308 93 1362 131
rect 1308 59 1318 93
rect 1352 59 1362 93
rect 1308 47 1362 59
rect 1392 93 1446 177
rect 1392 59 1402 93
rect 1436 59 1446 93
rect 1392 47 1446 59
rect 1476 165 1634 177
rect 1476 131 1486 165
rect 1520 131 1558 165
rect 1592 131 1634 165
rect 1476 93 1634 131
rect 1476 59 1486 93
rect 1520 59 1558 93
rect 1592 59 1634 93
rect 1476 47 1634 59
rect 1664 93 1718 177
rect 1664 59 1674 93
rect 1708 59 1718 93
rect 1664 47 1718 59
rect 1748 165 1802 177
rect 1748 131 1758 165
rect 1792 131 1802 165
rect 1748 93 1802 131
rect 1748 59 1758 93
rect 1792 59 1802 93
rect 1748 47 1802 59
rect 1832 93 1905 177
rect 1832 59 1851 93
rect 1885 59 1905 93
rect 1832 47 1905 59
rect 1935 165 1987 177
rect 1935 131 1945 165
rect 1979 131 1987 165
rect 1935 93 1987 131
rect 1935 59 1945 93
rect 1979 59 1987 93
rect 1935 47 1987 59
<< pdiff >>
rect 27 485 79 497
rect 27 451 35 485
rect 69 451 79 485
rect 27 417 79 451
rect 27 383 35 417
rect 69 383 79 417
rect 27 349 79 383
rect 27 315 35 349
rect 69 315 79 349
rect 27 297 79 315
rect 109 417 163 497
rect 109 383 119 417
rect 153 383 163 417
rect 109 349 163 383
rect 109 315 119 349
rect 153 315 163 349
rect 109 297 163 315
rect 193 485 247 497
rect 193 451 203 485
rect 237 451 247 485
rect 193 417 247 451
rect 193 383 203 417
rect 237 383 247 417
rect 193 297 247 383
rect 277 417 331 497
rect 277 383 287 417
rect 321 383 331 417
rect 277 349 331 383
rect 277 315 287 349
rect 321 315 331 349
rect 277 297 331 315
rect 361 451 418 497
rect 361 417 374 451
rect 408 417 418 451
rect 361 297 418 417
rect 448 485 502 497
rect 448 451 458 485
rect 492 451 502 485
rect 448 297 502 451
rect 532 469 586 497
rect 532 435 542 469
rect 576 435 586 469
rect 532 401 586 435
rect 532 367 542 401
rect 576 367 586 401
rect 532 297 586 367
rect 616 485 670 497
rect 616 451 626 485
rect 660 451 670 485
rect 616 297 670 451
rect 700 469 752 497
rect 700 435 710 469
rect 744 435 752 469
rect 700 401 752 435
rect 700 367 710 401
rect 744 367 752 401
rect 700 297 752 367
rect 806 485 858 497
rect 806 451 814 485
rect 848 451 858 485
rect 806 417 858 451
rect 806 383 814 417
rect 848 383 858 417
rect 806 297 858 383
rect 888 417 942 497
rect 888 383 898 417
rect 932 383 942 417
rect 888 349 942 383
rect 888 315 898 349
rect 932 315 942 349
rect 888 297 942 315
rect 972 485 1026 497
rect 972 451 982 485
rect 1016 451 1026 485
rect 972 417 1026 451
rect 972 383 982 417
rect 1016 383 1026 417
rect 972 297 1026 383
rect 1056 417 1110 497
rect 1056 383 1066 417
rect 1100 383 1110 417
rect 1056 349 1110 383
rect 1056 315 1066 349
rect 1100 315 1110 349
rect 1056 297 1110 315
rect 1140 485 1194 497
rect 1140 451 1150 485
rect 1184 451 1194 485
rect 1140 417 1194 451
rect 1140 383 1150 417
rect 1184 383 1194 417
rect 1140 297 1194 383
rect 1224 417 1278 497
rect 1224 383 1234 417
rect 1268 383 1278 417
rect 1224 349 1278 383
rect 1224 315 1234 349
rect 1268 315 1278 349
rect 1224 297 1278 315
rect 1308 485 1362 497
rect 1308 451 1318 485
rect 1352 451 1362 485
rect 1308 417 1362 451
rect 1308 383 1318 417
rect 1352 383 1362 417
rect 1308 297 1362 383
rect 1392 417 1446 497
rect 1392 383 1402 417
rect 1436 383 1446 417
rect 1392 349 1446 383
rect 1392 315 1402 349
rect 1436 315 1446 349
rect 1392 297 1446 315
rect 1476 485 1528 497
rect 1476 451 1486 485
rect 1520 451 1528 485
rect 1476 417 1528 451
rect 1476 383 1486 417
rect 1520 383 1528 417
rect 1476 297 1528 383
rect 1582 485 1634 497
rect 1582 451 1590 485
rect 1624 451 1634 485
rect 1582 417 1634 451
rect 1582 383 1590 417
rect 1624 383 1634 417
rect 1582 297 1634 383
rect 1664 485 1718 497
rect 1664 451 1674 485
rect 1708 451 1718 485
rect 1664 417 1718 451
rect 1664 383 1674 417
rect 1708 383 1718 417
rect 1664 349 1718 383
rect 1664 315 1674 349
rect 1708 315 1718 349
rect 1664 297 1718 315
rect 1748 485 1802 497
rect 1748 451 1758 485
rect 1792 451 1802 485
rect 1748 417 1802 451
rect 1748 383 1758 417
rect 1792 383 1802 417
rect 1748 297 1802 383
rect 1832 485 1905 497
rect 1832 451 1842 485
rect 1876 451 1905 485
rect 1832 417 1905 451
rect 1832 383 1842 417
rect 1876 383 1905 417
rect 1832 349 1905 383
rect 1832 315 1842 349
rect 1876 315 1905 349
rect 1832 297 1905 315
rect 1935 485 1987 497
rect 1935 451 1945 485
rect 1979 451 1987 485
rect 1935 417 1987 451
rect 1935 383 1945 417
rect 1979 383 1987 417
rect 1935 349 1987 383
rect 1935 315 1945 349
rect 1979 315 1987 349
rect 1935 297 1987 315
<< ndiffc >>
rect 35 127 69 161
rect 35 59 69 93
rect 119 131 153 165
rect 203 59 237 93
rect 287 131 321 165
rect 371 59 405 93
rect 458 131 492 165
rect 542 59 576 93
rect 626 131 660 165
rect 710 131 744 165
rect 710 59 744 93
rect 794 59 828 93
rect 878 131 912 165
rect 878 59 912 93
rect 978 59 1012 93
rect 1078 131 1112 165
rect 1146 131 1180 165
rect 1078 59 1112 93
rect 1146 59 1180 93
rect 1234 59 1268 93
rect 1318 131 1352 165
rect 1318 59 1352 93
rect 1402 59 1436 93
rect 1486 131 1520 165
rect 1558 131 1592 165
rect 1486 59 1520 93
rect 1558 59 1592 93
rect 1674 59 1708 93
rect 1758 131 1792 165
rect 1758 59 1792 93
rect 1851 59 1885 93
rect 1945 131 1979 165
rect 1945 59 1979 93
<< pdiffc >>
rect 35 451 69 485
rect 35 383 69 417
rect 35 315 69 349
rect 119 383 153 417
rect 119 315 153 349
rect 203 451 237 485
rect 203 383 237 417
rect 287 383 321 417
rect 287 315 321 349
rect 374 417 408 451
rect 458 451 492 485
rect 542 435 576 469
rect 542 367 576 401
rect 626 451 660 485
rect 710 435 744 469
rect 710 367 744 401
rect 814 451 848 485
rect 814 383 848 417
rect 898 383 932 417
rect 898 315 932 349
rect 982 451 1016 485
rect 982 383 1016 417
rect 1066 383 1100 417
rect 1066 315 1100 349
rect 1150 451 1184 485
rect 1150 383 1184 417
rect 1234 383 1268 417
rect 1234 315 1268 349
rect 1318 451 1352 485
rect 1318 383 1352 417
rect 1402 383 1436 417
rect 1402 315 1436 349
rect 1486 451 1520 485
rect 1486 383 1520 417
rect 1590 451 1624 485
rect 1590 383 1624 417
rect 1674 451 1708 485
rect 1674 383 1708 417
rect 1674 315 1708 349
rect 1758 451 1792 485
rect 1758 383 1792 417
rect 1842 451 1876 485
rect 1842 383 1876 417
rect 1842 315 1876 349
rect 1945 451 1979 485
rect 1945 383 1979 417
rect 1945 315 1979 349
<< poly >>
rect 79 497 109 523
rect 163 497 193 523
rect 247 497 277 523
rect 331 497 361 523
rect 418 497 448 523
rect 502 497 532 523
rect 586 497 616 523
rect 670 497 700 523
rect 858 497 888 523
rect 942 497 972 523
rect 1026 497 1056 523
rect 1110 497 1140 523
rect 1194 497 1224 523
rect 1278 497 1308 523
rect 1362 497 1392 523
rect 1446 497 1476 523
rect 1634 497 1664 523
rect 1718 497 1748 523
rect 1802 497 1832 523
rect 1905 497 1935 523
rect 79 261 109 297
rect 163 261 193 297
rect 247 261 277 297
rect 331 261 361 297
rect 22 249 361 261
rect 22 215 38 249
rect 72 215 119 249
rect 153 215 203 249
rect 237 215 287 249
rect 321 215 361 249
rect 22 203 361 215
rect 79 177 109 203
rect 163 177 193 203
rect 247 177 277 203
rect 331 177 361 203
rect 418 261 448 297
rect 502 261 532 297
rect 586 261 616 297
rect 670 261 700 297
rect 858 261 888 297
rect 942 261 972 297
rect 1026 261 1056 297
rect 1110 261 1140 297
rect 418 249 700 261
rect 418 215 457 249
rect 491 215 541 249
rect 575 215 626 249
rect 660 215 700 249
rect 418 203 700 215
rect 418 177 448 203
rect 502 177 532 203
rect 586 177 616 203
rect 670 177 700 203
rect 754 249 1140 261
rect 754 215 770 249
rect 804 215 854 249
rect 888 215 938 249
rect 972 215 1022 249
rect 1056 215 1140 249
rect 754 203 1140 215
rect 1194 261 1224 297
rect 1278 261 1308 297
rect 1362 261 1392 297
rect 1446 261 1476 297
rect 1194 249 1476 261
rect 1194 215 1234 249
rect 1268 215 1318 249
rect 1352 215 1402 249
rect 1436 215 1476 249
rect 1194 203 1476 215
rect 754 177 784 203
rect 838 177 868 203
rect 922 177 952 203
rect 1038 177 1068 203
rect 1194 177 1224 203
rect 1278 177 1308 203
rect 1362 177 1392 203
rect 1446 177 1476 203
rect 1634 261 1664 297
rect 1718 261 1748 297
rect 1802 261 1832 297
rect 1905 261 1935 297
rect 1634 249 1976 261
rect 1634 215 1674 249
rect 1708 215 1758 249
rect 1792 215 1842 249
rect 1876 215 1926 249
rect 1960 215 1976 249
rect 1634 203 1976 215
rect 1634 177 1664 203
rect 1718 177 1748 203
rect 1802 177 1832 203
rect 1905 177 1935 203
rect 79 21 109 47
rect 163 21 193 47
rect 247 21 277 47
rect 331 21 361 47
rect 418 21 448 47
rect 502 21 532 47
rect 586 21 616 47
rect 670 21 700 47
rect 754 21 784 47
rect 838 21 868 47
rect 922 21 952 47
rect 1038 21 1068 47
rect 1194 21 1224 47
rect 1278 21 1308 47
rect 1362 21 1392 47
rect 1446 21 1476 47
rect 1634 21 1664 47
rect 1718 21 1748 47
rect 1802 21 1832 47
rect 1905 21 1935 47
<< polycont >>
rect 38 215 72 249
rect 119 215 153 249
rect 203 215 237 249
rect 287 215 321 249
rect 457 215 491 249
rect 541 215 575 249
rect 626 215 660 249
rect 770 215 804 249
rect 854 215 888 249
rect 938 215 972 249
rect 1022 215 1056 249
rect 1234 215 1268 249
rect 1318 215 1352 249
rect 1402 215 1436 249
rect 1674 215 1708 249
rect 1758 215 1792 249
rect 1842 215 1876 249
rect 1926 215 1960 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2024 561
rect 18 485 408 493
rect 18 451 35 485
rect 69 451 203 485
rect 237 451 408 485
rect 18 417 69 451
rect 203 417 237 451
rect 442 485 508 527
rect 610 485 676 527
rect 442 451 458 485
rect 492 451 508 485
rect 442 435 508 451
rect 542 469 576 485
rect 610 451 626 485
rect 660 451 676 485
rect 610 435 676 451
rect 710 469 760 493
rect 744 435 760 469
rect 18 383 35 417
rect 18 349 69 383
rect 18 315 35 349
rect 18 299 69 315
rect 103 383 119 417
rect 153 383 169 417
rect 103 349 169 383
rect 203 367 237 383
rect 271 383 287 417
rect 321 383 340 417
rect 103 315 119 349
rect 153 333 169 349
rect 271 349 340 383
rect 374 401 408 417
rect 542 401 576 435
rect 710 401 760 435
rect 374 367 542 401
rect 576 367 710 401
rect 744 367 760 401
rect 798 485 1536 493
rect 798 451 814 485
rect 848 451 982 485
rect 1016 451 1150 485
rect 1184 451 1318 485
rect 1352 451 1486 485
rect 1520 451 1536 485
rect 798 417 848 451
rect 982 417 1016 451
rect 1150 417 1184 451
rect 1318 417 1352 451
rect 1486 417 1536 451
rect 798 383 814 417
rect 798 367 848 383
rect 882 383 898 417
rect 932 383 948 417
rect 271 333 287 349
rect 153 315 287 333
rect 321 333 340 349
rect 882 349 948 383
rect 982 367 1016 383
rect 1050 383 1066 417
rect 1100 383 1116 417
rect 882 333 898 349
rect 321 315 898 333
rect 932 333 948 349
rect 1050 349 1116 383
rect 1150 367 1184 383
rect 1218 383 1234 417
rect 1268 383 1284 417
rect 1050 333 1066 349
rect 932 315 1066 333
rect 1100 315 1116 349
rect 103 299 1116 315
rect 1218 349 1284 383
rect 1318 367 1352 383
rect 1386 383 1402 417
rect 1436 383 1452 417
rect 1218 315 1234 349
rect 1268 333 1284 349
rect 1386 349 1452 383
rect 1520 383 1536 417
rect 1486 367 1536 383
rect 1574 485 1624 527
rect 1574 451 1590 485
rect 1574 417 1624 451
rect 1574 383 1590 417
rect 1574 367 1624 383
rect 1658 485 1724 493
rect 1658 451 1674 485
rect 1708 451 1724 485
rect 1658 417 1724 451
rect 1658 383 1674 417
rect 1708 383 1724 417
rect 1386 333 1402 349
rect 1268 315 1402 333
rect 1436 333 1452 349
rect 1658 349 1724 383
rect 1758 485 1792 527
rect 1758 417 1792 451
rect 1758 367 1792 383
rect 1826 485 1892 493
rect 1826 451 1842 485
rect 1876 451 1892 485
rect 1826 417 1892 451
rect 1826 383 1842 417
rect 1876 383 1892 417
rect 1658 333 1674 349
rect 1436 315 1674 333
rect 1708 333 1724 349
rect 1826 349 1892 383
rect 1826 333 1842 349
rect 1708 315 1842 333
rect 1876 315 1892 349
rect 1218 299 1892 315
rect 1926 485 2007 527
rect 1926 451 1945 485
rect 1979 451 2007 485
rect 1926 417 2007 451
rect 1926 383 1945 417
rect 1979 383 2007 417
rect 1926 349 2007 383
rect 1926 315 1945 349
rect 1979 315 2007 349
rect 1926 299 2007 315
rect 22 249 337 255
rect 22 215 38 249
rect 72 215 119 249
rect 153 215 203 249
rect 237 215 287 249
rect 321 215 337 249
rect 371 181 407 299
rect 441 249 708 255
rect 441 215 457 249
rect 491 215 541 249
rect 575 215 626 249
rect 660 215 708 249
rect 754 249 1076 255
rect 754 215 770 249
rect 804 215 854 249
rect 888 215 938 249
rect 972 215 1022 249
rect 1056 215 1076 249
rect 1218 249 1452 255
rect 1218 215 1234 249
rect 1268 215 1318 249
rect 1352 215 1402 249
rect 1436 215 1452 249
rect 1658 249 2007 255
rect 1658 215 1674 249
rect 1708 215 1758 249
rect 1792 215 1842 249
rect 1876 215 1926 249
rect 1960 215 2007 249
rect 18 161 69 181
rect 18 127 35 161
rect 103 165 676 181
rect 103 131 119 165
rect 153 131 287 165
rect 321 131 458 165
rect 492 131 626 165
rect 660 131 676 165
rect 710 165 2007 181
rect 744 147 878 165
rect 744 131 760 147
rect 18 93 69 127
rect 710 93 760 131
rect 862 131 878 147
rect 912 147 1078 165
rect 912 131 928 147
rect 18 59 35 93
rect 69 59 203 93
rect 237 59 371 93
rect 405 59 542 93
rect 576 59 710 93
rect 744 59 760 93
rect 18 51 760 59
rect 794 93 828 109
rect 794 17 828 59
rect 862 93 928 131
rect 1062 131 1078 147
rect 1112 131 1146 165
rect 1180 147 1318 165
rect 1180 131 1196 147
rect 862 59 878 93
rect 912 59 928 93
rect 862 51 928 59
rect 962 93 1028 109
rect 962 59 978 93
rect 1012 59 1028 93
rect 962 17 1028 59
rect 1062 93 1196 131
rect 1302 131 1318 147
rect 1352 147 1486 165
rect 1352 131 1368 147
rect 1062 59 1078 93
rect 1112 59 1146 93
rect 1180 59 1196 93
rect 1062 51 1196 59
rect 1234 93 1268 109
rect 1234 17 1268 59
rect 1302 93 1368 131
rect 1470 131 1486 147
rect 1520 131 1558 165
rect 1592 147 1758 165
rect 1592 131 1608 147
rect 1302 59 1318 93
rect 1352 59 1368 93
rect 1302 51 1368 59
rect 1402 93 1436 109
rect 1402 17 1436 59
rect 1470 93 1608 131
rect 1742 131 1758 147
rect 1792 147 1945 165
rect 1792 131 1808 147
rect 1470 59 1486 93
rect 1520 59 1558 93
rect 1592 59 1608 93
rect 1470 51 1608 59
rect 1674 93 1708 109
rect 1674 17 1708 59
rect 1742 93 1808 131
rect 1929 131 1945 147
rect 1979 131 2007 165
rect 1742 59 1758 93
rect 1792 59 1808 93
rect 1742 51 1808 59
rect 1842 93 1894 109
rect 1842 59 1851 93
rect 1885 59 1894 93
rect 1842 17 1894 59
rect 1929 93 2007 131
rect 1929 59 1945 93
rect 1979 59 2007 93
rect 1929 51 2007 59
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2024 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 1593 527 1627 561
rect 1685 527 1719 561
rect 1777 527 1811 561
rect 1869 527 1903 561
rect 1961 527 1995 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1593 -17 1627 17
rect 1685 -17 1719 17
rect 1777 -17 1811 17
rect 1869 -17 1903 17
rect 1961 -17 1995 17
<< metal1 >>
rect 0 561 2024 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2024 561
rect 0 496 2024 527
rect 0 17 2024 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2024 17
rect 0 -48 2024 -17
<< labels >>
flabel locali s 1690 221 1724 255 0 FreeSans 250 0 0 0 A1
port 1 nsew signal input
flabel locali s 1782 221 1816 255 0 FreeSans 250 0 0 0 A1
port 1 nsew signal input
flabel locali s 1874 221 1908 255 0 FreeSans 250 0 0 0 A1
port 1 nsew signal input
flabel locali s 1966 221 2000 255 0 FreeSans 250 0 0 0 A1
port 1 nsew signal input
flabel locali s 1410 221 1444 255 0 FreeSans 250 0 0 0 A2
port 2 nsew signal input
flabel locali s 1318 221 1352 255 0 FreeSans 250 0 0 0 A2
port 2 nsew signal input
flabel locali s 1226 221 1260 255 0 FreeSans 250 0 0 0 A2
port 2 nsew signal input
flabel locali s 1042 221 1076 255 0 FreeSans 250 0 0 0 A3
port 3 nsew signal input
flabel locali s 950 221 984 255 0 FreeSans 250 0 0 0 A3
port 3 nsew signal input
flabel locali s 858 221 892 255 0 FreeSans 250 0 0 0 A3
port 3 nsew signal input
flabel locali s 766 221 800 255 0 FreeSans 250 0 0 0 A3
port 3 nsew signal input
flabel locali s 490 221 524 255 0 FreeSans 250 0 0 0 B1
port 4 nsew signal input
flabel locali s 582 221 616 255 0 FreeSans 250 0 0 0 B1
port 4 nsew signal input
flabel locali s 674 221 708 255 0 FreeSans 250 0 0 0 B1
port 4 nsew signal input
flabel locali s 306 357 340 391 0 FreeSans 250 0 0 0 Y
port 10 nsew signal output
flabel locali s 214 221 248 255 0 FreeSans 250 0 0 0 B2
port 5 nsew signal input
flabel locali s 122 221 156 255 0 FreeSans 250 0 0 0 B2
port 5 nsew signal input
flabel locali s 30 221 64 255 0 FreeSans 250 0 0 0 B2
port 5 nsew signal input
flabel pwell s 30 -17 64 17 0 FreeSans 200 0 0 0 VNB
port 7 nsew ground bidirectional
flabel nwell s 30 527 64 561 0 FreeSans 200 0 0 0 VPB
port 8 nsew power bidirectional
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 6 nsew ground bidirectional abutment
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 9 nsew power bidirectional abutment
rlabel comment s 0 0 0 0 4 o32ai_4
rlabel metal1 s 0 -48 2024 48 1 VGND
port 6 nsew ground bidirectional abutment
rlabel metal1 s 0 496 2024 592 1 VPWR
port 9 nsew power bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 2024 544
string GDS_END 1532130
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 1516152
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string path 0.000 0.000 10.120 0.000 
<< end >>
