magic
tech sky130B
magscale 1 2
timestamp 1649977179
<< metal4 >>
rect 0 13600 2000 18593
rect 0 12410 2000 13300
rect 0 11240 2000 12130
rect 0 10874 2000 10940
rect 0 10218 2000 10814
rect 0 9266 2000 9862
rect 0 9140 2000 9206
rect 0 7910 2000 8840
rect 0 6940 2000 7630
rect 0 5970 2000 6660
rect 0 4760 2000 5690
rect 0 3550 2000 4480
rect 0 2580 2000 3270
rect 0 1370 2000 2300
rect 0 0 2000 1090
<< obsm4 >>
rect 0 34750 2000 39593
rect 0 13380 2000 13520
rect 0 12210 2000 12330
rect 0 11020 2000 11160
rect 0 9922 2000 10158
<< metal5 >>
rect 0 34750 2000 39593
rect 0 13600 2000 18590
rect 0 12430 2000 13280
rect 0 11260 2000 12110
rect 0 9140 2000 10940
rect 0 7930 2000 8820
rect 0 6960 2000 7610
rect 0 5990 2000 6640
rect 0 4780 2000 5670
rect 0 3570 2000 4460
rect 0 2600 2000 3250
rect 0 1390 2000 2280
rect 0 20 2000 1070
<< labels >>
rlabel metal4 s 0 10218 2000 10814 6 AMUXBUS_A
port 1 nsew signal bidirectional
rlabel metal4 s 0 9266 2000 9862 6 AMUXBUS_B
port 2 nsew signal bidirectional
rlabel metal5 s 0 9140 2000 10940 6 VSSA
port 3 nsew ground bidirectional
rlabel metal4 s 0 10874 2000 10940 6 VSSA
port 3 nsew ground bidirectional
rlabel metal4 s 0 9140 2000 9206 6 VSSA
port 3 nsew ground bidirectional
rlabel metal5 s 0 6960 2000 7610 6 VSSA
port 3 nsew ground bidirectional
rlabel metal4 s 0 6940 2000 7630 6 VSSA
port 3 nsew ground bidirectional
rlabel metal5 s 0 2600 2000 3250 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 0 2580 2000 3270 6 VDDA
port 4 nsew power bidirectional
rlabel metal5 s 0 5990 2000 6640 6 VSWITCH
port 5 nsew power bidirectional
rlabel metal4 s 0 5970 2000 6660 6 VSWITCH
port 5 nsew power bidirectional
rlabel metal5 s 0 12430 2000 13280 6 VDDIO_Q
port 6 nsew power bidirectional
rlabel metal4 s 0 12410 2000 13300 6 VDDIO_Q
port 6 nsew power bidirectional
rlabel metal5 s 0 20 2000 1070 6 VCCHIB
port 7 nsew power bidirectional
rlabel metal4 s 0 0 2000 1090 6 VCCHIB
port 7 nsew power bidirectional
rlabel metal5 s 0 13600 2000 18590 6 VDDIO
port 8 nsew power bidirectional
rlabel metal4 s 0 13600 2000 18593 6 VDDIO
port 8 nsew power bidirectional
rlabel metal5 s 0 3570 2000 4460 6 VDDIO
port 8 nsew power bidirectional
rlabel metal4 s 0 3550 2000 4480 6 VDDIO
port 8 nsew power bidirectional
rlabel metal5 s 0 1390 2000 2280 6 VCCD
port 9 nsew power bidirectional
rlabel metal4 s 0 1370 2000 2300 6 VCCD
port 9 nsew power bidirectional
rlabel metal5 s 0 4780 2000 5670 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 0 4760 2000 5690 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal5 s 0 34750 2000 39593 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal5 s 0 7930 2000 8820 6 VSSD
port 11 nsew ground bidirectional
rlabel metal4 s 0 7910 2000 8840 6 VSSD
port 11 nsew ground bidirectional
rlabel metal5 s 0 11260 2000 12110 6 VSSIO_Q
port 12 nsew ground bidirectional
rlabel metal4 s 0 11240 2000 12130 6 VSSIO_Q
port 12 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 2000 39593
string LEFclass PAD SPACER
string LEFview TRUE
string GDS_END 2445150
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_ef_io.gds
string GDS_START 2435886
<< end >>
