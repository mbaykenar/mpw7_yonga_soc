magic
tech sky130B
magscale 12 1
timestamp 1598775307
<< metal5 >>
rect 0 70 40 75
rect 0 60 45 70
rect 30 45 45 60
rect 5 40 45 45
rect 0 30 45 40
rect 0 15 15 30
rect 30 15 45 30
rect 0 5 45 15
rect 5 0 45 5
<< properties >>
string FIXED_BBOX 0 -30 60 105
<< end >>
