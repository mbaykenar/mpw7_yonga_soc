magic
tech sky130B
magscale 1 2
timestamp 1649977179
<< metal3 >>
rect 100 8844 4900 8846
rect 100 8780 106 8844
rect 170 8780 187 8844
rect 251 8780 268 8844
rect 332 8780 349 8844
rect 413 8780 430 8844
rect 494 8780 510 8844
rect 574 8780 590 8844
rect 654 8780 670 8844
rect 734 8780 750 8844
rect 814 8780 830 8844
rect 894 8780 910 8844
rect 974 8780 990 8844
rect 1054 8780 1070 8844
rect 1134 8780 1150 8844
rect 1214 8780 1230 8844
rect 1294 8780 1310 8844
rect 1374 8780 1390 8844
rect 1454 8780 1470 8844
rect 1534 8780 1550 8844
rect 1614 8780 1630 8844
rect 1694 8780 1710 8844
rect 1774 8780 1790 8844
rect 1854 8780 1870 8844
rect 1934 8780 1950 8844
rect 2014 8780 2030 8844
rect 2094 8780 2110 8844
rect 2174 8780 2190 8844
rect 2254 8780 2270 8844
rect 2334 8780 2350 8844
rect 2414 8780 2430 8844
rect 2494 8780 2510 8844
rect 2574 8780 2590 8844
rect 2654 8780 2670 8844
rect 2734 8780 2750 8844
rect 2814 8780 2830 8844
rect 2894 8780 2910 8844
rect 2974 8780 2990 8844
rect 3054 8780 3070 8844
rect 3134 8780 3150 8844
rect 3214 8780 3230 8844
rect 3294 8780 3310 8844
rect 3374 8780 3390 8844
rect 3454 8780 3470 8844
rect 3534 8780 3550 8844
rect 3614 8780 3630 8844
rect 3694 8780 3710 8844
rect 3774 8780 3790 8844
rect 3854 8780 3870 8844
rect 3934 8780 3950 8844
rect 4014 8780 4030 8844
rect 4094 8780 4110 8844
rect 4174 8780 4190 8844
rect 4254 8780 4270 8844
rect 4334 8780 4350 8844
rect 4414 8780 4430 8844
rect 4494 8780 4510 8844
rect 4574 8780 4590 8844
rect 4654 8780 4670 8844
rect 4734 8780 4750 8844
rect 4814 8780 4830 8844
rect 4894 8780 4900 8844
rect 100 8758 4900 8780
rect 100 8694 106 8758
rect 170 8694 187 8758
rect 251 8694 268 8758
rect 332 8694 349 8758
rect 413 8694 430 8758
rect 494 8694 510 8758
rect 574 8694 590 8758
rect 654 8694 670 8758
rect 734 8694 750 8758
rect 814 8694 830 8758
rect 894 8694 910 8758
rect 974 8694 990 8758
rect 1054 8694 1070 8758
rect 1134 8694 1150 8758
rect 1214 8694 1230 8758
rect 1294 8694 1310 8758
rect 1374 8694 1390 8758
rect 1454 8694 1470 8758
rect 1534 8694 1550 8758
rect 1614 8694 1630 8758
rect 1694 8694 1710 8758
rect 1774 8694 1790 8758
rect 1854 8694 1870 8758
rect 1934 8694 1950 8758
rect 2014 8694 2030 8758
rect 2094 8694 2110 8758
rect 2174 8694 2190 8758
rect 2254 8694 2270 8758
rect 2334 8694 2350 8758
rect 2414 8694 2430 8758
rect 2494 8694 2510 8758
rect 2574 8694 2590 8758
rect 2654 8694 2670 8758
rect 2734 8694 2750 8758
rect 2814 8694 2830 8758
rect 2894 8694 2910 8758
rect 2974 8694 2990 8758
rect 3054 8694 3070 8758
rect 3134 8694 3150 8758
rect 3214 8694 3230 8758
rect 3294 8694 3310 8758
rect 3374 8694 3390 8758
rect 3454 8694 3470 8758
rect 3534 8694 3550 8758
rect 3614 8694 3630 8758
rect 3694 8694 3710 8758
rect 3774 8694 3790 8758
rect 3854 8694 3870 8758
rect 3934 8694 3950 8758
rect 4014 8694 4030 8758
rect 4094 8694 4110 8758
rect 4174 8694 4190 8758
rect 4254 8694 4270 8758
rect 4334 8694 4350 8758
rect 4414 8694 4430 8758
rect 4494 8694 4510 8758
rect 4574 8694 4590 8758
rect 4654 8694 4670 8758
rect 4734 8694 4750 8758
rect 4814 8694 4830 8758
rect 4894 8694 4900 8758
rect 100 8672 4900 8694
rect 100 8608 106 8672
rect 170 8608 187 8672
rect 251 8608 268 8672
rect 332 8608 349 8672
rect 413 8608 430 8672
rect 494 8608 510 8672
rect 574 8608 590 8672
rect 654 8608 670 8672
rect 734 8608 750 8672
rect 814 8608 830 8672
rect 894 8608 910 8672
rect 974 8608 990 8672
rect 1054 8608 1070 8672
rect 1134 8608 1150 8672
rect 1214 8608 1230 8672
rect 1294 8608 1310 8672
rect 1374 8608 1390 8672
rect 1454 8608 1470 8672
rect 1534 8608 1550 8672
rect 1614 8608 1630 8672
rect 1694 8608 1710 8672
rect 1774 8608 1790 8672
rect 1854 8608 1870 8672
rect 1934 8608 1950 8672
rect 2014 8608 2030 8672
rect 2094 8608 2110 8672
rect 2174 8608 2190 8672
rect 2254 8608 2270 8672
rect 2334 8608 2350 8672
rect 2414 8608 2430 8672
rect 2494 8608 2510 8672
rect 2574 8608 2590 8672
rect 2654 8608 2670 8672
rect 2734 8608 2750 8672
rect 2814 8608 2830 8672
rect 2894 8608 2910 8672
rect 2974 8608 2990 8672
rect 3054 8608 3070 8672
rect 3134 8608 3150 8672
rect 3214 8608 3230 8672
rect 3294 8608 3310 8672
rect 3374 8608 3390 8672
rect 3454 8608 3470 8672
rect 3534 8608 3550 8672
rect 3614 8608 3630 8672
rect 3694 8608 3710 8672
rect 3774 8608 3790 8672
rect 3854 8608 3870 8672
rect 3934 8608 3950 8672
rect 4014 8608 4030 8672
rect 4094 8608 4110 8672
rect 4174 8608 4190 8672
rect 4254 8608 4270 8672
rect 4334 8608 4350 8672
rect 4414 8608 4430 8672
rect 4494 8608 4510 8672
rect 4574 8608 4590 8672
rect 4654 8608 4670 8672
rect 4734 8608 4750 8672
rect 4814 8608 4830 8672
rect 4894 8608 4900 8672
rect 100 8586 4900 8608
rect 100 8522 106 8586
rect 170 8522 187 8586
rect 251 8522 268 8586
rect 332 8522 349 8586
rect 413 8522 430 8586
rect 494 8522 510 8586
rect 574 8522 590 8586
rect 654 8522 670 8586
rect 734 8522 750 8586
rect 814 8522 830 8586
rect 894 8522 910 8586
rect 974 8522 990 8586
rect 1054 8522 1070 8586
rect 1134 8522 1150 8586
rect 1214 8522 1230 8586
rect 1294 8522 1310 8586
rect 1374 8522 1390 8586
rect 1454 8522 1470 8586
rect 1534 8522 1550 8586
rect 1614 8522 1630 8586
rect 1694 8522 1710 8586
rect 1774 8522 1790 8586
rect 1854 8522 1870 8586
rect 1934 8522 1950 8586
rect 2014 8522 2030 8586
rect 2094 8522 2110 8586
rect 2174 8522 2190 8586
rect 2254 8522 2270 8586
rect 2334 8522 2350 8586
rect 2414 8522 2430 8586
rect 2494 8522 2510 8586
rect 2574 8522 2590 8586
rect 2654 8522 2670 8586
rect 2734 8522 2750 8586
rect 2814 8522 2830 8586
rect 2894 8522 2910 8586
rect 2974 8522 2990 8586
rect 3054 8522 3070 8586
rect 3134 8522 3150 8586
rect 3214 8522 3230 8586
rect 3294 8522 3310 8586
rect 3374 8522 3390 8586
rect 3454 8522 3470 8586
rect 3534 8522 3550 8586
rect 3614 8522 3630 8586
rect 3694 8522 3710 8586
rect 3774 8522 3790 8586
rect 3854 8522 3870 8586
rect 3934 8522 3950 8586
rect 4014 8522 4030 8586
rect 4094 8522 4110 8586
rect 4174 8522 4190 8586
rect 4254 8522 4270 8586
rect 4334 8522 4350 8586
rect 4414 8522 4430 8586
rect 4494 8522 4510 8586
rect 4574 8522 4590 8586
rect 4654 8522 4670 8586
rect 4734 8522 4750 8586
rect 4814 8522 4830 8586
rect 4894 8522 4900 8586
rect 100 8500 4900 8522
rect 100 8436 106 8500
rect 170 8436 187 8500
rect 251 8436 268 8500
rect 332 8436 349 8500
rect 413 8436 430 8500
rect 494 8436 510 8500
rect 574 8436 590 8500
rect 654 8436 670 8500
rect 734 8436 750 8500
rect 814 8436 830 8500
rect 894 8436 910 8500
rect 974 8436 990 8500
rect 1054 8436 1070 8500
rect 1134 8436 1150 8500
rect 1214 8436 1230 8500
rect 1294 8436 1310 8500
rect 1374 8436 1390 8500
rect 1454 8436 1470 8500
rect 1534 8436 1550 8500
rect 1614 8436 1630 8500
rect 1694 8436 1710 8500
rect 1774 8436 1790 8500
rect 1854 8436 1870 8500
rect 1934 8436 1950 8500
rect 2014 8436 2030 8500
rect 2094 8436 2110 8500
rect 2174 8436 2190 8500
rect 2254 8436 2270 8500
rect 2334 8436 2350 8500
rect 2414 8436 2430 8500
rect 2494 8436 2510 8500
rect 2574 8436 2590 8500
rect 2654 8436 2670 8500
rect 2734 8436 2750 8500
rect 2814 8436 2830 8500
rect 2894 8436 2910 8500
rect 2974 8436 2990 8500
rect 3054 8436 3070 8500
rect 3134 8436 3150 8500
rect 3214 8436 3230 8500
rect 3294 8436 3310 8500
rect 3374 8436 3390 8500
rect 3454 8436 3470 8500
rect 3534 8436 3550 8500
rect 3614 8436 3630 8500
rect 3694 8436 3710 8500
rect 3774 8436 3790 8500
rect 3854 8436 3870 8500
rect 3934 8436 3950 8500
rect 4014 8436 4030 8500
rect 4094 8436 4110 8500
rect 4174 8436 4190 8500
rect 4254 8436 4270 8500
rect 4334 8436 4350 8500
rect 4414 8436 4430 8500
rect 4494 8436 4510 8500
rect 4574 8436 4590 8500
rect 4654 8436 4670 8500
rect 4734 8436 4750 8500
rect 4814 8436 4830 8500
rect 4894 8436 4900 8500
rect 100 8414 4900 8436
rect 100 8350 106 8414
rect 170 8350 187 8414
rect 251 8350 268 8414
rect 332 8350 349 8414
rect 413 8350 430 8414
rect 494 8350 510 8414
rect 574 8350 590 8414
rect 654 8350 670 8414
rect 734 8350 750 8414
rect 814 8350 830 8414
rect 894 8350 910 8414
rect 974 8350 990 8414
rect 1054 8350 1070 8414
rect 1134 8350 1150 8414
rect 1214 8350 1230 8414
rect 1294 8350 1310 8414
rect 1374 8350 1390 8414
rect 1454 8350 1470 8414
rect 1534 8350 1550 8414
rect 1614 8350 1630 8414
rect 1694 8350 1710 8414
rect 1774 8350 1790 8414
rect 1854 8350 1870 8414
rect 1934 8350 1950 8414
rect 2014 8350 2030 8414
rect 2094 8350 2110 8414
rect 2174 8350 2190 8414
rect 2254 8350 2270 8414
rect 2334 8350 2350 8414
rect 2414 8350 2430 8414
rect 2494 8350 2510 8414
rect 2574 8350 2590 8414
rect 2654 8350 2670 8414
rect 2734 8350 2750 8414
rect 2814 8350 2830 8414
rect 2894 8350 2910 8414
rect 2974 8350 2990 8414
rect 3054 8350 3070 8414
rect 3134 8350 3150 8414
rect 3214 8350 3230 8414
rect 3294 8350 3310 8414
rect 3374 8350 3390 8414
rect 3454 8350 3470 8414
rect 3534 8350 3550 8414
rect 3614 8350 3630 8414
rect 3694 8350 3710 8414
rect 3774 8350 3790 8414
rect 3854 8350 3870 8414
rect 3934 8350 3950 8414
rect 4014 8350 4030 8414
rect 4094 8350 4110 8414
rect 4174 8350 4190 8414
rect 4254 8350 4270 8414
rect 4334 8350 4350 8414
rect 4414 8350 4430 8414
rect 4494 8350 4510 8414
rect 4574 8350 4590 8414
rect 4654 8350 4670 8414
rect 4734 8350 4750 8414
rect 4814 8350 4830 8414
rect 4894 8350 4900 8414
rect 100 8328 4900 8350
rect 100 8264 106 8328
rect 170 8264 187 8328
rect 251 8264 268 8328
rect 332 8264 349 8328
rect 413 8264 430 8328
rect 494 8264 510 8328
rect 574 8264 590 8328
rect 654 8264 670 8328
rect 734 8264 750 8328
rect 814 8264 830 8328
rect 894 8264 910 8328
rect 974 8264 990 8328
rect 1054 8264 1070 8328
rect 1134 8264 1150 8328
rect 1214 8264 1230 8328
rect 1294 8264 1310 8328
rect 1374 8264 1390 8328
rect 1454 8264 1470 8328
rect 1534 8264 1550 8328
rect 1614 8264 1630 8328
rect 1694 8264 1710 8328
rect 1774 8264 1790 8328
rect 1854 8264 1870 8328
rect 1934 8264 1950 8328
rect 2014 8264 2030 8328
rect 2094 8264 2110 8328
rect 2174 8264 2190 8328
rect 2254 8264 2270 8328
rect 2334 8264 2350 8328
rect 2414 8264 2430 8328
rect 2494 8264 2510 8328
rect 2574 8264 2590 8328
rect 2654 8264 2670 8328
rect 2734 8264 2750 8328
rect 2814 8264 2830 8328
rect 2894 8264 2910 8328
rect 2974 8264 2990 8328
rect 3054 8264 3070 8328
rect 3134 8264 3150 8328
rect 3214 8264 3230 8328
rect 3294 8264 3310 8328
rect 3374 8264 3390 8328
rect 3454 8264 3470 8328
rect 3534 8264 3550 8328
rect 3614 8264 3630 8328
rect 3694 8264 3710 8328
rect 3774 8264 3790 8328
rect 3854 8264 3870 8328
rect 3934 8264 3950 8328
rect 4014 8264 4030 8328
rect 4094 8264 4110 8328
rect 4174 8264 4190 8328
rect 4254 8264 4270 8328
rect 4334 8264 4350 8328
rect 4414 8264 4430 8328
rect 4494 8264 4510 8328
rect 4574 8264 4590 8328
rect 4654 8264 4670 8328
rect 4734 8264 4750 8328
rect 4814 8264 4830 8328
rect 4894 8264 4900 8328
rect 100 8242 4900 8264
rect 100 8178 106 8242
rect 170 8178 187 8242
rect 251 8178 268 8242
rect 332 8178 349 8242
rect 413 8178 430 8242
rect 494 8178 510 8242
rect 574 8178 590 8242
rect 654 8178 670 8242
rect 734 8178 750 8242
rect 814 8178 830 8242
rect 894 8178 910 8242
rect 974 8178 990 8242
rect 1054 8178 1070 8242
rect 1134 8178 1150 8242
rect 1214 8178 1230 8242
rect 1294 8178 1310 8242
rect 1374 8178 1390 8242
rect 1454 8178 1470 8242
rect 1534 8178 1550 8242
rect 1614 8178 1630 8242
rect 1694 8178 1710 8242
rect 1774 8178 1790 8242
rect 1854 8178 1870 8242
rect 1934 8178 1950 8242
rect 2014 8178 2030 8242
rect 2094 8178 2110 8242
rect 2174 8178 2190 8242
rect 2254 8178 2270 8242
rect 2334 8178 2350 8242
rect 2414 8178 2430 8242
rect 2494 8178 2510 8242
rect 2574 8178 2590 8242
rect 2654 8178 2670 8242
rect 2734 8178 2750 8242
rect 2814 8178 2830 8242
rect 2894 8178 2910 8242
rect 2974 8178 2990 8242
rect 3054 8178 3070 8242
rect 3134 8178 3150 8242
rect 3214 8178 3230 8242
rect 3294 8178 3310 8242
rect 3374 8178 3390 8242
rect 3454 8178 3470 8242
rect 3534 8178 3550 8242
rect 3614 8178 3630 8242
rect 3694 8178 3710 8242
rect 3774 8178 3790 8242
rect 3854 8178 3870 8242
rect 3934 8178 3950 8242
rect 4014 8178 4030 8242
rect 4094 8178 4110 8242
rect 4174 8178 4190 8242
rect 4254 8178 4270 8242
rect 4334 8178 4350 8242
rect 4414 8178 4430 8242
rect 4494 8178 4510 8242
rect 4574 8178 4590 8242
rect 4654 8178 4670 8242
rect 4734 8178 4750 8242
rect 4814 8178 4830 8242
rect 4894 8178 4900 8242
rect 100 8156 4900 8178
rect 100 8092 106 8156
rect 170 8092 187 8156
rect 251 8092 268 8156
rect 332 8092 349 8156
rect 413 8092 430 8156
rect 494 8092 510 8156
rect 574 8092 590 8156
rect 654 8092 670 8156
rect 734 8092 750 8156
rect 814 8092 830 8156
rect 894 8092 910 8156
rect 974 8092 990 8156
rect 1054 8092 1070 8156
rect 1134 8092 1150 8156
rect 1214 8092 1230 8156
rect 1294 8092 1310 8156
rect 1374 8092 1390 8156
rect 1454 8092 1470 8156
rect 1534 8092 1550 8156
rect 1614 8092 1630 8156
rect 1694 8092 1710 8156
rect 1774 8092 1790 8156
rect 1854 8092 1870 8156
rect 1934 8092 1950 8156
rect 2014 8092 2030 8156
rect 2094 8092 2110 8156
rect 2174 8092 2190 8156
rect 2254 8092 2270 8156
rect 2334 8092 2350 8156
rect 2414 8092 2430 8156
rect 2494 8092 2510 8156
rect 2574 8092 2590 8156
rect 2654 8092 2670 8156
rect 2734 8092 2750 8156
rect 2814 8092 2830 8156
rect 2894 8092 2910 8156
rect 2974 8092 2990 8156
rect 3054 8092 3070 8156
rect 3134 8092 3150 8156
rect 3214 8092 3230 8156
rect 3294 8092 3310 8156
rect 3374 8092 3390 8156
rect 3454 8092 3470 8156
rect 3534 8092 3550 8156
rect 3614 8092 3630 8156
rect 3694 8092 3710 8156
rect 3774 8092 3790 8156
rect 3854 8092 3870 8156
rect 3934 8092 3950 8156
rect 4014 8092 4030 8156
rect 4094 8092 4110 8156
rect 4174 8092 4190 8156
rect 4254 8092 4270 8156
rect 4334 8092 4350 8156
rect 4414 8092 4430 8156
rect 4494 8092 4510 8156
rect 4574 8092 4590 8156
rect 4654 8092 4670 8156
rect 4734 8092 4750 8156
rect 4814 8092 4830 8156
rect 4894 8092 4900 8156
rect 100 8070 4900 8092
rect 100 8006 106 8070
rect 170 8006 187 8070
rect 251 8006 268 8070
rect 332 8006 349 8070
rect 413 8006 430 8070
rect 494 8006 510 8070
rect 574 8006 590 8070
rect 654 8006 670 8070
rect 734 8006 750 8070
rect 814 8006 830 8070
rect 894 8006 910 8070
rect 974 8006 990 8070
rect 1054 8006 1070 8070
rect 1134 8006 1150 8070
rect 1214 8006 1230 8070
rect 1294 8006 1310 8070
rect 1374 8006 1390 8070
rect 1454 8006 1470 8070
rect 1534 8006 1550 8070
rect 1614 8006 1630 8070
rect 1694 8006 1710 8070
rect 1774 8006 1790 8070
rect 1854 8006 1870 8070
rect 1934 8006 1950 8070
rect 2014 8006 2030 8070
rect 2094 8006 2110 8070
rect 2174 8006 2190 8070
rect 2254 8006 2270 8070
rect 2334 8006 2350 8070
rect 2414 8006 2430 8070
rect 2494 8006 2510 8070
rect 2574 8006 2590 8070
rect 2654 8006 2670 8070
rect 2734 8006 2750 8070
rect 2814 8006 2830 8070
rect 2894 8006 2910 8070
rect 2974 8006 2990 8070
rect 3054 8006 3070 8070
rect 3134 8006 3150 8070
rect 3214 8006 3230 8070
rect 3294 8006 3310 8070
rect 3374 8006 3390 8070
rect 3454 8006 3470 8070
rect 3534 8006 3550 8070
rect 3614 8006 3630 8070
rect 3694 8006 3710 8070
rect 3774 8006 3790 8070
rect 3854 8006 3870 8070
rect 3934 8006 3950 8070
rect 4014 8006 4030 8070
rect 4094 8006 4110 8070
rect 4174 8006 4190 8070
rect 4254 8006 4270 8070
rect 4334 8006 4350 8070
rect 4414 8006 4430 8070
rect 4494 8006 4510 8070
rect 4574 8006 4590 8070
rect 4654 8006 4670 8070
rect 4734 8006 4750 8070
rect 4814 8006 4830 8070
rect 4894 8006 4900 8070
rect 100 7984 4900 8006
rect 100 7920 106 7984
rect 170 7920 187 7984
rect 251 7920 268 7984
rect 332 7920 349 7984
rect 413 7920 430 7984
rect 494 7920 510 7984
rect 574 7920 590 7984
rect 654 7920 670 7984
rect 734 7920 750 7984
rect 814 7920 830 7984
rect 894 7920 910 7984
rect 974 7920 990 7984
rect 1054 7920 1070 7984
rect 1134 7920 1150 7984
rect 1214 7920 1230 7984
rect 1294 7920 1310 7984
rect 1374 7920 1390 7984
rect 1454 7920 1470 7984
rect 1534 7920 1550 7984
rect 1614 7920 1630 7984
rect 1694 7920 1710 7984
rect 1774 7920 1790 7984
rect 1854 7920 1870 7984
rect 1934 7920 1950 7984
rect 2014 7920 2030 7984
rect 2094 7920 2110 7984
rect 2174 7920 2190 7984
rect 2254 7920 2270 7984
rect 2334 7920 2350 7984
rect 2414 7920 2430 7984
rect 2494 7920 2510 7984
rect 2574 7920 2590 7984
rect 2654 7920 2670 7984
rect 2734 7920 2750 7984
rect 2814 7920 2830 7984
rect 2894 7920 2910 7984
rect 2974 7920 2990 7984
rect 3054 7920 3070 7984
rect 3134 7920 3150 7984
rect 3214 7920 3230 7984
rect 3294 7920 3310 7984
rect 3374 7920 3390 7984
rect 3454 7920 3470 7984
rect 3534 7920 3550 7984
rect 3614 7920 3630 7984
rect 3694 7920 3710 7984
rect 3774 7920 3790 7984
rect 3854 7920 3870 7984
rect 3934 7920 3950 7984
rect 4014 7920 4030 7984
rect 4094 7920 4110 7984
rect 4174 7920 4190 7984
rect 4254 7920 4270 7984
rect 4334 7920 4350 7984
rect 4414 7920 4430 7984
rect 4494 7920 4510 7984
rect 4574 7920 4590 7984
rect 4654 7920 4670 7984
rect 4734 7920 4750 7984
rect 4814 7920 4830 7984
rect 4894 7920 4900 7984
rect 100 7918 4900 7920
rect 10151 8844 14940 8846
rect 10151 8780 10157 8844
rect 10221 8780 10239 8844
rect 10303 8780 10321 8844
rect 10385 8780 10403 8844
rect 10467 8780 10485 8844
rect 10549 8780 10567 8844
rect 10631 8780 10649 8844
rect 10713 8780 10731 8844
rect 10795 8780 10813 8844
rect 10877 8780 10895 8844
rect 10959 8780 10977 8844
rect 11041 8780 11059 8844
rect 11123 8780 11141 8844
rect 11205 8780 11223 8844
rect 11287 8780 11305 8844
rect 11369 8780 11387 8844
rect 11451 8780 11468 8844
rect 11532 8780 11549 8844
rect 11613 8780 11630 8844
rect 11694 8780 11711 8844
rect 11775 8780 11792 8844
rect 11856 8780 11873 8844
rect 11937 8780 11954 8844
rect 12018 8780 12035 8844
rect 12099 8780 12116 8844
rect 12180 8780 12197 8844
rect 12261 8780 12278 8844
rect 12342 8780 12359 8844
rect 12423 8780 12440 8844
rect 12504 8780 12521 8844
rect 12585 8780 12602 8844
rect 12666 8780 12683 8844
rect 12747 8780 12764 8844
rect 12828 8780 12845 8844
rect 12909 8780 12926 8844
rect 12990 8780 13007 8844
rect 13071 8780 13088 8844
rect 13152 8780 13169 8844
rect 13233 8780 13250 8844
rect 13314 8780 13331 8844
rect 13395 8780 13412 8844
rect 13476 8780 13493 8844
rect 13557 8780 13574 8844
rect 13638 8780 13655 8844
rect 13719 8780 13736 8844
rect 13800 8780 13817 8844
rect 13881 8780 13898 8844
rect 13962 8780 13979 8844
rect 14043 8780 14060 8844
rect 14124 8780 14141 8844
rect 14205 8780 14222 8844
rect 14286 8780 14303 8844
rect 14367 8780 14384 8844
rect 14448 8780 14465 8844
rect 14529 8780 14546 8844
rect 14610 8780 14627 8844
rect 14691 8780 14708 8844
rect 14772 8780 14789 8844
rect 14853 8780 14870 8844
rect 14934 8780 14940 8844
rect 10151 8758 14940 8780
rect 10151 8694 10157 8758
rect 10221 8694 10239 8758
rect 10303 8694 10321 8758
rect 10385 8694 10403 8758
rect 10467 8694 10485 8758
rect 10549 8694 10567 8758
rect 10631 8694 10649 8758
rect 10713 8694 10731 8758
rect 10795 8694 10813 8758
rect 10877 8694 10895 8758
rect 10959 8694 10977 8758
rect 11041 8694 11059 8758
rect 11123 8694 11141 8758
rect 11205 8694 11223 8758
rect 11287 8694 11305 8758
rect 11369 8694 11387 8758
rect 11451 8694 11468 8758
rect 11532 8694 11549 8758
rect 11613 8694 11630 8758
rect 11694 8694 11711 8758
rect 11775 8694 11792 8758
rect 11856 8694 11873 8758
rect 11937 8694 11954 8758
rect 12018 8694 12035 8758
rect 12099 8694 12116 8758
rect 12180 8694 12197 8758
rect 12261 8694 12278 8758
rect 12342 8694 12359 8758
rect 12423 8694 12440 8758
rect 12504 8694 12521 8758
rect 12585 8694 12602 8758
rect 12666 8694 12683 8758
rect 12747 8694 12764 8758
rect 12828 8694 12845 8758
rect 12909 8694 12926 8758
rect 12990 8694 13007 8758
rect 13071 8694 13088 8758
rect 13152 8694 13169 8758
rect 13233 8694 13250 8758
rect 13314 8694 13331 8758
rect 13395 8694 13412 8758
rect 13476 8694 13493 8758
rect 13557 8694 13574 8758
rect 13638 8694 13655 8758
rect 13719 8694 13736 8758
rect 13800 8694 13817 8758
rect 13881 8694 13898 8758
rect 13962 8694 13979 8758
rect 14043 8694 14060 8758
rect 14124 8694 14141 8758
rect 14205 8694 14222 8758
rect 14286 8694 14303 8758
rect 14367 8694 14384 8758
rect 14448 8694 14465 8758
rect 14529 8694 14546 8758
rect 14610 8694 14627 8758
rect 14691 8694 14708 8758
rect 14772 8694 14789 8758
rect 14853 8694 14870 8758
rect 14934 8694 14940 8758
rect 10151 8672 14940 8694
rect 10151 8608 10157 8672
rect 10221 8608 10239 8672
rect 10303 8608 10321 8672
rect 10385 8608 10403 8672
rect 10467 8608 10485 8672
rect 10549 8608 10567 8672
rect 10631 8608 10649 8672
rect 10713 8608 10731 8672
rect 10795 8608 10813 8672
rect 10877 8608 10895 8672
rect 10959 8608 10977 8672
rect 11041 8608 11059 8672
rect 11123 8608 11141 8672
rect 11205 8608 11223 8672
rect 11287 8608 11305 8672
rect 11369 8608 11387 8672
rect 11451 8608 11468 8672
rect 11532 8608 11549 8672
rect 11613 8608 11630 8672
rect 11694 8608 11711 8672
rect 11775 8608 11792 8672
rect 11856 8608 11873 8672
rect 11937 8608 11954 8672
rect 12018 8608 12035 8672
rect 12099 8608 12116 8672
rect 12180 8608 12197 8672
rect 12261 8608 12278 8672
rect 12342 8608 12359 8672
rect 12423 8608 12440 8672
rect 12504 8608 12521 8672
rect 12585 8608 12602 8672
rect 12666 8608 12683 8672
rect 12747 8608 12764 8672
rect 12828 8608 12845 8672
rect 12909 8608 12926 8672
rect 12990 8608 13007 8672
rect 13071 8608 13088 8672
rect 13152 8608 13169 8672
rect 13233 8608 13250 8672
rect 13314 8608 13331 8672
rect 13395 8608 13412 8672
rect 13476 8608 13493 8672
rect 13557 8608 13574 8672
rect 13638 8608 13655 8672
rect 13719 8608 13736 8672
rect 13800 8608 13817 8672
rect 13881 8608 13898 8672
rect 13962 8608 13979 8672
rect 14043 8608 14060 8672
rect 14124 8608 14141 8672
rect 14205 8608 14222 8672
rect 14286 8608 14303 8672
rect 14367 8608 14384 8672
rect 14448 8608 14465 8672
rect 14529 8608 14546 8672
rect 14610 8608 14627 8672
rect 14691 8608 14708 8672
rect 14772 8608 14789 8672
rect 14853 8608 14870 8672
rect 14934 8608 14940 8672
rect 10151 8586 14940 8608
rect 10151 8522 10157 8586
rect 10221 8522 10239 8586
rect 10303 8522 10321 8586
rect 10385 8522 10403 8586
rect 10467 8522 10485 8586
rect 10549 8522 10567 8586
rect 10631 8522 10649 8586
rect 10713 8522 10731 8586
rect 10795 8522 10813 8586
rect 10877 8522 10895 8586
rect 10959 8522 10977 8586
rect 11041 8522 11059 8586
rect 11123 8522 11141 8586
rect 11205 8522 11223 8586
rect 11287 8522 11305 8586
rect 11369 8522 11387 8586
rect 11451 8522 11468 8586
rect 11532 8522 11549 8586
rect 11613 8522 11630 8586
rect 11694 8522 11711 8586
rect 11775 8522 11792 8586
rect 11856 8522 11873 8586
rect 11937 8522 11954 8586
rect 12018 8522 12035 8586
rect 12099 8522 12116 8586
rect 12180 8522 12197 8586
rect 12261 8522 12278 8586
rect 12342 8522 12359 8586
rect 12423 8522 12440 8586
rect 12504 8522 12521 8586
rect 12585 8522 12602 8586
rect 12666 8522 12683 8586
rect 12747 8522 12764 8586
rect 12828 8522 12845 8586
rect 12909 8522 12926 8586
rect 12990 8522 13007 8586
rect 13071 8522 13088 8586
rect 13152 8522 13169 8586
rect 13233 8522 13250 8586
rect 13314 8522 13331 8586
rect 13395 8522 13412 8586
rect 13476 8522 13493 8586
rect 13557 8522 13574 8586
rect 13638 8522 13655 8586
rect 13719 8522 13736 8586
rect 13800 8522 13817 8586
rect 13881 8522 13898 8586
rect 13962 8522 13979 8586
rect 14043 8522 14060 8586
rect 14124 8522 14141 8586
rect 14205 8522 14222 8586
rect 14286 8522 14303 8586
rect 14367 8522 14384 8586
rect 14448 8522 14465 8586
rect 14529 8522 14546 8586
rect 14610 8522 14627 8586
rect 14691 8522 14708 8586
rect 14772 8522 14789 8586
rect 14853 8522 14870 8586
rect 14934 8522 14940 8586
rect 10151 8500 14940 8522
rect 10151 8436 10157 8500
rect 10221 8436 10239 8500
rect 10303 8436 10321 8500
rect 10385 8436 10403 8500
rect 10467 8436 10485 8500
rect 10549 8436 10567 8500
rect 10631 8436 10649 8500
rect 10713 8436 10731 8500
rect 10795 8436 10813 8500
rect 10877 8436 10895 8500
rect 10959 8436 10977 8500
rect 11041 8436 11059 8500
rect 11123 8436 11141 8500
rect 11205 8436 11223 8500
rect 11287 8436 11305 8500
rect 11369 8436 11387 8500
rect 11451 8436 11468 8500
rect 11532 8436 11549 8500
rect 11613 8436 11630 8500
rect 11694 8436 11711 8500
rect 11775 8436 11792 8500
rect 11856 8436 11873 8500
rect 11937 8436 11954 8500
rect 12018 8436 12035 8500
rect 12099 8436 12116 8500
rect 12180 8436 12197 8500
rect 12261 8436 12278 8500
rect 12342 8436 12359 8500
rect 12423 8436 12440 8500
rect 12504 8436 12521 8500
rect 12585 8436 12602 8500
rect 12666 8436 12683 8500
rect 12747 8436 12764 8500
rect 12828 8436 12845 8500
rect 12909 8436 12926 8500
rect 12990 8436 13007 8500
rect 13071 8436 13088 8500
rect 13152 8436 13169 8500
rect 13233 8436 13250 8500
rect 13314 8436 13331 8500
rect 13395 8436 13412 8500
rect 13476 8436 13493 8500
rect 13557 8436 13574 8500
rect 13638 8436 13655 8500
rect 13719 8436 13736 8500
rect 13800 8436 13817 8500
rect 13881 8436 13898 8500
rect 13962 8436 13979 8500
rect 14043 8436 14060 8500
rect 14124 8436 14141 8500
rect 14205 8436 14222 8500
rect 14286 8436 14303 8500
rect 14367 8436 14384 8500
rect 14448 8436 14465 8500
rect 14529 8436 14546 8500
rect 14610 8436 14627 8500
rect 14691 8436 14708 8500
rect 14772 8436 14789 8500
rect 14853 8436 14870 8500
rect 14934 8436 14940 8500
rect 10151 8414 14940 8436
rect 10151 8350 10157 8414
rect 10221 8350 10239 8414
rect 10303 8350 10321 8414
rect 10385 8350 10403 8414
rect 10467 8350 10485 8414
rect 10549 8350 10567 8414
rect 10631 8350 10649 8414
rect 10713 8350 10731 8414
rect 10795 8350 10813 8414
rect 10877 8350 10895 8414
rect 10959 8350 10977 8414
rect 11041 8350 11059 8414
rect 11123 8350 11141 8414
rect 11205 8350 11223 8414
rect 11287 8350 11305 8414
rect 11369 8350 11387 8414
rect 11451 8350 11468 8414
rect 11532 8350 11549 8414
rect 11613 8350 11630 8414
rect 11694 8350 11711 8414
rect 11775 8350 11792 8414
rect 11856 8350 11873 8414
rect 11937 8350 11954 8414
rect 12018 8350 12035 8414
rect 12099 8350 12116 8414
rect 12180 8350 12197 8414
rect 12261 8350 12278 8414
rect 12342 8350 12359 8414
rect 12423 8350 12440 8414
rect 12504 8350 12521 8414
rect 12585 8350 12602 8414
rect 12666 8350 12683 8414
rect 12747 8350 12764 8414
rect 12828 8350 12845 8414
rect 12909 8350 12926 8414
rect 12990 8350 13007 8414
rect 13071 8350 13088 8414
rect 13152 8350 13169 8414
rect 13233 8350 13250 8414
rect 13314 8350 13331 8414
rect 13395 8350 13412 8414
rect 13476 8350 13493 8414
rect 13557 8350 13574 8414
rect 13638 8350 13655 8414
rect 13719 8350 13736 8414
rect 13800 8350 13817 8414
rect 13881 8350 13898 8414
rect 13962 8350 13979 8414
rect 14043 8350 14060 8414
rect 14124 8350 14141 8414
rect 14205 8350 14222 8414
rect 14286 8350 14303 8414
rect 14367 8350 14384 8414
rect 14448 8350 14465 8414
rect 14529 8350 14546 8414
rect 14610 8350 14627 8414
rect 14691 8350 14708 8414
rect 14772 8350 14789 8414
rect 14853 8350 14870 8414
rect 14934 8350 14940 8414
rect 10151 8328 14940 8350
rect 10151 8264 10157 8328
rect 10221 8264 10239 8328
rect 10303 8264 10321 8328
rect 10385 8264 10403 8328
rect 10467 8264 10485 8328
rect 10549 8264 10567 8328
rect 10631 8264 10649 8328
rect 10713 8264 10731 8328
rect 10795 8264 10813 8328
rect 10877 8264 10895 8328
rect 10959 8264 10977 8328
rect 11041 8264 11059 8328
rect 11123 8264 11141 8328
rect 11205 8264 11223 8328
rect 11287 8264 11305 8328
rect 11369 8264 11387 8328
rect 11451 8264 11468 8328
rect 11532 8264 11549 8328
rect 11613 8264 11630 8328
rect 11694 8264 11711 8328
rect 11775 8264 11792 8328
rect 11856 8264 11873 8328
rect 11937 8264 11954 8328
rect 12018 8264 12035 8328
rect 12099 8264 12116 8328
rect 12180 8264 12197 8328
rect 12261 8264 12278 8328
rect 12342 8264 12359 8328
rect 12423 8264 12440 8328
rect 12504 8264 12521 8328
rect 12585 8264 12602 8328
rect 12666 8264 12683 8328
rect 12747 8264 12764 8328
rect 12828 8264 12845 8328
rect 12909 8264 12926 8328
rect 12990 8264 13007 8328
rect 13071 8264 13088 8328
rect 13152 8264 13169 8328
rect 13233 8264 13250 8328
rect 13314 8264 13331 8328
rect 13395 8264 13412 8328
rect 13476 8264 13493 8328
rect 13557 8264 13574 8328
rect 13638 8264 13655 8328
rect 13719 8264 13736 8328
rect 13800 8264 13817 8328
rect 13881 8264 13898 8328
rect 13962 8264 13979 8328
rect 14043 8264 14060 8328
rect 14124 8264 14141 8328
rect 14205 8264 14222 8328
rect 14286 8264 14303 8328
rect 14367 8264 14384 8328
rect 14448 8264 14465 8328
rect 14529 8264 14546 8328
rect 14610 8264 14627 8328
rect 14691 8264 14708 8328
rect 14772 8264 14789 8328
rect 14853 8264 14870 8328
rect 14934 8264 14940 8328
rect 10151 8242 14940 8264
rect 10151 8178 10157 8242
rect 10221 8178 10239 8242
rect 10303 8178 10321 8242
rect 10385 8178 10403 8242
rect 10467 8178 10485 8242
rect 10549 8178 10567 8242
rect 10631 8178 10649 8242
rect 10713 8178 10731 8242
rect 10795 8178 10813 8242
rect 10877 8178 10895 8242
rect 10959 8178 10977 8242
rect 11041 8178 11059 8242
rect 11123 8178 11141 8242
rect 11205 8178 11223 8242
rect 11287 8178 11305 8242
rect 11369 8178 11387 8242
rect 11451 8178 11468 8242
rect 11532 8178 11549 8242
rect 11613 8178 11630 8242
rect 11694 8178 11711 8242
rect 11775 8178 11792 8242
rect 11856 8178 11873 8242
rect 11937 8178 11954 8242
rect 12018 8178 12035 8242
rect 12099 8178 12116 8242
rect 12180 8178 12197 8242
rect 12261 8178 12278 8242
rect 12342 8178 12359 8242
rect 12423 8178 12440 8242
rect 12504 8178 12521 8242
rect 12585 8178 12602 8242
rect 12666 8178 12683 8242
rect 12747 8178 12764 8242
rect 12828 8178 12845 8242
rect 12909 8178 12926 8242
rect 12990 8178 13007 8242
rect 13071 8178 13088 8242
rect 13152 8178 13169 8242
rect 13233 8178 13250 8242
rect 13314 8178 13331 8242
rect 13395 8178 13412 8242
rect 13476 8178 13493 8242
rect 13557 8178 13574 8242
rect 13638 8178 13655 8242
rect 13719 8178 13736 8242
rect 13800 8178 13817 8242
rect 13881 8178 13898 8242
rect 13962 8178 13979 8242
rect 14043 8178 14060 8242
rect 14124 8178 14141 8242
rect 14205 8178 14222 8242
rect 14286 8178 14303 8242
rect 14367 8178 14384 8242
rect 14448 8178 14465 8242
rect 14529 8178 14546 8242
rect 14610 8178 14627 8242
rect 14691 8178 14708 8242
rect 14772 8178 14789 8242
rect 14853 8178 14870 8242
rect 14934 8178 14940 8242
rect 10151 8156 14940 8178
rect 10151 8092 10157 8156
rect 10221 8092 10239 8156
rect 10303 8092 10321 8156
rect 10385 8092 10403 8156
rect 10467 8092 10485 8156
rect 10549 8092 10567 8156
rect 10631 8092 10649 8156
rect 10713 8092 10731 8156
rect 10795 8092 10813 8156
rect 10877 8092 10895 8156
rect 10959 8092 10977 8156
rect 11041 8092 11059 8156
rect 11123 8092 11141 8156
rect 11205 8092 11223 8156
rect 11287 8092 11305 8156
rect 11369 8092 11387 8156
rect 11451 8092 11468 8156
rect 11532 8092 11549 8156
rect 11613 8092 11630 8156
rect 11694 8092 11711 8156
rect 11775 8092 11792 8156
rect 11856 8092 11873 8156
rect 11937 8092 11954 8156
rect 12018 8092 12035 8156
rect 12099 8092 12116 8156
rect 12180 8092 12197 8156
rect 12261 8092 12278 8156
rect 12342 8092 12359 8156
rect 12423 8092 12440 8156
rect 12504 8092 12521 8156
rect 12585 8092 12602 8156
rect 12666 8092 12683 8156
rect 12747 8092 12764 8156
rect 12828 8092 12845 8156
rect 12909 8092 12926 8156
rect 12990 8092 13007 8156
rect 13071 8092 13088 8156
rect 13152 8092 13169 8156
rect 13233 8092 13250 8156
rect 13314 8092 13331 8156
rect 13395 8092 13412 8156
rect 13476 8092 13493 8156
rect 13557 8092 13574 8156
rect 13638 8092 13655 8156
rect 13719 8092 13736 8156
rect 13800 8092 13817 8156
rect 13881 8092 13898 8156
rect 13962 8092 13979 8156
rect 14043 8092 14060 8156
rect 14124 8092 14141 8156
rect 14205 8092 14222 8156
rect 14286 8092 14303 8156
rect 14367 8092 14384 8156
rect 14448 8092 14465 8156
rect 14529 8092 14546 8156
rect 14610 8092 14627 8156
rect 14691 8092 14708 8156
rect 14772 8092 14789 8156
rect 14853 8092 14870 8156
rect 14934 8092 14940 8156
rect 10151 8070 14940 8092
rect 10151 8006 10157 8070
rect 10221 8006 10239 8070
rect 10303 8006 10321 8070
rect 10385 8006 10403 8070
rect 10467 8006 10485 8070
rect 10549 8006 10567 8070
rect 10631 8006 10649 8070
rect 10713 8006 10731 8070
rect 10795 8006 10813 8070
rect 10877 8006 10895 8070
rect 10959 8006 10977 8070
rect 11041 8006 11059 8070
rect 11123 8006 11141 8070
rect 11205 8006 11223 8070
rect 11287 8006 11305 8070
rect 11369 8006 11387 8070
rect 11451 8006 11468 8070
rect 11532 8006 11549 8070
rect 11613 8006 11630 8070
rect 11694 8006 11711 8070
rect 11775 8006 11792 8070
rect 11856 8006 11873 8070
rect 11937 8006 11954 8070
rect 12018 8006 12035 8070
rect 12099 8006 12116 8070
rect 12180 8006 12197 8070
rect 12261 8006 12278 8070
rect 12342 8006 12359 8070
rect 12423 8006 12440 8070
rect 12504 8006 12521 8070
rect 12585 8006 12602 8070
rect 12666 8006 12683 8070
rect 12747 8006 12764 8070
rect 12828 8006 12845 8070
rect 12909 8006 12926 8070
rect 12990 8006 13007 8070
rect 13071 8006 13088 8070
rect 13152 8006 13169 8070
rect 13233 8006 13250 8070
rect 13314 8006 13331 8070
rect 13395 8006 13412 8070
rect 13476 8006 13493 8070
rect 13557 8006 13574 8070
rect 13638 8006 13655 8070
rect 13719 8006 13736 8070
rect 13800 8006 13817 8070
rect 13881 8006 13898 8070
rect 13962 8006 13979 8070
rect 14043 8006 14060 8070
rect 14124 8006 14141 8070
rect 14205 8006 14222 8070
rect 14286 8006 14303 8070
rect 14367 8006 14384 8070
rect 14448 8006 14465 8070
rect 14529 8006 14546 8070
rect 14610 8006 14627 8070
rect 14691 8006 14708 8070
rect 14772 8006 14789 8070
rect 14853 8006 14870 8070
rect 14934 8006 14940 8070
rect 10151 7984 14940 8006
rect 10151 7920 10157 7984
rect 10221 7920 10239 7984
rect 10303 7920 10321 7984
rect 10385 7920 10403 7984
rect 10467 7920 10485 7984
rect 10549 7920 10567 7984
rect 10631 7920 10649 7984
rect 10713 7920 10731 7984
rect 10795 7920 10813 7984
rect 10877 7920 10895 7984
rect 10959 7920 10977 7984
rect 11041 7920 11059 7984
rect 11123 7920 11141 7984
rect 11205 7920 11223 7984
rect 11287 7920 11305 7984
rect 11369 7920 11387 7984
rect 11451 7920 11468 7984
rect 11532 7920 11549 7984
rect 11613 7920 11630 7984
rect 11694 7920 11711 7984
rect 11775 7920 11792 7984
rect 11856 7920 11873 7984
rect 11937 7920 11954 7984
rect 12018 7920 12035 7984
rect 12099 7920 12116 7984
rect 12180 7920 12197 7984
rect 12261 7920 12278 7984
rect 12342 7920 12359 7984
rect 12423 7920 12440 7984
rect 12504 7920 12521 7984
rect 12585 7920 12602 7984
rect 12666 7920 12683 7984
rect 12747 7920 12764 7984
rect 12828 7920 12845 7984
rect 12909 7920 12926 7984
rect 12990 7920 13007 7984
rect 13071 7920 13088 7984
rect 13152 7920 13169 7984
rect 13233 7920 13250 7984
rect 13314 7920 13331 7984
rect 13395 7920 13412 7984
rect 13476 7920 13493 7984
rect 13557 7920 13574 7984
rect 13638 7920 13655 7984
rect 13719 7920 13736 7984
rect 13800 7920 13817 7984
rect 13881 7920 13898 7984
rect 13962 7920 13979 7984
rect 14043 7920 14060 7984
rect 14124 7920 14141 7984
rect 14205 7920 14222 7984
rect 14286 7920 14303 7984
rect 14367 7920 14384 7984
rect 14448 7920 14465 7984
rect 14529 7920 14546 7984
rect 14610 7920 14627 7984
rect 14691 7920 14708 7984
rect 14772 7920 14789 7984
rect 14853 7920 14870 7984
rect 14934 7920 14940 7984
rect 10151 7918 14940 7920
<< via3 >>
rect 106 8780 170 8844
rect 187 8780 251 8844
rect 268 8780 332 8844
rect 349 8780 413 8844
rect 430 8780 494 8844
rect 510 8780 574 8844
rect 590 8780 654 8844
rect 670 8780 734 8844
rect 750 8780 814 8844
rect 830 8780 894 8844
rect 910 8780 974 8844
rect 990 8780 1054 8844
rect 1070 8780 1134 8844
rect 1150 8780 1214 8844
rect 1230 8780 1294 8844
rect 1310 8780 1374 8844
rect 1390 8780 1454 8844
rect 1470 8780 1534 8844
rect 1550 8780 1614 8844
rect 1630 8780 1694 8844
rect 1710 8780 1774 8844
rect 1790 8780 1854 8844
rect 1870 8780 1934 8844
rect 1950 8780 2014 8844
rect 2030 8780 2094 8844
rect 2110 8780 2174 8844
rect 2190 8780 2254 8844
rect 2270 8780 2334 8844
rect 2350 8780 2414 8844
rect 2430 8780 2494 8844
rect 2510 8780 2574 8844
rect 2590 8780 2654 8844
rect 2670 8780 2734 8844
rect 2750 8780 2814 8844
rect 2830 8780 2894 8844
rect 2910 8780 2974 8844
rect 2990 8780 3054 8844
rect 3070 8780 3134 8844
rect 3150 8780 3214 8844
rect 3230 8780 3294 8844
rect 3310 8780 3374 8844
rect 3390 8780 3454 8844
rect 3470 8780 3534 8844
rect 3550 8780 3614 8844
rect 3630 8780 3694 8844
rect 3710 8780 3774 8844
rect 3790 8780 3854 8844
rect 3870 8780 3934 8844
rect 3950 8780 4014 8844
rect 4030 8780 4094 8844
rect 4110 8780 4174 8844
rect 4190 8780 4254 8844
rect 4270 8780 4334 8844
rect 4350 8780 4414 8844
rect 4430 8780 4494 8844
rect 4510 8780 4574 8844
rect 4590 8780 4654 8844
rect 4670 8780 4734 8844
rect 4750 8780 4814 8844
rect 4830 8780 4894 8844
rect 106 8694 170 8758
rect 187 8694 251 8758
rect 268 8694 332 8758
rect 349 8694 413 8758
rect 430 8694 494 8758
rect 510 8694 574 8758
rect 590 8694 654 8758
rect 670 8694 734 8758
rect 750 8694 814 8758
rect 830 8694 894 8758
rect 910 8694 974 8758
rect 990 8694 1054 8758
rect 1070 8694 1134 8758
rect 1150 8694 1214 8758
rect 1230 8694 1294 8758
rect 1310 8694 1374 8758
rect 1390 8694 1454 8758
rect 1470 8694 1534 8758
rect 1550 8694 1614 8758
rect 1630 8694 1694 8758
rect 1710 8694 1774 8758
rect 1790 8694 1854 8758
rect 1870 8694 1934 8758
rect 1950 8694 2014 8758
rect 2030 8694 2094 8758
rect 2110 8694 2174 8758
rect 2190 8694 2254 8758
rect 2270 8694 2334 8758
rect 2350 8694 2414 8758
rect 2430 8694 2494 8758
rect 2510 8694 2574 8758
rect 2590 8694 2654 8758
rect 2670 8694 2734 8758
rect 2750 8694 2814 8758
rect 2830 8694 2894 8758
rect 2910 8694 2974 8758
rect 2990 8694 3054 8758
rect 3070 8694 3134 8758
rect 3150 8694 3214 8758
rect 3230 8694 3294 8758
rect 3310 8694 3374 8758
rect 3390 8694 3454 8758
rect 3470 8694 3534 8758
rect 3550 8694 3614 8758
rect 3630 8694 3694 8758
rect 3710 8694 3774 8758
rect 3790 8694 3854 8758
rect 3870 8694 3934 8758
rect 3950 8694 4014 8758
rect 4030 8694 4094 8758
rect 4110 8694 4174 8758
rect 4190 8694 4254 8758
rect 4270 8694 4334 8758
rect 4350 8694 4414 8758
rect 4430 8694 4494 8758
rect 4510 8694 4574 8758
rect 4590 8694 4654 8758
rect 4670 8694 4734 8758
rect 4750 8694 4814 8758
rect 4830 8694 4894 8758
rect 106 8608 170 8672
rect 187 8608 251 8672
rect 268 8608 332 8672
rect 349 8608 413 8672
rect 430 8608 494 8672
rect 510 8608 574 8672
rect 590 8608 654 8672
rect 670 8608 734 8672
rect 750 8608 814 8672
rect 830 8608 894 8672
rect 910 8608 974 8672
rect 990 8608 1054 8672
rect 1070 8608 1134 8672
rect 1150 8608 1214 8672
rect 1230 8608 1294 8672
rect 1310 8608 1374 8672
rect 1390 8608 1454 8672
rect 1470 8608 1534 8672
rect 1550 8608 1614 8672
rect 1630 8608 1694 8672
rect 1710 8608 1774 8672
rect 1790 8608 1854 8672
rect 1870 8608 1934 8672
rect 1950 8608 2014 8672
rect 2030 8608 2094 8672
rect 2110 8608 2174 8672
rect 2190 8608 2254 8672
rect 2270 8608 2334 8672
rect 2350 8608 2414 8672
rect 2430 8608 2494 8672
rect 2510 8608 2574 8672
rect 2590 8608 2654 8672
rect 2670 8608 2734 8672
rect 2750 8608 2814 8672
rect 2830 8608 2894 8672
rect 2910 8608 2974 8672
rect 2990 8608 3054 8672
rect 3070 8608 3134 8672
rect 3150 8608 3214 8672
rect 3230 8608 3294 8672
rect 3310 8608 3374 8672
rect 3390 8608 3454 8672
rect 3470 8608 3534 8672
rect 3550 8608 3614 8672
rect 3630 8608 3694 8672
rect 3710 8608 3774 8672
rect 3790 8608 3854 8672
rect 3870 8608 3934 8672
rect 3950 8608 4014 8672
rect 4030 8608 4094 8672
rect 4110 8608 4174 8672
rect 4190 8608 4254 8672
rect 4270 8608 4334 8672
rect 4350 8608 4414 8672
rect 4430 8608 4494 8672
rect 4510 8608 4574 8672
rect 4590 8608 4654 8672
rect 4670 8608 4734 8672
rect 4750 8608 4814 8672
rect 4830 8608 4894 8672
rect 106 8522 170 8586
rect 187 8522 251 8586
rect 268 8522 332 8586
rect 349 8522 413 8586
rect 430 8522 494 8586
rect 510 8522 574 8586
rect 590 8522 654 8586
rect 670 8522 734 8586
rect 750 8522 814 8586
rect 830 8522 894 8586
rect 910 8522 974 8586
rect 990 8522 1054 8586
rect 1070 8522 1134 8586
rect 1150 8522 1214 8586
rect 1230 8522 1294 8586
rect 1310 8522 1374 8586
rect 1390 8522 1454 8586
rect 1470 8522 1534 8586
rect 1550 8522 1614 8586
rect 1630 8522 1694 8586
rect 1710 8522 1774 8586
rect 1790 8522 1854 8586
rect 1870 8522 1934 8586
rect 1950 8522 2014 8586
rect 2030 8522 2094 8586
rect 2110 8522 2174 8586
rect 2190 8522 2254 8586
rect 2270 8522 2334 8586
rect 2350 8522 2414 8586
rect 2430 8522 2494 8586
rect 2510 8522 2574 8586
rect 2590 8522 2654 8586
rect 2670 8522 2734 8586
rect 2750 8522 2814 8586
rect 2830 8522 2894 8586
rect 2910 8522 2974 8586
rect 2990 8522 3054 8586
rect 3070 8522 3134 8586
rect 3150 8522 3214 8586
rect 3230 8522 3294 8586
rect 3310 8522 3374 8586
rect 3390 8522 3454 8586
rect 3470 8522 3534 8586
rect 3550 8522 3614 8586
rect 3630 8522 3694 8586
rect 3710 8522 3774 8586
rect 3790 8522 3854 8586
rect 3870 8522 3934 8586
rect 3950 8522 4014 8586
rect 4030 8522 4094 8586
rect 4110 8522 4174 8586
rect 4190 8522 4254 8586
rect 4270 8522 4334 8586
rect 4350 8522 4414 8586
rect 4430 8522 4494 8586
rect 4510 8522 4574 8586
rect 4590 8522 4654 8586
rect 4670 8522 4734 8586
rect 4750 8522 4814 8586
rect 4830 8522 4894 8586
rect 106 8436 170 8500
rect 187 8436 251 8500
rect 268 8436 332 8500
rect 349 8436 413 8500
rect 430 8436 494 8500
rect 510 8436 574 8500
rect 590 8436 654 8500
rect 670 8436 734 8500
rect 750 8436 814 8500
rect 830 8436 894 8500
rect 910 8436 974 8500
rect 990 8436 1054 8500
rect 1070 8436 1134 8500
rect 1150 8436 1214 8500
rect 1230 8436 1294 8500
rect 1310 8436 1374 8500
rect 1390 8436 1454 8500
rect 1470 8436 1534 8500
rect 1550 8436 1614 8500
rect 1630 8436 1694 8500
rect 1710 8436 1774 8500
rect 1790 8436 1854 8500
rect 1870 8436 1934 8500
rect 1950 8436 2014 8500
rect 2030 8436 2094 8500
rect 2110 8436 2174 8500
rect 2190 8436 2254 8500
rect 2270 8436 2334 8500
rect 2350 8436 2414 8500
rect 2430 8436 2494 8500
rect 2510 8436 2574 8500
rect 2590 8436 2654 8500
rect 2670 8436 2734 8500
rect 2750 8436 2814 8500
rect 2830 8436 2894 8500
rect 2910 8436 2974 8500
rect 2990 8436 3054 8500
rect 3070 8436 3134 8500
rect 3150 8436 3214 8500
rect 3230 8436 3294 8500
rect 3310 8436 3374 8500
rect 3390 8436 3454 8500
rect 3470 8436 3534 8500
rect 3550 8436 3614 8500
rect 3630 8436 3694 8500
rect 3710 8436 3774 8500
rect 3790 8436 3854 8500
rect 3870 8436 3934 8500
rect 3950 8436 4014 8500
rect 4030 8436 4094 8500
rect 4110 8436 4174 8500
rect 4190 8436 4254 8500
rect 4270 8436 4334 8500
rect 4350 8436 4414 8500
rect 4430 8436 4494 8500
rect 4510 8436 4574 8500
rect 4590 8436 4654 8500
rect 4670 8436 4734 8500
rect 4750 8436 4814 8500
rect 4830 8436 4894 8500
rect 106 8350 170 8414
rect 187 8350 251 8414
rect 268 8350 332 8414
rect 349 8350 413 8414
rect 430 8350 494 8414
rect 510 8350 574 8414
rect 590 8350 654 8414
rect 670 8350 734 8414
rect 750 8350 814 8414
rect 830 8350 894 8414
rect 910 8350 974 8414
rect 990 8350 1054 8414
rect 1070 8350 1134 8414
rect 1150 8350 1214 8414
rect 1230 8350 1294 8414
rect 1310 8350 1374 8414
rect 1390 8350 1454 8414
rect 1470 8350 1534 8414
rect 1550 8350 1614 8414
rect 1630 8350 1694 8414
rect 1710 8350 1774 8414
rect 1790 8350 1854 8414
rect 1870 8350 1934 8414
rect 1950 8350 2014 8414
rect 2030 8350 2094 8414
rect 2110 8350 2174 8414
rect 2190 8350 2254 8414
rect 2270 8350 2334 8414
rect 2350 8350 2414 8414
rect 2430 8350 2494 8414
rect 2510 8350 2574 8414
rect 2590 8350 2654 8414
rect 2670 8350 2734 8414
rect 2750 8350 2814 8414
rect 2830 8350 2894 8414
rect 2910 8350 2974 8414
rect 2990 8350 3054 8414
rect 3070 8350 3134 8414
rect 3150 8350 3214 8414
rect 3230 8350 3294 8414
rect 3310 8350 3374 8414
rect 3390 8350 3454 8414
rect 3470 8350 3534 8414
rect 3550 8350 3614 8414
rect 3630 8350 3694 8414
rect 3710 8350 3774 8414
rect 3790 8350 3854 8414
rect 3870 8350 3934 8414
rect 3950 8350 4014 8414
rect 4030 8350 4094 8414
rect 4110 8350 4174 8414
rect 4190 8350 4254 8414
rect 4270 8350 4334 8414
rect 4350 8350 4414 8414
rect 4430 8350 4494 8414
rect 4510 8350 4574 8414
rect 4590 8350 4654 8414
rect 4670 8350 4734 8414
rect 4750 8350 4814 8414
rect 4830 8350 4894 8414
rect 106 8264 170 8328
rect 187 8264 251 8328
rect 268 8264 332 8328
rect 349 8264 413 8328
rect 430 8264 494 8328
rect 510 8264 574 8328
rect 590 8264 654 8328
rect 670 8264 734 8328
rect 750 8264 814 8328
rect 830 8264 894 8328
rect 910 8264 974 8328
rect 990 8264 1054 8328
rect 1070 8264 1134 8328
rect 1150 8264 1214 8328
rect 1230 8264 1294 8328
rect 1310 8264 1374 8328
rect 1390 8264 1454 8328
rect 1470 8264 1534 8328
rect 1550 8264 1614 8328
rect 1630 8264 1694 8328
rect 1710 8264 1774 8328
rect 1790 8264 1854 8328
rect 1870 8264 1934 8328
rect 1950 8264 2014 8328
rect 2030 8264 2094 8328
rect 2110 8264 2174 8328
rect 2190 8264 2254 8328
rect 2270 8264 2334 8328
rect 2350 8264 2414 8328
rect 2430 8264 2494 8328
rect 2510 8264 2574 8328
rect 2590 8264 2654 8328
rect 2670 8264 2734 8328
rect 2750 8264 2814 8328
rect 2830 8264 2894 8328
rect 2910 8264 2974 8328
rect 2990 8264 3054 8328
rect 3070 8264 3134 8328
rect 3150 8264 3214 8328
rect 3230 8264 3294 8328
rect 3310 8264 3374 8328
rect 3390 8264 3454 8328
rect 3470 8264 3534 8328
rect 3550 8264 3614 8328
rect 3630 8264 3694 8328
rect 3710 8264 3774 8328
rect 3790 8264 3854 8328
rect 3870 8264 3934 8328
rect 3950 8264 4014 8328
rect 4030 8264 4094 8328
rect 4110 8264 4174 8328
rect 4190 8264 4254 8328
rect 4270 8264 4334 8328
rect 4350 8264 4414 8328
rect 4430 8264 4494 8328
rect 4510 8264 4574 8328
rect 4590 8264 4654 8328
rect 4670 8264 4734 8328
rect 4750 8264 4814 8328
rect 4830 8264 4894 8328
rect 106 8178 170 8242
rect 187 8178 251 8242
rect 268 8178 332 8242
rect 349 8178 413 8242
rect 430 8178 494 8242
rect 510 8178 574 8242
rect 590 8178 654 8242
rect 670 8178 734 8242
rect 750 8178 814 8242
rect 830 8178 894 8242
rect 910 8178 974 8242
rect 990 8178 1054 8242
rect 1070 8178 1134 8242
rect 1150 8178 1214 8242
rect 1230 8178 1294 8242
rect 1310 8178 1374 8242
rect 1390 8178 1454 8242
rect 1470 8178 1534 8242
rect 1550 8178 1614 8242
rect 1630 8178 1694 8242
rect 1710 8178 1774 8242
rect 1790 8178 1854 8242
rect 1870 8178 1934 8242
rect 1950 8178 2014 8242
rect 2030 8178 2094 8242
rect 2110 8178 2174 8242
rect 2190 8178 2254 8242
rect 2270 8178 2334 8242
rect 2350 8178 2414 8242
rect 2430 8178 2494 8242
rect 2510 8178 2574 8242
rect 2590 8178 2654 8242
rect 2670 8178 2734 8242
rect 2750 8178 2814 8242
rect 2830 8178 2894 8242
rect 2910 8178 2974 8242
rect 2990 8178 3054 8242
rect 3070 8178 3134 8242
rect 3150 8178 3214 8242
rect 3230 8178 3294 8242
rect 3310 8178 3374 8242
rect 3390 8178 3454 8242
rect 3470 8178 3534 8242
rect 3550 8178 3614 8242
rect 3630 8178 3694 8242
rect 3710 8178 3774 8242
rect 3790 8178 3854 8242
rect 3870 8178 3934 8242
rect 3950 8178 4014 8242
rect 4030 8178 4094 8242
rect 4110 8178 4174 8242
rect 4190 8178 4254 8242
rect 4270 8178 4334 8242
rect 4350 8178 4414 8242
rect 4430 8178 4494 8242
rect 4510 8178 4574 8242
rect 4590 8178 4654 8242
rect 4670 8178 4734 8242
rect 4750 8178 4814 8242
rect 4830 8178 4894 8242
rect 106 8092 170 8156
rect 187 8092 251 8156
rect 268 8092 332 8156
rect 349 8092 413 8156
rect 430 8092 494 8156
rect 510 8092 574 8156
rect 590 8092 654 8156
rect 670 8092 734 8156
rect 750 8092 814 8156
rect 830 8092 894 8156
rect 910 8092 974 8156
rect 990 8092 1054 8156
rect 1070 8092 1134 8156
rect 1150 8092 1214 8156
rect 1230 8092 1294 8156
rect 1310 8092 1374 8156
rect 1390 8092 1454 8156
rect 1470 8092 1534 8156
rect 1550 8092 1614 8156
rect 1630 8092 1694 8156
rect 1710 8092 1774 8156
rect 1790 8092 1854 8156
rect 1870 8092 1934 8156
rect 1950 8092 2014 8156
rect 2030 8092 2094 8156
rect 2110 8092 2174 8156
rect 2190 8092 2254 8156
rect 2270 8092 2334 8156
rect 2350 8092 2414 8156
rect 2430 8092 2494 8156
rect 2510 8092 2574 8156
rect 2590 8092 2654 8156
rect 2670 8092 2734 8156
rect 2750 8092 2814 8156
rect 2830 8092 2894 8156
rect 2910 8092 2974 8156
rect 2990 8092 3054 8156
rect 3070 8092 3134 8156
rect 3150 8092 3214 8156
rect 3230 8092 3294 8156
rect 3310 8092 3374 8156
rect 3390 8092 3454 8156
rect 3470 8092 3534 8156
rect 3550 8092 3614 8156
rect 3630 8092 3694 8156
rect 3710 8092 3774 8156
rect 3790 8092 3854 8156
rect 3870 8092 3934 8156
rect 3950 8092 4014 8156
rect 4030 8092 4094 8156
rect 4110 8092 4174 8156
rect 4190 8092 4254 8156
rect 4270 8092 4334 8156
rect 4350 8092 4414 8156
rect 4430 8092 4494 8156
rect 4510 8092 4574 8156
rect 4590 8092 4654 8156
rect 4670 8092 4734 8156
rect 4750 8092 4814 8156
rect 4830 8092 4894 8156
rect 106 8006 170 8070
rect 187 8006 251 8070
rect 268 8006 332 8070
rect 349 8006 413 8070
rect 430 8006 494 8070
rect 510 8006 574 8070
rect 590 8006 654 8070
rect 670 8006 734 8070
rect 750 8006 814 8070
rect 830 8006 894 8070
rect 910 8006 974 8070
rect 990 8006 1054 8070
rect 1070 8006 1134 8070
rect 1150 8006 1214 8070
rect 1230 8006 1294 8070
rect 1310 8006 1374 8070
rect 1390 8006 1454 8070
rect 1470 8006 1534 8070
rect 1550 8006 1614 8070
rect 1630 8006 1694 8070
rect 1710 8006 1774 8070
rect 1790 8006 1854 8070
rect 1870 8006 1934 8070
rect 1950 8006 2014 8070
rect 2030 8006 2094 8070
rect 2110 8006 2174 8070
rect 2190 8006 2254 8070
rect 2270 8006 2334 8070
rect 2350 8006 2414 8070
rect 2430 8006 2494 8070
rect 2510 8006 2574 8070
rect 2590 8006 2654 8070
rect 2670 8006 2734 8070
rect 2750 8006 2814 8070
rect 2830 8006 2894 8070
rect 2910 8006 2974 8070
rect 2990 8006 3054 8070
rect 3070 8006 3134 8070
rect 3150 8006 3214 8070
rect 3230 8006 3294 8070
rect 3310 8006 3374 8070
rect 3390 8006 3454 8070
rect 3470 8006 3534 8070
rect 3550 8006 3614 8070
rect 3630 8006 3694 8070
rect 3710 8006 3774 8070
rect 3790 8006 3854 8070
rect 3870 8006 3934 8070
rect 3950 8006 4014 8070
rect 4030 8006 4094 8070
rect 4110 8006 4174 8070
rect 4190 8006 4254 8070
rect 4270 8006 4334 8070
rect 4350 8006 4414 8070
rect 4430 8006 4494 8070
rect 4510 8006 4574 8070
rect 4590 8006 4654 8070
rect 4670 8006 4734 8070
rect 4750 8006 4814 8070
rect 4830 8006 4894 8070
rect 106 7920 170 7984
rect 187 7920 251 7984
rect 268 7920 332 7984
rect 349 7920 413 7984
rect 430 7920 494 7984
rect 510 7920 574 7984
rect 590 7920 654 7984
rect 670 7920 734 7984
rect 750 7920 814 7984
rect 830 7920 894 7984
rect 910 7920 974 7984
rect 990 7920 1054 7984
rect 1070 7920 1134 7984
rect 1150 7920 1214 7984
rect 1230 7920 1294 7984
rect 1310 7920 1374 7984
rect 1390 7920 1454 7984
rect 1470 7920 1534 7984
rect 1550 7920 1614 7984
rect 1630 7920 1694 7984
rect 1710 7920 1774 7984
rect 1790 7920 1854 7984
rect 1870 7920 1934 7984
rect 1950 7920 2014 7984
rect 2030 7920 2094 7984
rect 2110 7920 2174 7984
rect 2190 7920 2254 7984
rect 2270 7920 2334 7984
rect 2350 7920 2414 7984
rect 2430 7920 2494 7984
rect 2510 7920 2574 7984
rect 2590 7920 2654 7984
rect 2670 7920 2734 7984
rect 2750 7920 2814 7984
rect 2830 7920 2894 7984
rect 2910 7920 2974 7984
rect 2990 7920 3054 7984
rect 3070 7920 3134 7984
rect 3150 7920 3214 7984
rect 3230 7920 3294 7984
rect 3310 7920 3374 7984
rect 3390 7920 3454 7984
rect 3470 7920 3534 7984
rect 3550 7920 3614 7984
rect 3630 7920 3694 7984
rect 3710 7920 3774 7984
rect 3790 7920 3854 7984
rect 3870 7920 3934 7984
rect 3950 7920 4014 7984
rect 4030 7920 4094 7984
rect 4110 7920 4174 7984
rect 4190 7920 4254 7984
rect 4270 7920 4334 7984
rect 4350 7920 4414 7984
rect 4430 7920 4494 7984
rect 4510 7920 4574 7984
rect 4590 7920 4654 7984
rect 4670 7920 4734 7984
rect 4750 7920 4814 7984
rect 4830 7920 4894 7984
rect 10157 8780 10221 8844
rect 10239 8780 10303 8844
rect 10321 8780 10385 8844
rect 10403 8780 10467 8844
rect 10485 8780 10549 8844
rect 10567 8780 10631 8844
rect 10649 8780 10713 8844
rect 10731 8780 10795 8844
rect 10813 8780 10877 8844
rect 10895 8780 10959 8844
rect 10977 8780 11041 8844
rect 11059 8780 11123 8844
rect 11141 8780 11205 8844
rect 11223 8780 11287 8844
rect 11305 8780 11369 8844
rect 11387 8780 11451 8844
rect 11468 8780 11532 8844
rect 11549 8780 11613 8844
rect 11630 8780 11694 8844
rect 11711 8780 11775 8844
rect 11792 8780 11856 8844
rect 11873 8780 11937 8844
rect 11954 8780 12018 8844
rect 12035 8780 12099 8844
rect 12116 8780 12180 8844
rect 12197 8780 12261 8844
rect 12278 8780 12342 8844
rect 12359 8780 12423 8844
rect 12440 8780 12504 8844
rect 12521 8780 12585 8844
rect 12602 8780 12666 8844
rect 12683 8780 12747 8844
rect 12764 8780 12828 8844
rect 12845 8780 12909 8844
rect 12926 8780 12990 8844
rect 13007 8780 13071 8844
rect 13088 8780 13152 8844
rect 13169 8780 13233 8844
rect 13250 8780 13314 8844
rect 13331 8780 13395 8844
rect 13412 8780 13476 8844
rect 13493 8780 13557 8844
rect 13574 8780 13638 8844
rect 13655 8780 13719 8844
rect 13736 8780 13800 8844
rect 13817 8780 13881 8844
rect 13898 8780 13962 8844
rect 13979 8780 14043 8844
rect 14060 8780 14124 8844
rect 14141 8780 14205 8844
rect 14222 8780 14286 8844
rect 14303 8780 14367 8844
rect 14384 8780 14448 8844
rect 14465 8780 14529 8844
rect 14546 8780 14610 8844
rect 14627 8780 14691 8844
rect 14708 8780 14772 8844
rect 14789 8780 14853 8844
rect 14870 8780 14934 8844
rect 10157 8694 10221 8758
rect 10239 8694 10303 8758
rect 10321 8694 10385 8758
rect 10403 8694 10467 8758
rect 10485 8694 10549 8758
rect 10567 8694 10631 8758
rect 10649 8694 10713 8758
rect 10731 8694 10795 8758
rect 10813 8694 10877 8758
rect 10895 8694 10959 8758
rect 10977 8694 11041 8758
rect 11059 8694 11123 8758
rect 11141 8694 11205 8758
rect 11223 8694 11287 8758
rect 11305 8694 11369 8758
rect 11387 8694 11451 8758
rect 11468 8694 11532 8758
rect 11549 8694 11613 8758
rect 11630 8694 11694 8758
rect 11711 8694 11775 8758
rect 11792 8694 11856 8758
rect 11873 8694 11937 8758
rect 11954 8694 12018 8758
rect 12035 8694 12099 8758
rect 12116 8694 12180 8758
rect 12197 8694 12261 8758
rect 12278 8694 12342 8758
rect 12359 8694 12423 8758
rect 12440 8694 12504 8758
rect 12521 8694 12585 8758
rect 12602 8694 12666 8758
rect 12683 8694 12747 8758
rect 12764 8694 12828 8758
rect 12845 8694 12909 8758
rect 12926 8694 12990 8758
rect 13007 8694 13071 8758
rect 13088 8694 13152 8758
rect 13169 8694 13233 8758
rect 13250 8694 13314 8758
rect 13331 8694 13395 8758
rect 13412 8694 13476 8758
rect 13493 8694 13557 8758
rect 13574 8694 13638 8758
rect 13655 8694 13719 8758
rect 13736 8694 13800 8758
rect 13817 8694 13881 8758
rect 13898 8694 13962 8758
rect 13979 8694 14043 8758
rect 14060 8694 14124 8758
rect 14141 8694 14205 8758
rect 14222 8694 14286 8758
rect 14303 8694 14367 8758
rect 14384 8694 14448 8758
rect 14465 8694 14529 8758
rect 14546 8694 14610 8758
rect 14627 8694 14691 8758
rect 14708 8694 14772 8758
rect 14789 8694 14853 8758
rect 14870 8694 14934 8758
rect 10157 8608 10221 8672
rect 10239 8608 10303 8672
rect 10321 8608 10385 8672
rect 10403 8608 10467 8672
rect 10485 8608 10549 8672
rect 10567 8608 10631 8672
rect 10649 8608 10713 8672
rect 10731 8608 10795 8672
rect 10813 8608 10877 8672
rect 10895 8608 10959 8672
rect 10977 8608 11041 8672
rect 11059 8608 11123 8672
rect 11141 8608 11205 8672
rect 11223 8608 11287 8672
rect 11305 8608 11369 8672
rect 11387 8608 11451 8672
rect 11468 8608 11532 8672
rect 11549 8608 11613 8672
rect 11630 8608 11694 8672
rect 11711 8608 11775 8672
rect 11792 8608 11856 8672
rect 11873 8608 11937 8672
rect 11954 8608 12018 8672
rect 12035 8608 12099 8672
rect 12116 8608 12180 8672
rect 12197 8608 12261 8672
rect 12278 8608 12342 8672
rect 12359 8608 12423 8672
rect 12440 8608 12504 8672
rect 12521 8608 12585 8672
rect 12602 8608 12666 8672
rect 12683 8608 12747 8672
rect 12764 8608 12828 8672
rect 12845 8608 12909 8672
rect 12926 8608 12990 8672
rect 13007 8608 13071 8672
rect 13088 8608 13152 8672
rect 13169 8608 13233 8672
rect 13250 8608 13314 8672
rect 13331 8608 13395 8672
rect 13412 8608 13476 8672
rect 13493 8608 13557 8672
rect 13574 8608 13638 8672
rect 13655 8608 13719 8672
rect 13736 8608 13800 8672
rect 13817 8608 13881 8672
rect 13898 8608 13962 8672
rect 13979 8608 14043 8672
rect 14060 8608 14124 8672
rect 14141 8608 14205 8672
rect 14222 8608 14286 8672
rect 14303 8608 14367 8672
rect 14384 8608 14448 8672
rect 14465 8608 14529 8672
rect 14546 8608 14610 8672
rect 14627 8608 14691 8672
rect 14708 8608 14772 8672
rect 14789 8608 14853 8672
rect 14870 8608 14934 8672
rect 10157 8522 10221 8586
rect 10239 8522 10303 8586
rect 10321 8522 10385 8586
rect 10403 8522 10467 8586
rect 10485 8522 10549 8586
rect 10567 8522 10631 8586
rect 10649 8522 10713 8586
rect 10731 8522 10795 8586
rect 10813 8522 10877 8586
rect 10895 8522 10959 8586
rect 10977 8522 11041 8586
rect 11059 8522 11123 8586
rect 11141 8522 11205 8586
rect 11223 8522 11287 8586
rect 11305 8522 11369 8586
rect 11387 8522 11451 8586
rect 11468 8522 11532 8586
rect 11549 8522 11613 8586
rect 11630 8522 11694 8586
rect 11711 8522 11775 8586
rect 11792 8522 11856 8586
rect 11873 8522 11937 8586
rect 11954 8522 12018 8586
rect 12035 8522 12099 8586
rect 12116 8522 12180 8586
rect 12197 8522 12261 8586
rect 12278 8522 12342 8586
rect 12359 8522 12423 8586
rect 12440 8522 12504 8586
rect 12521 8522 12585 8586
rect 12602 8522 12666 8586
rect 12683 8522 12747 8586
rect 12764 8522 12828 8586
rect 12845 8522 12909 8586
rect 12926 8522 12990 8586
rect 13007 8522 13071 8586
rect 13088 8522 13152 8586
rect 13169 8522 13233 8586
rect 13250 8522 13314 8586
rect 13331 8522 13395 8586
rect 13412 8522 13476 8586
rect 13493 8522 13557 8586
rect 13574 8522 13638 8586
rect 13655 8522 13719 8586
rect 13736 8522 13800 8586
rect 13817 8522 13881 8586
rect 13898 8522 13962 8586
rect 13979 8522 14043 8586
rect 14060 8522 14124 8586
rect 14141 8522 14205 8586
rect 14222 8522 14286 8586
rect 14303 8522 14367 8586
rect 14384 8522 14448 8586
rect 14465 8522 14529 8586
rect 14546 8522 14610 8586
rect 14627 8522 14691 8586
rect 14708 8522 14772 8586
rect 14789 8522 14853 8586
rect 14870 8522 14934 8586
rect 10157 8436 10221 8500
rect 10239 8436 10303 8500
rect 10321 8436 10385 8500
rect 10403 8436 10467 8500
rect 10485 8436 10549 8500
rect 10567 8436 10631 8500
rect 10649 8436 10713 8500
rect 10731 8436 10795 8500
rect 10813 8436 10877 8500
rect 10895 8436 10959 8500
rect 10977 8436 11041 8500
rect 11059 8436 11123 8500
rect 11141 8436 11205 8500
rect 11223 8436 11287 8500
rect 11305 8436 11369 8500
rect 11387 8436 11451 8500
rect 11468 8436 11532 8500
rect 11549 8436 11613 8500
rect 11630 8436 11694 8500
rect 11711 8436 11775 8500
rect 11792 8436 11856 8500
rect 11873 8436 11937 8500
rect 11954 8436 12018 8500
rect 12035 8436 12099 8500
rect 12116 8436 12180 8500
rect 12197 8436 12261 8500
rect 12278 8436 12342 8500
rect 12359 8436 12423 8500
rect 12440 8436 12504 8500
rect 12521 8436 12585 8500
rect 12602 8436 12666 8500
rect 12683 8436 12747 8500
rect 12764 8436 12828 8500
rect 12845 8436 12909 8500
rect 12926 8436 12990 8500
rect 13007 8436 13071 8500
rect 13088 8436 13152 8500
rect 13169 8436 13233 8500
rect 13250 8436 13314 8500
rect 13331 8436 13395 8500
rect 13412 8436 13476 8500
rect 13493 8436 13557 8500
rect 13574 8436 13638 8500
rect 13655 8436 13719 8500
rect 13736 8436 13800 8500
rect 13817 8436 13881 8500
rect 13898 8436 13962 8500
rect 13979 8436 14043 8500
rect 14060 8436 14124 8500
rect 14141 8436 14205 8500
rect 14222 8436 14286 8500
rect 14303 8436 14367 8500
rect 14384 8436 14448 8500
rect 14465 8436 14529 8500
rect 14546 8436 14610 8500
rect 14627 8436 14691 8500
rect 14708 8436 14772 8500
rect 14789 8436 14853 8500
rect 14870 8436 14934 8500
rect 10157 8350 10221 8414
rect 10239 8350 10303 8414
rect 10321 8350 10385 8414
rect 10403 8350 10467 8414
rect 10485 8350 10549 8414
rect 10567 8350 10631 8414
rect 10649 8350 10713 8414
rect 10731 8350 10795 8414
rect 10813 8350 10877 8414
rect 10895 8350 10959 8414
rect 10977 8350 11041 8414
rect 11059 8350 11123 8414
rect 11141 8350 11205 8414
rect 11223 8350 11287 8414
rect 11305 8350 11369 8414
rect 11387 8350 11451 8414
rect 11468 8350 11532 8414
rect 11549 8350 11613 8414
rect 11630 8350 11694 8414
rect 11711 8350 11775 8414
rect 11792 8350 11856 8414
rect 11873 8350 11937 8414
rect 11954 8350 12018 8414
rect 12035 8350 12099 8414
rect 12116 8350 12180 8414
rect 12197 8350 12261 8414
rect 12278 8350 12342 8414
rect 12359 8350 12423 8414
rect 12440 8350 12504 8414
rect 12521 8350 12585 8414
rect 12602 8350 12666 8414
rect 12683 8350 12747 8414
rect 12764 8350 12828 8414
rect 12845 8350 12909 8414
rect 12926 8350 12990 8414
rect 13007 8350 13071 8414
rect 13088 8350 13152 8414
rect 13169 8350 13233 8414
rect 13250 8350 13314 8414
rect 13331 8350 13395 8414
rect 13412 8350 13476 8414
rect 13493 8350 13557 8414
rect 13574 8350 13638 8414
rect 13655 8350 13719 8414
rect 13736 8350 13800 8414
rect 13817 8350 13881 8414
rect 13898 8350 13962 8414
rect 13979 8350 14043 8414
rect 14060 8350 14124 8414
rect 14141 8350 14205 8414
rect 14222 8350 14286 8414
rect 14303 8350 14367 8414
rect 14384 8350 14448 8414
rect 14465 8350 14529 8414
rect 14546 8350 14610 8414
rect 14627 8350 14691 8414
rect 14708 8350 14772 8414
rect 14789 8350 14853 8414
rect 14870 8350 14934 8414
rect 10157 8264 10221 8328
rect 10239 8264 10303 8328
rect 10321 8264 10385 8328
rect 10403 8264 10467 8328
rect 10485 8264 10549 8328
rect 10567 8264 10631 8328
rect 10649 8264 10713 8328
rect 10731 8264 10795 8328
rect 10813 8264 10877 8328
rect 10895 8264 10959 8328
rect 10977 8264 11041 8328
rect 11059 8264 11123 8328
rect 11141 8264 11205 8328
rect 11223 8264 11287 8328
rect 11305 8264 11369 8328
rect 11387 8264 11451 8328
rect 11468 8264 11532 8328
rect 11549 8264 11613 8328
rect 11630 8264 11694 8328
rect 11711 8264 11775 8328
rect 11792 8264 11856 8328
rect 11873 8264 11937 8328
rect 11954 8264 12018 8328
rect 12035 8264 12099 8328
rect 12116 8264 12180 8328
rect 12197 8264 12261 8328
rect 12278 8264 12342 8328
rect 12359 8264 12423 8328
rect 12440 8264 12504 8328
rect 12521 8264 12585 8328
rect 12602 8264 12666 8328
rect 12683 8264 12747 8328
rect 12764 8264 12828 8328
rect 12845 8264 12909 8328
rect 12926 8264 12990 8328
rect 13007 8264 13071 8328
rect 13088 8264 13152 8328
rect 13169 8264 13233 8328
rect 13250 8264 13314 8328
rect 13331 8264 13395 8328
rect 13412 8264 13476 8328
rect 13493 8264 13557 8328
rect 13574 8264 13638 8328
rect 13655 8264 13719 8328
rect 13736 8264 13800 8328
rect 13817 8264 13881 8328
rect 13898 8264 13962 8328
rect 13979 8264 14043 8328
rect 14060 8264 14124 8328
rect 14141 8264 14205 8328
rect 14222 8264 14286 8328
rect 14303 8264 14367 8328
rect 14384 8264 14448 8328
rect 14465 8264 14529 8328
rect 14546 8264 14610 8328
rect 14627 8264 14691 8328
rect 14708 8264 14772 8328
rect 14789 8264 14853 8328
rect 14870 8264 14934 8328
rect 10157 8178 10221 8242
rect 10239 8178 10303 8242
rect 10321 8178 10385 8242
rect 10403 8178 10467 8242
rect 10485 8178 10549 8242
rect 10567 8178 10631 8242
rect 10649 8178 10713 8242
rect 10731 8178 10795 8242
rect 10813 8178 10877 8242
rect 10895 8178 10959 8242
rect 10977 8178 11041 8242
rect 11059 8178 11123 8242
rect 11141 8178 11205 8242
rect 11223 8178 11287 8242
rect 11305 8178 11369 8242
rect 11387 8178 11451 8242
rect 11468 8178 11532 8242
rect 11549 8178 11613 8242
rect 11630 8178 11694 8242
rect 11711 8178 11775 8242
rect 11792 8178 11856 8242
rect 11873 8178 11937 8242
rect 11954 8178 12018 8242
rect 12035 8178 12099 8242
rect 12116 8178 12180 8242
rect 12197 8178 12261 8242
rect 12278 8178 12342 8242
rect 12359 8178 12423 8242
rect 12440 8178 12504 8242
rect 12521 8178 12585 8242
rect 12602 8178 12666 8242
rect 12683 8178 12747 8242
rect 12764 8178 12828 8242
rect 12845 8178 12909 8242
rect 12926 8178 12990 8242
rect 13007 8178 13071 8242
rect 13088 8178 13152 8242
rect 13169 8178 13233 8242
rect 13250 8178 13314 8242
rect 13331 8178 13395 8242
rect 13412 8178 13476 8242
rect 13493 8178 13557 8242
rect 13574 8178 13638 8242
rect 13655 8178 13719 8242
rect 13736 8178 13800 8242
rect 13817 8178 13881 8242
rect 13898 8178 13962 8242
rect 13979 8178 14043 8242
rect 14060 8178 14124 8242
rect 14141 8178 14205 8242
rect 14222 8178 14286 8242
rect 14303 8178 14367 8242
rect 14384 8178 14448 8242
rect 14465 8178 14529 8242
rect 14546 8178 14610 8242
rect 14627 8178 14691 8242
rect 14708 8178 14772 8242
rect 14789 8178 14853 8242
rect 14870 8178 14934 8242
rect 10157 8092 10221 8156
rect 10239 8092 10303 8156
rect 10321 8092 10385 8156
rect 10403 8092 10467 8156
rect 10485 8092 10549 8156
rect 10567 8092 10631 8156
rect 10649 8092 10713 8156
rect 10731 8092 10795 8156
rect 10813 8092 10877 8156
rect 10895 8092 10959 8156
rect 10977 8092 11041 8156
rect 11059 8092 11123 8156
rect 11141 8092 11205 8156
rect 11223 8092 11287 8156
rect 11305 8092 11369 8156
rect 11387 8092 11451 8156
rect 11468 8092 11532 8156
rect 11549 8092 11613 8156
rect 11630 8092 11694 8156
rect 11711 8092 11775 8156
rect 11792 8092 11856 8156
rect 11873 8092 11937 8156
rect 11954 8092 12018 8156
rect 12035 8092 12099 8156
rect 12116 8092 12180 8156
rect 12197 8092 12261 8156
rect 12278 8092 12342 8156
rect 12359 8092 12423 8156
rect 12440 8092 12504 8156
rect 12521 8092 12585 8156
rect 12602 8092 12666 8156
rect 12683 8092 12747 8156
rect 12764 8092 12828 8156
rect 12845 8092 12909 8156
rect 12926 8092 12990 8156
rect 13007 8092 13071 8156
rect 13088 8092 13152 8156
rect 13169 8092 13233 8156
rect 13250 8092 13314 8156
rect 13331 8092 13395 8156
rect 13412 8092 13476 8156
rect 13493 8092 13557 8156
rect 13574 8092 13638 8156
rect 13655 8092 13719 8156
rect 13736 8092 13800 8156
rect 13817 8092 13881 8156
rect 13898 8092 13962 8156
rect 13979 8092 14043 8156
rect 14060 8092 14124 8156
rect 14141 8092 14205 8156
rect 14222 8092 14286 8156
rect 14303 8092 14367 8156
rect 14384 8092 14448 8156
rect 14465 8092 14529 8156
rect 14546 8092 14610 8156
rect 14627 8092 14691 8156
rect 14708 8092 14772 8156
rect 14789 8092 14853 8156
rect 14870 8092 14934 8156
rect 10157 8006 10221 8070
rect 10239 8006 10303 8070
rect 10321 8006 10385 8070
rect 10403 8006 10467 8070
rect 10485 8006 10549 8070
rect 10567 8006 10631 8070
rect 10649 8006 10713 8070
rect 10731 8006 10795 8070
rect 10813 8006 10877 8070
rect 10895 8006 10959 8070
rect 10977 8006 11041 8070
rect 11059 8006 11123 8070
rect 11141 8006 11205 8070
rect 11223 8006 11287 8070
rect 11305 8006 11369 8070
rect 11387 8006 11451 8070
rect 11468 8006 11532 8070
rect 11549 8006 11613 8070
rect 11630 8006 11694 8070
rect 11711 8006 11775 8070
rect 11792 8006 11856 8070
rect 11873 8006 11937 8070
rect 11954 8006 12018 8070
rect 12035 8006 12099 8070
rect 12116 8006 12180 8070
rect 12197 8006 12261 8070
rect 12278 8006 12342 8070
rect 12359 8006 12423 8070
rect 12440 8006 12504 8070
rect 12521 8006 12585 8070
rect 12602 8006 12666 8070
rect 12683 8006 12747 8070
rect 12764 8006 12828 8070
rect 12845 8006 12909 8070
rect 12926 8006 12990 8070
rect 13007 8006 13071 8070
rect 13088 8006 13152 8070
rect 13169 8006 13233 8070
rect 13250 8006 13314 8070
rect 13331 8006 13395 8070
rect 13412 8006 13476 8070
rect 13493 8006 13557 8070
rect 13574 8006 13638 8070
rect 13655 8006 13719 8070
rect 13736 8006 13800 8070
rect 13817 8006 13881 8070
rect 13898 8006 13962 8070
rect 13979 8006 14043 8070
rect 14060 8006 14124 8070
rect 14141 8006 14205 8070
rect 14222 8006 14286 8070
rect 14303 8006 14367 8070
rect 14384 8006 14448 8070
rect 14465 8006 14529 8070
rect 14546 8006 14610 8070
rect 14627 8006 14691 8070
rect 14708 8006 14772 8070
rect 14789 8006 14853 8070
rect 14870 8006 14934 8070
rect 10157 7920 10221 7984
rect 10239 7920 10303 7984
rect 10321 7920 10385 7984
rect 10403 7920 10467 7984
rect 10485 7920 10549 7984
rect 10567 7920 10631 7984
rect 10649 7920 10713 7984
rect 10731 7920 10795 7984
rect 10813 7920 10877 7984
rect 10895 7920 10959 7984
rect 10977 7920 11041 7984
rect 11059 7920 11123 7984
rect 11141 7920 11205 7984
rect 11223 7920 11287 7984
rect 11305 7920 11369 7984
rect 11387 7920 11451 7984
rect 11468 7920 11532 7984
rect 11549 7920 11613 7984
rect 11630 7920 11694 7984
rect 11711 7920 11775 7984
rect 11792 7920 11856 7984
rect 11873 7920 11937 7984
rect 11954 7920 12018 7984
rect 12035 7920 12099 7984
rect 12116 7920 12180 7984
rect 12197 7920 12261 7984
rect 12278 7920 12342 7984
rect 12359 7920 12423 7984
rect 12440 7920 12504 7984
rect 12521 7920 12585 7984
rect 12602 7920 12666 7984
rect 12683 7920 12747 7984
rect 12764 7920 12828 7984
rect 12845 7920 12909 7984
rect 12926 7920 12990 7984
rect 13007 7920 13071 7984
rect 13088 7920 13152 7984
rect 13169 7920 13233 7984
rect 13250 7920 13314 7984
rect 13331 7920 13395 7984
rect 13412 7920 13476 7984
rect 13493 7920 13557 7984
rect 13574 7920 13638 7984
rect 13655 7920 13719 7984
rect 13736 7920 13800 7984
rect 13817 7920 13881 7984
rect 13898 7920 13962 7984
rect 13979 7920 14043 7984
rect 14060 7920 14124 7984
rect 14141 7920 14205 7984
rect 14222 7920 14286 7984
rect 14303 7920 14367 7984
rect 14384 7920 14448 7984
rect 14465 7920 14529 7984
rect 14546 7920 14610 7984
rect 14627 7920 14691 7984
rect 14708 7920 14772 7984
rect 14789 7920 14853 7984
rect 14870 7920 14934 7984
<< metal4 >>
rect 0 34757 254 39600
rect 14746 34757 15000 39600
rect 0 13607 254 18600
rect 14746 13607 15000 18600
rect 0 12417 254 13307
rect 14746 12417 15000 13307
rect 0 11247 254 12137
rect 14746 11247 15000 12137
rect 0 10881 254 10947
rect 14746 10881 15000 10947
rect 0 10225 254 10821
rect 14746 10225 15000 10821
rect 0 9929 254 10165
rect 14746 9929 15000 10165
rect 0 9273 254 9869
rect 14746 9273 15000 9869
rect 0 9147 254 9213
rect 14746 9147 15000 9213
rect 0 8844 4895 8847
rect 0 8780 106 8844
rect 170 8780 187 8844
rect 251 8780 268 8844
rect 332 8780 349 8844
rect 413 8780 430 8844
rect 494 8780 510 8844
rect 574 8780 590 8844
rect 654 8780 670 8844
rect 734 8780 750 8844
rect 814 8780 830 8844
rect 894 8780 910 8844
rect 974 8780 990 8844
rect 1054 8780 1070 8844
rect 1134 8780 1150 8844
rect 1214 8780 1230 8844
rect 1294 8780 1310 8844
rect 1374 8780 1390 8844
rect 1454 8780 1470 8844
rect 1534 8780 1550 8844
rect 1614 8780 1630 8844
rect 1694 8780 1710 8844
rect 1774 8780 1790 8844
rect 1854 8780 1870 8844
rect 1934 8780 1950 8844
rect 2014 8780 2030 8844
rect 2094 8780 2110 8844
rect 2174 8780 2190 8844
rect 2254 8780 2270 8844
rect 2334 8780 2350 8844
rect 2414 8780 2430 8844
rect 2494 8780 2510 8844
rect 2574 8780 2590 8844
rect 2654 8780 2670 8844
rect 2734 8780 2750 8844
rect 2814 8780 2830 8844
rect 2894 8780 2910 8844
rect 2974 8780 2990 8844
rect 3054 8780 3070 8844
rect 3134 8780 3150 8844
rect 3214 8780 3230 8844
rect 3294 8780 3310 8844
rect 3374 8780 3390 8844
rect 3454 8780 3470 8844
rect 3534 8780 3550 8844
rect 3614 8780 3630 8844
rect 3694 8780 3710 8844
rect 3774 8780 3790 8844
rect 3854 8780 3870 8844
rect 3934 8780 3950 8844
rect 4014 8780 4030 8844
rect 4094 8780 4110 8844
rect 4174 8780 4190 8844
rect 4254 8780 4270 8844
rect 4334 8780 4350 8844
rect 4414 8780 4430 8844
rect 4494 8780 4510 8844
rect 4574 8780 4590 8844
rect 4654 8780 4670 8844
rect 4734 8780 4750 8844
rect 4814 8780 4830 8844
rect 4894 8780 4895 8844
rect 0 8758 4895 8780
rect 0 8694 106 8758
rect 170 8694 187 8758
rect 251 8694 268 8758
rect 332 8694 349 8758
rect 413 8694 430 8758
rect 494 8694 510 8758
rect 574 8694 590 8758
rect 654 8694 670 8758
rect 734 8694 750 8758
rect 814 8694 830 8758
rect 894 8694 910 8758
rect 974 8694 990 8758
rect 1054 8694 1070 8758
rect 1134 8694 1150 8758
rect 1214 8694 1230 8758
rect 1294 8694 1310 8758
rect 1374 8694 1390 8758
rect 1454 8694 1470 8758
rect 1534 8694 1550 8758
rect 1614 8694 1630 8758
rect 1694 8694 1710 8758
rect 1774 8694 1790 8758
rect 1854 8694 1870 8758
rect 1934 8694 1950 8758
rect 2014 8694 2030 8758
rect 2094 8694 2110 8758
rect 2174 8694 2190 8758
rect 2254 8694 2270 8758
rect 2334 8694 2350 8758
rect 2414 8694 2430 8758
rect 2494 8694 2510 8758
rect 2574 8694 2590 8758
rect 2654 8694 2670 8758
rect 2734 8694 2750 8758
rect 2814 8694 2830 8758
rect 2894 8694 2910 8758
rect 2974 8694 2990 8758
rect 3054 8694 3070 8758
rect 3134 8694 3150 8758
rect 3214 8694 3230 8758
rect 3294 8694 3310 8758
rect 3374 8694 3390 8758
rect 3454 8694 3470 8758
rect 3534 8694 3550 8758
rect 3614 8694 3630 8758
rect 3694 8694 3710 8758
rect 3774 8694 3790 8758
rect 3854 8694 3870 8758
rect 3934 8694 3950 8758
rect 4014 8694 4030 8758
rect 4094 8694 4110 8758
rect 4174 8694 4190 8758
rect 4254 8694 4270 8758
rect 4334 8694 4350 8758
rect 4414 8694 4430 8758
rect 4494 8694 4510 8758
rect 4574 8694 4590 8758
rect 4654 8694 4670 8758
rect 4734 8694 4750 8758
rect 4814 8694 4830 8758
rect 4894 8694 4895 8758
rect 0 8672 4895 8694
rect 0 8608 106 8672
rect 170 8608 187 8672
rect 251 8608 268 8672
rect 332 8608 349 8672
rect 413 8608 430 8672
rect 494 8608 510 8672
rect 574 8608 590 8672
rect 654 8608 670 8672
rect 734 8608 750 8672
rect 814 8608 830 8672
rect 894 8608 910 8672
rect 974 8608 990 8672
rect 1054 8608 1070 8672
rect 1134 8608 1150 8672
rect 1214 8608 1230 8672
rect 1294 8608 1310 8672
rect 1374 8608 1390 8672
rect 1454 8608 1470 8672
rect 1534 8608 1550 8672
rect 1614 8608 1630 8672
rect 1694 8608 1710 8672
rect 1774 8608 1790 8672
rect 1854 8608 1870 8672
rect 1934 8608 1950 8672
rect 2014 8608 2030 8672
rect 2094 8608 2110 8672
rect 2174 8608 2190 8672
rect 2254 8608 2270 8672
rect 2334 8608 2350 8672
rect 2414 8608 2430 8672
rect 2494 8608 2510 8672
rect 2574 8608 2590 8672
rect 2654 8608 2670 8672
rect 2734 8608 2750 8672
rect 2814 8608 2830 8672
rect 2894 8608 2910 8672
rect 2974 8608 2990 8672
rect 3054 8608 3070 8672
rect 3134 8608 3150 8672
rect 3214 8608 3230 8672
rect 3294 8608 3310 8672
rect 3374 8608 3390 8672
rect 3454 8608 3470 8672
rect 3534 8608 3550 8672
rect 3614 8608 3630 8672
rect 3694 8608 3710 8672
rect 3774 8608 3790 8672
rect 3854 8608 3870 8672
rect 3934 8608 3950 8672
rect 4014 8608 4030 8672
rect 4094 8608 4110 8672
rect 4174 8608 4190 8672
rect 4254 8608 4270 8672
rect 4334 8608 4350 8672
rect 4414 8608 4430 8672
rect 4494 8608 4510 8672
rect 4574 8608 4590 8672
rect 4654 8608 4670 8672
rect 4734 8608 4750 8672
rect 4814 8608 4830 8672
rect 4894 8608 4895 8672
rect 0 8586 4895 8608
rect 0 8522 106 8586
rect 170 8522 187 8586
rect 251 8522 268 8586
rect 332 8522 349 8586
rect 413 8522 430 8586
rect 494 8522 510 8586
rect 574 8522 590 8586
rect 654 8522 670 8586
rect 734 8522 750 8586
rect 814 8522 830 8586
rect 894 8522 910 8586
rect 974 8522 990 8586
rect 1054 8522 1070 8586
rect 1134 8522 1150 8586
rect 1214 8522 1230 8586
rect 1294 8522 1310 8586
rect 1374 8522 1390 8586
rect 1454 8522 1470 8586
rect 1534 8522 1550 8586
rect 1614 8522 1630 8586
rect 1694 8522 1710 8586
rect 1774 8522 1790 8586
rect 1854 8522 1870 8586
rect 1934 8522 1950 8586
rect 2014 8522 2030 8586
rect 2094 8522 2110 8586
rect 2174 8522 2190 8586
rect 2254 8522 2270 8586
rect 2334 8522 2350 8586
rect 2414 8522 2430 8586
rect 2494 8522 2510 8586
rect 2574 8522 2590 8586
rect 2654 8522 2670 8586
rect 2734 8522 2750 8586
rect 2814 8522 2830 8586
rect 2894 8522 2910 8586
rect 2974 8522 2990 8586
rect 3054 8522 3070 8586
rect 3134 8522 3150 8586
rect 3214 8522 3230 8586
rect 3294 8522 3310 8586
rect 3374 8522 3390 8586
rect 3454 8522 3470 8586
rect 3534 8522 3550 8586
rect 3614 8522 3630 8586
rect 3694 8522 3710 8586
rect 3774 8522 3790 8586
rect 3854 8522 3870 8586
rect 3934 8522 3950 8586
rect 4014 8522 4030 8586
rect 4094 8522 4110 8586
rect 4174 8522 4190 8586
rect 4254 8522 4270 8586
rect 4334 8522 4350 8586
rect 4414 8522 4430 8586
rect 4494 8522 4510 8586
rect 4574 8522 4590 8586
rect 4654 8522 4670 8586
rect 4734 8522 4750 8586
rect 4814 8522 4830 8586
rect 4894 8522 4895 8586
rect 0 8500 4895 8522
rect 0 8436 106 8500
rect 170 8436 187 8500
rect 251 8436 268 8500
rect 332 8436 349 8500
rect 413 8436 430 8500
rect 494 8436 510 8500
rect 574 8436 590 8500
rect 654 8436 670 8500
rect 734 8436 750 8500
rect 814 8436 830 8500
rect 894 8436 910 8500
rect 974 8436 990 8500
rect 1054 8436 1070 8500
rect 1134 8436 1150 8500
rect 1214 8436 1230 8500
rect 1294 8436 1310 8500
rect 1374 8436 1390 8500
rect 1454 8436 1470 8500
rect 1534 8436 1550 8500
rect 1614 8436 1630 8500
rect 1694 8436 1710 8500
rect 1774 8436 1790 8500
rect 1854 8436 1870 8500
rect 1934 8436 1950 8500
rect 2014 8436 2030 8500
rect 2094 8436 2110 8500
rect 2174 8436 2190 8500
rect 2254 8436 2270 8500
rect 2334 8436 2350 8500
rect 2414 8436 2430 8500
rect 2494 8436 2510 8500
rect 2574 8436 2590 8500
rect 2654 8436 2670 8500
rect 2734 8436 2750 8500
rect 2814 8436 2830 8500
rect 2894 8436 2910 8500
rect 2974 8436 2990 8500
rect 3054 8436 3070 8500
rect 3134 8436 3150 8500
rect 3214 8436 3230 8500
rect 3294 8436 3310 8500
rect 3374 8436 3390 8500
rect 3454 8436 3470 8500
rect 3534 8436 3550 8500
rect 3614 8436 3630 8500
rect 3694 8436 3710 8500
rect 3774 8436 3790 8500
rect 3854 8436 3870 8500
rect 3934 8436 3950 8500
rect 4014 8436 4030 8500
rect 4094 8436 4110 8500
rect 4174 8436 4190 8500
rect 4254 8436 4270 8500
rect 4334 8436 4350 8500
rect 4414 8436 4430 8500
rect 4494 8436 4510 8500
rect 4574 8436 4590 8500
rect 4654 8436 4670 8500
rect 4734 8436 4750 8500
rect 4814 8436 4830 8500
rect 4894 8436 4895 8500
rect 0 8414 4895 8436
rect 0 8350 106 8414
rect 170 8350 187 8414
rect 251 8350 268 8414
rect 332 8350 349 8414
rect 413 8350 430 8414
rect 494 8350 510 8414
rect 574 8350 590 8414
rect 654 8350 670 8414
rect 734 8350 750 8414
rect 814 8350 830 8414
rect 894 8350 910 8414
rect 974 8350 990 8414
rect 1054 8350 1070 8414
rect 1134 8350 1150 8414
rect 1214 8350 1230 8414
rect 1294 8350 1310 8414
rect 1374 8350 1390 8414
rect 1454 8350 1470 8414
rect 1534 8350 1550 8414
rect 1614 8350 1630 8414
rect 1694 8350 1710 8414
rect 1774 8350 1790 8414
rect 1854 8350 1870 8414
rect 1934 8350 1950 8414
rect 2014 8350 2030 8414
rect 2094 8350 2110 8414
rect 2174 8350 2190 8414
rect 2254 8350 2270 8414
rect 2334 8350 2350 8414
rect 2414 8350 2430 8414
rect 2494 8350 2510 8414
rect 2574 8350 2590 8414
rect 2654 8350 2670 8414
rect 2734 8350 2750 8414
rect 2814 8350 2830 8414
rect 2894 8350 2910 8414
rect 2974 8350 2990 8414
rect 3054 8350 3070 8414
rect 3134 8350 3150 8414
rect 3214 8350 3230 8414
rect 3294 8350 3310 8414
rect 3374 8350 3390 8414
rect 3454 8350 3470 8414
rect 3534 8350 3550 8414
rect 3614 8350 3630 8414
rect 3694 8350 3710 8414
rect 3774 8350 3790 8414
rect 3854 8350 3870 8414
rect 3934 8350 3950 8414
rect 4014 8350 4030 8414
rect 4094 8350 4110 8414
rect 4174 8350 4190 8414
rect 4254 8350 4270 8414
rect 4334 8350 4350 8414
rect 4414 8350 4430 8414
rect 4494 8350 4510 8414
rect 4574 8350 4590 8414
rect 4654 8350 4670 8414
rect 4734 8350 4750 8414
rect 4814 8350 4830 8414
rect 4894 8350 4895 8414
rect 0 8328 4895 8350
rect 0 8264 106 8328
rect 170 8264 187 8328
rect 251 8264 268 8328
rect 332 8264 349 8328
rect 413 8264 430 8328
rect 494 8264 510 8328
rect 574 8264 590 8328
rect 654 8264 670 8328
rect 734 8264 750 8328
rect 814 8264 830 8328
rect 894 8264 910 8328
rect 974 8264 990 8328
rect 1054 8264 1070 8328
rect 1134 8264 1150 8328
rect 1214 8264 1230 8328
rect 1294 8264 1310 8328
rect 1374 8264 1390 8328
rect 1454 8264 1470 8328
rect 1534 8264 1550 8328
rect 1614 8264 1630 8328
rect 1694 8264 1710 8328
rect 1774 8264 1790 8328
rect 1854 8264 1870 8328
rect 1934 8264 1950 8328
rect 2014 8264 2030 8328
rect 2094 8264 2110 8328
rect 2174 8264 2190 8328
rect 2254 8264 2270 8328
rect 2334 8264 2350 8328
rect 2414 8264 2430 8328
rect 2494 8264 2510 8328
rect 2574 8264 2590 8328
rect 2654 8264 2670 8328
rect 2734 8264 2750 8328
rect 2814 8264 2830 8328
rect 2894 8264 2910 8328
rect 2974 8264 2990 8328
rect 3054 8264 3070 8328
rect 3134 8264 3150 8328
rect 3214 8264 3230 8328
rect 3294 8264 3310 8328
rect 3374 8264 3390 8328
rect 3454 8264 3470 8328
rect 3534 8264 3550 8328
rect 3614 8264 3630 8328
rect 3694 8264 3710 8328
rect 3774 8264 3790 8328
rect 3854 8264 3870 8328
rect 3934 8264 3950 8328
rect 4014 8264 4030 8328
rect 4094 8264 4110 8328
rect 4174 8264 4190 8328
rect 4254 8264 4270 8328
rect 4334 8264 4350 8328
rect 4414 8264 4430 8328
rect 4494 8264 4510 8328
rect 4574 8264 4590 8328
rect 4654 8264 4670 8328
rect 4734 8264 4750 8328
rect 4814 8264 4830 8328
rect 4894 8264 4895 8328
rect 0 8242 4895 8264
rect 0 8178 106 8242
rect 170 8178 187 8242
rect 251 8178 268 8242
rect 332 8178 349 8242
rect 413 8178 430 8242
rect 494 8178 510 8242
rect 574 8178 590 8242
rect 654 8178 670 8242
rect 734 8178 750 8242
rect 814 8178 830 8242
rect 894 8178 910 8242
rect 974 8178 990 8242
rect 1054 8178 1070 8242
rect 1134 8178 1150 8242
rect 1214 8178 1230 8242
rect 1294 8178 1310 8242
rect 1374 8178 1390 8242
rect 1454 8178 1470 8242
rect 1534 8178 1550 8242
rect 1614 8178 1630 8242
rect 1694 8178 1710 8242
rect 1774 8178 1790 8242
rect 1854 8178 1870 8242
rect 1934 8178 1950 8242
rect 2014 8178 2030 8242
rect 2094 8178 2110 8242
rect 2174 8178 2190 8242
rect 2254 8178 2270 8242
rect 2334 8178 2350 8242
rect 2414 8178 2430 8242
rect 2494 8178 2510 8242
rect 2574 8178 2590 8242
rect 2654 8178 2670 8242
rect 2734 8178 2750 8242
rect 2814 8178 2830 8242
rect 2894 8178 2910 8242
rect 2974 8178 2990 8242
rect 3054 8178 3070 8242
rect 3134 8178 3150 8242
rect 3214 8178 3230 8242
rect 3294 8178 3310 8242
rect 3374 8178 3390 8242
rect 3454 8178 3470 8242
rect 3534 8178 3550 8242
rect 3614 8178 3630 8242
rect 3694 8178 3710 8242
rect 3774 8178 3790 8242
rect 3854 8178 3870 8242
rect 3934 8178 3950 8242
rect 4014 8178 4030 8242
rect 4094 8178 4110 8242
rect 4174 8178 4190 8242
rect 4254 8178 4270 8242
rect 4334 8178 4350 8242
rect 4414 8178 4430 8242
rect 4494 8178 4510 8242
rect 4574 8178 4590 8242
rect 4654 8178 4670 8242
rect 4734 8178 4750 8242
rect 4814 8178 4830 8242
rect 4894 8178 4895 8242
rect 0 8156 4895 8178
rect 0 8092 106 8156
rect 170 8092 187 8156
rect 251 8092 268 8156
rect 332 8092 349 8156
rect 413 8092 430 8156
rect 494 8092 510 8156
rect 574 8092 590 8156
rect 654 8092 670 8156
rect 734 8092 750 8156
rect 814 8092 830 8156
rect 894 8092 910 8156
rect 974 8092 990 8156
rect 1054 8092 1070 8156
rect 1134 8092 1150 8156
rect 1214 8092 1230 8156
rect 1294 8092 1310 8156
rect 1374 8092 1390 8156
rect 1454 8092 1470 8156
rect 1534 8092 1550 8156
rect 1614 8092 1630 8156
rect 1694 8092 1710 8156
rect 1774 8092 1790 8156
rect 1854 8092 1870 8156
rect 1934 8092 1950 8156
rect 2014 8092 2030 8156
rect 2094 8092 2110 8156
rect 2174 8092 2190 8156
rect 2254 8092 2270 8156
rect 2334 8092 2350 8156
rect 2414 8092 2430 8156
rect 2494 8092 2510 8156
rect 2574 8092 2590 8156
rect 2654 8092 2670 8156
rect 2734 8092 2750 8156
rect 2814 8092 2830 8156
rect 2894 8092 2910 8156
rect 2974 8092 2990 8156
rect 3054 8092 3070 8156
rect 3134 8092 3150 8156
rect 3214 8092 3230 8156
rect 3294 8092 3310 8156
rect 3374 8092 3390 8156
rect 3454 8092 3470 8156
rect 3534 8092 3550 8156
rect 3614 8092 3630 8156
rect 3694 8092 3710 8156
rect 3774 8092 3790 8156
rect 3854 8092 3870 8156
rect 3934 8092 3950 8156
rect 4014 8092 4030 8156
rect 4094 8092 4110 8156
rect 4174 8092 4190 8156
rect 4254 8092 4270 8156
rect 4334 8092 4350 8156
rect 4414 8092 4430 8156
rect 4494 8092 4510 8156
rect 4574 8092 4590 8156
rect 4654 8092 4670 8156
rect 4734 8092 4750 8156
rect 4814 8092 4830 8156
rect 4894 8092 4895 8156
rect 0 8070 4895 8092
rect 0 8006 106 8070
rect 170 8006 187 8070
rect 251 8006 268 8070
rect 332 8006 349 8070
rect 413 8006 430 8070
rect 494 8006 510 8070
rect 574 8006 590 8070
rect 654 8006 670 8070
rect 734 8006 750 8070
rect 814 8006 830 8070
rect 894 8006 910 8070
rect 974 8006 990 8070
rect 1054 8006 1070 8070
rect 1134 8006 1150 8070
rect 1214 8006 1230 8070
rect 1294 8006 1310 8070
rect 1374 8006 1390 8070
rect 1454 8006 1470 8070
rect 1534 8006 1550 8070
rect 1614 8006 1630 8070
rect 1694 8006 1710 8070
rect 1774 8006 1790 8070
rect 1854 8006 1870 8070
rect 1934 8006 1950 8070
rect 2014 8006 2030 8070
rect 2094 8006 2110 8070
rect 2174 8006 2190 8070
rect 2254 8006 2270 8070
rect 2334 8006 2350 8070
rect 2414 8006 2430 8070
rect 2494 8006 2510 8070
rect 2574 8006 2590 8070
rect 2654 8006 2670 8070
rect 2734 8006 2750 8070
rect 2814 8006 2830 8070
rect 2894 8006 2910 8070
rect 2974 8006 2990 8070
rect 3054 8006 3070 8070
rect 3134 8006 3150 8070
rect 3214 8006 3230 8070
rect 3294 8006 3310 8070
rect 3374 8006 3390 8070
rect 3454 8006 3470 8070
rect 3534 8006 3550 8070
rect 3614 8006 3630 8070
rect 3694 8006 3710 8070
rect 3774 8006 3790 8070
rect 3854 8006 3870 8070
rect 3934 8006 3950 8070
rect 4014 8006 4030 8070
rect 4094 8006 4110 8070
rect 4174 8006 4190 8070
rect 4254 8006 4270 8070
rect 4334 8006 4350 8070
rect 4414 8006 4430 8070
rect 4494 8006 4510 8070
rect 4574 8006 4590 8070
rect 4654 8006 4670 8070
rect 4734 8006 4750 8070
rect 4814 8006 4830 8070
rect 4894 8006 4895 8070
rect 0 7984 4895 8006
rect 0 7920 106 7984
rect 170 7920 187 7984
rect 251 7920 268 7984
rect 332 7920 349 7984
rect 413 7920 430 7984
rect 494 7920 510 7984
rect 574 7920 590 7984
rect 654 7920 670 7984
rect 734 7920 750 7984
rect 814 7920 830 7984
rect 894 7920 910 7984
rect 974 7920 990 7984
rect 1054 7920 1070 7984
rect 1134 7920 1150 7984
rect 1214 7920 1230 7984
rect 1294 7920 1310 7984
rect 1374 7920 1390 7984
rect 1454 7920 1470 7984
rect 1534 7920 1550 7984
rect 1614 7920 1630 7984
rect 1694 7920 1710 7984
rect 1774 7920 1790 7984
rect 1854 7920 1870 7984
rect 1934 7920 1950 7984
rect 2014 7920 2030 7984
rect 2094 7920 2110 7984
rect 2174 7920 2190 7984
rect 2254 7920 2270 7984
rect 2334 7920 2350 7984
rect 2414 7920 2430 7984
rect 2494 7920 2510 7984
rect 2574 7920 2590 7984
rect 2654 7920 2670 7984
rect 2734 7920 2750 7984
rect 2814 7920 2830 7984
rect 2894 7920 2910 7984
rect 2974 7920 2990 7984
rect 3054 7920 3070 7984
rect 3134 7920 3150 7984
rect 3214 7920 3230 7984
rect 3294 7920 3310 7984
rect 3374 7920 3390 7984
rect 3454 7920 3470 7984
rect 3534 7920 3550 7984
rect 3614 7920 3630 7984
rect 3694 7920 3710 7984
rect 3774 7920 3790 7984
rect 3854 7920 3870 7984
rect 3934 7920 3950 7984
rect 4014 7920 4030 7984
rect 4094 7920 4110 7984
rect 4174 7920 4190 7984
rect 4254 7920 4270 7984
rect 4334 7920 4350 7984
rect 4414 7920 4430 7984
rect 4494 7920 4510 7984
rect 4574 7920 4590 7984
rect 4654 7920 4670 7984
rect 4734 7920 4750 7984
rect 4814 7920 4830 7984
rect 4894 7920 4895 7984
rect 0 7917 4895 7920
rect 10156 8844 15000 8847
rect 10156 8780 10157 8844
rect 10221 8780 10239 8844
rect 10303 8780 10321 8844
rect 10385 8780 10403 8844
rect 10467 8780 10485 8844
rect 10549 8780 10567 8844
rect 10631 8780 10649 8844
rect 10713 8780 10731 8844
rect 10795 8780 10813 8844
rect 10877 8780 10895 8844
rect 10959 8780 10977 8844
rect 11041 8780 11059 8844
rect 11123 8780 11141 8844
rect 11205 8780 11223 8844
rect 11287 8780 11305 8844
rect 11369 8780 11387 8844
rect 11451 8780 11468 8844
rect 11532 8780 11549 8844
rect 11613 8780 11630 8844
rect 11694 8780 11711 8844
rect 11775 8780 11792 8844
rect 11856 8780 11873 8844
rect 11937 8780 11954 8844
rect 12018 8780 12035 8844
rect 12099 8780 12116 8844
rect 12180 8780 12197 8844
rect 12261 8780 12278 8844
rect 12342 8780 12359 8844
rect 12423 8780 12440 8844
rect 12504 8780 12521 8844
rect 12585 8780 12602 8844
rect 12666 8780 12683 8844
rect 12747 8780 12764 8844
rect 12828 8780 12845 8844
rect 12909 8780 12926 8844
rect 12990 8780 13007 8844
rect 13071 8780 13088 8844
rect 13152 8780 13169 8844
rect 13233 8780 13250 8844
rect 13314 8780 13331 8844
rect 13395 8780 13412 8844
rect 13476 8780 13493 8844
rect 13557 8780 13574 8844
rect 13638 8780 13655 8844
rect 13719 8780 13736 8844
rect 13800 8780 13817 8844
rect 13881 8780 13898 8844
rect 13962 8780 13979 8844
rect 14043 8780 14060 8844
rect 14124 8780 14141 8844
rect 14205 8780 14222 8844
rect 14286 8780 14303 8844
rect 14367 8780 14384 8844
rect 14448 8780 14465 8844
rect 14529 8780 14546 8844
rect 14610 8780 14627 8844
rect 14691 8780 14708 8844
rect 14772 8780 14789 8844
rect 14853 8780 14870 8844
rect 14934 8780 15000 8844
rect 10156 8758 15000 8780
rect 10156 8694 10157 8758
rect 10221 8694 10239 8758
rect 10303 8694 10321 8758
rect 10385 8694 10403 8758
rect 10467 8694 10485 8758
rect 10549 8694 10567 8758
rect 10631 8694 10649 8758
rect 10713 8694 10731 8758
rect 10795 8694 10813 8758
rect 10877 8694 10895 8758
rect 10959 8694 10977 8758
rect 11041 8694 11059 8758
rect 11123 8694 11141 8758
rect 11205 8694 11223 8758
rect 11287 8694 11305 8758
rect 11369 8694 11387 8758
rect 11451 8694 11468 8758
rect 11532 8694 11549 8758
rect 11613 8694 11630 8758
rect 11694 8694 11711 8758
rect 11775 8694 11792 8758
rect 11856 8694 11873 8758
rect 11937 8694 11954 8758
rect 12018 8694 12035 8758
rect 12099 8694 12116 8758
rect 12180 8694 12197 8758
rect 12261 8694 12278 8758
rect 12342 8694 12359 8758
rect 12423 8694 12440 8758
rect 12504 8694 12521 8758
rect 12585 8694 12602 8758
rect 12666 8694 12683 8758
rect 12747 8694 12764 8758
rect 12828 8694 12845 8758
rect 12909 8694 12926 8758
rect 12990 8694 13007 8758
rect 13071 8694 13088 8758
rect 13152 8694 13169 8758
rect 13233 8694 13250 8758
rect 13314 8694 13331 8758
rect 13395 8694 13412 8758
rect 13476 8694 13493 8758
rect 13557 8694 13574 8758
rect 13638 8694 13655 8758
rect 13719 8694 13736 8758
rect 13800 8694 13817 8758
rect 13881 8694 13898 8758
rect 13962 8694 13979 8758
rect 14043 8694 14060 8758
rect 14124 8694 14141 8758
rect 14205 8694 14222 8758
rect 14286 8694 14303 8758
rect 14367 8694 14384 8758
rect 14448 8694 14465 8758
rect 14529 8694 14546 8758
rect 14610 8694 14627 8758
rect 14691 8694 14708 8758
rect 14772 8694 14789 8758
rect 14853 8694 14870 8758
rect 14934 8694 15000 8758
rect 10156 8672 15000 8694
rect 10156 8608 10157 8672
rect 10221 8608 10239 8672
rect 10303 8608 10321 8672
rect 10385 8608 10403 8672
rect 10467 8608 10485 8672
rect 10549 8608 10567 8672
rect 10631 8608 10649 8672
rect 10713 8608 10731 8672
rect 10795 8608 10813 8672
rect 10877 8608 10895 8672
rect 10959 8608 10977 8672
rect 11041 8608 11059 8672
rect 11123 8608 11141 8672
rect 11205 8608 11223 8672
rect 11287 8608 11305 8672
rect 11369 8608 11387 8672
rect 11451 8608 11468 8672
rect 11532 8608 11549 8672
rect 11613 8608 11630 8672
rect 11694 8608 11711 8672
rect 11775 8608 11792 8672
rect 11856 8608 11873 8672
rect 11937 8608 11954 8672
rect 12018 8608 12035 8672
rect 12099 8608 12116 8672
rect 12180 8608 12197 8672
rect 12261 8608 12278 8672
rect 12342 8608 12359 8672
rect 12423 8608 12440 8672
rect 12504 8608 12521 8672
rect 12585 8608 12602 8672
rect 12666 8608 12683 8672
rect 12747 8608 12764 8672
rect 12828 8608 12845 8672
rect 12909 8608 12926 8672
rect 12990 8608 13007 8672
rect 13071 8608 13088 8672
rect 13152 8608 13169 8672
rect 13233 8608 13250 8672
rect 13314 8608 13331 8672
rect 13395 8608 13412 8672
rect 13476 8608 13493 8672
rect 13557 8608 13574 8672
rect 13638 8608 13655 8672
rect 13719 8608 13736 8672
rect 13800 8608 13817 8672
rect 13881 8608 13898 8672
rect 13962 8608 13979 8672
rect 14043 8608 14060 8672
rect 14124 8608 14141 8672
rect 14205 8608 14222 8672
rect 14286 8608 14303 8672
rect 14367 8608 14384 8672
rect 14448 8608 14465 8672
rect 14529 8608 14546 8672
rect 14610 8608 14627 8672
rect 14691 8608 14708 8672
rect 14772 8608 14789 8672
rect 14853 8608 14870 8672
rect 14934 8608 15000 8672
rect 10156 8586 15000 8608
rect 10156 8522 10157 8586
rect 10221 8522 10239 8586
rect 10303 8522 10321 8586
rect 10385 8522 10403 8586
rect 10467 8522 10485 8586
rect 10549 8522 10567 8586
rect 10631 8522 10649 8586
rect 10713 8522 10731 8586
rect 10795 8522 10813 8586
rect 10877 8522 10895 8586
rect 10959 8522 10977 8586
rect 11041 8522 11059 8586
rect 11123 8522 11141 8586
rect 11205 8522 11223 8586
rect 11287 8522 11305 8586
rect 11369 8522 11387 8586
rect 11451 8522 11468 8586
rect 11532 8522 11549 8586
rect 11613 8522 11630 8586
rect 11694 8522 11711 8586
rect 11775 8522 11792 8586
rect 11856 8522 11873 8586
rect 11937 8522 11954 8586
rect 12018 8522 12035 8586
rect 12099 8522 12116 8586
rect 12180 8522 12197 8586
rect 12261 8522 12278 8586
rect 12342 8522 12359 8586
rect 12423 8522 12440 8586
rect 12504 8522 12521 8586
rect 12585 8522 12602 8586
rect 12666 8522 12683 8586
rect 12747 8522 12764 8586
rect 12828 8522 12845 8586
rect 12909 8522 12926 8586
rect 12990 8522 13007 8586
rect 13071 8522 13088 8586
rect 13152 8522 13169 8586
rect 13233 8522 13250 8586
rect 13314 8522 13331 8586
rect 13395 8522 13412 8586
rect 13476 8522 13493 8586
rect 13557 8522 13574 8586
rect 13638 8522 13655 8586
rect 13719 8522 13736 8586
rect 13800 8522 13817 8586
rect 13881 8522 13898 8586
rect 13962 8522 13979 8586
rect 14043 8522 14060 8586
rect 14124 8522 14141 8586
rect 14205 8522 14222 8586
rect 14286 8522 14303 8586
rect 14367 8522 14384 8586
rect 14448 8522 14465 8586
rect 14529 8522 14546 8586
rect 14610 8522 14627 8586
rect 14691 8522 14708 8586
rect 14772 8522 14789 8586
rect 14853 8522 14870 8586
rect 14934 8522 15000 8586
rect 10156 8500 15000 8522
rect 10156 8436 10157 8500
rect 10221 8436 10239 8500
rect 10303 8436 10321 8500
rect 10385 8436 10403 8500
rect 10467 8436 10485 8500
rect 10549 8436 10567 8500
rect 10631 8436 10649 8500
rect 10713 8436 10731 8500
rect 10795 8436 10813 8500
rect 10877 8436 10895 8500
rect 10959 8436 10977 8500
rect 11041 8436 11059 8500
rect 11123 8436 11141 8500
rect 11205 8436 11223 8500
rect 11287 8436 11305 8500
rect 11369 8436 11387 8500
rect 11451 8436 11468 8500
rect 11532 8436 11549 8500
rect 11613 8436 11630 8500
rect 11694 8436 11711 8500
rect 11775 8436 11792 8500
rect 11856 8436 11873 8500
rect 11937 8436 11954 8500
rect 12018 8436 12035 8500
rect 12099 8436 12116 8500
rect 12180 8436 12197 8500
rect 12261 8436 12278 8500
rect 12342 8436 12359 8500
rect 12423 8436 12440 8500
rect 12504 8436 12521 8500
rect 12585 8436 12602 8500
rect 12666 8436 12683 8500
rect 12747 8436 12764 8500
rect 12828 8436 12845 8500
rect 12909 8436 12926 8500
rect 12990 8436 13007 8500
rect 13071 8436 13088 8500
rect 13152 8436 13169 8500
rect 13233 8436 13250 8500
rect 13314 8436 13331 8500
rect 13395 8436 13412 8500
rect 13476 8436 13493 8500
rect 13557 8436 13574 8500
rect 13638 8436 13655 8500
rect 13719 8436 13736 8500
rect 13800 8436 13817 8500
rect 13881 8436 13898 8500
rect 13962 8436 13979 8500
rect 14043 8436 14060 8500
rect 14124 8436 14141 8500
rect 14205 8436 14222 8500
rect 14286 8436 14303 8500
rect 14367 8436 14384 8500
rect 14448 8436 14465 8500
rect 14529 8436 14546 8500
rect 14610 8436 14627 8500
rect 14691 8436 14708 8500
rect 14772 8436 14789 8500
rect 14853 8436 14870 8500
rect 14934 8436 15000 8500
rect 10156 8414 15000 8436
rect 10156 8350 10157 8414
rect 10221 8350 10239 8414
rect 10303 8350 10321 8414
rect 10385 8350 10403 8414
rect 10467 8350 10485 8414
rect 10549 8350 10567 8414
rect 10631 8350 10649 8414
rect 10713 8350 10731 8414
rect 10795 8350 10813 8414
rect 10877 8350 10895 8414
rect 10959 8350 10977 8414
rect 11041 8350 11059 8414
rect 11123 8350 11141 8414
rect 11205 8350 11223 8414
rect 11287 8350 11305 8414
rect 11369 8350 11387 8414
rect 11451 8350 11468 8414
rect 11532 8350 11549 8414
rect 11613 8350 11630 8414
rect 11694 8350 11711 8414
rect 11775 8350 11792 8414
rect 11856 8350 11873 8414
rect 11937 8350 11954 8414
rect 12018 8350 12035 8414
rect 12099 8350 12116 8414
rect 12180 8350 12197 8414
rect 12261 8350 12278 8414
rect 12342 8350 12359 8414
rect 12423 8350 12440 8414
rect 12504 8350 12521 8414
rect 12585 8350 12602 8414
rect 12666 8350 12683 8414
rect 12747 8350 12764 8414
rect 12828 8350 12845 8414
rect 12909 8350 12926 8414
rect 12990 8350 13007 8414
rect 13071 8350 13088 8414
rect 13152 8350 13169 8414
rect 13233 8350 13250 8414
rect 13314 8350 13331 8414
rect 13395 8350 13412 8414
rect 13476 8350 13493 8414
rect 13557 8350 13574 8414
rect 13638 8350 13655 8414
rect 13719 8350 13736 8414
rect 13800 8350 13817 8414
rect 13881 8350 13898 8414
rect 13962 8350 13979 8414
rect 14043 8350 14060 8414
rect 14124 8350 14141 8414
rect 14205 8350 14222 8414
rect 14286 8350 14303 8414
rect 14367 8350 14384 8414
rect 14448 8350 14465 8414
rect 14529 8350 14546 8414
rect 14610 8350 14627 8414
rect 14691 8350 14708 8414
rect 14772 8350 14789 8414
rect 14853 8350 14870 8414
rect 14934 8350 15000 8414
rect 10156 8328 15000 8350
rect 10156 8264 10157 8328
rect 10221 8264 10239 8328
rect 10303 8264 10321 8328
rect 10385 8264 10403 8328
rect 10467 8264 10485 8328
rect 10549 8264 10567 8328
rect 10631 8264 10649 8328
rect 10713 8264 10731 8328
rect 10795 8264 10813 8328
rect 10877 8264 10895 8328
rect 10959 8264 10977 8328
rect 11041 8264 11059 8328
rect 11123 8264 11141 8328
rect 11205 8264 11223 8328
rect 11287 8264 11305 8328
rect 11369 8264 11387 8328
rect 11451 8264 11468 8328
rect 11532 8264 11549 8328
rect 11613 8264 11630 8328
rect 11694 8264 11711 8328
rect 11775 8264 11792 8328
rect 11856 8264 11873 8328
rect 11937 8264 11954 8328
rect 12018 8264 12035 8328
rect 12099 8264 12116 8328
rect 12180 8264 12197 8328
rect 12261 8264 12278 8328
rect 12342 8264 12359 8328
rect 12423 8264 12440 8328
rect 12504 8264 12521 8328
rect 12585 8264 12602 8328
rect 12666 8264 12683 8328
rect 12747 8264 12764 8328
rect 12828 8264 12845 8328
rect 12909 8264 12926 8328
rect 12990 8264 13007 8328
rect 13071 8264 13088 8328
rect 13152 8264 13169 8328
rect 13233 8264 13250 8328
rect 13314 8264 13331 8328
rect 13395 8264 13412 8328
rect 13476 8264 13493 8328
rect 13557 8264 13574 8328
rect 13638 8264 13655 8328
rect 13719 8264 13736 8328
rect 13800 8264 13817 8328
rect 13881 8264 13898 8328
rect 13962 8264 13979 8328
rect 14043 8264 14060 8328
rect 14124 8264 14141 8328
rect 14205 8264 14222 8328
rect 14286 8264 14303 8328
rect 14367 8264 14384 8328
rect 14448 8264 14465 8328
rect 14529 8264 14546 8328
rect 14610 8264 14627 8328
rect 14691 8264 14708 8328
rect 14772 8264 14789 8328
rect 14853 8264 14870 8328
rect 14934 8264 15000 8328
rect 10156 8242 15000 8264
rect 10156 8178 10157 8242
rect 10221 8178 10239 8242
rect 10303 8178 10321 8242
rect 10385 8178 10403 8242
rect 10467 8178 10485 8242
rect 10549 8178 10567 8242
rect 10631 8178 10649 8242
rect 10713 8178 10731 8242
rect 10795 8178 10813 8242
rect 10877 8178 10895 8242
rect 10959 8178 10977 8242
rect 11041 8178 11059 8242
rect 11123 8178 11141 8242
rect 11205 8178 11223 8242
rect 11287 8178 11305 8242
rect 11369 8178 11387 8242
rect 11451 8178 11468 8242
rect 11532 8178 11549 8242
rect 11613 8178 11630 8242
rect 11694 8178 11711 8242
rect 11775 8178 11792 8242
rect 11856 8178 11873 8242
rect 11937 8178 11954 8242
rect 12018 8178 12035 8242
rect 12099 8178 12116 8242
rect 12180 8178 12197 8242
rect 12261 8178 12278 8242
rect 12342 8178 12359 8242
rect 12423 8178 12440 8242
rect 12504 8178 12521 8242
rect 12585 8178 12602 8242
rect 12666 8178 12683 8242
rect 12747 8178 12764 8242
rect 12828 8178 12845 8242
rect 12909 8178 12926 8242
rect 12990 8178 13007 8242
rect 13071 8178 13088 8242
rect 13152 8178 13169 8242
rect 13233 8178 13250 8242
rect 13314 8178 13331 8242
rect 13395 8178 13412 8242
rect 13476 8178 13493 8242
rect 13557 8178 13574 8242
rect 13638 8178 13655 8242
rect 13719 8178 13736 8242
rect 13800 8178 13817 8242
rect 13881 8178 13898 8242
rect 13962 8178 13979 8242
rect 14043 8178 14060 8242
rect 14124 8178 14141 8242
rect 14205 8178 14222 8242
rect 14286 8178 14303 8242
rect 14367 8178 14384 8242
rect 14448 8178 14465 8242
rect 14529 8178 14546 8242
rect 14610 8178 14627 8242
rect 14691 8178 14708 8242
rect 14772 8178 14789 8242
rect 14853 8178 14870 8242
rect 14934 8178 15000 8242
rect 10156 8156 15000 8178
rect 10156 8092 10157 8156
rect 10221 8092 10239 8156
rect 10303 8092 10321 8156
rect 10385 8092 10403 8156
rect 10467 8092 10485 8156
rect 10549 8092 10567 8156
rect 10631 8092 10649 8156
rect 10713 8092 10731 8156
rect 10795 8092 10813 8156
rect 10877 8092 10895 8156
rect 10959 8092 10977 8156
rect 11041 8092 11059 8156
rect 11123 8092 11141 8156
rect 11205 8092 11223 8156
rect 11287 8092 11305 8156
rect 11369 8092 11387 8156
rect 11451 8092 11468 8156
rect 11532 8092 11549 8156
rect 11613 8092 11630 8156
rect 11694 8092 11711 8156
rect 11775 8092 11792 8156
rect 11856 8092 11873 8156
rect 11937 8092 11954 8156
rect 12018 8092 12035 8156
rect 12099 8092 12116 8156
rect 12180 8092 12197 8156
rect 12261 8092 12278 8156
rect 12342 8092 12359 8156
rect 12423 8092 12440 8156
rect 12504 8092 12521 8156
rect 12585 8092 12602 8156
rect 12666 8092 12683 8156
rect 12747 8092 12764 8156
rect 12828 8092 12845 8156
rect 12909 8092 12926 8156
rect 12990 8092 13007 8156
rect 13071 8092 13088 8156
rect 13152 8092 13169 8156
rect 13233 8092 13250 8156
rect 13314 8092 13331 8156
rect 13395 8092 13412 8156
rect 13476 8092 13493 8156
rect 13557 8092 13574 8156
rect 13638 8092 13655 8156
rect 13719 8092 13736 8156
rect 13800 8092 13817 8156
rect 13881 8092 13898 8156
rect 13962 8092 13979 8156
rect 14043 8092 14060 8156
rect 14124 8092 14141 8156
rect 14205 8092 14222 8156
rect 14286 8092 14303 8156
rect 14367 8092 14384 8156
rect 14448 8092 14465 8156
rect 14529 8092 14546 8156
rect 14610 8092 14627 8156
rect 14691 8092 14708 8156
rect 14772 8092 14789 8156
rect 14853 8092 14870 8156
rect 14934 8092 15000 8156
rect 10156 8070 15000 8092
rect 10156 8006 10157 8070
rect 10221 8006 10239 8070
rect 10303 8006 10321 8070
rect 10385 8006 10403 8070
rect 10467 8006 10485 8070
rect 10549 8006 10567 8070
rect 10631 8006 10649 8070
rect 10713 8006 10731 8070
rect 10795 8006 10813 8070
rect 10877 8006 10895 8070
rect 10959 8006 10977 8070
rect 11041 8006 11059 8070
rect 11123 8006 11141 8070
rect 11205 8006 11223 8070
rect 11287 8006 11305 8070
rect 11369 8006 11387 8070
rect 11451 8006 11468 8070
rect 11532 8006 11549 8070
rect 11613 8006 11630 8070
rect 11694 8006 11711 8070
rect 11775 8006 11792 8070
rect 11856 8006 11873 8070
rect 11937 8006 11954 8070
rect 12018 8006 12035 8070
rect 12099 8006 12116 8070
rect 12180 8006 12197 8070
rect 12261 8006 12278 8070
rect 12342 8006 12359 8070
rect 12423 8006 12440 8070
rect 12504 8006 12521 8070
rect 12585 8006 12602 8070
rect 12666 8006 12683 8070
rect 12747 8006 12764 8070
rect 12828 8006 12845 8070
rect 12909 8006 12926 8070
rect 12990 8006 13007 8070
rect 13071 8006 13088 8070
rect 13152 8006 13169 8070
rect 13233 8006 13250 8070
rect 13314 8006 13331 8070
rect 13395 8006 13412 8070
rect 13476 8006 13493 8070
rect 13557 8006 13574 8070
rect 13638 8006 13655 8070
rect 13719 8006 13736 8070
rect 13800 8006 13817 8070
rect 13881 8006 13898 8070
rect 13962 8006 13979 8070
rect 14043 8006 14060 8070
rect 14124 8006 14141 8070
rect 14205 8006 14222 8070
rect 14286 8006 14303 8070
rect 14367 8006 14384 8070
rect 14448 8006 14465 8070
rect 14529 8006 14546 8070
rect 14610 8006 14627 8070
rect 14691 8006 14708 8070
rect 14772 8006 14789 8070
rect 14853 8006 14870 8070
rect 14934 8006 15000 8070
rect 10156 7984 15000 8006
rect 10156 7920 10157 7984
rect 10221 7920 10239 7984
rect 10303 7920 10321 7984
rect 10385 7920 10403 7984
rect 10467 7920 10485 7984
rect 10549 7920 10567 7984
rect 10631 7920 10649 7984
rect 10713 7920 10731 7984
rect 10795 7920 10813 7984
rect 10877 7920 10895 7984
rect 10959 7920 10977 7984
rect 11041 7920 11059 7984
rect 11123 7920 11141 7984
rect 11205 7920 11223 7984
rect 11287 7920 11305 7984
rect 11369 7920 11387 7984
rect 11451 7920 11468 7984
rect 11532 7920 11549 7984
rect 11613 7920 11630 7984
rect 11694 7920 11711 7984
rect 11775 7920 11792 7984
rect 11856 7920 11873 7984
rect 11937 7920 11954 7984
rect 12018 7920 12035 7984
rect 12099 7920 12116 7984
rect 12180 7920 12197 7984
rect 12261 7920 12278 7984
rect 12342 7920 12359 7984
rect 12423 7920 12440 7984
rect 12504 7920 12521 7984
rect 12585 7920 12602 7984
rect 12666 7920 12683 7984
rect 12747 7920 12764 7984
rect 12828 7920 12845 7984
rect 12909 7920 12926 7984
rect 12990 7920 13007 7984
rect 13071 7920 13088 7984
rect 13152 7920 13169 7984
rect 13233 7920 13250 7984
rect 13314 7920 13331 7984
rect 13395 7920 13412 7984
rect 13476 7920 13493 7984
rect 13557 7920 13574 7984
rect 13638 7920 13655 7984
rect 13719 7920 13736 7984
rect 13800 7920 13817 7984
rect 13881 7920 13898 7984
rect 13962 7920 13979 7984
rect 14043 7920 14060 7984
rect 14124 7920 14141 7984
rect 14205 7920 14222 7984
rect 14286 7920 14303 7984
rect 14367 7920 14384 7984
rect 14448 7920 14465 7984
rect 14529 7920 14546 7984
rect 14610 7920 14627 7984
rect 14691 7920 14708 7984
rect 14772 7920 14789 7984
rect 14853 7920 14870 7984
rect 14934 7920 15000 7984
rect 10156 7917 15000 7920
rect 0 6947 254 7637
rect 14746 6947 15000 7637
rect 0 5977 254 6667
rect 14746 5977 15000 6667
rect 0 4767 254 5697
rect 14746 4767 15000 5697
rect 0 3557 254 4487
rect 14746 3557 15000 4487
rect 0 2587 193 3277
rect 14807 2587 15000 3277
rect 0 1377 254 2307
rect 14746 1377 15000 2307
rect 0 7 254 1097
rect 14746 7 15000 1097
<< metal5 >>
rect 0 34757 254 39600
rect 14746 34757 15000 39600
rect 0 13607 254 18597
rect 14746 13607 15000 18597
rect 0 12437 254 13287
rect 14746 12437 15000 13287
rect 0 11267 254 12117
rect 14746 11267 15000 12117
rect 0 9147 254 10947
rect 14746 9147 15000 10947
rect 0 7937 254 8827
rect 14746 7937 15000 8827
rect 0 6968 254 7617
rect 14746 6968 15000 7617
rect 0 5997 254 6647
rect 14746 5997 15000 6647
rect 0 4787 254 5677
rect 14746 4787 15000 5677
rect 0 3577 254 4467
rect 14746 3577 15000 4467
rect 0 2607 193 3257
rect 14807 2607 15000 3257
rect 0 1397 254 2287
rect 14746 1397 15000 2287
rect 0 27 254 1077
rect 14746 27 15000 1077
use sky130_fd_io__com_bus_hookup  sky130_fd_io__com_bus_hookup_0
timestamp 1649977179
transform 1 0 0 0 1 149
box 0 -142 15000 39451
<< labels >>
flabel metal5 s 0 9147 254 10947 3 FreeSans 520 0 0 0 VSSA
port 1 nsew ground bidirectional
flabel metal5 s 0 13607 254 18597 3 FreeSans 520 0 0 0 VDDIO
port 2 nsew power bidirectional
flabel metal5 s 0 12437 254 13287 3 FreeSans 520 0 0 0 VDDIO_Q
port 3 nsew power bidirectional
flabel metal5 s 0 6968 254 7617 3 FreeSans 520 0 0 0 VSSA
port 1 nsew ground bidirectional
flabel metal5 s 0 7937 254 8827 3 FreeSans 520 0 0 0 VSSD
port 4 nsew ground bidirectional
flabel metal5 s 0 4787 254 5677 3 FreeSans 520 0 0 0 VSSIO
port 5 nsew ground bidirectional
flabel metal5 s 0 5997 254 6647 3 FreeSans 520 0 0 0 VSWITCH
port 6 nsew power bidirectional
flabel metal5 s 0 11267 254 12117 3 FreeSans 520 0 0 0 VSSIO_Q
port 7 nsew ground bidirectional
flabel metal5 s 0 3577 254 4467 3 FreeSans 520 0 0 0 VDDIO
port 2 nsew power bidirectional
flabel metal5 s 0 2607 193 3257 3 FreeSans 520 0 0 0 VDDA
port 8 nsew power bidirectional
flabel metal5 s 0 1397 254 2287 3 FreeSans 520 0 0 0 VCCD
port 9 nsew power bidirectional
flabel metal5 s 0 27 254 1077 3 FreeSans 520 0 0 0 VCCHIB
port 10 nsew power bidirectional
flabel metal5 s 14746 9147 15000 10947 3 FreeSans 520 180 0 0 VSSA
port 1 nsew ground bidirectional
flabel metal5 s 14746 13607 15000 18597 3 FreeSans 520 180 0 0 VDDIO
port 2 nsew power bidirectional
flabel metal5 s 14746 12437 15000 13287 3 FreeSans 520 180 0 0 VDDIO_Q
port 3 nsew power bidirectional
flabel metal5 s 14746 6968 15000 7617 3 FreeSans 520 180 0 0 VSSA
port 1 nsew ground bidirectional
flabel metal5 s 14746 7937 15000 8827 3 FreeSans 520 180 0 0 VSSD
port 4 nsew ground bidirectional
flabel metal5 s 14746 4787 15000 5677 3 FreeSans 520 180 0 0 VSSIO
port 5 nsew ground bidirectional
flabel metal5 s 14746 5997 15000 6647 3 FreeSans 520 180 0 0 VSWITCH
port 6 nsew power bidirectional
flabel metal5 s 14746 11267 15000 12117 3 FreeSans 520 180 0 0 VSSIO_Q
port 7 nsew ground bidirectional
flabel metal5 s 14746 3577 15000 4467 3 FreeSans 520 180 0 0 VDDIO
port 2 nsew power bidirectional
flabel metal5 s 14807 2607 15000 3257 3 FreeSans 520 180 0 0 VDDA
port 8 nsew power bidirectional
flabel metal5 s 14746 1397 15000 2287 3 FreeSans 520 180 0 0 VCCD
port 9 nsew power bidirectional
flabel metal5 s 14746 27 15000 1077 3 FreeSans 520 180 0 0 VCCHIB
port 10 nsew power bidirectional
flabel metal5 s 14746 34757 15000 39600 3 FreeSans 520 180 0 0 VSSIO
port 5 nsew ground bidirectional
flabel metal5 s 0 34757 254 39600 3 FreeSans 520 0 0 0 VSSIO
port 5 nsew ground bidirectional
flabel metal4 s 0 3557 254 4487 3 FreeSans 520 0 0 0 VDDIO
port 2 nsew power bidirectional
flabel metal4 s 0 10881 254 10947 3 FreeSans 520 0 0 0 VSSA
port 1 nsew ground bidirectional
flabel metal4 s 0 5977 254 6667 3 FreeSans 520 0 0 0 VSWITCH
port 6 nsew power bidirectional
flabel metal4 s 0 4767 254 5697 3 FreeSans 520 0 0 0 VSSIO
port 5 nsew ground bidirectional
flabel metal4 s 0 11247 254 12137 3 FreeSans 520 0 0 0 VSSIO_Q
port 7 nsew ground bidirectional
flabel metal4 s 0 9147 254 9213 3 FreeSans 520 0 0 0 VSSA
port 1 nsew ground bidirectional
flabel metal4 s 0 9929 254 10165 3 FreeSans 520 0 0 0 VSSA
port 1 nsew ground bidirectional
flabel metal4 s 0 2587 193 3277 3 FreeSans 520 0 0 0 VDDA
port 8 nsew power bidirectional
flabel metal4 s 0 1377 254 2307 3 FreeSans 520 0 0 0 VCCD
port 9 nsew power bidirectional
flabel metal4 s 0 7 254 1097 3 FreeSans 520 0 0 0 VCCHIB
port 10 nsew power bidirectional
flabel metal4 s 0 9273 254 9869 3 FreeSans 520 0 0 0 AMUXBUS_B
port 11 nsew signal bidirectional
flabel metal4 s 0 12417 254 13307 3 FreeSans 520 0 0 0 VDDIO_Q
port 3 nsew power bidirectional
flabel metal4 s 0 7917 254 8847 3 FreeSans 520 0 0 0 VSSD
port 4 nsew ground bidirectional
flabel metal4 s 0 6947 254 7637 3 FreeSans 520 0 0 0 VSSA
port 1 nsew ground bidirectional
flabel metal4 s 0 10225 254 10821 3 FreeSans 520 0 0 0 AMUXBUS_A
port 12 nsew signal bidirectional
flabel metal4 s 0 13607 254 18600 3 FreeSans 520 0 0 0 VDDIO
port 2 nsew power bidirectional
flabel metal4 s 14746 3557 15000 4487 3 FreeSans 520 180 0 0 VDDIO
port 2 nsew power bidirectional
flabel metal4 s 14746 10881 15000 10947 3 FreeSans 520 180 0 0 VSSA
port 1 nsew ground bidirectional
flabel metal4 s 14746 5977 15000 6667 3 FreeSans 520 180 0 0 VSWITCH
port 6 nsew power bidirectional
flabel metal4 s 14746 4767 15000 5697 3 FreeSans 520 180 0 0 VSSIO
port 5 nsew ground bidirectional
flabel metal4 s 14746 11247 15000 12137 3 FreeSans 520 180 0 0 VSSIO_Q
port 7 nsew ground bidirectional
flabel metal4 s 14746 9147 15000 9213 3 FreeSans 520 180 0 0 VSSA
port 1 nsew ground bidirectional
flabel metal4 s 14746 9929 15000 10165 3 FreeSans 520 180 0 0 VSSA
port 1 nsew ground bidirectional
flabel metal4 s 14807 2587 15000 3277 3 FreeSans 520 180 0 0 VDDA
port 8 nsew power bidirectional
flabel metal4 s 14746 1377 15000 2307 3 FreeSans 520 180 0 0 VCCD
port 9 nsew power bidirectional
flabel metal4 s 14746 7 15000 1097 3 FreeSans 520 180 0 0 VCCHIB
port 10 nsew power bidirectional
flabel metal4 s 14746 9273 15000 9869 3 FreeSans 520 180 0 0 AMUXBUS_B
port 11 nsew signal bidirectional
flabel metal4 s 14746 12417 15000 13307 3 FreeSans 520 180 0 0 VDDIO_Q
port 3 nsew power bidirectional
flabel metal4 s 14746 7917 15000 8847 3 FreeSans 520 180 0 0 VSSD
port 4 nsew ground bidirectional
flabel metal4 s 14746 6947 15000 7637 3 FreeSans 520 180 0 0 VSSA
port 1 nsew ground bidirectional
flabel metal4 s 14746 10225 15000 10821 3 FreeSans 520 180 0 0 AMUXBUS_A
port 12 nsew signal bidirectional
flabel metal4 s 14746 13607 15000 18600 3 FreeSans 520 180 0 0 VDDIO
port 2 nsew power bidirectional
flabel metal4 s 14746 34757 15000 39600 3 FreeSans 520 180 0 0 VSSIO
port 5 nsew ground bidirectional
flabel metal4 s 14873 37932 14873 37932 3 FreeSans 520 180 0 0 VSSIO
port 5 nsew
flabel metal4 s 0 34757 254 39600 3 FreeSans 520 0 0 0 VSSIO
port 5 nsew ground bidirectional
flabel metal4 s 127 37932 127 37932 3 FreeSans 520 0 0 0 VSSIO
port 5 nsew
rlabel metal4 s 14746 10225 15000 10821 1 AMUXBUS_A
port 12 nsew signal bidirectional
rlabel metal4 s 14746 9273 15000 9869 1 AMUXBUS_B
port 11 nsew signal bidirectional
rlabel metal4 s 14746 1377 15000 2307 1 VCCD
port 9 nsew power bidirectional
rlabel metal5 s 0 1397 254 2287 1 VCCD
port 9 nsew power bidirectional
rlabel metal5 s 14746 1397 15000 2287 1 VCCD
port 9 nsew power bidirectional
rlabel metal4 s 14746 7 15000 1097 1 VCCHIB
port 10 nsew power bidirectional
rlabel metal5 s 0 27 254 1077 1 VCCHIB
port 10 nsew power bidirectional
rlabel metal5 s 14746 27 15000 1077 1 VCCHIB
port 10 nsew power bidirectional
rlabel metal4 s 14807 2587 15000 3277 1 VDDA
port 8 nsew power bidirectional
rlabel metal5 s 0 2607 193 3257 1 VDDA
port 8 nsew power bidirectional
rlabel metal5 s 14807 2607 15000 3257 1 VDDA
port 8 nsew power bidirectional
rlabel metal4 s 0 13607 254 18600 1 VDDIO
port 2 nsew power bidirectional
rlabel metal4 s 14746 3557 15000 4487 1 VDDIO
port 2 nsew power bidirectional
rlabel metal4 s 14746 13607 15000 18600 1 VDDIO
port 2 nsew power bidirectional
rlabel metal5 s 0 3577 254 4467 1 VDDIO
port 2 nsew power bidirectional
rlabel metal5 s 0 13607 254 18597 1 VDDIO
port 2 nsew power bidirectional
rlabel metal5 s 14746 3577 15000 4467 1 VDDIO
port 2 nsew power bidirectional
rlabel metal5 s 14746 13607 15000 18597 1 VDDIO
port 2 nsew power bidirectional
rlabel metal4 s 14746 12417 15000 13307 1 VDDIO_Q
port 3 nsew power bidirectional
rlabel metal5 s 0 12437 254 13287 1 VDDIO_Q
port 3 nsew power bidirectional
rlabel metal5 s 14746 12437 15000 13287 1 VDDIO_Q
port 3 nsew power bidirectional
rlabel metal4 s 0 9147 254 9213 1 VSSA
port 1 nsew ground bidirectional
rlabel metal4 s 0 9929 254 10165 1 VSSA
port 1 nsew ground bidirectional
rlabel metal4 s 0 10881 254 10947 1 VSSA
port 1 nsew ground bidirectional
rlabel metal4 s 14746 6947 15000 7637 1 VSSA
port 1 nsew ground bidirectional
rlabel metal4 s 14746 9147 15000 9213 1 VSSA
port 1 nsew ground bidirectional
rlabel metal4 s 14746 9929 15000 10165 1 VSSA
port 1 nsew ground bidirectional
rlabel metal4 s 14746 10881 15000 10947 1 VSSA
port 1 nsew ground bidirectional
rlabel metal5 s 0 6968 254 7617 1 VSSA
port 1 nsew ground bidirectional
rlabel metal5 s 0 9147 254 10947 1 VSSA
port 1 nsew ground bidirectional
rlabel metal5 s 14746 6968 15000 7617 1 VSSA
port 1 nsew ground bidirectional
rlabel metal5 s 14746 9147 15000 10947 1 VSSA
port 1 nsew ground bidirectional
rlabel metal3 s 10151 7918 14940 8846 1 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 0 7917 4895 8847 1 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 10156 7917 15000 8847 1 VSSD
port 4 nsew ground bidirectional
rlabel metal5 s 0 7937 254 8827 1 VSSD
port 4 nsew ground bidirectional
rlabel metal5 s 14746 7937 15000 8827 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 14882 8792 14922 8832 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 14882 8706 14922 8746 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 14882 8620 14922 8660 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 14882 8534 14922 8574 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 14882 8448 14922 8488 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 14882 8362 14922 8402 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 14882 8276 14922 8316 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 14882 8190 14922 8230 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 14882 8104 14922 8144 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 14882 8018 14922 8058 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 14882 7932 14922 7972 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 14801 8792 14841 8832 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 14801 8706 14841 8746 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 14801 8620 14841 8660 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 14801 8534 14841 8574 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 14801 8448 14841 8488 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 14801 8362 14841 8402 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 14801 8276 14841 8316 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 14801 8190 14841 8230 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 14801 8104 14841 8144 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 14801 8018 14841 8058 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 14801 7932 14841 7972 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 14720 8792 14760 8832 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 14720 8706 14760 8746 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 14720 8620 14760 8660 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 14720 8534 14760 8574 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 14720 8448 14760 8488 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 14720 8362 14760 8402 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 14720 8276 14760 8316 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 14720 8190 14760 8230 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 14720 8104 14760 8144 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 14720 8018 14760 8058 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 14720 7932 14760 7972 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 14639 8792 14679 8832 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 14639 8706 14679 8746 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 14639 8620 14679 8660 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 14639 8534 14679 8574 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 14639 8448 14679 8488 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 14639 8362 14679 8402 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 14639 8276 14679 8316 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 14639 8190 14679 8230 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 14639 8104 14679 8144 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 14639 8018 14679 8058 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 14639 7932 14679 7972 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 14558 8792 14598 8832 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 14558 8706 14598 8746 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 14558 8620 14598 8660 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 14558 8534 14598 8574 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 14558 8448 14598 8488 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 14558 8362 14598 8402 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 14558 8276 14598 8316 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 14558 8190 14598 8230 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 14558 8104 14598 8144 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 14558 8018 14598 8058 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 14558 7932 14598 7972 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 14477 8792 14517 8832 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 14477 8706 14517 8746 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 14477 8620 14517 8660 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 14477 8534 14517 8574 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 14477 8448 14517 8488 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 14477 8362 14517 8402 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 14477 8276 14517 8316 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 14477 8190 14517 8230 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 14477 8104 14517 8144 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 14477 8018 14517 8058 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 14477 7932 14517 7972 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 14396 8792 14436 8832 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 14396 8706 14436 8746 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 14396 8620 14436 8660 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 14396 8534 14436 8574 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 14396 8448 14436 8488 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 14396 8362 14436 8402 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 14396 8276 14436 8316 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 14396 8190 14436 8230 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 14396 8104 14436 8144 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 14396 8018 14436 8058 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 14396 7932 14436 7972 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 14315 8792 14355 8832 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 14315 8706 14355 8746 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 14315 8620 14355 8660 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 14315 8534 14355 8574 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 14315 8448 14355 8488 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 14315 8362 14355 8402 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 14315 8276 14355 8316 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 14315 8190 14355 8230 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 14315 8104 14355 8144 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 14315 8018 14355 8058 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 14315 7932 14355 7972 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 14234 8792 14274 8832 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 14234 8706 14274 8746 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 14234 8620 14274 8660 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 14234 8534 14274 8574 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 14234 8448 14274 8488 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 14234 8362 14274 8402 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 14234 8276 14274 8316 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 14234 8190 14274 8230 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 14234 8104 14274 8144 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 14234 8018 14274 8058 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 14234 7932 14274 7972 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 14153 8792 14193 8832 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 14153 8706 14193 8746 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 14153 8620 14193 8660 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 14153 8534 14193 8574 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 14153 8448 14193 8488 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 14153 8362 14193 8402 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 14153 8276 14193 8316 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 14153 8190 14193 8230 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 14153 8104 14193 8144 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 14153 8018 14193 8058 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 14153 7932 14193 7972 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 14072 8792 14112 8832 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 14072 8706 14112 8746 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 14072 8620 14112 8660 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 14072 8534 14112 8574 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 14072 8448 14112 8488 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 14072 8362 14112 8402 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 14072 8276 14112 8316 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 14072 8190 14112 8230 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 14072 8104 14112 8144 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 14072 8018 14112 8058 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 14072 7932 14112 7972 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13991 8792 14031 8832 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13991 8706 14031 8746 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13991 8620 14031 8660 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13991 8534 14031 8574 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13991 8448 14031 8488 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13991 8362 14031 8402 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13991 8276 14031 8316 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13991 8190 14031 8230 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13991 8104 14031 8144 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13991 8018 14031 8058 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13991 7932 14031 7972 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13910 8792 13950 8832 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13910 8706 13950 8746 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13910 8620 13950 8660 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13910 8534 13950 8574 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13910 8448 13950 8488 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13910 8362 13950 8402 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13910 8276 13950 8316 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13910 8190 13950 8230 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13910 8104 13950 8144 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13910 8018 13950 8058 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13910 7932 13950 7972 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13829 8792 13869 8832 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13829 8706 13869 8746 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13829 8620 13869 8660 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13829 8534 13869 8574 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13829 8448 13869 8488 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13829 8362 13869 8402 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13829 8276 13869 8316 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13829 8190 13869 8230 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13829 8104 13869 8144 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13829 8018 13869 8058 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13829 7932 13869 7972 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13748 8792 13788 8832 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13748 8706 13788 8746 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13748 8620 13788 8660 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13748 8534 13788 8574 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13748 8448 13788 8488 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13748 8362 13788 8402 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13748 8276 13788 8316 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13748 8190 13788 8230 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13748 8104 13788 8144 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13748 8018 13788 8058 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13748 7932 13788 7972 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13667 8792 13707 8832 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13667 8706 13707 8746 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13667 8620 13707 8660 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13667 8534 13707 8574 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13667 8448 13707 8488 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13667 8362 13707 8402 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13667 8276 13707 8316 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13667 8190 13707 8230 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13667 8104 13707 8144 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13667 8018 13707 8058 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13667 7932 13707 7972 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13586 8792 13626 8832 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13586 8706 13626 8746 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13586 8620 13626 8660 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13586 8534 13626 8574 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13586 8448 13626 8488 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13586 8362 13626 8402 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13586 8276 13626 8316 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13586 8190 13626 8230 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13586 8104 13626 8144 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13586 8018 13626 8058 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13586 7932 13626 7972 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13505 8792 13545 8832 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13505 8706 13545 8746 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13505 8620 13545 8660 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13505 8534 13545 8574 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13505 8448 13545 8488 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13505 8362 13545 8402 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13505 8276 13545 8316 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13505 8190 13545 8230 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13505 8104 13545 8144 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13505 8018 13545 8058 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13505 7932 13545 7972 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13424 8792 13464 8832 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13424 8706 13464 8746 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13424 8620 13464 8660 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13424 8534 13464 8574 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13424 8448 13464 8488 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13424 8362 13464 8402 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13424 8276 13464 8316 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13424 8190 13464 8230 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13424 8104 13464 8144 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13424 8018 13464 8058 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13424 7932 13464 7972 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13343 8792 13383 8832 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13343 8706 13383 8746 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13343 8620 13383 8660 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13343 8534 13383 8574 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13343 8448 13383 8488 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13343 8362 13383 8402 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13343 8276 13383 8316 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13343 8190 13383 8230 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13343 8104 13383 8144 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13343 8018 13383 8058 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13343 7932 13383 7972 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13262 8792 13302 8832 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13262 8706 13302 8746 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13262 8620 13302 8660 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13262 8534 13302 8574 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13262 8448 13302 8488 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13262 8362 13302 8402 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13262 8276 13302 8316 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13262 8190 13302 8230 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13262 8104 13302 8144 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13262 8018 13302 8058 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13262 7932 13302 7972 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13181 8792 13221 8832 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13181 8706 13221 8746 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13181 8620 13221 8660 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13181 8534 13221 8574 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13181 8448 13221 8488 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13181 8362 13221 8402 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13181 8276 13221 8316 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13181 8190 13221 8230 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13181 8104 13221 8144 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13181 8018 13221 8058 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13181 7932 13221 7972 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13100 8792 13140 8832 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13100 8706 13140 8746 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13100 8620 13140 8660 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13100 8534 13140 8574 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13100 8448 13140 8488 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13100 8362 13140 8402 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13100 8276 13140 8316 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13100 8190 13140 8230 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13100 8104 13140 8144 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13100 8018 13140 8058 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13100 7932 13140 7972 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13019 8792 13059 8832 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13019 8706 13059 8746 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13019 8620 13059 8660 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13019 8534 13059 8574 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13019 8448 13059 8488 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13019 8362 13059 8402 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13019 8276 13059 8316 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13019 8190 13059 8230 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13019 8104 13059 8144 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13019 8018 13059 8058 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 13019 7932 13059 7972 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 12938 8792 12978 8832 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 12938 8706 12978 8746 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 12938 8620 12978 8660 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 12938 8534 12978 8574 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 12938 8448 12978 8488 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 12938 8362 12978 8402 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 12938 8276 12978 8316 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 12938 8190 12978 8230 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 12938 8104 12978 8144 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 12938 8018 12978 8058 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 12938 7932 12978 7972 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 12857 8792 12897 8832 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 12857 8706 12897 8746 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 12857 8620 12897 8660 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 12857 8534 12897 8574 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 12857 8448 12897 8488 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 12857 8362 12897 8402 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 12857 8276 12897 8316 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 12857 8190 12897 8230 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 12857 8104 12897 8144 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 12857 8018 12897 8058 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 12857 7932 12897 7972 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 12776 8792 12816 8832 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 12776 8706 12816 8746 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 12776 8620 12816 8660 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 12776 8534 12816 8574 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 12776 8448 12816 8488 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 12776 8362 12816 8402 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 12776 8276 12816 8316 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 12776 8190 12816 8230 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 12776 8104 12816 8144 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 12776 8018 12816 8058 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 12776 7932 12816 7972 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 12695 8792 12735 8832 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 12695 8706 12735 8746 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 12695 8620 12735 8660 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 12695 8534 12735 8574 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 12695 8448 12735 8488 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 12695 8362 12735 8402 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 12695 8276 12735 8316 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 12695 8190 12735 8230 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 12695 8104 12735 8144 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 12695 8018 12735 8058 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 12695 7932 12735 7972 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 12614 8792 12654 8832 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 12614 8706 12654 8746 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 12614 8620 12654 8660 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 12614 8534 12654 8574 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 12614 8448 12654 8488 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 12614 8362 12654 8402 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 12614 8276 12654 8316 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 12614 8190 12654 8230 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 12614 8104 12654 8144 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 12614 8018 12654 8058 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 12614 7932 12654 7972 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 12533 8792 12573 8832 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 12533 8706 12573 8746 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 12533 8620 12573 8660 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 12533 8534 12573 8574 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 12533 8448 12573 8488 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 12533 8362 12573 8402 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 12533 8276 12573 8316 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 12533 8190 12573 8230 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 12533 8104 12573 8144 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 12533 8018 12573 8058 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 12533 7932 12573 7972 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 12452 8792 12492 8832 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 12452 8706 12492 8746 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 12452 8620 12492 8660 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 12452 8534 12492 8574 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 12452 8448 12492 8488 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 12452 8362 12492 8402 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 12452 8276 12492 8316 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 12452 8190 12492 8230 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 12452 8104 12492 8144 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 12452 8018 12492 8058 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 12452 7932 12492 7972 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 12371 8792 12411 8832 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 12371 8706 12411 8746 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 12371 8620 12411 8660 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 12371 8534 12411 8574 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 12371 8448 12411 8488 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 12371 8362 12411 8402 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 12371 8276 12411 8316 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 12371 8190 12411 8230 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 12371 8104 12411 8144 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 12371 8018 12411 8058 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 12371 7932 12411 7972 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 12290 8792 12330 8832 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 12290 8706 12330 8746 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 12290 8620 12330 8660 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 12290 8534 12330 8574 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 12290 8448 12330 8488 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 12290 8362 12330 8402 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 12290 8276 12330 8316 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 12290 8190 12330 8230 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 12290 8104 12330 8144 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 12290 8018 12330 8058 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 12290 7932 12330 7972 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 12209 8792 12249 8832 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 12209 8706 12249 8746 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 12209 8620 12249 8660 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 12209 8534 12249 8574 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 12209 8448 12249 8488 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 12209 8362 12249 8402 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 12209 8276 12249 8316 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 12209 8190 12249 8230 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 12209 8104 12249 8144 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 12209 8018 12249 8058 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 12209 7932 12249 7972 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 12128 8792 12168 8832 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 12128 8706 12168 8746 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 12128 8620 12168 8660 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 12128 8534 12168 8574 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 12128 8448 12168 8488 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 12128 8362 12168 8402 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 12128 8276 12168 8316 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 12128 8190 12168 8230 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 12128 8104 12168 8144 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 12128 8018 12168 8058 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 12128 7932 12168 7972 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 12047 8792 12087 8832 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 12047 8706 12087 8746 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 12047 8620 12087 8660 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 12047 8534 12087 8574 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 12047 8448 12087 8488 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 12047 8362 12087 8402 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 12047 8276 12087 8316 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 12047 8190 12087 8230 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 12047 8104 12087 8144 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 12047 8018 12087 8058 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 12047 7932 12087 7972 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 11966 8792 12006 8832 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 11966 8706 12006 8746 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 11966 8620 12006 8660 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 11966 8534 12006 8574 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 11966 8448 12006 8488 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 11966 8362 12006 8402 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 11966 8276 12006 8316 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 11966 8190 12006 8230 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 11966 8104 12006 8144 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 11966 8018 12006 8058 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 11966 7932 12006 7972 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 11885 8792 11925 8832 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 11885 8706 11925 8746 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 11885 8620 11925 8660 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 11885 8534 11925 8574 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 11885 8448 11925 8488 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 11885 8362 11925 8402 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 11885 8276 11925 8316 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 11885 8190 11925 8230 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 11885 8104 11925 8144 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 11885 8018 11925 8058 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 11885 7932 11925 7972 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 11804 8792 11844 8832 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 11804 8706 11844 8746 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 11804 8620 11844 8660 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 11804 8534 11844 8574 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 11804 8448 11844 8488 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 11804 8362 11844 8402 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 11804 8276 11844 8316 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 11804 8190 11844 8230 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 11804 8104 11844 8144 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 11804 8018 11844 8058 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 11804 7932 11844 7972 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 11723 8792 11763 8832 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 11723 8706 11763 8746 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 11723 8620 11763 8660 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 11723 8534 11763 8574 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 11723 8448 11763 8488 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 11723 8362 11763 8402 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 11723 8276 11763 8316 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 11723 8190 11763 8230 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 11723 8104 11763 8144 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 11723 8018 11763 8058 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 11723 7932 11763 7972 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 11642 8792 11682 8832 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 11642 8706 11682 8746 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 11642 8620 11682 8660 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 11642 8534 11682 8574 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 11642 8448 11682 8488 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 11642 8362 11682 8402 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 11642 8276 11682 8316 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 11642 8190 11682 8230 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 11642 8104 11682 8144 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 11642 8018 11682 8058 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 11642 7932 11682 7972 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 11561 8792 11601 8832 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 11561 8706 11601 8746 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 11561 8620 11601 8660 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 11561 8534 11601 8574 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 11561 8448 11601 8488 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 11561 8362 11601 8402 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 11561 8276 11601 8316 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 11561 8190 11601 8230 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 11561 8104 11601 8144 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 11561 8018 11601 8058 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 11561 7932 11601 7972 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 11480 8792 11520 8832 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 11480 8706 11520 8746 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 11480 8620 11520 8660 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 11480 8534 11520 8574 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 11480 8448 11520 8488 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 11480 8362 11520 8402 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 11480 8276 11520 8316 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 11480 8190 11520 8230 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 11480 8104 11520 8144 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 11480 8018 11520 8058 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 11480 7932 11520 7972 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 11399 8792 11439 8832 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 11399 8706 11439 8746 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 11399 8620 11439 8660 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 11399 8534 11439 8574 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 11399 8448 11439 8488 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 11399 8362 11439 8402 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 11399 8276 11439 8316 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 11399 8190 11439 8230 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 11399 8104 11439 8144 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 11399 8018 11439 8058 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 11399 7932 11439 7972 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 11317 8792 11357 8832 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 11317 8706 11357 8746 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 11317 8620 11357 8660 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 11317 8534 11357 8574 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 11317 8448 11357 8488 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 11317 8362 11357 8402 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 11317 8276 11357 8316 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 11317 8190 11357 8230 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 11317 8104 11357 8144 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 11317 8018 11357 8058 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 11317 7932 11357 7972 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 11235 8792 11275 8832 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 11235 8706 11275 8746 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 11235 8620 11275 8660 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 11235 8534 11275 8574 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 11235 8448 11275 8488 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 11235 8362 11275 8402 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 11235 8276 11275 8316 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 11235 8190 11275 8230 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 11235 8104 11275 8144 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 11235 8018 11275 8058 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 11235 7932 11275 7972 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 11153 8792 11193 8832 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 11153 8706 11193 8746 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 11153 8620 11193 8660 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 11153 8534 11193 8574 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 11153 8448 11193 8488 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 11153 8362 11193 8402 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 11153 8276 11193 8316 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 11153 8190 11193 8230 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 11153 8104 11193 8144 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 11153 8018 11193 8058 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 11153 7932 11193 7972 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 11071 8792 11111 8832 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 11071 8706 11111 8746 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 11071 8620 11111 8660 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 11071 8534 11111 8574 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 11071 8448 11111 8488 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 11071 8362 11111 8402 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 11071 8276 11111 8316 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 11071 8190 11111 8230 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 11071 8104 11111 8144 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 11071 8018 11111 8058 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 11071 7932 11111 7972 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 10989 8792 11029 8832 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 10989 8706 11029 8746 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 10989 8620 11029 8660 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 10989 8534 11029 8574 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 10989 8448 11029 8488 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 10989 8362 11029 8402 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 10989 8276 11029 8316 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 10989 8190 11029 8230 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 10989 8104 11029 8144 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 10989 8018 11029 8058 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 10989 7932 11029 7972 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 10907 8792 10947 8832 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 10907 8706 10947 8746 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 10907 8620 10947 8660 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 10907 8534 10947 8574 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 10907 8448 10947 8488 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 10907 8362 10947 8402 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 10907 8276 10947 8316 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 10907 8190 10947 8230 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 10907 8104 10947 8144 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 10907 8018 10947 8058 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 10907 7932 10947 7972 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 10825 8792 10865 8832 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 10825 8706 10865 8746 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 10825 8620 10865 8660 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 10825 8534 10865 8574 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 10825 8448 10865 8488 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 10825 8362 10865 8402 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 10825 8276 10865 8316 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 10825 8190 10865 8230 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 10825 8104 10865 8144 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 10825 8018 10865 8058 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 10825 7932 10865 7972 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 10743 8792 10783 8832 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 10743 8706 10783 8746 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 10743 8620 10783 8660 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 10743 8534 10783 8574 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 10743 8448 10783 8488 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 10743 8362 10783 8402 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 10743 8276 10783 8316 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 10743 8190 10783 8230 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 10743 8104 10783 8144 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 10743 8018 10783 8058 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 10743 7932 10783 7972 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 10661 8792 10701 8832 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 10661 8706 10701 8746 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 10661 8620 10701 8660 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 10661 8534 10701 8574 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 10661 8448 10701 8488 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 10661 8362 10701 8402 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 10661 8276 10701 8316 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 10661 8190 10701 8230 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 10661 8104 10701 8144 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 10661 8018 10701 8058 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 10661 7932 10701 7972 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 10579 8792 10619 8832 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 10579 8706 10619 8746 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 10579 8620 10619 8660 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 10579 8534 10619 8574 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 10579 8448 10619 8488 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 10579 8362 10619 8402 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 10579 8276 10619 8316 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 10579 8190 10619 8230 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 10579 8104 10619 8144 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 10579 8018 10619 8058 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 10579 7932 10619 7972 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 10497 8792 10537 8832 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 10497 8706 10537 8746 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 10497 8620 10537 8660 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 10497 8534 10537 8574 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 10497 8448 10537 8488 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 10497 8362 10537 8402 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 10497 8276 10537 8316 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 10497 8190 10537 8230 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 10497 8104 10537 8144 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 10497 8018 10537 8058 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 10497 7932 10537 7972 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 10415 8792 10455 8832 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 10415 8706 10455 8746 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 10415 8620 10455 8660 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 10415 8534 10455 8574 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 10415 8448 10455 8488 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 10415 8362 10455 8402 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 10415 8276 10455 8316 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 10415 8190 10455 8230 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 10415 8104 10455 8144 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 10415 8018 10455 8058 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 10415 7932 10455 7972 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 10333 8792 10373 8832 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 10333 8706 10373 8746 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 10333 8620 10373 8660 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 10333 8534 10373 8574 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 10333 8448 10373 8488 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 10333 8362 10373 8402 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 10333 8276 10373 8316 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 10333 8190 10373 8230 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 10333 8104 10373 8144 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 10333 8018 10373 8058 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 10333 7932 10373 7972 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 10251 8792 10291 8832 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 10251 8706 10291 8746 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 10251 8620 10291 8660 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 10251 8534 10291 8574 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 10251 8448 10291 8488 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 10251 8362 10291 8402 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 10251 8276 10291 8316 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 10251 8190 10291 8230 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 10251 8104 10291 8144 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 10251 8018 10291 8058 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 10251 7932 10291 7972 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 10169 8792 10209 8832 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 10169 8706 10209 8746 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 10169 8620 10209 8660 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 10169 8534 10209 8574 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 10169 8448 10209 8488 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 10169 8362 10209 8402 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 10169 8276 10209 8316 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 10169 8190 10209 8230 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 10169 8104 10209 8144 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 10169 8018 10209 8058 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 10169 7932 10209 7972 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 4842 8792 4882 8832 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 4842 8706 4882 8746 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 4842 8620 4882 8660 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 4842 8534 4882 8574 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 4842 8448 4882 8488 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 4842 8362 4882 8402 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 4842 8276 4882 8316 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 4842 8190 4882 8230 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 4842 8104 4882 8144 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 4842 8018 4882 8058 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 4842 7932 4882 7972 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 4762 8792 4802 8832 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 4762 8706 4802 8746 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 4762 8620 4802 8660 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 4762 8534 4802 8574 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 4762 8448 4802 8488 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 4762 8362 4802 8402 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 4762 8276 4802 8316 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 4762 8190 4802 8230 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 4762 8104 4802 8144 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 4762 8018 4802 8058 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 4762 7932 4802 7972 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 4682 8792 4722 8832 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 4682 8706 4722 8746 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 4682 8620 4722 8660 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 4682 8534 4722 8574 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 4682 8448 4722 8488 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 4682 8362 4722 8402 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 4682 8276 4722 8316 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 4682 8190 4722 8230 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 4682 8104 4722 8144 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 4682 8018 4722 8058 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 4682 7932 4722 7972 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 4602 8792 4642 8832 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 4602 8706 4642 8746 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 4602 8620 4642 8660 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 4602 8534 4642 8574 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 4602 8448 4642 8488 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 4602 8362 4642 8402 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 4602 8276 4642 8316 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 4602 8190 4642 8230 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 4602 8104 4642 8144 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 4602 8018 4642 8058 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 4602 7932 4642 7972 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 4522 8792 4562 8832 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 4522 8706 4562 8746 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 4522 8620 4562 8660 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 4522 8534 4562 8574 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 4522 8448 4562 8488 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 4522 8362 4562 8402 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 4522 8276 4562 8316 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 4522 8190 4562 8230 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 4522 8104 4562 8144 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 4522 8018 4562 8058 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 4522 7932 4562 7972 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 4442 8792 4482 8832 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 4442 8706 4482 8746 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 4442 8620 4482 8660 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 4442 8534 4482 8574 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 4442 8448 4482 8488 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 4442 8362 4482 8402 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 4442 8276 4482 8316 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 4442 8190 4482 8230 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 4442 8104 4482 8144 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 4442 8018 4482 8058 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 4442 7932 4482 7972 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 4362 8792 4402 8832 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 4362 8706 4402 8746 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 4362 8620 4402 8660 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 4362 8534 4402 8574 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 4362 8448 4402 8488 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 4362 8362 4402 8402 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 4362 8276 4402 8316 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 4362 8190 4402 8230 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 4362 8104 4402 8144 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 4362 8018 4402 8058 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 4362 7932 4402 7972 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 4282 8792 4322 8832 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 4282 8706 4322 8746 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 4282 8620 4322 8660 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 4282 8534 4322 8574 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 4282 8448 4322 8488 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 4282 8362 4322 8402 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 4282 8276 4322 8316 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 4282 8190 4322 8230 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 4282 8104 4322 8144 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 4282 8018 4322 8058 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 4282 7932 4322 7972 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 4202 8792 4242 8832 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 4202 8706 4242 8746 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 4202 8620 4242 8660 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 4202 8534 4242 8574 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 4202 8448 4242 8488 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 4202 8362 4242 8402 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 4202 8276 4242 8316 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 4202 8190 4242 8230 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 4202 8104 4242 8144 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 4202 8018 4242 8058 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 4202 7932 4242 7972 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 4122 8792 4162 8832 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 4122 8706 4162 8746 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 4122 8620 4162 8660 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 4122 8534 4162 8574 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 4122 8448 4162 8488 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 4122 8362 4162 8402 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 4122 8276 4162 8316 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 4122 8190 4162 8230 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 4122 8104 4162 8144 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 4122 8018 4162 8058 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 4122 7932 4162 7972 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 4042 8792 4082 8832 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 4042 8706 4082 8746 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 4042 8620 4082 8660 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 4042 8534 4082 8574 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 4042 8448 4082 8488 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 4042 8362 4082 8402 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 4042 8276 4082 8316 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 4042 8190 4082 8230 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 4042 8104 4082 8144 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 4042 8018 4082 8058 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 4042 7932 4082 7972 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3962 8792 4002 8832 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3962 8706 4002 8746 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3962 8620 4002 8660 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3962 8534 4002 8574 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3962 8448 4002 8488 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3962 8362 4002 8402 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3962 8276 4002 8316 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3962 8190 4002 8230 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3962 8104 4002 8144 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3962 8018 4002 8058 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3962 7932 4002 7972 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3882 8792 3922 8832 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3882 8706 3922 8746 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3882 8620 3922 8660 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3882 8534 3922 8574 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3882 8448 3922 8488 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3882 8362 3922 8402 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3882 8276 3922 8316 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3882 8190 3922 8230 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3882 8104 3922 8144 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3882 8018 3922 8058 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3882 7932 3922 7972 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3802 8792 3842 8832 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3802 8706 3842 8746 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3802 8620 3842 8660 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3802 8534 3842 8574 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3802 8448 3842 8488 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3802 8362 3842 8402 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3802 8276 3842 8316 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3802 8190 3842 8230 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3802 8104 3842 8144 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3802 8018 3842 8058 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3802 7932 3842 7972 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3722 8792 3762 8832 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3722 8706 3762 8746 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3722 8620 3762 8660 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3722 8534 3762 8574 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3722 8448 3762 8488 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3722 8362 3762 8402 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3722 8276 3762 8316 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3722 8190 3762 8230 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3722 8104 3762 8144 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3722 8018 3762 8058 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3722 7932 3762 7972 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3642 8792 3682 8832 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3642 8706 3682 8746 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3642 8620 3682 8660 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3642 8534 3682 8574 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3642 8448 3682 8488 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3642 8362 3682 8402 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3642 8276 3682 8316 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3642 8190 3682 8230 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3642 8104 3682 8144 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3642 8018 3682 8058 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3642 7932 3682 7972 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3562 8792 3602 8832 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3562 8706 3602 8746 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3562 8620 3602 8660 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3562 8534 3602 8574 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3562 8448 3602 8488 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3562 8362 3602 8402 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3562 8276 3602 8316 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3562 8190 3602 8230 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3562 8104 3602 8144 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3562 8018 3602 8058 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3562 7932 3602 7972 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3482 8792 3522 8832 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3482 8706 3522 8746 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3482 8620 3522 8660 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3482 8534 3522 8574 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3482 8448 3522 8488 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3482 8362 3522 8402 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3482 8276 3522 8316 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3482 8190 3522 8230 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3482 8104 3522 8144 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3482 8018 3522 8058 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3482 7932 3522 7972 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3402 8792 3442 8832 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3402 8706 3442 8746 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3402 8620 3442 8660 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3402 8534 3442 8574 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3402 8448 3442 8488 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3402 8362 3442 8402 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3402 8276 3442 8316 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3402 8190 3442 8230 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3402 8104 3442 8144 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3402 8018 3442 8058 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3402 7932 3442 7972 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3322 8792 3362 8832 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3322 8706 3362 8746 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3322 8620 3362 8660 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3322 8534 3362 8574 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3322 8448 3362 8488 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3322 8362 3362 8402 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3322 8276 3362 8316 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3322 8190 3362 8230 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3322 8104 3362 8144 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3322 8018 3362 8058 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3322 7932 3362 7972 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3242 8792 3282 8832 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3242 8706 3282 8746 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3242 8620 3282 8660 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3242 8534 3282 8574 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3242 8448 3282 8488 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3242 8362 3282 8402 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3242 8276 3282 8316 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3242 8190 3282 8230 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3242 8104 3282 8144 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3242 8018 3282 8058 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3242 7932 3282 7972 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3162 8792 3202 8832 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3162 8706 3202 8746 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3162 8620 3202 8660 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3162 8534 3202 8574 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3162 8448 3202 8488 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3162 8362 3202 8402 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3162 8276 3202 8316 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3162 8190 3202 8230 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3162 8104 3202 8144 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3162 8018 3202 8058 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3162 7932 3202 7972 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3082 8792 3122 8832 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3082 8706 3122 8746 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3082 8620 3122 8660 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3082 8534 3122 8574 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3082 8448 3122 8488 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3082 8362 3122 8402 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3082 8276 3122 8316 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3082 8190 3122 8230 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3082 8104 3122 8144 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3082 8018 3122 8058 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3082 7932 3122 7972 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3002 8792 3042 8832 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3002 8706 3042 8746 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3002 8620 3042 8660 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3002 8534 3042 8574 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3002 8448 3042 8488 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3002 8362 3042 8402 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3002 8276 3042 8316 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3002 8190 3042 8230 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3002 8104 3042 8144 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3002 8018 3042 8058 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 3002 7932 3042 7972 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 2922 8792 2962 8832 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 2922 8706 2962 8746 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 2922 8620 2962 8660 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 2922 8534 2962 8574 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 2922 8448 2962 8488 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 2922 8362 2962 8402 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 2922 8276 2962 8316 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 2922 8190 2962 8230 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 2922 8104 2962 8144 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 2922 8018 2962 8058 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 2922 7932 2962 7972 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 2842 8792 2882 8832 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 2842 8706 2882 8746 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 2842 8620 2882 8660 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 2842 8534 2882 8574 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 2842 8448 2882 8488 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 2842 8362 2882 8402 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 2842 8276 2882 8316 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 2842 8190 2882 8230 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 2842 8104 2882 8144 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 2842 8018 2882 8058 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 2842 7932 2882 7972 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 2762 8792 2802 8832 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 2762 8706 2802 8746 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 2762 8620 2802 8660 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 2762 8534 2802 8574 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 2762 8448 2802 8488 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 2762 8362 2802 8402 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 2762 8276 2802 8316 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 2762 8190 2802 8230 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 2762 8104 2802 8144 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 2762 8018 2802 8058 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 2762 7932 2802 7972 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 2682 8792 2722 8832 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 2682 8706 2722 8746 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 2682 8620 2722 8660 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 2682 8534 2722 8574 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 2682 8448 2722 8488 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 2682 8362 2722 8402 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 2682 8276 2722 8316 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 2682 8190 2722 8230 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 2682 8104 2722 8144 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 2682 8018 2722 8058 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 2682 7932 2722 7972 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 2602 8792 2642 8832 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 2602 8706 2642 8746 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 2602 8620 2642 8660 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 2602 8534 2642 8574 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 2602 8448 2642 8488 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 2602 8362 2642 8402 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 2602 8276 2642 8316 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 2602 8190 2642 8230 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 2602 8104 2642 8144 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 2602 8018 2642 8058 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 2602 7932 2642 7972 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 2522 8792 2562 8832 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 2522 8706 2562 8746 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 2522 8620 2562 8660 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 2522 8534 2562 8574 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 2522 8448 2562 8488 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 2522 8362 2562 8402 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 2522 8276 2562 8316 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 2522 8190 2562 8230 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 2522 8104 2562 8144 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 2522 8018 2562 8058 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 2522 7932 2562 7972 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 2442 8792 2482 8832 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 2442 8706 2482 8746 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 2442 8620 2482 8660 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 2442 8534 2482 8574 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 2442 8448 2482 8488 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 2442 8362 2482 8402 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 2442 8276 2482 8316 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 2442 8190 2482 8230 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 2442 8104 2482 8144 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 2442 8018 2482 8058 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 2442 7932 2482 7972 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 2362 8792 2402 8832 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 2362 8706 2402 8746 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 2362 8620 2402 8660 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 2362 8534 2402 8574 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 2362 8448 2402 8488 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 2362 8362 2402 8402 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 2362 8276 2402 8316 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 2362 8190 2402 8230 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 2362 8104 2402 8144 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 2362 8018 2402 8058 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 2362 7932 2402 7972 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 2282 8792 2322 8832 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 2282 8706 2322 8746 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 2282 8620 2322 8660 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 2282 8534 2322 8574 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 2282 8448 2322 8488 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 2282 8362 2322 8402 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 2282 8276 2322 8316 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 2282 8190 2322 8230 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 2282 8104 2322 8144 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 2282 8018 2322 8058 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 2282 7932 2322 7972 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 2202 8792 2242 8832 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 2202 8706 2242 8746 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 2202 8620 2242 8660 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 2202 8534 2242 8574 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 2202 8448 2242 8488 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 2202 8362 2242 8402 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 2202 8276 2242 8316 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 2202 8190 2242 8230 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 2202 8104 2242 8144 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 2202 8018 2242 8058 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 2202 7932 2242 7972 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 2122 8792 2162 8832 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 2122 8706 2162 8746 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 2122 8620 2162 8660 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 2122 8534 2162 8574 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 2122 8448 2162 8488 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 2122 8362 2162 8402 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 2122 8276 2162 8316 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 2122 8190 2162 8230 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 2122 8104 2162 8144 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 2122 8018 2162 8058 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 2122 7932 2162 7972 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 2042 8792 2082 8832 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 2042 8706 2082 8746 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 2042 8620 2082 8660 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 2042 8534 2082 8574 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 2042 8448 2082 8488 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 2042 8362 2082 8402 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 2042 8276 2082 8316 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 2042 8190 2082 8230 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 2042 8104 2082 8144 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 2042 8018 2082 8058 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 2042 7932 2082 7972 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1962 8792 2002 8832 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1962 8706 2002 8746 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1962 8620 2002 8660 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1962 8534 2002 8574 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1962 8448 2002 8488 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1962 8362 2002 8402 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1962 8276 2002 8316 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1962 8190 2002 8230 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1962 8104 2002 8144 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1962 8018 2002 8058 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1962 7932 2002 7972 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1882 8792 1922 8832 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1882 8706 1922 8746 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1882 8620 1922 8660 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1882 8534 1922 8574 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1882 8448 1922 8488 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1882 8362 1922 8402 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1882 8276 1922 8316 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1882 8190 1922 8230 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1882 8104 1922 8144 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1882 8018 1922 8058 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1882 7932 1922 7972 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1802 8792 1842 8832 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1802 8706 1842 8746 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1802 8620 1842 8660 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1802 8534 1842 8574 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1802 8448 1842 8488 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1802 8362 1842 8402 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1802 8276 1842 8316 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1802 8190 1842 8230 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1802 8104 1842 8144 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1802 8018 1842 8058 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1802 7932 1842 7972 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1722 8792 1762 8832 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1722 8706 1762 8746 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1722 8620 1762 8660 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1722 8534 1762 8574 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1722 8448 1762 8488 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1722 8362 1762 8402 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1722 8276 1762 8316 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1722 8190 1762 8230 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1722 8104 1762 8144 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1722 8018 1762 8058 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1722 7932 1762 7972 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1642 8792 1682 8832 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1642 8706 1682 8746 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1642 8620 1682 8660 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1642 8534 1682 8574 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1642 8448 1682 8488 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1642 8362 1682 8402 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1642 8276 1682 8316 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1642 8190 1682 8230 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1642 8104 1682 8144 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1642 8018 1682 8058 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1642 7932 1682 7972 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1562 8792 1602 8832 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1562 8706 1602 8746 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1562 8620 1602 8660 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1562 8534 1602 8574 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1562 8448 1602 8488 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1562 8362 1602 8402 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1562 8276 1602 8316 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1562 8190 1602 8230 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1562 8104 1602 8144 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1562 8018 1602 8058 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1562 7932 1602 7972 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1482 8792 1522 8832 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1482 8706 1522 8746 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1482 8620 1522 8660 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1482 8534 1522 8574 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1482 8448 1522 8488 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1482 8362 1522 8402 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1482 8276 1522 8316 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1482 8190 1522 8230 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1482 8104 1522 8144 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1482 8018 1522 8058 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1482 7932 1522 7972 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1402 8792 1442 8832 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1402 8706 1442 8746 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1402 8620 1442 8660 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1402 8534 1442 8574 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1402 8448 1442 8488 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1402 8362 1442 8402 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1402 8276 1442 8316 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1402 8190 1442 8230 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1402 8104 1442 8144 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1402 8018 1442 8058 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1402 7932 1442 7972 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1322 8792 1362 8832 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1322 8706 1362 8746 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1322 8620 1362 8660 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1322 8534 1362 8574 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1322 8448 1362 8488 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1322 8362 1362 8402 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1322 8276 1362 8316 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1322 8190 1362 8230 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1322 8104 1362 8144 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1322 8018 1362 8058 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1322 7932 1362 7972 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1242 8792 1282 8832 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1242 8706 1282 8746 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1242 8620 1282 8660 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1242 8534 1282 8574 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1242 8448 1282 8488 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1242 8362 1282 8402 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1242 8276 1282 8316 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1242 8190 1282 8230 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1242 8104 1282 8144 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1242 8018 1282 8058 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1242 7932 1282 7972 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1162 8792 1202 8832 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1162 8706 1202 8746 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1162 8620 1202 8660 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1162 8534 1202 8574 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1162 8448 1202 8488 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1162 8362 1202 8402 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1162 8276 1202 8316 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1162 8190 1202 8230 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1162 8104 1202 8144 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1162 8018 1202 8058 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1162 7932 1202 7972 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1082 8792 1122 8832 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1082 8706 1122 8746 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1082 8620 1122 8660 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1082 8534 1122 8574 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1082 8448 1122 8488 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1082 8362 1122 8402 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1082 8276 1122 8316 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1082 8190 1122 8230 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1082 8104 1122 8144 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1082 8018 1122 8058 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1082 7932 1122 7972 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1002 8792 1042 8832 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1002 8706 1042 8746 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1002 8620 1042 8660 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1002 8534 1042 8574 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1002 8448 1042 8488 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1002 8362 1042 8402 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1002 8276 1042 8316 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1002 8190 1042 8230 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1002 8104 1042 8144 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1002 8018 1042 8058 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 1002 7932 1042 7972 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 922 8792 962 8832 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 922 8706 962 8746 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 922 8620 962 8660 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 922 8534 962 8574 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 922 8448 962 8488 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 922 8362 962 8402 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 922 8276 962 8316 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 922 8190 962 8230 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 922 8104 962 8144 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 922 8018 962 8058 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 922 7932 962 7972 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 842 8792 882 8832 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 842 8706 882 8746 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 842 8620 882 8660 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 842 8534 882 8574 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 842 8448 882 8488 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 842 8362 882 8402 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 842 8276 882 8316 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 842 8190 882 8230 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 842 8104 882 8144 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 842 8018 882 8058 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 842 7932 882 7972 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 762 8792 802 8832 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 762 8706 802 8746 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 762 8620 802 8660 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 762 8534 802 8574 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 762 8448 802 8488 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 762 8362 802 8402 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 762 8276 802 8316 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 762 8190 802 8230 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 762 8104 802 8144 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 762 8018 802 8058 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 762 7932 802 7972 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 682 8792 722 8832 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 682 8706 722 8746 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 682 8620 722 8660 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 682 8534 722 8574 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 682 8448 722 8488 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 682 8362 722 8402 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 682 8276 722 8316 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 682 8190 722 8230 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 682 8104 722 8144 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 682 8018 722 8058 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 682 7932 722 7972 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 602 8792 642 8832 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 602 8706 642 8746 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 602 8620 642 8660 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 602 8534 642 8574 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 602 8448 642 8488 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 602 8362 642 8402 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 602 8276 642 8316 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 602 8190 642 8230 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 602 8104 642 8144 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 602 8018 642 8058 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 602 7932 642 7972 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 522 8792 562 8832 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 522 8706 562 8746 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 522 8620 562 8660 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 522 8534 562 8574 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 522 8448 562 8488 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 522 8362 562 8402 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 522 8276 562 8316 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 522 8190 562 8230 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 522 8104 562 8144 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 522 8018 562 8058 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 522 7932 562 7972 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 442 8792 482 8832 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 442 8706 482 8746 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 442 8620 482 8660 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 442 8534 482 8574 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 442 8448 482 8488 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 442 8362 482 8402 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 442 8276 482 8316 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 442 8190 482 8230 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 442 8104 482 8144 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 442 8018 482 8058 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 442 7932 482 7972 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 361 8792 401 8832 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 361 8706 401 8746 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 361 8620 401 8660 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 361 8534 401 8574 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 361 8448 401 8488 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 361 8362 401 8402 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 361 8276 401 8316 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 361 8190 401 8230 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 361 8104 401 8144 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 361 8018 401 8058 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 361 7932 401 7972 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 280 8792 320 8832 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 280 8706 320 8746 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 280 8620 320 8660 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 280 8534 320 8574 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 280 8448 320 8488 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 280 8362 320 8402 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 280 8276 320 8316 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 280 8190 320 8230 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 280 8104 320 8144 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 280 8018 320 8058 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 280 7932 320 7972 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 199 8792 239 8832 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 199 8706 239 8746 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 199 8620 239 8660 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 199 8534 239 8574 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 199 8448 239 8488 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 199 8362 239 8402 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 199 8276 239 8316 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 199 8190 239 8230 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 199 8104 239 8144 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 199 8018 239 8058 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 199 7932 239 7972 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 118 8792 158 8832 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 118 8706 158 8746 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 118 8620 158 8660 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 118 8534 158 8574 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 118 8448 158 8488 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 118 8362 158 8402 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 118 8276 158 8316 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 118 8190 158 8230 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 118 8104 158 8144 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 118 8018 158 8058 1 VSSD
port 4 nsew ground bidirectional
rlabel via3 s 118 7932 158 7972 1 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 14746 34757 15000 39600 1 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 14746 4767 15000 5697 1 VSSIO
port 5 nsew ground bidirectional
rlabel metal5 s 0 34757 254 39600 1 VSSIO
port 5 nsew ground bidirectional
rlabel metal5 s 0 4787 254 5677 1 VSSIO
port 5 nsew ground bidirectional
rlabel metal5 s 14746 34757 15000 39600 1 VSSIO
port 5 nsew ground bidirectional
rlabel metal5 s 14746 4787 15000 5677 1 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 14746 11247 15000 12137 1 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal5 s 0 11267 254 12117 1 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal5 s 14746 11267 15000 12117 1 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 14746 5977 15000 6667 1 VSWITCH
port 6 nsew power bidirectional
rlabel metal5 s 0 5997 254 6647 1 VSWITCH
port 6 nsew power bidirectional
rlabel metal5 s 14746 5997 15000 6647 1 VSWITCH
port 6 nsew power bidirectional
<< properties >>
string FIXED_BBOX 0 0 15000 39600
string GDS_END 2266656
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 2174144
string LEFclass PAD
string LEFsymmetry X Y R90
<< end >>
