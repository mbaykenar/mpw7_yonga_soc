magic
tech sky130B
magscale 1 2
timestamp 1649977179
use sky130_fd_pr__hvdfm1sd2__example_55959141808251  sky130_fd_pr__hvdfm1sd2__example_55959141808251_0
timestamp 1649977179
transform 1 0 30 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfm1sd2__example_55959141808251  sky130_fd_pr__hvdfm1sd2__example_55959141808251_1
timestamp 1649977179
transform 1 0 116 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfm1sd2__example_55959141808251  sky130_fd_pr__hvdfm1sd2__example_55959141808251_2
timestamp 1649977179
transform 1 0 202 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfm1sd2__example_55959141808251  sky130_fd_pr__hvdfm1sd2__example_55959141808251_3
timestamp 1649977179
transform 1 0 288 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfm1sd__example_55959141808250  sky130_fd_pr__hvdfm1sd__example_55959141808250_0
timestamp 1649977179
transform -1 0 0 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfm1sd__example_55959141808250  sky130_fd_pr__hvdfm1sd__example_55959141808250_1
timestamp 1649977179
transform 1 0 374 0 1 0
box 0 0 1 1
<< labels >>
flabel comment s 402 697 402 697 0 FreeSans 300 0 0 0 D
flabel comment s 316 697 316 697 0 FreeSans 300 0 0 0 S
flabel comment s 230 697 230 697 0 FreeSans 300 0 0 0 D
flabel comment s 144 697 144 697 0 FreeSans 300 0 0 0 S
flabel comment s 58 697 58 697 0 FreeSans 300 0 0 0 D
flabel comment s -28 697 -28 697 0 FreeSans 300 0 0 0 S
<< properties >>
string GDS_END 37227056
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 37224058
<< end >>
