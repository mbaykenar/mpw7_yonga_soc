magic
tech sky130B
magscale 1 2
timestamp 1649977179
<< nwell >>
rect -66 377 258 897
<< pwell >>
rect 4 43 188 317
rect -26 -43 218 43
<< mvpsubdiff >>
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 192 17
<< mvnsubdiff >>
rect 0 797 31 831
rect 65 797 127 831
rect 161 797 192 831
<< mvpsubdiffcont >>
rect 31 -17 65 17
rect 127 -17 161 17
<< mvnsubdiffcont >>
rect 31 797 65 831
rect 127 797 161 831
<< mvndiode >>
rect 30 279 162 291
rect 30 245 42 279
rect 76 245 116 279
rect 150 245 162 279
rect 30 153 162 245
rect 30 119 42 153
rect 76 119 116 153
rect 150 119 162 153
rect 30 107 162 119
<< mvndiodec >>
rect 42 245 76 279
rect 116 245 150 279
rect 42 119 76 153
rect 116 119 150 153
<< locali >>
rect 0 797 31 831
rect 65 797 127 831
rect 161 797 192 831
rect 21 279 171 656
rect 21 245 42 279
rect 76 245 116 279
rect 150 245 171 279
rect 21 153 171 245
rect 21 119 42 153
rect 76 119 116 153
rect 150 119 171 153
rect 21 103 171 119
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 192 17
<< viali >>
rect 31 797 65 831
rect 127 797 161 831
rect 31 -17 65 17
rect 127 -17 161 17
<< metal1 >>
rect 0 831 192 837
rect 0 797 31 831
rect 65 797 127 831
rect 161 797 192 831
rect 0 791 192 797
rect 0 689 192 763
rect 0 51 192 125
rect 0 17 192 23
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 192 17
rect 0 -23 192 -17
<< labels >>
flabel locali s 31 612 65 646 0 FreeSans 200 0 0 0 DIODE
port 1 nsew default input
flabel locali s 127 612 161 646 0 FreeSans 200 0 0 0 DIODE
port 1 nsew default input
flabel locali s 31 538 65 572 0 FreeSans 200 0 0 0 DIODE
port 1 nsew default input
flabel locali s 127 538 161 572 0 FreeSans 200 0 0 0 DIODE
port 1 nsew default input
flabel locali s 31 464 65 498 0 FreeSans 200 0 0 0 DIODE
port 1 nsew default input
flabel locali s 127 464 161 498 0 FreeSans 200 0 0 0 DIODE
port 1 nsew default input
flabel locali s 31 390 65 424 0 FreeSans 200 0 0 0 DIODE
port 1 nsew default input
flabel locali s 127 390 161 424 0 FreeSans 200 0 0 0 DIODE
port 1 nsew default input
flabel locali s 31 316 65 350 0 FreeSans 200 0 0 0 DIODE
port 1 nsew default input
flabel locali s 127 316 161 350 0 FreeSans 200 0 0 0 DIODE
port 1 nsew default input
flabel locali s 127 242 161 276 0 FreeSans 200 0 0 0 DIODE
port 1 nsew default input
flabel locali s 127 168 161 202 0 FreeSans 200 0 0 0 DIODE
port 1 nsew default input
flabel locali s 31 168 65 202 0 FreeSans 200 0 0 0 DIODE
port 1 nsew default input
flabel locali s 31 242 65 276 0 FreeSans 200 0 0 0 DIODE
port 1 nsew default input
rlabel comment s 0 0 0 0 4 diode_2
flabel metal1 s 0 51 192 125 0 FreeSans 340 0 0 0 VGND
port 2 nsew ground bidirectional
flabel metal1 s 0 0 192 23 0 FreeSans 340 0 0 0 VNB
port 3 nsew ground bidirectional
flabel metal1 s 96 11 96 11 0 FreeSans 340 0 0 0 VNB
port 3 nsew
flabel metal1 s 0 689 192 763 0 FreeSans 340 0 0 0 VPWR
port 5 nsew power bidirectional
flabel metal1 s 0 791 192 814 0 FreeSans 340 0 0 0 VPB
port 4 nsew power bidirectional
flabel metal1 s 96 802 96 802 0 FreeSans 340 0 0 0 VPB
port 4 nsew
<< properties >>
string FIXED_BBOX 0 0 192 814
string GDS_END 1159870
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hvl/gds/sky130_fd_sc_hvl.gds
string GDS_START 1154836
string LEFclass CORE ANTENNACELL
string LEFsite unithv
string LEFsymmetry X Y
<< end >>
