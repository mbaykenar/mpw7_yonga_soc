magic
tech sky130B
magscale 1 2
timestamp 1649977179
use sky130_fd_pr__hvdfm1sd__example_5595914180846  sky130_fd_pr__hvdfm1sd__example_5595914180846_0
timestamp 1649977179
transform -1 0 0 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfm1sd__example_5595914180846  sky130_fd_pr__hvdfm1sd__example_5595914180846_1
timestamp 1649977179
transform 1 0 100 0 1 0
box 0 0 1 1
<< labels >>
flabel comment s 128 985 128 985 0 FreeSans 300 0 0 0 D
flabel comment s -28 985 -28 985 0 FreeSans 300 0 0 0 S
<< properties >>
string GDS_END 47706744
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 47705690
<< end >>
