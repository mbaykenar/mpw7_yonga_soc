magic
tech sky130B
magscale 1 2
timestamp 1649977179
<< metal3 >>
rect 10151 7918 14940 8846
<< obsm3 >>
rect 100 7918 4900 8846
<< metal4 >>
rect 0 34757 254 39600
rect 14746 34757 15000 39600
rect 0 13607 254 18600
rect 14746 13607 15000 18600
rect 0 12417 254 13307
rect 14746 12417 15000 13307
rect 0 11247 254 12137
rect 14746 11247 15000 12137
rect 0 10881 15000 10947
rect 0 10225 15000 10821
rect 0 9929 254 10165
rect 14746 9929 15000 10165
rect 0 9273 15000 9869
rect 0 9147 15000 9213
rect 0 7917 254 8847
rect 268 8780 332 8844
rect 349 8780 413 8844
rect 430 8780 494 8844
rect 510 8780 574 8844
rect 590 8780 654 8844
rect 670 8780 734 8844
rect 750 8780 814 8844
rect 830 8780 894 8844
rect 910 8780 974 8844
rect 990 8780 1054 8844
rect 1070 8780 1134 8844
rect 1150 8780 1214 8844
rect 1230 8780 1294 8844
rect 1310 8780 1374 8844
rect 1390 8780 1454 8844
rect 1470 8780 1534 8844
rect 1550 8780 1614 8844
rect 1630 8780 1694 8844
rect 1710 8780 1774 8844
rect 1790 8780 1854 8844
rect 1870 8780 1934 8844
rect 1950 8780 2014 8844
rect 2030 8780 2094 8844
rect 2110 8780 2174 8844
rect 2190 8780 2254 8844
rect 2270 8780 2334 8844
rect 2350 8780 2414 8844
rect 2430 8780 2494 8844
rect 2510 8780 2574 8844
rect 2590 8780 2654 8844
rect 2670 8780 2734 8844
rect 2750 8780 2814 8844
rect 2830 8780 2894 8844
rect 2910 8780 2974 8844
rect 2990 8780 3054 8844
rect 3070 8780 3134 8844
rect 3150 8780 3214 8844
rect 3230 8780 3294 8844
rect 3310 8780 3374 8844
rect 3390 8780 3454 8844
rect 3470 8780 3534 8844
rect 3550 8780 3614 8844
rect 3630 8780 3694 8844
rect 3710 8780 3774 8844
rect 3790 8780 3854 8844
rect 3870 8780 3934 8844
rect 3950 8780 4014 8844
rect 4030 8780 4094 8844
rect 4110 8780 4174 8844
rect 4190 8780 4254 8844
rect 4270 8780 4334 8844
rect 4350 8780 4414 8844
rect 4430 8780 4494 8844
rect 4510 8780 4574 8844
rect 4590 8780 4654 8844
rect 4670 8780 4734 8844
rect 4750 8780 4814 8844
rect 4830 8780 4894 8844
rect 268 8694 332 8758
rect 349 8694 413 8758
rect 430 8694 494 8758
rect 510 8694 574 8758
rect 590 8694 654 8758
rect 670 8694 734 8758
rect 750 8694 814 8758
rect 830 8694 894 8758
rect 910 8694 974 8758
rect 990 8694 1054 8758
rect 1070 8694 1134 8758
rect 1150 8694 1214 8758
rect 1230 8694 1294 8758
rect 1310 8694 1374 8758
rect 1390 8694 1454 8758
rect 1470 8694 1534 8758
rect 1550 8694 1614 8758
rect 1630 8694 1694 8758
rect 1710 8694 1774 8758
rect 1790 8694 1854 8758
rect 1870 8694 1934 8758
rect 1950 8694 2014 8758
rect 2030 8694 2094 8758
rect 2110 8694 2174 8758
rect 2190 8694 2254 8758
rect 2270 8694 2334 8758
rect 2350 8694 2414 8758
rect 2430 8694 2494 8758
rect 2510 8694 2574 8758
rect 2590 8694 2654 8758
rect 2670 8694 2734 8758
rect 2750 8694 2814 8758
rect 2830 8694 2894 8758
rect 2910 8694 2974 8758
rect 2990 8694 3054 8758
rect 3070 8694 3134 8758
rect 3150 8694 3214 8758
rect 3230 8694 3294 8758
rect 3310 8694 3374 8758
rect 3390 8694 3454 8758
rect 3470 8694 3534 8758
rect 3550 8694 3614 8758
rect 3630 8694 3694 8758
rect 3710 8694 3774 8758
rect 3790 8694 3854 8758
rect 3870 8694 3934 8758
rect 3950 8694 4014 8758
rect 4030 8694 4094 8758
rect 4110 8694 4174 8758
rect 4190 8694 4254 8758
rect 4270 8694 4334 8758
rect 4350 8694 4414 8758
rect 4430 8694 4494 8758
rect 4510 8694 4574 8758
rect 4590 8694 4654 8758
rect 4670 8694 4734 8758
rect 4750 8694 4814 8758
rect 4830 8694 4894 8758
rect 268 8608 332 8672
rect 349 8608 413 8672
rect 430 8608 494 8672
rect 510 8608 574 8672
rect 590 8608 654 8672
rect 670 8608 734 8672
rect 750 8608 814 8672
rect 830 8608 894 8672
rect 910 8608 974 8672
rect 990 8608 1054 8672
rect 1070 8608 1134 8672
rect 1150 8608 1214 8672
rect 1230 8608 1294 8672
rect 1310 8608 1374 8672
rect 1390 8608 1454 8672
rect 1470 8608 1534 8672
rect 1550 8608 1614 8672
rect 1630 8608 1694 8672
rect 1710 8608 1774 8672
rect 1790 8608 1854 8672
rect 1870 8608 1934 8672
rect 1950 8608 2014 8672
rect 2030 8608 2094 8672
rect 2110 8608 2174 8672
rect 2190 8608 2254 8672
rect 2270 8608 2334 8672
rect 2350 8608 2414 8672
rect 2430 8608 2494 8672
rect 2510 8608 2574 8672
rect 2590 8608 2654 8672
rect 2670 8608 2734 8672
rect 2750 8608 2814 8672
rect 2830 8608 2894 8672
rect 2910 8608 2974 8672
rect 2990 8608 3054 8672
rect 3070 8608 3134 8672
rect 3150 8608 3214 8672
rect 3230 8608 3294 8672
rect 3310 8608 3374 8672
rect 3390 8608 3454 8672
rect 3470 8608 3534 8672
rect 3550 8608 3614 8672
rect 3630 8608 3694 8672
rect 3710 8608 3774 8672
rect 3790 8608 3854 8672
rect 3870 8608 3934 8672
rect 3950 8608 4014 8672
rect 4030 8608 4094 8672
rect 4110 8608 4174 8672
rect 4190 8608 4254 8672
rect 4270 8608 4334 8672
rect 4350 8608 4414 8672
rect 4430 8608 4494 8672
rect 4510 8608 4574 8672
rect 4590 8608 4654 8672
rect 4670 8608 4734 8672
rect 4750 8608 4814 8672
rect 4830 8608 4894 8672
rect 268 8522 332 8586
rect 349 8522 413 8586
rect 430 8522 494 8586
rect 510 8522 574 8586
rect 590 8522 654 8586
rect 670 8522 734 8586
rect 750 8522 814 8586
rect 830 8522 894 8586
rect 910 8522 974 8586
rect 990 8522 1054 8586
rect 1070 8522 1134 8586
rect 1150 8522 1214 8586
rect 1230 8522 1294 8586
rect 1310 8522 1374 8586
rect 1390 8522 1454 8586
rect 1470 8522 1534 8586
rect 1550 8522 1614 8586
rect 1630 8522 1694 8586
rect 1710 8522 1774 8586
rect 1790 8522 1854 8586
rect 1870 8522 1934 8586
rect 1950 8522 2014 8586
rect 2030 8522 2094 8586
rect 2110 8522 2174 8586
rect 2190 8522 2254 8586
rect 2270 8522 2334 8586
rect 2350 8522 2414 8586
rect 2430 8522 2494 8586
rect 2510 8522 2574 8586
rect 2590 8522 2654 8586
rect 2670 8522 2734 8586
rect 2750 8522 2814 8586
rect 2830 8522 2894 8586
rect 2910 8522 2974 8586
rect 2990 8522 3054 8586
rect 3070 8522 3134 8586
rect 3150 8522 3214 8586
rect 3230 8522 3294 8586
rect 3310 8522 3374 8586
rect 3390 8522 3454 8586
rect 3470 8522 3534 8586
rect 3550 8522 3614 8586
rect 3630 8522 3694 8586
rect 3710 8522 3774 8586
rect 3790 8522 3854 8586
rect 3870 8522 3934 8586
rect 3950 8522 4014 8586
rect 4030 8522 4094 8586
rect 4110 8522 4174 8586
rect 4190 8522 4254 8586
rect 4270 8522 4334 8586
rect 4350 8522 4414 8586
rect 4430 8522 4494 8586
rect 4510 8522 4574 8586
rect 4590 8522 4654 8586
rect 4670 8522 4734 8586
rect 4750 8522 4814 8586
rect 4830 8522 4894 8586
rect 268 8436 332 8500
rect 349 8436 413 8500
rect 430 8436 494 8500
rect 510 8436 574 8500
rect 590 8436 654 8500
rect 670 8436 734 8500
rect 750 8436 814 8500
rect 830 8436 894 8500
rect 910 8436 974 8500
rect 990 8436 1054 8500
rect 1070 8436 1134 8500
rect 1150 8436 1214 8500
rect 1230 8436 1294 8500
rect 1310 8436 1374 8500
rect 1390 8436 1454 8500
rect 1470 8436 1534 8500
rect 1550 8436 1614 8500
rect 1630 8436 1694 8500
rect 1710 8436 1774 8500
rect 1790 8436 1854 8500
rect 1870 8436 1934 8500
rect 1950 8436 2014 8500
rect 2030 8436 2094 8500
rect 2110 8436 2174 8500
rect 2190 8436 2254 8500
rect 2270 8436 2334 8500
rect 2350 8436 2414 8500
rect 2430 8436 2494 8500
rect 2510 8436 2574 8500
rect 2590 8436 2654 8500
rect 2670 8436 2734 8500
rect 2750 8436 2814 8500
rect 2830 8436 2894 8500
rect 2910 8436 2974 8500
rect 2990 8436 3054 8500
rect 3070 8436 3134 8500
rect 3150 8436 3214 8500
rect 3230 8436 3294 8500
rect 3310 8436 3374 8500
rect 3390 8436 3454 8500
rect 3470 8436 3534 8500
rect 3550 8436 3614 8500
rect 3630 8436 3694 8500
rect 3710 8436 3774 8500
rect 3790 8436 3854 8500
rect 3870 8436 3934 8500
rect 3950 8436 4014 8500
rect 4030 8436 4094 8500
rect 4110 8436 4174 8500
rect 4190 8436 4254 8500
rect 4270 8436 4334 8500
rect 4350 8436 4414 8500
rect 4430 8436 4494 8500
rect 4510 8436 4574 8500
rect 4590 8436 4654 8500
rect 4670 8436 4734 8500
rect 4750 8436 4814 8500
rect 4830 8436 4894 8500
rect 268 8350 332 8414
rect 349 8350 413 8414
rect 430 8350 494 8414
rect 510 8350 574 8414
rect 590 8350 654 8414
rect 670 8350 734 8414
rect 750 8350 814 8414
rect 830 8350 894 8414
rect 910 8350 974 8414
rect 990 8350 1054 8414
rect 1070 8350 1134 8414
rect 1150 8350 1214 8414
rect 1230 8350 1294 8414
rect 1310 8350 1374 8414
rect 1390 8350 1454 8414
rect 1470 8350 1534 8414
rect 1550 8350 1614 8414
rect 1630 8350 1694 8414
rect 1710 8350 1774 8414
rect 1790 8350 1854 8414
rect 1870 8350 1934 8414
rect 1950 8350 2014 8414
rect 2030 8350 2094 8414
rect 2110 8350 2174 8414
rect 2190 8350 2254 8414
rect 2270 8350 2334 8414
rect 2350 8350 2414 8414
rect 2430 8350 2494 8414
rect 2510 8350 2574 8414
rect 2590 8350 2654 8414
rect 2670 8350 2734 8414
rect 2750 8350 2814 8414
rect 2830 8350 2894 8414
rect 2910 8350 2974 8414
rect 2990 8350 3054 8414
rect 3070 8350 3134 8414
rect 3150 8350 3214 8414
rect 3230 8350 3294 8414
rect 3310 8350 3374 8414
rect 3390 8350 3454 8414
rect 3470 8350 3534 8414
rect 3550 8350 3614 8414
rect 3630 8350 3694 8414
rect 3710 8350 3774 8414
rect 3790 8350 3854 8414
rect 3870 8350 3934 8414
rect 3950 8350 4014 8414
rect 4030 8350 4094 8414
rect 4110 8350 4174 8414
rect 4190 8350 4254 8414
rect 4270 8350 4334 8414
rect 4350 8350 4414 8414
rect 4430 8350 4494 8414
rect 4510 8350 4574 8414
rect 4590 8350 4654 8414
rect 4670 8350 4734 8414
rect 4750 8350 4814 8414
rect 4830 8350 4894 8414
rect 268 8264 332 8328
rect 349 8264 413 8328
rect 430 8264 494 8328
rect 510 8264 574 8328
rect 590 8264 654 8328
rect 670 8264 734 8328
rect 750 8264 814 8328
rect 830 8264 894 8328
rect 910 8264 974 8328
rect 990 8264 1054 8328
rect 1070 8264 1134 8328
rect 1150 8264 1214 8328
rect 1230 8264 1294 8328
rect 1310 8264 1374 8328
rect 1390 8264 1454 8328
rect 1470 8264 1534 8328
rect 1550 8264 1614 8328
rect 1630 8264 1694 8328
rect 1710 8264 1774 8328
rect 1790 8264 1854 8328
rect 1870 8264 1934 8328
rect 1950 8264 2014 8328
rect 2030 8264 2094 8328
rect 2110 8264 2174 8328
rect 2190 8264 2254 8328
rect 2270 8264 2334 8328
rect 2350 8264 2414 8328
rect 2430 8264 2494 8328
rect 2510 8264 2574 8328
rect 2590 8264 2654 8328
rect 2670 8264 2734 8328
rect 2750 8264 2814 8328
rect 2830 8264 2894 8328
rect 2910 8264 2974 8328
rect 2990 8264 3054 8328
rect 3070 8264 3134 8328
rect 3150 8264 3214 8328
rect 3230 8264 3294 8328
rect 3310 8264 3374 8328
rect 3390 8264 3454 8328
rect 3470 8264 3534 8328
rect 3550 8264 3614 8328
rect 3630 8264 3694 8328
rect 3710 8264 3774 8328
rect 3790 8264 3854 8328
rect 3870 8264 3934 8328
rect 3950 8264 4014 8328
rect 4030 8264 4094 8328
rect 4110 8264 4174 8328
rect 4190 8264 4254 8328
rect 4270 8264 4334 8328
rect 4350 8264 4414 8328
rect 4430 8264 4494 8328
rect 4510 8264 4574 8328
rect 4590 8264 4654 8328
rect 4670 8264 4734 8328
rect 4750 8264 4814 8328
rect 4830 8264 4894 8328
rect 268 8178 332 8242
rect 349 8178 413 8242
rect 430 8178 494 8242
rect 510 8178 574 8242
rect 590 8178 654 8242
rect 670 8178 734 8242
rect 750 8178 814 8242
rect 830 8178 894 8242
rect 910 8178 974 8242
rect 990 8178 1054 8242
rect 1070 8178 1134 8242
rect 1150 8178 1214 8242
rect 1230 8178 1294 8242
rect 1310 8178 1374 8242
rect 1390 8178 1454 8242
rect 1470 8178 1534 8242
rect 1550 8178 1614 8242
rect 1630 8178 1694 8242
rect 1710 8178 1774 8242
rect 1790 8178 1854 8242
rect 1870 8178 1934 8242
rect 1950 8178 2014 8242
rect 2030 8178 2094 8242
rect 2110 8178 2174 8242
rect 2190 8178 2254 8242
rect 2270 8178 2334 8242
rect 2350 8178 2414 8242
rect 2430 8178 2494 8242
rect 2510 8178 2574 8242
rect 2590 8178 2654 8242
rect 2670 8178 2734 8242
rect 2750 8178 2814 8242
rect 2830 8178 2894 8242
rect 2910 8178 2974 8242
rect 2990 8178 3054 8242
rect 3070 8178 3134 8242
rect 3150 8178 3214 8242
rect 3230 8178 3294 8242
rect 3310 8178 3374 8242
rect 3390 8178 3454 8242
rect 3470 8178 3534 8242
rect 3550 8178 3614 8242
rect 3630 8178 3694 8242
rect 3710 8178 3774 8242
rect 3790 8178 3854 8242
rect 3870 8178 3934 8242
rect 3950 8178 4014 8242
rect 4030 8178 4094 8242
rect 4110 8178 4174 8242
rect 4190 8178 4254 8242
rect 4270 8178 4334 8242
rect 4350 8178 4414 8242
rect 4430 8178 4494 8242
rect 4510 8178 4574 8242
rect 4590 8178 4654 8242
rect 4670 8178 4734 8242
rect 4750 8178 4814 8242
rect 4830 8178 4894 8242
rect 268 8092 332 8156
rect 349 8092 413 8156
rect 430 8092 494 8156
rect 510 8092 574 8156
rect 590 8092 654 8156
rect 670 8092 734 8156
rect 750 8092 814 8156
rect 830 8092 894 8156
rect 910 8092 974 8156
rect 990 8092 1054 8156
rect 1070 8092 1134 8156
rect 1150 8092 1214 8156
rect 1230 8092 1294 8156
rect 1310 8092 1374 8156
rect 1390 8092 1454 8156
rect 1470 8092 1534 8156
rect 1550 8092 1614 8156
rect 1630 8092 1694 8156
rect 1710 8092 1774 8156
rect 1790 8092 1854 8156
rect 1870 8092 1934 8156
rect 1950 8092 2014 8156
rect 2030 8092 2094 8156
rect 2110 8092 2174 8156
rect 2190 8092 2254 8156
rect 2270 8092 2334 8156
rect 2350 8092 2414 8156
rect 2430 8092 2494 8156
rect 2510 8092 2574 8156
rect 2590 8092 2654 8156
rect 2670 8092 2734 8156
rect 2750 8092 2814 8156
rect 2830 8092 2894 8156
rect 2910 8092 2974 8156
rect 2990 8092 3054 8156
rect 3070 8092 3134 8156
rect 3150 8092 3214 8156
rect 3230 8092 3294 8156
rect 3310 8092 3374 8156
rect 3390 8092 3454 8156
rect 3470 8092 3534 8156
rect 3550 8092 3614 8156
rect 3630 8092 3694 8156
rect 3710 8092 3774 8156
rect 3790 8092 3854 8156
rect 3870 8092 3934 8156
rect 3950 8092 4014 8156
rect 4030 8092 4094 8156
rect 4110 8092 4174 8156
rect 4190 8092 4254 8156
rect 4270 8092 4334 8156
rect 4350 8092 4414 8156
rect 4430 8092 4494 8156
rect 4510 8092 4574 8156
rect 4590 8092 4654 8156
rect 4670 8092 4734 8156
rect 4750 8092 4814 8156
rect 4830 8092 4894 8156
rect 268 8006 332 8070
rect 349 8006 413 8070
rect 430 8006 494 8070
rect 510 8006 574 8070
rect 590 8006 654 8070
rect 670 8006 734 8070
rect 750 8006 814 8070
rect 830 8006 894 8070
rect 910 8006 974 8070
rect 990 8006 1054 8070
rect 1070 8006 1134 8070
rect 1150 8006 1214 8070
rect 1230 8006 1294 8070
rect 1310 8006 1374 8070
rect 1390 8006 1454 8070
rect 1470 8006 1534 8070
rect 1550 8006 1614 8070
rect 1630 8006 1694 8070
rect 1710 8006 1774 8070
rect 1790 8006 1854 8070
rect 1870 8006 1934 8070
rect 1950 8006 2014 8070
rect 2030 8006 2094 8070
rect 2110 8006 2174 8070
rect 2190 8006 2254 8070
rect 2270 8006 2334 8070
rect 2350 8006 2414 8070
rect 2430 8006 2494 8070
rect 2510 8006 2574 8070
rect 2590 8006 2654 8070
rect 2670 8006 2734 8070
rect 2750 8006 2814 8070
rect 2830 8006 2894 8070
rect 2910 8006 2974 8070
rect 2990 8006 3054 8070
rect 3070 8006 3134 8070
rect 3150 8006 3214 8070
rect 3230 8006 3294 8070
rect 3310 8006 3374 8070
rect 3390 8006 3454 8070
rect 3470 8006 3534 8070
rect 3550 8006 3614 8070
rect 3630 8006 3694 8070
rect 3710 8006 3774 8070
rect 3790 8006 3854 8070
rect 3870 8006 3934 8070
rect 3950 8006 4014 8070
rect 4030 8006 4094 8070
rect 4110 8006 4174 8070
rect 4190 8006 4254 8070
rect 4270 8006 4334 8070
rect 4350 8006 4414 8070
rect 4430 8006 4494 8070
rect 4510 8006 4574 8070
rect 4590 8006 4654 8070
rect 4670 8006 4734 8070
rect 4750 8006 4814 8070
rect 4830 8006 4894 8070
rect 268 7920 332 7984
rect 349 7920 413 7984
rect 430 7920 494 7984
rect 510 7920 574 7984
rect 590 7920 654 7984
rect 670 7920 734 7984
rect 750 7920 814 7984
rect 830 7920 894 7984
rect 910 7920 974 7984
rect 990 7920 1054 7984
rect 1070 7920 1134 7984
rect 1150 7920 1214 7984
rect 1230 7920 1294 7984
rect 1310 7920 1374 7984
rect 1390 7920 1454 7984
rect 1470 7920 1534 7984
rect 1550 7920 1614 7984
rect 1630 7920 1694 7984
rect 1710 7920 1774 7984
rect 1790 7920 1854 7984
rect 1870 7920 1934 7984
rect 1950 7920 2014 7984
rect 2030 7920 2094 7984
rect 2110 7920 2174 7984
rect 2190 7920 2254 7984
rect 2270 7920 2334 7984
rect 2350 7920 2414 7984
rect 2430 7920 2494 7984
rect 2510 7920 2574 7984
rect 2590 7920 2654 7984
rect 2670 7920 2734 7984
rect 2750 7920 2814 7984
rect 2830 7920 2894 7984
rect 2910 7920 2974 7984
rect 2990 7920 3054 7984
rect 3070 7920 3134 7984
rect 3150 7920 3214 7984
rect 3230 7920 3294 7984
rect 3310 7920 3374 7984
rect 3390 7920 3454 7984
rect 3470 7920 3534 7984
rect 3550 7920 3614 7984
rect 3630 7920 3694 7984
rect 3710 7920 3774 7984
rect 3790 7920 3854 7984
rect 3870 7920 3934 7984
rect 3950 7920 4014 7984
rect 4030 7920 4094 7984
rect 4110 7920 4174 7984
rect 4190 7920 4254 7984
rect 4270 7920 4334 7984
rect 4350 7920 4414 7984
rect 4430 7920 4494 7984
rect 4510 7920 4574 7984
rect 4590 7920 4654 7984
rect 4670 7920 4734 7984
rect 4750 7920 4814 7984
rect 4830 7920 4894 7984
rect 14746 7917 15000 8847
rect 0 6947 254 7637
rect 14746 6947 15000 7637
rect 0 5977 254 6667
rect 14746 5977 15000 6667
rect 0 4767 254 5697
rect 14746 4767 15000 5697
rect 0 3557 254 4487
rect 14746 3557 15000 4487
rect 0 2587 193 3277
rect 14807 2587 15000 3277
rect 0 1377 254 2307
rect 14746 1377 15000 2307
rect 0 7 254 1097
rect 14746 7 15000 1097
<< obsm4 >>
rect 334 34677 14666 39600
rect 193 18680 14807 34677
rect 334 13527 14666 18680
rect 193 13387 14807 13527
rect 334 12337 14666 13387
rect 193 12217 14807 12337
rect 334 11167 14666 12217
rect 193 11027 14807 11167
rect 334 9949 14666 10145
rect 193 8927 14807 9067
rect 334 8844 14666 8927
rect 334 8780 349 8844
rect 413 8780 430 8844
rect 494 8780 510 8844
rect 574 8780 590 8844
rect 654 8780 670 8844
rect 734 8780 750 8844
rect 814 8780 830 8844
rect 894 8780 910 8844
rect 974 8780 990 8844
rect 1054 8780 1070 8844
rect 1134 8780 1150 8844
rect 1214 8780 1230 8844
rect 1294 8780 1310 8844
rect 1374 8780 1390 8844
rect 1454 8780 1470 8844
rect 1534 8780 1550 8844
rect 1614 8780 1630 8844
rect 1694 8780 1710 8844
rect 1774 8780 1790 8844
rect 1854 8780 1870 8844
rect 1934 8780 1950 8844
rect 2014 8780 2030 8844
rect 2094 8780 2110 8844
rect 2174 8780 2190 8844
rect 2254 8780 2270 8844
rect 2334 8780 2350 8844
rect 2414 8780 2430 8844
rect 2494 8780 2510 8844
rect 2574 8780 2590 8844
rect 2654 8780 2670 8844
rect 2734 8780 2750 8844
rect 2814 8780 2830 8844
rect 2894 8780 2910 8844
rect 2974 8780 2990 8844
rect 3054 8780 3070 8844
rect 3134 8780 3150 8844
rect 3214 8780 3230 8844
rect 3294 8780 3310 8844
rect 3374 8780 3390 8844
rect 3454 8780 3470 8844
rect 3534 8780 3550 8844
rect 3614 8780 3630 8844
rect 3694 8780 3710 8844
rect 3774 8780 3790 8844
rect 3854 8780 3870 8844
rect 3934 8780 3950 8844
rect 4014 8780 4030 8844
rect 4094 8780 4110 8844
rect 4174 8780 4190 8844
rect 4254 8780 4270 8844
rect 4334 8780 4350 8844
rect 4414 8780 4430 8844
rect 4494 8780 4510 8844
rect 4574 8780 4590 8844
rect 4654 8780 4670 8844
rect 4734 8780 4750 8844
rect 4814 8780 4830 8844
rect 4894 8780 14666 8844
rect 334 8758 14666 8780
rect 334 8694 349 8758
rect 413 8694 430 8758
rect 494 8694 510 8758
rect 574 8694 590 8758
rect 654 8694 670 8758
rect 734 8694 750 8758
rect 814 8694 830 8758
rect 894 8694 910 8758
rect 974 8694 990 8758
rect 1054 8694 1070 8758
rect 1134 8694 1150 8758
rect 1214 8694 1230 8758
rect 1294 8694 1310 8758
rect 1374 8694 1390 8758
rect 1454 8694 1470 8758
rect 1534 8694 1550 8758
rect 1614 8694 1630 8758
rect 1694 8694 1710 8758
rect 1774 8694 1790 8758
rect 1854 8694 1870 8758
rect 1934 8694 1950 8758
rect 2014 8694 2030 8758
rect 2094 8694 2110 8758
rect 2174 8694 2190 8758
rect 2254 8694 2270 8758
rect 2334 8694 2350 8758
rect 2414 8694 2430 8758
rect 2494 8694 2510 8758
rect 2574 8694 2590 8758
rect 2654 8694 2670 8758
rect 2734 8694 2750 8758
rect 2814 8694 2830 8758
rect 2894 8694 2910 8758
rect 2974 8694 2990 8758
rect 3054 8694 3070 8758
rect 3134 8694 3150 8758
rect 3214 8694 3230 8758
rect 3294 8694 3310 8758
rect 3374 8694 3390 8758
rect 3454 8694 3470 8758
rect 3534 8694 3550 8758
rect 3614 8694 3630 8758
rect 3694 8694 3710 8758
rect 3774 8694 3790 8758
rect 3854 8694 3870 8758
rect 3934 8694 3950 8758
rect 4014 8694 4030 8758
rect 4094 8694 4110 8758
rect 4174 8694 4190 8758
rect 4254 8694 4270 8758
rect 4334 8694 4350 8758
rect 4414 8694 4430 8758
rect 4494 8694 4510 8758
rect 4574 8694 4590 8758
rect 4654 8694 4670 8758
rect 4734 8694 4750 8758
rect 4814 8694 4830 8758
rect 4894 8694 14666 8758
rect 334 8672 14666 8694
rect 334 8608 349 8672
rect 413 8608 430 8672
rect 494 8608 510 8672
rect 574 8608 590 8672
rect 654 8608 670 8672
rect 734 8608 750 8672
rect 814 8608 830 8672
rect 894 8608 910 8672
rect 974 8608 990 8672
rect 1054 8608 1070 8672
rect 1134 8608 1150 8672
rect 1214 8608 1230 8672
rect 1294 8608 1310 8672
rect 1374 8608 1390 8672
rect 1454 8608 1470 8672
rect 1534 8608 1550 8672
rect 1614 8608 1630 8672
rect 1694 8608 1710 8672
rect 1774 8608 1790 8672
rect 1854 8608 1870 8672
rect 1934 8608 1950 8672
rect 2014 8608 2030 8672
rect 2094 8608 2110 8672
rect 2174 8608 2190 8672
rect 2254 8608 2270 8672
rect 2334 8608 2350 8672
rect 2414 8608 2430 8672
rect 2494 8608 2510 8672
rect 2574 8608 2590 8672
rect 2654 8608 2670 8672
rect 2734 8608 2750 8672
rect 2814 8608 2830 8672
rect 2894 8608 2910 8672
rect 2974 8608 2990 8672
rect 3054 8608 3070 8672
rect 3134 8608 3150 8672
rect 3214 8608 3230 8672
rect 3294 8608 3310 8672
rect 3374 8608 3390 8672
rect 3454 8608 3470 8672
rect 3534 8608 3550 8672
rect 3614 8608 3630 8672
rect 3694 8608 3710 8672
rect 3774 8608 3790 8672
rect 3854 8608 3870 8672
rect 3934 8608 3950 8672
rect 4014 8608 4030 8672
rect 4094 8608 4110 8672
rect 4174 8608 4190 8672
rect 4254 8608 4270 8672
rect 4334 8608 4350 8672
rect 4414 8608 4430 8672
rect 4494 8608 4510 8672
rect 4574 8608 4590 8672
rect 4654 8608 4670 8672
rect 4734 8608 4750 8672
rect 4814 8608 4830 8672
rect 4894 8608 14666 8672
rect 334 8586 14666 8608
rect 334 8522 349 8586
rect 413 8522 430 8586
rect 494 8522 510 8586
rect 574 8522 590 8586
rect 654 8522 670 8586
rect 734 8522 750 8586
rect 814 8522 830 8586
rect 894 8522 910 8586
rect 974 8522 990 8586
rect 1054 8522 1070 8586
rect 1134 8522 1150 8586
rect 1214 8522 1230 8586
rect 1294 8522 1310 8586
rect 1374 8522 1390 8586
rect 1454 8522 1470 8586
rect 1534 8522 1550 8586
rect 1614 8522 1630 8586
rect 1694 8522 1710 8586
rect 1774 8522 1790 8586
rect 1854 8522 1870 8586
rect 1934 8522 1950 8586
rect 2014 8522 2030 8586
rect 2094 8522 2110 8586
rect 2174 8522 2190 8586
rect 2254 8522 2270 8586
rect 2334 8522 2350 8586
rect 2414 8522 2430 8586
rect 2494 8522 2510 8586
rect 2574 8522 2590 8586
rect 2654 8522 2670 8586
rect 2734 8522 2750 8586
rect 2814 8522 2830 8586
rect 2894 8522 2910 8586
rect 2974 8522 2990 8586
rect 3054 8522 3070 8586
rect 3134 8522 3150 8586
rect 3214 8522 3230 8586
rect 3294 8522 3310 8586
rect 3374 8522 3390 8586
rect 3454 8522 3470 8586
rect 3534 8522 3550 8586
rect 3614 8522 3630 8586
rect 3694 8522 3710 8586
rect 3774 8522 3790 8586
rect 3854 8522 3870 8586
rect 3934 8522 3950 8586
rect 4014 8522 4030 8586
rect 4094 8522 4110 8586
rect 4174 8522 4190 8586
rect 4254 8522 4270 8586
rect 4334 8522 4350 8586
rect 4414 8522 4430 8586
rect 4494 8522 4510 8586
rect 4574 8522 4590 8586
rect 4654 8522 4670 8586
rect 4734 8522 4750 8586
rect 4814 8522 4830 8586
rect 4894 8522 14666 8586
rect 334 8500 14666 8522
rect 334 8436 349 8500
rect 413 8436 430 8500
rect 494 8436 510 8500
rect 574 8436 590 8500
rect 654 8436 670 8500
rect 734 8436 750 8500
rect 814 8436 830 8500
rect 894 8436 910 8500
rect 974 8436 990 8500
rect 1054 8436 1070 8500
rect 1134 8436 1150 8500
rect 1214 8436 1230 8500
rect 1294 8436 1310 8500
rect 1374 8436 1390 8500
rect 1454 8436 1470 8500
rect 1534 8436 1550 8500
rect 1614 8436 1630 8500
rect 1694 8436 1710 8500
rect 1774 8436 1790 8500
rect 1854 8436 1870 8500
rect 1934 8436 1950 8500
rect 2014 8436 2030 8500
rect 2094 8436 2110 8500
rect 2174 8436 2190 8500
rect 2254 8436 2270 8500
rect 2334 8436 2350 8500
rect 2414 8436 2430 8500
rect 2494 8436 2510 8500
rect 2574 8436 2590 8500
rect 2654 8436 2670 8500
rect 2734 8436 2750 8500
rect 2814 8436 2830 8500
rect 2894 8436 2910 8500
rect 2974 8436 2990 8500
rect 3054 8436 3070 8500
rect 3134 8436 3150 8500
rect 3214 8436 3230 8500
rect 3294 8436 3310 8500
rect 3374 8436 3390 8500
rect 3454 8436 3470 8500
rect 3534 8436 3550 8500
rect 3614 8436 3630 8500
rect 3694 8436 3710 8500
rect 3774 8436 3790 8500
rect 3854 8436 3870 8500
rect 3934 8436 3950 8500
rect 4014 8436 4030 8500
rect 4094 8436 4110 8500
rect 4174 8436 4190 8500
rect 4254 8436 4270 8500
rect 4334 8436 4350 8500
rect 4414 8436 4430 8500
rect 4494 8436 4510 8500
rect 4574 8436 4590 8500
rect 4654 8436 4670 8500
rect 4734 8436 4750 8500
rect 4814 8436 4830 8500
rect 4894 8436 14666 8500
rect 334 8414 14666 8436
rect 334 8350 349 8414
rect 413 8350 430 8414
rect 494 8350 510 8414
rect 574 8350 590 8414
rect 654 8350 670 8414
rect 734 8350 750 8414
rect 814 8350 830 8414
rect 894 8350 910 8414
rect 974 8350 990 8414
rect 1054 8350 1070 8414
rect 1134 8350 1150 8414
rect 1214 8350 1230 8414
rect 1294 8350 1310 8414
rect 1374 8350 1390 8414
rect 1454 8350 1470 8414
rect 1534 8350 1550 8414
rect 1614 8350 1630 8414
rect 1694 8350 1710 8414
rect 1774 8350 1790 8414
rect 1854 8350 1870 8414
rect 1934 8350 1950 8414
rect 2014 8350 2030 8414
rect 2094 8350 2110 8414
rect 2174 8350 2190 8414
rect 2254 8350 2270 8414
rect 2334 8350 2350 8414
rect 2414 8350 2430 8414
rect 2494 8350 2510 8414
rect 2574 8350 2590 8414
rect 2654 8350 2670 8414
rect 2734 8350 2750 8414
rect 2814 8350 2830 8414
rect 2894 8350 2910 8414
rect 2974 8350 2990 8414
rect 3054 8350 3070 8414
rect 3134 8350 3150 8414
rect 3214 8350 3230 8414
rect 3294 8350 3310 8414
rect 3374 8350 3390 8414
rect 3454 8350 3470 8414
rect 3534 8350 3550 8414
rect 3614 8350 3630 8414
rect 3694 8350 3710 8414
rect 3774 8350 3790 8414
rect 3854 8350 3870 8414
rect 3934 8350 3950 8414
rect 4014 8350 4030 8414
rect 4094 8350 4110 8414
rect 4174 8350 4190 8414
rect 4254 8350 4270 8414
rect 4334 8350 4350 8414
rect 4414 8350 4430 8414
rect 4494 8350 4510 8414
rect 4574 8350 4590 8414
rect 4654 8350 4670 8414
rect 4734 8350 4750 8414
rect 4814 8350 4830 8414
rect 4894 8350 14666 8414
rect 334 8328 14666 8350
rect 334 8264 349 8328
rect 413 8264 430 8328
rect 494 8264 510 8328
rect 574 8264 590 8328
rect 654 8264 670 8328
rect 734 8264 750 8328
rect 814 8264 830 8328
rect 894 8264 910 8328
rect 974 8264 990 8328
rect 1054 8264 1070 8328
rect 1134 8264 1150 8328
rect 1214 8264 1230 8328
rect 1294 8264 1310 8328
rect 1374 8264 1390 8328
rect 1454 8264 1470 8328
rect 1534 8264 1550 8328
rect 1614 8264 1630 8328
rect 1694 8264 1710 8328
rect 1774 8264 1790 8328
rect 1854 8264 1870 8328
rect 1934 8264 1950 8328
rect 2014 8264 2030 8328
rect 2094 8264 2110 8328
rect 2174 8264 2190 8328
rect 2254 8264 2270 8328
rect 2334 8264 2350 8328
rect 2414 8264 2430 8328
rect 2494 8264 2510 8328
rect 2574 8264 2590 8328
rect 2654 8264 2670 8328
rect 2734 8264 2750 8328
rect 2814 8264 2830 8328
rect 2894 8264 2910 8328
rect 2974 8264 2990 8328
rect 3054 8264 3070 8328
rect 3134 8264 3150 8328
rect 3214 8264 3230 8328
rect 3294 8264 3310 8328
rect 3374 8264 3390 8328
rect 3454 8264 3470 8328
rect 3534 8264 3550 8328
rect 3614 8264 3630 8328
rect 3694 8264 3710 8328
rect 3774 8264 3790 8328
rect 3854 8264 3870 8328
rect 3934 8264 3950 8328
rect 4014 8264 4030 8328
rect 4094 8264 4110 8328
rect 4174 8264 4190 8328
rect 4254 8264 4270 8328
rect 4334 8264 4350 8328
rect 4414 8264 4430 8328
rect 4494 8264 4510 8328
rect 4574 8264 4590 8328
rect 4654 8264 4670 8328
rect 4734 8264 4750 8328
rect 4814 8264 4830 8328
rect 4894 8264 14666 8328
rect 334 8242 14666 8264
rect 334 8178 349 8242
rect 413 8178 430 8242
rect 494 8178 510 8242
rect 574 8178 590 8242
rect 654 8178 670 8242
rect 734 8178 750 8242
rect 814 8178 830 8242
rect 894 8178 910 8242
rect 974 8178 990 8242
rect 1054 8178 1070 8242
rect 1134 8178 1150 8242
rect 1214 8178 1230 8242
rect 1294 8178 1310 8242
rect 1374 8178 1390 8242
rect 1454 8178 1470 8242
rect 1534 8178 1550 8242
rect 1614 8178 1630 8242
rect 1694 8178 1710 8242
rect 1774 8178 1790 8242
rect 1854 8178 1870 8242
rect 1934 8178 1950 8242
rect 2014 8178 2030 8242
rect 2094 8178 2110 8242
rect 2174 8178 2190 8242
rect 2254 8178 2270 8242
rect 2334 8178 2350 8242
rect 2414 8178 2430 8242
rect 2494 8178 2510 8242
rect 2574 8178 2590 8242
rect 2654 8178 2670 8242
rect 2734 8178 2750 8242
rect 2814 8178 2830 8242
rect 2894 8178 2910 8242
rect 2974 8178 2990 8242
rect 3054 8178 3070 8242
rect 3134 8178 3150 8242
rect 3214 8178 3230 8242
rect 3294 8178 3310 8242
rect 3374 8178 3390 8242
rect 3454 8178 3470 8242
rect 3534 8178 3550 8242
rect 3614 8178 3630 8242
rect 3694 8178 3710 8242
rect 3774 8178 3790 8242
rect 3854 8178 3870 8242
rect 3934 8178 3950 8242
rect 4014 8178 4030 8242
rect 4094 8178 4110 8242
rect 4174 8178 4190 8242
rect 4254 8178 4270 8242
rect 4334 8178 4350 8242
rect 4414 8178 4430 8242
rect 4494 8178 4510 8242
rect 4574 8178 4590 8242
rect 4654 8178 4670 8242
rect 4734 8178 4750 8242
rect 4814 8178 4830 8242
rect 4894 8178 14666 8242
rect 334 8156 14666 8178
rect 334 8092 349 8156
rect 413 8092 430 8156
rect 494 8092 510 8156
rect 574 8092 590 8156
rect 654 8092 670 8156
rect 734 8092 750 8156
rect 814 8092 830 8156
rect 894 8092 910 8156
rect 974 8092 990 8156
rect 1054 8092 1070 8156
rect 1134 8092 1150 8156
rect 1214 8092 1230 8156
rect 1294 8092 1310 8156
rect 1374 8092 1390 8156
rect 1454 8092 1470 8156
rect 1534 8092 1550 8156
rect 1614 8092 1630 8156
rect 1694 8092 1710 8156
rect 1774 8092 1790 8156
rect 1854 8092 1870 8156
rect 1934 8092 1950 8156
rect 2014 8092 2030 8156
rect 2094 8092 2110 8156
rect 2174 8092 2190 8156
rect 2254 8092 2270 8156
rect 2334 8092 2350 8156
rect 2414 8092 2430 8156
rect 2494 8092 2510 8156
rect 2574 8092 2590 8156
rect 2654 8092 2670 8156
rect 2734 8092 2750 8156
rect 2814 8092 2830 8156
rect 2894 8092 2910 8156
rect 2974 8092 2990 8156
rect 3054 8092 3070 8156
rect 3134 8092 3150 8156
rect 3214 8092 3230 8156
rect 3294 8092 3310 8156
rect 3374 8092 3390 8156
rect 3454 8092 3470 8156
rect 3534 8092 3550 8156
rect 3614 8092 3630 8156
rect 3694 8092 3710 8156
rect 3774 8092 3790 8156
rect 3854 8092 3870 8156
rect 3934 8092 3950 8156
rect 4014 8092 4030 8156
rect 4094 8092 4110 8156
rect 4174 8092 4190 8156
rect 4254 8092 4270 8156
rect 4334 8092 4350 8156
rect 4414 8092 4430 8156
rect 4494 8092 4510 8156
rect 4574 8092 4590 8156
rect 4654 8092 4670 8156
rect 4734 8092 4750 8156
rect 4814 8092 4830 8156
rect 4894 8092 14666 8156
rect 334 8070 14666 8092
rect 334 8006 349 8070
rect 413 8006 430 8070
rect 494 8006 510 8070
rect 574 8006 590 8070
rect 654 8006 670 8070
rect 734 8006 750 8070
rect 814 8006 830 8070
rect 894 8006 910 8070
rect 974 8006 990 8070
rect 1054 8006 1070 8070
rect 1134 8006 1150 8070
rect 1214 8006 1230 8070
rect 1294 8006 1310 8070
rect 1374 8006 1390 8070
rect 1454 8006 1470 8070
rect 1534 8006 1550 8070
rect 1614 8006 1630 8070
rect 1694 8006 1710 8070
rect 1774 8006 1790 8070
rect 1854 8006 1870 8070
rect 1934 8006 1950 8070
rect 2014 8006 2030 8070
rect 2094 8006 2110 8070
rect 2174 8006 2190 8070
rect 2254 8006 2270 8070
rect 2334 8006 2350 8070
rect 2414 8006 2430 8070
rect 2494 8006 2510 8070
rect 2574 8006 2590 8070
rect 2654 8006 2670 8070
rect 2734 8006 2750 8070
rect 2814 8006 2830 8070
rect 2894 8006 2910 8070
rect 2974 8006 2990 8070
rect 3054 8006 3070 8070
rect 3134 8006 3150 8070
rect 3214 8006 3230 8070
rect 3294 8006 3310 8070
rect 3374 8006 3390 8070
rect 3454 8006 3470 8070
rect 3534 8006 3550 8070
rect 3614 8006 3630 8070
rect 3694 8006 3710 8070
rect 3774 8006 3790 8070
rect 3854 8006 3870 8070
rect 3934 8006 3950 8070
rect 4014 8006 4030 8070
rect 4094 8006 4110 8070
rect 4174 8006 4190 8070
rect 4254 8006 4270 8070
rect 4334 8006 4350 8070
rect 4414 8006 4430 8070
rect 4494 8006 4510 8070
rect 4574 8006 4590 8070
rect 4654 8006 4670 8070
rect 4734 8006 4750 8070
rect 4814 8006 4830 8070
rect 4894 8006 14666 8070
rect 334 7984 14666 8006
rect 334 7920 349 7984
rect 413 7920 430 7984
rect 494 7920 510 7984
rect 574 7920 590 7984
rect 654 7920 670 7984
rect 734 7920 750 7984
rect 814 7920 830 7984
rect 894 7920 910 7984
rect 974 7920 990 7984
rect 1054 7920 1070 7984
rect 1134 7920 1150 7984
rect 1214 7920 1230 7984
rect 1294 7920 1310 7984
rect 1374 7920 1390 7984
rect 1454 7920 1470 7984
rect 1534 7920 1550 7984
rect 1614 7920 1630 7984
rect 1694 7920 1710 7984
rect 1774 7920 1790 7984
rect 1854 7920 1870 7984
rect 1934 7920 1950 7984
rect 2014 7920 2030 7984
rect 2094 7920 2110 7984
rect 2174 7920 2190 7984
rect 2254 7920 2270 7984
rect 2334 7920 2350 7984
rect 2414 7920 2430 7984
rect 2494 7920 2510 7984
rect 2574 7920 2590 7984
rect 2654 7920 2670 7984
rect 2734 7920 2750 7984
rect 2814 7920 2830 7984
rect 2894 7920 2910 7984
rect 2974 7920 2990 7984
rect 3054 7920 3070 7984
rect 3134 7920 3150 7984
rect 3214 7920 3230 7984
rect 3294 7920 3310 7984
rect 3374 7920 3390 7984
rect 3454 7920 3470 7984
rect 3534 7920 3550 7984
rect 3614 7920 3630 7984
rect 3694 7920 3710 7984
rect 3774 7920 3790 7984
rect 3854 7920 3870 7984
rect 3934 7920 3950 7984
rect 4014 7920 4030 7984
rect 4094 7920 4110 7984
rect 4174 7920 4190 7984
rect 4254 7920 4270 7984
rect 4334 7920 4350 7984
rect 4414 7920 4430 7984
rect 4494 7920 4510 7984
rect 4574 7920 4590 7984
rect 4654 7920 4670 7984
rect 4734 7920 4750 7984
rect 4814 7920 4830 7984
rect 4894 7920 14666 7984
rect 334 7837 14666 7920
rect 193 7717 14807 7837
rect 334 6867 14666 7717
rect 193 6747 14807 6867
rect 334 5897 14666 6747
rect 193 5777 14807 5897
rect 334 4687 14666 5777
rect 193 4567 14807 4687
rect 334 3477 14666 4567
rect 193 3357 14807 3477
rect 273 2507 14727 3357
rect 193 2387 14807 2507
rect 334 1297 14666 2387
rect 193 1177 14807 1297
rect 334 7 14666 1177
<< metal5 >>
rect 0 34757 254 39600
rect 14746 34757 15000 39600
rect 0 13607 254 18597
rect 0 12437 254 13287
rect 0 11267 254 12117
rect 0 9147 254 10947
rect 0 7937 254 8827
rect 0 6968 254 7617
rect 14746 13607 15000 18597
rect 14746 12437 15000 13287
rect 14746 11267 15000 12117
rect 14746 9147 15000 10947
rect 14746 7937 15000 8827
rect 14746 6968 15000 7617
rect 0 5997 254 6647
rect 0 4787 254 5677
rect 0 3577 254 4467
rect 14746 5997 15000 6647
rect 14746 4787 15000 5677
rect 14746 3577 15000 4467
rect 0 2607 193 3257
rect 14807 2607 15000 3257
rect 0 1397 254 2287
rect 0 27 254 1077
rect 14746 1397 15000 2287
rect 14746 27 15000 1077
<< obsm5 >>
rect 574 34437 14426 39600
rect 0 18917 15000 34437
rect 574 6968 14426 18917
rect 0 6967 15000 6968
rect 574 3257 14426 6967
rect 513 2607 14487 3257
rect 574 27 14426 2607
<< labels >>
rlabel metal5 s 0 9147 254 10947 6 VSSA
port 1 nsew ground bidirectional
rlabel metal5 s 0 6968 254 7617 6 VSSA
port 1 nsew ground bidirectional
rlabel metal5 s 14746 9147 15000 10947 6 VSSA
port 1 nsew ground bidirectional
rlabel metal5 s 14746 6968 15000 7617 6 VSSA
port 1 nsew ground bidirectional
rlabel metal4 s 0 10881 15000 10947 6 VSSA
port 1 nsew ground bidirectional
rlabel metal4 s 0 9147 15000 9213 6 VSSA
port 1 nsew ground bidirectional
rlabel metal4 s 0 9929 254 10165 6 VSSA
port 1 nsew ground bidirectional
rlabel metal4 s 0 6947 254 7637 6 VSSA
port 1 nsew ground bidirectional
rlabel metal4 s 14746 9929 15000 10165 6 VSSA
port 1 nsew ground bidirectional
rlabel metal4 s 14746 6947 15000 7637 6 VSSA
port 1 nsew ground bidirectional
rlabel metal5 s 0 13607 254 18597 6 VDDIO
port 2 nsew power bidirectional
rlabel metal5 s 0 3577 254 4467 6 VDDIO
port 2 nsew power bidirectional
rlabel metal5 s 14746 13607 15000 18597 6 VDDIO
port 2 nsew power bidirectional
rlabel metal5 s 14746 3577 15000 4467 6 VDDIO
port 2 nsew power bidirectional
rlabel metal4 s 0 3557 254 4487 6 VDDIO
port 2 nsew power bidirectional
rlabel metal4 s 0 13607 254 18600 6 VDDIO
port 2 nsew power bidirectional
rlabel metal4 s 14746 3557 15000 4487 6 VDDIO
port 2 nsew power bidirectional
rlabel metal4 s 14746 13607 15000 18600 6 VDDIO
port 2 nsew power bidirectional
rlabel metal5 s 0 12437 254 13287 6 VDDIO_Q
port 3 nsew power bidirectional
rlabel metal5 s 14746 12437 15000 13287 6 VDDIO_Q
port 3 nsew power bidirectional
rlabel metal4 s 0 12417 254 13307 6 VDDIO_Q
port 3 nsew power bidirectional
rlabel metal4 s 14746 12417 15000 13307 6 VDDIO_Q
port 3 nsew power bidirectional
rlabel metal5 s 0 7937 254 8827 6 VSSD
port 4 nsew ground bidirectional
rlabel metal5 s 14746 7937 15000 8827 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 0 7917 254 8847 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 14746 7917 15000 8847 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 10151 7918 14940 8846 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 14882 8792 14922 8832 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 14882 8706 14922 8746 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 14882 8620 14922 8660 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 14882 8534 14922 8574 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 14882 8448 14922 8488 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 14882 8362 14922 8402 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 14882 8276 14922 8316 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 14882 8190 14922 8230 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 14882 8104 14922 8144 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 14882 8018 14922 8058 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 14882 7932 14922 7972 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 14801 8792 14841 8832 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 14801 8706 14841 8746 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 14801 8620 14841 8660 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 14801 8534 14841 8574 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 14801 8448 14841 8488 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 14801 8362 14841 8402 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 14801 8276 14841 8316 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 14801 8190 14841 8230 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 14801 8104 14841 8144 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 14801 8018 14841 8058 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 14801 7932 14841 7972 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 14720 8792 14760 8832 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 14720 8706 14760 8746 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 14720 8620 14760 8660 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 14720 8534 14760 8574 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 14720 8448 14760 8488 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 14720 8362 14760 8402 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 14720 8276 14760 8316 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 14720 8190 14760 8230 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 14720 8104 14760 8144 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 14720 8018 14760 8058 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 14720 7932 14760 7972 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 14639 8792 14679 8832 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 14639 8706 14679 8746 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 14639 8620 14679 8660 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 14639 8534 14679 8574 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 14639 8448 14679 8488 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 14639 8362 14679 8402 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 14639 8276 14679 8316 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 14639 8190 14679 8230 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 14639 8104 14679 8144 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 14639 8018 14679 8058 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 14639 7932 14679 7972 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 14558 8792 14598 8832 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 14558 8706 14598 8746 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 14558 8620 14598 8660 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 14558 8534 14598 8574 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 14558 8448 14598 8488 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 14558 8362 14598 8402 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 14558 8276 14598 8316 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 14558 8190 14598 8230 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 14558 8104 14598 8144 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 14558 8018 14598 8058 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 14558 7932 14598 7972 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 14477 8792 14517 8832 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 14477 8706 14517 8746 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 14477 8620 14517 8660 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 14477 8534 14517 8574 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 14477 8448 14517 8488 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 14477 8362 14517 8402 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 14477 8276 14517 8316 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 14477 8190 14517 8230 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 14477 8104 14517 8144 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 14477 8018 14517 8058 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 14477 7932 14517 7972 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 14396 8792 14436 8832 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 14396 8706 14436 8746 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 14396 8620 14436 8660 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 14396 8534 14436 8574 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 14396 8448 14436 8488 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 14396 8362 14436 8402 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 14396 8276 14436 8316 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 14396 8190 14436 8230 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 14396 8104 14436 8144 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 14396 8018 14436 8058 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 14396 7932 14436 7972 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 14315 8792 14355 8832 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 14315 8706 14355 8746 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 14315 8620 14355 8660 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 14315 8534 14355 8574 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 14315 8448 14355 8488 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 14315 8362 14355 8402 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 14315 8276 14355 8316 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 14315 8190 14355 8230 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 14315 8104 14355 8144 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 14315 8018 14355 8058 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 14315 7932 14355 7972 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 14234 8792 14274 8832 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 14234 8706 14274 8746 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 14234 8620 14274 8660 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 14234 8534 14274 8574 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 14234 8448 14274 8488 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 14234 8362 14274 8402 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 14234 8276 14274 8316 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 14234 8190 14274 8230 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 14234 8104 14274 8144 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 14234 8018 14274 8058 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 14234 7932 14274 7972 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 14153 8792 14193 8832 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 14153 8706 14193 8746 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 14153 8620 14193 8660 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 14153 8534 14193 8574 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 14153 8448 14193 8488 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 14153 8362 14193 8402 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 14153 8276 14193 8316 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 14153 8190 14193 8230 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 14153 8104 14193 8144 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 14153 8018 14193 8058 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 14153 7932 14193 7972 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 14072 8792 14112 8832 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 14072 8706 14112 8746 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 14072 8620 14112 8660 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 14072 8534 14112 8574 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 14072 8448 14112 8488 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 14072 8362 14112 8402 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 14072 8276 14112 8316 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 14072 8190 14112 8230 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 14072 8104 14112 8144 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 14072 8018 14112 8058 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 14072 7932 14112 7972 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13991 8792 14031 8832 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13991 8706 14031 8746 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13991 8620 14031 8660 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13991 8534 14031 8574 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13991 8448 14031 8488 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13991 8362 14031 8402 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13991 8276 14031 8316 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13991 8190 14031 8230 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13991 8104 14031 8144 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13991 8018 14031 8058 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13991 7932 14031 7972 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13910 8792 13950 8832 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13910 8706 13950 8746 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13910 8620 13950 8660 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13910 8534 13950 8574 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13910 8448 13950 8488 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13910 8362 13950 8402 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13910 8276 13950 8316 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13910 8190 13950 8230 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13910 8104 13950 8144 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13910 8018 13950 8058 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13910 7932 13950 7972 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13829 8792 13869 8832 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13829 8706 13869 8746 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13829 8620 13869 8660 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13829 8534 13869 8574 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13829 8448 13869 8488 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13829 8362 13869 8402 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13829 8276 13869 8316 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13829 8190 13869 8230 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13829 8104 13869 8144 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13829 8018 13869 8058 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13829 7932 13869 7972 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13748 8792 13788 8832 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13748 8706 13788 8746 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13748 8620 13788 8660 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13748 8534 13788 8574 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13748 8448 13788 8488 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13748 8362 13788 8402 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13748 8276 13788 8316 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13748 8190 13788 8230 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13748 8104 13788 8144 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13748 8018 13788 8058 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13748 7932 13788 7972 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13667 8792 13707 8832 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13667 8706 13707 8746 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13667 8620 13707 8660 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13667 8534 13707 8574 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13667 8448 13707 8488 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13667 8362 13707 8402 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13667 8276 13707 8316 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13667 8190 13707 8230 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13667 8104 13707 8144 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13667 8018 13707 8058 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13667 7932 13707 7972 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13586 8792 13626 8832 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13586 8706 13626 8746 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13586 8620 13626 8660 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13586 8534 13626 8574 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13586 8448 13626 8488 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13586 8362 13626 8402 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13586 8276 13626 8316 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13586 8190 13626 8230 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13586 8104 13626 8144 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13586 8018 13626 8058 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13586 7932 13626 7972 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13505 8792 13545 8832 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13505 8706 13545 8746 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13505 8620 13545 8660 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13505 8534 13545 8574 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13505 8448 13545 8488 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13505 8362 13545 8402 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13505 8276 13545 8316 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13505 8190 13545 8230 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13505 8104 13545 8144 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13505 8018 13545 8058 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13505 7932 13545 7972 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13424 8792 13464 8832 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13424 8706 13464 8746 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13424 8620 13464 8660 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13424 8534 13464 8574 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13424 8448 13464 8488 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13424 8362 13464 8402 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13424 8276 13464 8316 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13424 8190 13464 8230 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13424 8104 13464 8144 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13424 8018 13464 8058 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13424 7932 13464 7972 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13343 8792 13383 8832 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13343 8706 13383 8746 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13343 8620 13383 8660 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13343 8534 13383 8574 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13343 8448 13383 8488 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13343 8362 13383 8402 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13343 8276 13383 8316 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13343 8190 13383 8230 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13343 8104 13383 8144 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13343 8018 13383 8058 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13343 7932 13383 7972 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13262 8792 13302 8832 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13262 8706 13302 8746 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13262 8620 13302 8660 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13262 8534 13302 8574 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13262 8448 13302 8488 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13262 8362 13302 8402 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13262 8276 13302 8316 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13262 8190 13302 8230 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13262 8104 13302 8144 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13262 8018 13302 8058 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13262 7932 13302 7972 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13181 8792 13221 8832 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13181 8706 13221 8746 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13181 8620 13221 8660 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13181 8534 13221 8574 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13181 8448 13221 8488 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13181 8362 13221 8402 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13181 8276 13221 8316 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13181 8190 13221 8230 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13181 8104 13221 8144 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13181 8018 13221 8058 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13181 7932 13221 7972 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13100 8792 13140 8832 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13100 8706 13140 8746 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13100 8620 13140 8660 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13100 8534 13140 8574 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13100 8448 13140 8488 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13100 8362 13140 8402 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13100 8276 13140 8316 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13100 8190 13140 8230 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13100 8104 13140 8144 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13100 8018 13140 8058 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13100 7932 13140 7972 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13019 8792 13059 8832 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13019 8706 13059 8746 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13019 8620 13059 8660 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13019 8534 13059 8574 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13019 8448 13059 8488 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13019 8362 13059 8402 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13019 8276 13059 8316 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13019 8190 13059 8230 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13019 8104 13059 8144 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13019 8018 13059 8058 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 13019 7932 13059 7972 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 12938 8792 12978 8832 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 12938 8706 12978 8746 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 12938 8620 12978 8660 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 12938 8534 12978 8574 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 12938 8448 12978 8488 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 12938 8362 12978 8402 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 12938 8276 12978 8316 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 12938 8190 12978 8230 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 12938 8104 12978 8144 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 12938 8018 12978 8058 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 12938 7932 12978 7972 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 12857 8792 12897 8832 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 12857 8706 12897 8746 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 12857 8620 12897 8660 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 12857 8534 12897 8574 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 12857 8448 12897 8488 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 12857 8362 12897 8402 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 12857 8276 12897 8316 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 12857 8190 12897 8230 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 12857 8104 12897 8144 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 12857 8018 12897 8058 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 12857 7932 12897 7972 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 12776 8792 12816 8832 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 12776 8706 12816 8746 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 12776 8620 12816 8660 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 12776 8534 12816 8574 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 12776 8448 12816 8488 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 12776 8362 12816 8402 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 12776 8276 12816 8316 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 12776 8190 12816 8230 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 12776 8104 12816 8144 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 12776 8018 12816 8058 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 12776 7932 12816 7972 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 12695 8792 12735 8832 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 12695 8706 12735 8746 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 12695 8620 12735 8660 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 12695 8534 12735 8574 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 12695 8448 12735 8488 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 12695 8362 12735 8402 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 12695 8276 12735 8316 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 12695 8190 12735 8230 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 12695 8104 12735 8144 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 12695 8018 12735 8058 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 12695 7932 12735 7972 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 12614 8792 12654 8832 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 12614 8706 12654 8746 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 12614 8620 12654 8660 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 12614 8534 12654 8574 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 12614 8448 12654 8488 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 12614 8362 12654 8402 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 12614 8276 12654 8316 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 12614 8190 12654 8230 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 12614 8104 12654 8144 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 12614 8018 12654 8058 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 12614 7932 12654 7972 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 12533 8792 12573 8832 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 12533 8706 12573 8746 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 12533 8620 12573 8660 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 12533 8534 12573 8574 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 12533 8448 12573 8488 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 12533 8362 12573 8402 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 12533 8276 12573 8316 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 12533 8190 12573 8230 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 12533 8104 12573 8144 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 12533 8018 12573 8058 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 12533 7932 12573 7972 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 12452 8792 12492 8832 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 12452 8706 12492 8746 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 12452 8620 12492 8660 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 12452 8534 12492 8574 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 12452 8448 12492 8488 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 12452 8362 12492 8402 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 12452 8276 12492 8316 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 12452 8190 12492 8230 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 12452 8104 12492 8144 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 12452 8018 12492 8058 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 12452 7932 12492 7972 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 12371 8792 12411 8832 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 12371 8706 12411 8746 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 12371 8620 12411 8660 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 12371 8534 12411 8574 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 12371 8448 12411 8488 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 12371 8362 12411 8402 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 12371 8276 12411 8316 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 12371 8190 12411 8230 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 12371 8104 12411 8144 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 12371 8018 12411 8058 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 12371 7932 12411 7972 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 12290 8792 12330 8832 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 12290 8706 12330 8746 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 12290 8620 12330 8660 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 12290 8534 12330 8574 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 12290 8448 12330 8488 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 12290 8362 12330 8402 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 12290 8276 12330 8316 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 12290 8190 12330 8230 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 12290 8104 12330 8144 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 12290 8018 12330 8058 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 12290 7932 12330 7972 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 12209 8792 12249 8832 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 12209 8706 12249 8746 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 12209 8620 12249 8660 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 12209 8534 12249 8574 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 12209 8448 12249 8488 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 12209 8362 12249 8402 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 12209 8276 12249 8316 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 12209 8190 12249 8230 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 12209 8104 12249 8144 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 12209 8018 12249 8058 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 12209 7932 12249 7972 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 12128 8792 12168 8832 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 12128 8706 12168 8746 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 12128 8620 12168 8660 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 12128 8534 12168 8574 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 12128 8448 12168 8488 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 12128 8362 12168 8402 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 12128 8276 12168 8316 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 12128 8190 12168 8230 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 12128 8104 12168 8144 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 12128 8018 12168 8058 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 12128 7932 12168 7972 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 12047 8792 12087 8832 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 12047 8706 12087 8746 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 12047 8620 12087 8660 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 12047 8534 12087 8574 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 12047 8448 12087 8488 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 12047 8362 12087 8402 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 12047 8276 12087 8316 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 12047 8190 12087 8230 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 12047 8104 12087 8144 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 12047 8018 12087 8058 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 12047 7932 12087 7972 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 11966 8792 12006 8832 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 11966 8706 12006 8746 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 11966 8620 12006 8660 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 11966 8534 12006 8574 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 11966 8448 12006 8488 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 11966 8362 12006 8402 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 11966 8276 12006 8316 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 11966 8190 12006 8230 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 11966 8104 12006 8144 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 11966 8018 12006 8058 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 11966 7932 12006 7972 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 11885 8792 11925 8832 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 11885 8706 11925 8746 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 11885 8620 11925 8660 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 11885 8534 11925 8574 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 11885 8448 11925 8488 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 11885 8362 11925 8402 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 11885 8276 11925 8316 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 11885 8190 11925 8230 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 11885 8104 11925 8144 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 11885 8018 11925 8058 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 11885 7932 11925 7972 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 11804 8792 11844 8832 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 11804 8706 11844 8746 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 11804 8620 11844 8660 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 11804 8534 11844 8574 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 11804 8448 11844 8488 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 11804 8362 11844 8402 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 11804 8276 11844 8316 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 11804 8190 11844 8230 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 11804 8104 11844 8144 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 11804 8018 11844 8058 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 11804 7932 11844 7972 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 11723 8792 11763 8832 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 11723 8706 11763 8746 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 11723 8620 11763 8660 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 11723 8534 11763 8574 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 11723 8448 11763 8488 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 11723 8362 11763 8402 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 11723 8276 11763 8316 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 11723 8190 11763 8230 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 11723 8104 11763 8144 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 11723 8018 11763 8058 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 11723 7932 11763 7972 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 11642 8792 11682 8832 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 11642 8706 11682 8746 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 11642 8620 11682 8660 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 11642 8534 11682 8574 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 11642 8448 11682 8488 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 11642 8362 11682 8402 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 11642 8276 11682 8316 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 11642 8190 11682 8230 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 11642 8104 11682 8144 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 11642 8018 11682 8058 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 11642 7932 11682 7972 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 11561 8792 11601 8832 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 11561 8706 11601 8746 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 11561 8620 11601 8660 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 11561 8534 11601 8574 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 11561 8448 11601 8488 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 11561 8362 11601 8402 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 11561 8276 11601 8316 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 11561 8190 11601 8230 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 11561 8104 11601 8144 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 11561 8018 11601 8058 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 11561 7932 11601 7972 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 11480 8792 11520 8832 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 11480 8706 11520 8746 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 11480 8620 11520 8660 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 11480 8534 11520 8574 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 11480 8448 11520 8488 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 11480 8362 11520 8402 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 11480 8276 11520 8316 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 11480 8190 11520 8230 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 11480 8104 11520 8144 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 11480 8018 11520 8058 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 11480 7932 11520 7972 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 11399 8792 11439 8832 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 11399 8706 11439 8746 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 11399 8620 11439 8660 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 11399 8534 11439 8574 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 11399 8448 11439 8488 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 11399 8362 11439 8402 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 11399 8276 11439 8316 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 11399 8190 11439 8230 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 11399 8104 11439 8144 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 11399 8018 11439 8058 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 11399 7932 11439 7972 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 11317 8792 11357 8832 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 11317 8706 11357 8746 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 11317 8620 11357 8660 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 11317 8534 11357 8574 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 11317 8448 11357 8488 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 11317 8362 11357 8402 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 11317 8276 11357 8316 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 11317 8190 11357 8230 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 11317 8104 11357 8144 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 11317 8018 11357 8058 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 11317 7932 11357 7972 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 11235 8792 11275 8832 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 11235 8706 11275 8746 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 11235 8620 11275 8660 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 11235 8534 11275 8574 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 11235 8448 11275 8488 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 11235 8362 11275 8402 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 11235 8276 11275 8316 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 11235 8190 11275 8230 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 11235 8104 11275 8144 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 11235 8018 11275 8058 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 11235 7932 11275 7972 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 11153 8792 11193 8832 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 11153 8706 11193 8746 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 11153 8620 11193 8660 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 11153 8534 11193 8574 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 11153 8448 11193 8488 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 11153 8362 11193 8402 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 11153 8276 11193 8316 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 11153 8190 11193 8230 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 11153 8104 11193 8144 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 11153 8018 11193 8058 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 11153 7932 11193 7972 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 11071 8792 11111 8832 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 11071 8706 11111 8746 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 11071 8620 11111 8660 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 11071 8534 11111 8574 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 11071 8448 11111 8488 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 11071 8362 11111 8402 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 11071 8276 11111 8316 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 11071 8190 11111 8230 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 11071 8104 11111 8144 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 11071 8018 11111 8058 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 11071 7932 11111 7972 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 10989 8792 11029 8832 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 10989 8706 11029 8746 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 10989 8620 11029 8660 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 10989 8534 11029 8574 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 10989 8448 11029 8488 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 10989 8362 11029 8402 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 10989 8276 11029 8316 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 10989 8190 11029 8230 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 10989 8104 11029 8144 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 10989 8018 11029 8058 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 10989 7932 11029 7972 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 10907 8792 10947 8832 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 10907 8706 10947 8746 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 10907 8620 10947 8660 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 10907 8534 10947 8574 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 10907 8448 10947 8488 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 10907 8362 10947 8402 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 10907 8276 10947 8316 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 10907 8190 10947 8230 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 10907 8104 10947 8144 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 10907 8018 10947 8058 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 10907 7932 10947 7972 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 10825 8792 10865 8832 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 10825 8706 10865 8746 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 10825 8620 10865 8660 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 10825 8534 10865 8574 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 10825 8448 10865 8488 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 10825 8362 10865 8402 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 10825 8276 10865 8316 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 10825 8190 10865 8230 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 10825 8104 10865 8144 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 10825 8018 10865 8058 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 10825 7932 10865 7972 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 10743 8792 10783 8832 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 10743 8706 10783 8746 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 10743 8620 10783 8660 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 10743 8534 10783 8574 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 10743 8448 10783 8488 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 10743 8362 10783 8402 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 10743 8276 10783 8316 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 10743 8190 10783 8230 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 10743 8104 10783 8144 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 10743 8018 10783 8058 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 10743 7932 10783 7972 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 10661 8792 10701 8832 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 10661 8706 10701 8746 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 10661 8620 10701 8660 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 10661 8534 10701 8574 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 10661 8448 10701 8488 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 10661 8362 10701 8402 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 10661 8276 10701 8316 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 10661 8190 10701 8230 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 10661 8104 10701 8144 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 10661 8018 10701 8058 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 10661 7932 10701 7972 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 10579 8792 10619 8832 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 10579 8706 10619 8746 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 10579 8620 10619 8660 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 10579 8534 10619 8574 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 10579 8448 10619 8488 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 10579 8362 10619 8402 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 10579 8276 10619 8316 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 10579 8190 10619 8230 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 10579 8104 10619 8144 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 10579 8018 10619 8058 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 10579 7932 10619 7972 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 10497 8792 10537 8832 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 10497 8706 10537 8746 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 10497 8620 10537 8660 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 10497 8534 10537 8574 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 10497 8448 10537 8488 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 10497 8362 10537 8402 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 10497 8276 10537 8316 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 10497 8190 10537 8230 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 10497 8104 10537 8144 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 10497 8018 10537 8058 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 10497 7932 10537 7972 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 10415 8792 10455 8832 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 10415 8706 10455 8746 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 10415 8620 10455 8660 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 10415 8534 10455 8574 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 10415 8448 10455 8488 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 10415 8362 10455 8402 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 10415 8276 10455 8316 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 10415 8190 10455 8230 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 10415 8104 10455 8144 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 10415 8018 10455 8058 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 10415 7932 10455 7972 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 10333 8792 10373 8832 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 10333 8706 10373 8746 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 10333 8620 10373 8660 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 10333 8534 10373 8574 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 10333 8448 10373 8488 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 10333 8362 10373 8402 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 10333 8276 10373 8316 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 10333 8190 10373 8230 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 10333 8104 10373 8144 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 10333 8018 10373 8058 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 10333 7932 10373 7972 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 10251 8792 10291 8832 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 10251 8706 10291 8746 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 10251 8620 10291 8660 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 10251 8534 10291 8574 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 10251 8448 10291 8488 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 10251 8362 10291 8402 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 10251 8276 10291 8316 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 10251 8190 10291 8230 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 10251 8104 10291 8144 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 10251 8018 10291 8058 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 10251 7932 10291 7972 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 10169 8792 10209 8832 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 10169 8706 10209 8746 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 10169 8620 10209 8660 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 10169 8534 10209 8574 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 10169 8448 10209 8488 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 10169 8362 10209 8402 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 10169 8276 10209 8316 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 10169 8190 10209 8230 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 10169 8104 10209 8144 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 10169 8018 10209 8058 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 10169 7932 10209 7972 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 4830 8780 4894 8844 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 4830 8780 4894 8844 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 4830 8694 4894 8758 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 4830 8694 4894 8758 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 4830 8608 4894 8672 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 4830 8608 4894 8672 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 4830 8522 4894 8586 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 4830 8522 4894 8586 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 4830 8436 4894 8500 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 4830 8436 4894 8500 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 4830 8350 4894 8414 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 4830 8350 4894 8414 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 4830 8264 4894 8328 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 4830 8264 4894 8328 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 4830 8178 4894 8242 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 4830 8178 4894 8242 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 4830 8092 4894 8156 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 4830 8092 4894 8156 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 4830 8006 4894 8070 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 4830 8006 4894 8070 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 4830 7920 4894 7984 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 4830 7920 4894 7984 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 4750 8780 4814 8844 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 4750 8780 4814 8844 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 4750 8694 4814 8758 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 4750 8694 4814 8758 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 4750 8608 4814 8672 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 4750 8608 4814 8672 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 4750 8522 4814 8586 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 4750 8522 4814 8586 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 4750 8436 4814 8500 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 4750 8436 4814 8500 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 4750 8350 4814 8414 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 4750 8350 4814 8414 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 4750 8264 4814 8328 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 4750 8264 4814 8328 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 4750 8178 4814 8242 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 4750 8178 4814 8242 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 4750 8092 4814 8156 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 4750 8092 4814 8156 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 4750 8006 4814 8070 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 4750 8006 4814 8070 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 4750 7920 4814 7984 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 4750 7920 4814 7984 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 4670 8780 4734 8844 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 4670 8780 4734 8844 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 4670 8694 4734 8758 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 4670 8694 4734 8758 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 4670 8608 4734 8672 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 4670 8608 4734 8672 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 4670 8522 4734 8586 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 4670 8522 4734 8586 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 4670 8436 4734 8500 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 4670 8436 4734 8500 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 4670 8350 4734 8414 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 4670 8350 4734 8414 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 4670 8264 4734 8328 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 4670 8264 4734 8328 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 4670 8178 4734 8242 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 4670 8178 4734 8242 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 4670 8092 4734 8156 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 4670 8092 4734 8156 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 4670 8006 4734 8070 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 4670 8006 4734 8070 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 4670 7920 4734 7984 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 4670 7920 4734 7984 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 4590 8780 4654 8844 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 4590 8780 4654 8844 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 4590 8694 4654 8758 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 4590 8694 4654 8758 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 4590 8608 4654 8672 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 4590 8608 4654 8672 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 4590 8522 4654 8586 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 4590 8522 4654 8586 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 4590 8436 4654 8500 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 4590 8436 4654 8500 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 4590 8350 4654 8414 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 4590 8350 4654 8414 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 4590 8264 4654 8328 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 4590 8264 4654 8328 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 4590 8178 4654 8242 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 4590 8178 4654 8242 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 4590 8092 4654 8156 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 4590 8092 4654 8156 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 4590 8006 4654 8070 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 4590 8006 4654 8070 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 4590 7920 4654 7984 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 4590 7920 4654 7984 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 4510 8780 4574 8844 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 4510 8780 4574 8844 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 4510 8694 4574 8758 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 4510 8694 4574 8758 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 4510 8608 4574 8672 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 4510 8608 4574 8672 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 4510 8522 4574 8586 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 4510 8522 4574 8586 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 4510 8436 4574 8500 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 4510 8436 4574 8500 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 4510 8350 4574 8414 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 4510 8350 4574 8414 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 4510 8264 4574 8328 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 4510 8264 4574 8328 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 4510 8178 4574 8242 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 4510 8178 4574 8242 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 4510 8092 4574 8156 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 4510 8092 4574 8156 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 4510 8006 4574 8070 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 4510 8006 4574 8070 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 4510 7920 4574 7984 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 4510 7920 4574 7984 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 4430 8780 4494 8844 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 4430 8780 4494 8844 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 4430 8694 4494 8758 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 4430 8694 4494 8758 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 4430 8608 4494 8672 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 4430 8608 4494 8672 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 4430 8522 4494 8586 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 4430 8522 4494 8586 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 4430 8436 4494 8500 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 4430 8436 4494 8500 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 4430 8350 4494 8414 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 4430 8350 4494 8414 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 4430 8264 4494 8328 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 4430 8264 4494 8328 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 4430 8178 4494 8242 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 4430 8178 4494 8242 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 4430 8092 4494 8156 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 4430 8092 4494 8156 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 4430 8006 4494 8070 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 4430 8006 4494 8070 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 4430 7920 4494 7984 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 4430 7920 4494 7984 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 4350 8780 4414 8844 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 4350 8780 4414 8844 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 4350 8694 4414 8758 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 4350 8694 4414 8758 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 4350 8608 4414 8672 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 4350 8608 4414 8672 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 4350 8522 4414 8586 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 4350 8522 4414 8586 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 4350 8436 4414 8500 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 4350 8436 4414 8500 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 4350 8350 4414 8414 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 4350 8350 4414 8414 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 4350 8264 4414 8328 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 4350 8264 4414 8328 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 4350 8178 4414 8242 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 4350 8178 4414 8242 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 4350 8092 4414 8156 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 4350 8092 4414 8156 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 4350 8006 4414 8070 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 4350 8006 4414 8070 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 4350 7920 4414 7984 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 4350 7920 4414 7984 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 4270 8780 4334 8844 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 4270 8780 4334 8844 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 4270 8694 4334 8758 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 4270 8694 4334 8758 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 4270 8608 4334 8672 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 4270 8608 4334 8672 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 4270 8522 4334 8586 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 4270 8522 4334 8586 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 4270 8436 4334 8500 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 4270 8436 4334 8500 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 4270 8350 4334 8414 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 4270 8350 4334 8414 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 4270 8264 4334 8328 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 4270 8264 4334 8328 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 4270 8178 4334 8242 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 4270 8178 4334 8242 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 4270 8092 4334 8156 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 4270 8092 4334 8156 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 4270 8006 4334 8070 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 4270 8006 4334 8070 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 4270 7920 4334 7984 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 4270 7920 4334 7984 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 4190 8780 4254 8844 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 4190 8780 4254 8844 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 4190 8694 4254 8758 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 4190 8694 4254 8758 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 4190 8608 4254 8672 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 4190 8608 4254 8672 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 4190 8522 4254 8586 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 4190 8522 4254 8586 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 4190 8436 4254 8500 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 4190 8436 4254 8500 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 4190 8350 4254 8414 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 4190 8350 4254 8414 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 4190 8264 4254 8328 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 4190 8264 4254 8328 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 4190 8178 4254 8242 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 4190 8178 4254 8242 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 4190 8092 4254 8156 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 4190 8092 4254 8156 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 4190 8006 4254 8070 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 4190 8006 4254 8070 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 4190 7920 4254 7984 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 4190 7920 4254 7984 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 4110 8780 4174 8844 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 4110 8780 4174 8844 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 4110 8694 4174 8758 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 4110 8694 4174 8758 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 4110 8608 4174 8672 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 4110 8608 4174 8672 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 4110 8522 4174 8586 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 4110 8522 4174 8586 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 4110 8436 4174 8500 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 4110 8436 4174 8500 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 4110 8350 4174 8414 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 4110 8350 4174 8414 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 4110 8264 4174 8328 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 4110 8264 4174 8328 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 4110 8178 4174 8242 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 4110 8178 4174 8242 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 4110 8092 4174 8156 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 4110 8092 4174 8156 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 4110 8006 4174 8070 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 4110 8006 4174 8070 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 4110 7920 4174 7984 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 4110 7920 4174 7984 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 4030 8780 4094 8844 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 4030 8780 4094 8844 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 4030 8694 4094 8758 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 4030 8694 4094 8758 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 4030 8608 4094 8672 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 4030 8608 4094 8672 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 4030 8522 4094 8586 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 4030 8522 4094 8586 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 4030 8436 4094 8500 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 4030 8436 4094 8500 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 4030 8350 4094 8414 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 4030 8350 4094 8414 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 4030 8264 4094 8328 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 4030 8264 4094 8328 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 4030 8178 4094 8242 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 4030 8178 4094 8242 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 4030 8092 4094 8156 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 4030 8092 4094 8156 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 4030 8006 4094 8070 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 4030 8006 4094 8070 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 4030 7920 4094 7984 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 4030 7920 4094 7984 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 3950 8780 4014 8844 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 3950 8780 4014 8844 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 3950 8694 4014 8758 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 3950 8694 4014 8758 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 3950 8608 4014 8672 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 3950 8608 4014 8672 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 3950 8522 4014 8586 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 3950 8522 4014 8586 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 3950 8436 4014 8500 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 3950 8436 4014 8500 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 3950 8350 4014 8414 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 3950 8350 4014 8414 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 3950 8264 4014 8328 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 3950 8264 4014 8328 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 3950 8178 4014 8242 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 3950 8178 4014 8242 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 3950 8092 4014 8156 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 3950 8092 4014 8156 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 3950 8006 4014 8070 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 3950 8006 4014 8070 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 3950 7920 4014 7984 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 3950 7920 4014 7984 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 3870 8780 3934 8844 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 3870 8780 3934 8844 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 3870 8694 3934 8758 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 3870 8694 3934 8758 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 3870 8608 3934 8672 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 3870 8608 3934 8672 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 3870 8522 3934 8586 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 3870 8522 3934 8586 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 3870 8436 3934 8500 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 3870 8436 3934 8500 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 3870 8350 3934 8414 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 3870 8350 3934 8414 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 3870 8264 3934 8328 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 3870 8264 3934 8328 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 3870 8178 3934 8242 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 3870 8178 3934 8242 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 3870 8092 3934 8156 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 3870 8092 3934 8156 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 3870 8006 3934 8070 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 3870 8006 3934 8070 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 3870 7920 3934 7984 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 3870 7920 3934 7984 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 3790 8780 3854 8844 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 3790 8780 3854 8844 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 3790 8694 3854 8758 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 3790 8694 3854 8758 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 3790 8608 3854 8672 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 3790 8608 3854 8672 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 3790 8522 3854 8586 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 3790 8522 3854 8586 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 3790 8436 3854 8500 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 3790 8436 3854 8500 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 3790 8350 3854 8414 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 3790 8350 3854 8414 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 3790 8264 3854 8328 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 3790 8264 3854 8328 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 3790 8178 3854 8242 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 3790 8178 3854 8242 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 3790 8092 3854 8156 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 3790 8092 3854 8156 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 3790 8006 3854 8070 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 3790 8006 3854 8070 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 3790 7920 3854 7984 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 3790 7920 3854 7984 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 3710 8780 3774 8844 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 3710 8780 3774 8844 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 3710 8694 3774 8758 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 3710 8694 3774 8758 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 3710 8608 3774 8672 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 3710 8608 3774 8672 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 3710 8522 3774 8586 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 3710 8522 3774 8586 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 3710 8436 3774 8500 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 3710 8436 3774 8500 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 3710 8350 3774 8414 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 3710 8350 3774 8414 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 3710 8264 3774 8328 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 3710 8264 3774 8328 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 3710 8178 3774 8242 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 3710 8178 3774 8242 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 3710 8092 3774 8156 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 3710 8092 3774 8156 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 3710 8006 3774 8070 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 3710 8006 3774 8070 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 3710 7920 3774 7984 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 3710 7920 3774 7984 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 3630 8780 3694 8844 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 3630 8780 3694 8844 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 3630 8694 3694 8758 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 3630 8694 3694 8758 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 3630 8608 3694 8672 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 3630 8608 3694 8672 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 3630 8522 3694 8586 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 3630 8522 3694 8586 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 3630 8436 3694 8500 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 3630 8436 3694 8500 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 3630 8350 3694 8414 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 3630 8350 3694 8414 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 3630 8264 3694 8328 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 3630 8264 3694 8328 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 3630 8178 3694 8242 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 3630 8178 3694 8242 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 3630 8092 3694 8156 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 3630 8092 3694 8156 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 3630 8006 3694 8070 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 3630 8006 3694 8070 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 3630 7920 3694 7984 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 3630 7920 3694 7984 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 3550 8780 3614 8844 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 3550 8780 3614 8844 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 3550 8694 3614 8758 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 3550 8694 3614 8758 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 3550 8608 3614 8672 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 3550 8608 3614 8672 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 3550 8522 3614 8586 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 3550 8522 3614 8586 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 3550 8436 3614 8500 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 3550 8436 3614 8500 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 3550 8350 3614 8414 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 3550 8350 3614 8414 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 3550 8264 3614 8328 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 3550 8264 3614 8328 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 3550 8178 3614 8242 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 3550 8178 3614 8242 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 3550 8092 3614 8156 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 3550 8092 3614 8156 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 3550 8006 3614 8070 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 3550 8006 3614 8070 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 3550 7920 3614 7984 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 3550 7920 3614 7984 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 3470 8780 3534 8844 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 3470 8780 3534 8844 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 3470 8694 3534 8758 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 3470 8694 3534 8758 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 3470 8608 3534 8672 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 3470 8608 3534 8672 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 3470 8522 3534 8586 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 3470 8522 3534 8586 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 3470 8436 3534 8500 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 3470 8436 3534 8500 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 3470 8350 3534 8414 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 3470 8350 3534 8414 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 3470 8264 3534 8328 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 3470 8264 3534 8328 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 3470 8178 3534 8242 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 3470 8178 3534 8242 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 3470 8092 3534 8156 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 3470 8092 3534 8156 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 3470 8006 3534 8070 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 3470 8006 3534 8070 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 3470 7920 3534 7984 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 3470 7920 3534 7984 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 3390 8780 3454 8844 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 3390 8780 3454 8844 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 3390 8694 3454 8758 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 3390 8694 3454 8758 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 3390 8608 3454 8672 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 3390 8608 3454 8672 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 3390 8522 3454 8586 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 3390 8522 3454 8586 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 3390 8436 3454 8500 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 3390 8436 3454 8500 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 3390 8350 3454 8414 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 3390 8350 3454 8414 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 3390 8264 3454 8328 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 3390 8264 3454 8328 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 3390 8178 3454 8242 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 3390 8178 3454 8242 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 3390 8092 3454 8156 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 3390 8092 3454 8156 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 3390 8006 3454 8070 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 3390 8006 3454 8070 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 3390 7920 3454 7984 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 3390 7920 3454 7984 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 3310 8780 3374 8844 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 3310 8780 3374 8844 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 3310 8694 3374 8758 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 3310 8694 3374 8758 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 3310 8608 3374 8672 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 3310 8608 3374 8672 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 3310 8522 3374 8586 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 3310 8522 3374 8586 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 3310 8436 3374 8500 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 3310 8436 3374 8500 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 3310 8350 3374 8414 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 3310 8350 3374 8414 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 3310 8264 3374 8328 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 3310 8264 3374 8328 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 3310 8178 3374 8242 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 3310 8178 3374 8242 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 3310 8092 3374 8156 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 3310 8092 3374 8156 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 3310 8006 3374 8070 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 3310 8006 3374 8070 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 3310 7920 3374 7984 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 3310 7920 3374 7984 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 3230 8780 3294 8844 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 3230 8780 3294 8844 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 3230 8694 3294 8758 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 3230 8694 3294 8758 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 3230 8608 3294 8672 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 3230 8608 3294 8672 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 3230 8522 3294 8586 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 3230 8522 3294 8586 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 3230 8436 3294 8500 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 3230 8436 3294 8500 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 3230 8350 3294 8414 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 3230 8350 3294 8414 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 3230 8264 3294 8328 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 3230 8264 3294 8328 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 3230 8178 3294 8242 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 3230 8178 3294 8242 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 3230 8092 3294 8156 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 3230 8092 3294 8156 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 3230 8006 3294 8070 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 3230 8006 3294 8070 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 3230 7920 3294 7984 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 3230 7920 3294 7984 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 3150 8780 3214 8844 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 3150 8780 3214 8844 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 3150 8694 3214 8758 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 3150 8694 3214 8758 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 3150 8608 3214 8672 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 3150 8608 3214 8672 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 3150 8522 3214 8586 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 3150 8522 3214 8586 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 3150 8436 3214 8500 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 3150 8436 3214 8500 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 3150 8350 3214 8414 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 3150 8350 3214 8414 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 3150 8264 3214 8328 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 3150 8264 3214 8328 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 3150 8178 3214 8242 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 3150 8178 3214 8242 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 3150 8092 3214 8156 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 3150 8092 3214 8156 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 3150 8006 3214 8070 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 3150 8006 3214 8070 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 3150 7920 3214 7984 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 3150 7920 3214 7984 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 3070 8780 3134 8844 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 3070 8780 3134 8844 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 3070 8694 3134 8758 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 3070 8694 3134 8758 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 3070 8608 3134 8672 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 3070 8608 3134 8672 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 3070 8522 3134 8586 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 3070 8522 3134 8586 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 3070 8436 3134 8500 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 3070 8436 3134 8500 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 3070 8350 3134 8414 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 3070 8350 3134 8414 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 3070 8264 3134 8328 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 3070 8264 3134 8328 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 3070 8178 3134 8242 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 3070 8178 3134 8242 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 3070 8092 3134 8156 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 3070 8092 3134 8156 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 3070 8006 3134 8070 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 3070 8006 3134 8070 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 3070 7920 3134 7984 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 3070 7920 3134 7984 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2990 8780 3054 8844 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2990 8780 3054 8844 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2990 8694 3054 8758 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2990 8694 3054 8758 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2990 8608 3054 8672 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2990 8608 3054 8672 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2990 8522 3054 8586 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2990 8522 3054 8586 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2990 8436 3054 8500 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2990 8436 3054 8500 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2990 8350 3054 8414 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2990 8350 3054 8414 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2990 8264 3054 8328 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2990 8264 3054 8328 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2990 8178 3054 8242 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2990 8178 3054 8242 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2990 8092 3054 8156 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2990 8092 3054 8156 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2990 8006 3054 8070 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2990 8006 3054 8070 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2990 7920 3054 7984 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2990 7920 3054 7984 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2910 8780 2974 8844 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2910 8780 2974 8844 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2910 8694 2974 8758 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2910 8694 2974 8758 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2910 8608 2974 8672 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2910 8608 2974 8672 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2910 8522 2974 8586 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2910 8522 2974 8586 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2910 8436 2974 8500 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2910 8436 2974 8500 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2910 8350 2974 8414 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2910 8350 2974 8414 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2910 8264 2974 8328 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2910 8264 2974 8328 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2910 8178 2974 8242 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2910 8178 2974 8242 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2910 8092 2974 8156 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2910 8092 2974 8156 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2910 8006 2974 8070 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2910 8006 2974 8070 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2910 7920 2974 7984 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2910 7920 2974 7984 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2830 8780 2894 8844 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2830 8780 2894 8844 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2830 8694 2894 8758 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2830 8694 2894 8758 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2830 8608 2894 8672 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2830 8608 2894 8672 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2830 8522 2894 8586 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2830 8522 2894 8586 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2830 8436 2894 8500 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2830 8436 2894 8500 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2830 8350 2894 8414 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2830 8350 2894 8414 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2830 8264 2894 8328 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2830 8264 2894 8328 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2830 8178 2894 8242 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2830 8178 2894 8242 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2830 8092 2894 8156 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2830 8092 2894 8156 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2830 8006 2894 8070 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2830 8006 2894 8070 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2830 7920 2894 7984 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2830 7920 2894 7984 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2750 8780 2814 8844 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2750 8780 2814 8844 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2750 8694 2814 8758 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2750 8694 2814 8758 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2750 8608 2814 8672 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2750 8608 2814 8672 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2750 8522 2814 8586 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2750 8522 2814 8586 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2750 8436 2814 8500 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2750 8436 2814 8500 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2750 8350 2814 8414 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2750 8350 2814 8414 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2750 8264 2814 8328 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2750 8264 2814 8328 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2750 8178 2814 8242 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2750 8178 2814 8242 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2750 8092 2814 8156 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2750 8092 2814 8156 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2750 8006 2814 8070 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2750 8006 2814 8070 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2750 7920 2814 7984 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2750 7920 2814 7984 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2670 8780 2734 8844 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2670 8780 2734 8844 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2670 8694 2734 8758 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2670 8694 2734 8758 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2670 8608 2734 8672 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2670 8608 2734 8672 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2670 8522 2734 8586 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2670 8522 2734 8586 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2670 8436 2734 8500 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2670 8436 2734 8500 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2670 8350 2734 8414 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2670 8350 2734 8414 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2670 8264 2734 8328 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2670 8264 2734 8328 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2670 8178 2734 8242 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2670 8178 2734 8242 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2670 8092 2734 8156 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2670 8092 2734 8156 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2670 8006 2734 8070 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2670 8006 2734 8070 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2670 7920 2734 7984 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2670 7920 2734 7984 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2590 8780 2654 8844 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2590 8780 2654 8844 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2590 8694 2654 8758 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2590 8694 2654 8758 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2590 8608 2654 8672 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2590 8608 2654 8672 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2590 8522 2654 8586 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2590 8522 2654 8586 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2590 8436 2654 8500 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2590 8436 2654 8500 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2590 8350 2654 8414 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2590 8350 2654 8414 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2590 8264 2654 8328 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2590 8264 2654 8328 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2590 8178 2654 8242 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2590 8178 2654 8242 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2590 8092 2654 8156 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2590 8092 2654 8156 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2590 8006 2654 8070 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2590 8006 2654 8070 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2590 7920 2654 7984 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2590 7920 2654 7984 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2510 8780 2574 8844 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2510 8780 2574 8844 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2510 8694 2574 8758 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2510 8694 2574 8758 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2510 8608 2574 8672 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2510 8608 2574 8672 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2510 8522 2574 8586 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2510 8522 2574 8586 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2510 8436 2574 8500 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2510 8436 2574 8500 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2510 8350 2574 8414 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2510 8350 2574 8414 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2510 8264 2574 8328 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2510 8264 2574 8328 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2510 8178 2574 8242 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2510 8178 2574 8242 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2510 8092 2574 8156 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2510 8092 2574 8156 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2510 8006 2574 8070 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2510 8006 2574 8070 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2510 7920 2574 7984 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2510 7920 2574 7984 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2430 8780 2494 8844 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2430 8780 2494 8844 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2430 8694 2494 8758 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2430 8694 2494 8758 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2430 8608 2494 8672 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2430 8608 2494 8672 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2430 8522 2494 8586 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2430 8522 2494 8586 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2430 8436 2494 8500 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2430 8436 2494 8500 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2430 8350 2494 8414 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2430 8350 2494 8414 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2430 8264 2494 8328 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2430 8264 2494 8328 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2430 8178 2494 8242 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2430 8178 2494 8242 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2430 8092 2494 8156 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2430 8092 2494 8156 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2430 8006 2494 8070 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2430 8006 2494 8070 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2430 7920 2494 7984 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2430 7920 2494 7984 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2350 8780 2414 8844 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2350 8780 2414 8844 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2350 8694 2414 8758 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2350 8694 2414 8758 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2350 8608 2414 8672 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2350 8608 2414 8672 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2350 8522 2414 8586 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2350 8522 2414 8586 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2350 8436 2414 8500 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2350 8436 2414 8500 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2350 8350 2414 8414 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2350 8350 2414 8414 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2350 8264 2414 8328 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2350 8264 2414 8328 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2350 8178 2414 8242 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2350 8178 2414 8242 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2350 8092 2414 8156 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2350 8092 2414 8156 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2350 8006 2414 8070 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2350 8006 2414 8070 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2350 7920 2414 7984 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2350 7920 2414 7984 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2270 8780 2334 8844 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2270 8780 2334 8844 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2270 8694 2334 8758 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2270 8694 2334 8758 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2270 8608 2334 8672 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2270 8608 2334 8672 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2270 8522 2334 8586 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2270 8522 2334 8586 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2270 8436 2334 8500 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2270 8436 2334 8500 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2270 8350 2334 8414 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2270 8350 2334 8414 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2270 8264 2334 8328 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2270 8264 2334 8328 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2270 8178 2334 8242 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2270 8178 2334 8242 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2270 8092 2334 8156 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2270 8092 2334 8156 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2270 8006 2334 8070 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2270 8006 2334 8070 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2270 7920 2334 7984 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2270 7920 2334 7984 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2190 8780 2254 8844 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2190 8780 2254 8844 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2190 8694 2254 8758 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2190 8694 2254 8758 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2190 8608 2254 8672 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2190 8608 2254 8672 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2190 8522 2254 8586 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2190 8522 2254 8586 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2190 8436 2254 8500 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2190 8436 2254 8500 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2190 8350 2254 8414 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2190 8350 2254 8414 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2190 8264 2254 8328 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2190 8264 2254 8328 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2190 8178 2254 8242 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2190 8178 2254 8242 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2190 8092 2254 8156 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2190 8092 2254 8156 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2190 8006 2254 8070 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2190 8006 2254 8070 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2190 7920 2254 7984 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2190 7920 2254 7984 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2110 8780 2174 8844 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2110 8780 2174 8844 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2110 8694 2174 8758 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2110 8694 2174 8758 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2110 8608 2174 8672 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2110 8608 2174 8672 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2110 8522 2174 8586 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2110 8522 2174 8586 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2110 8436 2174 8500 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2110 8436 2174 8500 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2110 8350 2174 8414 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2110 8350 2174 8414 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2110 8264 2174 8328 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2110 8264 2174 8328 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2110 8178 2174 8242 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2110 8178 2174 8242 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2110 8092 2174 8156 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2110 8092 2174 8156 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2110 8006 2174 8070 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2110 8006 2174 8070 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2110 7920 2174 7984 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2110 7920 2174 7984 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2030 8780 2094 8844 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2030 8780 2094 8844 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2030 8694 2094 8758 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2030 8694 2094 8758 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2030 8608 2094 8672 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2030 8608 2094 8672 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2030 8522 2094 8586 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2030 8522 2094 8586 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2030 8436 2094 8500 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2030 8436 2094 8500 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2030 8350 2094 8414 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2030 8350 2094 8414 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2030 8264 2094 8328 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2030 8264 2094 8328 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2030 8178 2094 8242 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2030 8178 2094 8242 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2030 8092 2094 8156 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2030 8092 2094 8156 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2030 8006 2094 8070 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2030 8006 2094 8070 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 2030 7920 2094 7984 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 2030 7920 2094 7984 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1950 8780 2014 8844 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1950 8780 2014 8844 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1950 8694 2014 8758 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1950 8694 2014 8758 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1950 8608 2014 8672 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1950 8608 2014 8672 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1950 8522 2014 8586 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1950 8522 2014 8586 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1950 8436 2014 8500 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1950 8436 2014 8500 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1950 8350 2014 8414 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1950 8350 2014 8414 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1950 8264 2014 8328 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1950 8264 2014 8328 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1950 8178 2014 8242 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1950 8178 2014 8242 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1950 8092 2014 8156 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1950 8092 2014 8156 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1950 8006 2014 8070 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1950 8006 2014 8070 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1950 7920 2014 7984 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1950 7920 2014 7984 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1870 8780 1934 8844 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1870 8780 1934 8844 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1870 8694 1934 8758 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1870 8694 1934 8758 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1870 8608 1934 8672 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1870 8608 1934 8672 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1870 8522 1934 8586 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1870 8522 1934 8586 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1870 8436 1934 8500 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1870 8436 1934 8500 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1870 8350 1934 8414 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1870 8350 1934 8414 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1870 8264 1934 8328 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1870 8264 1934 8328 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1870 8178 1934 8242 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1870 8178 1934 8242 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1870 8092 1934 8156 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1870 8092 1934 8156 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1870 8006 1934 8070 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1870 8006 1934 8070 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1870 7920 1934 7984 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1870 7920 1934 7984 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1790 8780 1854 8844 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1790 8780 1854 8844 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1790 8694 1854 8758 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1790 8694 1854 8758 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1790 8608 1854 8672 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1790 8608 1854 8672 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1790 8522 1854 8586 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1790 8522 1854 8586 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1790 8436 1854 8500 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1790 8436 1854 8500 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1790 8350 1854 8414 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1790 8350 1854 8414 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1790 8264 1854 8328 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1790 8264 1854 8328 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1790 8178 1854 8242 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1790 8178 1854 8242 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1790 8092 1854 8156 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1790 8092 1854 8156 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1790 8006 1854 8070 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1790 8006 1854 8070 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1790 7920 1854 7984 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1790 7920 1854 7984 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1710 8780 1774 8844 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1710 8780 1774 8844 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1710 8694 1774 8758 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1710 8694 1774 8758 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1710 8608 1774 8672 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1710 8608 1774 8672 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1710 8522 1774 8586 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1710 8522 1774 8586 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1710 8436 1774 8500 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1710 8436 1774 8500 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1710 8350 1774 8414 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1710 8350 1774 8414 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1710 8264 1774 8328 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1710 8264 1774 8328 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1710 8178 1774 8242 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1710 8178 1774 8242 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1710 8092 1774 8156 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1710 8092 1774 8156 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1710 8006 1774 8070 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1710 8006 1774 8070 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1710 7920 1774 7984 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1710 7920 1774 7984 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1630 8780 1694 8844 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1630 8780 1694 8844 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1630 8694 1694 8758 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1630 8694 1694 8758 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1630 8608 1694 8672 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1630 8608 1694 8672 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1630 8522 1694 8586 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1630 8522 1694 8586 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1630 8436 1694 8500 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1630 8436 1694 8500 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1630 8350 1694 8414 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1630 8350 1694 8414 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1630 8264 1694 8328 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1630 8264 1694 8328 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1630 8178 1694 8242 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1630 8178 1694 8242 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1630 8092 1694 8156 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1630 8092 1694 8156 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1630 8006 1694 8070 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1630 8006 1694 8070 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1630 7920 1694 7984 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1630 7920 1694 7984 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1550 8780 1614 8844 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1550 8780 1614 8844 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1550 8694 1614 8758 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1550 8694 1614 8758 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1550 8608 1614 8672 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1550 8608 1614 8672 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1550 8522 1614 8586 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1550 8522 1614 8586 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1550 8436 1614 8500 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1550 8436 1614 8500 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1550 8350 1614 8414 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1550 8350 1614 8414 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1550 8264 1614 8328 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1550 8264 1614 8328 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1550 8178 1614 8242 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1550 8178 1614 8242 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1550 8092 1614 8156 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1550 8092 1614 8156 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1550 8006 1614 8070 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1550 8006 1614 8070 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1550 7920 1614 7984 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1550 7920 1614 7984 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1470 8780 1534 8844 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1470 8780 1534 8844 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1470 8694 1534 8758 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1470 8694 1534 8758 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1470 8608 1534 8672 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1470 8608 1534 8672 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1470 8522 1534 8586 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1470 8522 1534 8586 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1470 8436 1534 8500 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1470 8436 1534 8500 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1470 8350 1534 8414 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1470 8350 1534 8414 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1470 8264 1534 8328 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1470 8264 1534 8328 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1470 8178 1534 8242 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1470 8178 1534 8242 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1470 8092 1534 8156 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1470 8092 1534 8156 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1470 8006 1534 8070 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1470 8006 1534 8070 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1470 7920 1534 7984 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1470 7920 1534 7984 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1390 8780 1454 8844 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1390 8780 1454 8844 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1390 8694 1454 8758 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1390 8694 1454 8758 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1390 8608 1454 8672 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1390 8608 1454 8672 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1390 8522 1454 8586 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1390 8522 1454 8586 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1390 8436 1454 8500 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1390 8436 1454 8500 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1390 8350 1454 8414 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1390 8350 1454 8414 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1390 8264 1454 8328 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1390 8264 1454 8328 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1390 8178 1454 8242 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1390 8178 1454 8242 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1390 8092 1454 8156 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1390 8092 1454 8156 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1390 8006 1454 8070 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1390 8006 1454 8070 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1390 7920 1454 7984 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1390 7920 1454 7984 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1310 8780 1374 8844 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1310 8780 1374 8844 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1310 8694 1374 8758 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1310 8694 1374 8758 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1310 8608 1374 8672 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1310 8608 1374 8672 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1310 8522 1374 8586 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1310 8522 1374 8586 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1310 8436 1374 8500 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1310 8436 1374 8500 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1310 8350 1374 8414 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1310 8350 1374 8414 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1310 8264 1374 8328 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1310 8264 1374 8328 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1310 8178 1374 8242 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1310 8178 1374 8242 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1310 8092 1374 8156 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1310 8092 1374 8156 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1310 8006 1374 8070 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1310 8006 1374 8070 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1310 7920 1374 7984 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1310 7920 1374 7984 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1230 8780 1294 8844 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1230 8780 1294 8844 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1230 8694 1294 8758 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1230 8694 1294 8758 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1230 8608 1294 8672 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1230 8608 1294 8672 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1230 8522 1294 8586 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1230 8522 1294 8586 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1230 8436 1294 8500 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1230 8436 1294 8500 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1230 8350 1294 8414 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1230 8350 1294 8414 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1230 8264 1294 8328 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1230 8264 1294 8328 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1230 8178 1294 8242 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1230 8178 1294 8242 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1230 8092 1294 8156 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1230 8092 1294 8156 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1230 8006 1294 8070 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1230 8006 1294 8070 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1230 7920 1294 7984 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1230 7920 1294 7984 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1150 8780 1214 8844 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1150 8780 1214 8844 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1150 8694 1214 8758 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1150 8694 1214 8758 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1150 8608 1214 8672 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1150 8608 1214 8672 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1150 8522 1214 8586 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1150 8522 1214 8586 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1150 8436 1214 8500 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1150 8436 1214 8500 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1150 8350 1214 8414 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1150 8350 1214 8414 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1150 8264 1214 8328 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1150 8264 1214 8328 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1150 8178 1214 8242 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1150 8178 1214 8242 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1150 8092 1214 8156 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1150 8092 1214 8156 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1150 8006 1214 8070 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1150 8006 1214 8070 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1150 7920 1214 7984 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1150 7920 1214 7984 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1070 8780 1134 8844 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1070 8780 1134 8844 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1070 8694 1134 8758 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1070 8694 1134 8758 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1070 8608 1134 8672 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1070 8608 1134 8672 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1070 8522 1134 8586 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1070 8522 1134 8586 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1070 8436 1134 8500 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1070 8436 1134 8500 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1070 8350 1134 8414 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1070 8350 1134 8414 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1070 8264 1134 8328 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1070 8264 1134 8328 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1070 8178 1134 8242 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1070 8178 1134 8242 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1070 8092 1134 8156 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1070 8092 1134 8156 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1070 8006 1134 8070 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1070 8006 1134 8070 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 1070 7920 1134 7984 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 1070 7920 1134 7984 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 990 8780 1054 8844 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 990 8780 1054 8844 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 990 8694 1054 8758 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 990 8694 1054 8758 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 990 8608 1054 8672 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 990 8608 1054 8672 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 990 8522 1054 8586 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 990 8522 1054 8586 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 990 8436 1054 8500 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 990 8436 1054 8500 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 990 8350 1054 8414 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 990 8350 1054 8414 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 990 8264 1054 8328 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 990 8264 1054 8328 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 990 8178 1054 8242 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 990 8178 1054 8242 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 990 8092 1054 8156 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 990 8092 1054 8156 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 990 8006 1054 8070 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 990 8006 1054 8070 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 990 7920 1054 7984 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 990 7920 1054 7984 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 910 8780 974 8844 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 910 8780 974 8844 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 910 8694 974 8758 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 910 8694 974 8758 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 910 8608 974 8672 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 910 8608 974 8672 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 910 8522 974 8586 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 910 8522 974 8586 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 910 8436 974 8500 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 910 8436 974 8500 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 910 8350 974 8414 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 910 8350 974 8414 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 910 8264 974 8328 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 910 8264 974 8328 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 910 8178 974 8242 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 910 8178 974 8242 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 910 8092 974 8156 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 910 8092 974 8156 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 910 8006 974 8070 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 910 8006 974 8070 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 910 7920 974 7984 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 910 7920 974 7984 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 830 8780 894 8844 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 830 8780 894 8844 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 830 8694 894 8758 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 830 8694 894 8758 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 830 8608 894 8672 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 830 8608 894 8672 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 830 8522 894 8586 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 830 8522 894 8586 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 830 8436 894 8500 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 830 8436 894 8500 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 830 8350 894 8414 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 830 8350 894 8414 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 830 8264 894 8328 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 830 8264 894 8328 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 830 8178 894 8242 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 830 8178 894 8242 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 830 8092 894 8156 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 830 8092 894 8156 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 830 8006 894 8070 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 830 8006 894 8070 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 830 7920 894 7984 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 830 7920 894 7984 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 750 8780 814 8844 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 750 8780 814 8844 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 750 8694 814 8758 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 750 8694 814 8758 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 750 8608 814 8672 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 750 8608 814 8672 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 750 8522 814 8586 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 750 8522 814 8586 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 750 8436 814 8500 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 750 8436 814 8500 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 750 8350 814 8414 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 750 8350 814 8414 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 750 8264 814 8328 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 750 8264 814 8328 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 750 8178 814 8242 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 750 8178 814 8242 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 750 8092 814 8156 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 750 8092 814 8156 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 750 8006 814 8070 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 750 8006 814 8070 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 750 7920 814 7984 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 750 7920 814 7984 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 670 8780 734 8844 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 670 8780 734 8844 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 670 8694 734 8758 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 670 8694 734 8758 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 670 8608 734 8672 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 670 8608 734 8672 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 670 8522 734 8586 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 670 8522 734 8586 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 670 8436 734 8500 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 670 8436 734 8500 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 670 8350 734 8414 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 670 8350 734 8414 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 670 8264 734 8328 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 670 8264 734 8328 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 670 8178 734 8242 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 670 8178 734 8242 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 670 8092 734 8156 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 670 8092 734 8156 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 670 8006 734 8070 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 670 8006 734 8070 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 670 7920 734 7984 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 670 7920 734 7984 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 590 8780 654 8844 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 590 8780 654 8844 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 590 8694 654 8758 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 590 8694 654 8758 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 590 8608 654 8672 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 590 8608 654 8672 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 590 8522 654 8586 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 590 8522 654 8586 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 590 8436 654 8500 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 590 8436 654 8500 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 590 8350 654 8414 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 590 8350 654 8414 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 590 8264 654 8328 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 590 8264 654 8328 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 590 8178 654 8242 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 590 8178 654 8242 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 590 8092 654 8156 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 590 8092 654 8156 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 590 8006 654 8070 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 590 8006 654 8070 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 590 7920 654 7984 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 590 7920 654 7984 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 510 8780 574 8844 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 510 8780 574 8844 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 510 8694 574 8758 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 510 8694 574 8758 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 510 8608 574 8672 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 510 8608 574 8672 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 510 8522 574 8586 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 510 8522 574 8586 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 510 8436 574 8500 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 510 8436 574 8500 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 510 8350 574 8414 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 510 8350 574 8414 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 510 8264 574 8328 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 510 8264 574 8328 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 510 8178 574 8242 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 510 8178 574 8242 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 510 8092 574 8156 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 510 8092 574 8156 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 510 8006 574 8070 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 510 8006 574 8070 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 510 7920 574 7984 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 510 7920 574 7984 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 430 8780 494 8844 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 430 8780 494 8844 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 430 8694 494 8758 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 430 8694 494 8758 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 430 8608 494 8672 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 430 8608 494 8672 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 430 8522 494 8586 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 430 8522 494 8586 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 430 8436 494 8500 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 430 8436 494 8500 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 430 8350 494 8414 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 430 8350 494 8414 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 430 8264 494 8328 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 430 8264 494 8328 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 430 8178 494 8242 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 430 8178 494 8242 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 430 8092 494 8156 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 430 8092 494 8156 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 430 8006 494 8070 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 430 8006 494 8070 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 430 7920 494 7984 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 430 7920 494 7984 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 349 8780 413 8844 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 349 8780 413 8844 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 349 8694 413 8758 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 349 8694 413 8758 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 349 8608 413 8672 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 349 8608 413 8672 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 349 8522 413 8586 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 349 8522 413 8586 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 349 8436 413 8500 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 349 8436 413 8500 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 349 8350 413 8414 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 349 8350 413 8414 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 349 8264 413 8328 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 349 8264 413 8328 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 349 8178 413 8242 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 349 8178 413 8242 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 349 8092 413 8156 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 349 8092 413 8156 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 349 8006 413 8070 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 349 8006 413 8070 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 349 7920 413 7984 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 349 7920 413 7984 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 268 8780 332 8844 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 268 8780 332 8844 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 268 8694 332 8758 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 268 8694 332 8758 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 268 8608 332 8672 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 268 8608 332 8672 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 268 8522 332 8586 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 268 8522 332 8586 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 268 8436 332 8500 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 268 8436 332 8500 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 268 8350 332 8414 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 268 8350 332 8414 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 268 8264 332 8328 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 268 8264 332 8328 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 268 8178 332 8242 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 268 8178 332 8242 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 268 8092 332 8156 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 268 8092 332 8156 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 268 8006 332 8070 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 268 8006 332 8070 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 268 7920 332 7984 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 268 7920 332 7984 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 187 8780 251 8844 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 187 8694 251 8758 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 187 8608 251 8672 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 187 8522 251 8586 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 187 8436 251 8500 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 187 8350 251 8414 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 187 8264 251 8328 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 187 8178 251 8242 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 187 8092 251 8156 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 187 8006 251 8070 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 187 7920 251 7984 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 106 8780 170 8844 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 106 8694 170 8758 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 106 8608 170 8672 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 106 8522 170 8586 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 106 8436 170 8500 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 106 8350 170 8414 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 106 8264 170 8328 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 106 8178 170 8242 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 106 8092 170 8156 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 106 8006 170 8070 6 VSSD
port 4 nsew ground bidirectional
rlabel metal3 s 106 7920 170 7984 6 VSSD
port 4 nsew ground bidirectional
rlabel metal5 s 0 4787 254 5677 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal5 s 14746 4787 15000 5677 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal5 s 14746 34757 15000 39600 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal5 s 0 34757 254 39600 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 0 4767 254 5697 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 14746 4767 15000 5697 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 14746 34757 15000 39600 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 0 34757 254 39600 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal5 s 0 5997 254 6647 6 VSWITCH
port 6 nsew power bidirectional
rlabel metal5 s 14746 5997 15000 6647 6 VSWITCH
port 6 nsew power bidirectional
rlabel metal4 s 0 5977 254 6667 6 VSWITCH
port 6 nsew power bidirectional
rlabel metal4 s 14746 5977 15000 6667 6 VSWITCH
port 6 nsew power bidirectional
rlabel metal5 s 0 11267 254 12117 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal5 s 14746 11267 15000 12117 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 0 11247 254 12137 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 14746 11247 15000 12137 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal5 s 0 2607 193 3257 6 VDDA
port 8 nsew power bidirectional
rlabel metal5 s 14807 2607 15000 3257 6 VDDA
port 8 nsew power bidirectional
rlabel metal4 s 0 2587 193 3277 6 VDDA
port 8 nsew power bidirectional
rlabel metal4 s 14807 2587 15000 3277 6 VDDA
port 8 nsew power bidirectional
rlabel metal5 s 0 1397 254 2287 6 VCCD
port 9 nsew power bidirectional
rlabel metal5 s 14746 1397 15000 2287 6 VCCD
port 9 nsew power bidirectional
rlabel metal4 s 0 1377 254 2307 6 VCCD
port 9 nsew power bidirectional
rlabel metal4 s 14746 1377 15000 2307 6 VCCD
port 9 nsew power bidirectional
rlabel metal5 s 0 27 254 1077 6 VCCHIB
port 10 nsew power bidirectional
rlabel metal5 s 14746 27 15000 1077 6 VCCHIB
port 10 nsew power bidirectional
rlabel metal4 s 0 7 254 1097 6 VCCHIB
port 10 nsew power bidirectional
rlabel metal4 s 14746 7 15000 1097 6 VCCHIB
port 10 nsew power bidirectional
rlabel metal4 s 0 9273 15000 9869 6 AMUXBUS_B
port 11 nsew signal bidirectional
rlabel metal4 s 0 10225 15000 10821 6 AMUXBUS_A
port 12 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 15000 39600
string LEFclass PAD
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_END 2266656
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 2174144
<< end >>
