magic
tech sky130B
magscale 1 2
timestamp 1649977179
<< nwell >>
rect -38 261 1694 582
<< pwell >>
rect 1 21 1655 203
rect 30 -17 64 21
<< locali >>
rect 19 451 757 485
rect 19 97 64 451
rect 1152 285 1570 319
rect 112 221 248 265
rect 112 199 214 221
rect 391 199 710 265
rect 1152 258 1186 285
rect 769 215 1186 258
rect 19 63 757 97
rect 1536 199 1570 285
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1656 561
rect 795 451 861 527
rect 963 451 1029 527
rect 1131 451 1197 527
rect 1231 417 1265 493
rect 1299 451 1365 527
rect 1399 417 1433 493
rect 1487 451 1553 527
rect 439 383 1433 417
rect 1231 359 1265 383
rect 1399 359 1433 383
rect 1587 359 1639 493
rect 103 315 1116 349
rect 1346 215 1502 249
rect 271 165 340 187
rect 1230 181 1290 187
rect 103 131 340 165
rect 439 131 1097 165
rect 795 17 861 93
rect 895 51 929 131
rect 963 17 1029 93
rect 1063 51 1097 131
rect 1230 143 1433 181
rect 1131 17 1196 118
rect 1230 51 1265 143
rect 1309 17 1359 109
rect 1399 102 1433 143
rect 1468 165 1502 215
rect 1604 165 1639 359
rect 1468 131 1639 165
rect 1487 17 1553 93
rect 1587 51 1639 131
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1656 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 1593 527 1627 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1593 -17 1627 17
<< metal1 >>
rect 0 561 1656 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1656 561
rect 0 496 1656 527
rect 0 17 1656 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1656 17
rect 0 -48 1656 -17
<< obsm1 >>
rect 294 184 352 193
rect 1218 184 1276 193
rect 294 156 1276 184
rect 294 147 352 156
rect 1218 147 1276 156
<< labels >>
rlabel locali s 112 199 214 221 6 A0
port 1 nsew signal input
rlabel locali s 112 221 248 265 6 A0
port 1 nsew signal input
rlabel locali s 391 199 710 265 6 A1
port 2 nsew signal input
rlabel locali s 1536 199 1570 285 6 S
port 3 nsew signal input
rlabel locali s 769 215 1186 258 6 S
port 3 nsew signal input
rlabel locali s 1152 258 1186 285 6 S
port 3 nsew signal input
rlabel locali s 1152 285 1570 319 6 S
port 3 nsew signal input
rlabel metal1 s 0 -48 1656 48 8 VGND
port 4 nsew ground bidirectional abutment
rlabel pwell s 30 -17 64 21 6 VNB
port 5 nsew ground bidirectional
rlabel pwell s 1 21 1655 203 6 VNB
port 5 nsew ground bidirectional
rlabel nwell s -38 261 1694 582 6 VPB
port 6 nsew power bidirectional
rlabel metal1 s 0 496 1656 592 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 19 63 757 97 6 Y
port 8 nsew signal output
rlabel locali s 19 97 64 451 6 Y
port 8 nsew signal output
rlabel locali s 19 451 757 485 6 Y
port 8 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 1656 544
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_END 1743856
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 1731714
<< end >>
