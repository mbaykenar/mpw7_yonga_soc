magic
tech sky130A
magscale 1 2
timestamp 1649977179
<< nwell >>
rect -38 261 1694 582
<< pwell >>
rect 834 157 1655 203
rect 1 21 1655 157
rect 30 -17 64 21
<< scnmos >>
rect 79 47 109 131
rect 163 47 193 131
rect 351 47 381 131
rect 435 47 465 131
rect 543 47 573 119
rect 629 47 659 119
rect 724 47 754 131
rect 912 47 942 177
rect 998 47 1028 177
rect 1092 47 1122 177
rect 1180 47 1210 177
rect 1368 47 1398 131
rect 1463 47 1493 177
rect 1547 47 1577 177
<< scpmoshvt >>
rect 79 363 109 491
rect 163 363 193 491
rect 351 369 381 497
rect 435 369 465 497
rect 531 413 561 497
rect 615 413 645 497
rect 711 413 741 497
rect 912 297 942 497
rect 998 297 1028 497
rect 1092 297 1122 497
rect 1180 297 1210 497
rect 1368 369 1398 497
rect 1463 297 1493 497
rect 1547 297 1577 497
<< ndiff >>
rect 27 119 79 131
rect 27 85 35 119
rect 69 85 79 119
rect 27 47 79 85
rect 109 93 163 131
rect 109 59 119 93
rect 153 59 163 93
rect 109 47 163 59
rect 193 119 245 131
rect 193 85 203 119
rect 237 85 245 119
rect 193 47 245 85
rect 299 119 351 131
rect 299 85 307 119
rect 341 85 351 119
rect 299 47 351 85
rect 381 89 435 131
rect 381 55 391 89
rect 425 55 435 89
rect 381 47 435 55
rect 465 119 515 131
rect 860 133 912 177
rect 674 119 724 131
rect 465 47 543 119
rect 573 107 629 119
rect 573 73 584 107
rect 618 73 629 107
rect 573 47 629 73
rect 659 47 724 119
rect 754 106 806 131
rect 754 72 764 106
rect 798 72 806 106
rect 754 47 806 72
rect 860 99 868 133
rect 902 99 912 133
rect 860 47 912 99
rect 942 47 998 177
rect 1028 89 1092 177
rect 1028 55 1038 89
rect 1072 55 1092 89
rect 1028 47 1092 55
rect 1122 133 1180 177
rect 1122 99 1136 133
rect 1170 99 1180 133
rect 1122 47 1180 99
rect 1210 93 1262 177
rect 1413 131 1463 177
rect 1210 59 1220 93
rect 1254 59 1262 93
rect 1210 47 1262 59
rect 1316 119 1368 131
rect 1316 85 1324 119
rect 1358 85 1368 119
rect 1316 47 1368 85
rect 1398 93 1463 131
rect 1398 59 1418 93
rect 1452 59 1463 93
rect 1398 47 1463 59
rect 1493 129 1547 177
rect 1493 95 1503 129
rect 1537 95 1547 129
rect 1493 47 1547 95
rect 1577 161 1629 177
rect 1577 127 1587 161
rect 1621 127 1629 161
rect 1577 93 1629 127
rect 1577 59 1587 93
rect 1621 59 1629 93
rect 1577 47 1629 59
<< pdiff >>
rect 27 477 79 491
rect 27 443 35 477
rect 69 443 79 477
rect 27 409 79 443
rect 27 375 35 409
rect 69 375 79 409
rect 27 363 79 375
rect 109 461 163 491
rect 109 427 119 461
rect 153 427 163 461
rect 109 363 163 427
rect 193 477 245 491
rect 193 443 203 477
rect 237 443 245 477
rect 193 409 245 443
rect 193 375 203 409
rect 237 375 245 409
rect 193 363 245 375
rect 299 483 351 497
rect 299 449 307 483
rect 341 449 351 483
rect 299 415 351 449
rect 299 381 307 415
rect 341 381 351 415
rect 299 369 351 381
rect 381 485 435 497
rect 381 451 391 485
rect 425 451 435 485
rect 381 417 435 451
rect 381 383 391 417
rect 425 383 435 417
rect 381 369 435 383
rect 465 413 531 497
rect 561 485 615 497
rect 561 451 571 485
rect 605 451 615 485
rect 561 413 615 451
rect 645 413 711 497
rect 741 477 793 497
rect 741 443 751 477
rect 785 443 793 477
rect 741 413 793 443
rect 860 485 912 497
rect 860 451 868 485
rect 902 451 912 485
rect 465 369 515 413
rect 860 297 912 451
rect 942 471 998 497
rect 942 437 954 471
rect 988 437 998 471
rect 942 368 998 437
rect 942 334 954 368
rect 988 334 998 368
rect 942 297 998 334
rect 1028 489 1092 497
rect 1028 455 1038 489
rect 1072 455 1092 489
rect 1028 421 1092 455
rect 1028 387 1038 421
rect 1072 387 1092 421
rect 1028 297 1092 387
rect 1122 477 1180 497
rect 1122 443 1136 477
rect 1170 443 1180 477
rect 1122 409 1180 443
rect 1122 375 1136 409
rect 1170 375 1180 409
rect 1122 297 1180 375
rect 1210 485 1262 497
rect 1210 451 1220 485
rect 1254 451 1262 485
rect 1210 417 1262 451
rect 1210 383 1220 417
rect 1254 383 1262 417
rect 1210 297 1262 383
rect 1316 485 1368 497
rect 1316 451 1324 485
rect 1358 451 1368 485
rect 1316 417 1368 451
rect 1316 383 1324 417
rect 1358 383 1368 417
rect 1316 369 1368 383
rect 1398 485 1463 497
rect 1398 451 1418 485
rect 1452 451 1463 485
rect 1398 417 1463 451
rect 1398 383 1418 417
rect 1452 383 1463 417
rect 1398 369 1463 383
rect 1413 297 1463 369
rect 1493 449 1547 497
rect 1493 415 1503 449
rect 1537 415 1547 449
rect 1493 381 1547 415
rect 1493 347 1503 381
rect 1537 347 1547 381
rect 1493 297 1547 347
rect 1577 485 1629 497
rect 1577 451 1587 485
rect 1621 451 1629 485
rect 1577 417 1629 451
rect 1577 383 1587 417
rect 1621 383 1629 417
rect 1577 349 1629 383
rect 1577 315 1587 349
rect 1621 315 1629 349
rect 1577 297 1629 315
<< ndiffc >>
rect 35 85 69 119
rect 119 59 153 93
rect 203 85 237 119
rect 307 85 341 119
rect 391 55 425 89
rect 584 73 618 107
rect 764 72 798 106
rect 868 99 902 133
rect 1038 55 1072 89
rect 1136 99 1170 133
rect 1220 59 1254 93
rect 1324 85 1358 119
rect 1418 59 1452 93
rect 1503 95 1537 129
rect 1587 127 1621 161
rect 1587 59 1621 93
<< pdiffc >>
rect 35 443 69 477
rect 35 375 69 409
rect 119 427 153 461
rect 203 443 237 477
rect 203 375 237 409
rect 307 449 341 483
rect 307 381 341 415
rect 391 451 425 485
rect 391 383 425 417
rect 571 451 605 485
rect 751 443 785 477
rect 868 451 902 485
rect 954 437 988 471
rect 954 334 988 368
rect 1038 455 1072 489
rect 1038 387 1072 421
rect 1136 443 1170 477
rect 1136 375 1170 409
rect 1220 451 1254 485
rect 1220 383 1254 417
rect 1324 451 1358 485
rect 1324 383 1358 417
rect 1418 451 1452 485
rect 1418 383 1452 417
rect 1503 415 1537 449
rect 1503 347 1537 381
rect 1587 451 1621 485
rect 1587 383 1621 417
rect 1587 315 1621 349
<< poly >>
rect 79 491 109 517
rect 163 491 193 517
rect 351 497 381 523
rect 435 497 465 523
rect 531 497 561 523
rect 615 497 645 523
rect 711 497 741 523
rect 912 497 942 523
rect 998 497 1028 523
rect 1092 497 1122 523
rect 1180 497 1210 523
rect 1368 497 1398 523
rect 1463 497 1493 523
rect 1547 497 1577 523
rect 79 348 109 363
rect 46 318 109 348
rect 46 280 76 318
rect 21 264 76 280
rect 163 274 193 363
rect 21 230 32 264
rect 66 230 76 264
rect 21 214 76 230
rect 118 264 193 274
rect 118 230 134 264
rect 168 230 193 264
rect 351 241 381 369
rect 118 220 193 230
rect 46 176 76 214
rect 46 146 109 176
rect 79 131 109 146
rect 163 131 193 220
rect 298 225 381 241
rect 298 191 308 225
rect 342 191 381 225
rect 435 219 465 369
rect 531 337 561 413
rect 615 375 645 413
rect 507 321 561 337
rect 603 365 669 375
rect 603 331 619 365
rect 653 331 669 365
rect 603 321 669 331
rect 711 373 741 413
rect 711 357 812 373
rect 711 323 768 357
rect 802 323 812 357
rect 507 287 517 321
rect 551 287 561 321
rect 711 307 812 323
rect 507 279 561 287
rect 507 271 659 279
rect 531 249 659 271
rect 298 175 381 191
rect 351 131 381 175
rect 424 203 478 219
rect 424 169 434 203
rect 468 169 478 203
rect 424 153 478 169
rect 533 191 587 207
rect 533 157 543 191
rect 577 157 587 191
rect 435 131 465 153
rect 533 141 587 157
rect 543 119 573 141
rect 629 119 659 249
rect 724 131 754 307
rect 912 265 942 297
rect 998 265 1028 297
rect 1092 265 1122 297
rect 1180 265 1210 297
rect 1368 265 1398 369
rect 1463 265 1493 297
rect 796 249 942 265
rect 796 215 806 249
rect 840 215 942 249
rect 796 199 942 215
rect 984 249 1038 265
rect 984 215 994 249
rect 1028 215 1038 249
rect 984 199 1038 215
rect 1080 249 1398 265
rect 1080 215 1090 249
rect 1124 215 1398 249
rect 1080 199 1398 215
rect 1441 259 1493 265
rect 1547 259 1577 297
rect 1441 249 1577 259
rect 1441 215 1451 249
rect 1485 215 1577 249
rect 1441 205 1577 215
rect 1441 199 1493 205
rect 912 177 942 199
rect 998 177 1028 199
rect 1092 177 1122 199
rect 1180 177 1210 199
rect 1368 131 1398 199
rect 1463 177 1493 199
rect 1547 177 1577 205
rect 79 21 109 47
rect 163 21 193 47
rect 351 21 381 47
rect 435 21 465 47
rect 543 21 573 47
rect 629 21 659 47
rect 724 21 754 47
rect 912 21 942 47
rect 998 21 1028 47
rect 1092 21 1122 47
rect 1180 21 1210 47
rect 1368 21 1398 47
rect 1463 21 1493 47
rect 1547 21 1577 47
<< polycont >>
rect 32 230 66 264
rect 134 230 168 264
rect 308 191 342 225
rect 619 331 653 365
rect 768 323 802 357
rect 517 287 551 321
rect 434 169 468 203
rect 543 157 577 191
rect 806 215 840 249
rect 994 215 1028 249
rect 1090 215 1124 249
rect 1451 215 1485 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1656 561
rect 17 477 69 493
rect 17 443 35 477
rect 17 409 69 443
rect 103 461 169 527
rect 103 427 119 461
rect 153 427 169 461
rect 203 477 248 493
rect 391 485 454 527
rect 751 485 920 527
rect 1022 489 1098 527
rect 237 443 248 477
rect 17 375 35 409
rect 203 409 248 443
rect 69 375 156 393
rect 17 359 156 375
rect 17 264 66 325
rect 17 230 32 264
rect 17 197 66 230
rect 122 323 156 359
rect 122 280 156 289
rect 237 391 248 409
rect 203 357 214 375
rect 203 337 248 357
rect 291 449 307 483
rect 341 449 357 483
rect 291 415 357 449
rect 291 381 307 415
rect 341 381 357 415
rect 122 264 168 280
rect 122 230 134 264
rect 122 214 168 230
rect 122 161 156 214
rect 17 127 156 161
rect 17 119 69 127
rect 17 85 35 119
rect 203 119 237 337
rect 291 333 357 381
rect 425 451 454 485
rect 549 451 571 485
rect 605 451 717 485
rect 391 417 454 451
rect 654 425 717 451
rect 751 477 868 485
rect 785 451 868 477
rect 902 451 920 485
rect 785 443 920 451
rect 751 427 920 443
rect 954 471 988 487
rect 425 383 454 417
rect 661 415 717 425
rect 679 409 717 415
rect 679 403 721 409
rect 391 367 454 383
rect 585 391 625 399
rect 683 398 721 403
rect 684 395 721 398
rect 686 392 721 395
rect 585 357 586 391
rect 620 381 625 391
rect 620 365 653 381
rect 291 299 428 333
rect 292 225 358 265
rect 292 191 308 225
rect 342 191 358 225
rect 394 219 428 299
rect 494 323 551 337
rect 528 321 551 323
rect 494 287 517 289
rect 494 271 551 287
rect 585 331 619 357
rect 585 315 653 331
rect 394 203 468 219
rect 585 207 619 315
rect 687 265 721 392
rect 954 373 988 437
rect 1022 455 1038 489
rect 1072 455 1098 489
rect 1022 421 1098 455
rect 1022 387 1038 421
rect 1072 387 1098 421
rect 1022 375 1098 387
rect 1136 477 1186 493
rect 1170 443 1186 477
rect 1136 409 1186 443
rect 1170 375 1186 409
rect 768 368 988 373
rect 768 357 954 368
rect 802 334 954 357
rect 988 334 1102 341
rect 802 323 1102 334
rect 768 307 1102 323
rect 1064 265 1102 307
rect 1136 332 1186 375
rect 1220 485 1272 527
rect 1254 451 1272 485
rect 1220 417 1272 451
rect 1254 383 1272 417
rect 1220 366 1272 383
rect 1307 485 1374 493
rect 1307 451 1324 485
rect 1358 451 1374 485
rect 1307 417 1374 451
rect 1307 383 1324 417
rect 1358 383 1374 417
rect 1136 299 1213 332
rect 1158 265 1213 299
rect 1307 265 1374 383
rect 1409 485 1468 527
rect 1409 451 1418 485
rect 1452 451 1468 485
rect 1409 417 1468 451
rect 1409 383 1418 417
rect 1452 383 1468 417
rect 1409 367 1468 383
rect 1503 449 1553 493
rect 1537 415 1553 449
rect 1503 381 1553 415
rect 1537 347 1553 381
rect 1503 321 1553 347
rect 1519 265 1553 321
rect 1587 485 1639 527
rect 1621 451 1639 485
rect 1587 417 1639 451
rect 1621 383 1639 417
rect 1587 349 1639 383
rect 1621 315 1639 349
rect 1587 299 1639 315
rect 687 249 840 265
rect 687 233 806 249
rect 394 169 434 203
rect 394 157 468 169
rect 17 69 69 85
rect 103 59 119 93
rect 153 59 169 93
rect 203 69 237 85
rect 307 153 468 157
rect 543 191 619 207
rect 577 157 619 191
rect 307 123 428 153
rect 543 141 619 157
rect 666 215 806 233
rect 666 199 840 215
rect 880 249 1030 265
rect 880 215 994 249
rect 1028 215 1030 249
rect 880 199 1030 215
rect 1064 249 1124 265
rect 1064 215 1090 249
rect 1064 199 1124 215
rect 307 119 341 123
rect 666 107 700 199
rect 1064 165 1102 199
rect 1158 177 1272 265
rect 1307 249 1485 265
rect 1307 215 1451 249
rect 1307 199 1485 215
rect 1519 211 1639 265
rect 1158 167 1230 177
rect 307 69 341 85
rect 103 17 169 59
rect 375 55 391 89
rect 425 55 441 89
rect 554 73 584 107
rect 618 73 700 107
rect 854 133 1102 165
rect 375 17 441 55
rect 748 72 764 106
rect 798 72 814 106
rect 854 99 868 133
rect 902 131 1102 133
rect 1136 133 1230 167
rect 902 99 914 131
rect 854 83 914 99
rect 1022 89 1098 97
rect 748 17 814 72
rect 1022 55 1038 89
rect 1072 55 1098 89
rect 1136 66 1170 99
rect 1307 119 1373 199
rect 1519 165 1553 211
rect 1022 17 1098 55
rect 1204 59 1220 93
rect 1254 59 1272 93
rect 1204 17 1272 59
rect 1307 85 1324 119
rect 1358 85 1373 119
rect 1503 129 1553 165
rect 1307 51 1373 85
rect 1407 93 1468 109
rect 1407 59 1418 93
rect 1452 59 1468 93
rect 1407 17 1468 59
rect 1537 95 1553 129
rect 1503 51 1553 95
rect 1587 161 1639 177
rect 1621 127 1639 161
rect 1587 93 1639 127
rect 1621 59 1639 93
rect 1587 17 1639 59
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1656 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 1593 527 1627 561
rect 122 289 156 323
rect 214 375 237 391
rect 237 375 248 391
rect 214 357 248 375
rect 586 365 620 391
rect 586 357 619 365
rect 619 357 620 365
rect 494 321 528 323
rect 494 289 517 321
rect 517 289 528 321
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1593 -17 1627 17
<< metal1 >>
rect 0 561 1656 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1656 561
rect 0 496 1656 527
rect 202 391 260 397
rect 202 357 214 391
rect 248 388 260 391
rect 574 391 632 397
rect 574 388 586 391
rect 248 360 586 388
rect 248 357 260 360
rect 202 351 260 357
rect 574 357 586 360
rect 620 357 632 391
rect 574 351 632 357
rect 110 323 168 329
rect 110 289 122 323
rect 156 320 168 323
rect 482 323 540 329
rect 482 320 494 323
rect 156 292 494 320
rect 156 289 168 292
rect 110 283 168 289
rect 482 289 494 292
rect 528 289 540 323
rect 482 283 540 289
rect 0 17 1656 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1656 17
rect 0 -48 1656 -17
<< labels >>
flabel locali s 1138 425 1172 459 0 FreeSans 200 0 0 0 Q
port 8 nsew signal output
flabel locali s 1136 85 1170 119 0 FreeSans 200 0 0 0 Q
port 8 nsew signal output
flabel locali s 1230 221 1264 255 0 FreeSans 200 0 0 0 Q
port 8 nsew signal output
flabel locali s 960 221 994 255 0 FreeSans 200 0 0 0 RESET_B
port 3 nsew signal input
flabel locali s 1599 221 1633 255 0 FreeSans 400 0 0 0 Q_N
port 9 nsew signal output
flabel locali s 1507 425 1541 459 0 FreeSans 400 0 0 0 Q_N
port 9 nsew signal output
flabel locali s 1507 357 1541 391 0 FreeSans 400 0 0 0 Q_N
port 9 nsew signal output
flabel locali s 1507 85 1541 119 0 FreeSans 400 0 0 0 Q_N
port 9 nsew signal output
flabel locali s 310 221 344 255 0 FreeSans 200 0 0 0 D
port 1 nsew signal input
flabel locali s 30 221 64 255 0 FreeSans 200 0 0 0 GATE
port 2 nsew clock input
flabel locali s 30 289 64 323 0 FreeSans 200 0 0 0 GATE
port 2 nsew clock input
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 4 nsew ground bidirectional abutment
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 7 nsew power bidirectional abutment
flabel nwell s 30 527 64 561 0 FreeSans 200 0 0 0 VPB
port 6 nsew power bidirectional
flabel nwell s 47 544 47 544 0 FreeSans 200 0 0 0 VPB
port 6 nsew
flabel pwell s 30 -17 64 17 0 FreeSans 200 0 0 0 VNB
port 5 nsew ground bidirectional
flabel pwell s 47 0 47 0 0 FreeSans 200 0 0 0 VNB
port 5 nsew
rlabel comment s 0 0 0 0 4 dlrbp_2
rlabel metal1 s 0 -48 1656 48 1 VGND
port 4 nsew ground bidirectional abutment
rlabel metal1 s 0 496 1656 592 1 VPWR
port 7 nsew power bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 1656 544
string GDS_END 2724808
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 2709966
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string path 0.000 0.000 41.400 0.000 
<< end >>
