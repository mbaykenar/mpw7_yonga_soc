magic
tech sky130A
magscale 1 2
timestamp 1649977179
<< nwell >>
rect -38 261 2522 582
<< pwell >>
rect 1 201 610 203
rect 1019 201 2480 203
rect 1 23 2480 201
rect 1 21 1106 23
rect 2192 21 2480 23
rect 29 -17 63 21
<< scnmos >>
rect 79 47 109 177
rect 174 47 204 175
rect 362 49 392 177
rect 498 47 528 177
rect 689 47 719 175
rect 774 47 804 175
rect 978 47 1008 175
rect 1126 49 1156 177
rect 1314 49 1344 177
rect 1399 49 1429 177
rect 1587 49 1617 177
rect 1675 49 1705 177
rect 1941 49 1971 177
rect 2025 49 2055 177
rect 2272 47 2302 177
rect 2356 47 2386 177
<< scpmoshvt >>
rect 83 297 113 497
rect 173 297 203 497
rect 365 297 395 497
rect 478 297 508 497
rect 689 297 719 465
rect 774 297 804 465
rect 985 297 1015 465
rect 1082 322 1112 490
rect 1302 297 1332 465
rect 1386 297 1416 465
rect 1692 315 1722 483
rect 1776 315 1806 483
rect 1944 297 1974 497
rect 2028 297 2058 497
rect 2272 297 2302 497
rect 2356 297 2386 497
<< ndiff >>
rect 27 161 79 177
rect 27 127 35 161
rect 69 127 79 161
rect 27 93 79 127
rect 27 59 35 93
rect 69 59 79 93
rect 27 47 79 59
rect 109 175 159 177
rect 109 93 174 175
rect 109 59 119 93
rect 153 59 174 93
rect 109 47 174 59
rect 204 161 256 175
rect 204 127 214 161
rect 248 127 256 161
rect 204 93 256 127
rect 204 59 214 93
rect 248 59 256 93
rect 204 47 256 59
rect 310 163 362 177
rect 310 129 318 163
rect 352 129 362 163
rect 310 95 362 129
rect 310 61 318 95
rect 352 61 362 95
rect 310 49 362 61
rect 392 93 498 177
rect 392 59 402 93
rect 436 59 498 93
rect 392 49 498 59
rect 431 47 498 49
rect 528 169 584 177
rect 1045 175 1126 177
rect 528 135 538 169
rect 572 135 584 169
rect 528 127 584 135
rect 528 47 578 127
rect 639 104 689 175
rect 637 93 689 104
rect 637 59 645 93
rect 679 59 689 93
rect 637 47 689 59
rect 719 161 774 175
rect 719 127 730 161
rect 764 127 774 161
rect 719 47 774 127
rect 804 163 872 175
rect 804 129 830 163
rect 864 129 872 163
rect 804 47 872 129
rect 926 101 978 175
rect 926 67 934 101
rect 968 67 978 101
rect 926 47 978 67
rect 1008 169 1126 175
rect 1008 135 1070 169
rect 1104 135 1126 169
rect 1008 49 1126 135
rect 1156 113 1208 177
rect 1156 79 1166 113
rect 1200 79 1208 113
rect 1156 49 1208 79
rect 1262 114 1314 177
rect 1262 80 1270 114
rect 1304 80 1314 114
rect 1262 49 1314 80
rect 1344 169 1399 177
rect 1344 135 1354 169
rect 1388 135 1399 169
rect 1344 49 1399 135
rect 1429 153 1481 177
rect 1429 119 1439 153
rect 1473 119 1481 153
rect 1429 49 1481 119
rect 1535 149 1587 177
rect 1535 115 1543 149
rect 1577 115 1587 149
rect 1535 49 1587 115
rect 1617 169 1675 177
rect 1617 135 1631 169
rect 1665 135 1675 169
rect 1617 49 1675 135
rect 1705 169 1761 177
rect 1705 135 1715 169
rect 1749 135 1761 169
rect 1705 49 1761 135
rect 1887 103 1941 177
rect 1887 69 1897 103
rect 1931 69 1941 103
rect 1887 49 1941 69
rect 1971 97 2025 177
rect 1971 63 1981 97
rect 2015 63 2025 97
rect 1971 49 2025 63
rect 2055 165 2107 177
rect 2055 131 2065 165
rect 2099 131 2107 165
rect 2055 97 2107 131
rect 2055 63 2065 97
rect 2099 63 2107 97
rect 2055 49 2107 63
rect 2218 127 2272 177
rect 2218 93 2228 127
rect 2262 93 2272 127
rect 1008 47 1080 49
rect 2218 47 2272 93
rect 2302 163 2356 177
rect 2302 129 2312 163
rect 2346 129 2356 163
rect 2302 95 2356 129
rect 2302 61 2312 95
rect 2346 61 2356 95
rect 2302 47 2356 61
rect 2386 163 2454 177
rect 2386 129 2412 163
rect 2446 129 2454 163
rect 2386 95 2454 129
rect 2386 61 2412 95
rect 2446 61 2454 95
rect 2386 47 2454 61
<< pdiff >>
rect 27 477 83 497
rect 27 443 39 477
rect 73 443 83 477
rect 27 409 83 443
rect 27 375 39 409
rect 73 375 83 409
rect 27 341 83 375
rect 27 307 39 341
rect 73 307 83 341
rect 27 297 83 307
rect 113 486 173 497
rect 113 452 129 486
rect 163 452 173 486
rect 113 297 173 452
rect 203 343 255 497
rect 203 309 213 343
rect 247 309 255 343
rect 203 297 255 309
rect 310 345 365 497
rect 310 311 318 345
rect 352 311 365 345
rect 310 297 365 311
rect 395 481 478 497
rect 395 447 429 481
rect 463 447 478 481
rect 395 297 478 447
rect 508 343 560 497
rect 508 309 518 343
rect 552 309 560 343
rect 508 297 560 309
rect 617 493 674 505
rect 617 459 629 493
rect 663 465 674 493
rect 920 493 970 505
rect 663 459 689 465
rect 617 297 689 459
rect 719 341 774 465
rect 719 307 729 341
rect 763 307 774 341
rect 719 297 774 307
rect 804 425 856 465
rect 804 391 814 425
rect 848 391 856 425
rect 804 297 856 391
rect 920 459 928 493
rect 962 465 970 493
rect 1030 465 1082 490
rect 962 459 985 465
rect 920 341 985 459
rect 920 307 941 341
rect 975 307 985 341
rect 920 297 985 307
rect 1015 446 1082 465
rect 1015 412 1025 446
rect 1059 412 1082 446
rect 1015 322 1082 412
rect 1112 390 1164 490
rect 1821 497 1926 505
rect 1821 493 1944 497
rect 1821 483 1861 493
rect 1112 356 1122 390
rect 1156 356 1164 390
rect 1112 322 1164 356
rect 1241 341 1302 465
rect 1015 297 1067 322
rect 1241 307 1258 341
rect 1292 307 1302 341
rect 1241 297 1302 307
rect 1332 341 1386 465
rect 1332 307 1342 341
rect 1376 307 1386 341
rect 1332 297 1386 307
rect 1416 363 1584 465
rect 1640 425 1692 483
rect 1640 391 1648 425
rect 1682 391 1692 425
rect 1640 380 1692 391
rect 1416 352 1588 363
rect 1416 318 1546 352
rect 1580 318 1588 352
rect 1416 308 1588 318
rect 1642 315 1692 380
rect 1722 357 1776 483
rect 1722 323 1732 357
rect 1766 323 1776 357
rect 1722 315 1776 323
rect 1806 459 1861 483
rect 1895 459 1944 493
rect 1806 341 1944 459
rect 1806 315 1900 341
rect 1416 307 1587 308
rect 1416 297 1585 307
rect 1862 307 1900 315
rect 1934 307 1944 341
rect 1862 297 1944 307
rect 1974 489 2028 497
rect 1974 455 1984 489
rect 2018 455 2028 489
rect 1974 297 2028 455
rect 2058 431 2114 497
rect 2058 397 2069 431
rect 2103 397 2114 431
rect 2058 297 2114 397
rect 2220 480 2272 497
rect 2220 446 2228 480
rect 2262 446 2272 480
rect 2220 412 2272 446
rect 2220 378 2228 412
rect 2262 378 2272 412
rect 2220 344 2272 378
rect 2220 310 2228 344
rect 2262 310 2272 344
rect 2220 297 2272 310
rect 2302 475 2356 497
rect 2302 441 2312 475
rect 2346 441 2356 475
rect 2302 407 2356 441
rect 2302 373 2312 407
rect 2346 373 2356 407
rect 2302 297 2356 373
rect 2386 477 2443 497
rect 2386 443 2397 477
rect 2431 443 2443 477
rect 2386 409 2443 443
rect 2386 375 2397 409
rect 2431 375 2443 409
rect 2386 297 2443 375
<< ndiffc >>
rect 35 127 69 161
rect 35 59 69 93
rect 119 59 153 93
rect 214 127 248 161
rect 214 59 248 93
rect 318 129 352 163
rect 318 61 352 95
rect 402 59 436 93
rect 538 135 572 169
rect 645 59 679 93
rect 730 127 764 161
rect 830 129 864 163
rect 934 67 968 101
rect 1070 135 1104 169
rect 1166 79 1200 113
rect 1270 80 1304 114
rect 1354 135 1388 169
rect 1439 119 1473 153
rect 1543 115 1577 149
rect 1631 135 1665 169
rect 1715 135 1749 169
rect 1897 69 1931 103
rect 1981 63 2015 97
rect 2065 131 2099 165
rect 2065 63 2099 97
rect 2228 93 2262 127
rect 2312 129 2346 163
rect 2312 61 2346 95
rect 2412 129 2446 163
rect 2412 61 2446 95
<< pdiffc >>
rect 39 443 73 477
rect 39 375 73 409
rect 39 307 73 341
rect 129 452 163 486
rect 213 309 247 343
rect 318 311 352 345
rect 429 447 463 481
rect 518 309 552 343
rect 629 459 663 493
rect 729 307 763 341
rect 814 391 848 425
rect 928 459 962 493
rect 941 307 975 341
rect 1025 412 1059 446
rect 1122 356 1156 390
rect 1258 307 1292 341
rect 1342 307 1376 341
rect 1648 391 1682 425
rect 1546 318 1580 352
rect 1732 323 1766 357
rect 1861 459 1895 493
rect 1900 307 1934 341
rect 1984 455 2018 489
rect 2069 397 2103 431
rect 2228 446 2262 480
rect 2228 378 2262 412
rect 2228 310 2262 344
rect 2312 441 2346 475
rect 2312 373 2346 407
rect 2397 443 2431 477
rect 2397 375 2431 409
<< poly >>
rect 83 497 113 523
rect 173 497 203 523
rect 365 497 395 523
rect 478 497 508 523
rect 689 465 719 491
rect 774 465 804 491
rect 985 465 1015 491
rect 1082 490 1112 516
rect 1302 465 1332 491
rect 1386 465 1416 491
rect 1692 483 1722 509
rect 1776 483 1806 509
rect 1944 497 1974 523
rect 2028 497 2058 523
rect 2272 497 2302 523
rect 2356 497 2386 523
rect 83 265 113 297
rect 173 265 203 297
rect 365 265 395 297
rect 478 265 508 297
rect 689 265 719 297
rect 67 249 131 265
rect 67 215 85 249
rect 119 215 131 249
rect 67 199 131 215
rect 173 249 395 265
rect 173 215 218 249
rect 252 215 395 249
rect 173 199 395 215
rect 439 249 719 265
rect 439 215 449 249
rect 483 215 719 249
rect 439 199 719 215
rect 79 177 109 199
rect 174 175 204 199
rect 362 177 392 199
rect 498 177 528 199
rect 79 21 109 47
rect 174 21 204 47
rect 362 23 392 49
rect 689 175 719 199
rect 774 265 804 297
rect 985 265 1015 297
rect 1082 265 1112 322
rect 1692 300 1722 315
rect 1302 265 1332 297
rect 1386 265 1416 297
rect 1601 270 1722 300
rect 1601 265 1633 270
rect 774 249 1015 265
rect 774 215 830 249
rect 864 215 1015 249
rect 774 199 1015 215
rect 1080 249 1179 265
rect 1080 215 1135 249
rect 1169 215 1179 249
rect 1080 199 1179 215
rect 1227 249 1344 265
rect 1227 215 1237 249
rect 1271 215 1344 249
rect 1227 199 1344 215
rect 1386 249 1633 265
rect 1386 215 1490 249
rect 1524 215 1633 249
rect 1776 222 1806 315
rect 1944 265 1974 297
rect 2028 265 2058 297
rect 2272 265 2302 297
rect 2356 265 2386 297
rect 1386 199 1633 215
rect 1675 221 1806 222
rect 1901 249 1974 265
rect 774 175 804 199
rect 978 175 1008 199
rect 1126 177 1156 199
rect 1314 177 1344 199
rect 1399 177 1429 199
rect 1587 177 1617 199
rect 1675 192 1851 221
rect 1901 215 1911 249
rect 1945 215 1974 249
rect 1901 199 1974 215
rect 2025 249 2086 265
rect 2025 215 2036 249
rect 2070 215 2086 249
rect 2025 199 2086 215
rect 2228 249 2302 265
rect 2228 215 2242 249
rect 2276 215 2302 249
rect 2228 199 2302 215
rect 2344 249 2398 265
rect 2344 215 2354 249
rect 2388 215 2398 249
rect 2344 199 2398 215
rect 1675 177 1705 192
rect 1797 171 1851 192
rect 1941 177 1971 199
rect 2025 177 2055 199
rect 2272 177 2302 199
rect 2356 177 2386 199
rect 1797 137 1807 171
rect 1841 137 1851 171
rect 1797 121 1851 137
rect 498 21 528 47
rect 689 21 719 47
rect 774 21 804 47
rect 978 21 1008 47
rect 1126 23 1156 49
rect 1314 23 1344 49
rect 1399 23 1429 49
rect 1587 23 1617 49
rect 1675 21 1705 49
rect 1941 21 1971 49
rect 2025 21 2055 49
rect 2272 21 2302 47
rect 2356 21 2386 47
<< polycont >>
rect 85 215 119 249
rect 218 215 252 249
rect 449 215 483 249
rect 830 215 864 249
rect 1135 215 1169 249
rect 1237 215 1271 249
rect 1490 215 1524 249
rect 1911 215 1945 249
rect 2036 215 2070 249
rect 2242 215 2276 249
rect 2354 215 2388 249
rect 1807 137 1841 171
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2053 561
rect 2087 527 2145 561
rect 2179 527 2237 561
rect 2271 527 2329 561
rect 2363 527 2421 561
rect 2455 527 2484 561
rect 17 477 79 493
rect 17 443 39 477
rect 73 443 79 477
rect 113 486 186 527
rect 113 452 129 486
rect 163 452 186 486
rect 413 481 479 527
rect 413 447 429 481
rect 463 447 479 481
rect 527 459 629 493
rect 663 459 928 493
rect 962 459 990 493
rect 1025 459 1512 493
rect 17 413 79 443
rect 527 413 561 459
rect 17 409 561 413
rect 17 375 39 409
rect 73 379 561 409
rect 606 391 814 425
rect 848 391 864 425
rect 73 375 89 379
rect 17 341 89 375
rect 17 307 39 341
rect 73 307 89 341
rect 197 323 213 343
rect 17 300 89 307
rect 123 309 213 323
rect 247 309 263 343
rect 17 161 51 300
rect 123 291 263 309
rect 122 289 263 291
rect 298 311 318 345
rect 352 311 368 345
rect 298 300 368 311
rect 298 289 364 300
rect 122 276 163 289
rect 122 265 156 276
rect 85 249 156 265
rect 119 215 156 249
rect 190 249 288 255
rect 190 215 218 249
rect 252 215 288 249
rect 85 199 156 215
rect 119 181 156 199
rect 323 181 364 289
rect 403 282 438 345
rect 472 323 518 343
rect 472 289 490 323
rect 552 309 572 343
rect 524 289 572 309
rect 398 255 438 282
rect 432 249 499 255
rect 432 221 449 249
rect 398 215 449 221
rect 483 215 499 249
rect 119 161 264 181
rect 17 127 35 161
rect 69 127 85 161
rect 119 147 214 161
rect 17 93 85 127
rect 198 127 214 147
rect 248 127 264 161
rect 17 59 35 93
rect 69 59 85 93
rect 17 51 85 59
rect 119 93 153 109
rect 119 17 153 59
rect 198 93 264 127
rect 198 59 214 93
rect 248 59 264 93
rect 198 51 264 59
rect 300 177 364 181
rect 300 163 504 177
rect 300 129 318 163
rect 352 143 504 163
rect 352 129 368 143
rect 300 95 368 129
rect 300 61 318 95
rect 352 61 368 95
rect 300 51 368 61
rect 402 93 436 109
rect 402 17 436 59
rect 470 85 504 143
rect 538 169 572 289
rect 538 119 572 135
rect 606 93 640 391
rect 831 357 864 391
rect 674 341 763 357
rect 674 307 729 341
rect 941 341 975 459
rect 674 291 763 307
rect 674 187 708 291
rect 814 289 873 323
rect 814 249 907 289
rect 814 215 830 249
rect 864 232 907 249
rect 864 215 880 232
rect 941 185 975 307
rect 1025 446 1059 459
rect 1025 264 1059 412
rect 1095 391 1175 406
rect 1095 357 1114 391
rect 1148 390 1175 391
rect 1095 356 1122 357
rect 1156 356 1175 390
rect 1095 340 1175 356
rect 1258 391 1444 425
rect 1258 341 1292 391
rect 1221 289 1230 323
rect 1264 289 1292 307
rect 1342 341 1376 357
rect 1025 230 1101 264
rect 1064 185 1101 230
rect 1135 255 1185 265
rect 1342 255 1376 307
rect 1135 249 1136 255
rect 1170 221 1185 255
rect 1169 215 1185 221
rect 1135 199 1185 215
rect 1221 249 1287 255
rect 1221 215 1237 249
rect 1271 215 1287 249
rect 1221 187 1287 215
rect 896 181 1029 185
rect 814 163 1029 181
rect 1064 173 1104 185
rect 1067 169 1104 173
rect 1067 168 1070 169
rect 708 153 730 161
rect 674 127 730 153
rect 764 127 780 161
rect 814 129 830 163
rect 864 161 1029 163
rect 864 156 1031 161
rect 864 151 1034 156
rect 864 147 912 151
rect 985 148 1034 151
rect 985 147 1036 148
rect 864 129 880 147
rect 990 143 1036 147
rect 996 138 1036 143
rect 1000 131 1036 138
rect 930 101 968 117
rect 930 93 934 101
rect 606 85 645 93
rect 470 59 645 85
rect 679 67 934 93
rect 679 59 968 67
rect 470 51 968 59
rect 1002 85 1036 131
rect 1221 153 1230 187
rect 1264 153 1287 187
rect 1221 148 1287 153
rect 1356 221 1376 255
rect 1322 185 1376 221
rect 1410 235 1444 391
rect 1478 285 1512 459
rect 1546 459 1861 493
rect 1895 459 1931 493
rect 1546 352 1592 459
rect 1629 391 1648 425
rect 1682 391 1850 425
rect 1580 318 1592 352
rect 1546 302 1592 318
rect 1478 280 1515 285
rect 1478 275 1519 280
rect 1478 255 1524 275
rect 1490 249 1524 255
rect 1410 226 1449 235
rect 1410 212 1456 226
rect 1413 209 1456 212
rect 1418 202 1456 209
rect 1322 169 1388 185
rect 1322 151 1354 169
rect 1070 119 1104 135
rect 1354 119 1388 135
rect 1422 153 1456 202
rect 1490 199 1524 215
rect 1558 165 1592 302
rect 1645 323 1732 357
rect 1766 323 1782 357
rect 1645 289 1692 323
rect 1726 289 1782 323
rect 1645 185 1681 289
rect 1816 255 1850 357
rect 1884 341 1931 459
rect 1968 489 2035 527
rect 1968 455 1984 489
rect 2018 455 2035 489
rect 2069 431 2138 493
rect 2103 397 2138 431
rect 2069 391 2138 397
rect 2069 375 2104 391
rect 1884 307 1900 341
rect 1934 307 2070 341
rect 1884 299 2070 307
rect 1422 119 1439 153
rect 1473 119 1489 153
rect 1541 149 1592 165
rect 1541 115 1543 149
rect 1577 115 1592 149
rect 1631 169 1681 185
rect 1665 135 1681 169
rect 1631 119 1681 135
rect 1715 221 1850 255
rect 1895 249 1973 265
rect 1715 169 1749 221
rect 1895 215 1911 249
rect 1945 215 1973 249
rect 1938 187 1973 215
rect 2036 249 2070 299
rect 2036 199 2070 215
rect 1818 171 1860 187
rect 1784 137 1807 153
rect 1841 137 1860 171
rect 1938 147 2002 187
rect 2104 165 2138 357
rect 1715 119 1749 135
rect 2049 131 2065 165
rect 2099 131 2138 165
rect 1150 85 1166 113
rect 1002 79 1166 85
rect 1200 79 1220 113
rect 1002 51 1220 79
rect 1254 80 1270 114
rect 1304 85 1320 114
rect 1541 85 1592 115
rect 1880 85 1897 103
rect 1304 80 1897 85
rect 1254 69 1897 80
rect 1931 69 1947 103
rect 1254 51 1947 69
rect 1981 97 2015 113
rect 1981 17 2015 63
rect 2049 97 2138 131
rect 2049 63 2065 97
rect 2099 63 2138 97
rect 2049 57 2138 63
rect 2174 480 2278 493
rect 2174 446 2228 480
rect 2262 446 2278 480
rect 2174 412 2278 446
rect 2174 378 2228 412
rect 2262 378 2278 412
rect 2174 344 2278 378
rect 2312 475 2363 527
rect 2346 441 2363 475
rect 2312 407 2363 441
rect 2346 373 2363 407
rect 2312 357 2363 373
rect 2397 477 2467 493
rect 2431 443 2467 477
rect 2397 409 2467 443
rect 2431 375 2467 409
rect 2397 357 2467 375
rect 2174 310 2228 344
rect 2262 310 2278 344
rect 2174 299 2278 310
rect 2174 165 2208 299
rect 2326 289 2336 323
rect 2370 289 2388 323
rect 2242 255 2292 265
rect 2242 249 2244 255
rect 2278 221 2292 255
rect 2276 215 2292 221
rect 2242 199 2292 215
rect 2326 249 2388 289
rect 2326 215 2354 249
rect 2326 199 2388 215
rect 2422 165 2467 357
rect 2174 127 2262 165
rect 2174 93 2228 127
rect 2174 54 2262 93
rect 2296 163 2362 165
rect 2296 129 2312 163
rect 2346 129 2362 163
rect 2296 95 2362 129
rect 2296 61 2312 95
rect 2346 61 2362 95
rect 2296 17 2362 61
rect 2396 163 2467 165
rect 2396 129 2412 163
rect 2446 129 2467 163
rect 2396 95 2467 129
rect 2396 61 2412 95
rect 2446 61 2467 95
rect 2396 51 2467 61
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2053 17
rect 2087 -17 2145 17
rect 2179 -17 2237 17
rect 2271 -17 2329 17
rect 2363 -17 2421 17
rect 2455 -17 2484 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 1593 527 1627 561
rect 1685 527 1719 561
rect 1777 527 1811 561
rect 1869 527 1903 561
rect 1961 527 1995 561
rect 2053 527 2087 561
rect 2145 527 2179 561
rect 2237 527 2271 561
rect 2329 527 2363 561
rect 2421 527 2455 561
rect 490 309 518 323
rect 518 309 524 323
rect 490 289 524 309
rect 398 221 432 255
rect 797 357 831 391
rect 873 289 907 323
rect 674 153 708 187
rect 1114 390 1148 391
rect 1114 357 1122 390
rect 1122 357 1148 390
rect 1230 307 1258 323
rect 1258 307 1264 323
rect 1230 289 1264 307
rect 1136 249 1170 255
rect 1136 221 1169 249
rect 1169 221 1170 249
rect 1230 153 1264 187
rect 1322 221 1356 255
rect 1816 357 1850 391
rect 1692 289 1726 323
rect 2104 357 2138 391
rect 1784 171 1818 187
rect 1784 153 1807 171
rect 1807 153 1818 171
rect 2336 289 2370 323
rect 2244 249 2278 255
rect 2244 221 2276 249
rect 2276 221 2278 249
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1593 -17 1627 17
rect 1685 -17 1719 17
rect 1777 -17 1811 17
rect 1869 -17 1903 17
rect 1961 -17 1995 17
rect 2053 -17 2087 17
rect 2145 -17 2179 17
rect 2237 -17 2271 17
rect 2329 -17 2363 17
rect 2421 -17 2455 17
<< metal1 >>
rect 0 561 2484 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2053 561
rect 2087 527 2145 561
rect 2179 527 2237 561
rect 2271 527 2329 561
rect 2363 527 2421 561
rect 2455 527 2484 561
rect 0 496 2484 527
rect 785 391 843 397
rect 785 357 797 391
rect 831 388 843 391
rect 1102 391 1160 397
rect 1102 388 1114 391
rect 831 360 1114 388
rect 831 357 843 360
rect 785 351 843 357
rect 1102 357 1114 360
rect 1148 357 1160 391
rect 1102 351 1160 357
rect 1804 391 1862 397
rect 1804 357 1816 391
rect 1850 388 1862 391
rect 2092 391 2150 397
rect 2092 388 2104 391
rect 1850 360 2104 388
rect 1850 357 1862 360
rect 1804 351 1862 357
rect 2092 357 2104 360
rect 2138 357 2150 391
rect 2092 351 2150 357
rect 478 323 536 329
rect 478 289 490 323
rect 524 320 536 323
rect 861 323 919 329
rect 861 320 873 323
rect 524 292 873 320
rect 524 289 536 292
rect 478 283 536 289
rect 861 289 873 292
rect 907 320 919 323
rect 1218 323 1276 329
rect 1218 320 1230 323
rect 907 292 1230 320
rect 907 289 919 292
rect 861 283 919 289
rect 1218 289 1230 292
rect 1264 289 1276 323
rect 1218 283 1276 289
rect 1680 323 1738 329
rect 1680 289 1692 323
rect 1726 320 1738 323
rect 2324 323 2382 329
rect 2324 320 2336 323
rect 1726 292 2336 320
rect 1726 289 1738 292
rect 1680 283 1738 289
rect 2324 289 2336 292
rect 2370 289 2382 323
rect 2324 283 2382 289
rect 386 255 444 261
rect 386 221 398 255
rect 432 252 444 255
rect 1124 255 1182 261
rect 1124 252 1136 255
rect 432 224 1136 252
rect 432 221 444 224
rect 386 215 444 221
rect 1124 221 1136 224
rect 1170 221 1182 255
rect 1124 215 1182 221
rect 1310 255 1368 261
rect 1310 221 1322 255
rect 1356 252 1368 255
rect 2232 255 2290 261
rect 2232 252 2244 255
rect 1356 224 2244 252
rect 1356 221 1368 224
rect 1310 215 1368 221
rect 2232 221 2244 224
rect 2278 221 2290 255
rect 2232 215 2290 221
rect 662 187 720 193
rect 662 153 674 187
rect 708 184 720 187
rect 1218 187 1276 193
rect 1218 184 1230 187
rect 708 156 1230 184
rect 708 153 720 156
rect 662 147 720 153
rect 1218 153 1230 156
rect 1264 184 1276 187
rect 1772 187 1830 193
rect 1772 184 1784 187
rect 1264 156 1784 184
rect 1264 153 1276 156
rect 1218 147 1276 153
rect 1772 153 1784 156
rect 1818 153 1830 187
rect 1772 147 1830 153
rect 0 17 2484 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2053 17
rect 2087 -17 2145 17
rect 2179 -17 2237 17
rect 2271 -17 2329 17
rect 2363 -17 2421 17
rect 2455 -17 2484 17
rect 0 -48 2484 -17
<< labels >>
flabel locali s 2244 357 2278 391 0 FreeSans 300 0 0 0 COUT
port 8 nsew signal output
flabel locali s 398 221 432 255 0 FreeSans 300 0 0 0 B
port 2 nsew signal input
flabel locali s 213 221 247 255 0 FreeSans 300 180 0 0 A
port 1 nsew signal input
flabel locali s 2428 221 2462 255 0 FreeSans 300 0 0 0 SUM
port 9 nsew signal output
flabel locali s 1968 153 2002 187 0 FreeSans 340 0 0 0 CI
port 3 nsew signal input
flabel metal1 s 415 238 415 238 0 FreeSans 300 0 0 0 B
port 2 nsew
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 7 nsew power bidirectional abutment
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 4 nsew ground bidirectional abutment
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 5 nsew ground bidirectional
flabel nwell s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 6 nsew power bidirectional
rlabel comment s 0 0 0 0 4 fah_1
rlabel locali s 1135 199 1185 265 1 B
port 2 nsew signal input
rlabel metal1 s 1124 252 1182 261 1 B
port 2 nsew signal input
rlabel metal1 s 1124 215 1182 224 1 B
port 2 nsew signal input
rlabel metal1 s 386 252 444 261 1 B
port 2 nsew signal input
rlabel metal1 s 386 224 1182 252 1 B
port 2 nsew signal input
rlabel metal1 s 386 215 444 224 1 B
port 2 nsew signal input
rlabel metal1 s 0 -48 2484 48 1 VGND
port 4 nsew ground bidirectional abutment
rlabel metal1 s 0 496 2484 592 1 VPWR
port 7 nsew power bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 2484 544
string GDS_END 2113468
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 2094028
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string path 0.000 13.600 62.100 13.600 
<< end >>
