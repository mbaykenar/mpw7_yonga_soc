magic
tech sky130A
magscale 1 2
timestamp 1649977179
<< nwell >>
rect 106 836 1440 844
rect 1777 836 2135 844
rect 106 728 2445 836
rect 106 512 2459 728
<< pwell >>
rect 706 252 840 360
rect 2011 252 2145 360
rect 146 116 2339 252
rect 146 8 1258 116
rect 1451 8 2339 116
rect 146 0 424 8
rect 756 0 1034 8
rect 1451 0 1729 8
rect 2061 0 2339 8
<< mvnmos >>
rect 225 26 345 226
rect 511 142 711 226
rect 835 26 955 226
rect 1121 142 1321 226
rect 1530 26 1650 226
rect 1816 142 2016 226
rect 2140 26 2260 226
<< mvpmos >>
rect 225 578 425 662
rect 591 578 711 778
rect 835 578 1035 662
rect 1201 578 1321 778
rect 1530 578 1730 662
rect 1896 578 2016 778
rect 2140 578 2340 662
<< mvndiff >>
rect 172 208 225 226
rect 172 174 180 208
rect 214 174 225 208
rect 172 140 225 174
rect 172 106 180 140
rect 214 106 225 140
rect 172 72 225 106
rect 172 38 180 72
rect 214 38 225 72
rect 172 26 225 38
rect 345 208 398 226
rect 345 174 356 208
rect 390 174 398 208
rect 345 140 398 174
rect 458 214 511 226
rect 458 180 466 214
rect 500 180 511 214
rect 458 142 511 180
rect 711 214 835 226
rect 711 180 722 214
rect 756 180 790 214
rect 824 180 835 214
rect 711 146 835 180
rect 711 142 790 146
rect 345 106 356 140
rect 390 106 398 140
rect 345 72 398 106
rect 345 38 356 72
rect 390 38 398 72
rect 782 112 790 142
rect 824 112 835 146
rect 782 78 835 112
rect 345 26 398 38
rect 782 44 790 78
rect 824 44 835 78
rect 782 26 835 44
rect 955 214 1008 226
rect 955 180 966 214
rect 1000 180 1008 214
rect 955 146 1008 180
rect 955 112 966 146
rect 1000 112 1008 146
rect 1068 214 1121 226
rect 1068 180 1076 214
rect 1110 180 1121 214
rect 1068 142 1121 180
rect 1321 214 1374 226
rect 1321 180 1332 214
rect 1366 180 1374 214
rect 1321 142 1374 180
rect 1477 208 1530 226
rect 1477 174 1485 208
rect 1519 174 1530 208
rect 1477 140 1530 174
rect 955 78 1008 112
rect 955 44 966 78
rect 1000 44 1008 78
rect 1477 106 1485 140
rect 1519 106 1530 140
rect 1477 72 1530 106
rect 955 26 1008 44
rect 1477 38 1485 72
rect 1519 38 1530 72
rect 1477 26 1530 38
rect 1650 208 1703 226
rect 1650 174 1661 208
rect 1695 174 1703 208
rect 1650 140 1703 174
rect 1763 214 1816 226
rect 1763 180 1771 214
rect 1805 180 1816 214
rect 1763 142 1816 180
rect 2016 214 2140 226
rect 2016 180 2027 214
rect 2061 180 2095 214
rect 2129 180 2140 214
rect 2016 146 2140 180
rect 2016 142 2095 146
rect 1650 106 1661 140
rect 1695 106 1703 140
rect 1650 72 1703 106
rect 1650 38 1661 72
rect 1695 38 1703 72
rect 2087 112 2095 142
rect 2129 112 2140 146
rect 2087 78 2140 112
rect 1650 26 1703 38
rect 2087 44 2095 78
rect 2129 44 2140 78
rect 2087 26 2140 44
rect 2260 214 2313 226
rect 2260 180 2271 214
rect 2305 180 2313 214
rect 2260 146 2313 180
rect 2260 112 2271 146
rect 2305 112 2313 146
rect 2260 78 2313 112
rect 2260 44 2271 78
rect 2305 44 2313 78
rect 2260 26 2313 44
<< mvpdiff >>
rect 538 766 591 778
rect 538 732 546 766
rect 580 732 591 766
rect 538 698 591 732
rect 538 664 546 698
rect 580 664 591 698
rect 172 650 225 662
rect 172 616 180 650
rect 214 616 225 650
rect 172 578 225 616
rect 425 650 478 662
rect 425 616 436 650
rect 470 616 478 650
rect 425 578 478 616
rect 538 630 591 664
rect 538 596 546 630
rect 580 596 591 630
rect 538 578 591 596
rect 711 766 764 778
rect 711 732 722 766
rect 756 732 764 766
rect 1148 766 1201 778
rect 711 698 764 732
rect 711 664 722 698
rect 756 664 764 698
rect 1148 732 1156 766
rect 1190 732 1201 766
rect 1148 698 1201 732
rect 711 662 764 664
rect 1148 664 1156 698
rect 1190 664 1201 698
rect 711 650 835 662
rect 711 630 790 650
rect 711 596 722 630
rect 756 616 790 630
rect 824 616 835 650
rect 756 596 835 616
rect 711 578 835 596
rect 1035 650 1088 662
rect 1035 616 1046 650
rect 1080 616 1088 650
rect 1035 578 1088 616
rect 1148 630 1201 664
rect 1148 596 1156 630
rect 1190 596 1201 630
rect 1148 578 1201 596
rect 1321 766 1374 778
rect 1321 732 1332 766
rect 1366 732 1374 766
rect 1843 766 1896 778
rect 1321 698 1374 732
rect 1321 664 1332 698
rect 1366 664 1374 698
rect 1843 732 1851 766
rect 1885 732 1896 766
rect 1843 698 1896 732
rect 1321 630 1374 664
rect 1843 664 1851 698
rect 1885 664 1896 698
rect 1321 596 1332 630
rect 1366 596 1374 630
rect 1321 578 1374 596
rect 1477 650 1530 662
rect 1477 616 1485 650
rect 1519 616 1530 650
rect 1477 578 1530 616
rect 1730 650 1783 662
rect 1730 616 1741 650
rect 1775 616 1783 650
rect 1730 578 1783 616
rect 1843 630 1896 664
rect 1843 596 1851 630
rect 1885 596 1896 630
rect 1843 578 1896 596
rect 2016 766 2069 778
rect 2016 732 2027 766
rect 2061 732 2069 766
rect 2016 698 2069 732
rect 2016 664 2027 698
rect 2061 664 2069 698
rect 2016 662 2069 664
rect 2016 650 2140 662
rect 2016 630 2095 650
rect 2016 596 2027 630
rect 2061 616 2095 630
rect 2129 616 2140 650
rect 2061 596 2140 616
rect 2016 578 2140 596
rect 2340 650 2393 662
rect 2340 616 2351 650
rect 2385 616 2393 650
rect 2340 578 2393 616
<< mvndiffc >>
rect 180 174 214 208
rect 180 106 214 140
rect 180 38 214 72
rect 356 174 390 208
rect 466 180 500 214
rect 722 180 756 214
rect 790 180 824 214
rect 356 106 390 140
rect 356 38 390 72
rect 790 112 824 146
rect 790 44 824 78
rect 966 180 1000 214
rect 966 112 1000 146
rect 1076 180 1110 214
rect 1332 180 1366 214
rect 1485 174 1519 208
rect 966 44 1000 78
rect 1485 106 1519 140
rect 1485 38 1519 72
rect 1661 174 1695 208
rect 1771 180 1805 214
rect 2027 180 2061 214
rect 2095 180 2129 214
rect 1661 106 1695 140
rect 1661 38 1695 72
rect 2095 112 2129 146
rect 2095 44 2129 78
rect 2271 180 2305 214
rect 2271 112 2305 146
rect 2271 44 2305 78
<< mvpdiffc >>
rect 546 732 580 766
rect 546 664 580 698
rect 180 616 214 650
rect 436 616 470 650
rect 546 596 580 630
rect 722 732 756 766
rect 722 664 756 698
rect 1156 732 1190 766
rect 1156 664 1190 698
rect 722 596 756 630
rect 790 616 824 650
rect 1046 616 1080 650
rect 1156 596 1190 630
rect 1332 732 1366 766
rect 1332 664 1366 698
rect 1851 732 1885 766
rect 1851 664 1885 698
rect 1332 596 1366 630
rect 1485 616 1519 650
rect 1741 616 1775 650
rect 1851 596 1885 630
rect 2027 732 2061 766
rect 2027 664 2061 698
rect 2027 596 2061 630
rect 2095 616 2129 650
rect 2351 616 2385 650
<< psubdiff >>
rect 2037 300 2061 334
rect 2095 300 2119 334
rect 1777 34 1801 68
rect 1835 34 1929 68
rect 1963 34 1987 68
<< mvpsubdiff >>
rect 732 300 756 334
rect 790 300 814 334
rect 472 34 496 68
rect 530 34 624 68
rect 658 34 682 68
rect 1082 34 1106 68
rect 1140 34 1174 68
rect 1208 34 1232 68
<< mvnsubdiff >>
rect 186 736 210 770
rect 244 736 308 770
rect 342 736 406 770
rect 440 736 464 770
rect 838 736 862 770
rect 896 736 939 770
rect 973 736 1016 770
rect 1050 736 1074 770
rect 1491 736 1515 770
rect 1549 736 1613 770
rect 1647 736 1711 770
rect 1745 736 1769 770
rect 2143 736 2167 770
rect 2201 736 2244 770
rect 2278 736 2321 770
rect 2355 736 2379 770
<< psubdiffcont >>
rect 2061 300 2095 334
rect 1801 34 1835 68
rect 1929 34 1963 68
<< mvpsubdiffcont >>
rect 756 300 790 334
rect 496 34 530 68
rect 624 34 658 68
rect 1106 34 1140 68
rect 1174 34 1208 68
<< mvnsubdiffcont >>
rect 210 736 244 770
rect 308 736 342 770
rect 406 736 440 770
rect 862 736 896 770
rect 939 736 973 770
rect 1016 736 1050 770
rect 1515 736 1549 770
rect 1613 736 1647 770
rect 1711 736 1745 770
rect 2167 736 2201 770
rect 2244 736 2278 770
rect 2321 736 2355 770
<< poly >>
rect 591 778 711 804
rect 1201 778 1321 804
rect 1896 778 2016 804
rect 225 662 425 688
rect 835 662 1035 688
rect 1530 662 1730 688
rect 2140 662 2340 688
rect 225 552 425 578
rect 225 530 345 552
rect 225 496 274 530
rect 308 496 345 530
rect 591 504 711 578
rect 225 462 345 496
rect 225 428 274 462
rect 308 428 345 462
rect 225 226 345 428
rect 454 488 711 504
rect 835 552 1035 578
rect 835 498 955 552
rect 1201 504 1321 578
rect 454 454 470 488
rect 504 454 711 488
rect 454 420 711 454
rect 821 482 955 498
rect 821 448 837 482
rect 871 448 905 482
rect 939 448 955 482
rect 821 432 955 448
rect 454 386 470 420
rect 504 386 711 420
rect 454 370 711 386
rect 511 226 711 370
rect 835 226 955 432
rect 997 488 1321 504
rect 997 454 1013 488
rect 1047 454 1321 488
rect 997 420 1321 454
rect 997 386 1013 420
rect 1047 386 1321 420
rect 997 370 1321 386
rect 1121 226 1321 370
rect 1530 552 1730 578
rect 1530 530 1650 552
rect 1530 496 1579 530
rect 1613 496 1650 530
rect 1896 504 2016 578
rect 1530 462 1650 496
rect 1530 428 1579 462
rect 1613 428 1650 462
rect 1530 226 1650 428
rect 1759 488 2016 504
rect 2140 552 2340 578
rect 2140 498 2260 552
rect 1759 454 1775 488
rect 1809 454 2016 488
rect 1759 420 2016 454
rect 2126 482 2260 498
rect 2126 448 2142 482
rect 2176 448 2210 482
rect 2244 448 2260 482
rect 2126 432 2260 448
rect 1759 386 1775 420
rect 1809 386 2016 420
rect 1759 370 2016 386
rect 1816 226 2016 370
rect 2140 226 2260 432
rect 2302 488 2368 504
rect 2302 454 2318 488
rect 2352 454 2368 488
rect 2302 420 2368 454
rect 2302 386 2318 420
rect 2352 386 2368 420
rect 2302 370 2368 386
rect 511 116 711 142
rect 1121 116 1321 142
rect 1816 116 2016 142
rect 225 0 345 26
rect 835 0 955 26
rect 1530 0 1650 26
rect 2140 0 2260 26
<< polycont >>
rect 274 496 308 530
rect 274 428 308 462
rect 470 454 504 488
rect 837 448 871 482
rect 905 448 939 482
rect 470 386 504 420
rect 1013 454 1047 488
rect 1013 386 1047 420
rect 1579 496 1613 530
rect 1579 428 1613 462
rect 1775 454 1809 488
rect 2142 448 2176 482
rect 2210 448 2244 482
rect 1775 386 1809 420
rect 2318 454 2352 488
rect 2318 386 2352 420
<< locali >>
rect 180 770 464 782
rect 180 736 210 770
rect 244 736 308 770
rect 342 736 406 770
rect 440 736 464 770
rect 180 711 464 736
rect 180 677 241 711
rect 275 677 313 711
rect 347 706 464 711
rect 546 766 580 782
rect 180 650 347 677
rect 546 698 580 732
rect 214 616 347 650
rect 180 600 347 616
rect 398 650 470 666
rect 398 616 436 650
rect 398 600 470 616
rect 546 630 580 664
rect 232 496 274 530
rect 308 496 338 530
rect 232 462 338 496
rect 232 448 274 462
rect 308 448 338 462
rect 266 428 274 448
rect 266 414 304 428
rect 398 504 432 600
rect 398 498 504 504
rect 432 464 470 498
rect 398 454 470 464
rect 398 420 504 454
rect 180 160 214 174
rect 180 88 214 106
rect 180 22 214 38
rect 267 34 301 414
rect 398 386 470 420
rect 398 370 504 386
rect 546 482 580 596
rect 722 770 1074 782
rect 722 766 862 770
rect 756 736 862 766
rect 896 736 939 770
rect 973 736 1016 770
rect 1050 736 1074 770
rect 756 732 1074 736
rect 722 706 1074 732
rect 1122 766 1190 782
rect 1122 732 1156 766
rect 722 703 932 706
rect 722 698 740 703
rect 774 669 812 703
rect 846 669 884 703
rect 918 669 932 703
rect 756 664 932 669
rect 1122 698 1190 732
rect 722 650 932 664
rect 722 630 790 650
rect 756 616 790 630
rect 824 616 932 650
rect 756 596 932 616
rect 722 580 932 596
rect 1003 650 1088 666
rect 1003 616 1046 650
rect 1080 616 1088 650
rect 1003 600 1088 616
rect 1122 664 1156 698
rect 1122 630 1190 664
rect 1003 504 1037 600
rect 1122 596 1156 630
rect 1122 548 1190 596
rect 1260 766 1366 782
rect 1260 732 1332 766
rect 1260 711 1366 732
rect 1294 677 1332 711
rect 1260 664 1332 677
rect 1260 630 1366 664
rect 1260 596 1332 630
rect 1485 770 1769 782
rect 1485 736 1515 770
rect 1549 736 1613 770
rect 1647 736 1711 770
rect 1745 736 1769 770
rect 1485 711 1769 736
rect 1485 677 1546 711
rect 1580 677 1618 711
rect 1652 706 1769 711
rect 1851 766 1885 782
rect 1485 650 1652 677
rect 1851 698 1885 732
rect 1519 616 1652 650
rect 1485 600 1652 616
rect 1703 650 1775 666
rect 1703 616 1741 650
rect 1703 600 1775 616
rect 1851 630 1885 664
rect 1260 582 1366 596
rect 1332 580 1366 582
rect 1122 514 1128 548
rect 1162 514 1200 548
rect 1003 488 1060 504
rect 546 448 837 482
rect 871 448 905 482
rect 939 448 955 482
rect 1003 470 1013 488
rect 1047 454 1060 488
rect 546 414 564 448
rect 598 414 636 448
rect 1037 436 1060 454
rect 1003 420 1060 436
rect 398 224 432 370
rect 546 242 580 414
rect 821 368 859 402
rect 893 368 932 402
rect 356 208 432 224
rect 390 174 432 208
rect 356 140 432 174
rect 466 214 580 242
rect 500 180 580 214
rect 466 176 580 180
rect 620 318 756 334
rect 654 284 692 318
rect 726 300 756 318
rect 790 300 814 334
rect 726 284 814 300
rect 466 164 500 176
rect 390 106 432 140
rect 356 72 432 106
rect 390 38 432 72
rect 620 68 682 284
rect 356 22 432 38
rect 472 34 496 68
rect 530 34 624 68
rect 658 34 682 68
rect 722 214 756 230
rect 790 214 828 230
rect 756 180 790 198
rect 824 180 828 214
rect 722 160 828 180
rect 722 126 756 160
rect 790 146 828 160
rect 722 112 790 126
rect 824 112 828 146
rect 722 88 828 112
rect 862 103 932 368
rect 1003 398 1013 420
rect 1047 386 1060 420
rect 1037 370 1060 386
rect 1003 230 1037 364
rect 1122 230 1156 514
rect 1537 496 1579 530
rect 1613 496 1643 530
rect 1537 462 1643 496
rect 1537 448 1579 462
rect 1613 448 1643 462
rect 1571 428 1579 448
rect 1571 414 1609 428
rect 1703 504 1737 600
rect 1703 498 1809 504
rect 1737 464 1775 498
rect 1703 454 1775 464
rect 1703 420 1809 454
rect 966 214 1037 230
rect 1000 180 1037 214
rect 966 146 1037 180
rect 1076 214 1156 230
rect 1110 180 1156 214
rect 1076 164 1156 180
rect 1190 229 1224 324
rect 1000 112 1037 146
rect 722 54 756 88
rect 790 78 828 88
rect 722 44 790 54
rect 824 44 828 78
rect 722 28 828 44
rect 966 78 1037 112
rect 1000 44 1037 78
rect 1190 157 1224 195
rect 1190 68 1224 123
rect 1332 160 1366 180
rect 1332 88 1366 126
rect 966 28 1037 44
rect 1082 34 1106 68
rect 1140 34 1174 68
rect 1208 34 1232 68
rect 1485 160 1519 174
rect 1485 88 1519 106
rect 1485 22 1519 38
rect 1572 34 1606 414
rect 1703 386 1775 420
rect 1703 370 1809 386
rect 1851 482 1885 596
rect 2027 770 2379 782
rect 2027 766 2167 770
rect 2061 736 2167 766
rect 2201 736 2244 770
rect 2278 736 2321 770
rect 2355 736 2379 770
rect 2061 732 2379 736
rect 2027 706 2379 732
rect 2027 703 2237 706
rect 2027 698 2045 703
rect 2079 669 2117 703
rect 2151 669 2189 703
rect 2223 669 2237 703
rect 2061 664 2237 669
rect 2027 650 2237 664
rect 2027 630 2095 650
rect 2061 616 2095 630
rect 2129 616 2237 650
rect 2061 596 2237 616
rect 2027 580 2237 596
rect 2308 650 2393 666
rect 2308 616 2351 650
rect 2385 616 2393 650
rect 2308 600 2393 616
rect 2308 504 2342 600
rect 2529 506 2552 540
rect 2308 488 2365 504
rect 1851 448 2142 482
rect 2176 448 2210 482
rect 2244 448 2260 482
rect 2308 470 2318 488
rect 2352 454 2365 488
rect 1851 414 1869 448
rect 1903 414 1941 448
rect 2342 436 2365 454
rect 2308 420 2365 436
rect 1703 224 1737 370
rect 1851 242 1885 414
rect 2157 368 2195 402
rect 2308 398 2318 420
rect 2352 386 2365 420
rect 1661 208 1737 224
rect 1695 174 1737 208
rect 1661 140 1737 174
rect 1771 214 1885 242
rect 1805 180 1885 214
rect 1771 176 1885 180
rect 1925 318 2061 334
rect 1959 284 1997 318
rect 2031 300 2061 318
rect 2095 300 2119 334
rect 2031 284 2119 300
rect 1771 164 1805 176
rect 1695 106 1737 140
rect 1661 72 1737 106
rect 1695 38 1737 72
rect 1925 68 1987 284
rect 1661 22 1737 38
rect 1777 34 1801 68
rect 1835 34 1929 68
rect 1963 34 1987 68
rect 2027 214 2061 230
rect 2095 214 2133 230
rect 2061 180 2095 198
rect 2129 180 2133 214
rect 2027 160 2133 180
rect 2027 126 2061 160
rect 2095 146 2133 160
rect 2027 112 2095 126
rect 2129 112 2133 146
rect 2027 88 2133 112
rect 2027 54 2061 88
rect 2095 78 2133 88
rect 2027 44 2095 54
rect 2129 44 2133 78
rect 2167 73 2237 368
rect 2342 370 2365 386
rect 2495 468 2552 506
rect 2529 434 2552 468
rect 2495 396 2552 434
rect 2308 230 2342 364
rect 2271 214 2342 230
rect 2305 180 2342 214
rect 2271 146 2342 180
rect 2305 112 2342 146
rect 2271 78 2342 112
rect 2027 28 2133 44
rect 2305 44 2342 78
rect 2529 362 2552 396
rect 2495 324 2552 362
rect 2529 290 2552 324
rect 2495 68 2552 290
rect 2271 28 2342 44
<< viali >>
rect 241 677 275 711
rect 313 677 347 711
rect 232 414 266 448
rect 304 428 308 448
rect 308 428 338 448
rect 304 414 338 428
rect 398 464 432 498
rect 470 488 504 498
rect 470 464 504 488
rect 180 208 214 232
rect 180 198 214 208
rect 180 140 214 160
rect 180 126 214 140
rect 180 72 214 88
rect 180 54 214 72
rect 740 698 774 703
rect 740 669 756 698
rect 756 669 774 698
rect 812 669 846 703
rect 884 669 918 703
rect 1260 677 1294 711
rect 1332 698 1366 711
rect 1332 677 1366 698
rect 1546 677 1580 711
rect 1618 677 1652 711
rect 1128 514 1162 548
rect 1200 514 1234 548
rect 1003 454 1013 470
rect 1013 454 1037 470
rect 564 414 598 448
rect 636 414 670 448
rect 1003 436 1037 454
rect 787 368 821 402
rect 859 368 893 402
rect 620 284 654 318
rect 692 284 726 318
rect 756 198 790 232
rect 756 126 790 160
rect 1003 386 1013 398
rect 1013 386 1037 398
rect 1003 364 1037 386
rect 1537 414 1571 448
rect 1609 428 1613 448
rect 1613 428 1643 448
rect 1609 414 1643 428
rect 1703 464 1737 498
rect 1775 488 1809 498
rect 1775 464 1809 488
rect 1190 195 1224 229
rect 756 54 790 88
rect 1190 123 1224 157
rect 1332 214 1366 232
rect 1332 198 1366 214
rect 1332 126 1366 160
rect 1332 54 1366 88
rect 1485 208 1519 232
rect 1485 198 1519 208
rect 1485 140 1519 160
rect 1485 126 1519 140
rect 1485 72 1519 88
rect 1485 54 1519 72
rect 2045 698 2079 703
rect 2045 669 2061 698
rect 2061 669 2079 698
rect 2117 669 2151 703
rect 2189 669 2223 703
rect 2495 506 2529 540
rect 2308 454 2318 470
rect 2318 454 2342 470
rect 1869 414 1903 448
rect 1941 414 1975 448
rect 2308 436 2342 454
rect 2123 368 2157 402
rect 2195 368 2229 402
rect 2308 386 2318 398
rect 2318 386 2342 398
rect 1925 284 1959 318
rect 1997 284 2031 318
rect 2061 198 2095 232
rect 2061 126 2095 160
rect 2061 54 2095 88
rect 2308 364 2342 386
rect 2495 434 2529 468
rect 2495 362 2529 396
rect 2495 290 2529 324
<< metal1 >>
rect 235 711 2560 776
rect 235 677 241 711
rect 275 677 313 711
rect 347 703 1260 711
rect 347 677 740 703
rect 235 669 740 677
rect 774 669 812 703
rect 846 669 884 703
rect 918 677 1260 703
rect 1294 677 1332 711
rect 1366 677 1546 711
rect 1580 677 1618 711
rect 1652 703 2560 711
rect 1652 677 2045 703
rect 918 669 2045 677
rect 2079 669 2117 703
rect 2151 669 2189 703
rect 2223 669 2560 703
rect 235 588 2560 669
tri 1287 563 1312 588 ne
tri 253 548 265 560 se
rect 265 548 787 560
tri 245 540 253 548 se
rect 253 540 787 548
rect 245 532 787 540
rect 245 514 332 532
tri 332 514 350 532 nw
tri 552 514 570 532 ne
rect 570 514 664 532
tri 664 514 682 532 nw
tri 757 514 775 532 ne
rect 775 514 787 532
rect 245 509 327 514
tri 327 509 332 514 nw
tri 570 509 575 514 ne
rect 575 509 659 514
tri 659 509 664 514 nw
tri 775 509 780 514 ne
rect 780 509 787 514
rect 325 508 326 509
tri 326 508 327 509 nw
tri 575 508 576 509 ne
rect 576 508 577 509
rect 657 508 658 509
tri 658 508 659 509 nw
tri 780 508 781 509 ne
rect 781 508 787 509
rect 839 508 851 560
rect 903 510 1054 560
rect 1056 559 1084 560
rect 1055 511 1085 559
rect 1086 548 1240 560
rect 1086 514 1128 548
rect 1162 514 1200 548
rect 1234 520 1240 548
tri 1240 520 1248 528 sw
rect 1234 514 1248 520
rect 1056 510 1084 511
rect 1086 510 1248 514
rect 903 508 918 510
tri 918 508 920 510 nw
tri 1114 508 1116 510 ne
rect 1116 508 1248 510
rect 246 507 324 508
tri 325 507 326 508 nw
tri 576 507 577 508 ne
rect 578 507 656 508
tri 657 507 658 508 nw
tri 1116 507 1117 508 ne
rect 1117 507 1248 508
tri 1117 506 1118 507 ne
rect 1118 506 1248 507
tri 1248 506 1262 520 sw
tri 1118 504 1120 506 ne
rect 1120 504 1262 506
rect 386 498 516 504
tri 1120 502 1122 504 ne
rect 1122 502 1262 504
tri 1200 498 1204 502 ne
rect 1204 498 1262 502
tri 1262 498 1270 506 sw
rect 1312 500 1386 588
rect 1444 508 1450 560
rect 1502 508 1514 560
rect 1566 532 1962 560
rect 1566 508 1572 532
tri 1860 510 1882 532 ne
rect 1882 509 1962 532
rect 1883 507 1961 508
rect 2489 540 2535 552
rect 2489 506 2495 540
rect 2529 506 2535 540
rect 1691 498 1821 504
tri 230 464 245 479 se
rect 246 478 324 479
tri 325 478 326 479 sw
rect 325 477 326 478
tri 326 477 327 478 sw
rect 245 464 327 477
tri 327 464 340 477 sw
rect 386 464 398 498
rect 432 464 470 498
rect 504 464 516 498
tri 1204 482 1220 498 ne
rect 1220 482 1270 498
tri 995 480 997 482 se
rect 997 480 1043 482
tri 1220 480 1222 482 ne
rect 1222 480 1270 482
tri 1270 480 1288 498 sw
tri 568 470 577 479 se
rect 578 478 656 479
tri 657 478 658 479 sw
rect 657 477 658 478
tri 658 477 659 478 sw
rect 577 470 659 477
tri 659 470 666 477 sw
tri 220 454 230 464 se
rect 230 454 340 464
tri 340 454 350 464 sw
rect 386 458 516 464
tri 556 458 568 470 se
rect 568 458 666 470
tri 386 454 390 458 ne
rect 390 454 512 458
tri 512 454 516 458 nw
tri 552 454 556 458 se
rect 556 454 666 458
tri 666 454 682 470 sw
rect 220 448 350 454
tri 390 448 396 454 ne
rect 396 448 506 454
tri 506 448 512 454 nw
rect 552 448 682 454
rect 220 414 232 448
rect 266 414 304 448
rect 338 414 350 448
tri 396 433 411 448 ne
rect 411 435 493 448
tri 493 435 506 448 nw
rect 491 434 492 435
tri 492 434 493 435 nw
rect 412 433 490 434
tri 491 433 492 434 nw
rect 220 408 350 414
rect 552 414 564 448
rect 598 414 636 448
rect 670 414 682 448
rect 775 414 936 480
rect 938 479 966 480
rect 552 408 682 414
tri 772 405 774 407 se
rect 774 405 780 414
tri 408 402 411 405 se
rect 412 404 490 405
tri 491 404 492 405 sw
tri 771 404 772 405 se
rect 772 404 780 405
rect 491 403 492 404
tri 492 403 493 404 sw
tri 770 403 771 404 se
rect 771 403 780 404
rect 411 402 493 403
tri 493 402 494 403 sw
tri 769 402 770 403 se
rect 770 402 780 403
tri 386 380 408 402 se
rect 408 380 494 402
tri 494 380 516 402 sw
tri 747 380 769 402 se
rect 769 380 780 402
rect 386 362 780 380
rect 832 362 844 414
rect 896 362 936 414
rect 386 352 936 362
rect 937 353 967 479
rect 968 470 1043 480
rect 968 436 1003 470
rect 1037 436 1043 470
tri 1222 464 1238 480 ne
rect 1238 464 1288 480
tri 1288 464 1304 480 sw
rect 1691 464 1703 498
rect 1737 464 1775 498
rect 1809 464 1821 498
tri 1873 470 1882 479 se
rect 1883 478 1961 479
tri 1962 478 1963 479 sw
rect 1962 477 1963 478
tri 1963 477 1964 478 sw
rect 1882 470 1964 477
tri 1964 470 1971 477 sw
rect 2302 470 2348 482
tri 1238 454 1248 464 ne
rect 1248 454 1304 464
tri 1304 454 1314 464 sw
rect 1691 458 1821 464
tri 1861 458 1873 470 se
rect 1873 458 1971 470
tri 1691 454 1695 458 ne
rect 1695 454 1817 458
tri 1817 454 1821 458 nw
tri 1857 454 1861 458 se
rect 1861 454 1971 458
tri 1971 454 1987 470 sw
tri 1248 448 1254 454 ne
rect 1254 448 1655 454
tri 1695 448 1701 454 ne
rect 1701 448 1811 454
tri 1811 448 1817 454 nw
rect 1857 448 1987 454
rect 968 398 1043 436
tri 1254 414 1288 448 ne
rect 1288 414 1537 448
rect 1571 414 1609 448
rect 1643 414 1655 448
tri 1701 433 1716 448 ne
rect 1716 435 1798 448
tri 1798 435 1811 448 nw
rect 1796 434 1797 435
tri 1797 434 1798 435 nw
rect 1717 433 1795 434
tri 1796 433 1797 434 nw
tri 1288 408 1294 414 ne
rect 1294 408 1655 414
rect 1857 414 1869 448
rect 1903 414 1941 448
rect 1975 414 1987 448
rect 2302 436 2308 470
rect 2342 436 2348 470
tri 2283 414 2302 433 se
rect 2302 414 2348 436
rect 1857 408 1987 414
tri 2028 408 2034 414 se
rect 2034 408 2040 414
tri 2025 405 2028 408 se
rect 2028 405 2040 408
rect 968 364 1003 398
rect 1037 364 1043 398
rect 938 352 966 353
rect 968 352 1043 364
rect 1717 404 1795 405
tri 1796 404 1797 405 sw
tri 2024 404 2025 405 se
rect 2025 404 2040 405
rect 1796 403 1797 404
tri 1797 403 1798 404 sw
tri 2023 403 2024 404 se
rect 2024 403 2040 404
rect 1716 402 1798 403
tri 1798 402 1799 403 sw
tri 2022 402 2023 403 se
rect 2023 402 2040 403
rect 1716 380 1799 402
tri 1799 380 1821 402 sw
tri 2000 380 2022 402 se
rect 2022 380 2040 402
rect 1716 362 2040 380
rect 2092 362 2104 414
rect 2156 408 2162 414
tri 2277 408 2283 414 se
rect 2283 408 2348 414
rect 2156 402 2241 408
rect 2157 368 2195 402
rect 2229 368 2241 402
rect 2156 362 2241 368
rect 1716 352 2241 362
rect 2242 353 2243 407
rect 2271 353 2272 407
rect 2273 398 2348 408
rect 2273 364 2308 398
rect 2342 364 2348 398
rect 2273 352 2348 364
rect 2489 468 2535 506
rect 2489 434 2495 468
rect 2529 434 2535 468
rect 2489 396 2535 434
rect 2489 362 2495 396
rect 2529 362 2535 396
tri 2464 324 2489 349 se
rect 2489 324 2535 362
rect 220 318 1386 324
rect 220 284 620 318
rect 654 284 692 318
rect 726 284 1386 318
rect 220 278 1386 284
rect 1525 318 2495 324
rect 1525 284 1925 318
rect 1959 284 1997 318
rect 2031 290 2495 318
rect 2529 290 2535 324
rect 2031 284 2535 290
rect 1525 278 2535 284
rect 88 232 1386 250
rect 88 198 180 232
rect 214 198 756 232
rect 790 229 1332 232
rect 790 198 1190 229
rect 88 195 1190 198
rect 1224 198 1332 229
rect 1366 198 1386 232
rect 1224 195 1386 198
rect 88 160 1386 195
rect 88 126 180 160
rect 214 126 756 160
rect 790 157 1332 160
rect 790 126 1190 157
rect 88 123 1190 126
rect 1224 126 1332 157
rect 1366 126 1386 160
rect 1224 123 1386 126
rect 88 88 1386 123
rect 88 54 180 88
rect 214 54 756 88
rect 790 54 1332 88
rect 1366 54 1386 88
rect 88 48 1386 54
rect 1393 232 2560 250
rect 1393 198 1485 232
rect 1519 198 2061 232
rect 2095 198 2560 232
rect 1393 160 2560 198
rect 1393 126 1485 160
rect 1519 126 2061 160
rect 2095 126 2560 160
rect 1393 88 2560 126
rect 1393 54 1485 88
rect 1519 54 2061 88
rect 2095 54 2560 88
rect 1393 48 2560 54
<< rmetal1 >>
rect 245 508 325 509
rect 577 508 657 509
rect 1054 559 1056 560
rect 1084 559 1086 560
rect 1054 511 1055 559
rect 1085 511 1086 559
rect 1054 510 1056 511
rect 1084 510 1086 511
rect 245 507 246 508
rect 324 507 325 508
rect 577 507 578 508
rect 656 507 657 508
rect 1882 508 1962 509
rect 1882 507 1883 508
rect 1961 507 1962 508
rect 245 478 246 479
rect 324 478 325 479
rect 245 477 325 478
rect 577 478 578 479
rect 656 478 657 479
rect 577 477 657 478
rect 411 434 491 435
rect 411 433 412 434
rect 490 433 491 434
rect 936 479 938 480
rect 966 479 968 480
rect 411 404 412 405
rect 490 404 491 405
rect 411 403 491 404
rect 936 353 937 479
rect 967 353 968 479
rect 1882 478 1883 479
rect 1961 478 1962 479
rect 1882 477 1962 478
rect 1716 434 1796 435
rect 1716 433 1717 434
rect 1795 433 1796 434
rect 936 352 938 353
rect 966 352 968 353
rect 1716 404 1717 405
rect 1795 404 1796 405
rect 1716 403 1796 404
rect 2241 407 2243 408
rect 2241 353 2242 407
rect 2241 352 2243 353
rect 2271 407 2273 408
rect 2272 353 2273 407
rect 2271 352 2273 353
<< via1 >>
rect 787 508 839 560
rect 851 508 903 560
rect 1450 508 1502 560
rect 1514 508 1566 560
rect 780 402 832 414
rect 780 368 787 402
rect 787 368 821 402
rect 821 368 832 402
rect 780 362 832 368
rect 844 402 896 414
rect 844 368 859 402
rect 859 368 893 402
rect 893 368 896 402
rect 844 362 896 368
rect 2040 362 2092 414
rect 2104 402 2156 414
rect 2104 368 2123 402
rect 2123 368 2156 402
rect 2104 362 2156 368
<< metal2 >>
rect 781 508 787 560
rect 839 508 851 560
rect 903 508 1450 560
rect 1502 508 1514 560
rect 1566 508 1572 560
rect 774 362 780 414
rect 832 362 844 414
rect 896 362 2040 414
rect 2092 362 2104 414
rect 2156 362 2162 414
use sky130_fd_io__tk_em1o_b_cdns_55959141808131  sky130_fd_io__tk_em1o_b_cdns_55959141808131_0
timestamp 1649977179
transform 1 0 2189 0 -1 408
box 21 24 115 28
use sky130_fd_io__tk_em1o_b_cdns_55959141808132  sky130_fd_io__tk_em1o_b_cdns_55959141808132_0
timestamp 1649977179
transform 0 -1 1796 1 0 351
box 21 24 115 28
use sky130_fd_io__tk_em1o_b_cdns_55959141808132  sky130_fd_io__tk_em1o_b_cdns_55959141808132_1
timestamp 1649977179
transform 0 -1 1962 1 0 425
box 21 24 115 28
use sky130_fd_io__tk_em1o_b_cdns_55959141808132  sky130_fd_io__tk_em1o_b_cdns_55959141808132_2
timestamp 1649977179
transform 0 -1 657 1 0 425
box 21 24 115 28
use sky130_fd_io__tk_em1o_b_cdns_55959141808132  sky130_fd_io__tk_em1o_b_cdns_55959141808132_3
timestamp 1649977179
transform 0 -1 491 1 0 351
box 21 24 115 28
use sky130_fd_io__tk_em1o_b_cdns_55959141808132  sky130_fd_io__tk_em1o_b_cdns_55959141808132_4
timestamp 1649977179
transform 0 -1 325 1 0 425
box 21 24 115 28
use sky130_fd_io__tk_em1s_b_cdns_55959141808129  sky130_fd_io__tk_em1s_b_cdns_55959141808129_0
timestamp 1649977179
transform -1 0 1138 0 -1 560
box 24 24 110 28
use sky130_fd_io__tk_em1s_b_cdns_55959141808130  sky130_fd_io__tk_em1s_b_cdns_55959141808130_0
timestamp 1649977179
transform 1 0 884 0 -1 480
box 21 24 113 28
use sky130_fd_pr__nfet_01v8__example_55959141808133  sky130_fd_pr__nfet_01v8__example_55959141808133_0
timestamp 1649977179
transform -1 0 2016 0 -1 226
box -28 0 228 29
use sky130_fd_pr__nfet_01v8__example_55959141808133  sky130_fd_pr__nfet_01v8__example_55959141808133_1
timestamp 1649977179
transform -1 0 1321 0 -1 226
box -28 0 228 29
use sky130_fd_pr__nfet_01v8__example_55959141808133  sky130_fd_pr__nfet_01v8__example_55959141808133_2
timestamp 1649977179
transform -1 0 711 0 -1 226
box -28 0 228 29
use sky130_fd_pr__nfet_01v8__example_55959141808134  sky130_fd_pr__nfet_01v8__example_55959141808134_0
timestamp 1649977179
transform 1 0 1530 0 1 26
box -28 0 148 97
use sky130_fd_pr__nfet_01v8__example_55959141808134  sky130_fd_pr__nfet_01v8__example_55959141808134_1
timestamp 1649977179
transform 1 0 2140 0 -1 226
box -28 0 148 97
use sky130_fd_pr__nfet_01v8__example_55959141808134  sky130_fd_pr__nfet_01v8__example_55959141808134_2
timestamp 1649977179
transform 1 0 835 0 -1 226
box -28 0 148 97
use sky130_fd_pr__nfet_01v8__example_55959141808134  sky130_fd_pr__nfet_01v8__example_55959141808134_3
timestamp 1649977179
transform 1 0 225 0 1 26
box -28 0 148 97
use sky130_fd_pr__pfet_01v8__example_55959141808135  sky130_fd_pr__pfet_01v8__example_55959141808135_0
timestamp 1649977179
transform 1 0 1530 0 -1 662
box -28 0 228 29
use sky130_fd_pr__pfet_01v8__example_55959141808135  sky130_fd_pr__pfet_01v8__example_55959141808135_1
timestamp 1649977179
transform 1 0 225 0 -1 662
box -28 0 228 29
use sky130_fd_pr__pfet_01v8__example_55959141808136  sky130_fd_pr__pfet_01v8__example_55959141808136_0
timestamp 1649977179
transform -1 0 2016 0 -1 778
box -28 0 148 97
use sky130_fd_pr__pfet_01v8__example_55959141808136  sky130_fd_pr__pfet_01v8__example_55959141808136_1
timestamp 1649977179
transform -1 0 1321 0 -1 778
box -28 0 148 97
use sky130_fd_pr__pfet_01v8__example_55959141808136  sky130_fd_pr__pfet_01v8__example_55959141808136_2
timestamp 1649977179
transform -1 0 711 0 -1 778
box -28 0 148 97
use sky130_fd_pr__pfet_01v8__example_55959141808138  sky130_fd_pr__pfet_01v8__example_55959141808138_0
timestamp 1649977179
transform 1 0 2140 0 -1 662
box -28 0 228 29
use sky130_fd_pr__pfet_01v8__example_55959141808138  sky130_fd_pr__pfet_01v8__example_55959141808138_1
timestamp 1649977179
transform 1 0 835 0 -1 662
box -28 0 228 29
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_0
timestamp 1649977179
transform 0 -1 2342 -1 0 470
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_1
timestamp 1649977179
transform -1 0 1809 0 1 464
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_2
timestamp 1649977179
transform -1 0 1643 0 1 414
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_3
timestamp 1649977179
transform -1 0 1975 0 1 414
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_4
timestamp 1649977179
transform -1 0 2229 0 1 368
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_5
timestamp 1649977179
transform -1 0 2031 0 1 284
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_6
timestamp 1649977179
transform -1 0 726 0 1 284
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_7
timestamp 1649977179
transform 0 -1 1224 -1 0 229
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_8
timestamp 1649977179
transform -1 0 893 0 1 368
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_9
timestamp 1649977179
transform -1 0 670 0 1 414
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_10
timestamp 1649977179
transform -1 0 338 0 1 414
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_11
timestamp 1649977179
transform -1 0 504 0 1 464
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_12
timestamp 1649977179
transform 0 -1 1037 -1 0 470
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_5595914180878  sky130_fd_pr__via_l1m1__example_5595914180878_0
timestamp 1649977179
transform 0 -1 1652 1 0 677
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_5595914180878  sky130_fd_pr__via_l1m1__example_5595914180878_1
timestamp 1649977179
transform 0 -1 1234 1 0 514
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_5595914180878  sky130_fd_pr__via_l1m1__example_5595914180878_2
timestamp 1649977179
transform 0 1 1260 1 0 677
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_5595914180878  sky130_fd_pr__via_l1m1__example_5595914180878_3
timestamp 1649977179
transform 0 -1 347 1 0 677
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_55959141808127  sky130_fd_pr__via_l1m1__example_55959141808127_0
timestamp 1649977179
transform 0 -1 2529 1 0 290
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_55959141808128  sky130_fd_pr__via_l1m1__example_55959141808128_0
timestamp 1649977179
transform -1 0 2095 0 1 54
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_55959141808128  sky130_fd_pr__via_l1m1__example_55959141808128_1
timestamp 1649977179
transform -1 0 1519 0 1 54
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_55959141808128  sky130_fd_pr__via_l1m1__example_55959141808128_2
timestamp 1649977179
transform 0 -1 2223 1 0 669
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_55959141808128  sky130_fd_pr__via_l1m1__example_55959141808128_3
timestamp 1649977179
transform 0 -1 918 1 0 669
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_55959141808128  sky130_fd_pr__via_l1m1__example_55959141808128_4
timestamp 1649977179
transform -1 0 214 0 1 54
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_55959141808128  sky130_fd_pr__via_l1m1__example_55959141808128_5
timestamp 1649977179
transform -1 0 790 0 1 54
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_55959141808128  sky130_fd_pr__via_l1m1__example_55959141808128_6
timestamp 1649977179
transform -1 0 1366 0 1 54
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_559591418083  sky130_fd_pr__via_pol1__example_559591418083_0
timestamp 1649977179
transform 0 -1 1629 -1 0 546
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_559591418083  sky130_fd_pr__via_pol1__example_559591418083_1
timestamp 1649977179
transform 0 -1 324 -1 0 546
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_5595914180833  sky130_fd_pr__via_pol1__example_5595914180833_0
timestamp 1649977179
transform 1 0 1759 0 1 370
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_5595914180833  sky130_fd_pr__via_pol1__example_5595914180833_1
timestamp 1649977179
transform 0 1 2126 1 0 432
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_5595914180833  sky130_fd_pr__via_pol1__example_5595914180833_2
timestamp 1649977179
transform 1 0 2302 0 1 370
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_5595914180833  sky130_fd_pr__via_pol1__example_5595914180833_3
timestamp 1649977179
transform 1 0 997 0 1 370
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_5595914180833  sky130_fd_pr__via_pol1__example_5595914180833_4
timestamp 1649977179
transform 0 1 821 1 0 432
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_5595914180833  sky130_fd_pr__via_pol1__example_5595914180833_5
timestamp 1649977179
transform 1 0 454 0 1 370
box 0 0 1 1
<< labels >>
flabel locali s 267 34 301 48 0 FreeSans 200 0 0 0 IN
port 1 nsew
flabel locali s 1021 337 1021 337 0 FreeSans 200 0 0 0 A3
port 2 nsew
flabel locali s 414 337 414 337 0 FreeSans 200 0 0 0 A1
port 3 nsew
flabel locali s 735 465 735 465 0 FreeSans 200 0 0 0 A2
port 4 nsew
flabel locali s 2326 337 2326 337 0 FreeSans 200 0 0 0 A7
port 5 nsew
flabel locali s 1719 337 1719 337 0 FreeSans 200 0 0 0 A5
port 6 nsew
flabel locali s 2040 465 2040 465 0 FreeSans 200 0 0 0 A6
port 7 nsew
flabel metal1 s 517 361 551 375 0 FreeSans 200 0 0 0 OUT_N
port 8 nsew
flabel metal1 s 517 541 551 555 0 FreeSans 200 0 0 0 OUT
port 9 nsew
flabel metal1 s 1366 48 1386 250 0 FreeSans 200 0 0 0 VGND
port 10 nsew
flabel metal1 s 1366 278 1386 324 0 FreeSans 200 0 0 0 VGND
port 10 nsew
flabel metal1 s 235 588 264 776 0 FreeSans 200 0 0 0 VCC_IO
port 11 nsew
flabel metal1 s 1360 500 1386 776 0 FreeSans 200 0 0 0 VCC_IO
port 11 nsew
flabel metal1 s 220 278 250 324 0 FreeSans 200 0 0 0 VGND
port 10 nsew
<< properties >>
string GDS_END 39982008
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 39965082
<< end >>
