magic
tech sky130A
magscale 1 2
timestamp 1649977179
use sky130_fd_pr__hvdfm1sd2__example_55959141808719  sky130_fd_pr__hvdfm1sd2__example_55959141808719_0
timestamp 1649977179
transform -1 0 0 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfm1sd2__example_55959141808719  sky130_fd_pr__hvdfm1sd2__example_55959141808719_1
timestamp 1649977179
transform 1 0 200 0 1 0
box 0 0 1 1
<< labels >>
flabel comment s 228 265 228 265 0 FreeSans 300 0 0 0 D
flabel comment s -28 265 -28 265 0 FreeSans 300 0 0 0 S
<< properties >>
string GDS_END 31290532
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 31289474
<< end >>
