magic
tech sky130B
magscale 1 2
timestamp 1649977179
<< nwell >>
rect -38 261 2522 582
<< pwell >>
rect 1 201 610 203
rect 1019 201 2480 203
rect 1 23 2480 201
rect 1 21 1106 23
rect 2192 21 2480 23
rect 29 -17 63 21
<< locali >>
rect 190 215 288 255
rect 1895 215 1973 265
rect 1938 187 1973 215
rect 1938 147 2002 187
rect 2174 299 2278 493
rect 2397 357 2467 493
rect 2174 165 2208 299
rect 2422 165 2467 357
rect 2174 54 2262 165
rect 2396 51 2467 165
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2053 561
rect 2087 527 2145 561
rect 2179 527 2237 561
rect 2271 527 2329 561
rect 2363 527 2421 561
rect 2455 527 2484 561
rect 17 413 79 493
rect 113 452 186 527
rect 413 447 479 527
rect 527 459 990 493
rect 1025 459 1512 493
rect 527 413 561 459
rect 17 379 561 413
rect 606 391 864 425
rect 17 300 89 379
rect 197 323 263 343
rect 17 161 51 300
rect 123 291 263 323
rect 122 289 263 291
rect 298 300 368 345
rect 298 289 364 300
rect 122 276 163 289
rect 122 265 156 276
rect 85 199 156 265
rect 119 181 156 199
rect 323 181 364 289
rect 403 282 438 345
rect 472 289 572 343
rect 398 255 438 282
rect 432 221 499 255
rect 398 215 499 221
rect 17 51 85 161
rect 119 147 264 181
rect 119 17 153 109
rect 198 51 264 147
rect 300 177 364 181
rect 300 143 504 177
rect 300 51 368 143
rect 402 17 436 109
rect 470 85 504 143
rect 538 119 572 289
rect 606 93 640 391
rect 797 357 864 391
rect 674 291 763 357
rect 674 161 708 291
rect 814 232 907 323
rect 814 215 880 232
rect 941 185 975 459
rect 1025 264 1059 459
rect 1095 340 1175 406
rect 1258 391 1444 425
rect 1258 323 1292 391
rect 1221 289 1292 323
rect 1025 230 1101 264
rect 1064 185 1101 230
rect 1135 255 1185 265
rect 1342 255 1376 357
rect 1135 221 1136 255
rect 1170 221 1185 255
rect 1135 199 1185 221
rect 896 181 1029 185
rect 814 161 1029 181
rect 1064 173 1104 185
rect 1067 168 1104 173
rect 674 127 780 161
rect 814 156 1031 161
rect 814 151 1034 156
rect 814 147 912 151
rect 985 148 1034 151
rect 985 147 1036 148
rect 814 129 880 147
rect 990 143 1036 147
rect 996 138 1036 143
rect 1000 131 1036 138
rect 930 93 968 117
rect 606 85 968 93
rect 470 51 968 85
rect 1002 85 1036 131
rect 1070 119 1104 168
rect 1221 148 1287 255
rect 1322 185 1376 255
rect 1410 235 1444 391
rect 1478 285 1512 459
rect 1546 459 1931 493
rect 1546 302 1592 459
rect 1629 391 1850 425
rect 1478 280 1515 285
rect 1478 275 1519 280
rect 1478 255 1524 275
rect 1410 226 1449 235
rect 1410 212 1456 226
rect 1413 209 1456 212
rect 1418 202 1456 209
rect 1322 151 1388 185
rect 1354 119 1388 151
rect 1422 153 1456 202
rect 1490 199 1524 255
rect 1558 165 1592 302
rect 1645 289 1782 357
rect 1645 185 1681 289
rect 1816 255 1850 391
rect 1884 341 1931 459
rect 1968 455 2035 527
rect 2069 375 2138 493
rect 1884 299 2070 341
rect 1422 119 1489 153
rect 1150 85 1220 113
rect 1002 51 1220 85
rect 1254 85 1320 114
rect 1541 85 1592 165
rect 1631 119 1681 185
rect 1715 221 1850 255
rect 1715 119 1749 221
rect 2036 199 2070 299
rect 1784 137 1860 187
rect 2104 165 2138 375
rect 1880 85 1947 103
rect 1254 51 1947 85
rect 1981 17 2015 113
rect 2049 57 2138 165
rect 2312 357 2363 527
rect 2242 199 2292 265
rect 2326 199 2388 323
rect 2296 17 2362 165
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2053 17
rect 2087 -17 2145 17
rect 2179 -17 2237 17
rect 2271 -17 2329 17
rect 2363 -17 2421 17
rect 2455 -17 2484 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 1593 527 1627 561
rect 1685 527 1719 561
rect 1777 527 1811 561
rect 1869 527 1903 561
rect 1961 527 1995 561
rect 2053 527 2087 561
rect 2145 527 2179 561
rect 2237 527 2271 561
rect 2329 527 2363 561
rect 2421 527 2455 561
rect 398 221 432 255
rect 1136 221 1170 255
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1593 -17 1627 17
rect 1685 -17 1719 17
rect 1777 -17 1811 17
rect 1869 -17 1903 17
rect 1961 -17 1995 17
rect 2053 -17 2087 17
rect 2145 -17 2179 17
rect 2237 -17 2271 17
rect 2329 -17 2363 17
rect 2421 -17 2455 17
<< metal1 >>
rect 0 561 2484 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2053 561
rect 2087 527 2145 561
rect 2179 527 2237 561
rect 2271 527 2329 561
rect 2363 527 2421 561
rect 2455 527 2484 561
rect 0 496 2484 527
rect 386 255 444 261
rect 386 221 398 255
rect 432 252 444 255
rect 1124 255 1182 261
rect 1124 252 1136 255
rect 432 224 1136 252
rect 432 221 444 224
rect 386 215 444 221
rect 1124 221 1136 224
rect 1170 221 1182 255
rect 1124 215 1182 221
rect 0 17 2484 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2053 17
rect 2087 -17 2145 17
rect 2179 -17 2237 17
rect 2271 -17 2329 17
rect 2363 -17 2421 17
rect 2455 -17 2484 17
rect 0 -48 2484 -17
<< obsm1 >>
rect 785 388 843 397
rect 1102 388 1160 397
rect 785 360 1160 388
rect 785 351 843 360
rect 1102 351 1160 360
rect 1804 388 1862 397
rect 2092 388 2150 397
rect 1804 360 2150 388
rect 1804 351 1862 360
rect 2092 351 2150 360
rect 478 320 536 329
rect 861 320 919 329
rect 1218 320 1276 329
rect 478 292 1276 320
rect 478 283 536 292
rect 861 283 919 292
rect 1218 283 1276 292
rect 1680 320 1738 329
rect 2324 320 2382 329
rect 1680 292 2382 320
rect 1680 283 1738 292
rect 2324 283 2382 292
rect 1310 252 1368 261
rect 2232 252 2290 261
rect 1310 224 2290 252
rect 1310 215 1368 224
rect 2232 215 2290 224
rect 662 184 720 193
rect 1218 184 1276 193
rect 1772 184 1830 193
rect 662 156 1830 184
rect 662 147 720 156
rect 1218 147 1276 156
rect 1772 147 1830 156
<< labels >>
rlabel locali s 190 215 288 255 6 A
port 1 nsew signal input
rlabel metal1 s 1124 215 1182 224 6 B
port 2 nsew signal input
rlabel metal1 s 386 215 444 224 6 B
port 2 nsew signal input
rlabel metal1 s 386 224 1182 252 6 B
port 2 nsew signal input
rlabel metal1 s 1124 252 1182 261 6 B
port 2 nsew signal input
rlabel metal1 s 386 252 444 261 6 B
port 2 nsew signal input
rlabel locali s 1938 147 2002 187 6 CI
port 3 nsew signal input
rlabel locali s 1938 187 1973 215 6 CI
port 3 nsew signal input
rlabel locali s 1895 215 1973 265 6 CI
port 3 nsew signal input
rlabel metal1 s 0 -48 2484 48 8 VGND
port 4 nsew ground bidirectional abutment
rlabel pwell s 29 -17 63 21 6 VNB
port 5 nsew ground bidirectional
rlabel pwell s 2192 21 2480 23 6 VNB
port 5 nsew ground bidirectional
rlabel pwell s 1 21 1106 23 6 VNB
port 5 nsew ground bidirectional
rlabel pwell s 1 23 2480 201 6 VNB
port 5 nsew ground bidirectional
rlabel pwell s 1019 201 2480 203 6 VNB
port 5 nsew ground bidirectional
rlabel pwell s 1 201 610 203 6 VNB
port 5 nsew ground bidirectional
rlabel nwell s -38 261 2522 582 6 VPB
port 6 nsew power bidirectional
rlabel metal1 s 0 496 2484 592 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 2174 54 2262 165 6 COUT
port 8 nsew signal output
rlabel locali s 2174 165 2208 299 6 COUT
port 8 nsew signal output
rlabel locali s 2174 299 2278 493 6 COUT
port 8 nsew signal output
rlabel locali s 2396 51 2467 165 6 SUM
port 9 nsew signal output
rlabel locali s 2422 165 2467 357 6 SUM
port 9 nsew signal output
rlabel locali s 2397 357 2467 493 6 SUM
port 9 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 2484 544
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_END 2113468
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 2094028
<< end >>
