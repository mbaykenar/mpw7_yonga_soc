magic
tech sky130B
magscale 12 1
timestamp 1598768087
<< metal5 >>
rect 0 100 35 105
rect 0 95 40 100
rect 0 85 45 95
rect 0 50 15 85
rect 30 50 45 85
rect 0 40 45 50
rect 0 35 40 40
rect 0 30 35 35
rect 0 0 15 30
<< properties >>
string FIXED_BBOX 0 -30 60 105
<< end >>
