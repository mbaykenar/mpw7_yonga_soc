magic
tech sky130B
magscale 12 1
timestamp 1598777367
<< metal5 >>
rect 15 75 30 90
rect 0 60 45 75
rect 15 0 30 60
<< properties >>
string FIXED_BBOX 0 -30 60 105
<< end >>
