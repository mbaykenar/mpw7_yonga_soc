magic
tech sky130A
magscale 1 2
timestamp 1649977179
use sky130_fd_pr__dfl1sd2__example_5595914180884  sky130_fd_pr__dfl1sd2__example_5595914180884_0
timestamp 1649977179
transform 1 0 120 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfl1sd__example_5595914180819  sky130_fd_pr__dfl1sd__example_5595914180819_0
timestamp 1649977179
transform -1 0 0 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfl1sd__example_5595914180819  sky130_fd_pr__dfl1sd__example_5595914180819_1
timestamp 1649977179
transform 1 0 296 0 1 0
box 0 0 1 1
<< labels >>
flabel comment s 324 267 324 267 0 FreeSans 300 0 0 0 D
flabel comment s 148 267 148 267 0 FreeSans 300 0 0 0 S
flabel comment s -28 267 -28 267 0 FreeSans 300 0 0 0 D
<< properties >>
string GDS_END 7449828
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 7448392
<< end >>
