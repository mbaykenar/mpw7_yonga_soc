module user_project_wrapper (user_clock2,
    vccd1,
    vccd2,
    vdda1,
    vdda2,
    vssa1,
    vssa2,
    vssd1,
    vssd2,
    wb_clk_i,
    wb_rst_i,
    wbs_ack_o,
    wbs_cyc_i,
    wbs_stb_i,
    wbs_we_i,
    analog_io,
    io_in,
    io_oeb,
    io_out,
    la_data_in,
    la_data_out,
    la_oenb,
    user_irq,
    wbs_adr_i,
    wbs_dat_i,
    wbs_dat_o,
    wbs_sel_i);
 input user_clock2;
 input vccd1;
 input vccd2;
 input vdda1;
 input vdda2;
 input vssa1;
 input vssa2;
 input vssd1;
 input vssd2;
 input wb_clk_i;
 input wb_rst_i;
 output wbs_ack_o;
 input wbs_cyc_i;
 input wbs_stb_i;
 input wbs_we_i;
 inout [28:0] analog_io;
 input [37:0] io_in;
 output [37:0] io_oeb;
 output [37:0] io_out;
 input [127:0] la_data_in;
 output [127:0] la_data_out;
 input [127:0] la_oenb;
 output [2:0] user_irq;
 input [31:0] wbs_adr_i;
 input [31:0] wbs_dat_i;
 output [31:0] wbs_dat_o;
 input [3:0] wbs_sel_i;

 wire \boot_addr_int[0] ;
 wire \boot_addr_int[10] ;
 wire \boot_addr_int[11] ;
 wire \boot_addr_int[12] ;
 wire \boot_addr_int[13] ;
 wire \boot_addr_int[14] ;
 wire \boot_addr_int[15] ;
 wire \boot_addr_int[16] ;
 wire \boot_addr_int[17] ;
 wire \boot_addr_int[18] ;
 wire \boot_addr_int[19] ;
 wire \boot_addr_int[1] ;
 wire \boot_addr_int[20] ;
 wire \boot_addr_int[21] ;
 wire \boot_addr_int[22] ;
 wire \boot_addr_int[23] ;
 wire \boot_addr_int[24] ;
 wire \boot_addr_int[25] ;
 wire \boot_addr_int[26] ;
 wire \boot_addr_int[27] ;
 wire \boot_addr_int[28] ;
 wire \boot_addr_int[29] ;
 wire \boot_addr_int[2] ;
 wire \boot_addr_int[30] ;
 wire \boot_addr_int[31] ;
 wire \boot_addr_int[3] ;
 wire \boot_addr_int[4] ;
 wire \boot_addr_int[5] ;
 wire \boot_addr_int[6] ;
 wire \boot_addr_int[7] ;
 wire \boot_addr_int[8] ;
 wire \boot_addr_int[9] ;
 wire cfgack_fll_int;
 wire \cfgad_fll_int[0] ;
 wire \cfgad_fll_int[1] ;
 wire \cfgd_fll_int[0] ;
 wire \cfgd_fll_int[10] ;
 wire \cfgd_fll_int[11] ;
 wire \cfgd_fll_int[12] ;
 wire \cfgd_fll_int[13] ;
 wire \cfgd_fll_int[14] ;
 wire \cfgd_fll_int[15] ;
 wire \cfgd_fll_int[16] ;
 wire \cfgd_fll_int[17] ;
 wire \cfgd_fll_int[18] ;
 wire \cfgd_fll_int[19] ;
 wire \cfgd_fll_int[1] ;
 wire \cfgd_fll_int[20] ;
 wire \cfgd_fll_int[21] ;
 wire \cfgd_fll_int[22] ;
 wire \cfgd_fll_int[23] ;
 wire \cfgd_fll_int[24] ;
 wire \cfgd_fll_int[25] ;
 wire \cfgd_fll_int[26] ;
 wire \cfgd_fll_int[27] ;
 wire \cfgd_fll_int[28] ;
 wire \cfgd_fll_int[29] ;
 wire \cfgd_fll_int[2] ;
 wire \cfgd_fll_int[30] ;
 wire \cfgd_fll_int[31] ;
 wire \cfgd_fll_int[3] ;
 wire \cfgd_fll_int[4] ;
 wire \cfgd_fll_int[5] ;
 wire \cfgd_fll_int[6] ;
 wire \cfgd_fll_int[7] ;
 wire \cfgd_fll_int[8] ;
 wire \cfgd_fll_int[9] ;
 wire \cfgq_fll_int[0] ;
 wire \cfgq_fll_int[10] ;
 wire \cfgq_fll_int[11] ;
 wire \cfgq_fll_int[12] ;
 wire \cfgq_fll_int[13] ;
 wire \cfgq_fll_int[14] ;
 wire \cfgq_fll_int[15] ;
 wire \cfgq_fll_int[16] ;
 wire \cfgq_fll_int[17] ;
 wire \cfgq_fll_int[18] ;
 wire \cfgq_fll_int[19] ;
 wire \cfgq_fll_int[1] ;
 wire \cfgq_fll_int[20] ;
 wire \cfgq_fll_int[21] ;
 wire \cfgq_fll_int[22] ;
 wire \cfgq_fll_int[23] ;
 wire \cfgq_fll_int[24] ;
 wire \cfgq_fll_int[25] ;
 wire \cfgq_fll_int[26] ;
 wire \cfgq_fll_int[27] ;
 wire \cfgq_fll_int[28] ;
 wire \cfgq_fll_int[29] ;
 wire \cfgq_fll_int[2] ;
 wire \cfgq_fll_int[30] ;
 wire \cfgq_fll_int[31] ;
 wire \cfgq_fll_int[3] ;
 wire \cfgq_fll_int[4] ;
 wire \cfgq_fll_int[5] ;
 wire \cfgq_fll_int[6] ;
 wire \cfgq_fll_int[7] ;
 wire \cfgq_fll_int[8] ;
 wire \cfgq_fll_int[9] ;
 wire cfgreq_fll_int;
 wire cfgweb_n_fll_int;
 wire clk_gate_core_int;
 wire clk_int;
 wire core_busy_int;
 wire \data_ram_dout1[0] ;
 wire \data_ram_dout1[10] ;
 wire \data_ram_dout1[11] ;
 wire \data_ram_dout1[12] ;
 wire \data_ram_dout1[13] ;
 wire \data_ram_dout1[14] ;
 wire \data_ram_dout1[15] ;
 wire \data_ram_dout1[16] ;
 wire \data_ram_dout1[17] ;
 wire \data_ram_dout1[18] ;
 wire \data_ram_dout1[19] ;
 wire \data_ram_dout1[1] ;
 wire \data_ram_dout1[20] ;
 wire \data_ram_dout1[21] ;
 wire \data_ram_dout1[22] ;
 wire \data_ram_dout1[23] ;
 wire \data_ram_dout1[24] ;
 wire \data_ram_dout1[25] ;
 wire \data_ram_dout1[26] ;
 wire \data_ram_dout1[27] ;
 wire \data_ram_dout1[28] ;
 wire \data_ram_dout1[29] ;
 wire \data_ram_dout1[2] ;
 wire \data_ram_dout1[30] ;
 wire \data_ram_dout1[31] ;
 wire \data_ram_dout1[3] ;
 wire \data_ram_dout1[4] ;
 wire \data_ram_dout1[5] ;
 wire \data_ram_dout1[6] ;
 wire \data_ram_dout1[7] ;
 wire \data_ram_dout1[8] ;
 wire \data_ram_dout1[9] ;
 wire \debug_addr[0] ;
 wire \debug_addr[10] ;
 wire \debug_addr[11] ;
 wire \debug_addr[12] ;
 wire \debug_addr[13] ;
 wire \debug_addr[14] ;
 wire \debug_addr[1] ;
 wire \debug_addr[2] ;
 wire \debug_addr[3] ;
 wire \debug_addr[4] ;
 wire \debug_addr[5] ;
 wire \debug_addr[6] ;
 wire \debug_addr[7] ;
 wire \debug_addr[8] ;
 wire \debug_addr[9] ;
 wire debug_gnt;
 wire \debug_rdata[0] ;
 wire \debug_rdata[10] ;
 wire \debug_rdata[11] ;
 wire \debug_rdata[12] ;
 wire \debug_rdata[13] ;
 wire \debug_rdata[14] ;
 wire \debug_rdata[15] ;
 wire \debug_rdata[16] ;
 wire \debug_rdata[17] ;
 wire \debug_rdata[18] ;
 wire \debug_rdata[19] ;
 wire \debug_rdata[1] ;
 wire \debug_rdata[20] ;
 wire \debug_rdata[21] ;
 wire \debug_rdata[22] ;
 wire \debug_rdata[23] ;
 wire \debug_rdata[24] ;
 wire \debug_rdata[25] ;
 wire \debug_rdata[26] ;
 wire \debug_rdata[27] ;
 wire \debug_rdata[28] ;
 wire \debug_rdata[29] ;
 wire \debug_rdata[2] ;
 wire \debug_rdata[30] ;
 wire \debug_rdata[31] ;
 wire \debug_rdata[3] ;
 wire \debug_rdata[4] ;
 wire \debug_rdata[5] ;
 wire \debug_rdata[6] ;
 wire \debug_rdata[7] ;
 wire \debug_rdata[8] ;
 wire \debug_rdata[9] ;
 wire debug_req;
 wire debug_rvalid;
 wire \debug_wdata[0] ;
 wire \debug_wdata[10] ;
 wire \debug_wdata[11] ;
 wire \debug_wdata[12] ;
 wire \debug_wdata[13] ;
 wire \debug_wdata[14] ;
 wire \debug_wdata[15] ;
 wire \debug_wdata[16] ;
 wire \debug_wdata[17] ;
 wire \debug_wdata[18] ;
 wire \debug_wdata[19] ;
 wire \debug_wdata[1] ;
 wire \debug_wdata[20] ;
 wire \debug_wdata[21] ;
 wire \debug_wdata[22] ;
 wire \debug_wdata[23] ;
 wire \debug_wdata[24] ;
 wire \debug_wdata[25] ;
 wire \debug_wdata[26] ;
 wire \debug_wdata[27] ;
 wire \debug_wdata[28] ;
 wire \debug_wdata[29] ;
 wire \debug_wdata[2] ;
 wire \debug_wdata[30] ;
 wire \debug_wdata[31] ;
 wire \debug_wdata[3] ;
 wire \debug_wdata[4] ;
 wire \debug_wdata[5] ;
 wire \debug_wdata[6] ;
 wire \debug_wdata[7] ;
 wire \debug_wdata[8] ;
 wire \debug_wdata[9] ;
 wire debug_we;
 wire fetch_enable_int;
 wire \gpio_padcfg[0] ;
 wire \gpio_padcfg[100] ;
 wire \gpio_padcfg[101] ;
 wire \gpio_padcfg[102] ;
 wire \gpio_padcfg[103] ;
 wire \gpio_padcfg[104] ;
 wire \gpio_padcfg[105] ;
 wire \gpio_padcfg[106] ;
 wire \gpio_padcfg[107] ;
 wire \gpio_padcfg[108] ;
 wire \gpio_padcfg[109] ;
 wire \gpio_padcfg[10] ;
 wire \gpio_padcfg[110] ;
 wire \gpio_padcfg[111] ;
 wire \gpio_padcfg[112] ;
 wire \gpio_padcfg[113] ;
 wire \gpio_padcfg[114] ;
 wire \gpio_padcfg[115] ;
 wire \gpio_padcfg[116] ;
 wire \gpio_padcfg[117] ;
 wire \gpio_padcfg[118] ;
 wire \gpio_padcfg[119] ;
 wire \gpio_padcfg[11] ;
 wire \gpio_padcfg[120] ;
 wire \gpio_padcfg[121] ;
 wire \gpio_padcfg[122] ;
 wire \gpio_padcfg[123] ;
 wire \gpio_padcfg[124] ;
 wire \gpio_padcfg[125] ;
 wire \gpio_padcfg[126] ;
 wire \gpio_padcfg[127] ;
 wire \gpio_padcfg[128] ;
 wire \gpio_padcfg[129] ;
 wire \gpio_padcfg[12] ;
 wire \gpio_padcfg[130] ;
 wire \gpio_padcfg[131] ;
 wire \gpio_padcfg[132] ;
 wire \gpio_padcfg[133] ;
 wire \gpio_padcfg[134] ;
 wire \gpio_padcfg[135] ;
 wire \gpio_padcfg[136] ;
 wire \gpio_padcfg[137] ;
 wire \gpio_padcfg[138] ;
 wire \gpio_padcfg[139] ;
 wire \gpio_padcfg[13] ;
 wire \gpio_padcfg[140] ;
 wire \gpio_padcfg[141] ;
 wire \gpio_padcfg[142] ;
 wire \gpio_padcfg[143] ;
 wire \gpio_padcfg[144] ;
 wire \gpio_padcfg[145] ;
 wire \gpio_padcfg[146] ;
 wire \gpio_padcfg[147] ;
 wire \gpio_padcfg[148] ;
 wire \gpio_padcfg[149] ;
 wire \gpio_padcfg[14] ;
 wire \gpio_padcfg[150] ;
 wire \gpio_padcfg[151] ;
 wire \gpio_padcfg[152] ;
 wire \gpio_padcfg[153] ;
 wire \gpio_padcfg[154] ;
 wire \gpio_padcfg[155] ;
 wire \gpio_padcfg[156] ;
 wire \gpio_padcfg[157] ;
 wire \gpio_padcfg[158] ;
 wire \gpio_padcfg[159] ;
 wire \gpio_padcfg[15] ;
 wire \gpio_padcfg[160] ;
 wire \gpio_padcfg[161] ;
 wire \gpio_padcfg[162] ;
 wire \gpio_padcfg[163] ;
 wire \gpio_padcfg[164] ;
 wire \gpio_padcfg[165] ;
 wire \gpio_padcfg[166] ;
 wire \gpio_padcfg[167] ;
 wire \gpio_padcfg[168] ;
 wire \gpio_padcfg[169] ;
 wire \gpio_padcfg[16] ;
 wire \gpio_padcfg[170] ;
 wire \gpio_padcfg[171] ;
 wire \gpio_padcfg[172] ;
 wire \gpio_padcfg[173] ;
 wire \gpio_padcfg[174] ;
 wire \gpio_padcfg[175] ;
 wire \gpio_padcfg[176] ;
 wire \gpio_padcfg[177] ;
 wire \gpio_padcfg[178] ;
 wire \gpio_padcfg[179] ;
 wire \gpio_padcfg[17] ;
 wire \gpio_padcfg[180] ;
 wire \gpio_padcfg[181] ;
 wire \gpio_padcfg[182] ;
 wire \gpio_padcfg[183] ;
 wire \gpio_padcfg[184] ;
 wire \gpio_padcfg[185] ;
 wire \gpio_padcfg[186] ;
 wire \gpio_padcfg[187] ;
 wire \gpio_padcfg[188] ;
 wire \gpio_padcfg[189] ;
 wire \gpio_padcfg[18] ;
 wire \gpio_padcfg[190] ;
 wire \gpio_padcfg[191] ;
 wire \gpio_padcfg[19] ;
 wire \gpio_padcfg[1] ;
 wire \gpio_padcfg[20] ;
 wire \gpio_padcfg[21] ;
 wire \gpio_padcfg[22] ;
 wire \gpio_padcfg[23] ;
 wire \gpio_padcfg[24] ;
 wire \gpio_padcfg[25] ;
 wire \gpio_padcfg[26] ;
 wire \gpio_padcfg[27] ;
 wire \gpio_padcfg[28] ;
 wire \gpio_padcfg[29] ;
 wire \gpio_padcfg[2] ;
 wire \gpio_padcfg[30] ;
 wire \gpio_padcfg[31] ;
 wire \gpio_padcfg[32] ;
 wire \gpio_padcfg[33] ;
 wire \gpio_padcfg[34] ;
 wire \gpio_padcfg[35] ;
 wire \gpio_padcfg[36] ;
 wire \gpio_padcfg[37] ;
 wire \gpio_padcfg[38] ;
 wire \gpio_padcfg[39] ;
 wire \gpio_padcfg[3] ;
 wire \gpio_padcfg[40] ;
 wire \gpio_padcfg[41] ;
 wire \gpio_padcfg[42] ;
 wire \gpio_padcfg[43] ;
 wire \gpio_padcfg[44] ;
 wire \gpio_padcfg[45] ;
 wire \gpio_padcfg[46] ;
 wire \gpio_padcfg[47] ;
 wire \gpio_padcfg[48] ;
 wire \gpio_padcfg[49] ;
 wire \gpio_padcfg[4] ;
 wire \gpio_padcfg[50] ;
 wire \gpio_padcfg[51] ;
 wire \gpio_padcfg[52] ;
 wire \gpio_padcfg[53] ;
 wire \gpio_padcfg[54] ;
 wire \gpio_padcfg[55] ;
 wire \gpio_padcfg[56] ;
 wire \gpio_padcfg[57] ;
 wire \gpio_padcfg[58] ;
 wire \gpio_padcfg[59] ;
 wire \gpio_padcfg[5] ;
 wire \gpio_padcfg[60] ;
 wire \gpio_padcfg[61] ;
 wire \gpio_padcfg[62] ;
 wire \gpio_padcfg[63] ;
 wire \gpio_padcfg[64] ;
 wire \gpio_padcfg[65] ;
 wire \gpio_padcfg[66] ;
 wire \gpio_padcfg[67] ;
 wire \gpio_padcfg[68] ;
 wire \gpio_padcfg[69] ;
 wire \gpio_padcfg[6] ;
 wire \gpio_padcfg[70] ;
 wire \gpio_padcfg[71] ;
 wire \gpio_padcfg[72] ;
 wire \gpio_padcfg[73] ;
 wire \gpio_padcfg[74] ;
 wire \gpio_padcfg[75] ;
 wire \gpio_padcfg[76] ;
 wire \gpio_padcfg[77] ;
 wire \gpio_padcfg[78] ;
 wire \gpio_padcfg[79] ;
 wire \gpio_padcfg[7] ;
 wire \gpio_padcfg[80] ;
 wire \gpio_padcfg[81] ;
 wire \gpio_padcfg[82] ;
 wire \gpio_padcfg[83] ;
 wire \gpio_padcfg[84] ;
 wire \gpio_padcfg[85] ;
 wire \gpio_padcfg[86] ;
 wire \gpio_padcfg[87] ;
 wire \gpio_padcfg[88] ;
 wire \gpio_padcfg[89] ;
 wire \gpio_padcfg[8] ;
 wire \gpio_padcfg[90] ;
 wire \gpio_padcfg[91] ;
 wire \gpio_padcfg[92] ;
 wire \gpio_padcfg[93] ;
 wire \gpio_padcfg[94] ;
 wire \gpio_padcfg[95] ;
 wire \gpio_padcfg[96] ;
 wire \gpio_padcfg[97] ;
 wire \gpio_padcfg[98] ;
 wire \gpio_padcfg[99] ;
 wire \gpio_padcfg[9] ;
 wire \instr_ram_dout1[0] ;
 wire \instr_ram_dout1[10] ;
 wire \instr_ram_dout1[11] ;
 wire \instr_ram_dout1[12] ;
 wire \instr_ram_dout1[13] ;
 wire \instr_ram_dout1[14] ;
 wire \instr_ram_dout1[15] ;
 wire \instr_ram_dout1[16] ;
 wire \instr_ram_dout1[17] ;
 wire \instr_ram_dout1[18] ;
 wire \instr_ram_dout1[19] ;
 wire \instr_ram_dout1[1] ;
 wire \instr_ram_dout1[20] ;
 wire \instr_ram_dout1[21] ;
 wire \instr_ram_dout1[22] ;
 wire \instr_ram_dout1[23] ;
 wire \instr_ram_dout1[24] ;
 wire \instr_ram_dout1[25] ;
 wire \instr_ram_dout1[26] ;
 wire \instr_ram_dout1[27] ;
 wire \instr_ram_dout1[28] ;
 wire \instr_ram_dout1[29] ;
 wire \instr_ram_dout1[2] ;
 wire \instr_ram_dout1[30] ;
 wire \instr_ram_dout1[31] ;
 wire \instr_ram_dout1[3] ;
 wire \instr_ram_dout1[4] ;
 wire \instr_ram_dout1[5] ;
 wire \instr_ram_dout1[6] ;
 wire \instr_ram_dout1[7] ;
 wire \instr_ram_dout1[8] ;
 wire \instr_ram_dout1[9] ;
 wire \irq_to_core_int[0] ;
 wire \irq_to_core_int[10] ;
 wire \irq_to_core_int[11] ;
 wire \irq_to_core_int[12] ;
 wire \irq_to_core_int[13] ;
 wire \irq_to_core_int[14] ;
 wire \irq_to_core_int[15] ;
 wire \irq_to_core_int[16] ;
 wire \irq_to_core_int[17] ;
 wire \irq_to_core_int[18] ;
 wire \irq_to_core_int[19] ;
 wire \irq_to_core_int[1] ;
 wire \irq_to_core_int[20] ;
 wire \irq_to_core_int[21] ;
 wire \irq_to_core_int[22] ;
 wire \irq_to_core_int[23] ;
 wire \irq_to_core_int[24] ;
 wire \irq_to_core_int[25] ;
 wire \irq_to_core_int[26] ;
 wire \irq_to_core_int[27] ;
 wire \irq_to_core_int[28] ;
 wire \irq_to_core_int[29] ;
 wire \irq_to_core_int[2] ;
 wire \irq_to_core_int[30] ;
 wire \irq_to_core_int[31] ;
 wire \irq_to_core_int[3] ;
 wire \irq_to_core_int[4] ;
 wire \irq_to_core_int[5] ;
 wire \irq_to_core_int[6] ;
 wire \irq_to_core_int[7] ;
 wire \irq_to_core_int[8] ;
 wire \irq_to_core_int[9] ;
 wire lock_fll_int;
 wire \masters_00_ar_addr[0] ;
 wire \masters_00_ar_addr[10] ;
 wire \masters_00_ar_addr[11] ;
 wire \masters_00_ar_addr[12] ;
 wire \masters_00_ar_addr[13] ;
 wire \masters_00_ar_addr[14] ;
 wire \masters_00_ar_addr[15] ;
 wire \masters_00_ar_addr[16] ;
 wire \masters_00_ar_addr[17] ;
 wire \masters_00_ar_addr[18] ;
 wire \masters_00_ar_addr[19] ;
 wire \masters_00_ar_addr[1] ;
 wire \masters_00_ar_addr[20] ;
 wire \masters_00_ar_addr[21] ;
 wire \masters_00_ar_addr[22] ;
 wire \masters_00_ar_addr[23] ;
 wire \masters_00_ar_addr[24] ;
 wire \masters_00_ar_addr[25] ;
 wire \masters_00_ar_addr[26] ;
 wire \masters_00_ar_addr[27] ;
 wire \masters_00_ar_addr[28] ;
 wire \masters_00_ar_addr[29] ;
 wire \masters_00_ar_addr[2] ;
 wire \masters_00_ar_addr[30] ;
 wire \masters_00_ar_addr[31] ;
 wire \masters_00_ar_addr[3] ;
 wire \masters_00_ar_addr[4] ;
 wire \masters_00_ar_addr[5] ;
 wire \masters_00_ar_addr[6] ;
 wire \masters_00_ar_addr[7] ;
 wire \masters_00_ar_addr[8] ;
 wire \masters_00_ar_addr[9] ;
 wire \masters_00_ar_burst[0] ;
 wire \masters_00_ar_burst[1] ;
 wire \masters_00_ar_cache[0] ;
 wire \masters_00_ar_cache[1] ;
 wire \masters_00_ar_cache[2] ;
 wire \masters_00_ar_cache[3] ;
 wire \masters_00_ar_len[0] ;
 wire \masters_00_ar_len[1] ;
 wire \masters_00_ar_len[2] ;
 wire \masters_00_ar_len[3] ;
 wire \masters_00_ar_len[4] ;
 wire \masters_00_ar_len[5] ;
 wire \masters_00_ar_len[6] ;
 wire \masters_00_ar_len[7] ;
 wire masters_00_ar_lock;
 wire \masters_00_ar_prot[0] ;
 wire \masters_00_ar_prot[1] ;
 wire \masters_00_ar_prot[2] ;
 wire \masters_00_ar_qos[0] ;
 wire \masters_00_ar_qos[1] ;
 wire \masters_00_ar_qos[2] ;
 wire \masters_00_ar_qos[3] ;
 wire masters_00_ar_ready;
 wire \masters_00_ar_region[0] ;
 wire \masters_00_ar_region[1] ;
 wire \masters_00_ar_region[2] ;
 wire \masters_00_ar_region[3] ;
 wire \masters_00_ar_size[0] ;
 wire \masters_00_ar_size[1] ;
 wire \masters_00_ar_size[2] ;
 wire masters_00_ar_valid;
 wire \masters_00_aw_addr[0] ;
 wire \masters_00_aw_addr[10] ;
 wire \masters_00_aw_addr[11] ;
 wire \masters_00_aw_addr[12] ;
 wire \masters_00_aw_addr[13] ;
 wire \masters_00_aw_addr[14] ;
 wire \masters_00_aw_addr[15] ;
 wire \masters_00_aw_addr[16] ;
 wire \masters_00_aw_addr[17] ;
 wire \masters_00_aw_addr[18] ;
 wire \masters_00_aw_addr[19] ;
 wire \masters_00_aw_addr[1] ;
 wire \masters_00_aw_addr[20] ;
 wire \masters_00_aw_addr[21] ;
 wire \masters_00_aw_addr[22] ;
 wire \masters_00_aw_addr[23] ;
 wire \masters_00_aw_addr[24] ;
 wire \masters_00_aw_addr[25] ;
 wire \masters_00_aw_addr[26] ;
 wire \masters_00_aw_addr[27] ;
 wire \masters_00_aw_addr[28] ;
 wire \masters_00_aw_addr[29] ;
 wire \masters_00_aw_addr[2] ;
 wire \masters_00_aw_addr[30] ;
 wire \masters_00_aw_addr[31] ;
 wire \masters_00_aw_addr[3] ;
 wire \masters_00_aw_addr[4] ;
 wire \masters_00_aw_addr[5] ;
 wire \masters_00_aw_addr[6] ;
 wire \masters_00_aw_addr[7] ;
 wire \masters_00_aw_addr[8] ;
 wire \masters_00_aw_addr[9] ;
 wire \masters_00_aw_burst[0] ;
 wire \masters_00_aw_burst[1] ;
 wire \masters_00_aw_cache[0] ;
 wire \masters_00_aw_cache[1] ;
 wire \masters_00_aw_cache[2] ;
 wire \masters_00_aw_cache[3] ;
 wire \masters_00_aw_len[0] ;
 wire \masters_00_aw_len[1] ;
 wire \masters_00_aw_len[2] ;
 wire \masters_00_aw_len[3] ;
 wire \masters_00_aw_len[4] ;
 wire \masters_00_aw_len[5] ;
 wire \masters_00_aw_len[6] ;
 wire \masters_00_aw_len[7] ;
 wire masters_00_aw_lock;
 wire \masters_00_aw_prot[0] ;
 wire \masters_00_aw_prot[1] ;
 wire \masters_00_aw_prot[2] ;
 wire \masters_00_aw_qos[0] ;
 wire \masters_00_aw_qos[1] ;
 wire \masters_00_aw_qos[2] ;
 wire \masters_00_aw_qos[3] ;
 wire masters_00_aw_ready;
 wire \masters_00_aw_region[0] ;
 wire \masters_00_aw_region[1] ;
 wire \masters_00_aw_region[2] ;
 wire \masters_00_aw_region[3] ;
 wire \masters_00_aw_size[0] ;
 wire \masters_00_aw_size[1] ;
 wire \masters_00_aw_size[2] ;
 wire masters_00_aw_valid;
 wire masters_00_b_ready;
 wire \masters_00_b_resp[0] ;
 wire \masters_00_b_resp[1] ;
 wire masters_00_b_valid;
 wire \masters_00_r_data[0] ;
 wire \masters_00_r_data[10] ;
 wire \masters_00_r_data[11] ;
 wire \masters_00_r_data[12] ;
 wire \masters_00_r_data[13] ;
 wire \masters_00_r_data[14] ;
 wire \masters_00_r_data[15] ;
 wire \masters_00_r_data[16] ;
 wire \masters_00_r_data[17] ;
 wire \masters_00_r_data[18] ;
 wire \masters_00_r_data[19] ;
 wire \masters_00_r_data[1] ;
 wire \masters_00_r_data[20] ;
 wire \masters_00_r_data[21] ;
 wire \masters_00_r_data[22] ;
 wire \masters_00_r_data[23] ;
 wire \masters_00_r_data[24] ;
 wire \masters_00_r_data[25] ;
 wire \masters_00_r_data[26] ;
 wire \masters_00_r_data[27] ;
 wire \masters_00_r_data[28] ;
 wire \masters_00_r_data[29] ;
 wire \masters_00_r_data[2] ;
 wire \masters_00_r_data[30] ;
 wire \masters_00_r_data[31] ;
 wire \masters_00_r_data[3] ;
 wire \masters_00_r_data[4] ;
 wire \masters_00_r_data[5] ;
 wire \masters_00_r_data[6] ;
 wire \masters_00_r_data[7] ;
 wire \masters_00_r_data[8] ;
 wire \masters_00_r_data[9] ;
 wire masters_00_r_last;
 wire masters_00_r_ready;
 wire \masters_00_r_resp[0] ;
 wire \masters_00_r_resp[1] ;
 wire masters_00_r_valid;
 wire \masters_00_w_data[0] ;
 wire \masters_00_w_data[10] ;
 wire \masters_00_w_data[11] ;
 wire \masters_00_w_data[12] ;
 wire \masters_00_w_data[13] ;
 wire \masters_00_w_data[14] ;
 wire \masters_00_w_data[15] ;
 wire \masters_00_w_data[16] ;
 wire \masters_00_w_data[17] ;
 wire \masters_00_w_data[18] ;
 wire \masters_00_w_data[19] ;
 wire \masters_00_w_data[1] ;
 wire \masters_00_w_data[20] ;
 wire \masters_00_w_data[21] ;
 wire \masters_00_w_data[22] ;
 wire \masters_00_w_data[23] ;
 wire \masters_00_w_data[24] ;
 wire \masters_00_w_data[25] ;
 wire \masters_00_w_data[26] ;
 wire \masters_00_w_data[27] ;
 wire \masters_00_w_data[28] ;
 wire \masters_00_w_data[29] ;
 wire \masters_00_w_data[2] ;
 wire \masters_00_w_data[30] ;
 wire \masters_00_w_data[31] ;
 wire \masters_00_w_data[3] ;
 wire \masters_00_w_data[4] ;
 wire \masters_00_w_data[5] ;
 wire \masters_00_w_data[6] ;
 wire \masters_00_w_data[7] ;
 wire \masters_00_w_data[8] ;
 wire \masters_00_w_data[9] ;
 wire masters_00_w_last;
 wire masters_00_w_ready;
 wire \masters_00_w_strb[0] ;
 wire \masters_00_w_strb[1] ;
 wire \masters_00_w_strb[2] ;
 wire \masters_00_w_strb[3] ;
 wire masters_00_w_valid;
 wire \masters_01_ar_addr[0] ;
 wire \masters_01_ar_addr[10] ;
 wire \masters_01_ar_addr[11] ;
 wire \masters_01_ar_addr[12] ;
 wire \masters_01_ar_addr[13] ;
 wire \masters_01_ar_addr[14] ;
 wire \masters_01_ar_addr[15] ;
 wire \masters_01_ar_addr[16] ;
 wire \masters_01_ar_addr[17] ;
 wire \masters_01_ar_addr[18] ;
 wire \masters_01_ar_addr[19] ;
 wire \masters_01_ar_addr[1] ;
 wire \masters_01_ar_addr[20] ;
 wire \masters_01_ar_addr[21] ;
 wire \masters_01_ar_addr[22] ;
 wire \masters_01_ar_addr[23] ;
 wire \masters_01_ar_addr[24] ;
 wire \masters_01_ar_addr[25] ;
 wire \masters_01_ar_addr[26] ;
 wire \masters_01_ar_addr[27] ;
 wire \masters_01_ar_addr[28] ;
 wire \masters_01_ar_addr[29] ;
 wire \masters_01_ar_addr[2] ;
 wire \masters_01_ar_addr[30] ;
 wire \masters_01_ar_addr[31] ;
 wire \masters_01_ar_addr[3] ;
 wire \masters_01_ar_addr[4] ;
 wire \masters_01_ar_addr[5] ;
 wire \masters_01_ar_addr[6] ;
 wire \masters_01_ar_addr[7] ;
 wire \masters_01_ar_addr[8] ;
 wire \masters_01_ar_addr[9] ;
 wire \masters_01_ar_burst[0] ;
 wire \masters_01_ar_burst[1] ;
 wire \masters_01_ar_cache[0] ;
 wire \masters_01_ar_cache[1] ;
 wire \masters_01_ar_cache[2] ;
 wire \masters_01_ar_cache[3] ;
 wire \masters_01_ar_len[0] ;
 wire \masters_01_ar_len[1] ;
 wire \masters_01_ar_len[2] ;
 wire \masters_01_ar_len[3] ;
 wire \masters_01_ar_len[4] ;
 wire \masters_01_ar_len[5] ;
 wire \masters_01_ar_len[6] ;
 wire \masters_01_ar_len[7] ;
 wire masters_01_ar_lock;
 wire \masters_01_ar_prot[0] ;
 wire \masters_01_ar_prot[1] ;
 wire \masters_01_ar_prot[2] ;
 wire \masters_01_ar_qos[0] ;
 wire \masters_01_ar_qos[1] ;
 wire \masters_01_ar_qos[2] ;
 wire \masters_01_ar_qos[3] ;
 wire masters_01_ar_ready;
 wire \masters_01_ar_region[0] ;
 wire \masters_01_ar_region[1] ;
 wire \masters_01_ar_region[2] ;
 wire \masters_01_ar_region[3] ;
 wire \masters_01_ar_size[0] ;
 wire \masters_01_ar_size[1] ;
 wire \masters_01_ar_size[2] ;
 wire masters_01_ar_valid;
 wire \masters_01_aw_addr[0] ;
 wire \masters_01_aw_addr[10] ;
 wire \masters_01_aw_addr[11] ;
 wire \masters_01_aw_addr[12] ;
 wire \masters_01_aw_addr[13] ;
 wire \masters_01_aw_addr[14] ;
 wire \masters_01_aw_addr[15] ;
 wire \masters_01_aw_addr[16] ;
 wire \masters_01_aw_addr[17] ;
 wire \masters_01_aw_addr[18] ;
 wire \masters_01_aw_addr[19] ;
 wire \masters_01_aw_addr[1] ;
 wire \masters_01_aw_addr[20] ;
 wire \masters_01_aw_addr[21] ;
 wire \masters_01_aw_addr[22] ;
 wire \masters_01_aw_addr[23] ;
 wire \masters_01_aw_addr[24] ;
 wire \masters_01_aw_addr[25] ;
 wire \masters_01_aw_addr[26] ;
 wire \masters_01_aw_addr[27] ;
 wire \masters_01_aw_addr[28] ;
 wire \masters_01_aw_addr[29] ;
 wire \masters_01_aw_addr[2] ;
 wire \masters_01_aw_addr[30] ;
 wire \masters_01_aw_addr[31] ;
 wire \masters_01_aw_addr[3] ;
 wire \masters_01_aw_addr[4] ;
 wire \masters_01_aw_addr[5] ;
 wire \masters_01_aw_addr[6] ;
 wire \masters_01_aw_addr[7] ;
 wire \masters_01_aw_addr[8] ;
 wire \masters_01_aw_addr[9] ;
 wire \masters_01_aw_burst[0] ;
 wire \masters_01_aw_burst[1] ;
 wire \masters_01_aw_cache[0] ;
 wire \masters_01_aw_cache[1] ;
 wire \masters_01_aw_cache[2] ;
 wire \masters_01_aw_cache[3] ;
 wire \masters_01_aw_len[0] ;
 wire \masters_01_aw_len[1] ;
 wire \masters_01_aw_len[2] ;
 wire \masters_01_aw_len[3] ;
 wire \masters_01_aw_len[4] ;
 wire \masters_01_aw_len[5] ;
 wire \masters_01_aw_len[6] ;
 wire \masters_01_aw_len[7] ;
 wire masters_01_aw_lock;
 wire \masters_01_aw_prot[0] ;
 wire \masters_01_aw_prot[1] ;
 wire \masters_01_aw_prot[2] ;
 wire \masters_01_aw_qos[0] ;
 wire \masters_01_aw_qos[1] ;
 wire \masters_01_aw_qos[2] ;
 wire \masters_01_aw_qos[3] ;
 wire masters_01_aw_ready;
 wire \masters_01_aw_region[0] ;
 wire \masters_01_aw_region[1] ;
 wire \masters_01_aw_region[2] ;
 wire \masters_01_aw_region[3] ;
 wire \masters_01_aw_size[0] ;
 wire \masters_01_aw_size[1] ;
 wire \masters_01_aw_size[2] ;
 wire masters_01_aw_valid;
 wire masters_01_b_ready;
 wire \masters_01_b_resp[0] ;
 wire \masters_01_b_resp[1] ;
 wire masters_01_b_valid;
 wire \masters_01_r_data[0] ;
 wire \masters_01_r_data[10] ;
 wire \masters_01_r_data[11] ;
 wire \masters_01_r_data[12] ;
 wire \masters_01_r_data[13] ;
 wire \masters_01_r_data[14] ;
 wire \masters_01_r_data[15] ;
 wire \masters_01_r_data[16] ;
 wire \masters_01_r_data[17] ;
 wire \masters_01_r_data[18] ;
 wire \masters_01_r_data[19] ;
 wire \masters_01_r_data[1] ;
 wire \masters_01_r_data[20] ;
 wire \masters_01_r_data[21] ;
 wire \masters_01_r_data[22] ;
 wire \masters_01_r_data[23] ;
 wire \masters_01_r_data[24] ;
 wire \masters_01_r_data[25] ;
 wire \masters_01_r_data[26] ;
 wire \masters_01_r_data[27] ;
 wire \masters_01_r_data[28] ;
 wire \masters_01_r_data[29] ;
 wire \masters_01_r_data[2] ;
 wire \masters_01_r_data[30] ;
 wire \masters_01_r_data[31] ;
 wire \masters_01_r_data[3] ;
 wire \masters_01_r_data[4] ;
 wire \masters_01_r_data[5] ;
 wire \masters_01_r_data[6] ;
 wire \masters_01_r_data[7] ;
 wire \masters_01_r_data[8] ;
 wire \masters_01_r_data[9] ;
 wire masters_01_r_last;
 wire masters_01_r_ready;
 wire \masters_01_r_resp[0] ;
 wire \masters_01_r_resp[1] ;
 wire masters_01_r_valid;
 wire \masters_01_w_data[0] ;
 wire \masters_01_w_data[10] ;
 wire \masters_01_w_data[11] ;
 wire \masters_01_w_data[12] ;
 wire \masters_01_w_data[13] ;
 wire \masters_01_w_data[14] ;
 wire \masters_01_w_data[15] ;
 wire \masters_01_w_data[16] ;
 wire \masters_01_w_data[17] ;
 wire \masters_01_w_data[18] ;
 wire \masters_01_w_data[19] ;
 wire \masters_01_w_data[1] ;
 wire \masters_01_w_data[20] ;
 wire \masters_01_w_data[21] ;
 wire \masters_01_w_data[22] ;
 wire \masters_01_w_data[23] ;
 wire \masters_01_w_data[24] ;
 wire \masters_01_w_data[25] ;
 wire \masters_01_w_data[26] ;
 wire \masters_01_w_data[27] ;
 wire \masters_01_w_data[28] ;
 wire \masters_01_w_data[29] ;
 wire \masters_01_w_data[2] ;
 wire \masters_01_w_data[30] ;
 wire \masters_01_w_data[31] ;
 wire \masters_01_w_data[3] ;
 wire \masters_01_w_data[4] ;
 wire \masters_01_w_data[5] ;
 wire \masters_01_w_data[6] ;
 wire \masters_01_w_data[7] ;
 wire \masters_01_w_data[8] ;
 wire \masters_01_w_data[9] ;
 wire masters_01_w_last;
 wire masters_01_w_ready;
 wire \masters_01_w_strb[0] ;
 wire \masters_01_w_strb[1] ;
 wire \masters_01_w_strb[2] ;
 wire \masters_01_w_strb[3] ;
 wire masters_01_w_valid;
 wire \masters_02_ar_addr[0] ;
 wire \masters_02_ar_addr[10] ;
 wire \masters_02_ar_addr[11] ;
 wire \masters_02_ar_addr[12] ;
 wire \masters_02_ar_addr[13] ;
 wire \masters_02_ar_addr[14] ;
 wire \masters_02_ar_addr[15] ;
 wire \masters_02_ar_addr[16] ;
 wire \masters_02_ar_addr[17] ;
 wire \masters_02_ar_addr[18] ;
 wire \masters_02_ar_addr[19] ;
 wire \masters_02_ar_addr[1] ;
 wire \masters_02_ar_addr[20] ;
 wire \masters_02_ar_addr[21] ;
 wire \masters_02_ar_addr[22] ;
 wire \masters_02_ar_addr[23] ;
 wire \masters_02_ar_addr[24] ;
 wire \masters_02_ar_addr[25] ;
 wire \masters_02_ar_addr[26] ;
 wire \masters_02_ar_addr[27] ;
 wire \masters_02_ar_addr[28] ;
 wire \masters_02_ar_addr[29] ;
 wire \masters_02_ar_addr[2] ;
 wire \masters_02_ar_addr[30] ;
 wire \masters_02_ar_addr[31] ;
 wire \masters_02_ar_addr[3] ;
 wire \masters_02_ar_addr[4] ;
 wire \masters_02_ar_addr[5] ;
 wire \masters_02_ar_addr[6] ;
 wire \masters_02_ar_addr[7] ;
 wire \masters_02_ar_addr[8] ;
 wire \masters_02_ar_addr[9] ;
 wire \masters_02_ar_burst[0] ;
 wire \masters_02_ar_burst[1] ;
 wire \masters_02_ar_cache[0] ;
 wire \masters_02_ar_cache[1] ;
 wire \masters_02_ar_cache[2] ;
 wire \masters_02_ar_cache[3] ;
 wire \masters_02_ar_len[0] ;
 wire \masters_02_ar_len[1] ;
 wire \masters_02_ar_len[2] ;
 wire \masters_02_ar_len[3] ;
 wire \masters_02_ar_len[4] ;
 wire \masters_02_ar_len[5] ;
 wire \masters_02_ar_len[6] ;
 wire \masters_02_ar_len[7] ;
 wire masters_02_ar_lock;
 wire \masters_02_ar_prot[0] ;
 wire \masters_02_ar_prot[1] ;
 wire \masters_02_ar_prot[2] ;
 wire \masters_02_ar_qos[0] ;
 wire \masters_02_ar_qos[1] ;
 wire \masters_02_ar_qos[2] ;
 wire \masters_02_ar_qos[3] ;
 wire masters_02_ar_ready;
 wire \masters_02_ar_region[0] ;
 wire \masters_02_ar_region[1] ;
 wire \masters_02_ar_region[2] ;
 wire \masters_02_ar_region[3] ;
 wire \masters_02_ar_size[0] ;
 wire \masters_02_ar_size[1] ;
 wire \masters_02_ar_size[2] ;
 wire masters_02_ar_valid;
 wire \masters_02_aw_addr[0] ;
 wire \masters_02_aw_addr[10] ;
 wire \masters_02_aw_addr[11] ;
 wire \masters_02_aw_addr[12] ;
 wire \masters_02_aw_addr[13] ;
 wire \masters_02_aw_addr[14] ;
 wire \masters_02_aw_addr[15] ;
 wire \masters_02_aw_addr[16] ;
 wire \masters_02_aw_addr[17] ;
 wire \masters_02_aw_addr[18] ;
 wire \masters_02_aw_addr[19] ;
 wire \masters_02_aw_addr[1] ;
 wire \masters_02_aw_addr[20] ;
 wire \masters_02_aw_addr[21] ;
 wire \masters_02_aw_addr[22] ;
 wire \masters_02_aw_addr[23] ;
 wire \masters_02_aw_addr[24] ;
 wire \masters_02_aw_addr[25] ;
 wire \masters_02_aw_addr[26] ;
 wire \masters_02_aw_addr[27] ;
 wire \masters_02_aw_addr[28] ;
 wire \masters_02_aw_addr[29] ;
 wire \masters_02_aw_addr[2] ;
 wire \masters_02_aw_addr[30] ;
 wire \masters_02_aw_addr[31] ;
 wire \masters_02_aw_addr[3] ;
 wire \masters_02_aw_addr[4] ;
 wire \masters_02_aw_addr[5] ;
 wire \masters_02_aw_addr[6] ;
 wire \masters_02_aw_addr[7] ;
 wire \masters_02_aw_addr[8] ;
 wire \masters_02_aw_addr[9] ;
 wire \masters_02_aw_burst[0] ;
 wire \masters_02_aw_burst[1] ;
 wire \masters_02_aw_cache[0] ;
 wire \masters_02_aw_cache[1] ;
 wire \masters_02_aw_cache[2] ;
 wire \masters_02_aw_cache[3] ;
 wire \masters_02_aw_len[0] ;
 wire \masters_02_aw_len[1] ;
 wire \masters_02_aw_len[2] ;
 wire \masters_02_aw_len[3] ;
 wire \masters_02_aw_len[4] ;
 wire \masters_02_aw_len[5] ;
 wire \masters_02_aw_len[6] ;
 wire \masters_02_aw_len[7] ;
 wire masters_02_aw_lock;
 wire \masters_02_aw_prot[0] ;
 wire \masters_02_aw_prot[1] ;
 wire \masters_02_aw_prot[2] ;
 wire \masters_02_aw_qos[0] ;
 wire \masters_02_aw_qos[1] ;
 wire \masters_02_aw_qos[2] ;
 wire \masters_02_aw_qos[3] ;
 wire masters_02_aw_ready;
 wire \masters_02_aw_region[0] ;
 wire \masters_02_aw_region[1] ;
 wire \masters_02_aw_region[2] ;
 wire \masters_02_aw_region[3] ;
 wire \masters_02_aw_size[0] ;
 wire \masters_02_aw_size[1] ;
 wire \masters_02_aw_size[2] ;
 wire masters_02_aw_valid;
 wire masters_02_b_ready;
 wire \masters_02_b_resp[0] ;
 wire \masters_02_b_resp[1] ;
 wire masters_02_b_valid;
 wire \masters_02_r_data[0] ;
 wire \masters_02_r_data[10] ;
 wire \masters_02_r_data[11] ;
 wire \masters_02_r_data[12] ;
 wire \masters_02_r_data[13] ;
 wire \masters_02_r_data[14] ;
 wire \masters_02_r_data[15] ;
 wire \masters_02_r_data[16] ;
 wire \masters_02_r_data[17] ;
 wire \masters_02_r_data[18] ;
 wire \masters_02_r_data[19] ;
 wire \masters_02_r_data[1] ;
 wire \masters_02_r_data[20] ;
 wire \masters_02_r_data[21] ;
 wire \masters_02_r_data[22] ;
 wire \masters_02_r_data[23] ;
 wire \masters_02_r_data[24] ;
 wire \masters_02_r_data[25] ;
 wire \masters_02_r_data[26] ;
 wire \masters_02_r_data[27] ;
 wire \masters_02_r_data[28] ;
 wire \masters_02_r_data[29] ;
 wire \masters_02_r_data[2] ;
 wire \masters_02_r_data[30] ;
 wire \masters_02_r_data[31] ;
 wire \masters_02_r_data[3] ;
 wire \masters_02_r_data[4] ;
 wire \masters_02_r_data[5] ;
 wire \masters_02_r_data[6] ;
 wire \masters_02_r_data[7] ;
 wire \masters_02_r_data[8] ;
 wire \masters_02_r_data[9] ;
 wire masters_02_r_last;
 wire masters_02_r_ready;
 wire \masters_02_r_resp[0] ;
 wire \masters_02_r_resp[1] ;
 wire masters_02_r_valid;
 wire \masters_02_w_data[0] ;
 wire \masters_02_w_data[10] ;
 wire \masters_02_w_data[11] ;
 wire \masters_02_w_data[12] ;
 wire \masters_02_w_data[13] ;
 wire \masters_02_w_data[14] ;
 wire \masters_02_w_data[15] ;
 wire \masters_02_w_data[16] ;
 wire \masters_02_w_data[17] ;
 wire \masters_02_w_data[18] ;
 wire \masters_02_w_data[19] ;
 wire \masters_02_w_data[1] ;
 wire \masters_02_w_data[20] ;
 wire \masters_02_w_data[21] ;
 wire \masters_02_w_data[22] ;
 wire \masters_02_w_data[23] ;
 wire \masters_02_w_data[24] ;
 wire \masters_02_w_data[25] ;
 wire \masters_02_w_data[26] ;
 wire \masters_02_w_data[27] ;
 wire \masters_02_w_data[28] ;
 wire \masters_02_w_data[29] ;
 wire \masters_02_w_data[2] ;
 wire \masters_02_w_data[30] ;
 wire \masters_02_w_data[31] ;
 wire \masters_02_w_data[3] ;
 wire \masters_02_w_data[4] ;
 wire \masters_02_w_data[5] ;
 wire \masters_02_w_data[6] ;
 wire \masters_02_w_data[7] ;
 wire \masters_02_w_data[8] ;
 wire \masters_02_w_data[9] ;
 wire masters_02_w_last;
 wire masters_02_w_ready;
 wire \masters_02_w_strb[0] ;
 wire \masters_02_w_strb[1] ;
 wire \masters_02_w_strb[2] ;
 wire \masters_02_w_strb[3] ;
 wire masters_02_w_valid;
 wire \mba_data_mem_addr0_o[0] ;
 wire \mba_data_mem_addr0_o[10] ;
 wire \mba_data_mem_addr0_o[11] ;
 wire \mba_data_mem_addr0_o[12] ;
 wire \mba_data_mem_addr0_o[13] ;
 wire \mba_data_mem_addr0_o[14] ;
 wire \mba_data_mem_addr0_o[15] ;
 wire \mba_data_mem_addr0_o[16] ;
 wire \mba_data_mem_addr0_o[17] ;
 wire \mba_data_mem_addr0_o[18] ;
 wire \mba_data_mem_addr0_o[19] ;
 wire \mba_data_mem_addr0_o[1] ;
 wire \mba_data_mem_addr0_o[20] ;
 wire \mba_data_mem_addr0_o[21] ;
 wire \mba_data_mem_addr0_o[22] ;
 wire \mba_data_mem_addr0_o[23] ;
 wire \mba_data_mem_addr0_o[24] ;
 wire \mba_data_mem_addr0_o[25] ;
 wire \mba_data_mem_addr0_o[26] ;
 wire \mba_data_mem_addr0_o[27] ;
 wire \mba_data_mem_addr0_o[28] ;
 wire \mba_data_mem_addr0_o[29] ;
 wire \mba_data_mem_addr0_o[2] ;
 wire \mba_data_mem_addr0_o[30] ;
 wire \mba_data_mem_addr0_o[31] ;
 wire \mba_data_mem_addr0_o[3] ;
 wire \mba_data_mem_addr0_o[4] ;
 wire \mba_data_mem_addr0_o[5] ;
 wire \mba_data_mem_addr0_o[6] ;
 wire \mba_data_mem_addr0_o[7] ;
 wire \mba_data_mem_addr0_o[8] ;
 wire \mba_data_mem_addr0_o[9] ;
 wire \mba_data_mem_addr1_o[0] ;
 wire \mba_data_mem_addr1_o[10] ;
 wire \mba_data_mem_addr1_o[11] ;
 wire \mba_data_mem_addr1_o[12] ;
 wire \mba_data_mem_addr1_o[13] ;
 wire \mba_data_mem_addr1_o[14] ;
 wire \mba_data_mem_addr1_o[15] ;
 wire \mba_data_mem_addr1_o[16] ;
 wire \mba_data_mem_addr1_o[17] ;
 wire \mba_data_mem_addr1_o[18] ;
 wire \mba_data_mem_addr1_o[19] ;
 wire \mba_data_mem_addr1_o[1] ;
 wire \mba_data_mem_addr1_o[20] ;
 wire \mba_data_mem_addr1_o[21] ;
 wire \mba_data_mem_addr1_o[22] ;
 wire \mba_data_mem_addr1_o[23] ;
 wire \mba_data_mem_addr1_o[24] ;
 wire \mba_data_mem_addr1_o[25] ;
 wire \mba_data_mem_addr1_o[26] ;
 wire \mba_data_mem_addr1_o[27] ;
 wire \mba_data_mem_addr1_o[28] ;
 wire \mba_data_mem_addr1_o[29] ;
 wire \mba_data_mem_addr1_o[2] ;
 wire \mba_data_mem_addr1_o[30] ;
 wire \mba_data_mem_addr1_o[31] ;
 wire \mba_data_mem_addr1_o[3] ;
 wire \mba_data_mem_addr1_o[4] ;
 wire \mba_data_mem_addr1_o[5] ;
 wire \mba_data_mem_addr1_o[6] ;
 wire \mba_data_mem_addr1_o[7] ;
 wire \mba_data_mem_addr1_o[8] ;
 wire \mba_data_mem_addr1_o[9] ;
 wire mba_data_mem_csb0_o;
 wire mba_data_mem_csb1_o;
 wire \mba_data_mem_din0_o[0] ;
 wire \mba_data_mem_din0_o[10] ;
 wire \mba_data_mem_din0_o[11] ;
 wire \mba_data_mem_din0_o[12] ;
 wire \mba_data_mem_din0_o[13] ;
 wire \mba_data_mem_din0_o[14] ;
 wire \mba_data_mem_din0_o[15] ;
 wire \mba_data_mem_din0_o[16] ;
 wire \mba_data_mem_din0_o[17] ;
 wire \mba_data_mem_din0_o[18] ;
 wire \mba_data_mem_din0_o[19] ;
 wire \mba_data_mem_din0_o[1] ;
 wire \mba_data_mem_din0_o[20] ;
 wire \mba_data_mem_din0_o[21] ;
 wire \mba_data_mem_din0_o[22] ;
 wire \mba_data_mem_din0_o[23] ;
 wire \mba_data_mem_din0_o[24] ;
 wire \mba_data_mem_din0_o[25] ;
 wire \mba_data_mem_din0_o[26] ;
 wire \mba_data_mem_din0_o[27] ;
 wire \mba_data_mem_din0_o[28] ;
 wire \mba_data_mem_din0_o[29] ;
 wire \mba_data_mem_din0_o[2] ;
 wire \mba_data_mem_din0_o[30] ;
 wire \mba_data_mem_din0_o[31] ;
 wire \mba_data_mem_din0_o[3] ;
 wire \mba_data_mem_din0_o[4] ;
 wire \mba_data_mem_din0_o[5] ;
 wire \mba_data_mem_din0_o[6] ;
 wire \mba_data_mem_din0_o[7] ;
 wire \mba_data_mem_din0_o[8] ;
 wire \mba_data_mem_din0_o[9] ;
 wire \mba_data_mem_dout0_i[0] ;
 wire \mba_data_mem_dout0_i[10] ;
 wire \mba_data_mem_dout0_i[11] ;
 wire \mba_data_mem_dout0_i[12] ;
 wire \mba_data_mem_dout0_i[13] ;
 wire \mba_data_mem_dout0_i[14] ;
 wire \mba_data_mem_dout0_i[15] ;
 wire \mba_data_mem_dout0_i[16] ;
 wire \mba_data_mem_dout0_i[17] ;
 wire \mba_data_mem_dout0_i[18] ;
 wire \mba_data_mem_dout0_i[19] ;
 wire \mba_data_mem_dout0_i[1] ;
 wire \mba_data_mem_dout0_i[20] ;
 wire \mba_data_mem_dout0_i[21] ;
 wire \mba_data_mem_dout0_i[22] ;
 wire \mba_data_mem_dout0_i[23] ;
 wire \mba_data_mem_dout0_i[24] ;
 wire \mba_data_mem_dout0_i[25] ;
 wire \mba_data_mem_dout0_i[26] ;
 wire \mba_data_mem_dout0_i[27] ;
 wire \mba_data_mem_dout0_i[28] ;
 wire \mba_data_mem_dout0_i[29] ;
 wire \mba_data_mem_dout0_i[2] ;
 wire \mba_data_mem_dout0_i[30] ;
 wire \mba_data_mem_dout0_i[31] ;
 wire \mba_data_mem_dout0_i[3] ;
 wire \mba_data_mem_dout0_i[4] ;
 wire \mba_data_mem_dout0_i[5] ;
 wire \mba_data_mem_dout0_i[6] ;
 wire \mba_data_mem_dout0_i[7] ;
 wire \mba_data_mem_dout0_i[8] ;
 wire \mba_data_mem_dout0_i[9] ;
 wire mba_data_mem_web0_o;
 wire \mba_data_mem_wmask0_o[0] ;
 wire \mba_data_mem_wmask0_o[1] ;
 wire \mba_data_mem_wmask0_o[2] ;
 wire \mba_data_mem_wmask0_o[3] ;
 wire \mba_instr_mem_addr0_o[0] ;
 wire \mba_instr_mem_addr0_o[10] ;
 wire \mba_instr_mem_addr0_o[11] ;
 wire \mba_instr_mem_addr0_o[12] ;
 wire \mba_instr_mem_addr0_o[13] ;
 wire \mba_instr_mem_addr0_o[14] ;
 wire \mba_instr_mem_addr0_o[15] ;
 wire \mba_instr_mem_addr0_o[16] ;
 wire \mba_instr_mem_addr0_o[17] ;
 wire \mba_instr_mem_addr0_o[18] ;
 wire \mba_instr_mem_addr0_o[19] ;
 wire \mba_instr_mem_addr0_o[1] ;
 wire \mba_instr_mem_addr0_o[20] ;
 wire \mba_instr_mem_addr0_o[21] ;
 wire \mba_instr_mem_addr0_o[22] ;
 wire \mba_instr_mem_addr0_o[23] ;
 wire \mba_instr_mem_addr0_o[24] ;
 wire \mba_instr_mem_addr0_o[25] ;
 wire \mba_instr_mem_addr0_o[26] ;
 wire \mba_instr_mem_addr0_o[27] ;
 wire \mba_instr_mem_addr0_o[28] ;
 wire \mba_instr_mem_addr0_o[29] ;
 wire \mba_instr_mem_addr0_o[2] ;
 wire \mba_instr_mem_addr0_o[30] ;
 wire \mba_instr_mem_addr0_o[31] ;
 wire \mba_instr_mem_addr0_o[3] ;
 wire \mba_instr_mem_addr0_o[4] ;
 wire \mba_instr_mem_addr0_o[5] ;
 wire \mba_instr_mem_addr0_o[6] ;
 wire \mba_instr_mem_addr0_o[7] ;
 wire \mba_instr_mem_addr0_o[8] ;
 wire \mba_instr_mem_addr0_o[9] ;
 wire \mba_instr_mem_addr1_o[0] ;
 wire \mba_instr_mem_addr1_o[10] ;
 wire \mba_instr_mem_addr1_o[11] ;
 wire \mba_instr_mem_addr1_o[12] ;
 wire \mba_instr_mem_addr1_o[13] ;
 wire \mba_instr_mem_addr1_o[14] ;
 wire \mba_instr_mem_addr1_o[15] ;
 wire \mba_instr_mem_addr1_o[16] ;
 wire \mba_instr_mem_addr1_o[17] ;
 wire \mba_instr_mem_addr1_o[18] ;
 wire \mba_instr_mem_addr1_o[19] ;
 wire \mba_instr_mem_addr1_o[1] ;
 wire \mba_instr_mem_addr1_o[20] ;
 wire \mba_instr_mem_addr1_o[21] ;
 wire \mba_instr_mem_addr1_o[22] ;
 wire \mba_instr_mem_addr1_o[23] ;
 wire \mba_instr_mem_addr1_o[24] ;
 wire \mba_instr_mem_addr1_o[25] ;
 wire \mba_instr_mem_addr1_o[26] ;
 wire \mba_instr_mem_addr1_o[27] ;
 wire \mba_instr_mem_addr1_o[28] ;
 wire \mba_instr_mem_addr1_o[29] ;
 wire \mba_instr_mem_addr1_o[2] ;
 wire \mba_instr_mem_addr1_o[30] ;
 wire \mba_instr_mem_addr1_o[31] ;
 wire \mba_instr_mem_addr1_o[3] ;
 wire \mba_instr_mem_addr1_o[4] ;
 wire \mba_instr_mem_addr1_o[5] ;
 wire \mba_instr_mem_addr1_o[6] ;
 wire \mba_instr_mem_addr1_o[7] ;
 wire \mba_instr_mem_addr1_o[8] ;
 wire \mba_instr_mem_addr1_o[9] ;
 wire mba_instr_mem_csb0_o;
 wire mba_instr_mem_csb1_o;
 wire \mba_instr_mem_din0_o[0] ;
 wire \mba_instr_mem_din0_o[10] ;
 wire \mba_instr_mem_din0_o[11] ;
 wire \mba_instr_mem_din0_o[12] ;
 wire \mba_instr_mem_din0_o[13] ;
 wire \mba_instr_mem_din0_o[14] ;
 wire \mba_instr_mem_din0_o[15] ;
 wire \mba_instr_mem_din0_o[16] ;
 wire \mba_instr_mem_din0_o[17] ;
 wire \mba_instr_mem_din0_o[18] ;
 wire \mba_instr_mem_din0_o[19] ;
 wire \mba_instr_mem_din0_o[1] ;
 wire \mba_instr_mem_din0_o[20] ;
 wire \mba_instr_mem_din0_o[21] ;
 wire \mba_instr_mem_din0_o[22] ;
 wire \mba_instr_mem_din0_o[23] ;
 wire \mba_instr_mem_din0_o[24] ;
 wire \mba_instr_mem_din0_o[25] ;
 wire \mba_instr_mem_din0_o[26] ;
 wire \mba_instr_mem_din0_o[27] ;
 wire \mba_instr_mem_din0_o[28] ;
 wire \mba_instr_mem_din0_o[29] ;
 wire \mba_instr_mem_din0_o[2] ;
 wire \mba_instr_mem_din0_o[30] ;
 wire \mba_instr_mem_din0_o[31] ;
 wire \mba_instr_mem_din0_o[3] ;
 wire \mba_instr_mem_din0_o[4] ;
 wire \mba_instr_mem_din0_o[5] ;
 wire \mba_instr_mem_din0_o[6] ;
 wire \mba_instr_mem_din0_o[7] ;
 wire \mba_instr_mem_din0_o[8] ;
 wire \mba_instr_mem_din0_o[9] ;
 wire \mba_instr_mem_dout0_i[0] ;
 wire \mba_instr_mem_dout0_i[10] ;
 wire \mba_instr_mem_dout0_i[11] ;
 wire \mba_instr_mem_dout0_i[12] ;
 wire \mba_instr_mem_dout0_i[13] ;
 wire \mba_instr_mem_dout0_i[14] ;
 wire \mba_instr_mem_dout0_i[15] ;
 wire \mba_instr_mem_dout0_i[16] ;
 wire \mba_instr_mem_dout0_i[17] ;
 wire \mba_instr_mem_dout0_i[18] ;
 wire \mba_instr_mem_dout0_i[19] ;
 wire \mba_instr_mem_dout0_i[1] ;
 wire \mba_instr_mem_dout0_i[20] ;
 wire \mba_instr_mem_dout0_i[21] ;
 wire \mba_instr_mem_dout0_i[22] ;
 wire \mba_instr_mem_dout0_i[23] ;
 wire \mba_instr_mem_dout0_i[24] ;
 wire \mba_instr_mem_dout0_i[25] ;
 wire \mba_instr_mem_dout0_i[26] ;
 wire \mba_instr_mem_dout0_i[27] ;
 wire \mba_instr_mem_dout0_i[28] ;
 wire \mba_instr_mem_dout0_i[29] ;
 wire \mba_instr_mem_dout0_i[2] ;
 wire \mba_instr_mem_dout0_i[30] ;
 wire \mba_instr_mem_dout0_i[31] ;
 wire \mba_instr_mem_dout0_i[3] ;
 wire \mba_instr_mem_dout0_i[4] ;
 wire \mba_instr_mem_dout0_i[5] ;
 wire \mba_instr_mem_dout0_i[6] ;
 wire \mba_instr_mem_dout0_i[7] ;
 wire \mba_instr_mem_dout0_i[8] ;
 wire \mba_instr_mem_dout0_i[9] ;
 wire mba_instr_mem_web0_o;
 wire \mba_instr_mem_wmask0_o[0] ;
 wire \mba_instr_mem_wmask0_o[1] ;
 wire \mba_instr_mem_wmask0_o[2] ;
 wire \mba_instr_mem_wmask0_o[3] ;
 wire rstn_int;
 wire scan_o;
 wire scl_padoen_o;
 wire sda_padoen_o;
 wire \slaves_00_ar_addr[0] ;
 wire \slaves_00_ar_addr[10] ;
 wire \slaves_00_ar_addr[11] ;
 wire \slaves_00_ar_addr[12] ;
 wire \slaves_00_ar_addr[13] ;
 wire \slaves_00_ar_addr[14] ;
 wire \slaves_00_ar_addr[15] ;
 wire \slaves_00_ar_addr[16] ;
 wire \slaves_00_ar_addr[17] ;
 wire \slaves_00_ar_addr[18] ;
 wire \slaves_00_ar_addr[19] ;
 wire \slaves_00_ar_addr[1] ;
 wire \slaves_00_ar_addr[20] ;
 wire \slaves_00_ar_addr[21] ;
 wire \slaves_00_ar_addr[22] ;
 wire \slaves_00_ar_addr[23] ;
 wire \slaves_00_ar_addr[24] ;
 wire \slaves_00_ar_addr[25] ;
 wire \slaves_00_ar_addr[26] ;
 wire \slaves_00_ar_addr[27] ;
 wire \slaves_00_ar_addr[28] ;
 wire \slaves_00_ar_addr[29] ;
 wire \slaves_00_ar_addr[2] ;
 wire \slaves_00_ar_addr[30] ;
 wire \slaves_00_ar_addr[31] ;
 wire \slaves_00_ar_addr[3] ;
 wire \slaves_00_ar_addr[4] ;
 wire \slaves_00_ar_addr[5] ;
 wire \slaves_00_ar_addr[6] ;
 wire \slaves_00_ar_addr[7] ;
 wire \slaves_00_ar_addr[8] ;
 wire \slaves_00_ar_addr[9] ;
 wire \slaves_00_ar_burst[0] ;
 wire \slaves_00_ar_burst[1] ;
 wire \slaves_00_ar_cache[0] ;
 wire \slaves_00_ar_cache[1] ;
 wire \slaves_00_ar_cache[2] ;
 wire \slaves_00_ar_cache[3] ;
 wire \slaves_00_ar_len[0] ;
 wire \slaves_00_ar_len[1] ;
 wire \slaves_00_ar_len[2] ;
 wire \slaves_00_ar_len[3] ;
 wire \slaves_00_ar_len[4] ;
 wire \slaves_00_ar_len[5] ;
 wire \slaves_00_ar_len[6] ;
 wire \slaves_00_ar_len[7] ;
 wire slaves_00_ar_lock;
 wire \slaves_00_ar_prot[0] ;
 wire \slaves_00_ar_prot[1] ;
 wire \slaves_00_ar_prot[2] ;
 wire \slaves_00_ar_qos[0] ;
 wire \slaves_00_ar_qos[1] ;
 wire \slaves_00_ar_qos[2] ;
 wire \slaves_00_ar_qos[3] ;
 wire slaves_00_ar_ready;
 wire \slaves_00_ar_region[0] ;
 wire \slaves_00_ar_region[1] ;
 wire \slaves_00_ar_region[2] ;
 wire \slaves_00_ar_region[3] ;
 wire \slaves_00_ar_size[0] ;
 wire \slaves_00_ar_size[1] ;
 wire \slaves_00_ar_size[2] ;
 wire slaves_00_ar_valid;
 wire \slaves_00_aw_addr[0] ;
 wire \slaves_00_aw_addr[10] ;
 wire \slaves_00_aw_addr[11] ;
 wire \slaves_00_aw_addr[12] ;
 wire \slaves_00_aw_addr[13] ;
 wire \slaves_00_aw_addr[14] ;
 wire \slaves_00_aw_addr[15] ;
 wire \slaves_00_aw_addr[16] ;
 wire \slaves_00_aw_addr[17] ;
 wire \slaves_00_aw_addr[18] ;
 wire \slaves_00_aw_addr[19] ;
 wire \slaves_00_aw_addr[1] ;
 wire \slaves_00_aw_addr[20] ;
 wire \slaves_00_aw_addr[21] ;
 wire \slaves_00_aw_addr[22] ;
 wire \slaves_00_aw_addr[23] ;
 wire \slaves_00_aw_addr[24] ;
 wire \slaves_00_aw_addr[25] ;
 wire \slaves_00_aw_addr[26] ;
 wire \slaves_00_aw_addr[27] ;
 wire \slaves_00_aw_addr[28] ;
 wire \slaves_00_aw_addr[29] ;
 wire \slaves_00_aw_addr[2] ;
 wire \slaves_00_aw_addr[30] ;
 wire \slaves_00_aw_addr[31] ;
 wire \slaves_00_aw_addr[3] ;
 wire \slaves_00_aw_addr[4] ;
 wire \slaves_00_aw_addr[5] ;
 wire \slaves_00_aw_addr[6] ;
 wire \slaves_00_aw_addr[7] ;
 wire \slaves_00_aw_addr[8] ;
 wire \slaves_00_aw_addr[9] ;
 wire \slaves_00_aw_burst[0] ;
 wire \slaves_00_aw_burst[1] ;
 wire \slaves_00_aw_cache[0] ;
 wire \slaves_00_aw_cache[1] ;
 wire \slaves_00_aw_cache[2] ;
 wire \slaves_00_aw_cache[3] ;
 wire \slaves_00_aw_len[0] ;
 wire \slaves_00_aw_len[1] ;
 wire \slaves_00_aw_len[2] ;
 wire \slaves_00_aw_len[3] ;
 wire \slaves_00_aw_len[4] ;
 wire \slaves_00_aw_len[5] ;
 wire \slaves_00_aw_len[6] ;
 wire \slaves_00_aw_len[7] ;
 wire slaves_00_aw_lock;
 wire \slaves_00_aw_prot[0] ;
 wire \slaves_00_aw_prot[1] ;
 wire \slaves_00_aw_prot[2] ;
 wire \slaves_00_aw_qos[0] ;
 wire \slaves_00_aw_qos[1] ;
 wire \slaves_00_aw_qos[2] ;
 wire \slaves_00_aw_qos[3] ;
 wire slaves_00_aw_ready;
 wire \slaves_00_aw_region[0] ;
 wire \slaves_00_aw_region[1] ;
 wire \slaves_00_aw_region[2] ;
 wire \slaves_00_aw_region[3] ;
 wire \slaves_00_aw_size[0] ;
 wire \slaves_00_aw_size[1] ;
 wire \slaves_00_aw_size[2] ;
 wire slaves_00_aw_valid;
 wire slaves_00_b_ready;
 wire \slaves_00_b_resp[0] ;
 wire \slaves_00_b_resp[1] ;
 wire slaves_00_b_valid;
 wire \slaves_00_r_data[0] ;
 wire \slaves_00_r_data[10] ;
 wire \slaves_00_r_data[11] ;
 wire \slaves_00_r_data[12] ;
 wire \slaves_00_r_data[13] ;
 wire \slaves_00_r_data[14] ;
 wire \slaves_00_r_data[15] ;
 wire \slaves_00_r_data[16] ;
 wire \slaves_00_r_data[17] ;
 wire \slaves_00_r_data[18] ;
 wire \slaves_00_r_data[19] ;
 wire \slaves_00_r_data[1] ;
 wire \slaves_00_r_data[20] ;
 wire \slaves_00_r_data[21] ;
 wire \slaves_00_r_data[22] ;
 wire \slaves_00_r_data[23] ;
 wire \slaves_00_r_data[24] ;
 wire \slaves_00_r_data[25] ;
 wire \slaves_00_r_data[26] ;
 wire \slaves_00_r_data[27] ;
 wire \slaves_00_r_data[28] ;
 wire \slaves_00_r_data[29] ;
 wire \slaves_00_r_data[2] ;
 wire \slaves_00_r_data[30] ;
 wire \slaves_00_r_data[31] ;
 wire \slaves_00_r_data[3] ;
 wire \slaves_00_r_data[4] ;
 wire \slaves_00_r_data[5] ;
 wire \slaves_00_r_data[6] ;
 wire \slaves_00_r_data[7] ;
 wire \slaves_00_r_data[8] ;
 wire \slaves_00_r_data[9] ;
 wire slaves_00_r_last;
 wire slaves_00_r_ready;
 wire \slaves_00_r_resp[0] ;
 wire \slaves_00_r_resp[1] ;
 wire slaves_00_r_valid;
 wire \slaves_00_w_data[0] ;
 wire \slaves_00_w_data[10] ;
 wire \slaves_00_w_data[11] ;
 wire \slaves_00_w_data[12] ;
 wire \slaves_00_w_data[13] ;
 wire \slaves_00_w_data[14] ;
 wire \slaves_00_w_data[15] ;
 wire \slaves_00_w_data[16] ;
 wire \slaves_00_w_data[17] ;
 wire \slaves_00_w_data[18] ;
 wire \slaves_00_w_data[19] ;
 wire \slaves_00_w_data[1] ;
 wire \slaves_00_w_data[20] ;
 wire \slaves_00_w_data[21] ;
 wire \slaves_00_w_data[22] ;
 wire \slaves_00_w_data[23] ;
 wire \slaves_00_w_data[24] ;
 wire \slaves_00_w_data[25] ;
 wire \slaves_00_w_data[26] ;
 wire \slaves_00_w_data[27] ;
 wire \slaves_00_w_data[28] ;
 wire \slaves_00_w_data[29] ;
 wire \slaves_00_w_data[2] ;
 wire \slaves_00_w_data[30] ;
 wire \slaves_00_w_data[31] ;
 wire \slaves_00_w_data[3] ;
 wire \slaves_00_w_data[4] ;
 wire \slaves_00_w_data[5] ;
 wire \slaves_00_w_data[6] ;
 wire \slaves_00_w_data[7] ;
 wire \slaves_00_w_data[8] ;
 wire \slaves_00_w_data[9] ;
 wire slaves_00_w_last;
 wire slaves_00_w_ready;
 wire \slaves_00_w_strb[0] ;
 wire \slaves_00_w_strb[1] ;
 wire \slaves_00_w_strb[2] ;
 wire \slaves_00_w_strb[3] ;
 wire slaves_00_w_valid;
 wire \slaves_01_ar_addr[0] ;
 wire \slaves_01_ar_addr[10] ;
 wire \slaves_01_ar_addr[11] ;
 wire \slaves_01_ar_addr[12] ;
 wire \slaves_01_ar_addr[13] ;
 wire \slaves_01_ar_addr[14] ;
 wire \slaves_01_ar_addr[15] ;
 wire \slaves_01_ar_addr[16] ;
 wire \slaves_01_ar_addr[17] ;
 wire \slaves_01_ar_addr[18] ;
 wire \slaves_01_ar_addr[19] ;
 wire \slaves_01_ar_addr[1] ;
 wire \slaves_01_ar_addr[20] ;
 wire \slaves_01_ar_addr[21] ;
 wire \slaves_01_ar_addr[22] ;
 wire \slaves_01_ar_addr[23] ;
 wire \slaves_01_ar_addr[24] ;
 wire \slaves_01_ar_addr[25] ;
 wire \slaves_01_ar_addr[26] ;
 wire \slaves_01_ar_addr[27] ;
 wire \slaves_01_ar_addr[28] ;
 wire \slaves_01_ar_addr[29] ;
 wire \slaves_01_ar_addr[2] ;
 wire \slaves_01_ar_addr[30] ;
 wire \slaves_01_ar_addr[31] ;
 wire \slaves_01_ar_addr[3] ;
 wire \slaves_01_ar_addr[4] ;
 wire \slaves_01_ar_addr[5] ;
 wire \slaves_01_ar_addr[6] ;
 wire \slaves_01_ar_addr[7] ;
 wire \slaves_01_ar_addr[8] ;
 wire \slaves_01_ar_addr[9] ;
 wire \slaves_01_ar_burst[0] ;
 wire \slaves_01_ar_burst[1] ;
 wire \slaves_01_ar_cache[0] ;
 wire \slaves_01_ar_cache[1] ;
 wire \slaves_01_ar_cache[2] ;
 wire \slaves_01_ar_cache[3] ;
 wire \slaves_01_ar_len[0] ;
 wire \slaves_01_ar_len[1] ;
 wire \slaves_01_ar_len[2] ;
 wire \slaves_01_ar_len[3] ;
 wire \slaves_01_ar_len[4] ;
 wire \slaves_01_ar_len[5] ;
 wire \slaves_01_ar_len[6] ;
 wire \slaves_01_ar_len[7] ;
 wire slaves_01_ar_lock;
 wire \slaves_01_ar_prot[0] ;
 wire \slaves_01_ar_prot[1] ;
 wire \slaves_01_ar_prot[2] ;
 wire \slaves_01_ar_qos[0] ;
 wire \slaves_01_ar_qos[1] ;
 wire \slaves_01_ar_qos[2] ;
 wire \slaves_01_ar_qos[3] ;
 wire slaves_01_ar_ready;
 wire \slaves_01_ar_region[0] ;
 wire \slaves_01_ar_region[1] ;
 wire \slaves_01_ar_region[2] ;
 wire \slaves_01_ar_region[3] ;
 wire \slaves_01_ar_size[0] ;
 wire \slaves_01_ar_size[1] ;
 wire \slaves_01_ar_size[2] ;
 wire slaves_01_ar_valid;
 wire \slaves_01_aw_addr[0] ;
 wire \slaves_01_aw_addr[10] ;
 wire \slaves_01_aw_addr[11] ;
 wire \slaves_01_aw_addr[12] ;
 wire \slaves_01_aw_addr[13] ;
 wire \slaves_01_aw_addr[14] ;
 wire \slaves_01_aw_addr[15] ;
 wire \slaves_01_aw_addr[16] ;
 wire \slaves_01_aw_addr[17] ;
 wire \slaves_01_aw_addr[18] ;
 wire \slaves_01_aw_addr[19] ;
 wire \slaves_01_aw_addr[1] ;
 wire \slaves_01_aw_addr[20] ;
 wire \slaves_01_aw_addr[21] ;
 wire \slaves_01_aw_addr[22] ;
 wire \slaves_01_aw_addr[23] ;
 wire \slaves_01_aw_addr[24] ;
 wire \slaves_01_aw_addr[25] ;
 wire \slaves_01_aw_addr[26] ;
 wire \slaves_01_aw_addr[27] ;
 wire \slaves_01_aw_addr[28] ;
 wire \slaves_01_aw_addr[29] ;
 wire \slaves_01_aw_addr[2] ;
 wire \slaves_01_aw_addr[30] ;
 wire \slaves_01_aw_addr[31] ;
 wire \slaves_01_aw_addr[3] ;
 wire \slaves_01_aw_addr[4] ;
 wire \slaves_01_aw_addr[5] ;
 wire \slaves_01_aw_addr[6] ;
 wire \slaves_01_aw_addr[7] ;
 wire \slaves_01_aw_addr[8] ;
 wire \slaves_01_aw_addr[9] ;
 wire \slaves_01_aw_burst[0] ;
 wire \slaves_01_aw_burst[1] ;
 wire \slaves_01_aw_cache[0] ;
 wire \slaves_01_aw_cache[1] ;
 wire \slaves_01_aw_cache[2] ;
 wire \slaves_01_aw_cache[3] ;
 wire \slaves_01_aw_len[0] ;
 wire \slaves_01_aw_len[1] ;
 wire \slaves_01_aw_len[2] ;
 wire \slaves_01_aw_len[3] ;
 wire \slaves_01_aw_len[4] ;
 wire \slaves_01_aw_len[5] ;
 wire \slaves_01_aw_len[6] ;
 wire \slaves_01_aw_len[7] ;
 wire slaves_01_aw_lock;
 wire \slaves_01_aw_prot[0] ;
 wire \slaves_01_aw_prot[1] ;
 wire \slaves_01_aw_prot[2] ;
 wire \slaves_01_aw_qos[0] ;
 wire \slaves_01_aw_qos[1] ;
 wire \slaves_01_aw_qos[2] ;
 wire \slaves_01_aw_qos[3] ;
 wire slaves_01_aw_ready;
 wire \slaves_01_aw_region[0] ;
 wire \slaves_01_aw_region[1] ;
 wire \slaves_01_aw_region[2] ;
 wire \slaves_01_aw_region[3] ;
 wire \slaves_01_aw_size[0] ;
 wire \slaves_01_aw_size[1] ;
 wire \slaves_01_aw_size[2] ;
 wire slaves_01_aw_valid;
 wire slaves_01_b_ready;
 wire \slaves_01_b_resp[0] ;
 wire \slaves_01_b_resp[1] ;
 wire slaves_01_b_valid;
 wire \slaves_01_r_data[0] ;
 wire \slaves_01_r_data[10] ;
 wire \slaves_01_r_data[11] ;
 wire \slaves_01_r_data[12] ;
 wire \slaves_01_r_data[13] ;
 wire \slaves_01_r_data[14] ;
 wire \slaves_01_r_data[15] ;
 wire \slaves_01_r_data[16] ;
 wire \slaves_01_r_data[17] ;
 wire \slaves_01_r_data[18] ;
 wire \slaves_01_r_data[19] ;
 wire \slaves_01_r_data[1] ;
 wire \slaves_01_r_data[20] ;
 wire \slaves_01_r_data[21] ;
 wire \slaves_01_r_data[22] ;
 wire \slaves_01_r_data[23] ;
 wire \slaves_01_r_data[24] ;
 wire \slaves_01_r_data[25] ;
 wire \slaves_01_r_data[26] ;
 wire \slaves_01_r_data[27] ;
 wire \slaves_01_r_data[28] ;
 wire \slaves_01_r_data[29] ;
 wire \slaves_01_r_data[2] ;
 wire \slaves_01_r_data[30] ;
 wire \slaves_01_r_data[31] ;
 wire \slaves_01_r_data[3] ;
 wire \slaves_01_r_data[4] ;
 wire \slaves_01_r_data[5] ;
 wire \slaves_01_r_data[6] ;
 wire \slaves_01_r_data[7] ;
 wire \slaves_01_r_data[8] ;
 wire \slaves_01_r_data[9] ;
 wire slaves_01_r_last;
 wire slaves_01_r_ready;
 wire \slaves_01_r_resp[0] ;
 wire \slaves_01_r_resp[1] ;
 wire slaves_01_r_valid;
 wire \slaves_01_w_data[0] ;
 wire \slaves_01_w_data[10] ;
 wire \slaves_01_w_data[11] ;
 wire \slaves_01_w_data[12] ;
 wire \slaves_01_w_data[13] ;
 wire \slaves_01_w_data[14] ;
 wire \slaves_01_w_data[15] ;
 wire \slaves_01_w_data[16] ;
 wire \slaves_01_w_data[17] ;
 wire \slaves_01_w_data[18] ;
 wire \slaves_01_w_data[19] ;
 wire \slaves_01_w_data[1] ;
 wire \slaves_01_w_data[20] ;
 wire \slaves_01_w_data[21] ;
 wire \slaves_01_w_data[22] ;
 wire \slaves_01_w_data[23] ;
 wire \slaves_01_w_data[24] ;
 wire \slaves_01_w_data[25] ;
 wire \slaves_01_w_data[26] ;
 wire \slaves_01_w_data[27] ;
 wire \slaves_01_w_data[28] ;
 wire \slaves_01_w_data[29] ;
 wire \slaves_01_w_data[2] ;
 wire \slaves_01_w_data[30] ;
 wire \slaves_01_w_data[31] ;
 wire \slaves_01_w_data[3] ;
 wire \slaves_01_w_data[4] ;
 wire \slaves_01_w_data[5] ;
 wire \slaves_01_w_data[6] ;
 wire \slaves_01_w_data[7] ;
 wire \slaves_01_w_data[8] ;
 wire \slaves_01_w_data[9] ;
 wire slaves_01_w_last;
 wire slaves_01_w_ready;
 wire \slaves_01_w_strb[0] ;
 wire \slaves_01_w_strb[1] ;
 wire \slaves_01_w_strb[2] ;
 wire \slaves_01_w_strb[3] ;
 wire slaves_01_w_valid;
 wire \slaves_02_ar_addr[0] ;
 wire \slaves_02_ar_addr[10] ;
 wire \slaves_02_ar_addr[11] ;
 wire \slaves_02_ar_addr[12] ;
 wire \slaves_02_ar_addr[13] ;
 wire \slaves_02_ar_addr[14] ;
 wire \slaves_02_ar_addr[15] ;
 wire \slaves_02_ar_addr[16] ;
 wire \slaves_02_ar_addr[17] ;
 wire \slaves_02_ar_addr[18] ;
 wire \slaves_02_ar_addr[19] ;
 wire \slaves_02_ar_addr[1] ;
 wire \slaves_02_ar_addr[20] ;
 wire \slaves_02_ar_addr[21] ;
 wire \slaves_02_ar_addr[22] ;
 wire \slaves_02_ar_addr[23] ;
 wire \slaves_02_ar_addr[24] ;
 wire \slaves_02_ar_addr[25] ;
 wire \slaves_02_ar_addr[26] ;
 wire \slaves_02_ar_addr[27] ;
 wire \slaves_02_ar_addr[28] ;
 wire \slaves_02_ar_addr[29] ;
 wire \slaves_02_ar_addr[2] ;
 wire \slaves_02_ar_addr[30] ;
 wire \slaves_02_ar_addr[31] ;
 wire \slaves_02_ar_addr[3] ;
 wire \slaves_02_ar_addr[4] ;
 wire \slaves_02_ar_addr[5] ;
 wire \slaves_02_ar_addr[6] ;
 wire \slaves_02_ar_addr[7] ;
 wire \slaves_02_ar_addr[8] ;
 wire \slaves_02_ar_addr[9] ;
 wire \slaves_02_ar_burst[0] ;
 wire \slaves_02_ar_burst[1] ;
 wire \slaves_02_ar_cache[0] ;
 wire \slaves_02_ar_cache[1] ;
 wire \slaves_02_ar_cache[2] ;
 wire \slaves_02_ar_cache[3] ;
 wire \slaves_02_ar_len[0] ;
 wire \slaves_02_ar_len[1] ;
 wire \slaves_02_ar_len[2] ;
 wire \slaves_02_ar_len[3] ;
 wire \slaves_02_ar_len[4] ;
 wire \slaves_02_ar_len[5] ;
 wire \slaves_02_ar_len[6] ;
 wire \slaves_02_ar_len[7] ;
 wire slaves_02_ar_lock;
 wire \slaves_02_ar_prot[0] ;
 wire \slaves_02_ar_prot[1] ;
 wire \slaves_02_ar_prot[2] ;
 wire \slaves_02_ar_qos[0] ;
 wire \slaves_02_ar_qos[1] ;
 wire \slaves_02_ar_qos[2] ;
 wire \slaves_02_ar_qos[3] ;
 wire slaves_02_ar_ready;
 wire \slaves_02_ar_region[0] ;
 wire \slaves_02_ar_region[1] ;
 wire \slaves_02_ar_region[2] ;
 wire \slaves_02_ar_region[3] ;
 wire \slaves_02_ar_size[0] ;
 wire \slaves_02_ar_size[1] ;
 wire \slaves_02_ar_size[2] ;
 wire slaves_02_ar_valid;
 wire \slaves_02_aw_addr[0] ;
 wire \slaves_02_aw_addr[10] ;
 wire \slaves_02_aw_addr[11] ;
 wire \slaves_02_aw_addr[12] ;
 wire \slaves_02_aw_addr[13] ;
 wire \slaves_02_aw_addr[14] ;
 wire \slaves_02_aw_addr[15] ;
 wire \slaves_02_aw_addr[16] ;
 wire \slaves_02_aw_addr[17] ;
 wire \slaves_02_aw_addr[18] ;
 wire \slaves_02_aw_addr[19] ;
 wire \slaves_02_aw_addr[1] ;
 wire \slaves_02_aw_addr[20] ;
 wire \slaves_02_aw_addr[21] ;
 wire \slaves_02_aw_addr[22] ;
 wire \slaves_02_aw_addr[23] ;
 wire \slaves_02_aw_addr[24] ;
 wire \slaves_02_aw_addr[25] ;
 wire \slaves_02_aw_addr[26] ;
 wire \slaves_02_aw_addr[27] ;
 wire \slaves_02_aw_addr[28] ;
 wire \slaves_02_aw_addr[29] ;
 wire \slaves_02_aw_addr[2] ;
 wire \slaves_02_aw_addr[30] ;
 wire \slaves_02_aw_addr[31] ;
 wire \slaves_02_aw_addr[3] ;
 wire \slaves_02_aw_addr[4] ;
 wire \slaves_02_aw_addr[5] ;
 wire \slaves_02_aw_addr[6] ;
 wire \slaves_02_aw_addr[7] ;
 wire \slaves_02_aw_addr[8] ;
 wire \slaves_02_aw_addr[9] ;
 wire \slaves_02_aw_burst[0] ;
 wire \slaves_02_aw_burst[1] ;
 wire \slaves_02_aw_cache[0] ;
 wire \slaves_02_aw_cache[1] ;
 wire \slaves_02_aw_cache[2] ;
 wire \slaves_02_aw_cache[3] ;
 wire \slaves_02_aw_len[0] ;
 wire \slaves_02_aw_len[1] ;
 wire \slaves_02_aw_len[2] ;
 wire \slaves_02_aw_len[3] ;
 wire \slaves_02_aw_len[4] ;
 wire \slaves_02_aw_len[5] ;
 wire \slaves_02_aw_len[6] ;
 wire \slaves_02_aw_len[7] ;
 wire slaves_02_aw_lock;
 wire \slaves_02_aw_prot[0] ;
 wire \slaves_02_aw_prot[1] ;
 wire \slaves_02_aw_prot[2] ;
 wire \slaves_02_aw_qos[0] ;
 wire \slaves_02_aw_qos[1] ;
 wire \slaves_02_aw_qos[2] ;
 wire \slaves_02_aw_qos[3] ;
 wire slaves_02_aw_ready;
 wire \slaves_02_aw_region[0] ;
 wire \slaves_02_aw_region[1] ;
 wire \slaves_02_aw_region[2] ;
 wire \slaves_02_aw_region[3] ;
 wire \slaves_02_aw_size[0] ;
 wire \slaves_02_aw_size[1] ;
 wire \slaves_02_aw_size[2] ;
 wire slaves_02_aw_valid;
 wire slaves_02_b_ready;
 wire \slaves_02_b_resp[0] ;
 wire \slaves_02_b_resp[1] ;
 wire slaves_02_b_valid;
 wire \slaves_02_r_data[0] ;
 wire \slaves_02_r_data[10] ;
 wire \slaves_02_r_data[11] ;
 wire \slaves_02_r_data[12] ;
 wire \slaves_02_r_data[13] ;
 wire \slaves_02_r_data[14] ;
 wire \slaves_02_r_data[15] ;
 wire \slaves_02_r_data[16] ;
 wire \slaves_02_r_data[17] ;
 wire \slaves_02_r_data[18] ;
 wire \slaves_02_r_data[19] ;
 wire \slaves_02_r_data[1] ;
 wire \slaves_02_r_data[20] ;
 wire \slaves_02_r_data[21] ;
 wire \slaves_02_r_data[22] ;
 wire \slaves_02_r_data[23] ;
 wire \slaves_02_r_data[24] ;
 wire \slaves_02_r_data[25] ;
 wire \slaves_02_r_data[26] ;
 wire \slaves_02_r_data[27] ;
 wire \slaves_02_r_data[28] ;
 wire \slaves_02_r_data[29] ;
 wire \slaves_02_r_data[2] ;
 wire \slaves_02_r_data[30] ;
 wire \slaves_02_r_data[31] ;
 wire \slaves_02_r_data[3] ;
 wire \slaves_02_r_data[4] ;
 wire \slaves_02_r_data[5] ;
 wire \slaves_02_r_data[6] ;
 wire \slaves_02_r_data[7] ;
 wire \slaves_02_r_data[8] ;
 wire \slaves_02_r_data[9] ;
 wire slaves_02_r_last;
 wire slaves_02_r_ready;
 wire \slaves_02_r_resp[0] ;
 wire \slaves_02_r_resp[1] ;
 wire slaves_02_r_valid;
 wire \slaves_02_w_data[0] ;
 wire \slaves_02_w_data[10] ;
 wire \slaves_02_w_data[11] ;
 wire \slaves_02_w_data[12] ;
 wire \slaves_02_w_data[13] ;
 wire \slaves_02_w_data[14] ;
 wire \slaves_02_w_data[15] ;
 wire \slaves_02_w_data[16] ;
 wire \slaves_02_w_data[17] ;
 wire \slaves_02_w_data[18] ;
 wire \slaves_02_w_data[19] ;
 wire \slaves_02_w_data[1] ;
 wire \slaves_02_w_data[20] ;
 wire \slaves_02_w_data[21] ;
 wire \slaves_02_w_data[22] ;
 wire \slaves_02_w_data[23] ;
 wire \slaves_02_w_data[24] ;
 wire \slaves_02_w_data[25] ;
 wire \slaves_02_w_data[26] ;
 wire \slaves_02_w_data[27] ;
 wire \slaves_02_w_data[28] ;
 wire \slaves_02_w_data[29] ;
 wire \slaves_02_w_data[2] ;
 wire \slaves_02_w_data[30] ;
 wire \slaves_02_w_data[31] ;
 wire \slaves_02_w_data[3] ;
 wire \slaves_02_w_data[4] ;
 wire \slaves_02_w_data[5] ;
 wire \slaves_02_w_data[6] ;
 wire \slaves_02_w_data[7] ;
 wire \slaves_02_w_data[8] ;
 wire \slaves_02_w_data[9] ;
 wire slaves_02_w_last;
 wire slaves_02_w_ready;
 wire \slaves_02_w_strb[0] ;
 wire \slaves_02_w_strb[1] ;
 wire \slaves_02_w_strb[2] ;
 wire \slaves_02_w_strb[3] ;
 wire slaves_02_w_valid;
 wire spi_master_csn1;
 wire spi_master_csn2;
 wire spi_master_csn3;
 wire spi_master_sdo1;
 wire spi_master_sdo2;
 wire spi_master_sdo3;
 wire spi_sdo1_o;
 wire spi_sdo2_o;
 wire spi_sdo3_o;
 wire uart_dtr;
 wire uart_rts;

 axi_node_intf_wrap axi_interconnect_i (.clk(clk_int),
    .m00_ar_lock(slaves_00_ar_lock),
    .m00_ar_ready(slaves_00_ar_ready),
    .m00_ar_valid(slaves_00_ar_valid),
    .m00_aw_lock(slaves_00_aw_lock),
    .m00_aw_ready(slaves_00_aw_ready),
    .m00_aw_valid(slaves_00_aw_valid),
    .m00_b_ready(slaves_00_b_ready),
    .m00_b_valid(slaves_00_b_valid),
    .m00_r_last(slaves_00_r_last),
    .m00_r_ready(slaves_00_r_ready),
    .m00_r_valid(slaves_00_r_valid),
    .m00_w_last(slaves_00_w_last),
    .m00_w_ready(slaves_00_w_ready),
    .m00_w_valid(slaves_00_w_valid),
    .m01_ar_lock(slaves_01_ar_lock),
    .m01_ar_ready(slaves_01_ar_ready),
    .m01_ar_valid(slaves_01_ar_valid),
    .m01_aw_lock(slaves_01_aw_lock),
    .m01_aw_ready(slaves_01_aw_ready),
    .m01_aw_valid(slaves_01_aw_valid),
    .m01_b_ready(slaves_01_b_ready),
    .m01_b_valid(slaves_01_b_valid),
    .m01_r_last(slaves_01_r_last),
    .m01_r_ready(slaves_01_r_ready),
    .m01_r_valid(slaves_01_r_valid),
    .m01_w_last(slaves_01_w_last),
    .m01_w_ready(slaves_01_w_ready),
    .m01_w_valid(slaves_01_w_valid),
    .m02_ar_lock(slaves_02_ar_lock),
    .m02_ar_ready(slaves_02_ar_ready),
    .m02_ar_valid(slaves_02_ar_valid),
    .m02_aw_lock(slaves_02_aw_lock),
    .m02_aw_ready(slaves_02_aw_ready),
    .m02_aw_valid(slaves_02_aw_valid),
    .m02_b_ready(slaves_02_b_ready),
    .m02_b_valid(slaves_02_b_valid),
    .m02_r_last(slaves_02_r_last),
    .m02_r_ready(slaves_02_r_ready),
    .m02_r_valid(slaves_02_r_valid),
    .m02_w_last(slaves_02_w_last),
    .m02_w_ready(slaves_02_w_ready),
    .m02_w_valid(slaves_02_w_valid),
    .rst_n(rstn_int),
    .s00_ar_lock(masters_00_ar_lock),
    .s00_ar_ready(masters_00_ar_ready),
    .s00_ar_valid(masters_00_ar_valid),
    .s00_aw_lock(masters_00_aw_lock),
    .s00_aw_ready(masters_00_aw_ready),
    .s00_aw_valid(masters_00_aw_valid),
    .s00_b_ready(masters_00_b_ready),
    .s00_b_valid(masters_00_b_valid),
    .s00_r_last(masters_00_r_last),
    .s00_r_ready(masters_00_r_ready),
    .s00_r_valid(masters_00_r_valid),
    .s00_w_last(masters_00_w_last),
    .s00_w_ready(masters_00_w_ready),
    .s00_w_valid(masters_00_w_valid),
    .s01_ar_lock(masters_01_ar_lock),
    .s01_ar_ready(masters_01_ar_ready),
    .s01_ar_valid(masters_01_ar_valid),
    .s01_aw_lock(masters_01_aw_lock),
    .s01_aw_ready(masters_01_aw_ready),
    .s01_aw_valid(masters_01_aw_valid),
    .s01_b_ready(masters_01_b_ready),
    .s01_b_valid(masters_01_b_valid),
    .s01_r_last(masters_01_r_last),
    .s01_r_ready(masters_01_r_ready),
    .s01_r_valid(masters_01_r_valid),
    .s01_w_last(masters_01_w_last),
    .s01_w_ready(masters_01_w_ready),
    .s01_w_valid(masters_01_w_valid),
    .s02_ar_lock(masters_02_ar_lock),
    .s02_ar_ready(masters_02_ar_ready),
    .s02_ar_valid(masters_02_ar_valid),
    .s02_aw_lock(masters_02_aw_lock),
    .s02_aw_ready(masters_02_aw_ready),
    .s02_aw_valid(masters_02_aw_valid),
    .s02_b_ready(masters_02_b_ready),
    .s02_b_valid(masters_02_b_valid),
    .s02_r_last(masters_02_r_last),
    .s02_r_ready(masters_02_r_ready),
    .s02_r_valid(masters_02_r_valid),
    .s02_w_last(masters_02_w_last),
    .s02_w_ready(masters_02_w_ready),
    .s02_w_valid(masters_02_w_valid),
    .test_en_i(la_data_in[2]),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .m00_ar_addr({\slaves_00_ar_addr[31] ,
    \slaves_00_ar_addr[30] ,
    \slaves_00_ar_addr[29] ,
    \slaves_00_ar_addr[28] ,
    \slaves_00_ar_addr[27] ,
    \slaves_00_ar_addr[26] ,
    \slaves_00_ar_addr[25] ,
    \slaves_00_ar_addr[24] ,
    \slaves_00_ar_addr[23] ,
    \slaves_00_ar_addr[22] ,
    \slaves_00_ar_addr[21] ,
    \slaves_00_ar_addr[20] ,
    \slaves_00_ar_addr[19] ,
    \slaves_00_ar_addr[18] ,
    \slaves_00_ar_addr[17] ,
    \slaves_00_ar_addr[16] ,
    \slaves_00_ar_addr[15] ,
    \slaves_00_ar_addr[14] ,
    \slaves_00_ar_addr[13] ,
    \slaves_00_ar_addr[12] ,
    \slaves_00_ar_addr[11] ,
    \slaves_00_ar_addr[10] ,
    \slaves_00_ar_addr[9] ,
    \slaves_00_ar_addr[8] ,
    \slaves_00_ar_addr[7] ,
    \slaves_00_ar_addr[6] ,
    \slaves_00_ar_addr[5] ,
    \slaves_00_ar_addr[4] ,
    \slaves_00_ar_addr[3] ,
    \slaves_00_ar_addr[2] ,
    \slaves_00_ar_addr[1] ,
    \slaves_00_ar_addr[0] }),
    .m00_ar_burst({\slaves_00_ar_burst[1] ,
    \slaves_00_ar_burst[0] }),
    .m00_ar_cache({\slaves_00_ar_cache[3] ,
    \slaves_00_ar_cache[2] ,
    \slaves_00_ar_cache[1] ,
    \slaves_00_ar_cache[0] }),
    .m00_ar_id({_NC1,
    _NC2,
    _NC3,
    _NC4,
    _NC5,
    _NC6,
    _NC7,
    _NC8,
    _NC9,
    _NC10,
    _NC11,
    _NC12}),
    .m00_ar_len({\slaves_00_ar_len[7] ,
    \slaves_00_ar_len[6] ,
    \slaves_00_ar_len[5] ,
    \slaves_00_ar_len[4] ,
    \slaves_00_ar_len[3] ,
    \slaves_00_ar_len[2] ,
    \slaves_00_ar_len[1] ,
    \slaves_00_ar_len[0] }),
    .m00_ar_prot({\slaves_00_ar_prot[2] ,
    \slaves_00_ar_prot[1] ,
    \slaves_00_ar_prot[0] }),
    .m00_ar_qos({\slaves_00_ar_qos[3] ,
    \slaves_00_ar_qos[2] ,
    \slaves_00_ar_qos[1] ,
    \slaves_00_ar_qos[0] }),
    .m00_ar_region({\slaves_00_ar_region[3] ,
    \slaves_00_ar_region[2] ,
    \slaves_00_ar_region[1] ,
    \slaves_00_ar_region[0] }),
    .m00_ar_size({\slaves_00_ar_size[2] ,
    \slaves_00_ar_size[1] ,
    \slaves_00_ar_size[0] }),
    .m00_ar_user({_NC13,
    _NC14}),
    .m00_aw_addr({\slaves_00_aw_addr[31] ,
    \slaves_00_aw_addr[30] ,
    \slaves_00_aw_addr[29] ,
    \slaves_00_aw_addr[28] ,
    \slaves_00_aw_addr[27] ,
    \slaves_00_aw_addr[26] ,
    \slaves_00_aw_addr[25] ,
    \slaves_00_aw_addr[24] ,
    \slaves_00_aw_addr[23] ,
    \slaves_00_aw_addr[22] ,
    \slaves_00_aw_addr[21] ,
    \slaves_00_aw_addr[20] ,
    \slaves_00_aw_addr[19] ,
    \slaves_00_aw_addr[18] ,
    \slaves_00_aw_addr[17] ,
    \slaves_00_aw_addr[16] ,
    \slaves_00_aw_addr[15] ,
    \slaves_00_aw_addr[14] ,
    \slaves_00_aw_addr[13] ,
    \slaves_00_aw_addr[12] ,
    \slaves_00_aw_addr[11] ,
    \slaves_00_aw_addr[10] ,
    \slaves_00_aw_addr[9] ,
    \slaves_00_aw_addr[8] ,
    \slaves_00_aw_addr[7] ,
    \slaves_00_aw_addr[6] ,
    \slaves_00_aw_addr[5] ,
    \slaves_00_aw_addr[4] ,
    \slaves_00_aw_addr[3] ,
    \slaves_00_aw_addr[2] ,
    \slaves_00_aw_addr[1] ,
    \slaves_00_aw_addr[0] }),
    .m00_aw_burst({\slaves_00_aw_burst[1] ,
    \slaves_00_aw_burst[0] }),
    .m00_aw_cache({\slaves_00_aw_cache[3] ,
    \slaves_00_aw_cache[2] ,
    \slaves_00_aw_cache[1] ,
    \slaves_00_aw_cache[0] }),
    .m00_aw_id({_NC15,
    _NC16,
    _NC17,
    _NC18,
    _NC19,
    _NC20,
    _NC21,
    _NC22,
    _NC23,
    _NC24,
    _NC25,
    _NC26}),
    .m00_aw_len({\slaves_00_aw_len[7] ,
    \slaves_00_aw_len[6] ,
    \slaves_00_aw_len[5] ,
    \slaves_00_aw_len[4] ,
    \slaves_00_aw_len[3] ,
    \slaves_00_aw_len[2] ,
    \slaves_00_aw_len[1] ,
    \slaves_00_aw_len[0] }),
    .m00_aw_prot({\slaves_00_aw_prot[2] ,
    \slaves_00_aw_prot[1] ,
    \slaves_00_aw_prot[0] }),
    .m00_aw_qos({\slaves_00_aw_qos[3] ,
    \slaves_00_aw_qos[2] ,
    \slaves_00_aw_qos[1] ,
    \slaves_00_aw_qos[0] }),
    .m00_aw_region({\slaves_00_aw_region[3] ,
    \slaves_00_aw_region[2] ,
    \slaves_00_aw_region[1] ,
    \slaves_00_aw_region[0] }),
    .m00_aw_size({\slaves_00_aw_size[2] ,
    \slaves_00_aw_size[1] ,
    \slaves_00_aw_size[0] }),
    .m00_aw_user({_NC27,
    _NC28}),
    .m00_b_id({_NC29,
    _NC30,
    _NC31,
    _NC32,
    _NC33,
    _NC34,
    _NC35,
    _NC36,
    _NC37,
    _NC38,
    _NC39,
    _NC40}),
    .m00_b_resp({\slaves_00_b_resp[1] ,
    \slaves_00_b_resp[0] }),
    .m00_b_user({_NC41,
    _NC42}),
    .m00_r_data({\slaves_00_r_data[31] ,
    \slaves_00_r_data[30] ,
    \slaves_00_r_data[29] ,
    \slaves_00_r_data[28] ,
    \slaves_00_r_data[27] ,
    \slaves_00_r_data[26] ,
    \slaves_00_r_data[25] ,
    \slaves_00_r_data[24] ,
    \slaves_00_r_data[23] ,
    \slaves_00_r_data[22] ,
    \slaves_00_r_data[21] ,
    \slaves_00_r_data[20] ,
    \slaves_00_r_data[19] ,
    \slaves_00_r_data[18] ,
    \slaves_00_r_data[17] ,
    \slaves_00_r_data[16] ,
    \slaves_00_r_data[15] ,
    \slaves_00_r_data[14] ,
    \slaves_00_r_data[13] ,
    \slaves_00_r_data[12] ,
    \slaves_00_r_data[11] ,
    \slaves_00_r_data[10] ,
    \slaves_00_r_data[9] ,
    \slaves_00_r_data[8] ,
    \slaves_00_r_data[7] ,
    \slaves_00_r_data[6] ,
    \slaves_00_r_data[5] ,
    \slaves_00_r_data[4] ,
    \slaves_00_r_data[3] ,
    \slaves_00_r_data[2] ,
    \slaves_00_r_data[1] ,
    \slaves_00_r_data[0] }),
    .m00_r_id({_NC43,
    _NC44,
    _NC45,
    _NC46,
    _NC47,
    _NC48,
    _NC49,
    _NC50,
    _NC51,
    _NC52,
    _NC53,
    _NC54}),
    .m00_r_resp({\slaves_00_r_resp[1] ,
    \slaves_00_r_resp[0] }),
    .m00_r_user({_NC55,
    _NC56}),
    .m00_w_data({\slaves_00_w_data[31] ,
    \slaves_00_w_data[30] ,
    \slaves_00_w_data[29] ,
    \slaves_00_w_data[28] ,
    \slaves_00_w_data[27] ,
    \slaves_00_w_data[26] ,
    \slaves_00_w_data[25] ,
    \slaves_00_w_data[24] ,
    \slaves_00_w_data[23] ,
    \slaves_00_w_data[22] ,
    \slaves_00_w_data[21] ,
    \slaves_00_w_data[20] ,
    \slaves_00_w_data[19] ,
    \slaves_00_w_data[18] ,
    \slaves_00_w_data[17] ,
    \slaves_00_w_data[16] ,
    \slaves_00_w_data[15] ,
    \slaves_00_w_data[14] ,
    \slaves_00_w_data[13] ,
    \slaves_00_w_data[12] ,
    \slaves_00_w_data[11] ,
    \slaves_00_w_data[10] ,
    \slaves_00_w_data[9] ,
    \slaves_00_w_data[8] ,
    \slaves_00_w_data[7] ,
    \slaves_00_w_data[6] ,
    \slaves_00_w_data[5] ,
    \slaves_00_w_data[4] ,
    \slaves_00_w_data[3] ,
    \slaves_00_w_data[2] ,
    \slaves_00_w_data[1] ,
    \slaves_00_w_data[0] }),
    .m00_w_strb({\slaves_00_w_strb[3] ,
    \slaves_00_w_strb[2] ,
    \slaves_00_w_strb[1] ,
    \slaves_00_w_strb[0] }),
    .m00_w_user({_NC57,
    _NC58}),
    .m01_ar_addr({\slaves_01_ar_addr[31] ,
    \slaves_01_ar_addr[30] ,
    \slaves_01_ar_addr[29] ,
    \slaves_01_ar_addr[28] ,
    \slaves_01_ar_addr[27] ,
    \slaves_01_ar_addr[26] ,
    \slaves_01_ar_addr[25] ,
    \slaves_01_ar_addr[24] ,
    \slaves_01_ar_addr[23] ,
    \slaves_01_ar_addr[22] ,
    \slaves_01_ar_addr[21] ,
    \slaves_01_ar_addr[20] ,
    \slaves_01_ar_addr[19] ,
    \slaves_01_ar_addr[18] ,
    \slaves_01_ar_addr[17] ,
    \slaves_01_ar_addr[16] ,
    \slaves_01_ar_addr[15] ,
    \slaves_01_ar_addr[14] ,
    \slaves_01_ar_addr[13] ,
    \slaves_01_ar_addr[12] ,
    \slaves_01_ar_addr[11] ,
    \slaves_01_ar_addr[10] ,
    \slaves_01_ar_addr[9] ,
    \slaves_01_ar_addr[8] ,
    \slaves_01_ar_addr[7] ,
    \slaves_01_ar_addr[6] ,
    \slaves_01_ar_addr[5] ,
    \slaves_01_ar_addr[4] ,
    \slaves_01_ar_addr[3] ,
    \slaves_01_ar_addr[2] ,
    \slaves_01_ar_addr[1] ,
    \slaves_01_ar_addr[0] }),
    .m01_ar_burst({\slaves_01_ar_burst[1] ,
    \slaves_01_ar_burst[0] }),
    .m01_ar_cache({\slaves_01_ar_cache[3] ,
    \slaves_01_ar_cache[2] ,
    \slaves_01_ar_cache[1] ,
    \slaves_01_ar_cache[0] }),
    .m01_ar_id({_NC59,
    _NC60,
    _NC61,
    _NC62,
    _NC63,
    _NC64,
    _NC65,
    _NC66,
    _NC67,
    _NC68,
    _NC69,
    _NC70}),
    .m01_ar_len({\slaves_01_ar_len[7] ,
    \slaves_01_ar_len[6] ,
    \slaves_01_ar_len[5] ,
    \slaves_01_ar_len[4] ,
    \slaves_01_ar_len[3] ,
    \slaves_01_ar_len[2] ,
    \slaves_01_ar_len[1] ,
    \slaves_01_ar_len[0] }),
    .m01_ar_prot({\slaves_01_ar_prot[2] ,
    \slaves_01_ar_prot[1] ,
    \slaves_01_ar_prot[0] }),
    .m01_ar_qos({\slaves_01_ar_qos[3] ,
    \slaves_01_ar_qos[2] ,
    \slaves_01_ar_qos[1] ,
    \slaves_01_ar_qos[0] }),
    .m01_ar_region({\slaves_01_ar_region[3] ,
    \slaves_01_ar_region[2] ,
    \slaves_01_ar_region[1] ,
    \slaves_01_ar_region[0] }),
    .m01_ar_size({\slaves_01_ar_size[2] ,
    \slaves_01_ar_size[1] ,
    \slaves_01_ar_size[0] }),
    .m01_ar_user({_NC71,
    _NC72}),
    .m01_aw_addr({\slaves_01_aw_addr[31] ,
    \slaves_01_aw_addr[30] ,
    \slaves_01_aw_addr[29] ,
    \slaves_01_aw_addr[28] ,
    \slaves_01_aw_addr[27] ,
    \slaves_01_aw_addr[26] ,
    \slaves_01_aw_addr[25] ,
    \slaves_01_aw_addr[24] ,
    \slaves_01_aw_addr[23] ,
    \slaves_01_aw_addr[22] ,
    \slaves_01_aw_addr[21] ,
    \slaves_01_aw_addr[20] ,
    \slaves_01_aw_addr[19] ,
    \slaves_01_aw_addr[18] ,
    \slaves_01_aw_addr[17] ,
    \slaves_01_aw_addr[16] ,
    \slaves_01_aw_addr[15] ,
    \slaves_01_aw_addr[14] ,
    \slaves_01_aw_addr[13] ,
    \slaves_01_aw_addr[12] ,
    \slaves_01_aw_addr[11] ,
    \slaves_01_aw_addr[10] ,
    \slaves_01_aw_addr[9] ,
    \slaves_01_aw_addr[8] ,
    \slaves_01_aw_addr[7] ,
    \slaves_01_aw_addr[6] ,
    \slaves_01_aw_addr[5] ,
    \slaves_01_aw_addr[4] ,
    \slaves_01_aw_addr[3] ,
    \slaves_01_aw_addr[2] ,
    \slaves_01_aw_addr[1] ,
    \slaves_01_aw_addr[0] }),
    .m01_aw_burst({\slaves_01_aw_burst[1] ,
    \slaves_01_aw_burst[0] }),
    .m01_aw_cache({\slaves_01_aw_cache[3] ,
    \slaves_01_aw_cache[2] ,
    \slaves_01_aw_cache[1] ,
    \slaves_01_aw_cache[0] }),
    .m01_aw_id({_NC73,
    _NC74,
    _NC75,
    _NC76,
    _NC77,
    _NC78,
    _NC79,
    _NC80,
    _NC81,
    _NC82,
    _NC83,
    _NC84}),
    .m01_aw_len({\slaves_01_aw_len[7] ,
    \slaves_01_aw_len[6] ,
    \slaves_01_aw_len[5] ,
    \slaves_01_aw_len[4] ,
    \slaves_01_aw_len[3] ,
    \slaves_01_aw_len[2] ,
    \slaves_01_aw_len[1] ,
    \slaves_01_aw_len[0] }),
    .m01_aw_prot({\slaves_01_aw_prot[2] ,
    \slaves_01_aw_prot[1] ,
    \slaves_01_aw_prot[0] }),
    .m01_aw_qos({\slaves_01_aw_qos[3] ,
    \slaves_01_aw_qos[2] ,
    \slaves_01_aw_qos[1] ,
    \slaves_01_aw_qos[0] }),
    .m01_aw_region({\slaves_01_aw_region[3] ,
    \slaves_01_aw_region[2] ,
    \slaves_01_aw_region[1] ,
    \slaves_01_aw_region[0] }),
    .m01_aw_size({\slaves_01_aw_size[2] ,
    \slaves_01_aw_size[1] ,
    \slaves_01_aw_size[0] }),
    .m01_aw_user({_NC85,
    _NC86}),
    .m01_b_id({_NC87,
    _NC88,
    _NC89,
    _NC90,
    _NC91,
    _NC92,
    _NC93,
    _NC94,
    _NC95,
    _NC96,
    _NC97,
    _NC98}),
    .m01_b_resp({\slaves_01_b_resp[1] ,
    \slaves_01_b_resp[0] }),
    .m01_b_user({_NC99,
    _NC100}),
    .m01_r_data({\slaves_01_r_data[31] ,
    \slaves_01_r_data[30] ,
    \slaves_01_r_data[29] ,
    \slaves_01_r_data[28] ,
    \slaves_01_r_data[27] ,
    \slaves_01_r_data[26] ,
    \slaves_01_r_data[25] ,
    \slaves_01_r_data[24] ,
    \slaves_01_r_data[23] ,
    \slaves_01_r_data[22] ,
    \slaves_01_r_data[21] ,
    \slaves_01_r_data[20] ,
    \slaves_01_r_data[19] ,
    \slaves_01_r_data[18] ,
    \slaves_01_r_data[17] ,
    \slaves_01_r_data[16] ,
    \slaves_01_r_data[15] ,
    \slaves_01_r_data[14] ,
    \slaves_01_r_data[13] ,
    \slaves_01_r_data[12] ,
    \slaves_01_r_data[11] ,
    \slaves_01_r_data[10] ,
    \slaves_01_r_data[9] ,
    \slaves_01_r_data[8] ,
    \slaves_01_r_data[7] ,
    \slaves_01_r_data[6] ,
    \slaves_01_r_data[5] ,
    \slaves_01_r_data[4] ,
    \slaves_01_r_data[3] ,
    \slaves_01_r_data[2] ,
    \slaves_01_r_data[1] ,
    \slaves_01_r_data[0] }),
    .m01_r_id({_NC101,
    _NC102,
    _NC103,
    _NC104,
    _NC105,
    _NC106,
    _NC107,
    _NC108,
    _NC109,
    _NC110,
    _NC111,
    _NC112}),
    .m01_r_resp({\slaves_01_r_resp[1] ,
    \slaves_01_r_resp[0] }),
    .m01_r_user({_NC113,
    _NC114}),
    .m01_w_data({\slaves_01_w_data[31] ,
    \slaves_01_w_data[30] ,
    \slaves_01_w_data[29] ,
    \slaves_01_w_data[28] ,
    \slaves_01_w_data[27] ,
    \slaves_01_w_data[26] ,
    \slaves_01_w_data[25] ,
    \slaves_01_w_data[24] ,
    \slaves_01_w_data[23] ,
    \slaves_01_w_data[22] ,
    \slaves_01_w_data[21] ,
    \slaves_01_w_data[20] ,
    \slaves_01_w_data[19] ,
    \slaves_01_w_data[18] ,
    \slaves_01_w_data[17] ,
    \slaves_01_w_data[16] ,
    \slaves_01_w_data[15] ,
    \slaves_01_w_data[14] ,
    \slaves_01_w_data[13] ,
    \slaves_01_w_data[12] ,
    \slaves_01_w_data[11] ,
    \slaves_01_w_data[10] ,
    \slaves_01_w_data[9] ,
    \slaves_01_w_data[8] ,
    \slaves_01_w_data[7] ,
    \slaves_01_w_data[6] ,
    \slaves_01_w_data[5] ,
    \slaves_01_w_data[4] ,
    \slaves_01_w_data[3] ,
    \slaves_01_w_data[2] ,
    \slaves_01_w_data[1] ,
    \slaves_01_w_data[0] }),
    .m01_w_strb({\slaves_01_w_strb[3] ,
    \slaves_01_w_strb[2] ,
    \slaves_01_w_strb[1] ,
    \slaves_01_w_strb[0] }),
    .m01_w_user({_NC115,
    _NC116}),
    .m02_ar_addr({\slaves_02_ar_addr[31] ,
    \slaves_02_ar_addr[30] ,
    \slaves_02_ar_addr[29] ,
    \slaves_02_ar_addr[28] ,
    \slaves_02_ar_addr[27] ,
    \slaves_02_ar_addr[26] ,
    \slaves_02_ar_addr[25] ,
    \slaves_02_ar_addr[24] ,
    \slaves_02_ar_addr[23] ,
    \slaves_02_ar_addr[22] ,
    \slaves_02_ar_addr[21] ,
    \slaves_02_ar_addr[20] ,
    \slaves_02_ar_addr[19] ,
    \slaves_02_ar_addr[18] ,
    \slaves_02_ar_addr[17] ,
    \slaves_02_ar_addr[16] ,
    \slaves_02_ar_addr[15] ,
    \slaves_02_ar_addr[14] ,
    \slaves_02_ar_addr[13] ,
    \slaves_02_ar_addr[12] ,
    \slaves_02_ar_addr[11] ,
    \slaves_02_ar_addr[10] ,
    \slaves_02_ar_addr[9] ,
    \slaves_02_ar_addr[8] ,
    \slaves_02_ar_addr[7] ,
    \slaves_02_ar_addr[6] ,
    \slaves_02_ar_addr[5] ,
    \slaves_02_ar_addr[4] ,
    \slaves_02_ar_addr[3] ,
    \slaves_02_ar_addr[2] ,
    \slaves_02_ar_addr[1] ,
    \slaves_02_ar_addr[0] }),
    .m02_ar_burst({\slaves_02_ar_burst[1] ,
    \slaves_02_ar_burst[0] }),
    .m02_ar_cache({\slaves_02_ar_cache[3] ,
    \slaves_02_ar_cache[2] ,
    \slaves_02_ar_cache[1] ,
    \slaves_02_ar_cache[0] }),
    .m02_ar_id({_NC117,
    _NC118,
    _NC119,
    _NC120,
    _NC121,
    _NC122,
    _NC123,
    _NC124,
    _NC125,
    _NC126,
    _NC127,
    _NC128}),
    .m02_ar_len({\slaves_02_ar_len[7] ,
    \slaves_02_ar_len[6] ,
    \slaves_02_ar_len[5] ,
    \slaves_02_ar_len[4] ,
    \slaves_02_ar_len[3] ,
    \slaves_02_ar_len[2] ,
    \slaves_02_ar_len[1] ,
    \slaves_02_ar_len[0] }),
    .m02_ar_prot({\slaves_02_ar_prot[2] ,
    \slaves_02_ar_prot[1] ,
    \slaves_02_ar_prot[0] }),
    .m02_ar_qos({\slaves_02_ar_qos[3] ,
    \slaves_02_ar_qos[2] ,
    \slaves_02_ar_qos[1] ,
    \slaves_02_ar_qos[0] }),
    .m02_ar_region({\slaves_02_ar_region[3] ,
    \slaves_02_ar_region[2] ,
    \slaves_02_ar_region[1] ,
    \slaves_02_ar_region[0] }),
    .m02_ar_size({\slaves_02_ar_size[2] ,
    \slaves_02_ar_size[1] ,
    \slaves_02_ar_size[0] }),
    .m02_ar_user({_NC129,
    _NC130}),
    .m02_aw_addr({\slaves_02_aw_addr[31] ,
    \slaves_02_aw_addr[30] ,
    \slaves_02_aw_addr[29] ,
    \slaves_02_aw_addr[28] ,
    \slaves_02_aw_addr[27] ,
    \slaves_02_aw_addr[26] ,
    \slaves_02_aw_addr[25] ,
    \slaves_02_aw_addr[24] ,
    \slaves_02_aw_addr[23] ,
    \slaves_02_aw_addr[22] ,
    \slaves_02_aw_addr[21] ,
    \slaves_02_aw_addr[20] ,
    \slaves_02_aw_addr[19] ,
    \slaves_02_aw_addr[18] ,
    \slaves_02_aw_addr[17] ,
    \slaves_02_aw_addr[16] ,
    \slaves_02_aw_addr[15] ,
    \slaves_02_aw_addr[14] ,
    \slaves_02_aw_addr[13] ,
    \slaves_02_aw_addr[12] ,
    \slaves_02_aw_addr[11] ,
    \slaves_02_aw_addr[10] ,
    \slaves_02_aw_addr[9] ,
    \slaves_02_aw_addr[8] ,
    \slaves_02_aw_addr[7] ,
    \slaves_02_aw_addr[6] ,
    \slaves_02_aw_addr[5] ,
    \slaves_02_aw_addr[4] ,
    \slaves_02_aw_addr[3] ,
    \slaves_02_aw_addr[2] ,
    \slaves_02_aw_addr[1] ,
    \slaves_02_aw_addr[0] }),
    .m02_aw_burst({\slaves_02_aw_burst[1] ,
    \slaves_02_aw_burst[0] }),
    .m02_aw_cache({\slaves_02_aw_cache[3] ,
    \slaves_02_aw_cache[2] ,
    \slaves_02_aw_cache[1] ,
    \slaves_02_aw_cache[0] }),
    .m02_aw_id({_NC131,
    _NC132,
    _NC133,
    _NC134,
    _NC135,
    _NC136,
    _NC137,
    _NC138,
    _NC139,
    _NC140,
    _NC141,
    _NC142}),
    .m02_aw_len({\slaves_02_aw_len[7] ,
    \slaves_02_aw_len[6] ,
    \slaves_02_aw_len[5] ,
    \slaves_02_aw_len[4] ,
    \slaves_02_aw_len[3] ,
    \slaves_02_aw_len[2] ,
    \slaves_02_aw_len[1] ,
    \slaves_02_aw_len[0] }),
    .m02_aw_prot({\slaves_02_aw_prot[2] ,
    \slaves_02_aw_prot[1] ,
    \slaves_02_aw_prot[0] }),
    .m02_aw_qos({\slaves_02_aw_qos[3] ,
    \slaves_02_aw_qos[2] ,
    \slaves_02_aw_qos[1] ,
    \slaves_02_aw_qos[0] }),
    .m02_aw_region({\slaves_02_aw_region[3] ,
    \slaves_02_aw_region[2] ,
    \slaves_02_aw_region[1] ,
    \slaves_02_aw_region[0] }),
    .m02_aw_size({\slaves_02_aw_size[2] ,
    \slaves_02_aw_size[1] ,
    \slaves_02_aw_size[0] }),
    .m02_aw_user({_NC143,
    _NC144}),
    .m02_b_id({_NC145,
    _NC146,
    _NC147,
    _NC148,
    _NC149,
    _NC150,
    _NC151,
    _NC152,
    _NC153,
    _NC154,
    _NC155,
    _NC156}),
    .m02_b_resp({\slaves_02_b_resp[1] ,
    \slaves_02_b_resp[0] }),
    .m02_b_user({_NC157,
    _NC158}),
    .m02_r_data({\slaves_02_r_data[31] ,
    \slaves_02_r_data[30] ,
    \slaves_02_r_data[29] ,
    \slaves_02_r_data[28] ,
    \slaves_02_r_data[27] ,
    \slaves_02_r_data[26] ,
    \slaves_02_r_data[25] ,
    \slaves_02_r_data[24] ,
    \slaves_02_r_data[23] ,
    \slaves_02_r_data[22] ,
    \slaves_02_r_data[21] ,
    \slaves_02_r_data[20] ,
    \slaves_02_r_data[19] ,
    \slaves_02_r_data[18] ,
    \slaves_02_r_data[17] ,
    \slaves_02_r_data[16] ,
    \slaves_02_r_data[15] ,
    \slaves_02_r_data[14] ,
    \slaves_02_r_data[13] ,
    \slaves_02_r_data[12] ,
    \slaves_02_r_data[11] ,
    \slaves_02_r_data[10] ,
    \slaves_02_r_data[9] ,
    \slaves_02_r_data[8] ,
    \slaves_02_r_data[7] ,
    \slaves_02_r_data[6] ,
    \slaves_02_r_data[5] ,
    \slaves_02_r_data[4] ,
    \slaves_02_r_data[3] ,
    \slaves_02_r_data[2] ,
    \slaves_02_r_data[1] ,
    \slaves_02_r_data[0] }),
    .m02_r_id({_NC159,
    _NC160,
    _NC161,
    _NC162,
    _NC163,
    _NC164,
    _NC165,
    _NC166,
    _NC167,
    _NC168,
    _NC169,
    _NC170}),
    .m02_r_resp({\slaves_02_r_resp[1] ,
    \slaves_02_r_resp[0] }),
    .m02_r_user({_NC171,
    _NC172}),
    .m02_w_data({\slaves_02_w_data[31] ,
    \slaves_02_w_data[30] ,
    \slaves_02_w_data[29] ,
    \slaves_02_w_data[28] ,
    \slaves_02_w_data[27] ,
    \slaves_02_w_data[26] ,
    \slaves_02_w_data[25] ,
    \slaves_02_w_data[24] ,
    \slaves_02_w_data[23] ,
    \slaves_02_w_data[22] ,
    \slaves_02_w_data[21] ,
    \slaves_02_w_data[20] ,
    \slaves_02_w_data[19] ,
    \slaves_02_w_data[18] ,
    \slaves_02_w_data[17] ,
    \slaves_02_w_data[16] ,
    \slaves_02_w_data[15] ,
    \slaves_02_w_data[14] ,
    \slaves_02_w_data[13] ,
    \slaves_02_w_data[12] ,
    \slaves_02_w_data[11] ,
    \slaves_02_w_data[10] ,
    \slaves_02_w_data[9] ,
    \slaves_02_w_data[8] ,
    \slaves_02_w_data[7] ,
    \slaves_02_w_data[6] ,
    \slaves_02_w_data[5] ,
    \slaves_02_w_data[4] ,
    \slaves_02_w_data[3] ,
    \slaves_02_w_data[2] ,
    \slaves_02_w_data[1] ,
    \slaves_02_w_data[0] }),
    .m02_w_strb({\slaves_02_w_strb[3] ,
    \slaves_02_w_strb[2] ,
    \slaves_02_w_strb[1] ,
    \slaves_02_w_strb[0] }),
    .m02_w_user({_NC173,
    _NC174}),
    .s00_ar_addr({\masters_00_ar_addr[31] ,
    \masters_00_ar_addr[30] ,
    \masters_00_ar_addr[29] ,
    \masters_00_ar_addr[28] ,
    \masters_00_ar_addr[27] ,
    \masters_00_ar_addr[26] ,
    \masters_00_ar_addr[25] ,
    \masters_00_ar_addr[24] ,
    \masters_00_ar_addr[23] ,
    \masters_00_ar_addr[22] ,
    \masters_00_ar_addr[21] ,
    \masters_00_ar_addr[20] ,
    \masters_00_ar_addr[19] ,
    \masters_00_ar_addr[18] ,
    \masters_00_ar_addr[17] ,
    \masters_00_ar_addr[16] ,
    \masters_00_ar_addr[15] ,
    \masters_00_ar_addr[14] ,
    \masters_00_ar_addr[13] ,
    \masters_00_ar_addr[12] ,
    \masters_00_ar_addr[11] ,
    \masters_00_ar_addr[10] ,
    \masters_00_ar_addr[9] ,
    \masters_00_ar_addr[8] ,
    \masters_00_ar_addr[7] ,
    \masters_00_ar_addr[6] ,
    \masters_00_ar_addr[5] ,
    \masters_00_ar_addr[4] ,
    \masters_00_ar_addr[3] ,
    \masters_00_ar_addr[2] ,
    \masters_00_ar_addr[1] ,
    \masters_00_ar_addr[0] }),
    .s00_ar_burst({\masters_00_ar_burst[1] ,
    \masters_00_ar_burst[0] }),
    .s00_ar_cache({\masters_00_ar_cache[3] ,
    \masters_00_ar_cache[2] ,
    \masters_00_ar_cache[1] ,
    \masters_00_ar_cache[0] }),
    .s00_ar_id({_NC175,
    _NC176,
    _NC177,
    _NC178,
    _NC179,
    _NC180,
    _NC181,
    _NC182,
    _NC183,
    _NC184}),
    .s00_ar_len({\masters_00_ar_len[7] ,
    \masters_00_ar_len[6] ,
    \masters_00_ar_len[5] ,
    \masters_00_ar_len[4] ,
    \masters_00_ar_len[3] ,
    \masters_00_ar_len[2] ,
    \masters_00_ar_len[1] ,
    \masters_00_ar_len[0] }),
    .s00_ar_prot({\masters_00_ar_prot[2] ,
    \masters_00_ar_prot[1] ,
    \masters_00_ar_prot[0] }),
    .s00_ar_qos({\masters_00_ar_qos[3] ,
    \masters_00_ar_qos[2] ,
    \masters_00_ar_qos[1] ,
    \masters_00_ar_qos[0] }),
    .s00_ar_region({\masters_00_ar_region[3] ,
    \masters_00_ar_region[2] ,
    \masters_00_ar_region[1] ,
    \masters_00_ar_region[0] }),
    .s00_ar_size({\masters_00_ar_size[2] ,
    \masters_00_ar_size[1] ,
    \masters_00_ar_size[0] }),
    .s00_ar_user({_NC185,
    _NC186}),
    .s00_aw_addr({\masters_00_aw_addr[31] ,
    \masters_00_aw_addr[30] ,
    \masters_00_aw_addr[29] ,
    \masters_00_aw_addr[28] ,
    \masters_00_aw_addr[27] ,
    \masters_00_aw_addr[26] ,
    \masters_00_aw_addr[25] ,
    \masters_00_aw_addr[24] ,
    \masters_00_aw_addr[23] ,
    \masters_00_aw_addr[22] ,
    \masters_00_aw_addr[21] ,
    \masters_00_aw_addr[20] ,
    \masters_00_aw_addr[19] ,
    \masters_00_aw_addr[18] ,
    \masters_00_aw_addr[17] ,
    \masters_00_aw_addr[16] ,
    \masters_00_aw_addr[15] ,
    \masters_00_aw_addr[14] ,
    \masters_00_aw_addr[13] ,
    \masters_00_aw_addr[12] ,
    \masters_00_aw_addr[11] ,
    \masters_00_aw_addr[10] ,
    \masters_00_aw_addr[9] ,
    \masters_00_aw_addr[8] ,
    \masters_00_aw_addr[7] ,
    \masters_00_aw_addr[6] ,
    \masters_00_aw_addr[5] ,
    \masters_00_aw_addr[4] ,
    \masters_00_aw_addr[3] ,
    \masters_00_aw_addr[2] ,
    \masters_00_aw_addr[1] ,
    \masters_00_aw_addr[0] }),
    .s00_aw_burst({\masters_00_aw_burst[1] ,
    \masters_00_aw_burst[0] }),
    .s00_aw_cache({\masters_00_aw_cache[3] ,
    \masters_00_aw_cache[2] ,
    \masters_00_aw_cache[1] ,
    \masters_00_aw_cache[0] }),
    .s00_aw_id({_NC187,
    _NC188,
    _NC189,
    _NC190,
    _NC191,
    _NC192,
    _NC193,
    _NC194,
    _NC195,
    _NC196}),
    .s00_aw_len({\masters_00_aw_len[7] ,
    \masters_00_aw_len[6] ,
    \masters_00_aw_len[5] ,
    \masters_00_aw_len[4] ,
    \masters_00_aw_len[3] ,
    \masters_00_aw_len[2] ,
    \masters_00_aw_len[1] ,
    \masters_00_aw_len[0] }),
    .s00_aw_prot({\masters_00_aw_prot[2] ,
    \masters_00_aw_prot[1] ,
    \masters_00_aw_prot[0] }),
    .s00_aw_qos({\masters_00_aw_qos[3] ,
    \masters_00_aw_qos[2] ,
    \masters_00_aw_qos[1] ,
    \masters_00_aw_qos[0] }),
    .s00_aw_region({\masters_00_aw_region[3] ,
    \masters_00_aw_region[2] ,
    \masters_00_aw_region[1] ,
    \masters_00_aw_region[0] }),
    .s00_aw_size({\masters_00_aw_size[2] ,
    \masters_00_aw_size[1] ,
    \masters_00_aw_size[0] }),
    .s00_aw_user({_NC197,
    _NC198}),
    .s00_b_id({_NC199,
    _NC200,
    _NC201,
    _NC202,
    _NC203,
    _NC204,
    _NC205,
    _NC206,
    _NC207,
    _NC208}),
    .s00_b_resp({\masters_00_b_resp[1] ,
    \masters_00_b_resp[0] }),
    .s00_b_user({_NC209,
    _NC210}),
    .s00_r_data({\masters_00_r_data[31] ,
    \masters_00_r_data[30] ,
    \masters_00_r_data[29] ,
    \masters_00_r_data[28] ,
    \masters_00_r_data[27] ,
    \masters_00_r_data[26] ,
    \masters_00_r_data[25] ,
    \masters_00_r_data[24] ,
    \masters_00_r_data[23] ,
    \masters_00_r_data[22] ,
    \masters_00_r_data[21] ,
    \masters_00_r_data[20] ,
    \masters_00_r_data[19] ,
    \masters_00_r_data[18] ,
    \masters_00_r_data[17] ,
    \masters_00_r_data[16] ,
    \masters_00_r_data[15] ,
    \masters_00_r_data[14] ,
    \masters_00_r_data[13] ,
    \masters_00_r_data[12] ,
    \masters_00_r_data[11] ,
    \masters_00_r_data[10] ,
    \masters_00_r_data[9] ,
    \masters_00_r_data[8] ,
    \masters_00_r_data[7] ,
    \masters_00_r_data[6] ,
    \masters_00_r_data[5] ,
    \masters_00_r_data[4] ,
    \masters_00_r_data[3] ,
    \masters_00_r_data[2] ,
    \masters_00_r_data[1] ,
    \masters_00_r_data[0] }),
    .s00_r_id({_NC211,
    _NC212,
    _NC213,
    _NC214,
    _NC215,
    _NC216,
    _NC217,
    _NC218,
    _NC219,
    _NC220}),
    .s00_r_resp({\masters_00_r_resp[1] ,
    \masters_00_r_resp[0] }),
    .s00_r_user({_NC221,
    _NC222}),
    .s00_w_data({\masters_00_w_data[31] ,
    \masters_00_w_data[30] ,
    \masters_00_w_data[29] ,
    \masters_00_w_data[28] ,
    \masters_00_w_data[27] ,
    \masters_00_w_data[26] ,
    \masters_00_w_data[25] ,
    \masters_00_w_data[24] ,
    \masters_00_w_data[23] ,
    \masters_00_w_data[22] ,
    \masters_00_w_data[21] ,
    \masters_00_w_data[20] ,
    \masters_00_w_data[19] ,
    \masters_00_w_data[18] ,
    \masters_00_w_data[17] ,
    \masters_00_w_data[16] ,
    \masters_00_w_data[15] ,
    \masters_00_w_data[14] ,
    \masters_00_w_data[13] ,
    \masters_00_w_data[12] ,
    \masters_00_w_data[11] ,
    \masters_00_w_data[10] ,
    \masters_00_w_data[9] ,
    \masters_00_w_data[8] ,
    \masters_00_w_data[7] ,
    \masters_00_w_data[6] ,
    \masters_00_w_data[5] ,
    \masters_00_w_data[4] ,
    \masters_00_w_data[3] ,
    \masters_00_w_data[2] ,
    \masters_00_w_data[1] ,
    \masters_00_w_data[0] }),
    .s00_w_strb({\masters_00_w_strb[3] ,
    \masters_00_w_strb[2] ,
    \masters_00_w_strb[1] ,
    \masters_00_w_strb[0] }),
    .s00_w_user({_NC223,
    _NC224}),
    .s01_ar_addr({\masters_01_ar_addr[31] ,
    \masters_01_ar_addr[30] ,
    \masters_01_ar_addr[29] ,
    \masters_01_ar_addr[28] ,
    \masters_01_ar_addr[27] ,
    \masters_01_ar_addr[26] ,
    \masters_01_ar_addr[25] ,
    \masters_01_ar_addr[24] ,
    \masters_01_ar_addr[23] ,
    \masters_01_ar_addr[22] ,
    \masters_01_ar_addr[21] ,
    \masters_01_ar_addr[20] ,
    \masters_01_ar_addr[19] ,
    \masters_01_ar_addr[18] ,
    \masters_01_ar_addr[17] ,
    \masters_01_ar_addr[16] ,
    \masters_01_ar_addr[15] ,
    \masters_01_ar_addr[14] ,
    \masters_01_ar_addr[13] ,
    \masters_01_ar_addr[12] ,
    \masters_01_ar_addr[11] ,
    \masters_01_ar_addr[10] ,
    \masters_01_ar_addr[9] ,
    \masters_01_ar_addr[8] ,
    \masters_01_ar_addr[7] ,
    \masters_01_ar_addr[6] ,
    \masters_01_ar_addr[5] ,
    \masters_01_ar_addr[4] ,
    \masters_01_ar_addr[3] ,
    \masters_01_ar_addr[2] ,
    \masters_01_ar_addr[1] ,
    \masters_01_ar_addr[0] }),
    .s01_ar_burst({\masters_01_ar_burst[1] ,
    \masters_01_ar_burst[0] }),
    .s01_ar_cache({\masters_01_ar_cache[3] ,
    \masters_01_ar_cache[2] ,
    \masters_01_ar_cache[1] ,
    \masters_01_ar_cache[0] }),
    .s01_ar_id({_NC225,
    _NC226,
    _NC227,
    _NC228,
    _NC229,
    _NC230,
    _NC231,
    _NC232,
    _NC233,
    _NC234}),
    .s01_ar_len({\masters_01_ar_len[7] ,
    \masters_01_ar_len[6] ,
    \masters_01_ar_len[5] ,
    \masters_01_ar_len[4] ,
    \masters_01_ar_len[3] ,
    \masters_01_ar_len[2] ,
    \masters_01_ar_len[1] ,
    \masters_01_ar_len[0] }),
    .s01_ar_prot({\masters_01_ar_prot[2] ,
    \masters_01_ar_prot[1] ,
    \masters_01_ar_prot[0] }),
    .s01_ar_qos({\masters_01_ar_qos[3] ,
    \masters_01_ar_qos[2] ,
    \masters_01_ar_qos[1] ,
    \masters_01_ar_qos[0] }),
    .s01_ar_region({\masters_01_ar_region[3] ,
    \masters_01_ar_region[2] ,
    \masters_01_ar_region[1] ,
    \masters_01_ar_region[0] }),
    .s01_ar_size({\masters_01_ar_size[2] ,
    \masters_01_ar_size[1] ,
    \masters_01_ar_size[0] }),
    .s01_ar_user({_NC235,
    _NC236}),
    .s01_aw_addr({\masters_01_aw_addr[31] ,
    \masters_01_aw_addr[30] ,
    \masters_01_aw_addr[29] ,
    \masters_01_aw_addr[28] ,
    \masters_01_aw_addr[27] ,
    \masters_01_aw_addr[26] ,
    \masters_01_aw_addr[25] ,
    \masters_01_aw_addr[24] ,
    \masters_01_aw_addr[23] ,
    \masters_01_aw_addr[22] ,
    \masters_01_aw_addr[21] ,
    \masters_01_aw_addr[20] ,
    \masters_01_aw_addr[19] ,
    \masters_01_aw_addr[18] ,
    \masters_01_aw_addr[17] ,
    \masters_01_aw_addr[16] ,
    \masters_01_aw_addr[15] ,
    \masters_01_aw_addr[14] ,
    \masters_01_aw_addr[13] ,
    \masters_01_aw_addr[12] ,
    \masters_01_aw_addr[11] ,
    \masters_01_aw_addr[10] ,
    \masters_01_aw_addr[9] ,
    \masters_01_aw_addr[8] ,
    \masters_01_aw_addr[7] ,
    \masters_01_aw_addr[6] ,
    \masters_01_aw_addr[5] ,
    \masters_01_aw_addr[4] ,
    \masters_01_aw_addr[3] ,
    \masters_01_aw_addr[2] ,
    \masters_01_aw_addr[1] ,
    \masters_01_aw_addr[0] }),
    .s01_aw_burst({\masters_01_aw_burst[1] ,
    \masters_01_aw_burst[0] }),
    .s01_aw_cache({\masters_01_aw_cache[3] ,
    \masters_01_aw_cache[2] ,
    \masters_01_aw_cache[1] ,
    \masters_01_aw_cache[0] }),
    .s01_aw_id({_NC237,
    _NC238,
    _NC239,
    _NC240,
    _NC241,
    _NC242,
    _NC243,
    _NC244,
    _NC245,
    _NC246}),
    .s01_aw_len({\masters_01_aw_len[7] ,
    \masters_01_aw_len[6] ,
    \masters_01_aw_len[5] ,
    \masters_01_aw_len[4] ,
    \masters_01_aw_len[3] ,
    \masters_01_aw_len[2] ,
    \masters_01_aw_len[1] ,
    \masters_01_aw_len[0] }),
    .s01_aw_prot({\masters_01_aw_prot[2] ,
    \masters_01_aw_prot[1] ,
    \masters_01_aw_prot[0] }),
    .s01_aw_qos({\masters_01_aw_qos[3] ,
    \masters_01_aw_qos[2] ,
    \masters_01_aw_qos[1] ,
    \masters_01_aw_qos[0] }),
    .s01_aw_region({\masters_01_aw_region[3] ,
    \masters_01_aw_region[2] ,
    \masters_01_aw_region[1] ,
    \masters_01_aw_region[0] }),
    .s01_aw_size({\masters_01_aw_size[2] ,
    \masters_01_aw_size[1] ,
    \masters_01_aw_size[0] }),
    .s01_aw_user({_NC247,
    _NC248}),
    .s01_b_id({_NC249,
    _NC250,
    _NC251,
    _NC252,
    _NC253,
    _NC254,
    _NC255,
    _NC256,
    _NC257,
    _NC258}),
    .s01_b_resp({\masters_01_b_resp[1] ,
    \masters_01_b_resp[0] }),
    .s01_b_user({_NC259,
    _NC260}),
    .s01_r_data({\masters_01_r_data[31] ,
    \masters_01_r_data[30] ,
    \masters_01_r_data[29] ,
    \masters_01_r_data[28] ,
    \masters_01_r_data[27] ,
    \masters_01_r_data[26] ,
    \masters_01_r_data[25] ,
    \masters_01_r_data[24] ,
    \masters_01_r_data[23] ,
    \masters_01_r_data[22] ,
    \masters_01_r_data[21] ,
    \masters_01_r_data[20] ,
    \masters_01_r_data[19] ,
    \masters_01_r_data[18] ,
    \masters_01_r_data[17] ,
    \masters_01_r_data[16] ,
    \masters_01_r_data[15] ,
    \masters_01_r_data[14] ,
    \masters_01_r_data[13] ,
    \masters_01_r_data[12] ,
    \masters_01_r_data[11] ,
    \masters_01_r_data[10] ,
    \masters_01_r_data[9] ,
    \masters_01_r_data[8] ,
    \masters_01_r_data[7] ,
    \masters_01_r_data[6] ,
    \masters_01_r_data[5] ,
    \masters_01_r_data[4] ,
    \masters_01_r_data[3] ,
    \masters_01_r_data[2] ,
    \masters_01_r_data[1] ,
    \masters_01_r_data[0] }),
    .s01_r_id({_NC261,
    _NC262,
    _NC263,
    _NC264,
    _NC265,
    _NC266,
    _NC267,
    _NC268,
    _NC269,
    _NC270}),
    .s01_r_resp({\masters_01_r_resp[1] ,
    \masters_01_r_resp[0] }),
    .s01_r_user({_NC271,
    _NC272}),
    .s01_w_data({\masters_01_w_data[31] ,
    \masters_01_w_data[30] ,
    \masters_01_w_data[29] ,
    \masters_01_w_data[28] ,
    \masters_01_w_data[27] ,
    \masters_01_w_data[26] ,
    \masters_01_w_data[25] ,
    \masters_01_w_data[24] ,
    \masters_01_w_data[23] ,
    \masters_01_w_data[22] ,
    \masters_01_w_data[21] ,
    \masters_01_w_data[20] ,
    \masters_01_w_data[19] ,
    \masters_01_w_data[18] ,
    \masters_01_w_data[17] ,
    \masters_01_w_data[16] ,
    \masters_01_w_data[15] ,
    \masters_01_w_data[14] ,
    \masters_01_w_data[13] ,
    \masters_01_w_data[12] ,
    \masters_01_w_data[11] ,
    \masters_01_w_data[10] ,
    \masters_01_w_data[9] ,
    \masters_01_w_data[8] ,
    \masters_01_w_data[7] ,
    \masters_01_w_data[6] ,
    \masters_01_w_data[5] ,
    \masters_01_w_data[4] ,
    \masters_01_w_data[3] ,
    \masters_01_w_data[2] ,
    \masters_01_w_data[1] ,
    \masters_01_w_data[0] }),
    .s01_w_strb({\masters_01_w_strb[3] ,
    \masters_01_w_strb[2] ,
    \masters_01_w_strb[1] ,
    \masters_01_w_strb[0] }),
    .s01_w_user({_NC273,
    _NC274}),
    .s02_ar_addr({\masters_02_ar_addr[31] ,
    \masters_02_ar_addr[30] ,
    \masters_02_ar_addr[29] ,
    \masters_02_ar_addr[28] ,
    \masters_02_ar_addr[27] ,
    \masters_02_ar_addr[26] ,
    \masters_02_ar_addr[25] ,
    \masters_02_ar_addr[24] ,
    \masters_02_ar_addr[23] ,
    \masters_02_ar_addr[22] ,
    \masters_02_ar_addr[21] ,
    \masters_02_ar_addr[20] ,
    \masters_02_ar_addr[19] ,
    \masters_02_ar_addr[18] ,
    \masters_02_ar_addr[17] ,
    \masters_02_ar_addr[16] ,
    \masters_02_ar_addr[15] ,
    \masters_02_ar_addr[14] ,
    \masters_02_ar_addr[13] ,
    \masters_02_ar_addr[12] ,
    \masters_02_ar_addr[11] ,
    \masters_02_ar_addr[10] ,
    \masters_02_ar_addr[9] ,
    \masters_02_ar_addr[8] ,
    \masters_02_ar_addr[7] ,
    \masters_02_ar_addr[6] ,
    \masters_02_ar_addr[5] ,
    \masters_02_ar_addr[4] ,
    \masters_02_ar_addr[3] ,
    \masters_02_ar_addr[2] ,
    \masters_02_ar_addr[1] ,
    \masters_02_ar_addr[0] }),
    .s02_ar_burst({\masters_02_ar_burst[1] ,
    \masters_02_ar_burst[0] }),
    .s02_ar_cache({\masters_02_ar_cache[3] ,
    \masters_02_ar_cache[2] ,
    \masters_02_ar_cache[1] ,
    \masters_02_ar_cache[0] }),
    .s02_ar_id({_NC275,
    _NC276,
    _NC277,
    _NC278,
    _NC279,
    _NC280,
    _NC281,
    _NC282,
    _NC283,
    _NC284}),
    .s02_ar_len({\masters_02_ar_len[7] ,
    \masters_02_ar_len[6] ,
    \masters_02_ar_len[5] ,
    \masters_02_ar_len[4] ,
    \masters_02_ar_len[3] ,
    \masters_02_ar_len[2] ,
    \masters_02_ar_len[1] ,
    \masters_02_ar_len[0] }),
    .s02_ar_prot({\masters_02_ar_prot[2] ,
    \masters_02_ar_prot[1] ,
    \masters_02_ar_prot[0] }),
    .s02_ar_qos({\masters_02_ar_qos[3] ,
    \masters_02_ar_qos[2] ,
    \masters_02_ar_qos[1] ,
    \masters_02_ar_qos[0] }),
    .s02_ar_region({\masters_02_ar_region[3] ,
    \masters_02_ar_region[2] ,
    \masters_02_ar_region[1] ,
    \masters_02_ar_region[0] }),
    .s02_ar_size({\masters_02_ar_size[2] ,
    \masters_02_ar_size[1] ,
    \masters_02_ar_size[0] }),
    .s02_ar_user({_NC285,
    _NC286}),
    .s02_aw_addr({\masters_02_aw_addr[31] ,
    \masters_02_aw_addr[30] ,
    \masters_02_aw_addr[29] ,
    \masters_02_aw_addr[28] ,
    \masters_02_aw_addr[27] ,
    \masters_02_aw_addr[26] ,
    \masters_02_aw_addr[25] ,
    \masters_02_aw_addr[24] ,
    \masters_02_aw_addr[23] ,
    \masters_02_aw_addr[22] ,
    \masters_02_aw_addr[21] ,
    \masters_02_aw_addr[20] ,
    \masters_02_aw_addr[19] ,
    \masters_02_aw_addr[18] ,
    \masters_02_aw_addr[17] ,
    \masters_02_aw_addr[16] ,
    \masters_02_aw_addr[15] ,
    \masters_02_aw_addr[14] ,
    \masters_02_aw_addr[13] ,
    \masters_02_aw_addr[12] ,
    \masters_02_aw_addr[11] ,
    \masters_02_aw_addr[10] ,
    \masters_02_aw_addr[9] ,
    \masters_02_aw_addr[8] ,
    \masters_02_aw_addr[7] ,
    \masters_02_aw_addr[6] ,
    \masters_02_aw_addr[5] ,
    \masters_02_aw_addr[4] ,
    \masters_02_aw_addr[3] ,
    \masters_02_aw_addr[2] ,
    \masters_02_aw_addr[1] ,
    \masters_02_aw_addr[0] }),
    .s02_aw_burst({\masters_02_aw_burst[1] ,
    \masters_02_aw_burst[0] }),
    .s02_aw_cache({\masters_02_aw_cache[3] ,
    \masters_02_aw_cache[2] ,
    \masters_02_aw_cache[1] ,
    \masters_02_aw_cache[0] }),
    .s02_aw_id({_NC287,
    _NC288,
    _NC289,
    _NC290,
    _NC291,
    _NC292,
    _NC293,
    _NC294,
    _NC295,
    _NC296}),
    .s02_aw_len({\masters_02_aw_len[7] ,
    \masters_02_aw_len[6] ,
    \masters_02_aw_len[5] ,
    \masters_02_aw_len[4] ,
    \masters_02_aw_len[3] ,
    \masters_02_aw_len[2] ,
    \masters_02_aw_len[1] ,
    \masters_02_aw_len[0] }),
    .s02_aw_prot({\masters_02_aw_prot[2] ,
    \masters_02_aw_prot[1] ,
    \masters_02_aw_prot[0] }),
    .s02_aw_qos({\masters_02_aw_qos[3] ,
    \masters_02_aw_qos[2] ,
    \masters_02_aw_qos[1] ,
    \masters_02_aw_qos[0] }),
    .s02_aw_region({\masters_02_aw_region[3] ,
    \masters_02_aw_region[2] ,
    \masters_02_aw_region[1] ,
    \masters_02_aw_region[0] }),
    .s02_aw_size({\masters_02_aw_size[2] ,
    \masters_02_aw_size[1] ,
    \masters_02_aw_size[0] }),
    .s02_aw_user({_NC297,
    _NC298}),
    .s02_b_id({_NC299,
    _NC300,
    _NC301,
    _NC302,
    _NC303,
    _NC304,
    _NC305,
    _NC306,
    _NC307,
    _NC308}),
    .s02_b_resp({\masters_02_b_resp[1] ,
    \masters_02_b_resp[0] }),
    .s02_b_user({_NC309,
    _NC310}),
    .s02_r_data({\masters_02_r_data[31] ,
    \masters_02_r_data[30] ,
    \masters_02_r_data[29] ,
    \masters_02_r_data[28] ,
    \masters_02_r_data[27] ,
    \masters_02_r_data[26] ,
    \masters_02_r_data[25] ,
    \masters_02_r_data[24] ,
    \masters_02_r_data[23] ,
    \masters_02_r_data[22] ,
    \masters_02_r_data[21] ,
    \masters_02_r_data[20] ,
    \masters_02_r_data[19] ,
    \masters_02_r_data[18] ,
    \masters_02_r_data[17] ,
    \masters_02_r_data[16] ,
    \masters_02_r_data[15] ,
    \masters_02_r_data[14] ,
    \masters_02_r_data[13] ,
    \masters_02_r_data[12] ,
    \masters_02_r_data[11] ,
    \masters_02_r_data[10] ,
    \masters_02_r_data[9] ,
    \masters_02_r_data[8] ,
    \masters_02_r_data[7] ,
    \masters_02_r_data[6] ,
    \masters_02_r_data[5] ,
    \masters_02_r_data[4] ,
    \masters_02_r_data[3] ,
    \masters_02_r_data[2] ,
    \masters_02_r_data[1] ,
    \masters_02_r_data[0] }),
    .s02_r_id({_NC311,
    _NC312,
    _NC313,
    _NC314,
    _NC315,
    _NC316,
    _NC317,
    _NC318,
    _NC319,
    _NC320}),
    .s02_r_resp({\masters_02_r_resp[1] ,
    \masters_02_r_resp[0] }),
    .s02_r_user({_NC321,
    _NC322}),
    .s02_w_data({\masters_02_w_data[31] ,
    \masters_02_w_data[30] ,
    \masters_02_w_data[29] ,
    \masters_02_w_data[28] ,
    \masters_02_w_data[27] ,
    \masters_02_w_data[26] ,
    \masters_02_w_data[25] ,
    \masters_02_w_data[24] ,
    \masters_02_w_data[23] ,
    \masters_02_w_data[22] ,
    \masters_02_w_data[21] ,
    \masters_02_w_data[20] ,
    \masters_02_w_data[19] ,
    \masters_02_w_data[18] ,
    \masters_02_w_data[17] ,
    \masters_02_w_data[16] ,
    \masters_02_w_data[15] ,
    \masters_02_w_data[14] ,
    \masters_02_w_data[13] ,
    \masters_02_w_data[12] ,
    \masters_02_w_data[11] ,
    \masters_02_w_data[10] ,
    \masters_02_w_data[9] ,
    \masters_02_w_data[8] ,
    \masters_02_w_data[7] ,
    \masters_02_w_data[6] ,
    \masters_02_w_data[5] ,
    \masters_02_w_data[4] ,
    \masters_02_w_data[3] ,
    \masters_02_w_data[2] ,
    \masters_02_w_data[1] ,
    \masters_02_w_data[0] }),
    .s02_w_strb({\masters_02_w_strb[3] ,
    \masters_02_w_strb[2] ,
    \masters_02_w_strb[1] ,
    \masters_02_w_strb[0] }),
    .s02_w_user({_NC323,
    _NC324}));
 mba_core_region core_region_i (.clk(clk_int),
    .clock_gating_i(clk_gate_core_int),
    .core_busy_o(core_busy_int),
    .core_master_ar_lock(masters_00_ar_lock),
    .core_master_ar_ready(masters_00_ar_ready),
    .core_master_ar_valid(masters_00_ar_valid),
    .core_master_aw_lock(masters_00_aw_lock),
    .core_master_aw_ready(masters_00_aw_ready),
    .core_master_aw_valid(masters_00_aw_valid),
    .core_master_b_ready(masters_00_b_ready),
    .core_master_b_valid(masters_00_b_valid),
    .core_master_r_last(masters_00_r_last),
    .core_master_r_ready(masters_00_r_ready),
    .core_master_r_valid(masters_00_r_valid),
    .core_master_w_last(masters_00_w_last),
    .core_master_w_ready(masters_00_w_ready),
    .core_master_w_valid(masters_00_w_valid),
    .data_slave_ar_lock(slaves_01_ar_lock),
    .data_slave_ar_ready(slaves_01_ar_ready),
    .data_slave_ar_valid(slaves_01_ar_valid),
    .data_slave_aw_lock(slaves_01_aw_lock),
    .data_slave_aw_ready(slaves_01_aw_ready),
    .data_slave_aw_valid(slaves_01_aw_valid),
    .data_slave_b_ready(slaves_01_b_ready),
    .data_slave_b_valid(slaves_01_b_valid),
    .data_slave_r_last(slaves_01_r_last),
    .data_slave_r_ready(slaves_01_r_ready),
    .data_slave_r_valid(slaves_01_r_valid),
    .data_slave_w_last(slaves_01_w_last),
    .data_slave_w_ready(slaves_01_w_ready),
    .data_slave_w_valid(slaves_01_w_valid),
    .dbg_master_ar_lock(masters_01_ar_lock),
    .dbg_master_ar_ready(masters_01_ar_ready),
    .dbg_master_ar_valid(masters_01_ar_valid),
    .dbg_master_aw_lock(masters_01_aw_lock),
    .dbg_master_aw_ready(masters_01_aw_ready),
    .dbg_master_aw_valid(masters_01_aw_valid),
    .dbg_master_b_ready(masters_01_b_ready),
    .dbg_master_b_valid(masters_01_b_valid),
    .dbg_master_r_last(masters_01_r_last),
    .dbg_master_r_ready(masters_01_r_ready),
    .dbg_master_r_valid(masters_01_r_valid),
    .dbg_master_w_last(masters_01_w_last),
    .dbg_master_w_ready(masters_01_w_ready),
    .dbg_master_w_valid(masters_01_w_valid),
    .debug_gnt(debug_gnt),
    .debug_req(debug_req),
    .debug_rvalid(debug_rvalid),
    .debug_we(debug_we),
    .fetch_enable_i(fetch_enable_int),
    .instr_slave_ar_lock(slaves_00_ar_lock),
    .instr_slave_ar_ready(slaves_00_ar_ready),
    .instr_slave_ar_valid(slaves_00_ar_valid),
    .instr_slave_aw_lock(slaves_00_aw_lock),
    .instr_slave_aw_ready(slaves_00_aw_ready),
    .instr_slave_aw_valid(slaves_00_aw_valid),
    .instr_slave_b_ready(slaves_00_b_ready),
    .instr_slave_b_valid(slaves_00_b_valid),
    .instr_slave_r_last(slaves_00_r_last),
    .instr_slave_r_ready(slaves_00_r_ready),
    .instr_slave_r_valid(slaves_00_r_valid),
    .instr_slave_w_last(slaves_00_w_last),
    .instr_slave_w_ready(slaves_00_w_ready),
    .instr_slave_w_valid(slaves_00_w_valid),
    .mba_data_mem_csb0_o(mba_data_mem_csb0_o),
    .mba_data_mem_csb1_o(mba_data_mem_csb1_o),
    .mba_data_mem_web0_o(mba_data_mem_web0_o),
    .mba_instr_mem_csb0_o(mba_instr_mem_csb0_o),
    .mba_instr_mem_csb1_o(mba_instr_mem_csb1_o),
    .mba_instr_mem_web0_o(mba_instr_mem_web0_o),
    .rst_n(rstn_int),
    .tck_i(io_in[12]),
    .tdi_i(io_in[15]),
    .tdo_o(io_out[26]),
    .testmode_i(la_data_in[2]),
    .tms_i(io_in[14]),
    .trstn_i(io_in[13]),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .boot_addr_i({\boot_addr_int[31] ,
    \boot_addr_int[30] ,
    \boot_addr_int[29] ,
    \boot_addr_int[28] ,
    \boot_addr_int[27] ,
    \boot_addr_int[26] ,
    \boot_addr_int[25] ,
    \boot_addr_int[24] ,
    \boot_addr_int[23] ,
    \boot_addr_int[22] ,
    \boot_addr_int[21] ,
    \boot_addr_int[20] ,
    \boot_addr_int[19] ,
    \boot_addr_int[18] ,
    \boot_addr_int[17] ,
    \boot_addr_int[16] ,
    \boot_addr_int[15] ,
    \boot_addr_int[14] ,
    \boot_addr_int[13] ,
    \boot_addr_int[12] ,
    \boot_addr_int[11] ,
    \boot_addr_int[10] ,
    \boot_addr_int[9] ,
    \boot_addr_int[8] ,
    \boot_addr_int[7] ,
    \boot_addr_int[6] ,
    \boot_addr_int[5] ,
    \boot_addr_int[4] ,
    \boot_addr_int[3] ,
    \boot_addr_int[2] ,
    \boot_addr_int[1] ,
    \boot_addr_int[0] }),
    .core_master_ar_addr({\masters_00_ar_addr[31] ,
    \masters_00_ar_addr[30] ,
    \masters_00_ar_addr[29] ,
    \masters_00_ar_addr[28] ,
    \masters_00_ar_addr[27] ,
    \masters_00_ar_addr[26] ,
    \masters_00_ar_addr[25] ,
    \masters_00_ar_addr[24] ,
    \masters_00_ar_addr[23] ,
    \masters_00_ar_addr[22] ,
    \masters_00_ar_addr[21] ,
    \masters_00_ar_addr[20] ,
    \masters_00_ar_addr[19] ,
    \masters_00_ar_addr[18] ,
    \masters_00_ar_addr[17] ,
    \masters_00_ar_addr[16] ,
    \masters_00_ar_addr[15] ,
    \masters_00_ar_addr[14] ,
    \masters_00_ar_addr[13] ,
    \masters_00_ar_addr[12] ,
    \masters_00_ar_addr[11] ,
    \masters_00_ar_addr[10] ,
    \masters_00_ar_addr[9] ,
    \masters_00_ar_addr[8] ,
    \masters_00_ar_addr[7] ,
    \masters_00_ar_addr[6] ,
    \masters_00_ar_addr[5] ,
    \masters_00_ar_addr[4] ,
    \masters_00_ar_addr[3] ,
    \masters_00_ar_addr[2] ,
    \masters_00_ar_addr[1] ,
    \masters_00_ar_addr[0] }),
    .core_master_ar_burst({\masters_00_ar_burst[1] ,
    \masters_00_ar_burst[0] }),
    .core_master_ar_cache({\masters_00_ar_cache[3] ,
    \masters_00_ar_cache[2] ,
    \masters_00_ar_cache[1] ,
    \masters_00_ar_cache[0] }),
    .core_master_ar_id({_NC325,
    _NC326,
    _NC327,
    _NC328,
    _NC329,
    _NC330,
    _NC331,
    _NC332,
    _NC333,
    _NC334}),
    .core_master_ar_len({\masters_00_ar_len[7] ,
    \masters_00_ar_len[6] ,
    \masters_00_ar_len[5] ,
    \masters_00_ar_len[4] ,
    \masters_00_ar_len[3] ,
    \masters_00_ar_len[2] ,
    \masters_00_ar_len[1] ,
    \masters_00_ar_len[0] }),
    .core_master_ar_prot({\masters_00_ar_prot[2] ,
    \masters_00_ar_prot[1] ,
    \masters_00_ar_prot[0] }),
    .core_master_ar_qos({\masters_00_ar_qos[3] ,
    \masters_00_ar_qos[2] ,
    \masters_00_ar_qos[1] ,
    \masters_00_ar_qos[0] }),
    .core_master_ar_region({\masters_00_ar_region[3] ,
    \masters_00_ar_region[2] ,
    \masters_00_ar_region[1] ,
    \masters_00_ar_region[0] }),
    .core_master_ar_size({\masters_00_ar_size[2] ,
    \masters_00_ar_size[1] ,
    \masters_00_ar_size[0] }),
    .core_master_ar_user({_NC335,
    _NC336}),
    .core_master_aw_addr({\masters_00_aw_addr[31] ,
    \masters_00_aw_addr[30] ,
    \masters_00_aw_addr[29] ,
    \masters_00_aw_addr[28] ,
    \masters_00_aw_addr[27] ,
    \masters_00_aw_addr[26] ,
    \masters_00_aw_addr[25] ,
    \masters_00_aw_addr[24] ,
    \masters_00_aw_addr[23] ,
    \masters_00_aw_addr[22] ,
    \masters_00_aw_addr[21] ,
    \masters_00_aw_addr[20] ,
    \masters_00_aw_addr[19] ,
    \masters_00_aw_addr[18] ,
    \masters_00_aw_addr[17] ,
    \masters_00_aw_addr[16] ,
    \masters_00_aw_addr[15] ,
    \masters_00_aw_addr[14] ,
    \masters_00_aw_addr[13] ,
    \masters_00_aw_addr[12] ,
    \masters_00_aw_addr[11] ,
    \masters_00_aw_addr[10] ,
    \masters_00_aw_addr[9] ,
    \masters_00_aw_addr[8] ,
    \masters_00_aw_addr[7] ,
    \masters_00_aw_addr[6] ,
    \masters_00_aw_addr[5] ,
    \masters_00_aw_addr[4] ,
    \masters_00_aw_addr[3] ,
    \masters_00_aw_addr[2] ,
    \masters_00_aw_addr[1] ,
    \masters_00_aw_addr[0] }),
    .core_master_aw_burst({\masters_00_aw_burst[1] ,
    \masters_00_aw_burst[0] }),
    .core_master_aw_cache({\masters_00_aw_cache[3] ,
    \masters_00_aw_cache[2] ,
    \masters_00_aw_cache[1] ,
    \masters_00_aw_cache[0] }),
    .core_master_aw_id({_NC337,
    _NC338,
    _NC339,
    _NC340,
    _NC341,
    _NC342,
    _NC343,
    _NC344,
    _NC345,
    _NC346}),
    .core_master_aw_len({\masters_00_aw_len[7] ,
    \masters_00_aw_len[6] ,
    \masters_00_aw_len[5] ,
    \masters_00_aw_len[4] ,
    \masters_00_aw_len[3] ,
    \masters_00_aw_len[2] ,
    \masters_00_aw_len[1] ,
    \masters_00_aw_len[0] }),
    .core_master_aw_prot({\masters_00_aw_prot[2] ,
    \masters_00_aw_prot[1] ,
    \masters_00_aw_prot[0] }),
    .core_master_aw_qos({\masters_00_aw_qos[3] ,
    \masters_00_aw_qos[2] ,
    \masters_00_aw_qos[1] ,
    \masters_00_aw_qos[0] }),
    .core_master_aw_region({\masters_00_aw_region[3] ,
    \masters_00_aw_region[2] ,
    \masters_00_aw_region[1] ,
    \masters_00_aw_region[0] }),
    .core_master_aw_size({\masters_00_aw_size[2] ,
    \masters_00_aw_size[1] ,
    \masters_00_aw_size[0] }),
    .core_master_aw_user({_NC347,
    _NC348}),
    .core_master_b_id({_NC349,
    _NC350,
    _NC351,
    _NC352,
    _NC353,
    _NC354,
    _NC355,
    _NC356,
    _NC357,
    _NC358}),
    .core_master_b_resp({\masters_00_b_resp[1] ,
    \masters_00_b_resp[0] }),
    .core_master_b_user({_NC359,
    _NC360}),
    .core_master_r_data({_NC361,
    _NC362,
    _NC363,
    _NC364,
    _NC365,
    _NC366,
    _NC367,
    _NC368,
    _NC369,
    _NC370,
    _NC371,
    _NC372,
    _NC373,
    _NC374,
    _NC375,
    _NC376,
    _NC377,
    _NC378,
    _NC379,
    _NC380,
    _NC381,
    _NC382,
    _NC383,
    _NC384,
    _NC385,
    _NC386,
    _NC387,
    _NC388,
    _NC389,
    _NC390,
    _NC391,
    _NC392,
    _NC393,
    _NC394,
    _NC395,
    _NC396,
    _NC397,
    _NC398,
    _NC399,
    _NC400,
    _NC401,
    _NC402,
    _NC403,
    _NC404,
    _NC405,
    _NC406,
    _NC407,
    _NC408,
    _NC409,
    _NC410,
    _NC411,
    _NC412,
    _NC413,
    _NC414,
    _NC415,
    _NC416,
    _NC417,
    _NC418,
    _NC419,
    _NC420,
    _NC421,
    _NC422,
    _NC423,
    _NC424}),
    .core_master_r_id({_NC425,
    _NC426,
    _NC427,
    _NC428,
    _NC429,
    _NC430,
    _NC431,
    _NC432,
    _NC433,
    _NC434}),
    .core_master_r_resp({\masters_00_r_resp[1] ,
    \masters_00_r_resp[0] }),
    .core_master_r_user({_NC435,
    _NC436}),
    .core_master_w_data({_NC437,
    _NC438,
    _NC439,
    _NC440,
    _NC441,
    _NC442,
    _NC443,
    _NC444,
    _NC445,
    _NC446,
    _NC447,
    _NC448,
    _NC449,
    _NC450,
    _NC451,
    _NC452,
    _NC453,
    _NC454,
    _NC455,
    _NC456,
    _NC457,
    _NC458,
    _NC459,
    _NC460,
    _NC461,
    _NC462,
    _NC463,
    _NC464,
    _NC465,
    _NC466,
    _NC467,
    _NC468,
    _NC469,
    _NC470,
    _NC471,
    _NC472,
    _NC473,
    _NC474,
    _NC475,
    _NC476,
    _NC477,
    _NC478,
    _NC479,
    _NC480,
    _NC481,
    _NC482,
    _NC483,
    _NC484,
    _NC485,
    _NC486,
    _NC487,
    _NC488,
    _NC489,
    _NC490,
    _NC491,
    _NC492,
    _NC493,
    _NC494,
    _NC495,
    _NC496,
    _NC497,
    _NC498,
    _NC499,
    _NC500}),
    .core_master_w_strb({_NC501,
    _NC502,
    _NC503,
    _NC504,
    _NC505,
    _NC506,
    _NC507,
    _NC508}),
    .core_master_w_user({_NC509,
    _NC510}),
    .data_slave_ar_addr({\slaves_01_ar_addr[31] ,
    \slaves_01_ar_addr[30] ,
    \slaves_01_ar_addr[29] ,
    \slaves_01_ar_addr[28] ,
    \slaves_01_ar_addr[27] ,
    \slaves_01_ar_addr[26] ,
    \slaves_01_ar_addr[25] ,
    \slaves_01_ar_addr[24] ,
    \slaves_01_ar_addr[23] ,
    \slaves_01_ar_addr[22] ,
    \slaves_01_ar_addr[21] ,
    \slaves_01_ar_addr[20] ,
    \slaves_01_ar_addr[19] ,
    \slaves_01_ar_addr[18] ,
    \slaves_01_ar_addr[17] ,
    \slaves_01_ar_addr[16] ,
    \slaves_01_ar_addr[15] ,
    \slaves_01_ar_addr[14] ,
    \slaves_01_ar_addr[13] ,
    \slaves_01_ar_addr[12] ,
    \slaves_01_ar_addr[11] ,
    \slaves_01_ar_addr[10] ,
    \slaves_01_ar_addr[9] ,
    \slaves_01_ar_addr[8] ,
    \slaves_01_ar_addr[7] ,
    \slaves_01_ar_addr[6] ,
    \slaves_01_ar_addr[5] ,
    \slaves_01_ar_addr[4] ,
    \slaves_01_ar_addr[3] ,
    \slaves_01_ar_addr[2] ,
    \slaves_01_ar_addr[1] ,
    \slaves_01_ar_addr[0] }),
    .data_slave_ar_burst({\slaves_01_ar_burst[1] ,
    \slaves_01_ar_burst[0] }),
    .data_slave_ar_cache({\slaves_01_ar_cache[3] ,
    \slaves_01_ar_cache[2] ,
    \slaves_01_ar_cache[1] ,
    \slaves_01_ar_cache[0] }),
    .data_slave_ar_id({_NC511,
    _NC512,
    _NC513,
    _NC514,
    _NC515,
    _NC516,
    _NC517,
    _NC518,
    _NC519,
    _NC520}),
    .data_slave_ar_len({\slaves_01_ar_len[7] ,
    \slaves_01_ar_len[6] ,
    \slaves_01_ar_len[5] ,
    \slaves_01_ar_len[4] ,
    \slaves_01_ar_len[3] ,
    \slaves_01_ar_len[2] ,
    \slaves_01_ar_len[1] ,
    \slaves_01_ar_len[0] }),
    .data_slave_ar_prot({\slaves_01_ar_prot[2] ,
    \slaves_01_ar_prot[1] ,
    \slaves_01_ar_prot[0] }),
    .data_slave_ar_qos({\slaves_01_ar_qos[3] ,
    \slaves_01_ar_qos[2] ,
    \slaves_01_ar_qos[1] ,
    \slaves_01_ar_qos[0] }),
    .data_slave_ar_region({\slaves_01_ar_region[3] ,
    \slaves_01_ar_region[2] ,
    \slaves_01_ar_region[1] ,
    \slaves_01_ar_region[0] }),
    .data_slave_ar_size({\slaves_01_ar_size[2] ,
    \slaves_01_ar_size[1] ,
    \slaves_01_ar_size[0] }),
    .data_slave_ar_user({_NC521,
    _NC522}),
    .data_slave_aw_addr({\slaves_01_aw_addr[31] ,
    \slaves_01_aw_addr[30] ,
    \slaves_01_aw_addr[29] ,
    \slaves_01_aw_addr[28] ,
    \slaves_01_aw_addr[27] ,
    \slaves_01_aw_addr[26] ,
    \slaves_01_aw_addr[25] ,
    \slaves_01_aw_addr[24] ,
    \slaves_01_aw_addr[23] ,
    \slaves_01_aw_addr[22] ,
    \slaves_01_aw_addr[21] ,
    \slaves_01_aw_addr[20] ,
    \slaves_01_aw_addr[19] ,
    \slaves_01_aw_addr[18] ,
    \slaves_01_aw_addr[17] ,
    \slaves_01_aw_addr[16] ,
    \slaves_01_aw_addr[15] ,
    \slaves_01_aw_addr[14] ,
    \slaves_01_aw_addr[13] ,
    \slaves_01_aw_addr[12] ,
    \slaves_01_aw_addr[11] ,
    \slaves_01_aw_addr[10] ,
    \slaves_01_aw_addr[9] ,
    \slaves_01_aw_addr[8] ,
    \slaves_01_aw_addr[7] ,
    \slaves_01_aw_addr[6] ,
    \slaves_01_aw_addr[5] ,
    \slaves_01_aw_addr[4] ,
    \slaves_01_aw_addr[3] ,
    \slaves_01_aw_addr[2] ,
    \slaves_01_aw_addr[1] ,
    \slaves_01_aw_addr[0] }),
    .data_slave_aw_burst({\slaves_01_aw_burst[1] ,
    \slaves_01_aw_burst[0] }),
    .data_slave_aw_cache({\slaves_01_aw_cache[3] ,
    \slaves_01_aw_cache[2] ,
    \slaves_01_aw_cache[1] ,
    \slaves_01_aw_cache[0] }),
    .data_slave_aw_id({_NC523,
    _NC524,
    _NC525,
    _NC526,
    _NC527,
    _NC528,
    _NC529,
    _NC530,
    _NC531,
    _NC532}),
    .data_slave_aw_len({\slaves_01_aw_len[7] ,
    \slaves_01_aw_len[6] ,
    \slaves_01_aw_len[5] ,
    \slaves_01_aw_len[4] ,
    \slaves_01_aw_len[3] ,
    \slaves_01_aw_len[2] ,
    \slaves_01_aw_len[1] ,
    \slaves_01_aw_len[0] }),
    .data_slave_aw_prot({\slaves_01_aw_prot[2] ,
    \slaves_01_aw_prot[1] ,
    \slaves_01_aw_prot[0] }),
    .data_slave_aw_qos({\slaves_01_aw_qos[3] ,
    \slaves_01_aw_qos[2] ,
    \slaves_01_aw_qos[1] ,
    \slaves_01_aw_qos[0] }),
    .data_slave_aw_region({\slaves_01_aw_region[3] ,
    \slaves_01_aw_region[2] ,
    \slaves_01_aw_region[1] ,
    \slaves_01_aw_region[0] }),
    .data_slave_aw_size({\slaves_01_aw_size[2] ,
    \slaves_01_aw_size[1] ,
    \slaves_01_aw_size[0] }),
    .data_slave_aw_user({_NC533,
    _NC534}),
    .data_slave_b_id({_NC535,
    _NC536,
    _NC537,
    _NC538,
    _NC539,
    _NC540,
    _NC541,
    _NC542,
    _NC543,
    _NC544}),
    .data_slave_b_resp({\slaves_01_b_resp[1] ,
    \slaves_01_b_resp[0] }),
    .data_slave_b_user({_NC545,
    _NC546}),
    .data_slave_r_data({_NC547,
    _NC548,
    _NC549,
    _NC550,
    _NC551,
    _NC552,
    _NC553,
    _NC554,
    _NC555,
    _NC556,
    _NC557,
    _NC558,
    _NC559,
    _NC560,
    _NC561,
    _NC562,
    _NC563,
    _NC564,
    _NC565,
    _NC566,
    _NC567,
    _NC568,
    _NC569,
    _NC570,
    _NC571,
    _NC572,
    _NC573,
    _NC574,
    _NC575,
    _NC576,
    _NC577,
    _NC578,
    _NC579,
    _NC580,
    _NC581,
    _NC582,
    _NC583,
    _NC584,
    _NC585,
    _NC586,
    _NC587,
    _NC588,
    _NC589,
    _NC590,
    _NC591,
    _NC592,
    _NC593,
    _NC594,
    _NC595,
    _NC596,
    _NC597,
    _NC598,
    _NC599,
    _NC600,
    _NC601,
    _NC602,
    _NC603,
    _NC604,
    _NC605,
    _NC606,
    _NC607,
    _NC608,
    _NC609,
    _NC610}),
    .data_slave_r_id({_NC611,
    _NC612,
    _NC613,
    _NC614,
    _NC615,
    _NC616,
    _NC617,
    _NC618,
    _NC619,
    _NC620}),
    .data_slave_r_resp({\slaves_01_r_resp[1] ,
    \slaves_01_r_resp[0] }),
    .data_slave_r_user({_NC621,
    _NC622}),
    .data_slave_w_data({_NC623,
    _NC624,
    _NC625,
    _NC626,
    _NC627,
    _NC628,
    _NC629,
    _NC630,
    _NC631,
    _NC632,
    _NC633,
    _NC634,
    _NC635,
    _NC636,
    _NC637,
    _NC638,
    _NC639,
    _NC640,
    _NC641,
    _NC642,
    _NC643,
    _NC644,
    _NC645,
    _NC646,
    _NC647,
    _NC648,
    _NC649,
    _NC650,
    _NC651,
    _NC652,
    _NC653,
    _NC654,
    _NC655,
    _NC656,
    _NC657,
    _NC658,
    _NC659,
    _NC660,
    _NC661,
    _NC662,
    _NC663,
    _NC664,
    _NC665,
    _NC666,
    _NC667,
    _NC668,
    _NC669,
    _NC670,
    _NC671,
    _NC672,
    _NC673,
    _NC674,
    _NC675,
    _NC676,
    _NC677,
    _NC678,
    _NC679,
    _NC680,
    _NC681,
    _NC682,
    _NC683,
    _NC684,
    _NC685,
    _NC686}),
    .data_slave_w_strb({_NC687,
    _NC688,
    _NC689,
    _NC690,
    _NC691,
    _NC692,
    _NC693,
    _NC694}),
    .data_slave_w_user({_NC695,
    _NC696}),
    .dbg_master_ar_addr({\masters_01_ar_addr[31] ,
    \masters_01_ar_addr[30] ,
    \masters_01_ar_addr[29] ,
    \masters_01_ar_addr[28] ,
    \masters_01_ar_addr[27] ,
    \masters_01_ar_addr[26] ,
    \masters_01_ar_addr[25] ,
    \masters_01_ar_addr[24] ,
    \masters_01_ar_addr[23] ,
    \masters_01_ar_addr[22] ,
    \masters_01_ar_addr[21] ,
    \masters_01_ar_addr[20] ,
    \masters_01_ar_addr[19] ,
    \masters_01_ar_addr[18] ,
    \masters_01_ar_addr[17] ,
    \masters_01_ar_addr[16] ,
    \masters_01_ar_addr[15] ,
    \masters_01_ar_addr[14] ,
    \masters_01_ar_addr[13] ,
    \masters_01_ar_addr[12] ,
    \masters_01_ar_addr[11] ,
    \masters_01_ar_addr[10] ,
    \masters_01_ar_addr[9] ,
    \masters_01_ar_addr[8] ,
    \masters_01_ar_addr[7] ,
    \masters_01_ar_addr[6] ,
    \masters_01_ar_addr[5] ,
    \masters_01_ar_addr[4] ,
    \masters_01_ar_addr[3] ,
    \masters_01_ar_addr[2] ,
    \masters_01_ar_addr[1] ,
    \masters_01_ar_addr[0] }),
    .dbg_master_ar_burst({\masters_01_ar_burst[1] ,
    \masters_01_ar_burst[0] }),
    .dbg_master_ar_cache({\masters_01_ar_cache[3] ,
    \masters_01_ar_cache[2] ,
    \masters_01_ar_cache[1] ,
    \masters_01_ar_cache[0] }),
    .dbg_master_ar_id({_NC697,
    _NC698,
    _NC699,
    _NC700,
    _NC701,
    _NC702,
    _NC703,
    _NC704,
    _NC705,
    _NC706}),
    .dbg_master_ar_len({\masters_01_ar_len[7] ,
    \masters_01_ar_len[6] ,
    \masters_01_ar_len[5] ,
    \masters_01_ar_len[4] ,
    \masters_01_ar_len[3] ,
    \masters_01_ar_len[2] ,
    \masters_01_ar_len[1] ,
    \masters_01_ar_len[0] }),
    .dbg_master_ar_prot({\masters_01_ar_prot[2] ,
    \masters_01_ar_prot[1] ,
    \masters_01_ar_prot[0] }),
    .dbg_master_ar_qos({\masters_01_ar_qos[3] ,
    \masters_01_ar_qos[2] ,
    \masters_01_ar_qos[1] ,
    \masters_01_ar_qos[0] }),
    .dbg_master_ar_region({\masters_01_ar_region[3] ,
    \masters_01_ar_region[2] ,
    \masters_01_ar_region[1] ,
    \masters_01_ar_region[0] }),
    .dbg_master_ar_size({\masters_01_ar_size[2] ,
    \masters_01_ar_size[1] ,
    \masters_01_ar_size[0] }),
    .dbg_master_ar_user({_NC707,
    _NC708}),
    .dbg_master_aw_addr({\masters_01_aw_addr[31] ,
    \masters_01_aw_addr[30] ,
    \masters_01_aw_addr[29] ,
    \masters_01_aw_addr[28] ,
    \masters_01_aw_addr[27] ,
    \masters_01_aw_addr[26] ,
    \masters_01_aw_addr[25] ,
    \masters_01_aw_addr[24] ,
    \masters_01_aw_addr[23] ,
    \masters_01_aw_addr[22] ,
    \masters_01_aw_addr[21] ,
    \masters_01_aw_addr[20] ,
    \masters_01_aw_addr[19] ,
    \masters_01_aw_addr[18] ,
    \masters_01_aw_addr[17] ,
    \masters_01_aw_addr[16] ,
    \masters_01_aw_addr[15] ,
    \masters_01_aw_addr[14] ,
    \masters_01_aw_addr[13] ,
    \masters_01_aw_addr[12] ,
    \masters_01_aw_addr[11] ,
    \masters_01_aw_addr[10] ,
    \masters_01_aw_addr[9] ,
    \masters_01_aw_addr[8] ,
    \masters_01_aw_addr[7] ,
    \masters_01_aw_addr[6] ,
    \masters_01_aw_addr[5] ,
    \masters_01_aw_addr[4] ,
    \masters_01_aw_addr[3] ,
    \masters_01_aw_addr[2] ,
    \masters_01_aw_addr[1] ,
    \masters_01_aw_addr[0] }),
    .dbg_master_aw_burst({\masters_01_aw_burst[1] ,
    \masters_01_aw_burst[0] }),
    .dbg_master_aw_cache({\masters_01_aw_cache[3] ,
    \masters_01_aw_cache[2] ,
    \masters_01_aw_cache[1] ,
    \masters_01_aw_cache[0] }),
    .dbg_master_aw_id({_NC709,
    _NC710,
    _NC711,
    _NC712,
    _NC713,
    _NC714,
    _NC715,
    _NC716,
    _NC717,
    _NC718}),
    .dbg_master_aw_len({\masters_01_aw_len[7] ,
    \masters_01_aw_len[6] ,
    \masters_01_aw_len[5] ,
    \masters_01_aw_len[4] ,
    \masters_01_aw_len[3] ,
    \masters_01_aw_len[2] ,
    \masters_01_aw_len[1] ,
    \masters_01_aw_len[0] }),
    .dbg_master_aw_prot({\masters_01_aw_prot[2] ,
    \masters_01_aw_prot[1] ,
    \masters_01_aw_prot[0] }),
    .dbg_master_aw_qos({\masters_01_aw_qos[3] ,
    \masters_01_aw_qos[2] ,
    \masters_01_aw_qos[1] ,
    \masters_01_aw_qos[0] }),
    .dbg_master_aw_region({\masters_01_aw_region[3] ,
    \masters_01_aw_region[2] ,
    \masters_01_aw_region[1] ,
    \masters_01_aw_region[0] }),
    .dbg_master_aw_size({\masters_01_aw_size[2] ,
    \masters_01_aw_size[1] ,
    \masters_01_aw_size[0] }),
    .dbg_master_aw_user({_NC719,
    _NC720}),
    .dbg_master_b_id({_NC721,
    _NC722,
    _NC723,
    _NC724,
    _NC725,
    _NC726,
    _NC727,
    _NC728,
    _NC729,
    _NC730}),
    .dbg_master_b_resp({\masters_01_b_resp[1] ,
    \masters_01_b_resp[0] }),
    .dbg_master_b_user({_NC731,
    _NC732}),
    .dbg_master_r_data({_NC733,
    _NC734,
    _NC735,
    _NC736,
    _NC737,
    _NC738,
    _NC739,
    _NC740,
    _NC741,
    _NC742,
    _NC743,
    _NC744,
    _NC745,
    _NC746,
    _NC747,
    _NC748,
    _NC749,
    _NC750,
    _NC751,
    _NC752,
    _NC753,
    _NC754,
    _NC755,
    _NC756,
    _NC757,
    _NC758,
    _NC759,
    _NC760,
    _NC761,
    _NC762,
    _NC763,
    _NC764,
    _NC765,
    _NC766,
    _NC767,
    _NC768,
    _NC769,
    _NC770,
    _NC771,
    _NC772,
    _NC773,
    _NC774,
    _NC775,
    _NC776,
    _NC777,
    _NC778,
    _NC779,
    _NC780,
    _NC781,
    _NC782,
    _NC783,
    _NC784,
    _NC785,
    _NC786,
    _NC787,
    _NC788,
    _NC789,
    _NC790,
    _NC791,
    _NC792,
    _NC793,
    _NC794,
    _NC795,
    _NC796}),
    .dbg_master_r_id({_NC797,
    _NC798,
    _NC799,
    _NC800,
    _NC801,
    _NC802,
    _NC803,
    _NC804,
    _NC805,
    _NC806}),
    .dbg_master_r_resp({\masters_01_r_resp[1] ,
    \masters_01_r_resp[0] }),
    .dbg_master_r_user({_NC807,
    _NC808}),
    .dbg_master_w_data({_NC809,
    _NC810,
    _NC811,
    _NC812,
    _NC813,
    _NC814,
    _NC815,
    _NC816,
    _NC817,
    _NC818,
    _NC819,
    _NC820,
    _NC821,
    _NC822,
    _NC823,
    _NC824,
    _NC825,
    _NC826,
    _NC827,
    _NC828,
    _NC829,
    _NC830,
    _NC831,
    _NC832,
    _NC833,
    _NC834,
    _NC835,
    _NC836,
    _NC837,
    _NC838,
    _NC839,
    _NC840,
    _NC841,
    _NC842,
    _NC843,
    _NC844,
    _NC845,
    _NC846,
    _NC847,
    _NC848,
    _NC849,
    _NC850,
    _NC851,
    _NC852,
    _NC853,
    _NC854,
    _NC855,
    _NC856,
    _NC857,
    _NC858,
    _NC859,
    _NC860,
    _NC861,
    _NC862,
    _NC863,
    _NC864,
    _NC865,
    _NC866,
    _NC867,
    _NC868,
    _NC869,
    _NC870,
    _NC871,
    _NC872}),
    .dbg_master_w_strb({_NC873,
    _NC874,
    _NC875,
    _NC876,
    _NC877,
    _NC878,
    _NC879,
    _NC880}),
    .dbg_master_w_user({_NC881,
    _NC882}),
    .debug_addr({\debug_addr[14] ,
    \debug_addr[13] ,
    \debug_addr[12] ,
    \debug_addr[11] ,
    \debug_addr[10] ,
    \debug_addr[9] ,
    \debug_addr[8] ,
    \debug_addr[7] ,
    \debug_addr[6] ,
    \debug_addr[5] ,
    \debug_addr[4] ,
    \debug_addr[3] ,
    \debug_addr[2] ,
    \debug_addr[1] ,
    \debug_addr[0] }),
    .debug_rdata({\debug_rdata[31] ,
    \debug_rdata[30] ,
    \debug_rdata[29] ,
    \debug_rdata[28] ,
    \debug_rdata[27] ,
    \debug_rdata[26] ,
    \debug_rdata[25] ,
    \debug_rdata[24] ,
    \debug_rdata[23] ,
    \debug_rdata[22] ,
    \debug_rdata[21] ,
    \debug_rdata[20] ,
    \debug_rdata[19] ,
    \debug_rdata[18] ,
    \debug_rdata[17] ,
    \debug_rdata[16] ,
    \debug_rdata[15] ,
    \debug_rdata[14] ,
    \debug_rdata[13] ,
    \debug_rdata[12] ,
    \debug_rdata[11] ,
    \debug_rdata[10] ,
    \debug_rdata[9] ,
    \debug_rdata[8] ,
    \debug_rdata[7] ,
    \debug_rdata[6] ,
    \debug_rdata[5] ,
    \debug_rdata[4] ,
    \debug_rdata[3] ,
    \debug_rdata[2] ,
    \debug_rdata[1] ,
    \debug_rdata[0] }),
    .debug_wdata({\debug_wdata[31] ,
    \debug_wdata[30] ,
    \debug_wdata[29] ,
    \debug_wdata[28] ,
    \debug_wdata[27] ,
    \debug_wdata[26] ,
    \debug_wdata[25] ,
    \debug_wdata[24] ,
    \debug_wdata[23] ,
    \debug_wdata[22] ,
    \debug_wdata[21] ,
    \debug_wdata[20] ,
    \debug_wdata[19] ,
    \debug_wdata[18] ,
    \debug_wdata[17] ,
    \debug_wdata[16] ,
    \debug_wdata[15] ,
    \debug_wdata[14] ,
    \debug_wdata[13] ,
    \debug_wdata[12] ,
    \debug_wdata[11] ,
    \debug_wdata[10] ,
    \debug_wdata[9] ,
    \debug_wdata[8] ,
    \debug_wdata[7] ,
    \debug_wdata[6] ,
    \debug_wdata[5] ,
    \debug_wdata[4] ,
    \debug_wdata[3] ,
    \debug_wdata[2] ,
    \debug_wdata[1] ,
    \debug_wdata[0] }),
    .instr_slave_ar_addr({\slaves_00_ar_addr[31] ,
    \slaves_00_ar_addr[30] ,
    \slaves_00_ar_addr[29] ,
    \slaves_00_ar_addr[28] ,
    \slaves_00_ar_addr[27] ,
    \slaves_00_ar_addr[26] ,
    \slaves_00_ar_addr[25] ,
    \slaves_00_ar_addr[24] ,
    \slaves_00_ar_addr[23] ,
    \slaves_00_ar_addr[22] ,
    \slaves_00_ar_addr[21] ,
    \slaves_00_ar_addr[20] ,
    \slaves_00_ar_addr[19] ,
    \slaves_00_ar_addr[18] ,
    \slaves_00_ar_addr[17] ,
    \slaves_00_ar_addr[16] ,
    \slaves_00_ar_addr[15] ,
    \slaves_00_ar_addr[14] ,
    \slaves_00_ar_addr[13] ,
    \slaves_00_ar_addr[12] ,
    \slaves_00_ar_addr[11] ,
    \slaves_00_ar_addr[10] ,
    \slaves_00_ar_addr[9] ,
    \slaves_00_ar_addr[8] ,
    \slaves_00_ar_addr[7] ,
    \slaves_00_ar_addr[6] ,
    \slaves_00_ar_addr[5] ,
    \slaves_00_ar_addr[4] ,
    \slaves_00_ar_addr[3] ,
    \slaves_00_ar_addr[2] ,
    \slaves_00_ar_addr[1] ,
    \slaves_00_ar_addr[0] }),
    .instr_slave_ar_burst({\slaves_00_ar_burst[1] ,
    \slaves_00_ar_burst[0] }),
    .instr_slave_ar_cache({\slaves_00_ar_cache[3] ,
    \slaves_00_ar_cache[2] ,
    \slaves_00_ar_cache[1] ,
    \slaves_00_ar_cache[0] }),
    .instr_slave_ar_id({_NC883,
    _NC884,
    _NC885,
    _NC886,
    _NC887,
    _NC888,
    _NC889,
    _NC890,
    _NC891,
    _NC892}),
    .instr_slave_ar_len({\slaves_00_ar_len[7] ,
    \slaves_00_ar_len[6] ,
    \slaves_00_ar_len[5] ,
    \slaves_00_ar_len[4] ,
    \slaves_00_ar_len[3] ,
    \slaves_00_ar_len[2] ,
    \slaves_00_ar_len[1] ,
    \slaves_00_ar_len[0] }),
    .instr_slave_ar_prot({\slaves_00_ar_prot[2] ,
    \slaves_00_ar_prot[1] ,
    \slaves_00_ar_prot[0] }),
    .instr_slave_ar_qos({\slaves_00_ar_qos[3] ,
    \slaves_00_ar_qos[2] ,
    \slaves_00_ar_qos[1] ,
    \slaves_00_ar_qos[0] }),
    .instr_slave_ar_region({\slaves_00_ar_region[3] ,
    \slaves_00_ar_region[2] ,
    \slaves_00_ar_region[1] ,
    \slaves_00_ar_region[0] }),
    .instr_slave_ar_size({\slaves_00_ar_size[2] ,
    \slaves_00_ar_size[1] ,
    \slaves_00_ar_size[0] }),
    .instr_slave_ar_user({_NC893,
    _NC894}),
    .instr_slave_aw_addr({\slaves_00_aw_addr[31] ,
    \slaves_00_aw_addr[30] ,
    \slaves_00_aw_addr[29] ,
    \slaves_00_aw_addr[28] ,
    \slaves_00_aw_addr[27] ,
    \slaves_00_aw_addr[26] ,
    \slaves_00_aw_addr[25] ,
    \slaves_00_aw_addr[24] ,
    \slaves_00_aw_addr[23] ,
    \slaves_00_aw_addr[22] ,
    \slaves_00_aw_addr[21] ,
    \slaves_00_aw_addr[20] ,
    \slaves_00_aw_addr[19] ,
    \slaves_00_aw_addr[18] ,
    \slaves_00_aw_addr[17] ,
    \slaves_00_aw_addr[16] ,
    \slaves_00_aw_addr[15] ,
    \slaves_00_aw_addr[14] ,
    \slaves_00_aw_addr[13] ,
    \slaves_00_aw_addr[12] ,
    \slaves_00_aw_addr[11] ,
    \slaves_00_aw_addr[10] ,
    \slaves_00_aw_addr[9] ,
    \slaves_00_aw_addr[8] ,
    \slaves_00_aw_addr[7] ,
    \slaves_00_aw_addr[6] ,
    \slaves_00_aw_addr[5] ,
    \slaves_00_aw_addr[4] ,
    \slaves_00_aw_addr[3] ,
    \slaves_00_aw_addr[2] ,
    \slaves_00_aw_addr[1] ,
    \slaves_00_aw_addr[0] }),
    .instr_slave_aw_burst({\slaves_00_aw_burst[1] ,
    \slaves_00_aw_burst[0] }),
    .instr_slave_aw_cache({\slaves_00_aw_cache[3] ,
    \slaves_00_aw_cache[2] ,
    \slaves_00_aw_cache[1] ,
    \slaves_00_aw_cache[0] }),
    .instr_slave_aw_id({_NC895,
    _NC896,
    _NC897,
    _NC898,
    _NC899,
    _NC900,
    _NC901,
    _NC902,
    _NC903,
    _NC904}),
    .instr_slave_aw_len({\slaves_00_aw_len[7] ,
    \slaves_00_aw_len[6] ,
    \slaves_00_aw_len[5] ,
    \slaves_00_aw_len[4] ,
    \slaves_00_aw_len[3] ,
    \slaves_00_aw_len[2] ,
    \slaves_00_aw_len[1] ,
    \slaves_00_aw_len[0] }),
    .instr_slave_aw_prot({\slaves_00_aw_prot[2] ,
    \slaves_00_aw_prot[1] ,
    \slaves_00_aw_prot[0] }),
    .instr_slave_aw_qos({\slaves_00_aw_qos[3] ,
    \slaves_00_aw_qos[2] ,
    \slaves_00_aw_qos[1] ,
    \slaves_00_aw_qos[0] }),
    .instr_slave_aw_region({\slaves_00_aw_region[3] ,
    \slaves_00_aw_region[2] ,
    \slaves_00_aw_region[1] ,
    \slaves_00_aw_region[0] }),
    .instr_slave_aw_size({\slaves_00_aw_size[2] ,
    \slaves_00_aw_size[1] ,
    \slaves_00_aw_size[0] }),
    .instr_slave_aw_user({_NC905,
    _NC906}),
    .instr_slave_b_id({_NC907,
    _NC908,
    _NC909,
    _NC910,
    _NC911,
    _NC912,
    _NC913,
    _NC914,
    _NC915,
    _NC916}),
    .instr_slave_b_resp({\slaves_00_b_resp[1] ,
    \slaves_00_b_resp[0] }),
    .instr_slave_b_user({_NC917,
    _NC918}),
    .instr_slave_r_data({_NC919,
    _NC920,
    _NC921,
    _NC922,
    _NC923,
    _NC924,
    _NC925,
    _NC926,
    _NC927,
    _NC928,
    _NC929,
    _NC930,
    _NC931,
    _NC932,
    _NC933,
    _NC934,
    _NC935,
    _NC936,
    _NC937,
    _NC938,
    _NC939,
    _NC940,
    _NC941,
    _NC942,
    _NC943,
    _NC944,
    _NC945,
    _NC946,
    _NC947,
    _NC948,
    _NC949,
    _NC950,
    _NC951,
    _NC952,
    _NC953,
    _NC954,
    _NC955,
    _NC956,
    _NC957,
    _NC958,
    _NC959,
    _NC960,
    _NC961,
    _NC962,
    _NC963,
    _NC964,
    _NC965,
    _NC966,
    _NC967,
    _NC968,
    _NC969,
    _NC970,
    _NC971,
    _NC972,
    _NC973,
    _NC974,
    _NC975,
    _NC976,
    _NC977,
    _NC978,
    _NC979,
    _NC980,
    _NC981,
    _NC982}),
    .instr_slave_r_id({_NC983,
    _NC984,
    _NC985,
    _NC986,
    _NC987,
    _NC988,
    _NC989,
    _NC990,
    _NC991,
    _NC992}),
    .instr_slave_r_resp({\slaves_00_r_resp[1] ,
    \slaves_00_r_resp[0] }),
    .instr_slave_r_user({_NC993,
    _NC994}),
    .instr_slave_w_data({_NC995,
    _NC996,
    _NC997,
    _NC998,
    _NC999,
    _NC1000,
    _NC1001,
    _NC1002,
    _NC1003,
    _NC1004,
    _NC1005,
    _NC1006,
    _NC1007,
    _NC1008,
    _NC1009,
    _NC1010,
    _NC1011,
    _NC1012,
    _NC1013,
    _NC1014,
    _NC1015,
    _NC1016,
    _NC1017,
    _NC1018,
    _NC1019,
    _NC1020,
    _NC1021,
    _NC1022,
    _NC1023,
    _NC1024,
    _NC1025,
    _NC1026,
    _NC1027,
    _NC1028,
    _NC1029,
    _NC1030,
    _NC1031,
    _NC1032,
    _NC1033,
    _NC1034,
    _NC1035,
    _NC1036,
    _NC1037,
    _NC1038,
    _NC1039,
    _NC1040,
    _NC1041,
    _NC1042,
    _NC1043,
    _NC1044,
    _NC1045,
    _NC1046,
    _NC1047,
    _NC1048,
    _NC1049,
    _NC1050,
    _NC1051,
    _NC1052,
    _NC1053,
    _NC1054,
    _NC1055,
    _NC1056,
    _NC1057,
    _NC1058}),
    .instr_slave_w_strb({_NC1059,
    _NC1060,
    _NC1061,
    _NC1062,
    _NC1063,
    _NC1064,
    _NC1065,
    _NC1066}),
    .instr_slave_w_user({_NC1067,
    _NC1068}),
    .irq_i({\irq_to_core_int[31] ,
    \irq_to_core_int[30] ,
    \irq_to_core_int[29] ,
    \irq_to_core_int[28] ,
    \irq_to_core_int[27] ,
    \irq_to_core_int[26] ,
    \irq_to_core_int[25] ,
    \irq_to_core_int[24] ,
    \irq_to_core_int[23] ,
    \irq_to_core_int[22] ,
    \irq_to_core_int[21] ,
    \irq_to_core_int[20] ,
    \irq_to_core_int[19] ,
    \irq_to_core_int[18] ,
    \irq_to_core_int[17] ,
    \irq_to_core_int[16] ,
    \irq_to_core_int[15] ,
    \irq_to_core_int[14] ,
    \irq_to_core_int[13] ,
    \irq_to_core_int[12] ,
    \irq_to_core_int[11] ,
    \irq_to_core_int[10] ,
    \irq_to_core_int[9] ,
    \irq_to_core_int[8] ,
    \irq_to_core_int[7] ,
    \irq_to_core_int[6] ,
    \irq_to_core_int[5] ,
    \irq_to_core_int[4] ,
    \irq_to_core_int[3] ,
    \irq_to_core_int[2] ,
    \irq_to_core_int[1] ,
    \irq_to_core_int[0] }),
    .mba_data_mem_addr0_o({\mba_data_mem_addr0_o[31] ,
    \mba_data_mem_addr0_o[30] ,
    \mba_data_mem_addr0_o[29] ,
    \mba_data_mem_addr0_o[28] ,
    \mba_data_mem_addr0_o[27] ,
    \mba_data_mem_addr0_o[26] ,
    \mba_data_mem_addr0_o[25] ,
    \mba_data_mem_addr0_o[24] ,
    \mba_data_mem_addr0_o[23] ,
    \mba_data_mem_addr0_o[22] ,
    \mba_data_mem_addr0_o[21] ,
    \mba_data_mem_addr0_o[20] ,
    \mba_data_mem_addr0_o[19] ,
    \mba_data_mem_addr0_o[18] ,
    \mba_data_mem_addr0_o[17] ,
    \mba_data_mem_addr0_o[16] ,
    \mba_data_mem_addr0_o[15] ,
    \mba_data_mem_addr0_o[14] ,
    \mba_data_mem_addr0_o[13] ,
    \mba_data_mem_addr0_o[12] ,
    \mba_data_mem_addr0_o[11] ,
    \mba_data_mem_addr0_o[10] ,
    \mba_data_mem_addr0_o[9] ,
    \mba_data_mem_addr0_o[8] ,
    \mba_data_mem_addr0_o[7] ,
    \mba_data_mem_addr0_o[6] ,
    \mba_data_mem_addr0_o[5] ,
    \mba_data_mem_addr0_o[4] ,
    \mba_data_mem_addr0_o[3] ,
    \mba_data_mem_addr0_o[2] ,
    \mba_data_mem_addr0_o[1] ,
    \mba_data_mem_addr0_o[0] }),
    .mba_data_mem_addr1_o({\mba_data_mem_addr1_o[31] ,
    \mba_data_mem_addr1_o[30] ,
    \mba_data_mem_addr1_o[29] ,
    \mba_data_mem_addr1_o[28] ,
    \mba_data_mem_addr1_o[27] ,
    \mba_data_mem_addr1_o[26] ,
    \mba_data_mem_addr1_o[25] ,
    \mba_data_mem_addr1_o[24] ,
    \mba_data_mem_addr1_o[23] ,
    \mba_data_mem_addr1_o[22] ,
    \mba_data_mem_addr1_o[21] ,
    \mba_data_mem_addr1_o[20] ,
    \mba_data_mem_addr1_o[19] ,
    \mba_data_mem_addr1_o[18] ,
    \mba_data_mem_addr1_o[17] ,
    \mba_data_mem_addr1_o[16] ,
    \mba_data_mem_addr1_o[15] ,
    \mba_data_mem_addr1_o[14] ,
    \mba_data_mem_addr1_o[13] ,
    \mba_data_mem_addr1_o[12] ,
    \mba_data_mem_addr1_o[11] ,
    \mba_data_mem_addr1_o[10] ,
    \mba_data_mem_addr1_o[9] ,
    \mba_data_mem_addr1_o[8] ,
    \mba_data_mem_addr1_o[7] ,
    \mba_data_mem_addr1_o[6] ,
    \mba_data_mem_addr1_o[5] ,
    \mba_data_mem_addr1_o[4] ,
    \mba_data_mem_addr1_o[3] ,
    \mba_data_mem_addr1_o[2] ,
    \mba_data_mem_addr1_o[1] ,
    \mba_data_mem_addr1_o[0] }),
    .mba_data_mem_din0_o({\mba_data_mem_din0_o[31] ,
    \mba_data_mem_din0_o[30] ,
    \mba_data_mem_din0_o[29] ,
    \mba_data_mem_din0_o[28] ,
    \mba_data_mem_din0_o[27] ,
    \mba_data_mem_din0_o[26] ,
    \mba_data_mem_din0_o[25] ,
    \mba_data_mem_din0_o[24] ,
    \mba_data_mem_din0_o[23] ,
    \mba_data_mem_din0_o[22] ,
    \mba_data_mem_din0_o[21] ,
    \mba_data_mem_din0_o[20] ,
    \mba_data_mem_din0_o[19] ,
    \mba_data_mem_din0_o[18] ,
    \mba_data_mem_din0_o[17] ,
    \mba_data_mem_din0_o[16] ,
    \mba_data_mem_din0_o[15] ,
    \mba_data_mem_din0_o[14] ,
    \mba_data_mem_din0_o[13] ,
    \mba_data_mem_din0_o[12] ,
    \mba_data_mem_din0_o[11] ,
    \mba_data_mem_din0_o[10] ,
    \mba_data_mem_din0_o[9] ,
    \mba_data_mem_din0_o[8] ,
    \mba_data_mem_din0_o[7] ,
    \mba_data_mem_din0_o[6] ,
    \mba_data_mem_din0_o[5] ,
    \mba_data_mem_din0_o[4] ,
    \mba_data_mem_din0_o[3] ,
    \mba_data_mem_din0_o[2] ,
    \mba_data_mem_din0_o[1] ,
    \mba_data_mem_din0_o[0] }),
    .mba_data_mem_dout0_i({\mba_data_mem_dout0_i[31] ,
    \mba_data_mem_dout0_i[30] ,
    \mba_data_mem_dout0_i[29] ,
    \mba_data_mem_dout0_i[28] ,
    \mba_data_mem_dout0_i[27] ,
    \mba_data_mem_dout0_i[26] ,
    \mba_data_mem_dout0_i[25] ,
    \mba_data_mem_dout0_i[24] ,
    \mba_data_mem_dout0_i[23] ,
    \mba_data_mem_dout0_i[22] ,
    \mba_data_mem_dout0_i[21] ,
    \mba_data_mem_dout0_i[20] ,
    \mba_data_mem_dout0_i[19] ,
    \mba_data_mem_dout0_i[18] ,
    \mba_data_mem_dout0_i[17] ,
    \mba_data_mem_dout0_i[16] ,
    \mba_data_mem_dout0_i[15] ,
    \mba_data_mem_dout0_i[14] ,
    \mba_data_mem_dout0_i[13] ,
    \mba_data_mem_dout0_i[12] ,
    \mba_data_mem_dout0_i[11] ,
    \mba_data_mem_dout0_i[10] ,
    \mba_data_mem_dout0_i[9] ,
    \mba_data_mem_dout0_i[8] ,
    \mba_data_mem_dout0_i[7] ,
    \mba_data_mem_dout0_i[6] ,
    \mba_data_mem_dout0_i[5] ,
    \mba_data_mem_dout0_i[4] ,
    \mba_data_mem_dout0_i[3] ,
    \mba_data_mem_dout0_i[2] ,
    \mba_data_mem_dout0_i[1] ,
    \mba_data_mem_dout0_i[0] }),
    .mba_data_mem_wmask0_o({\mba_data_mem_wmask0_o[3] ,
    \mba_data_mem_wmask0_o[2] ,
    \mba_data_mem_wmask0_o[1] ,
    \mba_data_mem_wmask0_o[0] }),
    .mba_instr_mem_addr0_o({\mba_instr_mem_addr0_o[31] ,
    \mba_instr_mem_addr0_o[30] ,
    \mba_instr_mem_addr0_o[29] ,
    \mba_instr_mem_addr0_o[28] ,
    \mba_instr_mem_addr0_o[27] ,
    \mba_instr_mem_addr0_o[26] ,
    \mba_instr_mem_addr0_o[25] ,
    \mba_instr_mem_addr0_o[24] ,
    \mba_instr_mem_addr0_o[23] ,
    \mba_instr_mem_addr0_o[22] ,
    \mba_instr_mem_addr0_o[21] ,
    \mba_instr_mem_addr0_o[20] ,
    \mba_instr_mem_addr0_o[19] ,
    \mba_instr_mem_addr0_o[18] ,
    \mba_instr_mem_addr0_o[17] ,
    \mba_instr_mem_addr0_o[16] ,
    \mba_instr_mem_addr0_o[15] ,
    \mba_instr_mem_addr0_o[14] ,
    \mba_instr_mem_addr0_o[13] ,
    \mba_instr_mem_addr0_o[12] ,
    \mba_instr_mem_addr0_o[11] ,
    \mba_instr_mem_addr0_o[10] ,
    \mba_instr_mem_addr0_o[9] ,
    \mba_instr_mem_addr0_o[8] ,
    \mba_instr_mem_addr0_o[7] ,
    \mba_instr_mem_addr0_o[6] ,
    \mba_instr_mem_addr0_o[5] ,
    \mba_instr_mem_addr0_o[4] ,
    \mba_instr_mem_addr0_o[3] ,
    \mba_instr_mem_addr0_o[2] ,
    \mba_instr_mem_addr0_o[1] ,
    \mba_instr_mem_addr0_o[0] }),
    .mba_instr_mem_addr1_o({\mba_instr_mem_addr1_o[31] ,
    \mba_instr_mem_addr1_o[30] ,
    \mba_instr_mem_addr1_o[29] ,
    \mba_instr_mem_addr1_o[28] ,
    \mba_instr_mem_addr1_o[27] ,
    \mba_instr_mem_addr1_o[26] ,
    \mba_instr_mem_addr1_o[25] ,
    \mba_instr_mem_addr1_o[24] ,
    \mba_instr_mem_addr1_o[23] ,
    \mba_instr_mem_addr1_o[22] ,
    \mba_instr_mem_addr1_o[21] ,
    \mba_instr_mem_addr1_o[20] ,
    \mba_instr_mem_addr1_o[19] ,
    \mba_instr_mem_addr1_o[18] ,
    \mba_instr_mem_addr1_o[17] ,
    \mba_instr_mem_addr1_o[16] ,
    \mba_instr_mem_addr1_o[15] ,
    \mba_instr_mem_addr1_o[14] ,
    \mba_instr_mem_addr1_o[13] ,
    \mba_instr_mem_addr1_o[12] ,
    \mba_instr_mem_addr1_o[11] ,
    \mba_instr_mem_addr1_o[10] ,
    \mba_instr_mem_addr1_o[9] ,
    \mba_instr_mem_addr1_o[8] ,
    \mba_instr_mem_addr1_o[7] ,
    \mba_instr_mem_addr1_o[6] ,
    \mba_instr_mem_addr1_o[5] ,
    \mba_instr_mem_addr1_o[4] ,
    \mba_instr_mem_addr1_o[3] ,
    \mba_instr_mem_addr1_o[2] ,
    \mba_instr_mem_addr1_o[1] ,
    \mba_instr_mem_addr1_o[0] }),
    .mba_instr_mem_din0_o({\mba_instr_mem_din0_o[31] ,
    \mba_instr_mem_din0_o[30] ,
    \mba_instr_mem_din0_o[29] ,
    \mba_instr_mem_din0_o[28] ,
    \mba_instr_mem_din0_o[27] ,
    \mba_instr_mem_din0_o[26] ,
    \mba_instr_mem_din0_o[25] ,
    \mba_instr_mem_din0_o[24] ,
    \mba_instr_mem_din0_o[23] ,
    \mba_instr_mem_din0_o[22] ,
    \mba_instr_mem_din0_o[21] ,
    \mba_instr_mem_din0_o[20] ,
    \mba_instr_mem_din0_o[19] ,
    \mba_instr_mem_din0_o[18] ,
    \mba_instr_mem_din0_o[17] ,
    \mba_instr_mem_din0_o[16] ,
    \mba_instr_mem_din0_o[15] ,
    \mba_instr_mem_din0_o[14] ,
    \mba_instr_mem_din0_o[13] ,
    \mba_instr_mem_din0_o[12] ,
    \mba_instr_mem_din0_o[11] ,
    \mba_instr_mem_din0_o[10] ,
    \mba_instr_mem_din0_o[9] ,
    \mba_instr_mem_din0_o[8] ,
    \mba_instr_mem_din0_o[7] ,
    \mba_instr_mem_din0_o[6] ,
    \mba_instr_mem_din0_o[5] ,
    \mba_instr_mem_din0_o[4] ,
    \mba_instr_mem_din0_o[3] ,
    \mba_instr_mem_din0_o[2] ,
    \mba_instr_mem_din0_o[1] ,
    \mba_instr_mem_din0_o[0] }),
    .mba_instr_mem_dout0_i({\mba_instr_mem_dout0_i[31] ,
    \mba_instr_mem_dout0_i[30] ,
    \mba_instr_mem_dout0_i[29] ,
    \mba_instr_mem_dout0_i[28] ,
    \mba_instr_mem_dout0_i[27] ,
    \mba_instr_mem_dout0_i[26] ,
    \mba_instr_mem_dout0_i[25] ,
    \mba_instr_mem_dout0_i[24] ,
    \mba_instr_mem_dout0_i[23] ,
    \mba_instr_mem_dout0_i[22] ,
    \mba_instr_mem_dout0_i[21] ,
    \mba_instr_mem_dout0_i[20] ,
    \mba_instr_mem_dout0_i[19] ,
    \mba_instr_mem_dout0_i[18] ,
    \mba_instr_mem_dout0_i[17] ,
    \mba_instr_mem_dout0_i[16] ,
    \mba_instr_mem_dout0_i[15] ,
    \mba_instr_mem_dout0_i[14] ,
    \mba_instr_mem_dout0_i[13] ,
    \mba_instr_mem_dout0_i[12] ,
    \mba_instr_mem_dout0_i[11] ,
    \mba_instr_mem_dout0_i[10] ,
    \mba_instr_mem_dout0_i[9] ,
    \mba_instr_mem_dout0_i[8] ,
    \mba_instr_mem_dout0_i[7] ,
    \mba_instr_mem_dout0_i[6] ,
    \mba_instr_mem_dout0_i[5] ,
    \mba_instr_mem_dout0_i[4] ,
    \mba_instr_mem_dout0_i[3] ,
    \mba_instr_mem_dout0_i[2] ,
    \mba_instr_mem_dout0_i[1] ,
    \mba_instr_mem_dout0_i[0] }),
    .mba_instr_mem_wmask0_o({\mba_instr_mem_wmask0_o[3] ,
    \mba_instr_mem_wmask0_o[2] ,
    \mba_instr_mem_wmask0_o[1] ,
    \mba_instr_mem_wmask0_o[0] }));
 sky130_sram_2kbyte_1rw1r_32x512_8 data_ram (.csb0(mba_data_mem_csb0_o),
    .csb1(mba_data_mem_csb1_o),
    .web0(mba_data_mem_web0_o),
    .clk0(clk_int),
    .clk1(io_in[21]),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .addr0({\mba_data_mem_addr0_o[10] ,
    \mba_data_mem_addr0_o[9] ,
    \mba_data_mem_addr0_o[8] ,
    \mba_data_mem_addr0_o[7] ,
    \mba_data_mem_addr0_o[6] ,
    \mba_data_mem_addr0_o[5] ,
    \mba_data_mem_addr0_o[4] ,
    \mba_data_mem_addr0_o[3] ,
    \mba_data_mem_addr0_o[2] }),
    .addr1({\mba_data_mem_addr1_o[10] ,
    \mba_data_mem_addr1_o[9] ,
    \mba_data_mem_addr1_o[8] ,
    \mba_data_mem_addr1_o[7] ,
    \mba_data_mem_addr1_o[6] ,
    \mba_data_mem_addr1_o[5] ,
    \mba_data_mem_addr1_o[4] ,
    \mba_data_mem_addr1_o[3] ,
    \mba_data_mem_addr1_o[2] }),
    .din0({\mba_data_mem_din0_o[31] ,
    \mba_data_mem_din0_o[30] ,
    \mba_data_mem_din0_o[29] ,
    \mba_data_mem_din0_o[28] ,
    \mba_data_mem_din0_o[27] ,
    \mba_data_mem_din0_o[26] ,
    \mba_data_mem_din0_o[25] ,
    \mba_data_mem_din0_o[24] ,
    \mba_data_mem_din0_o[23] ,
    \mba_data_mem_din0_o[22] ,
    \mba_data_mem_din0_o[21] ,
    \mba_data_mem_din0_o[20] ,
    \mba_data_mem_din0_o[19] ,
    \mba_data_mem_din0_o[18] ,
    \mba_data_mem_din0_o[17] ,
    \mba_data_mem_din0_o[16] ,
    \mba_data_mem_din0_o[15] ,
    \mba_data_mem_din0_o[14] ,
    \mba_data_mem_din0_o[13] ,
    \mba_data_mem_din0_o[12] ,
    \mba_data_mem_din0_o[11] ,
    \mba_data_mem_din0_o[10] ,
    \mba_data_mem_din0_o[9] ,
    \mba_data_mem_din0_o[8] ,
    \mba_data_mem_din0_o[7] ,
    \mba_data_mem_din0_o[6] ,
    \mba_data_mem_din0_o[5] ,
    \mba_data_mem_din0_o[4] ,
    \mba_data_mem_din0_o[3] ,
    \mba_data_mem_din0_o[2] ,
    \mba_data_mem_din0_o[1] ,
    \mba_data_mem_din0_o[0] }),
    .dout0({\mba_data_mem_dout0_i[31] ,
    \mba_data_mem_dout0_i[30] ,
    \mba_data_mem_dout0_i[29] ,
    \mba_data_mem_dout0_i[28] ,
    \mba_data_mem_dout0_i[27] ,
    \mba_data_mem_dout0_i[26] ,
    \mba_data_mem_dout0_i[25] ,
    \mba_data_mem_dout0_i[24] ,
    \mba_data_mem_dout0_i[23] ,
    \mba_data_mem_dout0_i[22] ,
    \mba_data_mem_dout0_i[21] ,
    \mba_data_mem_dout0_i[20] ,
    \mba_data_mem_dout0_i[19] ,
    \mba_data_mem_dout0_i[18] ,
    \mba_data_mem_dout0_i[17] ,
    \mba_data_mem_dout0_i[16] ,
    \mba_data_mem_dout0_i[15] ,
    \mba_data_mem_dout0_i[14] ,
    \mba_data_mem_dout0_i[13] ,
    \mba_data_mem_dout0_i[12] ,
    \mba_data_mem_dout0_i[11] ,
    \mba_data_mem_dout0_i[10] ,
    \mba_data_mem_dout0_i[9] ,
    \mba_data_mem_dout0_i[8] ,
    \mba_data_mem_dout0_i[7] ,
    \mba_data_mem_dout0_i[6] ,
    \mba_data_mem_dout0_i[5] ,
    \mba_data_mem_dout0_i[4] ,
    \mba_data_mem_dout0_i[3] ,
    \mba_data_mem_dout0_i[2] ,
    \mba_data_mem_dout0_i[1] ,
    \mba_data_mem_dout0_i[0] }),
    .dout1({\data_ram_dout1[31] ,
    \data_ram_dout1[30] ,
    \data_ram_dout1[29] ,
    \data_ram_dout1[28] ,
    \data_ram_dout1[27] ,
    \data_ram_dout1[26] ,
    \data_ram_dout1[25] ,
    \data_ram_dout1[24] ,
    \data_ram_dout1[23] ,
    \data_ram_dout1[22] ,
    \data_ram_dout1[21] ,
    \data_ram_dout1[20] ,
    \data_ram_dout1[19] ,
    \data_ram_dout1[18] ,
    \data_ram_dout1[17] ,
    \data_ram_dout1[16] ,
    \data_ram_dout1[15] ,
    \data_ram_dout1[14] ,
    \data_ram_dout1[13] ,
    \data_ram_dout1[12] ,
    \data_ram_dout1[11] ,
    \data_ram_dout1[10] ,
    \data_ram_dout1[9] ,
    \data_ram_dout1[8] ,
    \data_ram_dout1[7] ,
    \data_ram_dout1[6] ,
    \data_ram_dout1[5] ,
    \data_ram_dout1[4] ,
    \data_ram_dout1[3] ,
    \data_ram_dout1[2] ,
    \data_ram_dout1[1] ,
    \data_ram_dout1[0] }),
    .wmask0({\mba_data_mem_wmask0_o[3] ,
    \mba_data_mem_wmask0_o[2] ,
    \mba_data_mem_wmask0_o[1] ,
    \mba_data_mem_wmask0_o[0] }));
 sky130_sram_2kbyte_1rw1r_32x512_8 instr_ram (.csb0(mba_instr_mem_csb0_o),
    .csb1(mba_instr_mem_csb1_o),
    .web0(mba_instr_mem_web0_o),
    .clk0(clk_int),
    .clk1(io_in[21]),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .addr0({\mba_instr_mem_addr0_o[10] ,
    \mba_instr_mem_addr0_o[9] ,
    \mba_instr_mem_addr0_o[8] ,
    \mba_instr_mem_addr0_o[7] ,
    \mba_instr_mem_addr0_o[6] ,
    \mba_instr_mem_addr0_o[5] ,
    \mba_instr_mem_addr0_o[4] ,
    \mba_instr_mem_addr0_o[3] ,
    \mba_instr_mem_addr0_o[2] }),
    .addr1({\mba_instr_mem_addr1_o[10] ,
    \mba_instr_mem_addr1_o[9] ,
    \mba_instr_mem_addr1_o[8] ,
    \mba_instr_mem_addr1_o[7] ,
    \mba_instr_mem_addr1_o[6] ,
    \mba_instr_mem_addr1_o[5] ,
    \mba_instr_mem_addr1_o[4] ,
    \mba_instr_mem_addr1_o[3] ,
    \mba_instr_mem_addr1_o[2] }),
    .din0({\mba_instr_mem_din0_o[31] ,
    \mba_instr_mem_din0_o[30] ,
    \mba_instr_mem_din0_o[29] ,
    \mba_instr_mem_din0_o[28] ,
    \mba_instr_mem_din0_o[27] ,
    \mba_instr_mem_din0_o[26] ,
    \mba_instr_mem_din0_o[25] ,
    \mba_instr_mem_din0_o[24] ,
    \mba_instr_mem_din0_o[23] ,
    \mba_instr_mem_din0_o[22] ,
    \mba_instr_mem_din0_o[21] ,
    \mba_instr_mem_din0_o[20] ,
    \mba_instr_mem_din0_o[19] ,
    \mba_instr_mem_din0_o[18] ,
    \mba_instr_mem_din0_o[17] ,
    \mba_instr_mem_din0_o[16] ,
    \mba_instr_mem_din0_o[15] ,
    \mba_instr_mem_din0_o[14] ,
    \mba_instr_mem_din0_o[13] ,
    \mba_instr_mem_din0_o[12] ,
    \mba_instr_mem_din0_o[11] ,
    \mba_instr_mem_din0_o[10] ,
    \mba_instr_mem_din0_o[9] ,
    \mba_instr_mem_din0_o[8] ,
    \mba_instr_mem_din0_o[7] ,
    \mba_instr_mem_din0_o[6] ,
    \mba_instr_mem_din0_o[5] ,
    \mba_instr_mem_din0_o[4] ,
    \mba_instr_mem_din0_o[3] ,
    \mba_instr_mem_din0_o[2] ,
    \mba_instr_mem_din0_o[1] ,
    \mba_instr_mem_din0_o[0] }),
    .dout0({\mba_instr_mem_dout0_i[31] ,
    \mba_instr_mem_dout0_i[30] ,
    \mba_instr_mem_dout0_i[29] ,
    \mba_instr_mem_dout0_i[28] ,
    \mba_instr_mem_dout0_i[27] ,
    \mba_instr_mem_dout0_i[26] ,
    \mba_instr_mem_dout0_i[25] ,
    \mba_instr_mem_dout0_i[24] ,
    \mba_instr_mem_dout0_i[23] ,
    \mba_instr_mem_dout0_i[22] ,
    \mba_instr_mem_dout0_i[21] ,
    \mba_instr_mem_dout0_i[20] ,
    \mba_instr_mem_dout0_i[19] ,
    \mba_instr_mem_dout0_i[18] ,
    \mba_instr_mem_dout0_i[17] ,
    \mba_instr_mem_dout0_i[16] ,
    \mba_instr_mem_dout0_i[15] ,
    \mba_instr_mem_dout0_i[14] ,
    \mba_instr_mem_dout0_i[13] ,
    \mba_instr_mem_dout0_i[12] ,
    \mba_instr_mem_dout0_i[11] ,
    \mba_instr_mem_dout0_i[10] ,
    \mba_instr_mem_dout0_i[9] ,
    \mba_instr_mem_dout0_i[8] ,
    \mba_instr_mem_dout0_i[7] ,
    \mba_instr_mem_dout0_i[6] ,
    \mba_instr_mem_dout0_i[5] ,
    \mba_instr_mem_dout0_i[4] ,
    \mba_instr_mem_dout0_i[3] ,
    \mba_instr_mem_dout0_i[2] ,
    \mba_instr_mem_dout0_i[1] ,
    \mba_instr_mem_dout0_i[0] }),
    .dout1({\instr_ram_dout1[31] ,
    \instr_ram_dout1[30] ,
    \instr_ram_dout1[29] ,
    \instr_ram_dout1[28] ,
    \instr_ram_dout1[27] ,
    \instr_ram_dout1[26] ,
    \instr_ram_dout1[25] ,
    \instr_ram_dout1[24] ,
    \instr_ram_dout1[23] ,
    \instr_ram_dout1[22] ,
    \instr_ram_dout1[21] ,
    \instr_ram_dout1[20] ,
    \instr_ram_dout1[19] ,
    \instr_ram_dout1[18] ,
    \instr_ram_dout1[17] ,
    \instr_ram_dout1[16] ,
    \instr_ram_dout1[15] ,
    \instr_ram_dout1[14] ,
    \instr_ram_dout1[13] ,
    \instr_ram_dout1[12] ,
    \instr_ram_dout1[11] ,
    \instr_ram_dout1[10] ,
    \instr_ram_dout1[9] ,
    \instr_ram_dout1[8] ,
    \instr_ram_dout1[7] ,
    \instr_ram_dout1[6] ,
    \instr_ram_dout1[5] ,
    \instr_ram_dout1[4] ,
    \instr_ram_dout1[3] ,
    \instr_ram_dout1[2] ,
    \instr_ram_dout1[1] ,
    \instr_ram_dout1[0] }),
    .wmask0({\mba_instr_mem_wmask0_o[3] ,
    \mba_instr_mem_wmask0_o[2] ,
    \mba_instr_mem_wmask0_o[1] ,
    \mba_instr_mem_wmask0_o[0] }));
 peripherals peripherals_i (.axi_spi_master_ar_lock(masters_02_ar_lock),
    .axi_spi_master_ar_ready(masters_02_ar_ready),
    .axi_spi_master_ar_valid(masters_02_ar_valid),
    .axi_spi_master_aw_lock(masters_02_aw_lock),
    .axi_spi_master_aw_ready(masters_02_aw_ready),
    .axi_spi_master_aw_valid(masters_02_aw_valid),
    .axi_spi_master_b_ready(masters_02_b_ready),
    .axi_spi_master_b_valid(masters_02_b_valid),
    .axi_spi_master_r_last(masters_02_r_last),
    .axi_spi_master_r_ready(masters_02_r_ready),
    .axi_spi_master_r_valid(masters_02_r_valid),
    .axi_spi_master_w_last(masters_02_w_last),
    .axi_spi_master_w_ready(masters_02_w_ready),
    .axi_spi_master_w_valid(masters_02_w_valid),
    .clk_gate_core_o(clk_gate_core_int),
    .clk_i(clk_int),
    .clk_i_pll(user_clock2),
    .clk_o_pll(clk_int),
    .clk_sel_i_pll(la_data_in[0]),
    .clk_standalone_i_pll(la_data_in[1]),
    .core_busy_i(core_busy_int),
    .debug_gnt(debug_gnt),
    .debug_req(debug_req),
    .debug_rvalid(debug_rvalid),
    .debug_we(debug_we),
    .fetch_enable_i(la_data_in[6]),
    .fetch_enable_o(fetch_enable_int),
    .fll1_ack_i(cfgack_fll_int),
    .fll1_lock_i(lock_fll_int),
    .fll1_req_o(cfgreq_fll_int),
    .fll1_wrn_o(cfgweb_n_fll_int),
    .fll_ack_o_pll(cfgack_fll_int),
    .fll_lock_o_pll(lock_fll_int),
    .fll_req_i_pll(cfgreq_fll_int),
    .fll_wrn_i_pll(cfgweb_n_fll_int),
    .rst_n(rstn_int),
    .rstn_i_pll(wb_rst_i),
    .rstn_o_pll(rstn_int),
    .scan_en_i_pll(la_data_in[3]),
    .scan_i_pll(io_in[21]),
    .scan_o_pll(scan_o),
    .scl_pad_i(io_in[22]),
    .scl_pad_o(io_out[28]),
    .scl_padoen_o(scl_padoen_o),
    .sda_pad_i(io_in[23]),
    .sda_pad_o(io_out[27]),
    .sda_padoen_o(sda_padoen_o),
    .slave_ar_lock(slaves_02_ar_lock),
    .slave_ar_ready(slaves_02_ar_ready),
    .slave_ar_valid(slaves_02_ar_valid),
    .slave_aw_lock(slaves_02_aw_lock),
    .slave_aw_ready(slaves_02_aw_ready),
    .slave_aw_valid(slaves_02_aw_valid),
    .slave_b_ready(slaves_02_b_ready),
    .slave_b_valid(slaves_02_b_valid),
    .slave_r_last(slaves_02_r_last),
    .slave_r_ready(slaves_02_r_ready),
    .slave_r_valid(slaves_02_r_valid),
    .slave_w_last(slaves_02_w_last),
    .slave_w_ready(slaves_02_w_ready),
    .slave_w_valid(slaves_02_w_valid),
    .spi_clk_i(io_in[17]),
    .spi_cs_i(io_in[18]),
    .spi_master_clk(io_out[33]),
    .spi_master_csn0(io_out[32]),
    .spi_master_csn1(spi_master_csn1),
    .spi_master_csn2(spi_master_csn2),
    .spi_master_csn3(spi_master_csn3),
    .spi_master_sdi0(io_in[21]),
    .spi_master_sdi1(io_in[21]),
    .spi_master_sdi2(io_in[21]),
    .spi_master_sdi3(io_in[21]),
    .spi_master_sdo0(io_out[29]),
    .spi_master_sdo1(spi_master_sdo1),
    .spi_master_sdo2(spi_master_sdo2),
    .spi_master_sdo3(spi_master_sdo3),
    .spi_sdi0_i(io_in[19]),
    .spi_sdi1_i(io_in[21]),
    .spi_sdi2_i(io_in[21]),
    .spi_sdi3_i(io_in[21]),
    .spi_sdo0_o(io_out[35]),
    .spi_sdo1_o(spi_sdo1_o),
    .spi_sdo2_o(spi_sdo2_o),
    .spi_sdo3_o(spi_sdo3_o),
    .testmode_i(la_data_in[2]),
    .testmode_i_pll(la_data_in[2]),
    .uart_cts(la_data_in[4]),
    .uart_dsr(la_data_in[5]),
    .uart_dtr(uart_dtr),
    .uart_rts(uart_rts),
    .uart_rx(io_in[20]),
    .uart_tx(io_out[34]),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .wbs_ack_o_pll(wbs_ack_o),
    .axi_spi_master_ar_addr({\masters_02_ar_addr[31] ,
    \masters_02_ar_addr[30] ,
    \masters_02_ar_addr[29] ,
    \masters_02_ar_addr[28] ,
    \masters_02_ar_addr[27] ,
    \masters_02_ar_addr[26] ,
    \masters_02_ar_addr[25] ,
    \masters_02_ar_addr[24] ,
    \masters_02_ar_addr[23] ,
    \masters_02_ar_addr[22] ,
    \masters_02_ar_addr[21] ,
    \masters_02_ar_addr[20] ,
    \masters_02_ar_addr[19] ,
    \masters_02_ar_addr[18] ,
    \masters_02_ar_addr[17] ,
    \masters_02_ar_addr[16] ,
    \masters_02_ar_addr[15] ,
    \masters_02_ar_addr[14] ,
    \masters_02_ar_addr[13] ,
    \masters_02_ar_addr[12] ,
    \masters_02_ar_addr[11] ,
    \masters_02_ar_addr[10] ,
    \masters_02_ar_addr[9] ,
    \masters_02_ar_addr[8] ,
    \masters_02_ar_addr[7] ,
    \masters_02_ar_addr[6] ,
    \masters_02_ar_addr[5] ,
    \masters_02_ar_addr[4] ,
    \masters_02_ar_addr[3] ,
    \masters_02_ar_addr[2] ,
    \masters_02_ar_addr[1] ,
    \masters_02_ar_addr[0] }),
    .axi_spi_master_ar_burst({\masters_02_ar_burst[1] ,
    \masters_02_ar_burst[0] }),
    .axi_spi_master_ar_cache({\masters_02_ar_cache[3] ,
    \masters_02_ar_cache[2] ,
    \masters_02_ar_cache[1] ,
    \masters_02_ar_cache[0] }),
    .axi_spi_master_ar_id({_NC1069,
    _NC1070,
    _NC1071,
    _NC1072,
    _NC1073,
    _NC1074}),
    .axi_spi_master_ar_len({\masters_02_ar_len[7] ,
    \masters_02_ar_len[6] ,
    \masters_02_ar_len[5] ,
    \masters_02_ar_len[4] ,
    \masters_02_ar_len[3] ,
    \masters_02_ar_len[2] ,
    \masters_02_ar_len[1] ,
    \masters_02_ar_len[0] }),
    .axi_spi_master_ar_prot({\masters_02_ar_prot[2] ,
    \masters_02_ar_prot[1] ,
    \masters_02_ar_prot[0] }),
    .axi_spi_master_ar_qos({\masters_02_ar_qos[3] ,
    \masters_02_ar_qos[2] ,
    \masters_02_ar_qos[1] ,
    \masters_02_ar_qos[0] }),
    .axi_spi_master_ar_region({\masters_02_ar_region[3] ,
    \masters_02_ar_region[2] ,
    \masters_02_ar_region[1] ,
    \masters_02_ar_region[0] }),
    .axi_spi_master_ar_size({\masters_02_ar_size[2] ,
    \masters_02_ar_size[1] ,
    \masters_02_ar_size[0] }),
    .axi_spi_master_ar_user({_NC1075,
    _NC1076,
    _NC1077,
    _NC1078,
    _NC1079,
    _NC1080}),
    .axi_spi_master_aw_addr({\masters_02_aw_addr[31] ,
    \masters_02_aw_addr[30] ,
    \masters_02_aw_addr[29] ,
    \masters_02_aw_addr[28] ,
    \masters_02_aw_addr[27] ,
    \masters_02_aw_addr[26] ,
    \masters_02_aw_addr[25] ,
    \masters_02_aw_addr[24] ,
    \masters_02_aw_addr[23] ,
    \masters_02_aw_addr[22] ,
    \masters_02_aw_addr[21] ,
    \masters_02_aw_addr[20] ,
    \masters_02_aw_addr[19] ,
    \masters_02_aw_addr[18] ,
    \masters_02_aw_addr[17] ,
    \masters_02_aw_addr[16] ,
    \masters_02_aw_addr[15] ,
    \masters_02_aw_addr[14] ,
    \masters_02_aw_addr[13] ,
    \masters_02_aw_addr[12] ,
    \masters_02_aw_addr[11] ,
    \masters_02_aw_addr[10] ,
    \masters_02_aw_addr[9] ,
    \masters_02_aw_addr[8] ,
    \masters_02_aw_addr[7] ,
    \masters_02_aw_addr[6] ,
    \masters_02_aw_addr[5] ,
    \masters_02_aw_addr[4] ,
    \masters_02_aw_addr[3] ,
    \masters_02_aw_addr[2] ,
    \masters_02_aw_addr[1] ,
    \masters_02_aw_addr[0] }),
    .axi_spi_master_aw_burst({\masters_02_aw_burst[1] ,
    \masters_02_aw_burst[0] }),
    .axi_spi_master_aw_cache({\masters_02_aw_cache[3] ,
    \masters_02_aw_cache[2] ,
    \masters_02_aw_cache[1] ,
    \masters_02_aw_cache[0] }),
    .axi_spi_master_aw_id({_NC1081,
    _NC1082,
    _NC1083,
    _NC1084,
    _NC1085,
    _NC1086}),
    .axi_spi_master_aw_len({\masters_02_aw_len[7] ,
    \masters_02_aw_len[6] ,
    \masters_02_aw_len[5] ,
    \masters_02_aw_len[4] ,
    \masters_02_aw_len[3] ,
    \masters_02_aw_len[2] ,
    \masters_02_aw_len[1] ,
    \masters_02_aw_len[0] }),
    .axi_spi_master_aw_prot({\masters_02_aw_prot[2] ,
    \masters_02_aw_prot[1] ,
    \masters_02_aw_prot[0] }),
    .axi_spi_master_aw_qos({\masters_02_aw_qos[3] ,
    \masters_02_aw_qos[2] ,
    \masters_02_aw_qos[1] ,
    \masters_02_aw_qos[0] }),
    .axi_spi_master_aw_region({\masters_02_aw_region[3] ,
    \masters_02_aw_region[2] ,
    \masters_02_aw_region[1] ,
    \masters_02_aw_region[0] }),
    .axi_spi_master_aw_size({\masters_02_aw_size[2] ,
    \masters_02_aw_size[1] ,
    \masters_02_aw_size[0] }),
    .axi_spi_master_aw_user({_NC1087,
    _NC1088,
    _NC1089,
    _NC1090,
    _NC1091,
    _NC1092}),
    .axi_spi_master_b_id({_NC1093,
    _NC1094,
    _NC1095,
    _NC1096,
    _NC1097,
    _NC1098}),
    .axi_spi_master_b_resp({\masters_02_b_resp[1] ,
    \masters_02_b_resp[0] }),
    .axi_spi_master_b_user({_NC1099,
    _NC1100,
    _NC1101,
    _NC1102,
    _NC1103,
    _NC1104}),
    .axi_spi_master_r_data({_NC1105,
    _NC1106,
    _NC1107,
    _NC1108,
    _NC1109,
    _NC1110,
    _NC1111,
    _NC1112,
    _NC1113,
    _NC1114,
    _NC1115,
    _NC1116,
    _NC1117,
    _NC1118,
    _NC1119,
    _NC1120,
    _NC1121,
    _NC1122,
    _NC1123,
    _NC1124,
    _NC1125,
    _NC1126,
    _NC1127,
    _NC1128,
    _NC1129,
    _NC1130,
    _NC1131,
    _NC1132,
    _NC1133,
    _NC1134,
    _NC1135,
    _NC1136,
    _NC1137,
    _NC1138,
    _NC1139,
    _NC1140,
    _NC1141,
    _NC1142,
    _NC1143,
    _NC1144,
    _NC1145,
    _NC1146,
    _NC1147,
    _NC1148,
    _NC1149,
    _NC1150,
    _NC1151,
    _NC1152,
    _NC1153,
    _NC1154,
    _NC1155,
    _NC1156,
    _NC1157,
    _NC1158,
    _NC1159,
    _NC1160,
    _NC1161,
    _NC1162,
    _NC1163,
    _NC1164,
    _NC1165,
    _NC1166,
    _NC1167,
    _NC1168}),
    .axi_spi_master_r_id({_NC1169,
    _NC1170,
    _NC1171,
    _NC1172,
    _NC1173,
    _NC1174}),
    .axi_spi_master_r_resp({\masters_02_r_resp[1] ,
    \masters_02_r_resp[0] }),
    .axi_spi_master_r_user({_NC1175,
    _NC1176,
    _NC1177,
    _NC1178,
    _NC1179,
    _NC1180}),
    .axi_spi_master_w_data({_NC1181,
    _NC1182,
    _NC1183,
    _NC1184,
    _NC1185,
    _NC1186,
    _NC1187,
    _NC1188,
    _NC1189,
    _NC1190,
    _NC1191,
    _NC1192,
    _NC1193,
    _NC1194,
    _NC1195,
    _NC1196,
    _NC1197,
    _NC1198,
    _NC1199,
    _NC1200,
    _NC1201,
    _NC1202,
    _NC1203,
    _NC1204,
    _NC1205,
    _NC1206,
    _NC1207,
    _NC1208,
    _NC1209,
    _NC1210,
    _NC1211,
    _NC1212,
    _NC1213,
    _NC1214,
    _NC1215,
    _NC1216,
    _NC1217,
    _NC1218,
    _NC1219,
    _NC1220,
    _NC1221,
    _NC1222,
    _NC1223,
    _NC1224,
    _NC1225,
    _NC1226,
    _NC1227,
    _NC1228,
    _NC1229,
    _NC1230,
    _NC1231,
    _NC1232,
    _NC1233,
    _NC1234,
    _NC1235,
    _NC1236,
    _NC1237,
    _NC1238,
    _NC1239,
    _NC1240,
    _NC1241,
    _NC1242,
    _NC1243,
    _NC1244}),
    .axi_spi_master_w_strb({_NC1245,
    _NC1246,
    _NC1247,
    _NC1248,
    _NC1249,
    _NC1250,
    _NC1251,
    _NC1252}),
    .axi_spi_master_w_user({_NC1253,
    _NC1254,
    _NC1255,
    _NC1256,
    _NC1257,
    _NC1258}),
    .boot_addr_o({\boot_addr_int[31] ,
    \boot_addr_int[30] ,
    \boot_addr_int[29] ,
    \boot_addr_int[28] ,
    \boot_addr_int[27] ,
    \boot_addr_int[26] ,
    \boot_addr_int[25] ,
    \boot_addr_int[24] ,
    \boot_addr_int[23] ,
    \boot_addr_int[22] ,
    \boot_addr_int[21] ,
    \boot_addr_int[20] ,
    \boot_addr_int[19] ,
    \boot_addr_int[18] ,
    \boot_addr_int[17] ,
    \boot_addr_int[16] ,
    \boot_addr_int[15] ,
    \boot_addr_int[14] ,
    \boot_addr_int[13] ,
    \boot_addr_int[12] ,
    \boot_addr_int[11] ,
    \boot_addr_int[10] ,
    \boot_addr_int[9] ,
    \boot_addr_int[8] ,
    \boot_addr_int[7] ,
    \boot_addr_int[6] ,
    \boot_addr_int[5] ,
    \boot_addr_int[4] ,
    \boot_addr_int[3] ,
    \boot_addr_int[2] ,
    \boot_addr_int[1] ,
    \boot_addr_int[0] }),
    .debug_addr({\debug_addr[14] ,
    \debug_addr[13] ,
    \debug_addr[12] ,
    \debug_addr[11] ,
    \debug_addr[10] ,
    \debug_addr[9] ,
    \debug_addr[8] ,
    \debug_addr[7] ,
    \debug_addr[6] ,
    \debug_addr[5] ,
    \debug_addr[4] ,
    \debug_addr[3] ,
    \debug_addr[2] ,
    \debug_addr[1] ,
    \debug_addr[0] }),
    .debug_rdata({\debug_rdata[31] ,
    \debug_rdata[30] ,
    \debug_rdata[29] ,
    \debug_rdata[28] ,
    \debug_rdata[27] ,
    \debug_rdata[26] ,
    \debug_rdata[25] ,
    \debug_rdata[24] ,
    \debug_rdata[23] ,
    \debug_rdata[22] ,
    \debug_rdata[21] ,
    \debug_rdata[20] ,
    \debug_rdata[19] ,
    \debug_rdata[18] ,
    \debug_rdata[17] ,
    \debug_rdata[16] ,
    \debug_rdata[15] ,
    \debug_rdata[14] ,
    \debug_rdata[13] ,
    \debug_rdata[12] ,
    \debug_rdata[11] ,
    \debug_rdata[10] ,
    \debug_rdata[9] ,
    \debug_rdata[8] ,
    \debug_rdata[7] ,
    \debug_rdata[6] ,
    \debug_rdata[5] ,
    \debug_rdata[4] ,
    \debug_rdata[3] ,
    \debug_rdata[2] ,
    \debug_rdata[1] ,
    \debug_rdata[0] }),
    .debug_wdata({\debug_wdata[31] ,
    \debug_wdata[30] ,
    \debug_wdata[29] ,
    \debug_wdata[28] ,
    \debug_wdata[27] ,
    \debug_wdata[26] ,
    \debug_wdata[25] ,
    \debug_wdata[24] ,
    \debug_wdata[23] ,
    \debug_wdata[22] ,
    \debug_wdata[21] ,
    \debug_wdata[20] ,
    \debug_wdata[19] ,
    \debug_wdata[18] ,
    \debug_wdata[17] ,
    \debug_wdata[16] ,
    \debug_wdata[15] ,
    \debug_wdata[14] ,
    \debug_wdata[13] ,
    \debug_wdata[12] ,
    \debug_wdata[11] ,
    \debug_wdata[10] ,
    \debug_wdata[9] ,
    \debug_wdata[8] ,
    \debug_wdata[7] ,
    \debug_wdata[6] ,
    \debug_wdata[5] ,
    \debug_wdata[4] ,
    \debug_wdata[3] ,
    \debug_wdata[2] ,
    \debug_wdata[1] ,
    \debug_wdata[0] }),
    .fll1_add_o({\cfgad_fll_int[1] ,
    \cfgad_fll_int[0] }),
    .fll1_rdata_i({\cfgq_fll_int[31] ,
    \cfgq_fll_int[30] ,
    \cfgq_fll_int[29] ,
    \cfgq_fll_int[28] ,
    \cfgq_fll_int[27] ,
    \cfgq_fll_int[26] ,
    \cfgq_fll_int[25] ,
    \cfgq_fll_int[24] ,
    \cfgq_fll_int[23] ,
    \cfgq_fll_int[22] ,
    \cfgq_fll_int[21] ,
    \cfgq_fll_int[20] ,
    \cfgq_fll_int[19] ,
    \cfgq_fll_int[18] ,
    \cfgq_fll_int[17] ,
    \cfgq_fll_int[16] ,
    \cfgq_fll_int[15] ,
    \cfgq_fll_int[14] ,
    \cfgq_fll_int[13] ,
    \cfgq_fll_int[12] ,
    \cfgq_fll_int[11] ,
    \cfgq_fll_int[10] ,
    \cfgq_fll_int[9] ,
    \cfgq_fll_int[8] ,
    \cfgq_fll_int[7] ,
    \cfgq_fll_int[6] ,
    \cfgq_fll_int[5] ,
    \cfgq_fll_int[4] ,
    \cfgq_fll_int[3] ,
    \cfgq_fll_int[2] ,
    \cfgq_fll_int[1] ,
    \cfgq_fll_int[0] }),
    .fll1_wdata_o({\cfgd_fll_int[31] ,
    \cfgd_fll_int[30] ,
    \cfgd_fll_int[29] ,
    \cfgd_fll_int[28] ,
    \cfgd_fll_int[27] ,
    \cfgd_fll_int[26] ,
    \cfgd_fll_int[25] ,
    \cfgd_fll_int[24] ,
    \cfgd_fll_int[23] ,
    \cfgd_fll_int[22] ,
    \cfgd_fll_int[21] ,
    \cfgd_fll_int[20] ,
    \cfgd_fll_int[19] ,
    \cfgd_fll_int[18] ,
    \cfgd_fll_int[17] ,
    \cfgd_fll_int[16] ,
    \cfgd_fll_int[15] ,
    \cfgd_fll_int[14] ,
    \cfgd_fll_int[13] ,
    \cfgd_fll_int[12] ,
    \cfgd_fll_int[11] ,
    \cfgd_fll_int[10] ,
    \cfgd_fll_int[9] ,
    \cfgd_fll_int[8] ,
    \cfgd_fll_int[7] ,
    \cfgd_fll_int[6] ,
    \cfgd_fll_int[5] ,
    \cfgd_fll_int[4] ,
    \cfgd_fll_int[3] ,
    \cfgd_fll_int[2] ,
    \cfgd_fll_int[1] ,
    \cfgd_fll_int[0] }),
    .fll_add_i_pll({\cfgad_fll_int[1] ,
    \cfgad_fll_int[0] }),
    .fll_data_i_pll({\cfgd_fll_int[31] ,
    \cfgd_fll_int[30] ,
    \cfgd_fll_int[29] ,
    \cfgd_fll_int[28] ,
    \cfgd_fll_int[27] ,
    \cfgd_fll_int[26] ,
    \cfgd_fll_int[25] ,
    \cfgd_fll_int[24] ,
    \cfgd_fll_int[23] ,
    \cfgd_fll_int[22] ,
    \cfgd_fll_int[21] ,
    \cfgd_fll_int[20] ,
    \cfgd_fll_int[19] ,
    \cfgd_fll_int[18] ,
    \cfgd_fll_int[17] ,
    \cfgd_fll_int[16] ,
    \cfgd_fll_int[15] ,
    \cfgd_fll_int[14] ,
    \cfgd_fll_int[13] ,
    \cfgd_fll_int[12] ,
    \cfgd_fll_int[11] ,
    \cfgd_fll_int[10] ,
    \cfgd_fll_int[9] ,
    \cfgd_fll_int[8] ,
    \cfgd_fll_int[7] ,
    \cfgd_fll_int[6] ,
    \cfgd_fll_int[5] ,
    \cfgd_fll_int[4] ,
    \cfgd_fll_int[3] ,
    \cfgd_fll_int[2] ,
    \cfgd_fll_int[1] ,
    \cfgd_fll_int[0] }),
    .fll_r_data_o_pll({\cfgq_fll_int[31] ,
    \cfgq_fll_int[30] ,
    \cfgq_fll_int[29] ,
    \cfgq_fll_int[28] ,
    \cfgq_fll_int[27] ,
    \cfgq_fll_int[26] ,
    \cfgq_fll_int[25] ,
    \cfgq_fll_int[24] ,
    \cfgq_fll_int[23] ,
    \cfgq_fll_int[22] ,
    \cfgq_fll_int[21] ,
    \cfgq_fll_int[20] ,
    \cfgq_fll_int[19] ,
    \cfgq_fll_int[18] ,
    \cfgq_fll_int[17] ,
    \cfgq_fll_int[16] ,
    \cfgq_fll_int[15] ,
    \cfgq_fll_int[14] ,
    \cfgq_fll_int[13] ,
    \cfgq_fll_int[12] ,
    \cfgq_fll_int[11] ,
    \cfgq_fll_int[10] ,
    \cfgq_fll_int[9] ,
    \cfgq_fll_int[8] ,
    \cfgq_fll_int[7] ,
    \cfgq_fll_int[6] ,
    \cfgq_fll_int[5] ,
    \cfgq_fll_int[4] ,
    \cfgq_fll_int[3] ,
    \cfgq_fll_int[2] ,
    \cfgq_fll_int[1] ,
    \cfgq_fll_int[0] }),
    .gpio_dir({la_data_out[127],
    la_data_out[126],
    la_data_out[125],
    la_data_out[124],
    la_data_out[123],
    la_data_out[122],
    la_data_out[121],
    la_data_out[120],
    la_data_out[119],
    la_data_out[118],
    la_data_out[117],
    la_data_out[116],
    la_data_out[115],
    la_data_out[114],
    la_data_out[113],
    la_data_out[112],
    la_data_out[111],
    la_data_out[110],
    la_data_out[109],
    la_data_out[108],
    la_data_out[107],
    la_data_out[106],
    la_data_out[105],
    la_data_out[104],
    la_data_out[103],
    la_data_out[102],
    la_data_out[101],
    la_data_out[100],
    la_data_out[99],
    la_data_out[98],
    la_data_out[97],
    la_data_out[96]}),
    .gpio_in({la_data_in[38],
    la_data_in[37],
    la_data_in[36],
    la_data_in[35],
    la_data_in[34],
    la_data_in[33],
    la_data_in[32],
    la_data_in[31],
    la_data_in[30],
    la_data_in[29],
    la_data_in[28],
    la_data_in[27],
    la_data_in[26],
    la_data_in[25],
    la_data_in[24],
    la_data_in[23],
    la_data_in[22],
    la_data_in[21],
    la_data_in[20],
    la_data_in[19],
    la_data_in[18],
    la_data_in[17],
    la_data_in[16],
    la_data_in[15],
    la_data_in[14],
    la_data_in[13],
    la_data_in[12],
    la_data_in[11],
    la_data_in[10],
    la_data_in[9],
    la_data_in[8],
    la_data_in[7]}),
    .gpio_out({la_data_out[95],
    la_data_out[94],
    la_data_out[93],
    la_data_out[92],
    la_data_out[91],
    la_data_out[90],
    la_data_out[89],
    la_data_out[88],
    la_data_out[87],
    la_data_out[86],
    la_data_out[85],
    la_data_out[84],
    la_data_out[83],
    la_data_out[82],
    la_data_out[81],
    la_data_out[80],
    la_data_out[79],
    la_data_out[78],
    la_data_out[77],
    la_data_out[76],
    la_data_out[75],
    la_data_out[74],
    la_data_out[73],
    la_data_out[72],
    la_data_out[71],
    la_data_out[70],
    la_data_out[69],
    la_data_out[68],
    la_data_out[67],
    la_data_out[66],
    la_data_out[65],
    la_data_out[64]}),
    .gpio_padcfg({\gpio_padcfg[191] ,
    \gpio_padcfg[190] ,
    \gpio_padcfg[189] ,
    \gpio_padcfg[188] ,
    \gpio_padcfg[187] ,
    \gpio_padcfg[186] ,
    \gpio_padcfg[185] ,
    \gpio_padcfg[184] ,
    \gpio_padcfg[183] ,
    \gpio_padcfg[182] ,
    \gpio_padcfg[181] ,
    \gpio_padcfg[180] ,
    \gpio_padcfg[179] ,
    \gpio_padcfg[178] ,
    \gpio_padcfg[177] ,
    \gpio_padcfg[176] ,
    \gpio_padcfg[175] ,
    \gpio_padcfg[174] ,
    \gpio_padcfg[173] ,
    \gpio_padcfg[172] ,
    \gpio_padcfg[171] ,
    \gpio_padcfg[170] ,
    \gpio_padcfg[169] ,
    \gpio_padcfg[168] ,
    \gpio_padcfg[167] ,
    \gpio_padcfg[166] ,
    \gpio_padcfg[165] ,
    \gpio_padcfg[164] ,
    \gpio_padcfg[163] ,
    \gpio_padcfg[162] ,
    \gpio_padcfg[161] ,
    \gpio_padcfg[160] ,
    \gpio_padcfg[159] ,
    \gpio_padcfg[158] ,
    \gpio_padcfg[157] ,
    \gpio_padcfg[156] ,
    \gpio_padcfg[155] ,
    \gpio_padcfg[154] ,
    \gpio_padcfg[153] ,
    \gpio_padcfg[152] ,
    \gpio_padcfg[151] ,
    \gpio_padcfg[150] ,
    \gpio_padcfg[149] ,
    \gpio_padcfg[148] ,
    \gpio_padcfg[147] ,
    \gpio_padcfg[146] ,
    \gpio_padcfg[145] ,
    \gpio_padcfg[144] ,
    \gpio_padcfg[143] ,
    \gpio_padcfg[142] ,
    \gpio_padcfg[141] ,
    \gpio_padcfg[140] ,
    \gpio_padcfg[139] ,
    \gpio_padcfg[138] ,
    \gpio_padcfg[137] ,
    \gpio_padcfg[136] ,
    \gpio_padcfg[135] ,
    \gpio_padcfg[134] ,
    \gpio_padcfg[133] ,
    \gpio_padcfg[132] ,
    \gpio_padcfg[131] ,
    \gpio_padcfg[130] ,
    \gpio_padcfg[129] ,
    \gpio_padcfg[128] ,
    \gpio_padcfg[127] ,
    \gpio_padcfg[126] ,
    \gpio_padcfg[125] ,
    \gpio_padcfg[124] ,
    \gpio_padcfg[123] ,
    \gpio_padcfg[122] ,
    \gpio_padcfg[121] ,
    \gpio_padcfg[120] ,
    \gpio_padcfg[119] ,
    \gpio_padcfg[118] ,
    \gpio_padcfg[117] ,
    \gpio_padcfg[116] ,
    \gpio_padcfg[115] ,
    \gpio_padcfg[114] ,
    \gpio_padcfg[113] ,
    \gpio_padcfg[112] ,
    \gpio_padcfg[111] ,
    \gpio_padcfg[110] ,
    \gpio_padcfg[109] ,
    \gpio_padcfg[108] ,
    \gpio_padcfg[107] ,
    \gpio_padcfg[106] ,
    \gpio_padcfg[105] ,
    \gpio_padcfg[104] ,
    \gpio_padcfg[103] ,
    \gpio_padcfg[102] ,
    \gpio_padcfg[101] ,
    \gpio_padcfg[100] ,
    \gpio_padcfg[99] ,
    \gpio_padcfg[98] ,
    \gpio_padcfg[97] ,
    \gpio_padcfg[96] ,
    \gpio_padcfg[95] ,
    \gpio_padcfg[94] ,
    \gpio_padcfg[93] ,
    \gpio_padcfg[92] ,
    \gpio_padcfg[91] ,
    \gpio_padcfg[90] ,
    \gpio_padcfg[89] ,
    \gpio_padcfg[88] ,
    \gpio_padcfg[87] ,
    \gpio_padcfg[86] ,
    \gpio_padcfg[85] ,
    \gpio_padcfg[84] ,
    \gpio_padcfg[83] ,
    \gpio_padcfg[82] ,
    \gpio_padcfg[81] ,
    \gpio_padcfg[80] ,
    \gpio_padcfg[79] ,
    \gpio_padcfg[78] ,
    \gpio_padcfg[77] ,
    \gpio_padcfg[76] ,
    \gpio_padcfg[75] ,
    \gpio_padcfg[74] ,
    \gpio_padcfg[73] ,
    \gpio_padcfg[72] ,
    \gpio_padcfg[71] ,
    \gpio_padcfg[70] ,
    \gpio_padcfg[69] ,
    \gpio_padcfg[68] ,
    \gpio_padcfg[67] ,
    \gpio_padcfg[66] ,
    \gpio_padcfg[65] ,
    \gpio_padcfg[64] ,
    \gpio_padcfg[63] ,
    \gpio_padcfg[62] ,
    \gpio_padcfg[61] ,
    \gpio_padcfg[60] ,
    \gpio_padcfg[59] ,
    \gpio_padcfg[58] ,
    \gpio_padcfg[57] ,
    \gpio_padcfg[56] ,
    \gpio_padcfg[55] ,
    \gpio_padcfg[54] ,
    \gpio_padcfg[53] ,
    \gpio_padcfg[52] ,
    \gpio_padcfg[51] ,
    \gpio_padcfg[50] ,
    \gpio_padcfg[49] ,
    \gpio_padcfg[48] ,
    \gpio_padcfg[47] ,
    \gpio_padcfg[46] ,
    \gpio_padcfg[45] ,
    \gpio_padcfg[44] ,
    \gpio_padcfg[43] ,
    \gpio_padcfg[42] ,
    \gpio_padcfg[41] ,
    \gpio_padcfg[40] ,
    \gpio_padcfg[39] ,
    \gpio_padcfg[38] ,
    \gpio_padcfg[37] ,
    \gpio_padcfg[36] ,
    \gpio_padcfg[35] ,
    \gpio_padcfg[34] ,
    \gpio_padcfg[33] ,
    \gpio_padcfg[32] ,
    \gpio_padcfg[31] ,
    \gpio_padcfg[30] ,
    \gpio_padcfg[29] ,
    \gpio_padcfg[28] ,
    \gpio_padcfg[27] ,
    \gpio_padcfg[26] ,
    \gpio_padcfg[25] ,
    \gpio_padcfg[24] ,
    \gpio_padcfg[23] ,
    \gpio_padcfg[22] ,
    \gpio_padcfg[21] ,
    \gpio_padcfg[20] ,
    \gpio_padcfg[19] ,
    \gpio_padcfg[18] ,
    \gpio_padcfg[17] ,
    \gpio_padcfg[16] ,
    \gpio_padcfg[15] ,
    \gpio_padcfg[14] ,
    \gpio_padcfg[13] ,
    \gpio_padcfg[12] ,
    \gpio_padcfg[11] ,
    \gpio_padcfg[10] ,
    \gpio_padcfg[9] ,
    \gpio_padcfg[8] ,
    \gpio_padcfg[7] ,
    \gpio_padcfg[6] ,
    \gpio_padcfg[5] ,
    \gpio_padcfg[4] ,
    \gpio_padcfg[3] ,
    \gpio_padcfg[2] ,
    \gpio_padcfg[1] ,
    \gpio_padcfg[0] }),
    .io_oeb_pll({io_oeb[37],
    io_oeb[36],
    io_oeb[35],
    io_oeb[34],
    io_oeb[33],
    io_oeb[32],
    io_oeb[31],
    io_oeb[30],
    io_oeb[29],
    io_oeb[28],
    io_oeb[27],
    io_oeb[26],
    io_oeb[25],
    io_oeb[24],
    io_oeb[23],
    io_oeb[22],
    io_oeb[21],
    io_oeb[20],
    io_oeb[19],
    io_oeb[18],
    io_oeb[17],
    io_oeb[16],
    io_oeb[15],
    io_oeb[14],
    io_oeb[13],
    io_oeb[12],
    io_oeb[11],
    io_oeb[10],
    io_oeb[9],
    io_oeb[8],
    io_oeb[7],
    io_oeb[6],
    io_oeb[5],
    io_oeb[4],
    io_oeb[3],
    io_oeb[2],
    io_oeb[1],
    io_oeb[0]}),
    .io_out_pll({io_out[25],
    io_out[24],
    io_out[23],
    io_out[22],
    io_out[21],
    io_out[20],
    io_out[19],
    io_out[18],
    io_out[17],
    io_out[16],
    io_out[15],
    io_out[14],
    io_out[13],
    io_out[12],
    io_out[11],
    io_out[10],
    io_out[9],
    io_out[8],
    io_out[7],
    io_out[6],
    io_out[5],
    io_out[4],
    io_out[3],
    io_out[2],
    io_out[1],
    io_out[0]}),
    .irq_o({\irq_to_core_int[31] ,
    \irq_to_core_int[30] ,
    \irq_to_core_int[29] ,
    \irq_to_core_int[28] ,
    \irq_to_core_int[27] ,
    \irq_to_core_int[26] ,
    \irq_to_core_int[25] ,
    \irq_to_core_int[24] ,
    \irq_to_core_int[23] ,
    \irq_to_core_int[22] ,
    \irq_to_core_int[21] ,
    \irq_to_core_int[20] ,
    \irq_to_core_int[19] ,
    \irq_to_core_int[18] ,
    \irq_to_core_int[17] ,
    \irq_to_core_int[16] ,
    \irq_to_core_int[15] ,
    \irq_to_core_int[14] ,
    \irq_to_core_int[13] ,
    \irq_to_core_int[12] ,
    \irq_to_core_int[11] ,
    \irq_to_core_int[10] ,
    \irq_to_core_int[9] ,
    \irq_to_core_int[8] ,
    \irq_to_core_int[7] ,
    \irq_to_core_int[6] ,
    \irq_to_core_int[5] ,
    \irq_to_core_int[4] ,
    \irq_to_core_int[3] ,
    \irq_to_core_int[2] ,
    \irq_to_core_int[1] ,
    \irq_to_core_int[0] }),
    .la_data_out_pll({la_data_out[63],
    la_data_out[62],
    la_data_out[61],
    la_data_out[60],
    la_data_out[59],
    la_data_out[58],
    la_data_out[57],
    la_data_out[56],
    la_data_out[55],
    la_data_out[54],
    la_data_out[53],
    la_data_out[52],
    la_data_out[51],
    la_data_out[50],
    la_data_out[49],
    la_data_out[48],
    la_data_out[47],
    la_data_out[46],
    la_data_out[45],
    la_data_out[44],
    la_data_out[43],
    la_data_out[42],
    la_data_out[41],
    la_data_out[40],
    la_data_out[39],
    la_data_out[38],
    la_data_out[37],
    la_data_out[36],
    la_data_out[35],
    la_data_out[34],
    la_data_out[33],
    la_data_out[32],
    la_data_out[31],
    la_data_out[30],
    la_data_out[29],
    la_data_out[28],
    la_data_out[27],
    la_data_out[26],
    la_data_out[25],
    la_data_out[24],
    la_data_out[23],
    la_data_out[22],
    la_data_out[21],
    la_data_out[20],
    la_data_out[19],
    la_data_out[18],
    la_data_out[17],
    la_data_out[16],
    la_data_out[15],
    la_data_out[14],
    la_data_out[13],
    la_data_out[12],
    la_data_out[11],
    la_data_out[10],
    la_data_out[9],
    la_data_out[8],
    la_data_out[7],
    la_data_out[6],
    la_data_out[5],
    la_data_out[4],
    la_data_out[3],
    la_data_out[2],
    la_data_out[1],
    la_data_out[0]}),
    .slave_ar_addr({\slaves_02_ar_addr[31] ,
    \slaves_02_ar_addr[30] ,
    \slaves_02_ar_addr[29] ,
    \slaves_02_ar_addr[28] ,
    \slaves_02_ar_addr[27] ,
    \slaves_02_ar_addr[26] ,
    \slaves_02_ar_addr[25] ,
    \slaves_02_ar_addr[24] ,
    \slaves_02_ar_addr[23] ,
    \slaves_02_ar_addr[22] ,
    \slaves_02_ar_addr[21] ,
    \slaves_02_ar_addr[20] ,
    \slaves_02_ar_addr[19] ,
    \slaves_02_ar_addr[18] ,
    \slaves_02_ar_addr[17] ,
    \slaves_02_ar_addr[16] ,
    \slaves_02_ar_addr[15] ,
    \slaves_02_ar_addr[14] ,
    \slaves_02_ar_addr[13] ,
    \slaves_02_ar_addr[12] ,
    \slaves_02_ar_addr[11] ,
    \slaves_02_ar_addr[10] ,
    \slaves_02_ar_addr[9] ,
    \slaves_02_ar_addr[8] ,
    \slaves_02_ar_addr[7] ,
    \slaves_02_ar_addr[6] ,
    \slaves_02_ar_addr[5] ,
    \slaves_02_ar_addr[4] ,
    \slaves_02_ar_addr[3] ,
    \slaves_02_ar_addr[2] ,
    \slaves_02_ar_addr[1] ,
    \slaves_02_ar_addr[0] }),
    .slave_ar_burst({\slaves_02_ar_burst[1] ,
    \slaves_02_ar_burst[0] }),
    .slave_ar_cache({\slaves_02_ar_cache[3] ,
    \slaves_02_ar_cache[2] ,
    \slaves_02_ar_cache[1] ,
    \slaves_02_ar_cache[0] }),
    .slave_ar_id({_NC1259,
    _NC1260,
    _NC1261,
    _NC1262,
    _NC1263,
    _NC1264}),
    .slave_ar_len({\slaves_02_ar_len[7] ,
    \slaves_02_ar_len[6] ,
    \slaves_02_ar_len[5] ,
    \slaves_02_ar_len[4] ,
    \slaves_02_ar_len[3] ,
    \slaves_02_ar_len[2] ,
    \slaves_02_ar_len[1] ,
    \slaves_02_ar_len[0] }),
    .slave_ar_prot({\slaves_02_ar_prot[2] ,
    \slaves_02_ar_prot[1] ,
    \slaves_02_ar_prot[0] }),
    .slave_ar_qos({\slaves_02_ar_qos[3] ,
    \slaves_02_ar_qos[2] ,
    \slaves_02_ar_qos[1] ,
    \slaves_02_ar_qos[0] }),
    .slave_ar_region({\slaves_02_ar_region[3] ,
    \slaves_02_ar_region[2] ,
    \slaves_02_ar_region[1] ,
    \slaves_02_ar_region[0] }),
    .slave_ar_size({\slaves_02_ar_size[2] ,
    \slaves_02_ar_size[1] ,
    \slaves_02_ar_size[0] }),
    .slave_ar_user({_NC1265,
    _NC1266,
    _NC1267,
    _NC1268,
    _NC1269,
    _NC1270}),
    .slave_aw_addr({\slaves_02_aw_addr[31] ,
    \slaves_02_aw_addr[30] ,
    \slaves_02_aw_addr[29] ,
    \slaves_02_aw_addr[28] ,
    \slaves_02_aw_addr[27] ,
    \slaves_02_aw_addr[26] ,
    \slaves_02_aw_addr[25] ,
    \slaves_02_aw_addr[24] ,
    \slaves_02_aw_addr[23] ,
    \slaves_02_aw_addr[22] ,
    \slaves_02_aw_addr[21] ,
    \slaves_02_aw_addr[20] ,
    \slaves_02_aw_addr[19] ,
    \slaves_02_aw_addr[18] ,
    \slaves_02_aw_addr[17] ,
    \slaves_02_aw_addr[16] ,
    \slaves_02_aw_addr[15] ,
    \slaves_02_aw_addr[14] ,
    \slaves_02_aw_addr[13] ,
    \slaves_02_aw_addr[12] ,
    \slaves_02_aw_addr[11] ,
    \slaves_02_aw_addr[10] ,
    \slaves_02_aw_addr[9] ,
    \slaves_02_aw_addr[8] ,
    \slaves_02_aw_addr[7] ,
    \slaves_02_aw_addr[6] ,
    \slaves_02_aw_addr[5] ,
    \slaves_02_aw_addr[4] ,
    \slaves_02_aw_addr[3] ,
    \slaves_02_aw_addr[2] ,
    \slaves_02_aw_addr[1] ,
    \slaves_02_aw_addr[0] }),
    .slave_aw_burst({\slaves_02_aw_burst[1] ,
    \slaves_02_aw_burst[0] }),
    .slave_aw_cache({\slaves_02_aw_cache[3] ,
    \slaves_02_aw_cache[2] ,
    \slaves_02_aw_cache[1] ,
    \slaves_02_aw_cache[0] }),
    .slave_aw_id({_NC1271,
    _NC1272,
    _NC1273,
    _NC1274,
    _NC1275,
    _NC1276}),
    .slave_aw_len({\slaves_02_aw_len[7] ,
    \slaves_02_aw_len[6] ,
    \slaves_02_aw_len[5] ,
    \slaves_02_aw_len[4] ,
    \slaves_02_aw_len[3] ,
    \slaves_02_aw_len[2] ,
    \slaves_02_aw_len[1] ,
    \slaves_02_aw_len[0] }),
    .slave_aw_prot({\slaves_02_aw_prot[2] ,
    \slaves_02_aw_prot[1] ,
    \slaves_02_aw_prot[0] }),
    .slave_aw_qos({\slaves_02_aw_qos[3] ,
    \slaves_02_aw_qos[2] ,
    \slaves_02_aw_qos[1] ,
    \slaves_02_aw_qos[0] }),
    .slave_aw_region({\slaves_02_aw_region[3] ,
    \slaves_02_aw_region[2] ,
    \slaves_02_aw_region[1] ,
    \slaves_02_aw_region[0] }),
    .slave_aw_size({\slaves_02_aw_size[2] ,
    \slaves_02_aw_size[1] ,
    \slaves_02_aw_size[0] }),
    .slave_aw_user({_NC1277,
    _NC1278,
    _NC1279,
    _NC1280,
    _NC1281,
    _NC1282}),
    .slave_b_id({_NC1283,
    _NC1284,
    _NC1285,
    _NC1286,
    _NC1287,
    _NC1288}),
    .slave_b_resp({\slaves_02_b_resp[1] ,
    \slaves_02_b_resp[0] }),
    .slave_b_user({_NC1289,
    _NC1290,
    _NC1291,
    _NC1292,
    _NC1293,
    _NC1294}),
    .slave_r_data({_NC1295,
    _NC1296,
    _NC1297,
    _NC1298,
    _NC1299,
    _NC1300,
    _NC1301,
    _NC1302,
    _NC1303,
    _NC1304,
    _NC1305,
    _NC1306,
    _NC1307,
    _NC1308,
    _NC1309,
    _NC1310,
    _NC1311,
    _NC1312,
    _NC1313,
    _NC1314,
    _NC1315,
    _NC1316,
    _NC1317,
    _NC1318,
    _NC1319,
    _NC1320,
    _NC1321,
    _NC1322,
    _NC1323,
    _NC1324,
    _NC1325,
    _NC1326,
    _NC1327,
    _NC1328,
    _NC1329,
    _NC1330,
    _NC1331,
    _NC1332,
    _NC1333,
    _NC1334,
    _NC1335,
    _NC1336,
    _NC1337,
    _NC1338,
    _NC1339,
    _NC1340,
    _NC1341,
    _NC1342,
    _NC1343,
    _NC1344,
    _NC1345,
    _NC1346,
    _NC1347,
    _NC1348,
    _NC1349,
    _NC1350,
    _NC1351,
    _NC1352,
    _NC1353,
    _NC1354,
    _NC1355,
    _NC1356,
    _NC1357,
    _NC1358}),
    .slave_r_id({_NC1359,
    _NC1360,
    _NC1361,
    _NC1362,
    _NC1363,
    _NC1364}),
    .slave_r_resp({\slaves_02_r_resp[1] ,
    \slaves_02_r_resp[0] }),
    .slave_r_user({_NC1365,
    _NC1366,
    _NC1367,
    _NC1368,
    _NC1369,
    _NC1370}),
    .slave_w_data({_NC1371,
    _NC1372,
    _NC1373,
    _NC1374,
    _NC1375,
    _NC1376,
    _NC1377,
    _NC1378,
    _NC1379,
    _NC1380,
    _NC1381,
    _NC1382,
    _NC1383,
    _NC1384,
    _NC1385,
    _NC1386,
    _NC1387,
    _NC1388,
    _NC1389,
    _NC1390,
    _NC1391,
    _NC1392,
    _NC1393,
    _NC1394,
    _NC1395,
    _NC1396,
    _NC1397,
    _NC1398,
    _NC1399,
    _NC1400,
    _NC1401,
    _NC1402,
    _NC1403,
    _NC1404,
    _NC1405,
    _NC1406,
    _NC1407,
    _NC1408,
    _NC1409,
    _NC1410,
    _NC1411,
    _NC1412,
    _NC1413,
    _NC1414,
    _NC1415,
    _NC1416,
    _NC1417,
    _NC1418,
    _NC1419,
    _NC1420,
    _NC1421,
    _NC1422,
    _NC1423,
    _NC1424,
    _NC1425,
    _NC1426,
    _NC1427,
    _NC1428,
    _NC1429,
    _NC1430,
    _NC1431,
    _NC1432,
    _NC1433,
    _NC1434}),
    .slave_w_strb({_NC1435,
    _NC1436,
    _NC1437,
    _NC1438,
    _NC1439,
    _NC1440,
    _NC1441,
    _NC1442}),
    .slave_w_user({_NC1443,
    _NC1444,
    _NC1445,
    _NC1446,
    _NC1447,
    _NC1448}),
    .spi_master_mode({io_out[31],
    io_out[30]}),
    .spi_mode_o({io_out[37],
    io_out[36]}),
    .user_irq_pll({user_irq[2],
    user_irq[1],
    user_irq[0]}),
    .wbs_dat_o_pll({wbs_dat_o[31],
    wbs_dat_o[30],
    wbs_dat_o[29],
    wbs_dat_o[28],
    wbs_dat_o[27],
    wbs_dat_o[26],
    wbs_dat_o[25],
    wbs_dat_o[24],
    wbs_dat_o[23],
    wbs_dat_o[22],
    wbs_dat_o[21],
    wbs_dat_o[20],
    wbs_dat_o[19],
    wbs_dat_o[18],
    wbs_dat_o[17],
    wbs_dat_o[16],
    wbs_dat_o[15],
    wbs_dat_o[14],
    wbs_dat_o[13],
    wbs_dat_o[12],
    wbs_dat_o[11],
    wbs_dat_o[10],
    wbs_dat_o[9],
    wbs_dat_o[8],
    wbs_dat_o[7],
    wbs_dat_o[6],
    wbs_dat_o[5],
    wbs_dat_o[4],
    wbs_dat_o[3],
    wbs_dat_o[2],
    wbs_dat_o[1],
    wbs_dat_o[0]}));
endmodule
