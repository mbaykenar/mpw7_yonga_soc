magic
tech sky130B
magscale 12 1
timestamp 1598773327
<< metal5 >>
rect 20 100 90 105
rect 15 95 95 100
rect 10 90 100 95
rect 5 85 30 90
rect 80 85 105 90
rect 0 80 25 85
rect 85 80 105 85
rect 0 75 20 80
rect 0 0 15 75
rect 40 70 65 75
rect 35 65 70 70
rect 30 55 75 65
rect 30 20 45 55
rect 60 20 75 55
rect 90 20 105 80
rect 30 10 105 20
rect 35 5 100 10
rect 40 0 60 5
rect 75 0 95 5
rect 0 -5 20 0
rect 0 -10 25 -5
rect 5 -15 30 -10
rect 10 -20 90 -15
rect 15 -25 90 -20
rect 20 -30 90 -25
<< properties >>
string FIXED_BBOX 0 -30 120 105
<< end >>
