* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

* SKY130 Spice File.
.param sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre = 0.0
.param sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre = 0.0
.param sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre = 0.0
.param sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre = 0.0
* statistics {
*   process {
*   }
*   mismatch {
*     vary sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre dist=gauss std = 1.0
*     vary sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre dist=gauss std = 1.0
*     vary sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre dist=gauss std = 1.0
*     vary sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre dist=gauss std = 1.0
*   }
* }
.subckt  sky130_fd_pr__pfet_01v8_lvt d g s b
+ 
.param  l = 1 w = 1 nf = 1.0 ad = 0 as = 0 pd = 0 ps = 0 nrd = 0 nrs = 0 sa = 0 sb = 0 sd = 0 mult = 1
msky130_fd_pr__pfet_01v8_lvt d g s b sky130_fd_pr__pfet_01v8_lvt__model l = {l} w = {w} nf = {nf} ad = {ad} as = {as} pd = {pd} ps = {ps} nrd = {nrd} nrs = {nrs} sa = {sa} sb = {sb} sd = {sd}
.model sky130_fd_pr__pfet_01v8_lvt__model.0 pmos
* DC IV MOS Parameters
+ lmin = 2.0e-05 lmax = 1.0e-04 wmin = 7e-06 wmax = 1.0e-4
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 2.8e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 7.476e-9
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -7.916e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25000000.0
+ tnoib = 0.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.23e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-0.450452+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.64774
+ k2 = -0.0458948
+ k3 = 3.39
+ dvt0 = 2.4422
+ dvt1 = 0.16136
+ dvt2 = 0.026237
+ dvt0w = 0.5
+ dvt1w = 1928100.0
+ dvt2w = -0.032
+ w0 = 1.0e-8
+ k3b = 1.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 123760.0
+ ua = -3.0054e-9
+ ub = 3.0419e-18
+ uc = 4.9353e-11
+ rdsw = 484.7
+ prwb = 0.1
+ prwg = 0.052
+ wr = 1.0
+ u0 = 0.0025272667
+ a0 = 1.78166
+ keta = -0.01258
+ a1 = 0.0
+ a2 = 0.46703705
+ ags = 0.390807
+ b0 = 0.0
+ b1 = 2.1073e-24
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.1819+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))}
+ nfactor = {3.9789+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -6.393105e-11
+ cdsc = 2.8125e-7
+ cdscb = 1.0e-4
+ cdscd = 1.0e-10
+ eta0 = 0.2
+ etab = -0.00025
+ dsub = 1.0
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.030097
+ pdiblc1 = 0.0
+ pdiblc2 = 0.0018466
+ pdiblcb = -0.025
+ drout = 0.43496
+ pscbe1 = 800000000.0
+ pscbe2 = 8.6797e-9
+ pvag = 0.0
+ delta = 0.01363
+ alpha0 = 5.0449517e-13
+ alpha1 = -4.0583656e-18
+ beta0 = 6.2016506
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -1.07085
+ kt2 = -0.055045
+ at = 285600.0
+ ute = -0.22271
+ ua1 = 6.8217e-10
+ ub1 = -1.4864e-19
+ uc1 = -9.961e-12
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+41
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 1.4472e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 2.0e-11
+ cgso = 2.0e-11
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 0.0
+ cgdl = 0.0
+ cf = 0.0
+ clc = 7.0e-8
+ cle = 0.492
+ dlc = -1.2e-8
+ dwc = 0.0
+ vfbcv = -1.0
+ acde = 0.44
+ moin = 8.7
+ noff = 2.6123
+ voffcv = 0.112
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007653568198
+ mjs = 0.3362
+ pbs = 0.6587
+ cjsws = 9.1602368e-11
+ mjsws = 0.2659
+ pbsws = 0.7418
+ cjswgs = 2.39155046e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.1 pmos
* DC IV MOS Parameters
+ lmin = 8e-06 lmax = 2.0e-05 wmin = 7e-06 wmax = 1.0e-4
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 2.8e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 7.476e-9
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -7.916e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25000000.0
+ tnoib = 0.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.23e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-0.450452+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.64774
+ k2 = -0.0458948
+ k3 = 3.39
+ dvt0 = 2.4422
+ dvt1 = 0.16136
+ dvt2 = 0.026237
+ dvt0w = 0.5
+ dvt1w = 1928100.0
+ dvt2w = -0.032
+ w0 = 1.0e-8
+ k3b = 1.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 123760.0
+ ua = -3.0054e-9
+ ub = 3.0419e-18
+ uc = 4.9353e-11
+ rdsw = 484.7
+ prwb = 0.1
+ prwg = 0.052
+ wr = 1.0
+ u0 = 0.0025272667
+ a0 = 1.78166
+ keta = -0.01258
+ a1 = 0.0
+ a2 = 0.46703705
+ ags = 0.390807
+ b0 = 0.0
+ b1 = 2.1073e-24
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.1819+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))}
+ nfactor = {3.9789+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -6.393105e-11
+ cdsc = 2.8125e-7
+ cdscb = 1.0e-4
+ cdscd = 1.0e-10
+ eta0 = 0.2
+ etab = -0.00025
+ dsub = 1.0
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.030097
+ pdiblc1 = 0.0
+ pdiblc2 = 0.0018466
+ pdiblcb = -0.025
+ drout = 0.43496
+ pscbe1 = 800000000.0
+ pscbe2 = 8.6797e-9
+ pvag = 0.0
+ delta = 0.01363
+ alpha0 = 5.0449517e-13
+ alpha1 = -4.0583656e-18
+ beta0 = 6.2016506
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -1.07085
+ kt2 = -0.055045
+ at = 285600.0
+ ute = -0.22271
+ ua1 = 6.8217e-10
+ ub1 = -1.4864e-19
+ uc1 = -9.961e-12
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+41
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 1.4472e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 2.0e-11
+ cgso = 2.0e-11
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 0.0
+ cgdl = 0.0
+ cf = 0.0
+ clc = 7.0e-8
+ cle = 0.492
+ dlc = -1.2e-8
+ dwc = 0.0
+ vfbcv = -1.0
+ acde = 0.44
+ moin = 8.7
+ noff = 2.6123
+ voffcv = 0.112
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007653568198
+ mjs = 0.3362
+ pbs = 0.6587
+ cjsws = 9.1602368e-11
+ mjsws = 0.2659
+ pbsws = 0.7418
+ cjswgs = 2.39155046e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.2 pmos
* DC IV MOS Parameters
+ lmin = 4e-06 lmax = 8e-06 wmin = 7e-06 wmax = 1.0e-4
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 2.8e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 7.476e-9
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -7.916e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25000000.0
+ tnoib = 0.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.23e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-4.586515046e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 6.555011957e-8
+ k1 = 0.64774
+ k2 = -4.616172578e-02 lk2 = 2.133911456e-9
+ k3 = 3.39
+ dvt0 = 2.4422
+ dvt1 = 0.16136
+ dvt2 = 0.026237
+ dvt0w = 0.5
+ dvt1w = 1928100.0
+ dvt2w = -0.032
+ w0 = 1.0e-8
+ k3b = 1.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 123760.0
+ ua = -3.064217540e-09 lua = 4.702109418e-16
+ ub = 3.130975120e-18 lub = -7.121021393e-25
+ uc = 3.779220780e-11 luc = 9.242159716e-17
+ rdsw = 484.7
+ prwb = 0.1
+ prwg = 0.052
+ wr = 1.0
+ u0 = 2.442647034e-03 lu0 = 6.764834609e-10
+ a0 = 1.880980756e+00 la0 = -7.940098518e-7
+ keta = -0.01258
+ a1 = 0.0
+ a2 = 0.46703705
+ ags = 3.751948876e-01 lags = 1.248094714e-7
+ b0 = 0.0
+ b1 = 2.1073e-24
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.1819+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))}
+ nfactor = {4.450349046e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -3.768952253e-06 wnfactor = -6.776263578e-21
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -6.393105e-11
+ cdsc = 2.8125e-7
+ cdscb = 1.0e-4
+ cdscd = 1.0e-10
+ eta0 = 0.2
+ etab = -0.00025
+ dsub = 1.0
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.030097
+ pdiblc1 = 0.0
+ pdiblc2 = 7.488388000e-05 lpdiblc2 = 1.416380735e-8
+ pdiblcb = -0.025
+ drout = 0.43496
+ pscbe1 = 800000000.0
+ pscbe2 = 8.6797e-9
+ pvag = 0.0
+ delta = 5.859893400e-03 ldelta = 6.211734020e-8
+ alpha0 = 5.0449517e-13
+ alpha1 = -4.0583656e-18
+ beta0 = 6.2016506
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -1.134350974e+00 lkt1 = 5.076521865e-7
+ kt2 = -0.055045
+ at = 2.991709740e+05 lat = -1.084917945e-1
+ ute = -3.123143780e-01 lute = 7.163332395e-7
+ ua1 = 6.682694880e-10 lua1 = 1.111262531e-16
+ ub1 = -1.753625360e-19 lub1 = 2.136306418e-25
+ uc1 = -9.961e-12
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+41
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 1.4472e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 2.0e-11
+ cgso = 2.0e-11
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 0.0
+ cgdl = 0.0
+ cf = 0.0
+ clc = 7.0e-8
+ cle = 0.492
+ dlc = -1.2e-8
+ dwc = 0.0
+ vfbcv = -1.0
+ acde = 0.44
+ moin = 8.7
+ noff = 2.6123
+ voffcv = 0.112
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007653568198
+ mjs = 0.3362
+ pbs = 0.6587
+ cjsws = 9.1602368e-11
+ mjsws = 0.2659
+ pbsws = 0.7418
+ cjswgs = 2.39155046e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.3 pmos
* DC IV MOS Parameters
+ lmin = 2e-06 lmax = 4e-06 wmin = 7e-06 wmax = 1.0e-4
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 2.8e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 7.476e-9
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -7.916e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25000000.0
+ tnoib = 0.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.23e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-4.217136380e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -8.199449477e-8
+ k1 = 0.64774
+ k2 = -3.880974332e-02 lk2 = -2.723284728e-8
+ k3 = 3.39
+ dvt0 = 2.4422
+ dvt1 = 0.16136
+ dvt2 = 0.026237
+ dvt0w = 0.5
+ dvt1w = 1928100.0
+ dvt2w = -0.032
+ w0 = 1.0e-8
+ k3b = 1.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 1.566795664e+05 lvsat = -1.314939160e-1
+ ua = -3.113132120e-09 lua = 6.655953401e-16
+ ub = 3.175873360e-18 lub = -8.914436692e-25
+ uc = 6.136577640e-11 luc = -1.740665252e-18
+ rdsw = 484.7
+ prwb = 0.1
+ prwg = 0.052
+ wr = 1.0
+ u0 = 2.318823015e-03 lu0 = 1.171086123e-9
+ a0 = 2.278057913e+00 la0 = -2.380094848e-6
+ keta = -0.01258
+ a1 = 0.0
+ a2 = 0.46703705
+ ags = 4.214498572e-01 lags = -5.995137920e-8
+ b0 = 0.0
+ b1 = 2.1073e-24
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.1819+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))}
+ nfactor = {3.358197228e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 5.935389685e-7
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -6.393105e-11
+ cdsc = 2.8125e-7
+ cdscb = 1.0e-4
+ cdscd = 1.0e-10
+ eta0 = 0.2
+ etab = -0.00025
+ dsub = 1.0
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.030097
+ pdiblc1 = 0.0
+ pdiblc2 = 2.638259200e-04 lpdiblc2 = 1.340909727e-8
+ pdiblcb = -0.025
+ drout = 0.43496
+ pscbe1 = 800000000.0
+ pscbe2 = 8.6797e-9
+ pvag = 0.0
+ delta = 1.967986080e-02 ldelta = 6.914862420e-9
+ alpha0 = 5.0449517e-13
+ alpha1 = -4.0583656e-18
+ beta0 = 6.2016506
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -1.049800552e+00 lkt1 = 1.699239809e-7
+ kt2 = -0.055045
+ at = 3.780323040e+05 lat = -4.234954911e-1
+ ute = -0.13298
+ ua1 = 6.9609e-10
+ ub1 = -1.571260340e-19 lub1 = 1.407867582e-25
+ uc1 = -9.961e-12
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+41
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 1.4472e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 2.0e-11
+ cgso = 2.0e-11
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 0.0
+ cgdl = 0.0
+ cf = 0.0
+ clc = 7.0e-8
+ cle = 0.492
+ dlc = -1.2e-8
+ dwc = 0.0
+ vfbcv = -1.0
+ acde = 0.44
+ moin = 8.7
+ noff = 2.6123
+ voffcv = 0.112
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007653568198
+ mjs = 0.3362
+ pbs = 0.6587
+ cjsws = 9.1602368e-11
+ mjsws = 0.2659
+ pbsws = 0.7418
+ cjswgs = 2.39155046e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.4 pmos
* DC IV MOS Parameters
+ lmin = 1.5e-06 lmax = 2e-06 wmin = 7e-06 wmax = 1.0e-4
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 2.8e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 7.476e-9
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -7.916e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25000000.0
+ tnoib = 0.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.23e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-4.682476832e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 1.081300497e-8
+ k1 = 0.64774
+ k2 = -4.457785344e-02 lk2 = -1.572892846e-8
+ k3 = 3.39
+ dvt0 = 2.4422
+ dvt1 = 0.16136
+ dvt2 = 0.026237
+ dvt0w = 0.5
+ dvt1w = 1928100.0
+ dvt2w = -0.032
+ w0 = 1.0e-8
+ k3b = 1.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 90748.0
+ ua = -2.234840640e-09 lua = -1.086069188e-15
+ ub = 1.831961120e-18 lub = 1.788854902e-24
+ uc = 2.748768160e-11 luc = 6.582580702e-17
+ rdsw = 484.7
+ prwb = 0.1
+ prwg = 0.052
+ wr = 1.0
+ u0 = 3.149729505e-03 lu0 = -4.860737818e-10
+ a0 = 1.084274478e+00 la0 = 7.868338790e-10
+ keta = -0.01258
+ a1 = 0.0
+ a2 = 0.46703705
+ ags = 1.599373280e-01 lags = 4.616092090e-7
+ b0 = 0.0
+ b1 = 2.1073e-24
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.1819+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))}
+ nfactor = {5.160541248e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -3.001055945e-6
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -6.393105e-11
+ cdsc = 2.8125e-7
+ cdscb = 1.0e-4
+ cdscd = 1.0e-10
+ eta0 = 0.2
+ etab = -0.00025
+ dsub = 1.0
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.030097
+ pdiblc1 = 0.0
+ pdiblc2 = -3.278730240e-03 lpdiblc2 = 2.047437127e-8
+ pdiblcb = -0.025
+ drout = 0.43496
+ pscbe1 = 800000000.0
+ pscbe2 = 8.6797e-9
+ pvag = 0.0
+ delta = 1.696915040e-02 ldelta = 1.232110324e-8
+ alpha0 = 5.0449517e-13
+ alpha1 = -4.0583656e-18
+ beta0 = 6.2016506
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -9.697706240e-01 lkt1 = 1.031229251e-8
+ kt2 = -0.055045
+ at = 2.058295840e+05 lat = -8.005438633e-2
+ ute = -0.13298
+ ua1 = 8.001002400e-10 lua1 = -2.074380227e-16
+ ub1 = -3.124733360e-19 lub1 = 4.506114173e-25
+ uc1 = -9.961e-12
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+41
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 1.4472e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 2.0e-11
+ cgso = 2.0e-11
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 0.0
+ cgdl = 0.0
+ cf = 0.0
+ clc = 7.0e-8
+ cle = 0.492
+ dlc = -1.2e-8
+ dwc = 0.0
+ vfbcv = -1.0
+ acde = 0.44
+ moin = 8.7
+ noff = 2.6123
+ voffcv = 0.112
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007653568198
+ mjs = 0.3362
+ pbs = 0.6587
+ cjsws = 9.1602368e-11
+ mjsws = 0.2659
+ pbsws = 0.7418
+ cjswgs = 2.39155046e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.5 pmos
* DC IV MOS Parameters
+ lmin = 1e-06 lmax = 1.5e-06 wmin = 7e-06 wmax = 1.0e-4
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 2.8e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 7.476e-9
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -7.916e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25000000.0
+ tnoib = 0.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.23e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-4.471281872e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -2.074796985e-8
+ k1 = 0.64774
+ k2 = -4.888670784e-02 lk2 = -9.289776444e-9
+ k3 = 3.39
+ dvt0 = 2.4422
+ dvt1 = 0.16136
+ dvt2 = 0.026237
+ dvt0w = 0.5
+ dvt1w = 1928100.0
+ dvt2w = -0.032
+ w0 = 1.0e-8
+ k3b = 1.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 9.002606560e+04 lvsat = 1.078858767e-3
+ ua = -3.153121440e-09 lua = 2.862096399e-16
+ ub = 3.140969440e-18 lub = -1.673271311e-25
+ uc = 6.937218560e-11 luc = 3.233604239e-18
+ rdsw = 484.7
+ prwb = 0.1
+ prwg = 0.052
+ wr = 1.0
+ u0 = 2.023902403e-03 lu0 = 1.196362239e-9
+ a0 = 9.850964896e-01 la0 = 1.489984203e-7
+ keta = -0.01258
+ a1 = 0.0
+ a2 = 0.46703705
+ ags = 3.280548800e-02 lags = 6.515950307e-7
+ b0 = 0.0
+ b1 = 2.1073e-24
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-1.529629600e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = -4.324351258e-8
+ nfactor = {4.406944648e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -1.874881186e-6
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -6.393105e-11
+ cdsc = 2.8125e-7
+ cdscb = 1.0e-4
+ cdscd = 1.0e-10
+ eta0 = 0.2
+ etab = -0.00025
+ dsub = 1.0
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.030097
+ pdiblc1 = 0.0
+ pdiblc2 = 5.973280000e-04 lpdiblc2 = 1.468198984e-8
+ pdiblcb = -0.025
+ drout = 0.43496
+ pscbe1 = 800000000.0
+ pscbe2 = 8.6797e-9
+ pvag = 0.0
+ delta = 1.023634720e-02 ldelta = 2.238260434e-8
+ alpha0 = 5.0449517e-13
+ alpha1 = -4.0583656e-18
+ beta0 = 6.2016506
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -1.093733040e+00 lkt1 = 1.955617270e-7
+ kt2 = -9.336122080e-02 lkt2 = 5.725976036e-8
+ at = 2.043466720e+05 lat = -7.783832264e-2
+ ute = 5.615488000e-02 lute = -2.826431647e-7
+ ua1 = 6.6129e-10
+ ub1 = -1.050445280e-20 lub1 = -6.508817357e-28
+ uc1 = -9.961e-12
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+41
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 1.4472e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 2.0e-11
+ cgso = 2.0e-11
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 0.0
+ cgdl = 0.0
+ cf = 0.0
+ clc = 7.0e-8
+ cle = 0.492
+ dlc = -1.2e-8
+ dwc = 0.0
+ vfbcv = -1.0
+ acde = 0.44
+ moin = 8.7
+ noff = 2.6123
+ voffcv = 0.112
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007653568198
+ mjs = 0.3362
+ pbs = 0.6587
+ cjsws = 9.1602368e-11
+ mjsws = 0.2659
+ pbsws = 0.7418
+ cjswgs = 2.39155046e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 2.74e-6
+ sbref = 2.74e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.6 pmos
* DC IV MOS Parameters
+ lmin = 5e-07 lmax = 1e-06 wmin = 7e-06 wmax = 1.0e-4
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 2.8e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 7.476e-9
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -7.916e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25000000.0
+ tnoib = 0.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.23e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope2/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-4.736924432e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 5.667526318e-9
+ k1 = 0.64774
+ k2 = -6.468823488e-02 lk2 = 6.423262045e-9
+ k3 = 3.39
+ dvt0 = 2.4422
+ dvt1 = 0.16136
+ dvt2 = 0.026237
+ dvt0w = 0.5
+ dvt1w = 1928100.0
+ dvt2w = -0.032
+ w0 = 1.0e-8
+ k3b = 1.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 6.320409760e+04 lvsat = 2.775062375e-2
+ ua = -2.789854560e-09 lua = -7.502294554e-17
+ ub = 2.825072160e-18 lub = 1.468011241e-25
+ uc = 7.576047360e-11 luc = -3.118909348e-18
+ rdsw = 484.7
+ prwb = 0.1
+ prwg = 0.052
+ wr = 1.0
+ u0 = 3.245856438e-03 lu0 = -1.874885354e-11
+ a0 = 1.201400147e+00 la0 = -6.609393678e-8
+ keta = -0.01258
+ a1 = 0.0
+ a2 = 0.46703705
+ ags = 9.522773600e-01 lags = -2.627277988e-7
+ b0 = 7.305551040e-07 lb0 = -7.264639954e-13
+ b1 = 2.1073e-24
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-2.108370400e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = 1.430647258e-8
+ nfactor = {1.451035064e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 1.064475304e-6
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -6.393105e-11
+ cdsc = 2.8125e-7
+ cdscb = 1.0e-4
+ cdscd = 1.0e-10
+ eta0 = 0.2
+ etab = -0.00025
+ dsub = 1.0
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.030097
+ pdiblc1 = 0.0
+ pdiblc2 = -2.274734080e-02 lpdiblc2 = 3.789592849e-08 ppdiblc2 = 2.524354897e-29
+ pdiblcb = -0.025
+ drout = 0.43496
+ pscbe1 = 800000000.0
+ pscbe2 = 8.6797e-9
+ pvag = 0.0
+ delta = 2.136885600e-02 ldelta = 1.131243759e-8
+ alpha0 = 5.0449517e-13
+ alpha1 = -4.0583656e-18
+ beta0 = 6.2016506
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -8.993837920e-01 lkt1 = 2.300834765e-9
+ kt2 = -1.576964320e-02 lkt2 = -1.989730440e-8
+ at = 1.920565792e+05 lat = -6.561705436e-2
+ ute = -5.958848000e-02 lute = -1.675479675e-7
+ ua1 = 4.288626720e-10 lua1 = 2.311257350e-16
+ ub1 = 5.703157168e-19 lub1 = -5.782184584e-25 wub1 = 2.295887404e-40 pub1 = 2.299005293e-46
+ uc1 = -2.284941472e-11 luc1 = 1.281623960e-17
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+41
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 1.4472e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 2.0e-11
+ cgso = 2.0e-11
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 0.0
+ cgdl = 0.0
+ cf = 0.0
+ clc = 7.0e-8
+ cle = 0.492
+ dlc = -1.2e-8
+ dwc = 0.0
+ vfbcv = -1.0
+ acde = 0.44
+ moin = 8.7
+ noff = 2.6123
+ voffcv = 0.112
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007653568198
+ mjs = 0.3362
+ pbs = 0.6587
+ cjsws = 9.1602368e-11
+ mjsws = 0.2659
+ pbsws = 0.7418
+ cjswgs = 2.39155046e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 1.74e-6
+ sbref = 1.74e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.7 pmos
* DC IV MOS Parameters
+ lmin = 3.5e-07 lmax = 5e-07 wmin = 7e-06 wmax = 1.0e-4
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 2.8e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 7.476e-9
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -7.916e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25000000.0
+ tnoib = 0.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.23e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope3/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-4.495229360e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope1/sqrt(l*w*mult))} lvth0 = -6.281878042e-9
+ k1 = 0.64774
+ k2 = -5.754312472e-02 lk2 = 2.890719582e-9
+ k3 = 3.39
+ dvt0 = 2.4422
+ dvt1 = 0.16136
+ dvt2 = 0.026237
+ dvt0w = 0.5
+ dvt1w = 1928100.0
+ dvt2w = -0.032
+ w0 = 1.0e-8
+ k3b = 1.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 1.517833680e+05 lvsat = -1.604296754e-2
+ ua = -3.074079200e-09 lua = 6.549771648e-17
+ ub = 3.030160000e-18 lub = 4.540569600e-26
+ uc = 8.394894400e-11 luc = -7.167289114e-18
+ rdsw = 484.7
+ prwb = 0.1
+ prwg = 0.052
+ wr = 1.0
+ u0 = 2.306985896e-03 lu0 = 4.454287426e-10
+ a0 = 1.223188640e+00 la0 = -7.686616762e-8
+ keta = -0.01258
+ a1 = 0.0
+ a2 = 0.46703705
+ ags = 4.111120000e-01 lags = 4.824355200e-9
+ b0 = -2.435183680e-06 lb0 = 8.386772594e-13
+ b1 = 2.1073e-24
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {1.575636000e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = -1.678308038e-7
+ nfactor = {9.168616000e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 1.328570665e-6
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -6.393105e-11
+ cdsc = 2.8125e-7
+ cdscb = 1.0e-4
+ cdscd = 1.0e-10
+ eta0 = 0.2
+ etab = -0.00025
+ dsub = 1.0
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.030097
+ pdiblc1 = 0.0
+ pdiblc2 = -8.848803200e-02 lpdiblc2 = 7.039812622e-8
+ pdiblcb = -0.025
+ drout = 0.43496
+ pscbe1 = 800000000.0
+ pscbe2 = 8.6797e-9
+ pvag = 0.0
+ delta = 2.489701600e-02 ldelta = 9.568115290e-9
+ alpha0 = 5.0449517e-13
+ alpha1 = -4.0583656e-18
+ beta0 = 6.2016506
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -1.111334640e+00 lkt1 = 1.070893340e-7
+ kt2 = -0.056015
+ at = 1.376778160e+05 lat = -3.873219383e-2
+ ute = -0.39848
+ ua1 = 8.9635e-10
+ ub1 = -5.9922e-19
+ uc1 = 3.0734e-12
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+41
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 1.4472e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 2.0e-11
+ cgso = 2.0e-11
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 0.0
+ cgdl = 0.0
+ cf = 0.0
+ clc = 7.0e-8
+ cle = 0.492
+ dlc = -1.2e-8
+ dwc = 0.0
+ vfbcv = -1.0
+ acde = 0.44
+ moin = 8.7
+ noff = 2.6123
+ voffcv = 0.112
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007653568198
+ mjs = 0.3362
+ pbs = 0.6587
+ cjsws = 9.1602368e-11
+ mjsws = 0.2659
+ pbsws = 0.7418
+ cjswgs = 2.39155046e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 1.44e-6
+ sbref = 1.44e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.8 pmos
* DC IV MOS Parameters
+ lmin = 2.0e-05 lmax = 1.0e-04 wmin = 5.0e-06 wmax = 7.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 2.8e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 7.476e-9
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -7.916e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25000000.0
+ tnoib = 0.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.23e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-4.864066587e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} wvth0 = 2.511450168e-7
+ k1 = 0.64774
+ k2 = -5.162411567e-02 wk2 = 4.001954494e-8
+ k3 = 3.39
+ dvt0 = 2.4422
+ dvt1 = 0.16136
+ dvt2 = 0.026237
+ dvt0w = 0.5
+ dvt1w = 1928100.0
+ dvt2w = -0.032
+ w0 = 1.0e-8
+ k3b = 1.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 123760.0
+ ua = -3.121800871e-09 wua = 8.130656698e-16
+ ub = 3.232079581e-18 wub = -1.328413503e-24
+ uc = 5.087094712e-11 wuc = -1.060293347e-17
+ rdsw = 484.7
+ prwb = 0.1
+ prwg = 0.052
+ wr = 1.0
+ u0 = 2.601261512e-03 wu0 = -5.168573152e-10
+ a0 = 1.735423680e+00 wa0 = 3.229629159e-7
+ keta = -0.01258
+ a1 = 0.0
+ a2 = 0.46703705
+ ags = 4.347676458e-01 wags = -3.070672209e-7
+ b0 = 0.0
+ b1 = 2.1073e-24
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.1819+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))}
+ nfactor = {3.619727292e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} wnfactor = 2.508838608e-6
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -6.393105e-11
+ cdsc = 2.8125e-7
+ cdscb = 1.0e-4
+ cdscd = 1.0e-10
+ eta0 = 0.2
+ etab = -0.00025
+ dsub = 1.0
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.030097
+ pdiblc1 = 0.0
+ pdiblc2 = 2.350837605e-03 wpdiblc2 = -3.522123876e-9
+ pdiblcb = -0.025
+ drout = 0.43496
+ pscbe1 = 800000000.0
+ pscbe2 = 8.6797e-9
+ pvag = 0.0
+ delta = 3.485427320e-03 wdelta = 7.086032711e-8
+ alpha0 = 5.0449517e-13
+ alpha1 = -4.0583656e-18
+ beta0 = 6.2016506
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -7.937810322e-01 wkt1 = -1.935340040e-6
+ kt2 = -0.055045
+ at = 285600.0
+ ute = -0.22271
+ ua1 = 6.8217e-10
+ ub1 = -1.4864e-19
+ uc1 = -9.961e-12
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+41
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 1.4472e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 2.0e-11
+ cgso = 2.0e-11
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 0.0
+ cgdl = 0.0
+ cf = 0.0
+ clc = 7.0e-8
+ cle = 0.492
+ dlc = -1.2e-8
+ dwc = 0.0
+ vfbcv = -1.0
+ acde = 0.44
+ moin = 8.7
+ noff = 2.6123
+ voffcv = 0.112
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007653568198
+ mjs = 0.3362
+ pbs = 0.6587
+ cjsws = 9.1602368e-11
+ mjsws = 0.2659
+ pbsws = 0.7418
+ cjswgs = 2.39155046e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.9 pmos
* DC IV MOS Parameters
+ lmin = 8e-06 lmax = 2.0e-05 wmin = 5.0e-06 wmax = 7.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 2.8e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 7.476e-9
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -7.916e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25000000.0
+ tnoib = 0.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.23e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-4.864066587e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} wvth0 = 2.511450168e-7
+ k1 = 0.64774
+ k2 = -5.162411567e-02 wk2 = 4.001954494e-8
+ k3 = 3.39
+ dvt0 = 2.4422
+ dvt1 = 0.16136
+ dvt2 = 0.026237
+ dvt0w = 0.5
+ dvt1w = 1928100.0
+ dvt2w = -0.032
+ w0 = 1.0e-8
+ k3b = 1.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 123760.0
+ ua = -3.121800871e-09 wua = 8.130656698e-16
+ ub = 3.232079581e-18 wub = -1.328413503e-24
+ uc = 5.087094712e-11 wuc = -1.060293347e-17
+ rdsw = 484.7
+ prwb = 0.1
+ prwg = 0.052
+ wr = 1.0
+ u0 = 2.601261512e-03 wu0 = -5.168573152e-10
+ a0 = 1.735423680e+00 wa0 = 3.229629159e-7
+ keta = -0.01258
+ a1 = 0.0
+ a2 = 0.46703705
+ ags = 4.347676458e-01 wags = -3.070672209e-7
+ b0 = 0.0
+ b1 = 2.1073e-24
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.1819+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))}
+ nfactor = {3.619727292e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} wnfactor = 2.508838608e-6
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -6.393105e-11
+ cdsc = 2.8125e-7
+ cdscb = 1.0e-4
+ cdscd = 1.0e-10
+ eta0 = 0.2
+ etab = -0.00025
+ dsub = 1.0
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.030097
+ pdiblc1 = 0.0
+ pdiblc2 = 2.350837605e-03 wpdiblc2 = -3.522123876e-9
+ pdiblcb = -0.025
+ drout = 0.43496
+ pscbe1 = 800000000.0
+ pscbe2 = 8.6797e-9
+ pvag = 0.0
+ delta = 3.485427320e-03 wdelta = 7.086032711e-8
+ alpha0 = 5.0449517e-13
+ alpha1 = -4.0583656e-18
+ beta0 = 6.2016506
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -7.937810322e-01 wkt1 = -1.935340040e-6
+ kt2 = -0.055045
+ at = 285600.0
+ ute = -0.22271
+ ua1 = 6.8217e-10
+ ub1 = -1.4864e-19
+ uc1 = -9.961e-12
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+41
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 1.4472e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 2.0e-11
+ cgso = 2.0e-11
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 0.0
+ cgdl = 0.0
+ cf = 0.0
+ clc = 7.0e-8
+ cle = 0.492
+ dlc = -1.2e-8
+ dwc = 0.0
+ vfbcv = -1.0
+ acde = 0.44
+ moin = 8.7
+ noff = 2.6123
+ voffcv = 0.112
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007653568198
+ mjs = 0.3362
+ pbs = 0.6587
+ cjsws = 9.1602368e-11
+ mjsws = 0.2659
+ pbsws = 0.7418
+ cjswgs = 2.39155046e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.10 pmos
* DC IV MOS Parameters
+ lmin = 4e-06 lmax = 8e-06 wmin = 5.0e-06 wmax = 7.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 2.8e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 7.476e-9
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -7.916e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25000000.0
+ tnoib = 0.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.23e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-4.976203840e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 8.964700585e-08 wvth0 = 2.721994934e-07 pvth0 = -1.683179073e-13
+ k1 = 0.64774
+ k2 = -5.633546139e-02 lk2 = 3.766438225e-08 wk2 = 7.106403157e-08 pk2 = -2.481820440e-13
+ k3 = 3.39
+ dvt0 = 2.4422
+ dvt1 = 0.16136
+ dvt2 = 0.026237
+ dvt0w = 0.5
+ dvt1w = 1928100.0
+ dvt2w = -0.032
+ w0 = 1.0e-8
+ k3b = 1.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 123760.0
+ ua = -3.327222541e-09 lua = 1.642222999e-15 wua = 1.837102555e-15 pua = -8.186560478e-21
+ ub = 3.543176576e-18 lub = -2.487033812e-24 wub = -2.879246953e-24 pub = 1.239798293e-29
+ uc = 1.049460290e-11 luc = 3.227846462e-16 wuc = 1.906750805e-16 puc = -1.609096955e-21
+ rdsw = 484.7
+ prwb = 0.1
+ prwg = 0.052
+ wr = 1.0
+ u0 = 2.367015281e-03 lu0 = 1.872658069e-09 wu0 = 5.282914208e-10 pu0 = -8.355337055e-15
+ a0 = 2.052385610e+00 la0 = -2.533920451e-06 wa0 = -1.197271129e-06 pa0 = 1.215335905e-11
+ keta = -0.01258
+ a1 = 0.0
+ a2 = 0.46703705
+ ags = 4.830764275e-01 lags = -3.861997247e-07 wags = -7.535577347e-07 pags = 3.569423763e-12
+ b0 = 0.0
+ b1 = 2.1073e-24
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.1819+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))}
+ nfactor = {4.037686987e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -3.341336988e-06 wnfactor = 2.882464290e-06 pnfactor = -2.986913152e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -6.393105e-11
+ cdsc = 2.8125e-7
+ cdscb = 1.0e-4
+ cdscd = 1.0e-10
+ eta0 = 0.2
+ etab = -0.00025
+ dsub = 1.0
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.030097
+ pdiblc1 = 0.0
+ pdiblc2 = -1.270175929e-04 lpdiblc2 = 1.980896560e-08 wpdiblc2 = 1.410291480e-09 ppdiblc2 = -3.943170132e-14
+ pdiblcb = -0.025
+ drout = 0.43496
+ pscbe1 = 800000000.0
+ pscbe2 = 8.6797e-9
+ pvag = 0.0
+ delta = -1.193099316e-02 ldelta = 1.232450319e-07 wdelta = 1.242701966e-07 pdelta = -4.269798606e-13
+ alpha0 = 5.0449517e-13
+ alpha1 = -4.0583656e-18
+ beta0 = 6.2016506
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -5.778878873e-01 lkt1 = -1.725936157e-06 wkt1 = -3.886921371e-06 pkt1 = 1.560172179e-11
+ kt2 = -0.055045
+ at = 2.991709740e+05 lat = -1.084917945e-1
+ ute = -3.123143780e-01 lute = 7.163332395e-7
+ ua1 = 6.682694880e-10 lua1 = 1.111262531e-16
+ ub1 = -1.753625360e-19 lub1 = 2.136306418e-25
+ uc1 = -9.961e-12
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+41
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 1.4472e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 2.0e-11
+ cgso = 2.0e-11
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 0.0
+ cgdl = 0.0
+ cf = 0.0
+ clc = 7.0e-8
+ cle = 0.492
+ dlc = -1.2e-8
+ dwc = 0.0
+ vfbcv = -1.0
+ acde = 0.44
+ moin = 8.7
+ noff = 2.6123
+ voffcv = 0.112
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007653568198
+ mjs = 0.3362
+ pbs = 0.6587
+ cjsws = 9.1602368e-11
+ mjsws = 0.2659
+ pbsws = 0.7418
+ cjswgs = 2.39155046e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.11 pmos
* DC IV MOS Parameters
+ lmin = 2e-06 lmax = 4e-06 wmin = 5.0e-06 wmax = 7.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 2.8e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 7.476e-9
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -7.916e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25000000.0
+ tnoib = 0.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.23e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-4.007508083e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -2.972888276e-07 wvth0 = -1.464263719e-07 pvth0 = 1.503841249e-12
+ k1 = 0.64774
+ k2 = -2.728337775e-02 lk2 = -7.838126065e-08 wk2 = -8.051221679e-08 pk2 = 3.572741225e-13
+ k3 = 3.39
+ dvt0 = 2.4422
+ dvt1 = 0.16136
+ dvt2 = 0.026237
+ dvt0w = 0.5
+ dvt1w = 1928100.0
+ dvt2w = -0.032
+ w0 = 1.0e-8
+ k3b = 1.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 2.387323757e+05 lvsat = -4.592456576e-01 wvsat = -5.731428116e-01 pvsat = 2.289361647e-6
+ ua = -3.645202145e-09 lua = 2.912360732e-15 wua = 3.716534667e-15 pua = -1.569376411e-20
+ ub = 3.994770385e-18 lub = -4.290880126e-24 wub = -5.720035029e-24 pub = 2.374522682e-29
+ uc = 1.110001615e-10 luc = -7.867475726e-17 wuc = -3.466985627e-16 puc = 5.373883255e-22
+ rdsw = 484.7
+ prwb = 0.1
+ prwg = 0.052
+ wr = 1.0
+ u0 = 1.838762253e-03 lu0 = 3.982711963e-09 wu0 = 3.353247459e-09 pu0 = -1.963934145e-14
+ a0 = 3.436131446e+00 la0 = -8.061154820e-06 wa0 = -8.089199214e-06 pa0 = 3.968247659e-11
+ keta = -0.01258
+ a1 = 0.0
+ a2 = 0.46703705
+ ags = 6.590416397e-01 lags = -1.089075168e-06 wags = -1.659590005e-06 pags = 7.188479064e-12
+ b0 = 0.0
+ b1 = 2.1073e-24
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.1819+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))}
+ nfactor = {9.338606487e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 9.056586937e-06 wnfactor = 1.693410737e-05 pnfactor = -5.911479629e-11
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -6.393105e-11
+ cdsc = 2.8125e-7
+ cdscb = 1.0e-4
+ cdscd = 1.0e-10
+ eta0 = 0.2
+ etab = -0.00025
+ dsub = 1.0
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.030097
+ pdiblc1 = 0.0
+ pdiblc2 = 2.375208404e-03 lpdiblc2 = 9.814074073e-09 wpdiblc2 = -1.474810800e-08 ppdiblc2 = 2.511140956e-14
+ pdiblcb = -0.025
+ drout = 0.43496
+ pscbe1 = 800000000.0
+ pscbe2 = 8.6797e-9
+ pvag = 0.0
+ delta = 3.346518452e-02 ldelta = -5.808546025e-08 wdelta = -9.629114790e-08 pdelta = 4.540303739e-13
+ alpha0 = 5.0449517e-13
+ alpha1 = -4.0583656e-18
+ beta0 = 6.2016506
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -1.041581005e+00 lkt1 = 1.262396339e-07 wkt1 = -5.741392715e-08 pkt1 = 3.051372606e-13
+ kt2 = -0.055045
+ at = 5.814493013e+05 lat = -1.236024345e+00 wat = -1.420877490e+00 pat = 5.675553047e-6
+ ute = -0.13298
+ ua1 = 6.9609e-10
+ ub1 = -2.449776196e-19 lub1 = 4.917011319e-25 wub1 = 6.136475426e-25 pub1 = -2.451153744e-30
+ uc1 = -9.961e-12
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+41
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 1.4472e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 2.0e-11
+ cgso = 2.0e-11
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 0.0
+ cgdl = 0.0
+ cf = 0.0
+ clc = 7.0e-8
+ cle = 0.492
+ dlc = -1.2e-8
+ dwc = 0.0
+ vfbcv = -1.0
+ acde = 0.44
+ moin = 8.7
+ noff = 2.6123
+ voffcv = 0.112
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007653568198
+ mjs = 0.3362
+ pbs = 0.6587
+ cjsws = 9.1602368e-11
+ mjsws = 0.2659
+ pbsws = 0.7418
+ cjswgs = 2.39155046e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.12 pmos
* DC IV MOS Parameters
+ lmin = 1.5e-06 lmax = 2e-06 wmin = 5.0e-06 wmax = 7.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 2.8e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 7.476e-9
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -7.916e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25000000.0
+ tnoib = 0.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.23e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-6.227728571e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 1.455119467e-07 wvth0 = 1.079365757e-06 pvth0 = -9.408785732e-13
+ k1 = 0.64774
+ k2 = -5.030940708e-02 lk2 = -3.245814775e-08 wk2 = 4.003517730e-08 pk2 = 1.168543997e-13
+ k3 = 3.39
+ dvt0 = 2.4422
+ dvt1 = 0.16136
+ dvt2 = 0.026237
+ dvt0w = 0.5
+ dvt1w = 1928100.0
+ dvt2w = -0.032
+ w0 = 1.0e-8
+ k3b = 1.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = -3.876929948e+05 lvsat = 7.900971013e-01 wvsat = 3.341933314e+00 pvsat = -5.518866177e-6
+ ua = -4.901468211e-10 lua = -3.380081607e-15 wua = -1.218677007e-14 pua = 1.602378686e-20
+ ub = -8.162212032e-19 lub = 5.304161498e-24 wub = 1.849768064e-23 pub = -2.455458531e-29
+ uc = 5.303659099e-11 luc = 3.692778787e-17 wuc = -1.784603584e-16 puc = 2.018540508e-22
+ rdsw = 484.7
+ prwb = 0.1
+ prwg = 0.052
+ wr = 1.0
+ u0 = 5.325683390e-03 lu0 = -2.971603552e-09 wu0 = -1.519914233e-08 pu0 = 1.736154475e-14
+ a0 = -8.494784464e-01 la0 = 4.860655492e-07 wa0 = 1.350735700e-05 pa0 = -3.389695120e-12
+ keta = -0.01258
+ a1 = 0.0
+ a2 = 0.46703705
+ ags = 3.380521997e-01 lags = -4.488938291e-07 wags = -1.244140928e-06 pags = 6.359907426e-12
+ b0 = 0.0
+ b1 = 2.1073e-24
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.1819+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))}
+ nfactor = {9.971838909e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -8.968756906e-06 wnfactor = -3.360714511e-05 pnfactor = 4.168467766e-11
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -6.393105e-11
+ cdsc = 2.8125e-7
+ cdscb = 1.0e-4
+ cdscd = 1.0e-10
+ eta0 = 0.2
+ etab = -0.00025
+ dsub = 1.0
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.030097
+ pdiblc1 = 0.0
+ pdiblc2 = -6.755076593e-03 lpdiblc2 = 2.802351447e-08 wpdiblc2 = 2.428244614e-08 ppdiblc2 = -5.273112762e-14
+ pdiblcb = -0.025
+ drout = 0.43496
+ pscbe1 = 800000000.0
+ pscbe2 = 8.6797e-9
+ pvag = 0.0
+ delta = -6.396132487e-03 ldelta = 2.141395040e-08 wdelta = 1.632076225e-07 pdelta = -6.351397383e-14
+ alpha0 = 5.0449517e-13
+ alpha1 = -4.0583656e-18
+ beta0 = 6.2016506
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -9.231123693e-01 lkt1 = -1.100342140e-07 wkt1 = -3.259101484e-07 pkt1 = 8.406261243e-13
+ kt2 = -2.067721383e-01 lkt2 = 3.026046046e-07 wkt2 = 1.059821344e-06 pkt2 = -2.113707688e-12
+ at = -8.460038989e+05 lat = 1.610888317e+00 wat = 7.347107366e+00 pat = -1.181131595e-5
+ ute = -0.13298
+ ua1 = 8.464370986e-10 lua1 = -2.998522535e-16 wua1 = -3.236651818e-16 pua1 = 6.455178386e-22
+ ub1 = 3.893300660e-20 lub1 = -7.453022106e-26 wub1 = -2.454590171e-24 pub1 = 3.668139551e-30
+ uc1 = -9.961e-12
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+41
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 1.4472e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 2.0e-11
+ cgso = 2.0e-11
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 0.0
+ cgdl = 0.0
+ cf = 0.0
+ clc = 7.0e-8
+ cle = 0.492
+ dlc = -1.2e-8
+ dwc = 0.0
+ vfbcv = -1.0
+ acde = 0.44
+ moin = 8.7
+ noff = 2.6123
+ voffcv = 0.112
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007653568198
+ mjs = 0.3362
+ pbs = 0.6587
+ cjsws = 9.1602368e-11
+ mjsws = 0.2659
+ pbsws = 0.7418
+ cjswgs = 2.39155046e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.13 pmos
* DC IV MOS Parameters
+ lmin = 1e-06 lmax = 1.5e-06 wmin = 5.0e-06 wmax = 7.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 2.8e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 7.476e-9
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -7.916e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25000000.0
+ tnoib = 0.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.23e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-4.935826571e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -4.754988830e-08 wvth0 = 3.244867020e-07 pvth0 = 1.872126869e-13
+ k1 = 0.64774
+ k2 = -4.988764066e-02 lk2 = -3.308843548e-08 wk2 = 6.991563826e-09 pk2 = 1.662347757e-13
+ k3 = 3.39
+ dvt0 = 2.4422
+ dvt1 = 0.16136
+ dvt2 = 0.026237
+ dvt0w = 0.5
+ dvt1w = 1928100.0
+ dvt2w = -0.032
+ w0 = 1.0e-8
+ k3b = 1.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 4.247553090e+05 lvsat = -4.240256438e-01 wvsat = -2.338099832e+00 pvsat = 2.969375355e-6
+ ua = -3.222586688e-09 lua = 7.032765301e-16 wua = 4.852180921e-16 pua = -2.913232247e-21
+ ub = 3.124193358e-18 lub = -5.843940213e-25 wub = 1.171817404e-25 pub = 2.913232247e-30
+ uc = 1.040374915e-10 luc = -3.928795792e-17 wuc = -2.421388260e-16 puc = 2.970151527e-22
+ rdsw = 484.7
+ prwb = 0.1
+ prwg = 0.052
+ wr = 1.0
+ u0 = 1.749608033e-03 lu0 = 2.372483462e-09 wu0 = 1.915959340e-09 pu0 = -8.215263193e-15
+ a0 = -1.962563685e+00 la0 = 2.149460130e-06 wa0 = 2.058954781e-05 pa0 = -1.397332106e-11
+ keta = -0.01258
+ a1 = 0.0
+ a2 = 0.46703705
+ ags = -1.641173666e+00 lags = 2.508861305e-06 wags = 1.169282474e-05 pags = -1.297309407e-11
+ b0 = 0.0
+ b1 = 2.1073e-24
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-8.083669331e-02+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = -1.510290055e-07 wvoff = -5.038054349e-07 pvoff = 7.528868419e-13
+ nfactor = {6.503925356e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -3.786306893e-06 wnfactor = -1.464751090e-05 pnfactor = 1.335140031e-11
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -6.393105e-11
+ cdsc = 2.8125e-7
+ cdscb = 1.0e-4
+ cdscd = 1.0e-10
+ eta0 = 0.2
+ etab = -0.00025
+ dsub = 1.0
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.030097
+ pdiblc1 = 0.0
+ pdiblc2 = 1.739099758e-02 lpdiblc2 = -8.060378777e-09 wpdiblc2 = -1.173045881e-07 ppdiblc2 = 1.588565364e-13
+ pdiblcb = -0.025
+ drout = 0.43496
+ pscbe1 = 800000000.0
+ pscbe2 = 8.6797e-9
+ pvag = 0.0
+ delta = 5.502178720e-03 ldelta = 3.633114129e-09 wdelta = 3.306839408e-08 pdelta = 1.309660891e-13
+ alpha0 = 5.0449517e-13
+ alpha1 = -4.0583656e-18
+ beta0 = 6.2016506
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -1.170931772e+00 lkt1 = 2.603071021e-07 wkt1 = 5.392368520e-07 pkt1 = -4.522495531e-13
+ kt2 = 5.836591748e-02 lkt2 = -9.361770594e-08 wkt2 = -1.059821344e-06 pkt2 = 1.053886344e-12
+ at = 9.371843412e+05 lat = -1.053908189e+00 wat = -5.118906295e+00 pat = 6.817894865e-6
+ ute = 3.430240933e-01 lute = -7.113405170e-07 wute = -2.003795225e-06 pute = 2.994471584e-12
+ ua1 = 5.166036478e-10 lua1 = 1.930508554e-16 wua1 = 1.010641115e-15 pua1 = -1.348469491e-21
+ ub1 = -9.418840951e-21 lub1 = -2.273220083e-27 wub1 = -7.583050876e-27 pub1 = 1.133211123e-32
+ uc1 = -9.961e-12
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+41
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 1.4472e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 2.0e-11
+ cgso = 2.0e-11
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 0.0
+ cgdl = 0.0
+ cf = 0.0
+ clc = 7.0e-8
+ cle = 0.492
+ dlc = -1.2e-8
+ dwc = 0.0
+ vfbcv = -1.0
+ acde = 0.44
+ moin = 8.7
+ noff = 2.6123
+ voffcv = 0.112
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007653568198
+ mjs = 0.3362
+ pbs = 0.6587
+ cjsws = 9.1602368e-11
+ mjsws = 0.2659
+ pbsws = 0.7418
+ cjswgs = 2.39155046e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 2.74e-6
+ sbref = 2.74e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.14 pmos
* DC IV MOS Parameters
+ lmin = 5e-07 lmax = 1e-06 wmin = 5.0e-06 wmax = 7.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 2.8e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 7.476e-9
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -7.916e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25000000.0
+ tnoib = 0.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.23e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope2/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-5.711617328e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 2.959474459e-08 wvth0 = 6.808276664e-07 pvth0 = -1.671327682e-13
+ k1 = 0.64774
+ k2 = -1.133864848e-01 lk2 = 3.005481509e-08 wk2 = 3.401596130e-07 pk2 = -1.650675323e-13
+ k3 = 3.39
+ dvt0 = 2.4422
+ dvt1 = 0.16136
+ dvt2 = 0.026237
+ dvt0w = 0.5
+ dvt1w = 1928100.0
+ dvt2w = -0.032
+ w0 = 1.0e-8
+ k3b = 1.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 9.656614278e+03 lvsat = -1.125150179e-02 wvsat = 3.740317413e-01 pvsat = 2.724317190e-7
+ ua = -1.775445946e-09 lua = -7.357602237e-16 wua = -7.085692860e-15 pua = 4.615281603e-21
+ ub = 1.488559256e-18 lub = 1.042080530e-24 wub = 9.335606789e-24 pub = -6.253569621e-30
+ uc = 3.651704314e-11 luc = 2.785437597e-17 wuc = 2.741172454e-16 puc = -2.163498847e-22
+ rdsw = 484.7
+ prwb = 0.1
+ prwg = 0.052
+ wr = 1.0
+ u0 = 5.225760367e-03 lu0 = -1.084202419e-09 wu0 = -1.382972398e-08 pu0 = 7.442244299e-15
+ a0 = 9.222606696e-01 la0 = -7.192092085e-07 wa0 = 1.949802650e-06 pa0 = 4.562041523e-12
+ keta = -0.01258
+ a1 = 0.0
+ a2 = 0.46703705
+ ags = 1.140259026e+00 lags = -2.569953637e-07 wags = -1.313060957e-06 pags = -4.004133409e-14
+ b0 = -5.063575781e-07 lb0 = 5.035219756e-13 wb0 = 8.639894456e-12 pb0 = -8.591511047e-18
+ b1 = 2.1073e-24
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-2.829633067e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = 4.996569883e-08 wvoff = 5.038054349e-07 pvoff = -2.490814070e-13
+ nfactor = {1.252649687e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 1.435561633e-06 wnfactor = 1.385731381e-06 pnfactor = -2.592055819e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -6.393105e-11
+ cdsc = 2.8125e-7
+ cdscb = 1.0e-4
+ cdscd = 1.0e-10
+ eta0 = 0.2
+ etab = -0.00025
+ dsub = 1.0
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.030097
+ pdiblc1 = 0.0
+ pdiblc2 = -4.153656099e-02 lpdiblc2 = 5.053718547e-08 wpdiblc2 = 1.312436049e-07 ppdiblc2 = -8.829978676e-14
+ pdiblcb = -0.025
+ drout = 0.43496
+ pscbe1 = 800000000.0
+ pscbe2 = 8.6797e-9
+ pvag = 0.0
+ delta = 4.106256910e-03 ldelta = 5.021218777e-09 wdelta = 1.205800832e-07 pdelta = 4.394446541e-14
+ alpha0 = 5.0449517e-13
+ alpha1 = -4.0583656e-18
+ beta0 = 6.2016506
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -9.049659690e-01 lkt1 = -4.169292885e-09 wkt1 = 3.899177422e-08 pkt1 = 4.519415220e-14
+ kt2 = -1.576964320e-02 lkt2 = -1.989730440e-8
+ at = -3.026155963e+05 lat = 1.789488692e-01 wat = 3.455308890e+00 pat = -1.708304715e-6
+ ute = -3.464576933e-01 lute = -2.571982844e-08 wute = 2.003795225e-06 pute = -9.906763590e-13
+ ua1 = 5.272121655e-10 lua1 = 1.825017454e-16 wua1 = -6.869759332e-16 pua1 = 3.396409014e-22
+ ub1 = 5.692301050e-19 lub1 = -5.776817319e-25 wub1 = 7.583050876e-27 pub1 = -3.749060353e-33
+ uc1 = -2.284941472e-11 luc1 = 1.281623960e-17
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+41
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 1.4472e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 2.0e-11
+ cgso = 2.0e-11
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 0.0
+ cgdl = 0.0
+ cf = 0.0
+ clc = 7.0e-8
+ cle = 0.492
+ dlc = -1.2e-8
+ dwc = 0.0
+ vfbcv = -1.0
+ acde = 0.44
+ moin = 8.7
+ noff = 2.6123
+ voffcv = 0.112
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007653568198
+ mjs = 0.3362
+ pbs = 0.6587
+ cjsws = 9.1602368e-11
+ mjsws = 0.2659
+ pbsws = 0.7418
+ cjswgs = 2.39155046e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 1.74e-6
+ sbref = 1.74e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.15 pmos
* DC IV MOS Parameters
+ lmin = 3.5e-07 lmax = 5e-07 wmin = 5.0e-06 wmax = 7.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 2.8e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 7.476e-9
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -7.916e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25000000.0
+ tnoib = 0.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.23e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope3/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-5.083989650e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -1.435167788e-09 wvth0 = 4.112518889e-07 pvth0 = -3.385450377e-14
+ k1 = 0.64774
+ k2 = -4.397542706e-02 lk2 = -4.262011839e-09 wk2 = -9.477101943e-08 pk2 = 4.996217230e-14
+ k3 = 3.39
+ dvt0 = 2.4422
+ dvt1 = 0.16136
+ dvt2 = 0.026237
+ dvt0w = 0.5
+ dvt1w = 1928100.0
+ dvt2w = -0.032
+ w0 = 1.0e-8
+ k3b = 1.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = -2.762935712e+05 lvsat = 1.301222699e-01 wvsat = 2.990137968e+00 pvsat = -1.020971199e-6
+ ua = -4.135503596e-09 lua = 4.310522785e-16 wua = 7.414100356e-15 pua = -2.553416163e-21
+ ub = 4.593542837e-18 lub = -4.930233532e-25 wub = -1.092030416e-23 pub = 3.760952753e-30
+ uc = 1.610911660e-10 luc = -3.373507037e-17 wuc = -5.388421234e-16 puc = 1.855772273e-22
+ rdsw = 484.7
+ prwb = 0.1
+ prwg = 0.052
+ wr = 1.0
+ u0 = 1.155112769e-03 lu0 = 9.283257532e-10 wu0 = 8.045889083e-09 pu0 = -3.373058798e-15
+ a0 = -4.050956890e+00 la0 = 1.739549553e-06 wa0 = 3.684015968e-05 pa0 = -1.268775100e-11
+ keta = -0.01258
+ a1 = 0.0
+ a2 = 0.46703705
+ ags = 1.093466766e+00 lags = -2.338612706e-07 wags = -4.766280794e-06 pags = 1.667230553e-12
+ b0 = 1.687858594e-06 lb0 = -5.812984996e-13 wb0 = -2.879964819e-11 pb0 = 9.918598835e-18
+ b1 = 2.1073e-24
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {1.643848634e-02+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = -9.805854764e-08 wvoff = 9.857656930e-07 pvoff = -4.873625586e-13
+ nfactor = {-1.746376765e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 2.918280311e-06 wnfactor = 1.860284781e-05 pnfactor = -1.110419818e-11
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -6.393105e-11
+ cdsc = 2.8125e-7
+ cdscb = 1.0e-4
+ cdscd = 1.0e-10
+ eta0 = 0.2
+ etab = -0.00025
+ dsub = 1.0
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.030097
+ pdiblc1 = 0.0
+ pdiblc2 = -1.576217744e-01 lpdiblc2 = 1.079297150e-07 wpdiblc2 = 4.829025089e-07 ppdiblc2 = -2.621599489e-13
+ pdiblcb = -0.025
+ drout = 0.43496
+ pscbe1 = 800000000.0
+ pscbe2 = 8.6797e-9
+ pvag = 0.0
+ delta = 1.427768939e-03 ldelta = 6.345463229e-09 wdelta = 1.639338172e-07 pdelta = 2.251037933e-14
+ alpha0 = 5.0449517e-13
+ alpha1 = -4.0583656e-18
+ beta0 = 6.2016506
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -1.278453987e+00 lkt1 = 1.804831834e-07 wkt1 = 1.167336663e-06 pkt1 = -5.126595608e-13
+ kt2 = -0.056015
+ at = 1.376778160e+05 lat = -3.873219383e-2
+ ute = -0.39848
+ ua1 = 8.9635e-10
+ ub1 = -5.9922e-19
+ uc1 = 3.0734e-12
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+41
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 1.4472e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 2.0e-11
+ cgso = 2.0e-11
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 0.0
+ cgdl = 0.0
+ cf = 0.0
+ clc = 7.0e-8
+ cle = 0.492
+ dlc = -1.2e-8
+ dwc = 0.0
+ vfbcv = -1.0
+ acde = 0.44
+ moin = 8.7
+ noff = 2.6123
+ voffcv = 0.112
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007653568198
+ mjs = 0.3362
+ pbs = 0.6587
+ cjsws = 9.1602368e-11
+ mjsws = 0.2659
+ pbsws = 0.7418
+ cjswgs = 2.39155046e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 1.44e-6
+ sbref = 1.44e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.16 pmos
* DC IV MOS Parameters
+ lmin = 2.0e-05 lmax = 1.0e-04 wmin = 3.0e-06 wmax = 5.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 2.8e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 7.476e-9
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -7.916e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25000000.0
+ tnoib = 0.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.23e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-4.439836454e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} wvth0 = 3.966425946e-8
+ k1 = 0.64774
+ k2 = -4.300262321e-02 wk2 = -2.959008814e-9
+ k3 = 3.39
+ dvt0 = 2.4422
+ dvt1 = 0.16136
+ dvt2 = 0.026237
+ dvt0w = 0.5
+ dvt1w = 1928100.0
+ dvt2w = -0.032
+ w0 = 1.0e-8
+ k3b = 1.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 123760.0
+ ua = -3.107952400e-09 wua = 7.440303781e-16
+ ub = 3.070076680e-18 wub = -5.208212647e-25
+ uc = 3.055610254e-11 wuc = 9.066754188e-17
+ rdsw = 484.7
+ prwb = 0.1
+ prwg = 0.052
+ wr = 1.0
+ u0 = 2.147941328e-03 wu0 = 1.742965564e-9
+ a0 = 1.797971214e+00 wa0 = 1.116045567e-8
+ keta = -0.01258
+ a1 = 0.0
+ a2 = 0.46703705
+ ags = 3.804833676e-01 wags = -3.645748853e-8
+ b0 = 0.0
+ b1 = 2.1073e-24
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.1819+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))}
+ nfactor = {3.669720461e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} wnfactor = 2.259620258e-6
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -6.393105e-11
+ cdsc = 2.8125e-7
+ cdscb = 1.0e-4
+ cdscd = 1.0e-10
+ eta0 = 0.2
+ etab = -0.00025
+ dsub = 1.0
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.030097
+ pdiblc1 = 0.0
+ pdiblc2 = 7.438602708e-04 wpdiblc2 = 4.488735271e-9
+ pdiblcb = -0.025
+ drout = 0.43496
+ pscbe1 = 800000000.0
+ pscbe2 = 8.6797e-9
+ pvag = 0.0
+ delta = 1.327168129e-02 wdelta = 2.207538132e-8
+ alpha0 = 5.0449517e-13
+ alpha1 = -4.0583656e-18
+ beta0 = 6.2016506
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -1.359142748e+00 wkt1 = 8.830152527e-7
+ kt2 = -0.055045
+ at = 2.898686186e+05 wat = -2.127926881e-2
+ ute = -1.196661430e-01 wute = -5.136785731e-7
+ ua1 = 6.8217e-10
+ ub1 = -1.464161392e-19 wub1 = -1.108605263e-26
+ uc1 = -9.961e-12
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+41
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 1.4472e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 2.0e-11
+ cgso = 2.0e-11
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 0.0
+ cgdl = 0.0
+ cf = 0.0
+ clc = 7.0e-8
+ cle = 0.492
+ dlc = -1.2e-8
+ dwc = 0.0
+ vfbcv = -1.0
+ acde = 0.44
+ moin = 8.7
+ noff = 2.6123
+ voffcv = 0.112
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007653568198
+ mjs = 0.3362
+ pbs = 0.6587
+ cjsws = 9.1602368e-11
+ mjsws = 0.2659
+ pbsws = 0.7418
+ cjswgs = 2.39155046e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.17 pmos
* DC IV MOS Parameters
+ lmin = 8e-06 lmax = 2.0e-05 wmin = 3.0e-06 wmax = 5.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 2.8e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 7.476e-9
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -7.916e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25000000.0
+ tnoib = 0.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.23e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-4.439836454e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} wvth0 = 3.966425946e-8
+ k1 = 0.64774
+ k2 = -4.300262321e-02 wk2 = -2.959008814e-9
+ k3 = 3.39
+ dvt0 = 2.4422
+ dvt1 = 0.16136
+ dvt2 = 0.026237
+ dvt0w = 0.5
+ dvt1w = 1928100.0
+ dvt2w = -0.032
+ w0 = 1.0e-8
+ k3b = 1.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 123760.0
+ ua = -3.107952400e-09 wua = 7.440303781e-16
+ ub = 3.070076680e-18 wub = -5.208212647e-25
+ uc = 3.055610254e-11 wuc = 9.066754188e-17
+ rdsw = 484.7
+ prwb = 0.1
+ prwg = 0.052
+ wr = 1.0
+ u0 = 2.147941328e-03 wu0 = 1.742965564e-9
+ a0 = 1.797971214e+00 wa0 = 1.116045567e-8
+ keta = -0.01258
+ a1 = 0.0
+ a2 = 0.46703705
+ ags = 3.804833676e-01 wags = -3.645748853e-8
+ b0 = 0.0
+ b1 = 2.1073e-24
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.1819+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))}
+ nfactor = {3.669720461e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} wnfactor = 2.259620258e-6
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -6.393105e-11
+ cdsc = 2.8125e-7
+ cdscb = 1.0e-4
+ cdscd = 1.0e-10
+ eta0 = 0.2
+ etab = -0.00025
+ dsub = 1.0
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.030097
+ pdiblc1 = 0.0
+ pdiblc2 = 7.438602708e-04 wpdiblc2 = 4.488735271e-9
+ pdiblcb = -0.025
+ drout = 0.43496
+ pscbe1 = 800000000.0
+ pscbe2 = 8.6797e-9
+ pvag = 0.0
+ delta = 1.327168129e-02 wdelta = 2.207538132e-8
+ alpha0 = 5.0449517e-13
+ alpha1 = -4.0583656e-18
+ beta0 = 6.2016506
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -1.359142748e+00 wkt1 = 8.830152527e-7
+ kt2 = -0.055045
+ at = 2.898686186e+05 wat = -2.127926881e-2
+ ute = -1.196661430e-01 wute = -5.136785731e-7
+ ua1 = 6.8217e-10
+ ub1 = -1.464161392e-19 wub1 = -1.108605263e-26
+ uc1 = -9.961e-12
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+41
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 1.4472e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 2.0e-11
+ cgso = 2.0e-11
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 0.0
+ cgdl = 0.0
+ cf = 0.0
+ clc = 7.0e-8
+ cle = 0.492
+ dlc = -1.2e-8
+ dwc = 0.0
+ vfbcv = -1.0
+ acde = 0.44
+ moin = 8.7
+ noff = 2.6123
+ voffcv = 0.112
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007653568198
+ mjs = 0.3362
+ pbs = 0.6587
+ cjsws = 9.1602368e-11
+ mjsws = 0.2659
+ pbsws = 0.7418
+ cjswgs = 2.39155046e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.18 pmos
* DC IV MOS Parameters
+ lmin = 4e-06 lmax = 8e-06 wmin = 3.0e-06 wmax = 5.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 2.8e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 7.476e-9
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -7.916e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25000000.0
+ tnoib = 0.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.23e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-4.377462396e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -4.986431764e-08 wvth0 = -2.627599083e-08 pvth0 = 5.271527369e-13
+ k1 = 0.64774
+ k2 = -3.569000014e-02 lk2 = -5.846003382e-08 wk2 = -3.185458373e-08 pk2 = 2.310027841e-13
+ k3 = 3.39
+ dvt0 = 2.4422
+ dvt1 = 0.16136
+ dvt2 = 0.026237
+ dvt0w = 0.5
+ dvt1w = 1928100.0
+ dvt2w = -0.032
+ w0 = 1.0e-8
+ k3b = 1.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 123760.0
+ ua = -3.152665434e-09 lua = 3.574538789e-16 wua = 9.669269988e-16 pua = -1.781924744e-21
+ ub = 3.070076680e-18 wub = -5.208212647e-25
+ uc = 3.055610254e-11 wuc = 9.066754188e-17
+ rdsw = 484.7
+ prwb = 0.1
+ prwg = 0.052
+ wr = 1.0
+ u0 = 1.895562740e-03 lu0 = 2.017615381e-09 wu0 = 2.878504968e-09 pu0 = -9.077956212e-15
+ a0 = 1.878579084e+00 la0 = -6.444115598e-07 wa0 = -3.308372593e-07 pa0 = 2.734066533e-12
+ keta = -0.01258
+ a1 = 0.0
+ a2 = 0.46703705
+ ags = 3.328546013e-01 lags = 3.807634097e-07 wags = -4.694720081e-09 pags = -2.539242761e-13
+ b0 = 0.0
+ b1 = 2.1073e-24
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.1819+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))}
+ nfactor = {3.624284492e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 3.632333127e-07 wnfactor = 4.943295571e-06 pnfactor = -2.145437392e-11
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -6.393105e-11
+ cdsc = 2.8125e-7
+ cdscb = 1.0e-4
+ cdscd = 1.0e-10
+ eta0 = 0.2
+ etab = -0.00025
+ dsub = 1.0
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.030097
+ pdiblc1 = 0.0
+ pdiblc2 = -1.497520522e-03 lpdiblc2 = 1.791849461e-08 wpdiblc2 = 8.242314363e-09 ppdiblc2 = -3.000761269e-14
+ pdiblcb = -0.025
+ drout = 0.43496
+ pscbe1 = 800000000.0
+ pscbe2 = 8.6797e-9
+ pvag = 0.0
+ delta = 1.181842103e-02 ldelta = 1.161794385e-08 wdelta = 5.878226883e-09 pdelta = 1.294865314e-13
+ alpha0 = 5.0449517e-13
+ alpha1 = -4.0583656e-18
+ beta0 = 6.2016506
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -1.706598571e+00 lkt1 = 2.777700826e-06 wkt1 = 1.739755564e-06 pkt1 = -6.849124742e-12
+ kt2 = -0.055045
+ at = 3.077022352e+05 lat = -1.425690643e-01 wat = -4.252874665e-02 pat = 1.698768256e-7
+ ute = -1.063709255e-01 lute = -1.062872873e-07 wute = -1.026637996e-06 pute = 4.100802812e-12
+ ua1 = 6.682694880e-10 lua1 = 1.111262531e-16
+ ub1 = -1.709179279e-19 lub1 = 1.958770991e-25 wub1 = -2.215658479e-26 pub1 = 8.850226230e-32
+ uc1 = -9.961e-12
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+41
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 1.4472e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 2.0e-11
+ cgso = 2.0e-11
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 0.0
+ cgdl = 0.0
+ cf = 0.0
+ clc = 7.0e-8
+ cle = 0.492
+ dlc = -1.2e-8
+ dwc = 0.0
+ vfbcv = -1.0
+ acde = 0.44
+ moin = 8.7
+ noff = 2.6123
+ voffcv = 0.112
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007653568198
+ mjs = 0.3362
+ pbs = 0.6587
+ cjsws = 9.1602368e-11
+ mjsws = 0.2659
+ pbsws = 0.7418
+ cjswgs = 2.39155046e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.19 pmos
* DC IV MOS Parameters
+ lmin = 2e-06 lmax = 4e-06 wmin = 3.0e-06 wmax = 5.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 2.8e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 7.476e-9
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -7.916e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25000000.0
+ tnoib = 0.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.23e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-4.446857209e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -2.214525354e-08 wvth0 = 7.259127622e-08 pvth0 = 1.322373254e-13
+ k1 = 0.64774
+ k2 = -5.331628715e-02 lk2 = 1.194640699e-08 wk2 = 4.926308614e-08 pk2 = -9.301363641e-14
+ k3 = 3.39
+ dvt0 = 2.4422
+ dvt1 = 0.16136
+ dvt2 = 0.026237
+ dvt0w = 0.5
+ dvt1w = 1928100.0
+ dvt2w = -0.032
+ w0 = 1.0e-8
+ k3b = 1.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 123760.0
+ ua = -2.916032420e-09 lua = -5.877530322e-16 wua = 8.158858559e-17 pua = 1.754471013e-21
+ ub = 2.775291051e-18 lub = 1.177491717e-24 wub = 3.591279877e-25 pub = -3.514869294e-30
+ uc = -2.128076763e-12 luc = 1.305536858e-16 wuc = 2.172511354e-16 puc = -5.056255061e-22
+ rdsw = 484.7
+ prwb = 0.1
+ prwg = 0.052
+ wr = 1.0
+ u0 = 2.369411897e-03 lu0 = 1.248723090e-10 wu0 = 7.079335152e-10 pu0 = -4.078256016e-16
+ a0 = 1.434169437e+00 la0 = 1.130738336e-06 wa0 = 1.890677495e-06 pa0 = -6.139552002e-12
+ keta = -0.01258
+ a1 = 0.0
+ a2 = 0.46703705
+ ags = 2.308081771e-01 lags = 7.883776463e-07 wags = 4.751743611e-07 pags = -2.170713334e-12
+ b0 = 0.0
+ b1 = 2.1073e-24
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.1819+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))}
+ nfactor = {4.383396073e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -2.668961986e-06 wnfactor = -2.619922921e-07 pnfactor = -6.623720802e-13
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -6.393105e-11
+ cdsc = 2.8125e-7
+ cdscb = 1.0e-4
+ cdscd = 1.0e-10
+ eta0 = 0.2
+ etab = -0.00025
+ dsub = 1.0
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.030097
+ pdiblc1 = 0.0
+ pdiblc2 = -1.467300553e-03 lpdiblc2 = 1.779778396e-08 wpdiblc2 = 4.406983594e-09 ppdiblc2 = -1.468776747e-14
+ pdiblcb = -0.025
+ drout = 0.43496
+ pscbe1 = 800000000.0
+ pscbe2 = 8.6797e-9
+ pvag = 0.0
+ delta = 1.266017464e-02 ldelta = 8.255643234e-09 wdelta = 7.422825020e-09 pdelta = 1.233167886e-13
+ alpha0 = 5.0449517e-13
+ alpha1 = -4.0583656e-18
+ beta0 = 6.2016506
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -1.036457736e+00 lkt1 = 1.008902747e-07 wkt1 = -8.295367301e-08 pkt1 = 4.315050330e-13
+ kt2 = -0.055045
+ at = 2.853630531e+05 lat = -5.333743550e-02 wat = 5.512666901e-02 pat = -2.201979667e-7
+ ute = -0.13298
+ ua1 = 6.9609e-10
+ ub1 = -1.2188e-19
+ uc1 = -9.961e-12
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+41
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 1.4472e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 2.0e-11
+ cgso = 2.0e-11
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 0.0
+ cgdl = 0.0
+ cf = 0.0
+ clc = 7.0e-8
+ cle = 0.492
+ dlc = -1.2e-8
+ dwc = 0.0
+ vfbcv = -1.0
+ acde = 0.44
+ moin = 8.7
+ noff = 2.6123
+ voffcv = 0.112
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007653568198
+ mjs = 0.3362
+ pbs = 0.6587
+ cjsws = 9.1602368e-11
+ mjsws = 0.2659
+ pbsws = 0.7418
+ cjswgs = 2.39155046e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.20 pmos
* DC IV MOS Parameters
+ lmin = 1.5e-06 lmax = 2e-06 wmin = 3.0e-06 wmax = 5.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 2.8e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 7.476e-9
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -7.916e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25000000.0
+ tnoib = 0.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.23e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-4.365235225e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -3.842394188e-08 wvth0 = 1.509038842e-07 pvth0 = -2.394933989e-14
+ k1 = 0.64774
+ k2 = -5.033887716e-02 lk2 = 6.008260522e-09 wk2 = 4.018208708e-08 pk2 = -7.490249188e-14
+ k3 = 3.39
+ dvt0 = 2.4422
+ dvt1 = 0.16136
+ dvt2 = 0.026237
+ dvt0w = 0.5
+ dvt1w = 1928100.0
+ dvt2w = -0.032
+ w0 = 1.0e-8
+ k3b = 1.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 5.199177925e+05 lvsat = -7.900971013e-01 wvsat = -1.182550026e+00 pvsat = 2.358477772e-6
+ ua = -3.003633671e-09 lua = -4.130410963e-16 wua = 3.430825262e-16 pua = 1.232947498e-21
+ ub = 2.892636887e-18 lub = 9.434571803e-25 wub = 8.845033135e-27 pub = -2.816264969e-30
+ uc = -3.342407414e-11 luc = 1.929704230e-16 wuc = 2.525502073e-16 puc = -5.760259751e-22
+ rdsw = 484.7
+ prwb = 0.1
+ prwg = 0.052
+ wr = 1.0
+ u0 = 1.914892719e-03 lu0 = 1.031365357e-09 wu0 = 1.803812880e-09 pu0 = -2.593447407e-15
+ a0 = 1.909251612e+00 la0 = 1.832344456e-07 wa0 = -2.450447622e-07 pa0 = -1.880067532e-12
+ keta = -0.01258
+ a1 = 0.0
+ a2 = 0.46703705
+ ags = -1.030969534e-01 lags = 1.454318039e-06 wags = 9.550087750e-07 pags = -3.127695089e-12
+ b0 = 0.0
+ b1 = 2.1073e-24
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.1819+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))}
+ nfactor = {4.783503782e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -3.466936801e-06 wnfactor = -7.743045456e-06 pnfactor = 1.425784035e-11
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -6.393105e-11
+ cdsc = 2.8125e-7
+ cdscb = 1.0e-4
+ cdscd = 1.0e-10
+ eta0 = 0.2
+ etab = -0.00025
+ dsub = 1.0
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.030097
+ pdiblc1 = 0.0
+ pdiblc2 = -7.423973215e-03 lpdiblc2 = 2.967777192e-08 wpdiblc2 = 2.761692791e-08 ppdiblc2 = -6.097768041e-14
+ pdiblcb = -0.025
+ drout = 0.43496
+ pscbe1 = 800000000.0
+ pscbe2 = 8.6797e-9
+ pvag = 0.0
+ delta = -1.440346889e-02 ldelta = 6.223137389e-08 wdelta = 2.031245788e-07 pdelta = -2.669907892e-13
+ alpha0 = 5.0449517e-13
+ alpha1 = -4.0583656e-18
+ beta0 = 6.2016506
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -1.054327956e+00 lkt1 = 1.365306412e-07 wkt1 = 3.282058471e-07 pkt1 = -3.885115138e-13
+ kt2 = 9.668213828e-02 lkt2 = -3.026046046e-07 wkt2 = -4.529127907e-07 pkt2 = 9.032892697e-13
+ at = 1.110114556e+06 lat = -1.698221833e+00 wat = -2.404237026e+00 pat = 4.684756987e-6
+ ute = -0.13298
+ ua1 = 9.090011608e-10 lua1 = -4.246300191e-16 wua1 = -6.355500347e-16 pua1 = 1.267540989e-21
+ ub1 = -9.483448068e-19 lub1 = 1.648301411e-24 wub1 = 2.467037119e-24 pub1 = -4.920258829e-30
+ uc1 = -9.961e-12
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+41
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 1.4472e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 2.0e-11
+ cgso = 2.0e-11
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 0.0
+ cgdl = 0.0
+ cf = 0.0
+ clc = 7.0e-8
+ cle = 0.492
+ dlc = -1.2e-8
+ dwc = 0.0
+ vfbcv = -1.0
+ acde = 0.44
+ moin = 8.7
+ noff = 2.6123
+ voffcv = 0.112
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007653568198
+ mjs = 0.3362
+ pbs = 0.6587
+ cjsws = 9.1602368e-11
+ mjsws = 0.2659
+ pbsws = 0.7418
+ cjswgs = 2.39155046e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.21 pmos
* DC IV MOS Parameters
+ lmin = 1e-06 lmax = 1.5e-06 wmin = 3.0e-06 wmax = 5.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 2.8e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 7.476e-9
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -7.916e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25000000.0
+ tnoib = 0.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.23e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-5.539146859e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 1.370054127e-07 wvth0 = 6.252447616e-07 pvth0 = -7.328043472e-13
+ k1 = 0.64774
+ k2 = -6.256346140e-02 lk2 = 2.427667921e-08 wk2 = 7.018113864e-08 pk2 = -1.197330745e-13
+ k3 = 3.39
+ dvt0 = 2.4422
+ dvt1 = 0.16136
+ dvt2 = 0.026237
+ dvt0w = 0.5
+ dvt1w = 1928100.0
+ dvt2w = -0.032
+ w0 = 1.0e-8
+ k3b = 1.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = -2.950518845e+05 lvsat = 4.277935839e-01 wvsat = 1.250173578e+00 pvsat = -1.276984382e-6
+ ua = -3.161590542e-09 lua = -1.769903496e-16 wua = 1.811493738e-16 pua = 1.474940401e-21
+ ub = 3.631122076e-18 lub = -1.601350853e-25 wub = -2.409882253e-24 pub = 7.982810867e-31
+ uc = 1.588360267e-10 luc = -9.434307180e-17 wuc = -5.153121542e-16 puc = 5.714675381e-22
+ rdsw = 484.7
+ prwb = 0.1
+ prwg = 0.052
+ wr = 1.0
+ u0 = 4.130860645e-03 lu0 = -2.280177112e-09 wu0 = -9.954699231e-09 pu0 = 1.497847309e-14
+ a0 = 1.123363260e+00 la0 = 1.357666000e-06 wa0 = 5.206053863e-06 pa0 = -1.002618932e-11
+ keta = -0.01258
+ a1 = 0.0
+ a2 = 0.46703705
+ ags = -1.106845905e-01 lags = 1.465657003e-06 wags = 4.063263237e-06 pags = -7.772670558e-12
+ b0 = 0.0
+ b1 = 2.1073e-24
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.1819+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))}
+ nfactor = {5.198205985e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -4.086667773e-06 wnfactor = -8.138437163e-06 pnfactor = 1.484871372e-11
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -6.393105e-11
+ cdsc = 2.8125e-7
+ cdscb = 1.0e-4
+ cdscd = 1.0e-10
+ eta0 = 0.2
+ etab = -0.00025
+ dsub = 1.0
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.030097
+ pdiblc1 = 0.0
+ pdiblc2 = -1.483574667e-02 lpdiblc2 = 4.075392618e-08 wpdiblc2 = 4.334727888e-08 ppdiblc2 = -8.448511689e-14
+ pdiblcb = -0.025
+ drout = 0.43496
+ pscbe1 = 800000000.0
+ pscbe2 = 8.6797e-9
+ pvag = 0.0
+ delta = 3.774569402e-02 ldelta = -1.570033516e-08 wdelta = -1.276670774e-07 pdelta = 2.273442618e-13
+ alpha0 = 5.0449517e-13
+ alpha1 = -4.0583656e-18
+ beta0 = 6.2016506
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -1.369243615e+00 lkt1 = 6.071406028e-07 wkt1 = 1.527830906e-06 pkt1 = -2.181231202e-12
+ kt2 = -2.450883591e-01 lkt2 = 2.081372267e-07 wkt2 = 4.529127907e-07 pkt2 = -4.503764790e-13
+ at = -6.458038851e+05 lat = 9.258226854e-01 wat = 2.772365996e+00 pat = -3.051158569e-6
+ ute = -6.691962966e-01 lute = 8.013216337e-07 wute = 3.042172006e-06 pute = -4.546221845e-12
+ ua1 = 5.918468712e-10 lua1 = 4.932535128e-17 wua1 = 6.355500347e-16 pua1 = -6.319909545e-22
+ ub1 = 4.839473348e-19 lub1 = -4.921159657e-25 wub1 = -2.467037119e-24 pub1 = 2.453221711e-30
+ uc1 = -9.961e-12
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+41
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 1.4472e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 2.0e-11
+ cgso = 2.0e-11
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 0.0
+ cgdl = 0.0
+ cf = 0.0
+ clc = 7.0e-8
+ cle = 0.492
+ dlc = -1.2e-8
+ dwc = 0.0
+ vfbcv = -1.0
+ acde = 0.44
+ moin = 8.7
+ noff = 2.6123
+ voffcv = 0.112
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007653568198
+ mjs = 0.3362
+ pbs = 0.6587
+ cjsws = 9.1602368e-11
+ mjsws = 0.2659
+ pbsws = 0.7418
+ cjswgs = 2.39155046e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 2.74e-6
+ sbref = 2.74e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.22 pmos
* DC IV MOS Parameters
+ lmin = 5e-07 lmax = 1e-06 wmin = 3.0e-06 wmax = 5.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 2.8e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 7.476e-9
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -7.916e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25000000.0
+ tnoib = 0.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.23e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope2/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-3.592433361e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -5.657577757e-08 wvth0 = -3.755957132e-07 pvth0 = 2.624314210e-13
+ k1 = 0.64774
+ k2 = -2.313517308e-02 lk2 = -1.493081070e-08 wk2 = -1.097475078e-07 pk2 = 5.918797152e-14
+ k3 = 3.39
+ dvt0 = 2.4422
+ dvt1 = 0.16136
+ dvt2 = 0.026237
+ dvt0w = 0.5
+ dvt1w = 1928100.0
+ dvt2w = -0.032
+ w0 = 1.0e-8
+ k3b = 1.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 1.467496214e+04 lvsat = 1.198012077e-01 wvsat = 3.490150363e-01 pvsat = -3.808723281e-7
+ ua = -3.860260525e-09 lua = 5.177670821e-16 wua = 3.307207888e-15 pua = -1.633612185e-21
+ ub = 4.002440454e-18 lub = -5.293740804e-25 wub = -3.196211651e-24 pub = 1.580207040e-30
+ uc = 7.475688874e-11 luc = -1.073477697e-17 wuc = 8.348977963e-17 puc = -2.398110499e-23
+ rdsw = 484.7
+ prwb = 0.1
+ prwg = 0.052
+ wr = 1.0
+ u0 = 2.268095256e-04 lu0 = 1.602011322e-09 wu0 = 1.109028592e-08 pu0 = -5.948660139e-15
+ a0 = 3.054728792e+00 la0 = -5.628838859e-07 wa0 = -8.680653301e-06 pa0 = 3.782752286e-12
+ keta = -0.01258
+ a1 = 0.0
+ a2 = 0.46703705
+ ags = 2.322695764e+00 lags = -9.540964206e-07 wags = -7.207564853e-06 pags = 3.435040895e-12
+ b0 = 1.436664019e-06 lb0 = -1.428618701e-12 wb0 = -1.046161472e-12 pb0 = 1.040302968e-18
+ b1 = 2.1073e-24
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.1819+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))}
+ nfactor = {-1.206471899e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 2.282143915e-06 wnfactor = 1.364457053e-05 pnfactor = -6.812309128e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -6.393105e-11
+ cdsc = 2.8125e-7
+ cdscb = 1.0e-4
+ cdscd = 1.0e-10
+ eta0 = 0.2
+ etab = -0.00025
+ dsub = 1.0
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.030097
+ pdiblc1 = 0.0
+ pdiblc2 = -9.804184284e-03 lpdiblc2 = 3.575054054e-08 wpdiblc2 = -2.694381612e-08 ppdiblc2 = -1.458765203e-14
+ pdiblcb = -0.025
+ drout = 0.43496
+ pscbe1 = 800000000.0
+ pscbe2 = 8.6797e-9
+ pvag = 0.0
+ delta = 2.953963187e-03 ldelta = 1.889656198e-08 wdelta = 1.263243228e-07 pdelta = -2.522478645e-14
+ alpha0 = 5.0449517e-13
+ alpha1 = -4.0583656e-18
+ beta0 = 6.2016506
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -6.643157576e-01 lkt1 = -9.383965868e-08 wkt1 = -1.160661081e-06 pkt1 = 4.922052299e-13
+ kt2 = -8.330096427e-03 lkt2 = -2.729518971e-08 wkt2 = -3.708649776e-08 pkt2 = 3.687881337e-14
+ at = 5.138530430e+05 lat = -2.273401638e-01 wat = -6.148264673e-01 pat = 3.170656163e-7
+ ute = 6.128402314e-01 lute = -4.735354898e-07 wute = -2.778350976e-06 pute = 1.241706208e-12
+ ua1 = 3.894048800e-10 lua1 = 2.506336673e-16
+ ub1 = 5.176959761e-19 lub1 = -5.256756146e-25 wub1 = 2.644831570e-25 pub1 = -2.630020513e-31
+ uc1 = -2.284941472e-11 luc1 = 1.281623960e-17 wuc1 = 2.465190329e-32 puc1 = 1.175494351e-38
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+41
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 1.4472e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 2.0e-11
+ cgso = 2.0e-11
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 0.0
+ cgdl = 0.0
+ cf = 0.0
+ clc = 7.0e-8
+ cle = 0.492
+ dlc = -1.2e-8
+ dwc = 0.0
+ vfbcv = -1.0
+ acde = 0.44
+ moin = 8.7
+ noff = 2.6123
+ voffcv = 0.112
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007653568198
+ mjs = 0.3362
+ pbs = 0.6587
+ cjsws = 9.1602368e-11
+ mjsws = 0.2659
+ pbsws = 0.7418
+ cjswgs = 2.39155046e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 1.74e-6
+ sbref = 1.74e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.23 pmos
* DC IV MOS Parameters
+ lmin = 3.5e-07 lmax = 5e-07 wmin = 3.0e-06 wmax = 5.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 2.8e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 7.476e-9
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -7.916e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25000000.0
+ tnoib = 0.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.23e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope3/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-3.797897142e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope1/sqrt(l*w*mult))} lvth0 = -4.641764822e-08 wvth0 = -2.298713995e-07 pvth0 = 1.903853203e-13
+ k1 = 0.64774
+ k2 = -3.815933590e-02 lk2 = -7.502864603e-09 wk2 = -1.237645130e-07 pk2 = 6.611797889e-14
+ k3 = 3.39
+ dvt0 = 2.4422
+ dvt1 = 0.16136
+ dvt2 = 0.026237
+ dvt0w = 0.5
+ dvt1w = 1928100.0
+ dvt2w = -0.032
+ w0 = 1.0e-8
+ k3b = 1.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 6.669693164e+05 lvsat = -2.026931211e-01 wvsat = -1.712072803e+00 pvsat = 6.381294998e-7
+ ua = -2.883571214e-09 lua = 3.489188677e-17 wua = 1.173157339e-15 pua = -5.785375939e-22
+ ub = 2.725739067e-18 lub = 1.018270854e-25 wub = -1.609212711e-24 pub = 7.955947642e-31
+ uc = -1.338483519e-11 luc = 3.284249134e-17 wuc = 3.309291173e-16 puc = -1.463151135e-22
+ rdsw = 484.7
+ prwb = 0.1
+ prwg = 0.052
+ wr = 1.0
+ u0 = 2.374327408e-03 lu0 = 5.402784810e-10 wu0 = 1.968045586e-09 pu0 = -1.438624520e-15
+ a0 = 5.712683402e+00 la0 = -1.876976645e-06 wa0 = -1.183205582e-05 pa0 = 5.340805693e-12
+ keta = -0.01258
+ a1 = 0.0
+ a2 = 0.46703705
+ ags = -1.142113310e-01 lags = 2.507104469e-07 wags = 1.254052488e-06 pags = -7.483827182e-13
+ b0 = -4.788880065e-06 lb0 = 1.649290294e-12 wb0 = 3.487204908e-12 pb0 = -1.200993370e-18
+ b1 = 2.1073e-24
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {3.865527657e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = -2.810430474e-07 wvoff = -8.592717553e-07 pvoff = 4.248239558e-13
+ nfactor = {4.066283568e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -3.247063882e-07 wnfactor = -1.037354295e-05 pnfactor = 5.062246176e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -6.393105e-11
+ cdsc = 2.8125e-7
+ cdscb = 1.0e-4
+ cdscd = 1.0e-10
+ eta0 = 0.2
+ etab = -0.00025
+ dsub = 1.0
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.030097
+ pdiblc1 = 0.0
+ pdiblc2 = -3.097773221e-02 lpdiblc2 = 4.621874263e-08 wpdiblc2 = -1.484241202e-07 ppdiblc2 = 4.547221030e-14
+ pdiblcb = -0.025
+ drout = 0.43496
+ pscbe1 = 800000000.0
+ pscbe2 = 8.6797e-9
+ pvag = 0.0
+ delta = 5.923589745e-02 ldelta = -8.929226321e-09 wdelta = -1.242424782e-07 pdelta = 9.865543992e-14
+ alpha0 = 5.0449517e-13
+ alpha1 = -4.0583656e-18
+ beta0 = 6.2016506
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -1.016307545e+00 lkt1 = 8.018508107e-08 wkt1 = -1.394759347e-07 pkt1 = -1.266870644e-14
+ kt2 = -8.081348924e-02 lkt2 = 8.540599695e-09 wkt2 = 1.236216592e-07 pkt2 = -4.257529943e-14
+ at = 1.201648976e+05 lat = -3.270074473e-02 wat = 8.730273890e-02 pat = -3.006706328e-8
+ ute = -2.220717825e-01 lute = -6.075499010e-08 wute = -8.794034317e-07 pute = 3.028665419e-13
+ ua1 = 8.9635e-10
+ ub1 = -4.223690402e-19 lub1 = -6.090747055e-26 wub1 = -8.816105234e-25 pub1 = 3.036266643e-31
+ uc1 = 3.0734e-12
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+41
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 1.4472e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 2.0e-11
+ cgso = 2.0e-11
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 0.0
+ cgdl = 0.0
+ cf = 0.0
+ clc = 7.0e-8
+ cle = 0.492
+ dlc = -1.2e-8
+ dwc = 0.0
+ vfbcv = -1.0
+ acde = 0.44
+ moin = 8.7
+ noff = 2.6123
+ voffcv = 0.112
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007653568198
+ mjs = 0.3362
+ pbs = 0.6587
+ cjsws = 9.1602368e-11
+ mjsws = 0.2659
+ pbsws = 0.7418
+ cjswgs = 2.39155046e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 1.44e-6
+ sbref = 1.44e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.24 pmos
* DC IV MOS Parameters
+ lmin = 2.0e-05 lmax = 1.0e-04 wmin = 1e-06 wmax = 3.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 2.8e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 7.476e-9
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -7.916e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25000000.0
+ tnoib = 0.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.23e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-4.478565212e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} wvth0 = 5.122497951e-8
+ k1 = 0.64774
+ k2 = -4.916126480e-02 wk2 = 1.542483196e-8
+ k3 = 3.39
+ dvt0 = 2.4422
+ dvt1 = 0.16136
+ dvt2 = 0.026237
+ dvt0w = 0.5
+ dvt1w = 1928100.0
+ dvt2w = -0.032
+ w0 = 1.0e-8
+ k3b = 1.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 123760.0
+ ua = -2.845106338e-09 wua = -4.057773476e-17
+ ub = 2.873731934e-18 wub = 6.527722548e-26
+ uc = 5.912933226e-11 wuc = 5.375079648e-18
+ rdsw = 484.7
+ prwb = 0.1
+ prwg = 0.052
+ wr = 1.0
+ u0 = 2.826979137e-03 wu0 = -2.839948914e-10
+ a0 = 1.946068784e+00 wa0 = -4.309179007e-7
+ keta = -0.01258
+ a1 = 0.0
+ a2 = 0.46703705
+ ags = 4.115234577e-01 wags = -1.291136473e-7
+ b0 = 0.0
+ b1 = 2.1073e-24
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.1819+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))}
+ nfactor = {4.035734449e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} wnfactor = 1.167050937e-6
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -6.393105e-11
+ cdsc = 2.8125e-7
+ cdscb = 1.0e-4
+ cdscd = 1.0e-10
+ eta0 = 0.2
+ etab = -0.00025
+ dsub = 1.0
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.030097
+ pdiblc1 = 0.0
+ pdiblc2 = 2.668905030e-03 wpdiblc2 = -1.257615736e-9
+ pdiblcb = -0.025
+ drout = 0.43496
+ pscbe1 = 800000000.0
+ pscbe2 = 8.6797e-9
+ pvag = 0.0
+ delta = 2.448898624e-02 wdelta = -1.140881238e-8
+ alpha0 = 5.0449517e-13
+ alpha1 = -4.0583656e-18
+ beta0 = 6.2016506
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -9.727942383e-01 wkt1 = -2.702535943e-7
+ kt2 = -0.055045
+ at = 2.869166035e+05 wat = -1.246736198e-2
+ ute = -0.29175
+ ua1 = 6.8217e-10
+ ub1 = -1.5013e-19
+ uc1 = -9.961e-12
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+41
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 1.4472e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 2.0e-11
+ cgso = 2.0e-11
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 0.0
+ cgdl = 0.0
+ cf = 0.0
+ clc = 7.0e-8
+ cle = 0.492
+ dlc = -1.2e-8
+ dwc = 0.0
+ vfbcv = -1.0
+ acde = 0.44
+ moin = 8.7
+ noff = 2.6123
+ voffcv = 0.112
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007653568198
+ mjs = 0.3362
+ pbs = 0.6587
+ cjsws = 9.1602368e-11
+ mjsws = 0.2659
+ pbsws = 0.7418
+ cjswgs = 2.39155046e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.25 pmos
* DC IV MOS Parameters
+ lmin = 8e-06 lmax = 2.0e-05 wmin = 1e-06 wmax = 3.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 2.8e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 7.476e-9
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -7.916e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25000000.0
+ tnoib = 0.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.23e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-4.478565212e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} wvth0 = 5.122497951e-8
+ k1 = 0.64774
+ k2 = -4.916126480e-02 wk2 = 1.542483196e-8
+ k3 = 3.39
+ dvt0 = 2.4422
+ dvt1 = 0.16136
+ dvt2 = 0.026237
+ dvt0w = 0.5
+ dvt1w = 1928100.0
+ dvt2w = -0.032
+ w0 = 1.0e-8
+ k3b = 1.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 123760.0
+ ua = -2.845106338e-09 wua = -4.057773476e-17
+ ub = 2.873731934e-18 wub = 6.527722548e-26
+ uc = 5.912933226e-11 wuc = 5.375079648e-18
+ rdsw = 484.7
+ prwb = 0.1
+ prwg = 0.052
+ wr = 1.0
+ u0 = 2.826979137e-03 wu0 = -2.839948914e-10
+ a0 = 1.946068784e+00 wa0 = -4.309179007e-7
+ keta = -0.01258
+ a1 = 0.0
+ a2 = 0.46703705
+ ags = 4.115234577e-01 wags = -1.291136473e-7
+ b0 = 0.0
+ b1 = 2.1073e-24
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.1819+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))}
+ nfactor = {4.035734449e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} wnfactor = 1.167050937e-6
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -6.393105e-11
+ cdsc = 2.8125e-7
+ cdscb = 1.0e-4
+ cdscd = 1.0e-10
+ eta0 = 0.2
+ etab = -0.00025
+ dsub = 1.0
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.030097
+ pdiblc1 = 0.0
+ pdiblc2 = 2.668905030e-03 wpdiblc2 = -1.257615736e-9
+ pdiblcb = -0.025
+ drout = 0.43496
+ pscbe1 = 800000000.0
+ pscbe2 = 8.6797e-9
+ pvag = 0.0
+ delta = 2.448898624e-02 wdelta = -1.140881238e-8
+ alpha0 = 5.0449517e-13
+ alpha1 = -4.0583656e-18
+ beta0 = 6.2016506
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -9.727942383e-01 wkt1 = -2.702535943e-7
+ kt2 = -0.055045
+ at = 2.869166035e+05 wat = -1.246736198e-2
+ ute = -0.29175
+ ua1 = 6.8217e-10
+ ub1 = -1.5013e-19
+ uc1 = -9.961e-12
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+41
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 1.4472e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 2.0e-11
+ cgso = 2.0e-11
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 0.0
+ cgdl = 0.0
+ cf = 0.0
+ clc = 7.0e-8
+ cle = 0.492
+ dlc = -1.2e-8
+ dwc = 0.0
+ vfbcv = -1.0
+ acde = 0.44
+ moin = 8.7
+ noff = 2.6123
+ voffcv = 0.112
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007653568198
+ mjs = 0.3362
+ pbs = 0.6587
+ cjsws = 9.1602368e-11
+ mjsws = 0.2659
+ pbsws = 0.7418
+ cjswgs = 2.39155046e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.26 pmos
* DC IV MOS Parameters
+ lmin = 4e-06 lmax = 8e-06 wmin = 1e-06 wmax = 3.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 2.8e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 7.476e-9
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -7.916e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25000000.0
+ tnoib = 0.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.23e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-4.651056143e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 1.378961495e-07 wvth0 = 5.539305591e-08 pvth0 = -3.332126999e-14
+ k1 = 0.64774
+ k2 = -5.229020380e-02 lk2 = 2.501398995e-08 wk2 = 1.769782100e-08 pk2 = -1.817118359e-14
+ k3 = 3.39
+ dvt0 = 2.4422
+ dvt1 = 0.16136
+ dvt2 = 0.026237
+ dvt0w = 0.5
+ dvt1w = 1928100.0
+ dvt2w = -0.032
+ w0 = 1.0e-8
+ k3b = 1.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 123760.0
+ ua = -2.824985027e-09 lua = -1.608578060e-16 wua = -1.121474495e-17 pua = -2.347394857e-22
+ ub = 2.914554195e-18 lub = -3.263494810e-25 wub = -5.657918221e-26 pub = 9.741688656e-31
+ uc = 5.912933226e-11 wuc = 5.375079648e-18
+ rdsw = 484.7
+ prwb = 0.1
+ prwg = 0.052
+ wr = 1.0
+ u0 = 3.023006004e-03 lu0 = -1.567117185e-09 wu0 = -4.869672925e-10 pu0 = 1.622642563e-15
+ a0 = 1.942108301e+00 la0 = 3.166168969e-08 wa0 = -5.204750196e-07 pa0 = 7.159554314e-13
+ keta = -0.01258
+ a1 = 0.0
+ a2 = 0.46703705
+ ags = 3.806134040e-01 lags = 2.471073330e-07 wags = -1.472570387e-07 pags = 1.450455282e-13
+ b0 = 0.0
+ b1 = 2.1073e-24
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.1819+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))}
+ nfactor = {5.207603812e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -9.368392437e-06 wnfactor = 2.170114015e-07 pnfactor = 7.594996060e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -6.393105e-11
+ cdsc = 2.8125e-7
+ cdscb = 1.0e-4
+ cdscd = 1.0e-10
+ eta0 = 0.2
+ etab = -0.00025
+ dsub = 1.0
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.030097
+ pdiblc1 = 0.0
+ pdiblc2 = 2.767954761e-03 lpdiblc2 = -7.918431740e-10 wpdiblc2 = -4.490334099e-09 ppdiblc2 = 2.584364368e-14
+ pdiblcb = -0.025
+ drout = 0.43496
+ pscbe1 = 800000000.0
+ pscbe2 = 8.6797e-9
+ pvag = 0.0
+ delta = 1.901431008e-02 ldelta = 4.376675113e-08 wdelta = -1.560184733e-08 pdelta = 3.352079856e-14
+ alpha0 = 5.0449517e-13
+ alpha1 = -4.0583656e-18
+ beta0 = 6.2016506
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -9.633645737e-01 lkt1 = -7.538451101e-08 wkt1 = -4.788335924e-07 pkt1 = 1.667471937e-12
+ kt2 = -0.055045
+ at = 3.018023378e+05 lat = -1.190025141e-01 wat = -2.491726966e-02 pat = 9.952954194e-8
+ ute = -4.502977220e-01 lute = 1.267493909e-6
+ ua1 = 6.682694880e-10 lua1 = 1.111262531e-16
+ ub1 = -1.537629899e-19 lub1 = 2.904357429e-26 wub1 = -7.336489818e-26 pub1 = 5.865083420e-31
+ uc1 = -9.961e-12
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+41
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 1.4472e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 2.0e-11
+ cgso = 2.0e-11
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 0.0
+ cgdl = 0.0
+ cf = 0.0
+ clc = 7.0e-8
+ cle = 0.492
+ dlc = -1.2e-8
+ dwc = 0.0
+ vfbcv = -1.0
+ acde = 0.44
+ moin = 8.7
+ noff = 2.6123
+ voffcv = 0.112
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007653568198
+ mjs = 0.3362
+ pbs = 0.6587
+ cjsws = 9.1602368e-11
+ mjsws = 0.2659
+ pbsws = 0.7418
+ cjswgs = 2.39155046e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.27 pmos
* DC IV MOS Parameters
+ lmin = 2e-06 lmax = 4e-06 wmin = 1e-06 wmax = 3.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 2.8e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 7.476e-9
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -7.916e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25000000.0
+ tnoib = 0.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.23e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-4.430233822e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 4.969088194e-08 wvth0 = 6.762911569e-08 pvth0 = -8.219698718e-14
+ k1 = 0.64774
+ k2 = -4.255793417e-02 lk2 = -1.386058786e-08 wk2 = 1.714888611e-08 pk2 = -1.597851806e-14
+ k3 = 3.39
+ dvt0 = 2.4422
+ dvt1 = 0.16136
+ dvt2 = 0.026237
+ dvt0w = 0.5
+ dvt1w = 1928100.0
+ dvt2w = -0.032
+ w0 = 1.0e-8
+ k3b = 1.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 123760.0
+ ua = -2.840698611e-09 lua = -9.809146598e-17 wua = -1.432864504e-16 pua = 2.928077343e-22
+ ub = 2.803138174e-18 lub = 1.186906738e-25 wub = 2.760029889e-25 pub = -3.542973585e-31
+ uc = 7.363920701e-11 luc = -5.795824370e-17 wuc = -8.917843455e-18 puc = 5.709165204e-23
+ rdsw = 484.7
+ prwb = 0.1
+ prwg = 0.052
+ wr = 1.0
+ u0 = 2.692808046e-03 lu0 = -2.481744612e-10 wu0 = -2.574195131e-10 pu0 = 7.057369136e-16
+ a0 = 2.243536499e+00 la0 = -1.172363106e-06 wa0 = -5.253220353e-07 pa0 = 7.353163509e-13
+ keta = -0.01258
+ a1 = 0.0
+ a2 = 0.46703705
+ ags = 4.534420017e-01 lags = -4.379921770e-08 wags = -1.893982918e-07 pags = 3.133745496e-13
+ b0 = 0.0
+ b1 = 2.1073e-24
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.1819+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))}
+ nfactor = {3.377341142e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -2.057591227e-06 wnfactor = 2.741129968e-06 pnfactor = -2.487343142e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -6.393105e-11
+ cdsc = 2.8125e-7
+ cdscb = 1.0e-4
+ cdscd = 1.0e-10
+ eta0 = 0.2
+ etab = -0.00025
+ dsub = 1.0
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.030097
+ pdiblc1 = 0.0
+ pdiblc2 = 7.195206015e-06 lpdiblc2 = 1.023573479e-08 wpdiblc2 = 5.542977376e-12 ppdiblc2 = 7.885312286e-15
+ pdiblcb = -0.025
+ drout = 0.43496
+ pscbe1 = 800000000.0
+ pscbe2 = 8.6797e-9
+ pvag = 0.0
+ delta = 1.213994084e-02 ldelta = 7.122573161e-08 wdelta = 8.975747882e-09 pdelta = -6.465194774e-14
+ alpha0 = 5.0449517e-13
+ alpha1 = -4.0583656e-18
+ beta0 = 6.2016506
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -1.064057279e+00 lkt1 = 3.268224304e-07 wkt1 = -5.677119134e-10 pkt1 = -2.429132964e-13
+ kt2 = -0.055045
+ at = 3.038306520e+05 lat = -1.271044123e-1
+ ute = -1.434315642e-01 lute = 4.174772792e-08 wute = 3.119842072e-08 pute = -1.246189717e-13
+ ua1 = 6.9609e-10
+ ub1 = -1.710349202e-19 lub1 = 9.803457293e-26 wub1 = 1.467297964e-25 pub1 = -2.926379059e-31
+ uc1 = -9.961e-12
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+41
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 1.4472e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 2.0e-11
+ cgso = 2.0e-11
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 0.0
+ cgdl = 0.0
+ cf = 0.0
+ clc = 7.0e-8
+ cle = 0.492
+ dlc = -1.2e-8
+ dwc = 0.0
+ vfbcv = -1.0
+ acde = 0.44
+ moin = 8.7
+ noff = 2.6123
+ voffcv = 0.112
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007653568198
+ mjs = 0.3362
+ pbs = 0.6587
+ cjsws = 9.1602368e-11
+ mjsws = 0.2659
+ pbsws = 0.7418
+ cjswgs = 2.39155046e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.28 pmos
* DC IV MOS Parameters
+ lmin = 1.5e-06 lmax = 2e-06 wmin = 1e-06 wmax = 3.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 2.8e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 7.476e-9
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -7.916e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25000000.0
+ tnoib = 0.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.23e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-3.833491909e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -6.932332538e-08 wvth0 = -7.824048267e-09 pvth0 = 6.828680302e-14
+ k1 = 0.64774
+ k2 = -3.522581170e-02 lk2 = -2.848377291e-08 wk2 = -4.931138764e-09 pk2 = 2.805788354e-14
+ k3 = 3.39
+ dvt0 = 2.4422
+ dvt1 = 0.16136
+ dvt2 = 0.026237
+ dvt0w = 0.5
+ dvt1w = 1928100.0
+ dvt2w = -0.032
+ w0 = 1.0e-8
+ k3b = 1.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 123760.0
+ ua = -2.889882058e-09 wua = 3.528498675e-18
+ ub = 2.862650144e-18 wub = 9.835690056e-26
+ uc = 4.457871578e-11 wuc = 1.970813531e-17
+ rdsw = 484.7
+ prwb = 0.1
+ prwg = 0.052
+ wr = 1.0
+ u0 = 2.446724860e-03 lu0 = 2.426138454e-10 wu0 = 2.162684114e-10 pu0 = -2.389862832e-16
+ a0 = 1.989920802e+00 la0 = -6.665519585e-07 wa0 = -4.858461642e-07 pa0 = 6.565856737e-13
+ keta = -0.01258
+ a1 = 0.0
+ a2 = 0.46703705
+ ags = 1.272505409e-01 lags = 6.067570317e-07 wags = 2.674104477e-07 pags = -5.976848006e-13
+ b0 = 0.0
+ b1 = 2.1073e-24
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.1819+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))}
+ nfactor = {1.365696025e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 1.954433794e-06 wnfactor = 2.459274752e-06 pnfactor = -1.925211100e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -6.393105e-11
+ cdsc = 2.8125e-7
+ cdscb = 1.0e-4
+ cdscd = 1.0e-10
+ eta0 = 0.2
+ etab = -0.00025
+ dsub = 1.0
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.030097
+ pdiblc1 = 0.0
+ pdiblc2 = -1.782923056e-03 lpdiblc2 = 1.380594665e-08 wpdiblc2 = 1.077812241e-08 ppdiblc2 = -1.359952014e-14
+ pdiblcb = -0.025
+ drout = 0.43496
+ pscbe1 = 800000000.0
+ pscbe2 = 8.6797e-9
+ pvag = 0.0
+ delta = 6.821660907e-02 ldelta = -4.061357551e-08 wdelta = -4.350031964e-08 pdelta = 4.000632133e-14
+ alpha0 = 5.0449517e-13
+ alpha1 = -4.0583656e-18
+ beta0 = 6.2016506
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -9.049603431e-01 lkt1 = 9.519501817e-09 wkt1 = -1.176636456e-07 pkt1 = -9.377166226e-15
+ kt2 = -0.055045
+ at = 3.364990924e+05 lat = -1.922583498e-01 wat = -9.495773312e-02 pat = 1.893837029e-7
+ ute = -1.224990893e-01 wute = -3.128602158e-8
+ ua1 = 6.9609e-10
+ ub1 = -1.2188e-19
+ uc1 = -9.961e-12
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+41
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 1.4472e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 2.0e-11
+ cgso = 2.0e-11
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 0.0
+ cgdl = 0.0
+ cf = 0.0
+ clc = 7.0e-8
+ cle = 0.492
+ dlc = -1.2e-8
+ dwc = 0.0
+ vfbcv = -1.0
+ acde = 0.44
+ moin = 8.7
+ noff = 2.6123
+ voffcv = 0.112
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007653568198
+ mjs = 0.3362
+ pbs = 0.6587
+ cjsws = 9.1602368e-11
+ mjsws = 0.2659
+ pbsws = 0.7418
+ cjswgs = 2.39155046e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.29 pmos
* DC IV MOS Parameters
+ lmin = 1e-06 lmax = 1.5e-06 wmin = 1e-06 wmax = 3.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 2.8e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 7.476e-9
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -7.916e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25000000.0
+ tnoib = 0.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.23e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-2.999067500e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -1.940197090e-07 wvth0 = -1.329811195e-07 pvth0 = 2.553215302e-13
+ k1 = 0.64774
+ k2 = -3.429769272e-02 lk2 = -2.987075392e-08 wk2 = -1.419353764e-08 pk2 = 4.189961243e-14
+ k3 = 3.39
+ dvt0 = 2.4422
+ dvt1 = 0.16136
+ dvt2 = 0.026237
+ dvt0w = 0.5
+ dvt1w = 1928100.0
+ dvt2w = -0.032
+ w0 = 1.0e-8
+ k3b = 1.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 123760.0
+ ua = -3.206603053e-09 lua = 4.733078560e-16 wua = 3.155138821e-16 pua = -4.662309569e-22
+ ub = 2.755493369e-18 lub = 1.601350853e-25 wub = 2.039114679e-25 pub = -1.577407455e-31
+ uc = -5.239965021e-11 luc = 1.449244701e-16 wuc = 1.152364808e-16 puc = -1.427575595e-22
+ rdsw = 484.7
+ prwb = 0.1
+ prwg = 0.052
+ wr = 1.0
+ u0 = -1.112394704e-04 lu0 = 4.065235741e-09 wu0 = 2.708173235e-09 pu0 = -3.962888852e-15
+ a0 = 3.219306597e+00 la0 = -2.503746091e-06 wa0 = -1.050437603e-06 pa0 = 1.500311120e-12
+ keta = -0.01258
+ a1 = 0.0
+ a2 = 0.46703705
+ ags = 1.596156188e+00 lags = -1.588375568e-06 wags = -1.031738416e-06 pags = 1.343763261e-12
+ b0 = 0.0
+ b1 = 2.1073e-24
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.1819+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))}
+ nfactor = {-9.864541955e-02+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 4.142745649e-06 wnfactor = 7.672918529e-06 pnfactor = -9.716480359e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -6.393105e-11
+ cdsc = 2.8125e-7
+ cdscb = 1.0e-4
+ cdscd = 1.0e-10
+ eta0 = 0.2
+ etab = -0.00025
+ dsub = 1.0
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.030097
+ pdiblc1 = 0.0
+ pdiblc2 = 3.452987237e-03 lpdiblc2 = 5.981402313e-09 wpdiblc2 = -1.124546971e-08 ppdiblc2 = 1.931253593e-14
+ pdiblcb = -0.025
+ drout = 0.43496
+ pscbe1 = 800000000.0
+ pscbe2 = 8.6797e-9
+ pvag = 0.0
+ delta = 2.891008018e-03 ldelta = 5.700900270e-08 wdelta = -2.362416664e-08 pdelta = 1.030339828e-14
+ alpha0 = 5.0449517e-13
+ alpha1 = -4.0583656e-18
+ beta0 = 6.2016506
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -6.506881010e-01 lkt1 = -3.704649368e-07 wkt1 = -6.170917940e-07 pkt1 = 7.369682586e-13
+ kt2 = -9.336122080e-02 lkt2 = 5.725976036e-8
+ at = 2.299094310e+05 lat = -3.297075991e-02 wat = 1.583197130e-01 pat = -1.891141126e-7
+ ute = 5.937751710e-01 lute = -1.070400255e-06 wute = -7.278584479e-07 pute = 1.040957834e-12
+ ua1 = 8.047580320e-10 lua1 = -1.623935070e-16
+ ub1 = -3.425174720e-19 lub1 = 3.297206382e-25
+ uc1 = -9.961e-12
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+41
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 1.4472e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 2.0e-11
+ cgso = 2.0e-11
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 0.0
+ cgdl = 0.0
+ cf = 0.0
+ clc = 7.0e-8
+ cle = 0.492
+ dlc = -1.2e-8
+ dwc = 0.0
+ vfbcv = -1.0
+ acde = 0.44
+ moin = 8.7
+ noff = 2.6123
+ voffcv = 0.112
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007653568198
+ mjs = 0.3362
+ pbs = 0.6587
+ cjsws = 9.1602368e-11
+ mjsws = 0.2659
+ pbsws = 0.7418
+ cjswgs = 2.39155046e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 2.74e-6
+ sbref = 2.74e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.30 pmos
* DC IV MOS Parameters
+ lmin = 5e-07 lmax = 1e-06 wmin = 1e-06 wmax = 3.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 2.8e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 7.476e-9
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -7.916e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25000000.0
+ tnoib = 0.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.23e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope2/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-5.372551247e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 4.199951477e-08 wvth0 = 1.557780202e-07 pvth0 = -3.182055825e-14
+ k1 = 0.64774
+ k2 = -7.216546204e-02 lk2 = 7.784955895e-09 wk2 = 3.661025815e-08 pk2 = -8.619682112e-15
+ k3 = 3.39
+ dvt0 = 2.4422
+ dvt1 = 0.16136
+ dvt2 = 0.026237
+ dvt0w = 0.5
+ dvt1w = 1928100.0
+ dvt2w = -0.032
+ w0 = 1.0e-8
+ k3b = 1.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 1.260937315e+05 lvsat = -2.320662595e-03 wvsat = 1.642466170e-02 pvsat = -1.633268359e-8
+ ua = -2.705835824e-09 lua = -2.465507672e-17 wua = -1.388052570e-16 pua = -1.445600502e-23
+ ub = 2.955490879e-18 lub = -3.874243903e-26 wub = -7.101691666e-26 pub = 1.156480401e-31
+ uc = 1.177368754e-10 luc = -2.425929097e-17 wuc = -4.480754372e-17 puc = 1.639021849e-23
+ rdsw = 484.7
+ prwb = 0.1
+ prwg = 0.052
+ wr = 1.0
+ u0 = 4.536510405e-03 lu0 = -5.564867355e-10 wu0 = -1.774378074e-09 pu0 = 4.945601701e-16
+ a0 = -3.576855774e-01 la0 = 1.053214927e-06 wa0 = 1.505567389e-06 pa0 = -1.041380244e-12
+ keta = -0.01258
+ a1 = 0.0
+ a2 = 0.46703705
+ ags = -3.286237866e-01 lags = 3.256256393e-07 wags = 7.067512675e-07 pags = -3.849908801e-13
+ b0 = 1.567506541e-06 lb0 = -1.558728504e-12 wb0 = -1.436732679e-12 pb0 = 1.428686976e-18
+ b1 = 5.445233443e-08 lb1 = -5.414740135e-14 wb1 = -1.625428320e-13 pb1 = 1.616325921e-19
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.1819+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))}
+ nfactor = {4.294385596e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -2.256843930e-07 wnfactor = -2.775753138e-06 pnfactor = 6.736787459e-13
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -6.393105e-11
+ cdsc = 2.8125e-7
+ cdscb = 1.0e-4
+ cdscd = 1.0e-10
+ eta0 = 0.2
+ etab = -0.00025
+ dsub = 1.0
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.030097
+ pdiblc1 = 0.0
+ pdiblc2 = -2.138041016e-02 lpdiblc2 = 3.067573269e-08 wpdiblc2 = 7.611773787e-09 ppdiblc2 = 5.608929947e-16
+ pdiblcb = -0.025
+ drout = 0.43496
+ pscbe1 = 800000000.0
+ pscbe2 = 8.6797e-9
+ pvag = 0.0
+ delta = 5.188371922e-02 ldelta = 8.290650686e-09 wdelta = -1.973334761e-08 pdelta = 6.434367834e-15
+ alpha0 = 5.0449517e-13
+ alpha1 = -4.0583656e-18
+ beta0 = 6.2016506
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -1.109952835e+00 lkt1 = 8.622791464e-08 wkt1 = 1.695869856e-07 pkt1 = -4.530511973e-14
+ kt2 = -2.075418400e-02 lkt2 = -1.494067703e-8
+ at = 3.280447319e+05 lat = -1.305565031e-01 wat = -6.017973988e-02 pat = 2.816174338e-8
+ ute = -4.331209124e-01 lute = -4.925478926e-08 wute = 3.438932441e-07 pute = -2.479204861e-14
+ ua1 = 3.894048800e-10 lua1 = 2.506336673e-16
+ ub1 = 6.062986240e-19 lub1 = -6.137820877e-25 wub1 = -7.461634063e-41 pub1 = -1.094764425e-47
+ uc1 = -2.284941472e-11 luc1 = 1.281623960e-17
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+41
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 1.4472e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 2.0e-11
+ cgso = 2.0e-11
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 0.0
+ cgdl = 0.0
+ cf = 0.0
+ clc = 7.0e-8
+ cle = 0.492
+ dlc = -1.2e-8
+ dwc = 0.0
+ vfbcv = -1.0
+ acde = 0.44
+ moin = 8.7
+ noff = 2.6123
+ voffcv = 0.112
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007653568198
+ mjs = 0.3362
+ pbs = 0.6587
+ cjsws = 9.1602368e-11
+ mjsws = 0.2659
+ pbsws = 0.7418
+ cjswgs = 2.39155046e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 1.74e-6
+ sbref = 1.74e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.31 pmos
* DC IV MOS Parameters
+ lmin = 3.5e-07 lmax = 5e-07 wmin = 1e-06 wmax = 3.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 2.8e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 7.476e-9
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -7.916e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25000000.0
+ tnoib = 0.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.23e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope3/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-5.367761371e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 4.176270331e-08 wvth0 = 2.387406080e-07 pvth0 = -7.283726164e-14
+ k1 = 0.64774
+ k2 = -9.194721654e-02 lk2 = 1.756505532e-08 wk2 = 3.679489249e-08 pk2 = -8.710965330e-15
+ k3 = 3.39
+ dvt0 = 2.4422
+ dvt1 = 0.16136
+ dvt2 = 0.026237
+ dvt0w = 0.5
+ dvt1w = 1928100.0
+ dvt2w = -0.032
+ w0 = 1.0e-8
+ k3b = 1.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 8.859795159e+04 lvsat = 1.621725099e-02 wvsat = 1.439348237e-02 pvsat = -1.532846853e-8
+ ua = -2.321180996e-09 lua = -2.148284235e-16 wua = -5.056044559e-16 pua = 1.668895189e-22
+ ub = 2.016844244e-18 lub = 4.253244576e-25 wub = 5.068723631e-25 pub = -1.700604198e-31
+ uc = 1.174942768e-10 luc = -2.413935022e-17 wuc = -5.975131428e-17 puc = 2.377841866e-23
+ rdsw = 484.7
+ prwb = 0.1
+ prwg = 0.052
+ wr = 1.0
+ u0 = 3.507390567e-03 lu0 = -4.768988784e-11 wu0 = -1.414202333e-09 pu0 = 3.164892837e-16
+ a0 = 2.037631515e+00 la0 = -1.310298433e-07 wa0 = -8.618495389e-07 pa0 = 1.290706850e-13
+ keta = -1.172621950e-02 lketa = -4.221090809e-10 wketa = -2.548575784e-09 pketa = 1.260015868e-15
+ a1 = 0.0
+ a2 = 0.46703705
+ ags = 3.300041246e-01 wags = -7.195196881e-8
+ b0 = -5.423438130e-06 lb0 = 1.897594541e-12 wb0 = 5.381391191e-12 pb0 = -1.942193465e-18
+ b1 = 5.127462474e-08 lb1 = -5.257634168e-14 wb1 = -1.530572160e-13 pb1 = 1.569429036e-19
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {7.006141517e-02+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = -1.245697237e-07 wvoff = 8.547011770e-08 pvoff = -4.225642619e-14
+ nfactor = {2.443188824e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 6.895472911e-07 wnfactor = -5.528527233e-06 pnfactor = 2.034650259e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -6.393105e-11
+ cdsc = 2.8125e-7
+ cdscb = 1.0e-4
+ cdscd = 1.0e-10
+ eta0 = 0.2
+ etab = -0.00025
+ dsub = 1.0
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.030097
+ pdiblc1 = 0.0
+ pdiblc2 = -9.666541752e-02 lpdiblc2 = 6.789664033e-08 wpdiblc2 = 4.765677346e-08 ppdiblc2 = -1.923735485e-14
+ pdiblcb = -0.025
+ drout = 0.43496
+ pscbe1 = 800000000.0
+ pscbe2 = 8.6797e-9
+ pvag = 0.0
+ delta = -1.535133613e-02 ldelta = 4.153166205e-08 wdelta = 9.840399425e-08 pdelta = -5.197273398e-14
+ alpha0 = 5.0449517e-13
+ alpha1 = -4.0583656e-18
+ beta0 = 6.2016506
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -1.169220456e+00 lkt1 = 1.155298266e-07 wkt1 = 3.169764448e-07 pkt1 = -1.181744683e-13
+ kt2 = -7.256047259e-02 lkt2 = 1.067235205e-08 wkt2 = 9.898600835e-08 pkt2 = -4.893868253e-14
+ at = 1.510890536e+05 lat = -4.306961576e-02 wat = -5.007351278e-03 pat = 8.845144503e-10
+ ute = -6.305393711e-01 lute = 4.834889671e-08 wute = 3.398919266e-07 pute = -2.281379724e-14
+ ua1 = 7.005119767e-10 lua1 = 9.682231872e-17 wua1 = 5.845858998e-16 pua1 = -2.890192689e-22
+ ub1 = -3.029774256e-19 lub1 = -1.642360088e-25 wub1 = -1.238000224e-24 pub1 = 6.120673106e-31
+ uc1 = 3.352294451e-11 luc1 = -1.505425481e-17 wuc1 = -9.089335194e-17 puc1 = 4.493767320e-23
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+41
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 1.4472e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 2.0e-11
+ cgso = 2.0e-11
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 0.0
+ cgdl = 0.0
+ cf = 0.0
+ clc = 7.0e-8
+ cle = 0.492
+ dlc = -1.2e-8
+ dwc = 0.0
+ vfbcv = -1.0
+ acde = 0.44
+ moin = 8.7
+ noff = 2.6123
+ voffcv = 0.112
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007653568198
+ mjs = 0.3362
+ pbs = 0.6587
+ cjsws = 9.1602368e-11
+ mjsws = 0.2659
+ pbsws = 0.7418
+ cjswgs = 2.39155046e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 1.44e-6
+ sbref = 1.44e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.32 pmos
* DC IV MOS Parameters
+ lmin = 2.0e-05 lmax = 1.0e-04 wmin = 5.5e-07 wmax = 1.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 2.8e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 7.476e-9
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -7.916e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25000000.0
+ tnoib = 0.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.23e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-4.310444637e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} wvth0 = 3.466429585e-8
+ k1 = 0.64774
+ k2 = -4.768499569e-02 wk2 = 1.397063602e-8
+ k3 = 3.39
+ dvt0 = 2.4422
+ dvt1 = 0.16136
+ dvt2 = 0.026237
+ dvt0w = 0.5
+ dvt1w = 1928100.0
+ dvt2w = -0.032
+ w0 = 1.0e-8
+ k3b = 1.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 123760.0
+ ua = -2.714727941e-09 wua = -1.690067132e-16
+ ub = 2.777107609e-18 wub = 1.604568241e-25
+ uc = 6.996144891e-11 wuc = -5.295075195e-18
+ rdsw = 484.7
+ prwb = 0.1
+ prwg = 0.052
+ wr = 1.0
+ u0 = 2.892886571e-03 wu0 = -3.489168776e-10
+ a0 = 1.252631147e+00 wa0 = 2.521514573e-7
+ keta = -0.01258
+ a1 = 0.0
+ a2 = 0.46703705
+ ags = 2.992836896e-01 wags = -1.855208827e-8
+ b0 = 1.088133063e-07 wb0 = -1.071863297e-13
+ b1 = -3.709309435e-07 wb1 = 3.653847840e-13
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.1819+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))}
+ nfactor = {4.962725764e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} wnfactor = 2.539199961e-7
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -6.393105e-11
+ cdsc = 2.8125e-7
+ cdscb = 1.0e-4
+ cdscd = 1.0e-10
+ eta0 = 0.2
+ etab = -0.00025
+ dsub = 1.0
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.030097
+ pdiblc1 = 0.0
+ pdiblc2 = 2.532779657e-03 wpdiblc2 = -1.123525710e-9
+ pdiblcb = -0.025
+ drout = 0.43496
+ pscbe1 = 800000000.0
+ pscbe2 = 8.6797e-9
+ pvag = 0.0
+ delta = 1.211393996e-02 wdelta = 7.812022019e-10
+ alpha0 = 5.0449517e-13
+ alpha1 = -4.0583656e-18
+ beta0 = 6.2016506
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -1.376952645e+00 wkt1 = 1.278618357e-7
+ kt2 = -0.055045
+ at = 2.648074853e+05 wat = 9.311180667e-3
+ ute = -2.986818441e-01 wute = 6.828199156e-9
+ ua1 = 6.8217e-10
+ ub1 = -1.5013e-19
+ uc1 = -9.961e-12
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+41
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 1.4472e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 2.0e-11
+ cgso = 2.0e-11
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 0.0
+ cgdl = 0.0
+ cf = 0.0
+ clc = 7.0e-8
+ cle = 0.492
+ dlc = -1.2e-8
+ dwc = 0.0
+ vfbcv = -1.0
+ acde = 0.44
+ moin = 8.7
+ noff = 2.6123
+ voffcv = 0.112
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007653568198
+ mjs = 0.3362
+ pbs = 0.6587
+ cjsws = 9.1602368e-11
+ mjsws = 0.2659
+ pbsws = 0.7418
+ cjswgs = 2.39155046e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.33 pmos
* DC IV MOS Parameters
+ lmin = 8e-06 lmax = 2.0e-05 wmin = 5.5e-07 wmax = 1.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 2.8e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 7.476e-9
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -7.916e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25000000.0
+ tnoib = 0.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.23e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-4.310444637e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope1/sqrt(l*w*mult))} wvth0 = 3.466429585e-8
+ k1 = 0.64774
+ k2 = -4.768499569e-02 wk2 = 1.397063602e-8
+ k3 = 3.39
+ dvt0 = 2.4422
+ dvt1 = 0.16136
+ dvt2 = 0.026237
+ dvt0w = 0.5
+ dvt1w = 1928100.0
+ dvt2w = -0.032
+ w0 = 1.0e-8
+ k3b = 1.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 123760.0
+ ua = -2.714727941e-09 wua = -1.690067132e-16
+ ub = 2.777107609e-18 wub = 1.604568241e-25
+ uc = 6.996144891e-11 wuc = -5.295075195e-18
+ rdsw = 484.7
+ prwb = 0.1
+ prwg = 0.052
+ wr = 1.0
+ u0 = 2.892886571e-03 wu0 = -3.489168776e-10
+ a0 = 1.252631147e+00 wa0 = 2.521514573e-7
+ keta = -0.01258
+ a1 = 0.0
+ a2 = 0.46703705
+ ags = 2.992836896e-01 wags = -1.855208827e-8
+ b0 = 1.088133063e-07 wb0 = -1.071863297e-13
+ b1 = -3.709309435e-07 wb1 = 3.653847840e-13
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.1819+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))}
+ nfactor = {4.962725764e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} wnfactor = 2.539199961e-7
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -6.393105e-11
+ cdsc = 2.8125e-7
+ cdscb = 1.0e-4
+ cdscd = 1.0e-10
+ eta0 = 0.2
+ etab = -0.00025
+ dsub = 1.0
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.030097
+ pdiblc1 = 0.0
+ pdiblc2 = 2.532779657e-03 wpdiblc2 = -1.123525710e-9
+ pdiblcb = -0.025
+ drout = 0.43496
+ pscbe1 = 800000000.0
+ pscbe2 = 8.6797e-9
+ pvag = 0.0
+ delta = 1.211393996e-02 wdelta = 7.812022019e-10
+ alpha0 = 5.0449517e-13
+ alpha1 = -4.0583656e-18
+ beta0 = 6.2016506
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -1.376952645e+00 wkt1 = 1.278618357e-7
+ kt2 = -0.055045
+ at = 2.648074853e+05 wat = 9.311180667e-3
+ ute = -2.986818441e-01 wute = 6.828199156e-9
+ ua1 = 6.8217e-10
+ ub1 = -1.5013e-19
+ uc1 = -9.961e-12
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+41
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 1.4472e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 2.0e-11
+ cgso = 2.0e-11
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 0.0
+ cgdl = 0.0
+ cf = 0.0
+ clc = 7.0e-8
+ cle = 0.492
+ dlc = -1.2e-8
+ dwc = 0.0
+ vfbcv = -1.0
+ acde = 0.44
+ moin = 8.7
+ noff = 2.6123
+ voffcv = 0.112
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007653568198
+ mjs = 0.3362
+ pbs = 0.6587
+ cjsws = 9.1602368e-11
+ mjsws = 0.2659
+ pbsws = 0.7418
+ cjswgs = 2.39155046e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.34 pmos
* DC IV MOS Parameters
+ lmin = 4e-06 lmax = 8e-06 wmin = 5.5e-07 wmax = 1.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 2.8e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 7.476e-9
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -7.916e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25000000.0
+ tnoib = 0.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.23e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-4.570656245e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope1/sqrt(l*w*mult))} lvth0 = 2.080235681e-07 wvth0 = 4.747328007e-08 pvth0 = -1.024001435e-13
+ k1 = 0.64774
+ k2 = -5.170463872e-02 lk2 = 3.213463431e-08 wk2 = 1.712101129e-08 pk2 = -2.518536007e-14
+ k3 = 3.39
+ dvt0 = 2.4422
+ dvt1 = 0.16136
+ dvt2 = 0.026237
+ dvt0w = 0.5
+ dvt1w = 1928100.0
+ dvt2w = -0.032
+ w0 = 1.0e-8
+ k3b = 1.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 123760.0
+ ua = -2.653280831e-09 lua = -4.912327788e-16 wua = -1.803516197e-16 pua = 9.069572049e-23
+ ub = 2.632245133e-18 lub = 1.158088580e-24 wub = 2.215087951e-25 pub = -4.880738773e-31
+ uc = 6.354273773e-11 luc = 5.131374465e-17 wuc = 1.027663415e-18 puc = -5.054650154e-23
+ rdsw = 484.7
+ prwb = 0.1
+ prwg = 0.052
+ wr = 1.0
+ u0 = 2.779025898e-03 lu0 = 9.102477651e-10 wu0 = -2.466351772e-10 pu0 = -8.176808257e-16
+ a0 = 1.003982928e+00 la0 = 1.987793321e-06 wa0 = 4.036235027e-07 pa0 = -1.210928120e-12
+ keta = -0.01258
+ a1 = 0.0
+ a2 = 0.46703705
+ ags = 1.598862947e-01 lags = 1.114398534e-06 wags = 7.016975883e-08 pags = -7.092779345e-13
+ b0 = 1.615043601e-08 lb0 = 7.407840499e-13 wb0 = -1.590895469e-14 pb0 = -7.297078468e-19
+ b1 = -3.704560111e-07 lb1 = -3.796799456e-15 wb1 = 3.649169528e-13 pb1 = 3.740029711e-21
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.1819+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))}
+ nfactor = {3.922606342e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 8.315130704e-06 wnfactor = 1.482795589e-06 pnfactor = -9.824123043e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -6.393105e-11
+ cdsc = 2.8125e-7
+ cdscb = 1.0e-4
+ cdscd = 1.0e-10
+ eta0 = 0.2
+ etab = -0.00025
+ dsub = 1.0
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.030097
+ pdiblc1 = 0.0
+ pdiblc2 = -1.294702722e-03 lpdiblc2 = 3.059842513e-08 wpdiblc2 = -4.884214698e-10 ppdiblc2 = -5.077277334e-15
+ pdiblcb = -0.025
+ drout = 0.43496
+ pscbe1 = 800000000.0
+ pscbe2 = 8.6797e-9
+ pvag = 0.0
+ delta = -3.869901880e-03 ldelta = 1.277812252e-07 wdelta = 6.940199893e-09 pdelta = -4.923749114e-14
+ alpha0 = 5.0449517e-13
+ alpha1 = -4.0583656e-18
+ beta0 = 6.2016506
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -1.760800036e+00 lkt1 = 3.068629581e-06 wkt1 = 3.066786144e-07 pkt1 = -1.429532856e-12
+ kt2 = -0.055045
+ at = 2.543498940e+05 lat = 8.360216782e-02 wat = 2.182566515e-02 pat = -1.000457948e-7
+ ute = -4.199426246e-01 lute = 9.694071834e-07 wute = -2.990122802e-08 pute = 2.936297326e-13
+ ua1 = 6.682694880e-10 lua1 = 1.111262531e-16
+ ub1 = -2.875736061e-19 lub1 = 1.098779165e-24 wub1 = 5.844498170e-26 pub1 = -4.672325617e-31
+ uc1 = -9.961e-12
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+41
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 1.4472e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 2.0e-11
+ cgso = 2.0e-11
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 0.0
+ cgdl = 0.0
+ cf = 0.0
+ clc = 7.0e-8
+ cle = 0.492
+ dlc = -1.2e-8
+ dwc = 0.0
+ vfbcv = -1.0
+ acde = 0.44
+ moin = 8.7
+ noff = 2.6123
+ voffcv = 0.112
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007653568198
+ mjs = 0.3362
+ pbs = 0.6587
+ cjsws = 9.1602368e-11
+ mjsws = 0.2659
+ pbsws = 0.7418
+ cjswgs = 2.39155046e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.35 pmos
* DC IV MOS Parameters
+ lmin = 2e-06 lmax = 4e-06 wmin = 5.5e-07 wmax = 1.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 2.8e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 7.476e-9
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -7.916e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25000000.0
+ tnoib = 0.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.23e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-3.737729407e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope1/sqrt(l*w*mult))} lvth0 = -1.246807279e-07 wvth0 = -5.858932187e-10 pvth0 = 8.956741831e-14
+ k1 = 0.64774
+ k2 = -2.911305667e-02 lk2 = -5.810518105e-08 wk2 = 3.905036416e-09 pk2 = 2.760452997e-14
+ k3 = 3.39
+ dvt0 = 2.4422
+ dvt1 = 0.16136
+ dvt2 = 0.026237
+ dvt0w = 0.5
+ dvt1w = 1928100.0
+ dvt2w = -0.032
+ w0 = 1.0e-8
+ k3b = 1.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 123760.0
+ ua = -2.897261180e-09 lua = 4.833223284e-16 wua = -8.756960455e-17 pua = -2.799127610e-22
+ ub = 3.077949920e-18 lub = -6.222346207e-25 wub = 5.300228552e-27 pub = 3.755496210e-31
+ uc = 7.638915888e-11 wuc = -1.162667805e-17
+ rdsw = 484.7
+ prwb = 0.1
+ prwg = 0.052
+ wr = 1.0
+ u0 = 2.800208761e-03 lu0 = 8.256349392e-10 wu0 = -3.632143723e-10 pu0 = -3.520168887e-16
+ a0 = 1.735020033e+00 la0 = -9.322612927e-07 wa0 = -2.440890758e-08 pa0 = 4.988045401e-13
+ keta = -0.01258
+ a1 = 0.0
+ a2 = 0.46703705
+ ags = 3.845415478e-01 lags = 2.170355909e-07 wags = -1.215280375e-07 pags = 5.643974304e-14
+ b0 = 2.721888053e-07 lb0 = -2.819356123e-13 wb0 = -2.681190383e-13 pb0 = 2.777201110e-19
+ b1 = -4.647777682e-07 lb1 = 3.729620271e-13 wb1 = 4.578284110e-13 pb1 = -3.673854988e-19
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.1819+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))}
+ nfactor = {7.356939409e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -5.402969298e-06 wnfactor = -1.178965346e-06 pnfactor = 8.080148368e-13
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -6.393105e-11
+ cdsc = 2.8125e-7
+ cdscb = 1.0e-4
+ cdscd = 1.0e-10
+ eta0 = 0.2
+ etab = -0.00025
+ dsub = 1.0
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.030097
+ pdiblc1 = 0.0
+ pdiblc2 = 1.212501191e-03 lpdiblc2 = 2.058364982e-08 wpdiblc2 = -1.181741272e-09 ppdiblc2 = -2.307880715e-15
+ pdiblcb = -0.025
+ drout = 0.43496
+ pscbe1 = 800000000.0
+ pscbe2 = 8.6797e-9
+ pvag = 0.0
+ delta = 3.276109190e-02 ldelta = -1.853761633e-08 wdelta = -1.133707573e-08 pdelta = 2.376925862e-14
+ alpha0 = 5.0449517e-13
+ alpha1 = -4.0583656e-18
+ beta0 = 6.2016506
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -8.903018098e-01 lkt1 = -4.084885324e-07 wkt1 = -1.717251892e-07 pkt1 = 4.814032968e-13
+ kt2 = -0.055045
+ at = 3.008993547e+05 lat = -1.023349977e-01 wat = 2.887468569e-03 pat = -2.439906233e-8
+ ute = -1.307996642e-01 lute = -1.855454574e-07 wute = 1.875539293e-08 pute = 9.927572590e-14
+ ua1 = 6.9609e-10
+ ub1 = 9.658631218e-20 lub1 = -4.357092130e-25 wub1 = -1.168899634e-25 pub1 = 2.331253430e-31
+ uc1 = -9.961e-12
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+41
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 1.4472e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 2.0e-11
+ cgso = 2.0e-11
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 0.0
+ cgdl = 0.0
+ cf = 0.0
+ clc = 7.0e-8
+ cle = 0.492
+ dlc = -1.2e-8
+ dwc = 0.0
+ vfbcv = -1.0
+ acde = 0.44
+ moin = 8.7
+ noff = 2.6123
+ voffcv = 0.112
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007653568198
+ mjs = 0.3362
+ pbs = 0.6587
+ cjsws = 9.1602368e-11
+ mjsws = 0.2659
+ pbsws = 0.7418
+ cjswgs = 2.39155046e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.36 pmos
* DC IV MOS Parameters
+ lmin = 1.5e-06 lmax = 2e-06 wmin = 5.5e-07 wmax = 1.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 2.8e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 7.476e-9
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -7.916e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25000000.0
+ tnoib = 0.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.23e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-4.362883478e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope1/sqrt(l*w*mult))} wvth0 = 4.432356241e-8
+ k1 = 0.64774
+ k2 = -5.824722286e-02 wk2 = 1.774605626e-8
+ k3 = 3.39
+ dvt0 = 2.4422
+ dvt1 = 0.16136
+ dvt2 = 0.026237
+ dvt0w = 0.5
+ dvt1w = 1928100.0
+ dvt2w = -0.032
+ w0 = 1.0e-8
+ k3b = 1.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 123760.0
+ ua = -2.654921465e-09 wua = -2.279189633e-16
+ ub = 2.765959035e-18 wub = 1.936022848e-25
+ uc = 7.638915888e-11 wuc = -1.162667805e-17
+ rdsw = 484.7
+ prwb = 0.1
+ prwg = 0.052
+ wr = 1.0
+ u0 = 3.214185365e-03 wu0 = -5.397170241e-10
+ a0 = 1.267580556e+00 wa0 = 2.256936496e-7
+ keta = -0.01258
+ a1 = 0.0
+ a2 = 0.46703705
+ ags = 4.933640462e-01 wags = -9.322892844e-8
+ b0 = 1.308251810e-07 wb0 = -1.288690829e-13
+ b1 = -2.777731417e-07 wb1 = 2.736198777e-13
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.1819+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))}
+ nfactor = {4.647869364e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} wnfactor = -7.738235304e-7
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -6.393105e-11
+ cdsc = 2.8125e-7
+ cdscb = 1.0e-4
+ cdscd = 1.0e-10
+ eta0 = 0.2
+ etab = -0.00025
+ dsub = 1.0
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.030097
+ pdiblc1 = 0.0
+ pdiblc2 = 1.153322412e-02 wpdiblc2 = -2.338921735e-9
+ pdiblcb = -0.025
+ drout = 0.43496
+ pscbe1 = 800000000.0
+ pscbe2 = 8.6797e-9
+ pvag = 0.0
+ delta = 2.346625820e-02 wdelta = 5.809239762e-10
+ alpha0 = 5.0449517e-13
+ alpha1 = -4.0583656e-18
+ beta0 = 6.2016506
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -1.095119566e+00 wkt1 = 6.965231626e-8
+ kt2 = -0.055045
+ at = 2.495881845e+05 wat = -9.346317198e-3
+ ute = -2.238328859e-01 wute = 6.853263215e-8
+ ua1 = 6.9609e-10
+ ub1 = -1.2188e-19
+ uc1 = -9.961e-12
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+41
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 1.4472e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 2.0e-11
+ cgso = 2.0e-11
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 0.0
+ cgdl = 0.0
+ cf = 0.0
+ clc = 7.0e-8
+ cle = 0.492
+ dlc = -1.2e-8
+ dwc = 0.0
+ vfbcv = -1.0
+ acde = 0.44
+ moin = 8.7
+ noff = 2.6123
+ voffcv = 0.112
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007653568198
+ mjs = 0.3362
+ pbs = 0.6587
+ cjsws = 9.1602368e-11
+ mjsws = 0.2659
+ pbsws = 0.7418
+ cjswgs = 2.39155046e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.37 pmos
* DC IV MOS Parameters
+ lmin = 1e-06 lmax = 1.5e-06 wmin = 5.5e-07 wmax = 1.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 2.8e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 7.476e-9
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -7.916e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25000000.0
+ tnoib = 0.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.23e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-5.645526352e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope1/sqrt(l*w*mult))} lvth0 = 1.916781510e-07 wvth0 = 1.277077804e-07 pvth0 = -1.246093754e-13
+ k1 = 0.64774
+ k2 = -9.970197314e-02 lk2 = 6.194997882e-08 wk2 = 5.023281798e-08 pk2 = -4.854821672e-14
+ k3 = 3.39
+ dvt0 = 2.4422
+ dvt1 = 0.16136
+ dvt2 = 0.026237
+ dvt0w = 0.5
+ dvt1w = 1928100.0
+ dvt2w = -0.032
+ w0 = 1.0e-8
+ k3b = 1.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 5.213874296e+04 lvsat = 1.070308065e-01 wvsat = 7.055037601e-02 pvsat = -1.054304819e-7
+ ua = -1.915487792e-09 lua = -1.105009680e-15 wua = -9.562966236e-16 pua = 1.088487576e-21
+ ub = 1.970246112e-18 lub = 1.189113391e-24 wub = 9.774177076e-25 pub = -1.171333768e-30
+ uc = 1.198636970e-10 luc = -6.496834977e-17 wuc = -5.445118488e-17 puc = 6.399694301e-23
+ rdsw = 484.7
+ prwb = 0.1
+ prwg = 0.052
+ wr = 1.0
+ u0 = 4.869747491e-03 lu0 = -2.474072041e-09 wu0 = -2.198338009e-09 pu0 = 2.478643200e-15
+ a0 = 1.826995236e+00 la0 = -8.359892973e-07 wa0 = 3.210559183e-07 pa0 = -1.425093743e-13
+ keta = -1.079467086e-02 lketa = -2.667995871e-09 wketa = -1.758634901e-09 pketa = 2.628103996e-15
+ a1 = 0.0
+ a2 = 0.46703705
+ ags = 1.178576573e+00 lags = -1.023981600e-06 wags = -6.204024509e-07 pags = 7.878081120e-13
+ b0 = 3.426243341e-07 lb0 = -3.165126545e-13 wb0 = -3.375014151e-13 pb0 = 3.117801573e-19
+ b1 = -4.416923684e-07 lb1 = 2.449608924e-13 wb1 = 4.350881841e-13 pb1 = -2.412982371e-19
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.1819+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))}
+ nfactor = {1.202686792e+01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -1.102717544e-05 wnfactor = -4.271294132e-06 pnfactor = 5.226620067e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -6.393105e-11
+ cdsc = 2.8125e-7
+ cdscb = 1.0e-4
+ cdscd = 1.0e-10
+ eta0 = 0.2
+ etab = -0.00025
+ dsub = 1.0
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.030097
+ pdiblc1 = 0.0
+ pdiblc2 = 4.858378491e-03 lpdiblc2 = 9.974889315e-09 wpdiblc2 = -1.262984755e-08 ppdiblc2 = 1.537875954e-14
+ pdiblcb = -0.025
+ drout = 0.43496
+ pscbe1 = 800000000.0
+ pscbe2 = 8.6797e-9
+ pvag = 0.0
+ delta = -5.925143684e-02 ldelta = 1.236133235e-07 wdelta = 3.758912439e-08 pdelta = -5.530505469e-14
+ alpha0 = 5.0449517e-13
+ alpha1 = -4.0583656e-18
+ beta0 = 6.2016506
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -1.490517074e+00 lkt1 = 5.908820362e-07 wkt1 = 2.101800561e-07 pkt1 = -2.100046544e-13
+ kt2 = -2.105544821e-01 lkt2 = 2.323933701e-07 wkt2 = 1.154409877e-07 pkt2 = -1.725150120e-13
+ at = 2.918183708e+05 lat = -6.310879036e-02 wat = 9.733643574e-02 pat = -1.594267060e-7
+ ute = -2.139097634e-01 lute = -1.482911439e-08 wute = 6.774998138e-08 pute = 1.169593302e-15
+ ua1 = 9.979992208e-10 lua1 = -4.511731395e-16 wua1 = -1.903518465e-16 pua1 = 2.844617994e-22
+ ub1 = -5.388043613e-19 lub1 = 6.230517656e-25 wub1 = 1.933520078e-25 pub1 = -2.889452404e-31
+ uc1 = 8.453375214e-11 luc1 = -1.412129576e-16 wuc1 = -9.308186660e-17 puc1 = 1.391015414e-22
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+41
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 1.4472e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 2.0e-11
+ cgso = 2.0e-11
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 0.0
+ cgdl = 0.0
+ cf = 0.0
+ clc = 7.0e-8
+ cle = 0.492
+ dlc = -1.2e-8
+ dwc = 0.0
+ vfbcv = -1.0
+ acde = 0.44
+ moin = 8.7
+ noff = 2.6123
+ voffcv = 0.112
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007653568198
+ mjs = 0.3362
+ pbs = 0.6587
+ cjsws = 9.1602368e-11
+ mjsws = 0.2659
+ pbsws = 0.7418
+ cjswgs = 2.39155046e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 2.74e-6
+ sbref = 2.74e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.38 pmos
* DC IV MOS Parameters
+ lmin = 5e-07 lmax = 1e-06 wmin = 5.5e-07 wmax = 1.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 2.8e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 7.476e-9
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -7.916e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25000000.0
+ tnoib = 0.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.23e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope2/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-4.187973341e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope1/sqrt(l*w*mult))} lvth0 = 4.673907961e-08 wvth0 = 3.909141047e-08 pvth0 = -3.648925711e-14
+ k1 = 0.64774
+ k2 = -3.596466925e-02 lk2 = -1.430396165e-09 wk2 = 9.507396173e-10 pk2 = 4.578820029e-16
+ k3 = 3.39
+ dvt0 = 2.4422
+ dvt1 = 0.16136
+ dvt2 = 0.026237
+ dvt0w = 0.5
+ dvt1w = 1928100.0
+ dvt2w = -0.032
+ w0 = 1.0e-8
+ k3b = 1.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 1.863842903e+05 lvsat = -2.646296575e-02 wvsat = -4.296443268e-02 pvsat = 7.448643851e-9
+ ua = -3.101914627e-09 lua = 7.477316359e-17 wua = 2.513513751e-16 pua = -1.123975943e-22
+ ub = 3.331728366e-18 lub = -1.647445622e-25 wub = -4.416289008e-25 pub = 2.397661796e-31
+ uc = 6.494258832e-11 luc = -1.035479929e-17 wuc = 7.197363225e-18 puc = 2.693626773e-24
+ rdsw = 484.7
+ prwb = 0.1
+ prwg = 0.052
+ wr = 1.0
+ u0 = 2.503055668e-03 lu0 = -1.206336922e-10 wu0 = 2.286724479e-10 pu0 = 6.522400151e-17
+ a0 = 8.118717710e-01 la0 = 1.734494764e-07 wa0 = 3.534972617e-07 pa0 = -1.747690462e-13
+ keta = -1.347769164e-02 wketa = 8.842693590e-10
+ a1 = 0.0
+ a2 = 0.46703705
+ ags = 3.276448171e-01 lags = -1.778150620e-07 wags = 6.029519200e-08 pags = 1.109223759e-13
+ b0 = 7.610056454e-08 lb0 = -5.148141799e-14 wb0 = 3.237379506e-14 pb0 = -5.602375171e-20
+ b1 = -1.463818407e-07 lb1 = -4.869589637e-14 wb1 = 3.528847055e-14 pb1 = 1.562625980e-19
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.1819+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))}
+ nfactor = {7.391799567e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 1.973014698e-07 wnfactor = 7.262950667e-07 pnfactor = 2.570173677e-13
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -6.393105e-11
+ cdsc = 2.8125e-7
+ cdscb = 1.0e-4
+ cdscd = 1.0e-10
+ eta0 = 0.2
+ etab = -0.00025
+ dsub = 1.0
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.030097
+ pdiblc1 = 0.0
+ pdiblc2 = 1.300374711e-02 lpdiblc2 = 1.875134762e-09 wpdiblc2 = -2.625827157e-08 ppdiblc2 = 2.893086438e-14
+ pdiblcb = -0.025
+ drout = 0.43496
+ pscbe1 = 800000000.0
+ pscbe2 = 8.6797e-9
+ pvag = 0.0
+ delta = 3.609779515e-02 ldelta = 2.879804718e-08 wdelta = -4.183454679e-09 pdelta = -1.376640207e-14
+ alpha0 = 5.0449517e-13
+ alpha1 = -4.0583656e-18
+ beta0 = 6.2016506
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -1.051092167e+00 lkt1 = 1.539179087e-07 wkt1 = 1.116064022e-07 pkt1 = -1.119830130e-13
+ kt2 = 5.603687518e-02 lkt2 = -3.270507562e-08 wkt2 = -7.564287926e-08 pkt2 = 1.749878530e-14
+ at = 4.406018237e+05 lat = -2.110590560e-01 wat = -1.710538781e-01 pat = 1.074606221e-7
+ ute = -6.499298767e-02 lute = -1.629119561e-07 wute = -1.873043193e-08 pute = 8.716571630e-14
+ ua1 = -7.440364279e-12 lua1 = 5.486359839e-16 wua1 = 3.909116142e-16 pua1 = -2.935465859e-22
+ ub1 = 1.221374061e-18 lub1 = -1.127269657e-24 wub1 = -6.058788287e-25 pub1 = 5.058099033e-31
+ uc1 = -8.568713394e-11 luc1 = 2.805469152e-17 wuc1 = 6.189816964e-17 puc1 = -1.501060659e-23
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+41
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 1.4472e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 2.0e-11
+ cgso = 2.0e-11
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 0.0
+ cgdl = 0.0
+ cf = 0.0
+ clc = 7.0e-8
+ cle = 0.492
+ dlc = -1.2e-8
+ dwc = 0.0
+ vfbcv = -1.0
+ acde = 0.44
+ moin = 8.7
+ noff = 2.6123
+ voffcv = 0.112
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007653568198
+ mjs = 0.3362
+ pbs = 0.6587
+ cjsws = 9.1602368e-11
+ mjsws = 0.2659
+ pbsws = 0.7418
+ cjswgs = 2.39155046e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 1.74e-6
+ sbref = 1.74e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.39 pmos
* DC IV MOS Parameters
+ lmin = 3.5e-07 lmax = 5e-07 wmin = 5.5e-07 wmax = 1.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 2.8e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 7.476e-9
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -7.916e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25000000.0
+ tnoib = 0.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.23e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope3/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-1.495123461e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope1/sqrt(l*w*mult))} lvth0 = -8.639541843e-08 wvth0 = -1.427328148e-07 pvth0 = 5.340463987e-14
+ k1 = 0.64774
+ k2 = -4.285005839e-02 lk2 = 1.973740224e-09 wk2 = -1.156816495e-08 pk2 = 6.647228421e-15
+ k3 = 3.39
+ dvt0 = 2.4422
+ dvt1 = 0.16136
+ dvt2 = 0.026237
+ dvt0w = 0.5
+ dvt1w = 1928100.0
+ dvt2w = -0.032
+ w0 = 1.0e-8
+ k3b = 1.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 1.637122457e+05 lvsat = -1.525390691e-02 wvsat = -5.959770282e-02 pvsat = 1.567213261e-8
+ ua = -3.076683126e-09 lua = 6.229870963e-17 wua = 2.386014056e-16 pua = -1.060940094e-22
+ ub = 2.612994519e-18 lub = 1.905974519e-25 wub = -8.036427329e-26 pub = 6.115694775e-32
+ uc = 1.607392219e-11 luc = 1.380586924e-17 wuc = 4.015260322e-17 puc = -1.359944388e-23
+ rdsw = 484.7
+ prwb = 0.1
+ prwg = 0.052
+ wr = 1.0
+ u0 = 8.659502652e-04 lu0 = 6.887512189e-10 wu0 = 1.187743154e-09 pu0 = -4.089405556e-16
+ a0 = 1.1627
+ keta = -1.727227166e-02 lketa = 1.876040360e-09 wketa = 2.914551807e-09 pketa = -1.003771642e-15
+ a1 = 0.0
+ a2 = 0.46703705
+ ags = -7.446080985e-01 lags = 3.523067795e-07 wags = 9.865926523e-07 pags = -3.470390885e-13
+ b0 = 7.894683512e-07 lb0 = -4.041704517e-13 wb0 = -7.386199123e-13 pb0 = 3.251555372e-19
+ b1 = -1.841702328e-06 lb1 = 7.894705525e-13 wb1 = 1.711615945e-12 pb1 = -6.725137054e-19
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {2.231116726e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = -2.002377709e-07 wvoff = -6.529173224e-08 pvoff = 3.228023242e-14
+ nfactor = {-9.890587250e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 5.452658377e-06 wnfactor = 6.620834220e-06 pnfactor = -2.657242790e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -6.393105e-11
+ cdsc = 2.8125e-7
+ cdscb = 1.0e-4
+ cdscd = 1.0e-10
+ eta0 = 0.2
+ etab = -0.00025
+ dsub = 1.0
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.030097
+ pdiblc1 = 0.0
+ pdiblc2 = -2.703778191e-03 lpdiblc2 = 9.640935270e-09 wpdiblc2 = -4.489995143e-08 ppdiblc2 = 3.814731091e-14
+ pdiblcb = -0.025
+ drout = 0.43496
+ pscbe1 = 800000000.0
+ pscbe2 = 8.6797e-9
+ pvag = 0.0
+ delta = 1.509909476e-01 ldelta = -2.800512739e-08 wdelta = -6.545113965e-08 pdelta = 1.652434138e-14
+ alpha0 = 5.0449517e-13
+ alpha1 = -4.0583656e-18
+ beta0 = 6.2016506
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -1.217657857e-01 lkt1 = -3.055410542e-07 wkt1 = -7.148166835e-07 pkt1 = 2.966005606e-13
+ kt2 = 1.626020472e-01 lkt2 = -8.539089664e-08 wkt2 = -1.326603614e-07 pkt2 = 4.568822846e-14
+ at = -4.433949910e+04 lat = 2.869593405e-02 wat = 1.874991537e-01 pat = -6.980799686e-8
+ ute = -8.127409949e-01 lute = 2.067746586e-07 wute = 5.193692717e-07 pute = -1.788707772e-13
+ ua1 = 1.972651465e-09 lua1 = -4.303214166e-16 wua1 = -6.685325589e-16 pua1 = 2.302426133e-22
+ ub1 = -2.955731024e-18 lub1 = 9.378910967e-25 wub1 = 1.375089403e-24 pub1 = -4.735807904e-31
+ uc1 = -1.642735167e-10 luc1 = 6.690779914e-17 wuc1 = 1.039456565e-16 puc1 = -3.579888411e-23
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+41
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 1.4472e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 2.0e-11
+ cgso = 2.0e-11
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 0.0
+ cgdl = 0.0
+ cf = 0.0
+ clc = 7.0e-8
+ cle = 0.492
+ dlc = -1.2e-8
+ dwc = 0.0
+ vfbcv = -1.0
+ acde = 0.44
+ moin = 8.7
+ noff = 2.6123
+ voffcv = 0.112
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007653568198
+ mjs = 0.3362
+ pbs = 0.6587
+ cjsws = 9.1602368e-11
+ mjsws = 0.2659
+ pbsws = 0.7418
+ cjswgs = 2.39155046e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 1.44e-6
+ sbref = 1.44e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.40 pmos
* DC IV MOS Parameters
+ lmin = 2.0e-05 lmax = 1.0e-04 wmin = 4.2e-07 wmax = 5.5e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 2.8e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 7.476e-9
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -7.916e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25000000.0
+ tnoib = 0.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.23e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-2.796856678e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope1/sqrt(l*w*mult))} wvth0 = -4.631992516e-8
+ k1 = 0.64774
+ k2 = 9.844950209e-03 wk2 = -1.681064647e-8
+ k3 = 3.39
+ dvt0 = 2.4422
+ dvt1 = 0.16136
+ dvt2 = 0.026237
+ dvt0w = 0.5
+ dvt1w = 1928100.0
+ dvt2w = -0.032
+ w0 = 1.0e-8
+ k3b = 1.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 123760.0
+ ua = -3.354638400e-09 wua = 1.733760978e-16
+ ub = 3.679898369e-18 wub = -3.225795667e-25
+ uc = 5.987805477e-11 wuc = 1.000246718e-19
+ rdsw = 484.7
+ prwb = 0.1
+ prwg = 0.052
+ wr = 1.0
+ u0 = 1.887468671e-03 wu0 = 1.890299590e-10
+ a0 = 2.042018468e+00 wa0 = -1.702086499e-7
+ keta = -0.01258
+ a1 = 0.0
+ a2 = 0.46703705
+ ags = 6.141664240e-01 wags = -1.870294655e-7
+ b0 = 2.402889743e-07 wb0 = -1.775321230e-13
+ b1 = -2.216963188e-07 wb1 = 2.855370965e-13
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {2.746825686e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} wvoff = -2.442935902e-7
+ nfactor = {1.084687183e+01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} wnfactor = -2.894380587e-6
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -6.393105e-11
+ cdsc = 2.8125e-7
+ cdscb = 1.0e-4
+ cdscd = 1.0e-10
+ eta0 = 0.2
+ etab = -0.00025
+ dsub = 1.0
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -4.524491454e-01 wpclm = 2.581853500e-7
+ pdiblc1 = 0.0
+ pdiblc2 = 1.367614996e-03 wpdiblc2 = -5.001066884e-10
+ pdiblcb = -0.025
+ drout = 4.620670585e-01 wdrout = -1.450357742e-8
+ pscbe1 = 800000000.0
+ pscbe2 = 8.6797e-9
+ pvag = 0.0
+ delta = 1.031492148e-02 wdelta = 1.743763446e-9
+ alpha0 = 5.0449517e-13
+ alpha1 = -4.0583656e-18
+ beta0 = 6.2016506
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -2.268687071e+00 wkt1 = 6.049825568e-7
+ kt2 = -0.055045
+ at = 2.574397569e+05 wat = 1.325326902e-2
+ ute = -6.244466554e-01 wute = 1.811280099e-7
+ ua1 = 6.8217e-10
+ ub1 = -7.061596185e-20 wub1 = -4.254382709e-26
+ uc1 = -9.961e-12
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+41
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 1.4472e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 2.0e-11
+ cgso = 2.0e-11
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 0.0
+ cgdl = 0.0
+ cf = 0.0
+ clc = 7.0e-8
+ cle = 0.492
+ dlc = -1.2e-8
+ dwc = 0.0
+ vfbcv = -1.0
+ acde = 0.44
+ moin = 8.7
+ noff = 2.6123
+ voffcv = 0.112
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007653568198
+ mjs = 0.3362
+ pbs = 0.6587
+ cjsws = 9.1602368e-11
+ mjsws = 0.2659
+ pbsws = 0.7418
+ cjswgs = 2.39155046e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.41 pmos
* DC IV MOS Parameters
+ lmin = 8e-06 lmax = 2.0e-05 wmin = 4.2e-07 wmax = 5.5e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 2.8e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 7.476e-9
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -7.916e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25000000.0
+ tnoib = 0.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.23e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-2.303075165e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope1/sqrt(l*w*mult))} lvth0 = -9.872865089e-07 wvth0 = -7.273960627e-08 pvth0 = 5.282456720e-13
+ k1 = 0.64774
+ k2 = 2.518753693e-02 lk2 = -3.067658159e-07 wk2 = -2.501966681e-08 pk2 = 1.641344363e-13
+ k3 = 3.39
+ dvt0 = 2.4422
+ dvt1 = 0.16136
+ dvt2 = 0.026237
+ dvt0w = 0.5
+ dvt1w = 1928100.0
+ dvt2w = -0.032
+ w0 = 1.0e-8
+ k3b = 1.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 123760.0
+ ua = -3.354638400e-09 wua = 1.733760978e-16
+ ub = 3.679898369e-18 wub = -3.225795667e-25
+ uc = 5.987805477e-11 wuc = 1.000246718e-19
+ rdsw = 484.7
+ prwb = 0.1
+ prwg = 0.052
+ wr = 1.0
+ u0 = 1.911005206e-03 lu0 = -4.705988913e-10 wu0 = 1.764367831e-10 pu0 = 2.517929956e-16
+ a0 = 1.691430168e+00 la0 = 7.009802693e-06 wa0 = 1.737291849e-08 pa0 = -3.750580911e-12
+ keta = -0.01258
+ a1 = 0.0
+ a2 = 0.46703705
+ ags = 6.141664240e-01 wags = -1.870294655e-7
+ b0 = 5.683038708e-07 lb0 = -6.558461045e-12 wb0 = -3.530358373e-13 pb0 = 3.509091465e-18
+ b1 = -1.020502107e-06 lb1 = 1.597164245e-11 wb1 = 7.129365358e-13 pb1 = -8.545595348e-18
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {5.788578758e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = -6.081802763e-06 wvoff = -4.070419799e-07 pvoff = 3.254056404e-12
+ nfactor = {1.359968534e+01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -5.504085454e-05 wnfactor = -4.367267953e-06 pnfactor = 2.944949914e-11
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -6.393105e-11
+ cdsc = 2.8125e-7
+ cdscb = 1.0e-4
+ cdscd = 1.0e-10
+ eta0 = 0.2
+ etab = -0.00025
+ dsub = 1.0
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -4.524491454e-01 wpclm = 2.581853500e-7
+ pdiblc1 = 0.0
+ pdiblc2 = 3.630289878e-03 lpdiblc2 = -4.524082665e-08 wpdiblc2 = -1.710746358e-09 ppdiblc2 = 2.420601382e-14
+ pdiblcb = -0.025
+ drout = 4.620670585e-01 wdrout = -1.450357742e-8
+ pscbe1 = 800000000.0
+ pscbe2 = 8.6797e-9
+ pvag = 0.0
+ delta = 2.189948808e-02 ldelta = -2.316264584e-07 wdelta = -4.454535745e-09 pdelta = 1.239312733e-13
+ alpha0 = 5.0449517e-13
+ alpha1 = -4.0583656e-18
+ beta0 = 6.2016506
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -3.039586943e+00 lkt1 = 1.541368041e-05 wkt1 = 1.017450992e-06 pkt1 = -8.247058879e-12
+ kt2 = -0.055045
+ at = 2.233565131e+05 lat = 6.814740096e-01 wat = 3.148944044e-02 pat = -3.646213059e-7
+ ute = -6.244466554e-01 wute = 1.811280099e-7
+ ua1 = 6.8217e-10
+ ub1 = -1.764370963e-20 lub1 = -1.059148400e-24 wub1 = -7.088652469e-26 pub1 = 5.666952330e-31
+ uc1 = -9.961e-12
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+41
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 1.4472e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 2.0e-11
+ cgso = 2.0e-11
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 0.0
+ cgdl = 0.0
+ cf = 0.0
+ clc = 7.0e-8
+ cle = 0.492
+ dlc = -1.2e-8
+ dwc = 0.0
+ vfbcv = -1.0
+ acde = 0.44
+ moin = 8.7
+ noff = 2.6123
+ voffcv = 0.112
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007653568198
+ mjs = 0.3362
+ pbs = 0.6587
+ cjsws = 9.1602368e-11
+ mjsws = 0.2659
+ pbsws = 0.7418
+ cjswgs = 2.39155046e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.42 pmos
* DC IV MOS Parameters
+ lmin = 4e-06 lmax = 8e-06 wmin = 4.2e-07 wmax = 5.5e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 2.8e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 7.476e-9
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -7.916e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25000000.0
+ tnoib = 0.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.23e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope2/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-3.949477174e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope1/sqrt(l*w*mult))} lvth0 = 3.289131133e-07 wvth0 = 1.423721812e-08 pvth0 = -1.670818528e-13
+ k1 = 0.64774
+ k2 = -1.887788126e-02 lk2 = 4.551076326e-08 wk2 = -4.428796362e-10 pk2 = -3.234223111e-14
+ k3 = 3.39
+ dvt0 = 2.4422
+ dvt1 = 0.16136
+ dvt2 = 0.026237
+ dvt0w = 0.5
+ dvt1w = 1928100.0
+ dvt2w = -0.032
+ w0 = 1.0e-8
+ k3b = 1.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 123760.0
+ ua = -3.406803156e-09 lua = 4.170259269e-16 wua = 2.228189933e-16 pua = -3.952662835e-22
+ ub = 4.024686478e-18 lub = -2.756374060e-24 wub = -5.235141620e-25 pub = 1.606351529e-30
+ uc = 1.008054692e-10 luc = -3.271901221e-16 wuc = -1.890968655e-17 puc = 1.519712354e-22
+ rdsw = 484.7
+ prwb = 0.1
+ prwg = 0.052
+ wr = 1.0
+ u0 = 2.499764223e-03 lu0 = -5.177373973e-09 wu0 = -9.721677621e-11 pu0 = 2.439489010e-15
+ a0 = 2.920394094e+00 la0 = -2.815026516e-06 wa0 = -6.217484589e-07 pa0 = 1.358811028e-12
+ keta = -0.01258
+ a1 = 0.0
+ a2 = 0.46703705
+ ags = 7.229168068e-01 lags = -8.693940601e-07 wags = -2.310785906e-07 pags = 3.521463253e-13
+ b0 = -2.852271971e-07 lb0 = 2.650077240e-13 wb0 = 1.453425452e-13 pb0 = -4.751446752e-19
+ b1 = 1.949399093e-06 lb1 = -7.770935701e-12 wb1 = -8.763168808e-13 pb1 = 4.159532165e-18
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.1819+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))}
+ nfactor = {8.691373377e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -1.580184536e-05 wnfactor = -1.068723675e-06 pnfactor = 3.079616767e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -6.393105e-11
+ cdsc = 2.8125e-7
+ cdscb = 1.0e-4
+ cdscd = 1.0e-10
+ eta0 = 0.2
+ etab = -0.00025
+ dsub = 1.0
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -4.524491454e-01 wpclm = 2.581853500e-7
+ pdiblc1 = 0.0
+ pdiblc2 = 1.563549316e-03 lpdiblc2 = -2.871847591e-08 wpdiblc2 = -2.017723507e-09 ppdiblc2 = 2.666011193e-14
+ pdiblcb = -0.025
+ drout = 4.620670585e-01 wdrout = -1.450357742e-8
+ pscbe1 = 800000000.0
+ pscbe2 = 8.6797e-9
+ pvag = 0.0
+ delta = -4.113715150e-03 ldelta = -2.366650655e-08 wdelta = 7.070651696e-09 pdelta = 3.179431485e-14
+ alpha0 = 5.0449517e-13
+ alpha1 = -4.0583656e-18
+ beta0 = 6.2016506
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -8.833203689e-01 lkt1 = -1.824377089e-06 wkt1 = -1.628151262e-07 pkt1 = 1.188460576e-12
+ kt2 = -0.055045
+ at = 3.478857935e+05 lat = -3.140628697e-01 wat = -2.822053080e-02 pat = 1.127240882e-7
+ ute = -1.152407130e+00 lute = 4.220727217e-06 wute = 3.620024406e-07 pute = -1.445982549e-12
+ ua1 = 6.682694880e-10 lua1 = 1.111262531e-16
+ ub1 = -1.783404500e-19 lub1 = 2.255256215e-25
+ uc1 = -9.961e-12
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+41
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 1.4472e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 2.0e-11
+ cgso = 2.0e-11
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 0.0
+ cgdl = 0.0
+ cf = 0.0
+ clc = 7.0e-8
+ cle = 0.492
+ dlc = -1.2e-8
+ dwc = 0.0
+ vfbcv = -1.0
+ acde = 0.44
+ moin = 8.7
+ noff = 2.6123
+ voffcv = 0.112
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007653568198
+ mjs = 0.3362
+ pbs = 0.6587
+ cjsws = 9.1602368e-11
+ mjsws = 0.2659
+ pbsws = 0.7418
+ cjswgs = 2.39155046e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.43 pmos
* DC IV MOS Parameters
+ lmin = 2e-06 lmax = 4e-06 wmin = 4.2e-07 wmax = 5.5e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 2.8e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 7.476e-9
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -7.916e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25000000.0
+ tnoib = 0.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.23e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-3.469840158e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope1/sqrt(l*w*mult))} lvth0 = 1.373269035e-07 wvth0 = -1.491925395e-08 pvth0 = -5.061924083e-14
+ k1 = 0.64774
+ k2 = -7.819635061e-03 lk2 = 1.339704638e-09 wk2 = -7.487966229e-09 pk2 = -4.201337226e-15
+ k3 = 3.39
+ dvt0 = 2.4422
+ dvt1 = 0.16136
+ dvt2 = 0.026237
+ dvt0w = 0.5
+ dvt1w = 1928100.0
+ dvt2w = -0.032
+ w0 = 1.0e-8
+ k3b = 1.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 123760.0
+ ua = -3.261358213e-09 lua = -1.639393526e-16 wua = 1.072397848e-16 pua = 6.640330687e-23
+ ub = 3.252542285e-18 lub = 3.278787051e-25 wub = -8.811506757e-26 pub = -1.328066137e-31
+ uc = 1.889326160e-11 wuc = 1.913638680e-17
+ rdsw = 484.7
+ prwb = 0.1
+ prwg = 0.052
+ wr = 1.0
+ u0 = 1.192469579e-03 lu0 = 4.448375222e-11 wu0 = 4.970032615e-10 pu0 = 6.593649162e-17
+ a0 = 2.005615615e+00 la0 = 8.389646433e-07 wa0 = -1.691905321e-07 pa0 = -4.488863545e-13
+ keta = -0.01258
+ a1 = 0.0
+ a2 = 0.46703705
+ ags = 3.434268171e-01 lags = 6.464407545e-07 wags = -9.952968307e-08 pags = -1.733126309e-13
+ b0 = -1.414928926e-07 lb0 = -3.091245819e-13 wb0 = -4.677947317e-14 pb0 = 2.922675149e-19
+ b1 = -1.324640600e-06 lb1 = 5.306888446e-12 wb1 = 9.178962993e-13 pb1 = -3.007272962e-18
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.1819+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))}
+ nfactor = {7.479701334e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -1.096194255e-05 wnfactor = -1.244648869e-06 pnfactor = 3.782332359e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -6.393105e-11
+ cdsc = 2.8125e-7
+ cdscb = 1.0e-4
+ cdscd = 1.0e-10
+ eta0 = 0.2
+ etab = -0.00025
+ dsub = 1.0
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -4.524491454e-01 wpclm = 2.581853500e-7
+ pdiblc1 = 0.0
+ pdiblc2 = -1.691889235e-02 lpdiblc2 = 4.510778909e-08 wpdiblc2 = 8.519424580e-09 ppdiblc2 = -1.542947238e-14
+ pdiblcb = -0.025
+ drout = 4.620670585e-01 wdrout = -1.450357742e-8
+ pscbe1 = 800000000.0
+ pscbe2 = 8.6797e-9
+ pvag = 0.0
+ delta = -4.848766842e-02 ldelta = 1.535808124e-07 wdelta = 3.213491098e-08 pdelta = -6.832236244e-14
+ alpha0 = 5.0449517e-13
+ alpha1 = -4.0583656e-18
+ beta0 = 6.2016506
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -1.824013459e+00 lkt1 = 1.933127390e-06 wkt1 = 3.278553613e-07 pkt1 = -7.714736192e-13
+ kt2 = -0.055045
+ at = 3.062960080e+05 lat = -1.479366304e-1
+ ute = -1.433581237e-01 lute = 1.901818668e-07 wute = 2.547477154e-08 pute = -1.017564275e-13
+ ua1 = 6.9609e-10
+ ub1 = -1.2188e-19
+ uc1 = -9.961e-12
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+41
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 1.4472e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 2.0e-11
+ cgso = 2.0e-11
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 0.0
+ cgdl = 0.0
+ cf = 0.0
+ clc = 7.0e-8
+ cle = 0.492
+ dlc = -1.2e-8
+ dwc = 0.0
+ vfbcv = -1.0
+ acde = 0.44
+ moin = 8.7
+ noff = 2.6123
+ voffcv = 0.112
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007653568198
+ mjs = 0.3362
+ pbs = 0.6587
+ cjsws = 9.1602368e-11
+ mjsws = 0.2659
+ pbsws = 0.7418
+ cjswgs = 2.39155046e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.44 pmos
* DC IV MOS Parameters
+ lmin = 1.5e-06 lmax = 2e-06 wmin = 4.2e-07 wmax = 5.5e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 2.8e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 7.476e-9
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -7.916e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25000000.0
+ tnoib = 0.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.23e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-2.781277665e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope1/sqrt(l*w*mult))} wvth0 = -4.029994028e-8
+ k1 = 0.64774
+ k2 = -7.147901889e-03 wk2 = -9.594533230e-9
+ k3 = 3.39
+ dvt0 = 2.4422
+ dvt1 = 0.16136
+ dvt2 = 0.026237
+ dvt0w = 0.5
+ dvt1w = 1928100.0
+ dvt2w = -0.032
+ w0 = 1.0e-8
+ k3b = 1.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 123760.0
+ ua = -3.343558049e-09 wua = 1.405346639e-16
+ ub = 3.416941957e-18 wub = -1.547048258e-25
+ uc = 1.889326160e-11 wuc = 1.913638680e-17
+ rdsw = 484.7
+ prwb = 0.1
+ prwg = 0.052
+ wr = 1.0
+ u0 = 1.214773907e-03 wu0 = 5.300640776e-10
+ a0 = 2.426275785e+00 wa0 = -3.942639148e-7
+ keta = -0.01258
+ a1 = 0.0
+ a2 = 0.46703705
+ ags = 6.675547526e-01 wags = -1.864293175e-7
+ b0 = -2.964891732e-07 wb0 = 9.976460769e-14
+ b1 = 1.336254129e-06 wb1 = -5.899621852e-13
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.1819+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))}
+ nfactor = {1.983340246e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} wnfactor = 6.518274448e-7
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -6.393105e-11
+ cdsc = 2.8125e-7
+ cdscb = 1.0e-4
+ cdscd = 1.0e-10
+ eta0 = 0.2
+ etab = -0.00025
+ dsub = 1.0
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -4.524491454e-01 wpclm = 2.581853500e-7
+ pdiblc1 = 0.0
+ pdiblc2 = 5.698330418e-03 wpdiblc2 = 7.830264727e-10
+ pdiblcb = -0.025
+ drout = 4.620670585e-01 wdrout = -1.450357742e-8
+ pscbe1 = 800000000.0
+ pscbe2 = 8.6797e-9
+ pvag = 0.0
+ delta = 2.851835465e-02 wdelta = -2.122190121e-9
+ alpha0 = 5.0449517e-13
+ alpha1 = -4.0583656e-18
+ beta0 = 6.2016506
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -8.547357865e-01 wkt1 = -5.896454405e-8
+ kt2 = -0.055045
+ at = 232120.0
+ ute = -4.800018806e-02 wute = -2.554630119e-8
+ ua1 = 6.9609e-10
+ ub1 = -1.2188e-19
+ uc1 = -9.961e-12
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+41
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 1.4472e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 2.0e-11
+ cgso = 2.0e-11
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 0.0
+ cgdl = 0.0
+ cf = 0.0
+ clc = 7.0e-8
+ cle = 0.492
+ dlc = -1.2e-8
+ dwc = 0.0
+ vfbcv = -1.0
+ acde = 0.44
+ moin = 8.7
+ noff = 2.6123
+ voffcv = 0.112
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007653568198
+ mjs = 0.3362
+ pbs = 0.6587
+ cjsws = 9.1602368e-11
+ mjsws = 0.2659
+ pbsws = 0.7418
+ cjswgs = 2.39155046e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.45 pmos
* DC IV MOS Parameters
+ lmin = 1e-06 lmax = 1.5e-06 wmin = 4.2e-07 wmax = 5.5e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 2.8e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 7.476e-9
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -7.916e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25000000.0
+ tnoib = 0.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.23e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-2.100546892e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope1/sqrt(l*w*mult))} lvth0 = -1.017284067e-07 wvth0 = -6.196563655e-08 pvth0 = 3.237721651e-14
+ k1 = 0.64774
+ k2 = 1.793033905e-02 lk2 = -3.747692326e-08 wk2 = -1.270611539e-08 pk2 = 4.649948382e-15
+ k3 = 3.39
+ dvt0 = 2.4422
+ dvt1 = 0.16136
+ dvt2 = 0.026237
+ dvt0w = 0.5
+ dvt1w = 1928100.0
+ dvt2w = -0.032
+ w0 = 1.0e-8
+ k3b = 1.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 3.716797359e+05 lvsat = -3.704912534e-01 wvsat = -1.004193932e-01 pvsat = 1.500667412e-7
+ ua = -4.494026749e-09 lua = 1.719260425e-15 wua = 4.233454880e-16 pua = -4.226324955e-22
+ ub = 5.192268265e-18 lub = -2.653047635e-24 wub = -7.465188011e-25 pub = 8.844068047e-31
+ uc = -7.809398269e-11 luc = 1.449377379e-16 wuc = 5.146567573e-17 puc = -4.831288937e-23
+ rdsw = 484.7
+ prwb = 0.1
+ prwg = 0.052
+ wr = 1.0
+ u0 = 2.468516546e-04 lu0 = 1.446463014e-09 wu0 = 2.751331623e-10 pu0 = 3.809687598e-16
+ a0 = 4.443521928e+00 la0 = -3.014572636e-06 wa0 = -1.078911455e-06 pa0 = 1.023137284e-12
+ keta = -1.875998549e-02 lketa = 9.235370321e-09 wketa = 2.503190764e-09 pketa = -3.740768278e-15
+ a1 = 0.0
+ a2 = 0.46703705
+ ags = -9.074681559e-01 lags = 2.353714235e-06 wags = 4.957316092e-07 pags = -1.019421289e-12
+ b0 = -1.976643399e-06 lb0 = 2.510822475e-12 wb0 = 9.034181468e-13 pb0 = -1.200979849e-18
+ b1 = 5.746681201e-06 lb1 = -6.590942217e-12 wb1 = -2.875988717e-12 pb1 = 3.416238050e-18
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.1819+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))}
+ nfactor = {2.693733159e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -1.061611169e-06 wnfactor = 7.223809540e-07 pnfactor = -1.054351642e-13
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -6.393105e-11
+ cdsc = 2.8125e-7
+ cdscb = 1.0e-4
+ cdscd = 1.0e-10
+ eta0 = 0.2
+ etab = -0.00025
+ dsub = 1.0
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -4.524491454e-01 wpclm = 2.581853500e-7
+ pdiblc1 = 0.0
+ pdiblc2 = -4.490180179e-02 lpdiblc2 = 7.561683757e-08 wpdiblc2 = 1.399423738e-08 ppdiblc2 = -1.974283358e-14
+ pdiblcb = -0.025
+ drout = 4.620670585e-01 wdrout = -1.450357742e-8
+ pscbe1 = 800000000.0
+ pscbe2 = 8.6797e-9
+ pvag = 0.0
+ delta = 1.936825423e-02 ldelta = 1.367391006e-08 wdelta = -4.476184084e-09 pdelta = 3.517808579e-15
+ alpha0 = 5.0449517e-13
+ alpha1 = -4.0583656e-18
+ beta0 = 6.2016506
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -8.726649800e-01 lkt1 = 2.679338684e-08 wkt1 = -1.204004710e-07 pkt1 = 9.180984925e-14
+ kt2 = 5.203707200e-03 lkt2 = -9.003566804e-8
+ at = 9.767182471e+05 lat = -1.112727620e+00 wat = -2.691178733e-01 pat = 4.021697498e-7
+ ute = -1.800541895e-01 lute = 1.973414998e-07 wute = 4.963562433e-08 pute = -1.123518695e-13
+ ua1 = 3.733623339e-10 lua1 = 4.822842242e-16 wua1 = 1.438588705e-16 pua1 = -2.149826961e-22
+ ub1 = -4.568487561e-19 lub1 = 5.005773090e-25 wub1 = 1.495018251e-25 pub1 = -2.234155274e-31
+ uc1 = -8.943543680e-11 luc1 = 1.187665984e-16 wuc1 = -6.162975822e-33 puc1 = 1.175494351e-38
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+41
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 1.4472e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 2.0e-11
+ cgso = 2.0e-11
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 0.0
+ cgdl = 0.0
+ cf = 0.0
+ clc = 7.0e-8
+ cle = 0.492
+ dlc = -1.2e-8
+ dwc = 0.0
+ vfbcv = -1.0
+ acde = 0.44
+ moin = 8.7
+ noff = 2.6123
+ voffcv = 0.112
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007653568198
+ mjs = 0.3362
+ pbs = 0.6587
+ cjsws = 9.1602368e-11
+ mjsws = 0.2659
+ pbsws = 0.7418
+ cjswgs = 2.39155046e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 2.74e-6
+ sbref = 2.74e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.46 pmos
* DC IV MOS Parameters
+ lmin = 5e-07 lmax = 1e-06 wmin = 4.2e-07 wmax = 5.5e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 2.8e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 7.476e-9
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -7.916e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25000000.0
+ tnoib = 0.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.23e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope2/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-1.630336006e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope2/sqrt(l*w*mult))} lvth0 = -1.484861773e-07 wvth0 = -9.775446360e-08 pvth0 = 6.796562613e-14
+ k1 = 0.64774
+ k2 = 1.717679989e-02 lk2 = -3.672760392e-08 wk2 = -2.748249716e-08 pk2 = 1.934358242e-14
+ k3 = 3.39
+ dvt0 = 2.4422
+ dvt1 = 0.16136
+ dvt2 = 0.026237
+ dvt0w = 0.5
+ dvt1w = 1928100.0
+ dvt2w = -0.032
+ w0 = 1.0e-8
+ k3b = 1.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 1.375857016e+05 lvsat = -1.377081456e-01 wvsat = -1.685484537e-02 pvsat = 6.697015484e-8
+ ua = -2.759653720e-09 lua = -5.400115163e-18 wua = 6.822536163e-17 pua = -6.950104183e-23
+ ub = 2.124083669e-18 lub = 3.979551280e-25 wub = 2.045189795e-25 pub = -6.130516426e-32
+ uc = 8.818359686e-11 luc = -2.040868724e-17 wuc = -5.237691916e-18 puc = 8.072939411e-24
+ rdsw = 484.7
+ prwb = 0.1
+ prwg = 0.052
+ wr = 1.0
+ u0 = 5.427889941e-04 lu0 = 1.152182924e-09 wu0 = 1.277509211e-09 pu0 = -6.157939832e-16
+ a0 = 3.281140972e+00 la0 = -1.858701013e-06 wa0 = -9.676802856e-07 pa0 = 9.125290091e-13
+ keta = -9.472605846e-03 wketa = -1.258643787e-9
+ a1 = 0.0
+ a2 = 0.46703705
+ ags = 1.337411384e+00 lags = 1.214060196e-07 wags = -4.799783903e-07 pags = -4.917526545e-14
+ b0 = 1.236065455e-06 lb0 = -6.838952092e-13 wb0 = -5.882630995e-13 pb0 = 2.823479824e-19
+ b1 = -2.776613885e-06 lb1 = 1.884622416e-12 wb1 = 1.442588865e-12 pb1 = -8.781554986e-19
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.1819+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))}
+ nfactor = {-2.118325902e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 3.723500362e-06 wnfactor = 2.255197861e-06 pnfactor = -1.629668297e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -6.393105e-11
+ cdsc = 2.8125e-7
+ cdscb = 1.0e-4
+ cdscd = 1.0e-10
+ eta0 = 0.2
+ etab = -0.00025
+ dsub = 1.0
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -8.285602172e-01 lpclm = 3.740048498e-07 wpclm = 4.594228267e-07 ppclm = -2.001105469e-13
+ pdiblc1 = 0.0
+ pdiblc2 = -1.252641263e-01 lpdiblc2 = 1.555291331e-07 wpdiblc2 = 4.772167757e-08 ppdiblc2 = -5.328140011e-14
+ pdiblcb = -0.025
+ drout = 4.620670585e-01 wdrout = -1.450357742e-8
+ pscbe1 = 800000000.0
+ pscbe2 = 8.6797e-9
+ pvag = 0.0
+ delta = 9.424127375e-02 ldelta = -6.077982055e-08 wdelta = -3.529300662e-08 pdelta = 3.416205691e-14
+ alpha0 = 5.0449517e-13
+ alpha1 = -4.0583656e-18
+ beta0 = 6.2016506
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -5.637117044e-01 lkt1 = -2.804297504e-07 wkt1 = -1.491655395e-07 pkt1 = 1.204138333e-13
+ kt2 = -0.085339
+ at = -3.012027963e+05 lat = 1.580370651e-01 wat = 2.258472002e-01 pat = -9.002351928e-8
+ ute = 1.354712275e-01 lute = -1.164169749e-07 wute = -1.259884093e-07 pute = 6.228866957e-14
+ ua1 = 9.029117574e-10 lua1 = -4.429972254e-17 wua1 = -9.617046783e-17 pua1 = 2.370247795e-23
+ ub1 = 8.905531727e-19 lub1 = -8.392791689e-25 wub1 = -4.288737743e-25 pub1 = 3.517211686e-31
+ uc1 = 3.0e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+41
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 1.4472e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 2.0e-11
+ cgso = 2.0e-11
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 0.0
+ cgdl = 0.0
+ cf = 0.0
+ clc = 7.0e-8
+ cle = 0.492
+ dlc = -1.2e-8
+ dwc = 0.0
+ vfbcv = -1.0
+ acde = 0.44
+ moin = 8.7
+ noff = 2.6123
+ voffcv = 0.112
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007653568198
+ mjs = 0.3362
+ pbs = 0.6587
+ cjsws = 9.1602368e-11
+ mjsws = 0.2659
+ pbsws = 0.7418
+ cjswgs = 2.39155046e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 1.74e-6
+ sbref = 1.74e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.47 pmos
* DC IV MOS Parameters
+ lmin = 3.5e-07 lmax = 5e-07 wmin = 4.2e-07 wmax = 5.5e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 2.8e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 7.476e-9
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -7.916e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25000000.0
+ tnoib = 0.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.23e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope3/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-2.669101785e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope1/sqrt(l*w*mult))} lvth0 = -9.712959711e-08 wvth0 = -7.991933937e-08 pvth0 = 5.914794071e-14
+ k1 = 0.64774
+ k2 = -3.082103431e-02 lk2 = -1.299747469e-08 wk2 = -1.800427022e-08 pk2 = 1.465754702e-14
+ k3 = 3.39
+ dvt0 = 2.4422
+ dvt1 = 0.16136
+ dvt2 = 0.026237
+ dvt0w = 0.5
+ dvt1w = 1928100.0
+ dvt2w = -0.032
+ w0 = 1.0e-8
+ k3b = 1.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = -5.062851338e+05 lvsat = 1.806215954e-01 wvsat = 2.988830551e-01 pvsat = -8.913066314e-8
+ ua = -2.073443004e-09 lua = -3.446626931e-16 wua = -2.981802150e-16 pua = 1.116498753e-22
+ ub = 1.320790852e-18 lub = 7.951030964e-25 wub = 6.110267143e-25 pub = -2.622825884e-31
+ uc = 7.979688230e-11 luc = -1.626229556e-17 wuc = 6.057760859e-18 puc = 2.488467559e-24
+ rdsw = 484.7
+ prwb = 0.1
+ prwg = 0.052
+ wr = 1.0
+ u0 = 2.729224958e-03 lu0 = 7.120898296e-11 wu0 = 1.908017560e-10 pu0 = -7.852581736e-17
+ a0 = -4.783675508e-01 wa0 = 8.780499109e-7
+ keta = -9.472605846e-03 wketa = -1.258643787e-9
+ a1 = 0.0
+ a2 = 0.46703705
+ ags = 4.049647402e+00 lags = -1.219523467e-06 wags = -1.578564165e-06 pags = 4.939655414e-13
+ b0 = -4.852296558e-07 lb0 = 1.671130935e-13 wb0 = -5.659529299e-14 pb0 = 1.949141890e-20
+ b1 = 3.412430078e-06 lb1 = -1.175240919e-12 wb1 = -1.099597091e-12 pb1 = 3.787012380e-19
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {5.367323361e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = -3.552918269e-07 wvoff = -2.330938410e-07 pvoff = 1.152415950e-13
+ nfactor = {1.930965099e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 1.721530890e-06 wnfactor = 2.957362789e-07 pnfactor = -6.609104905e-13
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -6.393105e-11
+ cdsc = 2.8125e-7
+ cdscb = 1.0e-4
+ cdscd = 1.0e-10
+ eta0 = 0.2
+ etab = -0.00025
+ dsub = 1.0
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -7.207791588e-02 wpclm = 5.466848439e-8
+ pdiblc1 = 0.0
+ pdiblc2 = -7.566071834e-02 lpdiblc2 = 1.310052082e-07 wpdiblc2 = -5.864486519e-09 ppdiblc2 = -2.678840058e-14
+ pdiblcb = -0.025
+ drout = 4.620670585e-01 wdrout = -1.450357742e-8
+ pscbe1 = 800000000.0
+ pscbe2 = 8.6797e-9
+ pvag = 0.0
+ delta = 1.275507657e-01 ldelta = -7.724803336e-08 wdelta = -5.290951719e-08 pdelta = 4.287165974e-14
+ alpha0 = 5.0449517e-13
+ alpha1 = -4.0583656e-18
+ beta0 = 6.2016506
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -2.228086217e+00 lkt1 = 5.424370084e-07 wkt1 = 4.121658505e-07 pkt1 = -1.571084059e-13
+ kt2 = -0.085339
+ at = 3.651974523e+04 lat = -8.932959457e-03 wat = 1.442355768e-01 pat = -4.967473264e-8
+ ute = 1.579556000e-01 lute = -1.275332486e-7
+ ua1 = 1.020267349e-09 lua1 = -1.023203270e-16 wua1 = -1.589613423e-16 pua1 = 5.474628630e-23
+ ub1 = -2.126180082e-18 lub1 = 6.521937523e-25 wub1 = 9.312398306e-25 pub1 = -3.207189977e-31
+ uc1 = 3.0e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+41
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 1.4472e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 2.0e-11
+ cgso = 2.0e-11
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 0.0
+ cgdl = 0.0
+ cf = 0.0
+ clc = 7.0e-8
+ cle = 0.492
+ dlc = -1.2e-8
+ dwc = 0.0
+ vfbcv = -1.0
+ acde = 0.44
+ moin = 8.7
+ noff = 2.6123
+ voffcv = 0.112
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007653568198
+ mjs = 0.3362
+ pbs = 0.6587
+ cjsws = 9.1602368e-11
+ mjsws = 0.2659
+ pbsws = 0.7418
+ cjswgs = 2.39155046e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 1.44e-6
+ sbref = 1.44e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.ends sky130_fd_pr__pfet_01v8_lvt
