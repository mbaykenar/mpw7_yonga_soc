magic
tech sky130A
magscale 1 2
timestamp 1649977179
<< nwell >>
rect 2301 20338 3262 20816
rect 26300 19944 26966 20818
rect 3418 17147 4118 19651
rect 3418 17032 4139 17147
rect 3418 17006 3458 17032
rect 2884 16334 3458 16360
rect 3727 16334 4139 17032
rect 2884 16246 4139 16334
rect 2884 15334 3798 16246
rect 7789 15315 8341 16378
rect 21644 7946 22063 8677
<< pwell >>
rect 50 38005 258 39950
rect 24043 37567 27047 37703
rect 193 35941 365 37534
rect 243 32342 365 35941
rect 22797 37221 27047 37567
rect 243 31731 938 32342
rect 243 31679 1339 31731
rect 253 23855 358 31679
rect 973 27129 1339 31679
rect 17996 30731 18468 33357
rect 973 23855 1784 27129
rect 253 23803 1784 23855
rect 254 23566 1784 23803
rect 254 22263 1528 23566
rect 17996 23474 19038 30731
rect 688 16196 1046 22263
rect 22797 22089 23661 37221
rect 3458 16334 3727 17032
rect 200 11442 1252 12998
rect 19650 11648 25554 11655
rect 6720 11501 25554 11648
rect 6720 11358 19709 11501
rect 25074 11381 25554 11501
rect 6720 11320 19408 11358
rect 6720 11122 10354 11320
rect 14040 11290 19408 11320
rect 6720 9615 7272 11122
rect 10023 9615 10245 11122
rect 16259 11086 19408 11290
rect 25074 11227 26309 11381
rect 16259 10999 19676 11086
rect 6720 9553 10245 9615
rect 6720 9343 10633 9553
rect 16537 9508 16827 10305
rect 19522 9811 19676 10999
rect 26223 10396 26309 11227
rect 26223 9834 27879 10396
rect 142 8209 1872 8887
rect 6720 8471 7272 9343
rect 10423 8491 10633 9343
rect 23829 9032 24094 9460
rect 21668 8968 22888 8974
rect 20758 8916 22888 8968
rect 23540 8946 24094 9032
rect 20758 8780 22949 8916
rect 23820 8882 24094 8946
rect 20758 8536 21564 8780
rect 142 6175 872 8209
rect 7062 7254 7272 8471
rect 22144 8558 22949 8780
rect 27521 8404 27879 9834
rect 27244 7630 27879 8404
rect 14231 6956 15119 7063
rect 13004 6264 15119 6956
rect 142 4978 382 6175
rect 142 4182 434 4978
rect 142 4151 1074 4182
rect 142 3895 2146 4151
rect 142 3115 694 3895
rect 1313 3259 2146 3895
rect 1313 3115 3159 3259
rect 142 2507 3159 3115
rect 25786 1714 27906 2060
<< psubdiff >>
rect 76 39900 232 39924
rect 110 39866 198 39900
rect 76 39831 232 39866
rect 110 39797 198 39831
rect 76 39762 232 39797
rect 110 39728 198 39762
rect 76 39693 232 39728
rect 110 39659 198 39693
rect 76 39624 232 39659
rect 110 39590 198 39624
rect 76 39555 232 39590
rect 110 39521 198 39555
rect 76 39486 232 39521
rect 110 39452 198 39486
rect 76 39417 232 39452
rect 110 39383 198 39417
rect 76 39348 232 39383
rect 110 39314 198 39348
rect 76 39279 232 39314
rect 110 39245 198 39279
rect 76 39209 232 39245
rect 110 39175 198 39209
rect 76 39139 232 39175
rect 110 39105 198 39139
rect 76 39069 232 39105
rect 110 39035 198 39069
rect 76 38999 232 39035
rect 110 38965 198 38999
rect 76 38929 232 38965
rect 110 38895 198 38929
rect 76 38859 232 38895
rect 110 38825 198 38859
rect 76 38789 232 38825
rect 110 38755 198 38789
rect 76 38719 232 38755
rect 110 38685 198 38719
rect 76 38649 232 38685
rect 110 38615 198 38649
rect 76 38579 232 38615
rect 110 38545 198 38579
rect 76 38509 232 38545
rect 110 38475 198 38509
rect 76 38439 232 38475
rect 110 38405 198 38439
rect 76 38369 232 38405
rect 110 38335 198 38369
rect 76 38299 232 38335
rect 110 38265 198 38299
rect 76 38229 232 38265
rect 110 38195 198 38229
rect 76 38159 232 38195
rect 110 38125 198 38159
rect 76 38089 232 38125
rect 110 38055 198 38089
rect 76 38031 232 38055
rect 226 12948 1226 12972
rect 226 12914 233 12948
rect 267 12914 301 12948
rect 335 12914 369 12948
rect 403 12914 437 12948
rect 471 12914 505 12948
rect 539 12914 573 12948
rect 607 12914 641 12948
rect 675 12914 709 12948
rect 743 12914 777 12948
rect 811 12914 845 12948
rect 879 12914 913 12948
rect 947 12914 981 12948
rect 1015 12914 1049 12948
rect 1083 12914 1117 12948
rect 1151 12914 1185 12948
rect 1219 12914 1226 12948
rect 226 12877 1226 12914
rect 226 12843 233 12877
rect 267 12843 301 12877
rect 335 12843 369 12877
rect 403 12843 437 12877
rect 471 12843 505 12877
rect 539 12843 573 12877
rect 607 12843 641 12877
rect 675 12843 709 12877
rect 743 12843 777 12877
rect 811 12843 845 12877
rect 879 12843 913 12877
rect 947 12843 981 12877
rect 1015 12843 1049 12877
rect 1083 12843 1117 12877
rect 1151 12843 1185 12877
rect 1219 12843 1226 12877
rect 226 12806 1226 12843
rect 226 12772 233 12806
rect 267 12772 301 12806
rect 335 12772 369 12806
rect 403 12772 437 12806
rect 471 12772 505 12806
rect 539 12772 573 12806
rect 607 12772 641 12806
rect 675 12772 709 12806
rect 743 12772 777 12806
rect 811 12772 845 12806
rect 879 12772 913 12806
rect 947 12772 981 12806
rect 1015 12772 1049 12806
rect 1083 12772 1117 12806
rect 1151 12772 1185 12806
rect 1219 12772 1226 12806
rect 226 12735 1226 12772
rect 226 12701 233 12735
rect 267 12701 301 12735
rect 335 12701 369 12735
rect 403 12701 437 12735
rect 471 12701 505 12735
rect 539 12701 573 12735
rect 607 12701 641 12735
rect 675 12701 709 12735
rect 743 12701 777 12735
rect 811 12701 845 12735
rect 879 12701 913 12735
rect 947 12701 981 12735
rect 1015 12701 1049 12735
rect 1083 12701 1117 12735
rect 1151 12701 1185 12735
rect 1219 12701 1226 12735
rect 226 12664 1226 12701
rect 226 12630 233 12664
rect 267 12630 301 12664
rect 335 12630 369 12664
rect 403 12630 437 12664
rect 471 12630 505 12664
rect 539 12630 573 12664
rect 607 12630 641 12664
rect 675 12630 709 12664
rect 743 12630 777 12664
rect 811 12630 845 12664
rect 879 12630 913 12664
rect 947 12630 981 12664
rect 1015 12630 1049 12664
rect 1083 12630 1117 12664
rect 1151 12630 1185 12664
rect 1219 12630 1226 12664
rect 226 12593 1226 12630
rect 226 12559 233 12593
rect 267 12559 301 12593
rect 335 12559 369 12593
rect 403 12559 437 12593
rect 471 12559 505 12593
rect 539 12559 573 12593
rect 607 12559 641 12593
rect 675 12559 709 12593
rect 743 12559 777 12593
rect 811 12559 845 12593
rect 879 12559 913 12593
rect 947 12559 981 12593
rect 1015 12559 1049 12593
rect 1083 12559 1117 12593
rect 1151 12559 1185 12593
rect 1219 12559 1226 12593
rect 226 12522 1226 12559
rect 226 12488 233 12522
rect 267 12488 301 12522
rect 335 12488 369 12522
rect 403 12488 437 12522
rect 471 12488 505 12522
rect 539 12488 573 12522
rect 607 12488 641 12522
rect 675 12488 709 12522
rect 743 12488 777 12522
rect 811 12488 845 12522
rect 879 12488 913 12522
rect 947 12488 981 12522
rect 1015 12488 1049 12522
rect 1083 12488 1117 12522
rect 1151 12488 1185 12522
rect 1219 12488 1226 12522
rect 226 12451 1226 12488
rect 226 12417 233 12451
rect 267 12417 301 12451
rect 335 12417 369 12451
rect 403 12417 437 12451
rect 471 12417 505 12451
rect 539 12417 573 12451
rect 607 12417 641 12451
rect 675 12417 709 12451
rect 743 12417 777 12451
rect 811 12417 845 12451
rect 879 12417 913 12451
rect 947 12417 981 12451
rect 1015 12417 1049 12451
rect 1083 12417 1117 12451
rect 1151 12417 1185 12451
rect 1219 12417 1226 12451
rect 226 12380 1226 12417
rect 226 12346 233 12380
rect 267 12346 301 12380
rect 335 12346 369 12380
rect 403 12346 437 12380
rect 471 12346 505 12380
rect 539 12346 573 12380
rect 607 12346 641 12380
rect 675 12346 709 12380
rect 743 12346 777 12380
rect 811 12346 845 12380
rect 879 12346 913 12380
rect 947 12346 981 12380
rect 1015 12346 1049 12380
rect 1083 12346 1117 12380
rect 1151 12346 1185 12380
rect 1219 12346 1226 12380
rect 226 12309 1226 12346
rect 226 12275 233 12309
rect 267 12275 301 12309
rect 335 12275 369 12309
rect 403 12275 437 12309
rect 471 12275 505 12309
rect 539 12275 573 12309
rect 607 12275 641 12309
rect 675 12275 709 12309
rect 743 12275 777 12309
rect 811 12275 845 12309
rect 879 12275 913 12309
rect 947 12275 981 12309
rect 1015 12275 1049 12309
rect 1083 12275 1117 12309
rect 1151 12275 1185 12309
rect 1219 12275 1226 12309
rect 226 12238 1226 12275
rect 226 12204 233 12238
rect 267 12204 301 12238
rect 335 12204 369 12238
rect 403 12204 437 12238
rect 471 12204 505 12238
rect 539 12204 573 12238
rect 607 12204 641 12238
rect 675 12204 709 12238
rect 743 12204 777 12238
rect 811 12204 845 12238
rect 879 12204 913 12238
rect 947 12204 981 12238
rect 1015 12204 1049 12238
rect 1083 12204 1117 12238
rect 1151 12204 1185 12238
rect 1219 12204 1226 12238
rect 226 12167 1226 12204
rect 226 12133 233 12167
rect 267 12133 301 12167
rect 335 12133 369 12167
rect 403 12133 437 12167
rect 471 12133 505 12167
rect 539 12133 573 12167
rect 607 12133 641 12167
rect 675 12133 709 12167
rect 743 12133 777 12167
rect 811 12133 845 12167
rect 879 12133 913 12167
rect 947 12133 981 12167
rect 1015 12133 1049 12167
rect 1083 12133 1117 12167
rect 1151 12133 1185 12167
rect 1219 12133 1226 12167
rect 226 12096 1226 12133
rect 226 12062 233 12096
rect 267 12062 301 12096
rect 335 12062 369 12096
rect 403 12062 437 12096
rect 471 12062 505 12096
rect 539 12062 573 12096
rect 607 12062 641 12096
rect 675 12062 709 12096
rect 743 12062 777 12096
rect 811 12062 845 12096
rect 879 12062 913 12096
rect 947 12062 981 12096
rect 1015 12062 1049 12096
rect 1083 12062 1117 12096
rect 1151 12062 1185 12096
rect 1219 12062 1226 12096
rect 226 12025 1226 12062
rect 226 11991 233 12025
rect 267 11991 301 12025
rect 335 11991 369 12025
rect 403 11991 437 12025
rect 471 11991 505 12025
rect 539 11991 573 12025
rect 607 11991 641 12025
rect 675 11991 709 12025
rect 743 11991 777 12025
rect 811 11991 845 12025
rect 879 11991 913 12025
rect 947 11991 981 12025
rect 1015 11991 1049 12025
rect 1083 11991 1117 12025
rect 1151 11991 1185 12025
rect 1219 11991 1226 12025
rect 226 11954 1226 11991
rect 226 11920 233 11954
rect 267 11920 301 11954
rect 335 11920 369 11954
rect 403 11920 437 11954
rect 471 11920 505 11954
rect 539 11920 573 11954
rect 607 11920 641 11954
rect 675 11920 709 11954
rect 743 11920 777 11954
rect 811 11920 845 11954
rect 879 11920 913 11954
rect 947 11920 981 11954
rect 1015 11920 1049 11954
rect 1083 11920 1117 11954
rect 1151 11920 1185 11954
rect 1219 11920 1226 11954
rect 226 11883 1226 11920
rect 226 11849 233 11883
rect 267 11849 301 11883
rect 335 11849 369 11883
rect 403 11849 437 11883
rect 471 11849 505 11883
rect 539 11849 573 11883
rect 607 11849 641 11883
rect 675 11849 709 11883
rect 743 11849 777 11883
rect 811 11849 845 11883
rect 879 11849 913 11883
rect 947 11849 981 11883
rect 1015 11849 1049 11883
rect 1083 11849 1117 11883
rect 1151 11849 1185 11883
rect 1219 11849 1226 11883
rect 226 11812 1226 11849
rect 226 11778 233 11812
rect 267 11778 301 11812
rect 335 11778 369 11812
rect 403 11778 437 11812
rect 471 11778 505 11812
rect 539 11778 573 11812
rect 607 11778 641 11812
rect 675 11778 709 11812
rect 743 11778 777 11812
rect 811 11778 845 11812
rect 879 11778 913 11812
rect 947 11778 981 11812
rect 1015 11778 1049 11812
rect 1083 11778 1117 11812
rect 1151 11778 1185 11812
rect 1219 11778 1226 11812
rect 226 11741 1226 11778
rect 226 11707 233 11741
rect 267 11707 301 11741
rect 335 11707 369 11741
rect 403 11707 437 11741
rect 471 11707 505 11741
rect 539 11707 573 11741
rect 607 11707 641 11741
rect 675 11707 709 11741
rect 743 11707 777 11741
rect 811 11707 845 11741
rect 879 11707 913 11741
rect 947 11707 981 11741
rect 1015 11707 1049 11741
rect 1083 11707 1117 11741
rect 1151 11707 1185 11741
rect 1219 11707 1226 11741
rect 226 11670 1226 11707
rect 226 11636 233 11670
rect 267 11636 301 11670
rect 335 11636 369 11670
rect 403 11636 437 11670
rect 471 11636 505 11670
rect 539 11636 573 11670
rect 607 11636 641 11670
rect 675 11636 709 11670
rect 743 11636 777 11670
rect 811 11636 845 11670
rect 879 11636 913 11670
rect 947 11636 981 11670
rect 1015 11636 1049 11670
rect 1083 11636 1117 11670
rect 1151 11636 1185 11670
rect 1219 11636 1226 11670
rect 226 11598 1226 11636
rect 226 11564 233 11598
rect 267 11564 301 11598
rect 335 11564 369 11598
rect 403 11564 437 11598
rect 471 11564 505 11598
rect 539 11564 573 11598
rect 607 11564 641 11598
rect 675 11564 709 11598
rect 743 11564 777 11598
rect 811 11564 845 11598
rect 879 11564 913 11598
rect 947 11564 981 11598
rect 1015 11564 1049 11598
rect 1083 11564 1117 11598
rect 1151 11564 1185 11598
rect 1219 11564 1226 11598
rect 226 11526 1226 11564
rect 226 11492 233 11526
rect 267 11492 301 11526
rect 335 11492 369 11526
rect 403 11492 437 11526
rect 471 11492 505 11526
rect 539 11492 573 11526
rect 607 11492 641 11526
rect 675 11492 709 11526
rect 743 11492 777 11526
rect 811 11492 845 11526
rect 879 11492 913 11526
rect 947 11492 981 11526
rect 1015 11492 1049 11526
rect 1083 11492 1117 11526
rect 1151 11492 1185 11526
rect 1219 11492 1226 11526
rect 226 11468 1226 11492
rect 16285 11062 19382 11076
rect 16285 11028 16319 11062
rect 16353 11028 16388 11062
rect 16422 11028 16457 11062
rect 16491 11028 16526 11062
rect 16560 11028 16594 11062
rect 16628 11028 16662 11062
rect 16696 11028 16730 11062
rect 16764 11028 16798 11062
rect 16832 11028 16866 11062
rect 16900 11028 16934 11062
rect 16968 11028 17002 11062
rect 17036 11028 17070 11062
rect 17104 11028 17138 11062
rect 17172 11028 17206 11062
rect 17240 11028 17274 11062
rect 17308 11028 17342 11062
rect 17376 11028 17410 11062
rect 17444 11028 17478 11062
rect 17512 11028 17546 11062
rect 17580 11028 17614 11062
rect 17648 11028 17682 11062
rect 17716 11028 17750 11062
rect 17784 11028 17818 11062
rect 17852 11028 17886 11062
rect 17920 11028 17954 11062
rect 17988 11028 18022 11062
rect 18056 11028 18090 11062
rect 18124 11028 18158 11062
rect 18192 11028 18226 11062
rect 18260 11028 18294 11062
rect 18328 11028 18362 11062
rect 18396 11028 18430 11062
rect 18464 11028 18498 11062
rect 18532 11028 18566 11062
rect 18600 11028 18634 11062
rect 18668 11028 18702 11062
rect 18736 11028 18770 11062
rect 18804 11028 18838 11062
rect 18872 11028 18906 11062
rect 18940 11028 18974 11062
rect 19008 11028 19042 11062
rect 19076 11028 19110 11062
rect 19144 11028 19178 11062
rect 19212 11028 19246 11062
rect 19280 11028 19314 11062
rect 19348 11028 19382 11062
rect 16285 11025 19382 11028
rect 19548 11036 19650 11060
rect 19582 11002 19616 11036
rect 19548 10933 19650 11002
rect 19582 10899 19616 10933
rect 19548 10830 19650 10899
rect 19582 10796 19616 10830
rect 19548 10727 19650 10796
rect 19582 10693 19616 10727
rect 19548 10623 19650 10693
rect 19582 10589 19616 10623
rect 19548 10519 19650 10589
rect 19582 10485 19616 10519
rect 19548 10415 19650 10485
rect 19582 10381 19616 10415
rect 19548 10311 19650 10381
rect 16563 10255 16801 10279
rect 16597 10221 16631 10255
rect 16665 10221 16699 10255
rect 16733 10221 16767 10255
rect 16563 10182 16801 10221
rect 16597 10148 16631 10182
rect 16665 10148 16699 10182
rect 16733 10148 16767 10182
rect 16563 10109 16801 10148
rect 16597 10075 16631 10109
rect 16665 10075 16699 10109
rect 16733 10075 16767 10109
rect 16563 10036 16801 10075
rect 16597 10002 16631 10036
rect 16665 10002 16699 10036
rect 16733 10002 16767 10036
rect 16563 9962 16801 10002
rect 16597 9928 16631 9962
rect 16665 9928 16699 9962
rect 16733 9928 16767 9962
rect 16563 9888 16801 9928
rect 16597 9854 16631 9888
rect 16665 9854 16699 9888
rect 16733 9854 16767 9888
rect 16563 9814 16801 9854
rect 19582 10277 19616 10311
rect 19548 10207 19650 10277
rect 19582 10173 19616 10207
rect 19548 10103 19650 10173
rect 19582 10069 19616 10103
rect 19548 9999 19650 10069
rect 19582 9965 19616 9999
rect 19548 9895 19650 9965
rect 19582 9861 19616 9895
rect 19548 9837 19650 9861
rect 16597 9780 16631 9814
rect 16665 9780 16699 9814
rect 16733 9780 16767 9814
rect 16563 9740 16801 9780
rect 16597 9706 16631 9740
rect 16665 9706 16699 9740
rect 16733 9706 16767 9740
rect 16563 9666 16801 9706
rect 16597 9632 16631 9666
rect 16665 9632 16699 9666
rect 16733 9632 16767 9666
rect 16563 9592 16801 9632
rect 16597 9558 16631 9592
rect 16665 9558 16699 9592
rect 16733 9558 16767 9592
rect 16563 9534 16801 9558
rect 23566 8972 23590 9006
rect 23624 8972 23654 9006
<< nsubdiff >>
rect 3484 16360 3701 17006
<< mvpsubdiff >>
rect 24069 37674 27021 37677
rect 24069 37640 24093 37674
rect 24127 37640 24162 37674
rect 24196 37640 24231 37674
rect 24265 37640 24300 37674
rect 24334 37640 24369 37674
rect 24403 37640 24438 37674
rect 24472 37640 24507 37674
rect 24541 37640 24576 37674
rect 24610 37640 24645 37674
rect 24679 37640 24714 37674
rect 24748 37640 24783 37674
rect 24817 37640 24852 37674
rect 24886 37640 24921 37674
rect 24955 37640 24990 37674
rect 25024 37640 25059 37674
rect 25093 37640 25127 37674
rect 25161 37640 25195 37674
rect 25229 37640 25263 37674
rect 25297 37640 25331 37674
rect 25365 37640 25399 37674
rect 25433 37640 25467 37674
rect 25501 37640 25535 37674
rect 25569 37640 25603 37674
rect 25637 37640 25671 37674
rect 25705 37640 25739 37674
rect 25773 37640 25807 37674
rect 25841 37640 25875 37674
rect 25909 37640 25943 37674
rect 25977 37640 26011 37674
rect 26045 37640 26079 37674
rect 26113 37640 26147 37674
rect 26181 37640 26215 37674
rect 26249 37640 26283 37674
rect 26317 37640 26351 37674
rect 26385 37640 26419 37674
rect 26453 37640 26487 37674
rect 26521 37640 26555 37674
rect 26589 37640 26623 37674
rect 26657 37640 26691 37674
rect 26725 37640 26759 37674
rect 26793 37640 26827 37674
rect 26861 37640 26895 37674
rect 26929 37640 26963 37674
rect 26997 37640 27021 37674
rect 24069 37596 27021 37640
rect 24069 37562 24093 37596
rect 24127 37562 24162 37596
rect 24196 37562 24231 37596
rect 24265 37562 24300 37596
rect 24334 37562 24369 37596
rect 24403 37562 24438 37596
rect 24472 37562 24507 37596
rect 24541 37562 24576 37596
rect 24610 37562 24645 37596
rect 24679 37562 24714 37596
rect 24748 37562 24783 37596
rect 24817 37562 24852 37596
rect 24886 37562 24921 37596
rect 24955 37562 24990 37596
rect 25024 37562 25059 37596
rect 25093 37562 25127 37596
rect 25161 37562 25195 37596
rect 25229 37562 25263 37596
rect 25297 37562 25331 37596
rect 25365 37562 25399 37596
rect 25433 37562 25467 37596
rect 25501 37562 25535 37596
rect 25569 37562 25603 37596
rect 25637 37562 25671 37596
rect 25705 37562 25739 37596
rect 25773 37562 25807 37596
rect 25841 37562 25875 37596
rect 25909 37562 25943 37596
rect 25977 37562 26011 37596
rect 26045 37562 26079 37596
rect 26113 37562 26147 37596
rect 26181 37562 26215 37596
rect 26249 37562 26283 37596
rect 26317 37562 26351 37596
rect 26385 37562 26419 37596
rect 26453 37562 26487 37596
rect 26521 37562 26555 37596
rect 26589 37562 26623 37596
rect 26657 37562 26691 37596
rect 26725 37562 26759 37596
rect 26793 37562 26827 37596
rect 26861 37562 26895 37596
rect 26929 37562 26963 37596
rect 26997 37562 27021 37596
rect 24069 37541 27021 37562
rect 22823 37540 27021 37541
rect 22823 37517 23711 37540
rect 219 37484 339 37508
rect 253 37450 305 37484
rect 219 37415 339 37450
rect 253 37381 305 37415
rect 219 37346 339 37381
rect 253 37312 305 37346
rect 219 37277 339 37312
rect 253 37243 305 37277
rect 219 37208 339 37243
rect 253 37174 305 37208
rect 219 37139 339 37174
rect 253 37105 305 37139
rect 219 37070 339 37105
rect 253 37036 305 37070
rect 219 37001 339 37036
rect 253 36967 305 37001
rect 219 36932 339 36967
rect 253 36898 305 36932
rect 219 36863 339 36898
rect 253 36829 305 36863
rect 219 36794 339 36829
rect 253 36760 305 36794
rect 219 36725 339 36760
rect 253 36691 305 36725
rect 219 36655 339 36691
rect 253 36621 305 36655
rect 219 36585 339 36621
rect 253 36551 305 36585
rect 219 36515 339 36551
rect 253 36481 305 36515
rect 219 36445 339 36481
rect 253 36411 305 36445
rect 219 36375 339 36411
rect 253 36341 305 36375
rect 219 36305 339 36341
rect 253 36271 305 36305
rect 219 36235 339 36271
rect 253 36201 305 36235
rect 219 36165 339 36201
rect 253 36131 305 36165
rect 219 36095 339 36131
rect 253 36061 305 36095
rect 219 36025 339 36061
rect 253 35991 305 36025
rect 219 35967 339 35991
rect 269 35891 339 35967
rect 269 35857 278 35891
rect 312 35857 339 35891
rect 269 35823 339 35857
rect 269 35789 278 35823
rect 312 35789 339 35823
rect 269 35755 339 35789
rect 269 35721 278 35755
rect 312 35721 339 35755
rect 269 35687 339 35721
rect 269 35653 278 35687
rect 312 35653 339 35687
rect 269 35619 339 35653
rect 269 35585 278 35619
rect 312 35585 339 35619
rect 269 35551 339 35585
rect 269 35517 278 35551
rect 312 35517 339 35551
rect 269 35483 339 35517
rect 269 35449 278 35483
rect 312 35449 339 35483
rect 269 35415 339 35449
rect 269 35381 278 35415
rect 312 35381 339 35415
rect 269 35347 339 35381
rect 269 35313 278 35347
rect 312 35313 339 35347
rect 269 35279 339 35313
rect 269 35245 278 35279
rect 312 35245 339 35279
rect 269 35211 339 35245
rect 269 35177 278 35211
rect 312 35177 339 35211
rect 269 35143 339 35177
rect 269 35109 278 35143
rect 312 35109 339 35143
rect 269 35075 339 35109
rect 269 35041 278 35075
rect 312 35041 339 35075
rect 269 35006 339 35041
rect 269 34972 278 35006
rect 312 34972 339 35006
rect 269 34937 339 34972
rect 269 34903 278 34937
rect 312 34903 339 34937
rect 269 34868 339 34903
rect 269 34834 278 34868
rect 312 34834 339 34868
rect 269 34799 339 34834
rect 269 34765 278 34799
rect 312 34765 339 34799
rect 269 34730 339 34765
rect 269 34696 278 34730
rect 312 34696 339 34730
rect 269 34661 339 34696
rect 269 34627 278 34661
rect 312 34627 339 34661
rect 269 34592 339 34627
rect 269 34558 278 34592
rect 312 34558 339 34592
rect 269 34523 339 34558
rect 269 34489 278 34523
rect 312 34489 339 34523
rect 269 34454 339 34489
rect 269 34420 278 34454
rect 312 34420 339 34454
rect 269 34385 339 34420
rect 269 34351 278 34385
rect 312 34351 339 34385
rect 269 34316 339 34351
rect 269 34282 278 34316
rect 312 34282 339 34316
rect 269 34247 339 34282
rect 269 34213 278 34247
rect 312 34213 339 34247
rect 269 34178 339 34213
rect 269 34144 278 34178
rect 312 34144 339 34178
rect 269 34109 339 34144
rect 269 34075 278 34109
rect 312 34075 339 34109
rect 269 34040 339 34075
rect 269 34006 278 34040
rect 312 34006 339 34040
rect 269 33971 339 34006
rect 269 33937 278 33971
rect 312 33937 339 33971
rect 269 33902 339 33937
rect 269 33868 278 33902
rect 312 33868 339 33902
rect 269 33833 339 33868
rect 269 33799 278 33833
rect 312 33799 339 33833
rect 269 33764 339 33799
rect 269 33730 278 33764
rect 312 33730 339 33764
rect 269 33695 339 33730
rect 269 33661 278 33695
rect 312 33661 339 33695
rect 269 33626 339 33661
rect 269 33592 278 33626
rect 312 33592 339 33626
rect 269 33557 339 33592
rect 269 33523 278 33557
rect 312 33523 339 33557
rect 269 33488 339 33523
rect 269 33454 278 33488
rect 312 33454 339 33488
rect 269 33419 339 33454
rect 269 33385 278 33419
rect 312 33385 339 33419
rect 269 33350 339 33385
rect 269 33316 278 33350
rect 312 33316 339 33350
rect 22823 37483 22827 37517
rect 22861 37483 22897 37517
rect 22931 37483 22967 37517
rect 23001 37483 23037 37517
rect 23071 37483 23107 37517
rect 23141 37483 23177 37517
rect 23211 37483 23247 37517
rect 23281 37483 23317 37517
rect 23351 37483 23387 37517
rect 23421 37483 23457 37517
rect 23491 37483 23527 37517
rect 23561 37483 23597 37517
rect 23631 37506 23711 37517
rect 23745 37506 23794 37540
rect 23828 37506 23877 37540
rect 23911 37506 23959 37540
rect 23993 37518 27021 37540
rect 23993 37506 24093 37518
rect 23631 37484 24093 37506
rect 24127 37484 24162 37518
rect 24196 37484 24231 37518
rect 24265 37484 24300 37518
rect 24334 37484 24369 37518
rect 24403 37484 24438 37518
rect 24472 37484 24507 37518
rect 24541 37484 24576 37518
rect 24610 37484 24645 37518
rect 24679 37484 24714 37518
rect 24748 37484 24783 37518
rect 24817 37484 24852 37518
rect 24886 37484 24921 37518
rect 24955 37484 24990 37518
rect 25024 37484 25059 37518
rect 25093 37484 25127 37518
rect 25161 37484 25195 37518
rect 25229 37484 25263 37518
rect 25297 37484 25331 37518
rect 25365 37484 25399 37518
rect 25433 37484 25467 37518
rect 25501 37484 25535 37518
rect 25569 37484 25603 37518
rect 25637 37484 25671 37518
rect 25705 37484 25739 37518
rect 25773 37484 25807 37518
rect 25841 37484 25875 37518
rect 25909 37484 25943 37518
rect 25977 37484 26011 37518
rect 26045 37484 26079 37518
rect 26113 37484 26147 37518
rect 26181 37484 26215 37518
rect 26249 37484 26283 37518
rect 26317 37484 26351 37518
rect 26385 37484 26419 37518
rect 26453 37484 26487 37518
rect 26521 37484 26555 37518
rect 26589 37484 26623 37518
rect 26657 37484 26691 37518
rect 26725 37484 26759 37518
rect 26793 37484 26827 37518
rect 26861 37484 26895 37518
rect 26929 37484 26963 37518
rect 26997 37484 27021 37518
rect 23631 37483 27021 37484
rect 22823 37454 27021 37483
rect 22823 37449 23711 37454
rect 22823 37415 22827 37449
rect 22861 37415 22897 37449
rect 22931 37415 22967 37449
rect 23001 37415 23037 37449
rect 23071 37415 23107 37449
rect 23141 37415 23177 37449
rect 23211 37415 23247 37449
rect 23281 37415 23317 37449
rect 23351 37415 23387 37449
rect 23421 37415 23457 37449
rect 23491 37415 23527 37449
rect 23561 37415 23597 37449
rect 23631 37420 23711 37449
rect 23745 37420 23794 37454
rect 23828 37420 23877 37454
rect 23911 37420 23959 37454
rect 23993 37440 27021 37454
rect 23993 37420 24093 37440
rect 23631 37415 24093 37420
rect 22823 37406 24093 37415
rect 24127 37406 24162 37440
rect 24196 37406 24231 37440
rect 24265 37406 24300 37440
rect 24334 37406 24369 37440
rect 24403 37406 24438 37440
rect 24472 37406 24507 37440
rect 24541 37406 24576 37440
rect 24610 37406 24645 37440
rect 24679 37406 24714 37440
rect 24748 37406 24783 37440
rect 24817 37406 24852 37440
rect 24886 37406 24921 37440
rect 24955 37406 24990 37440
rect 25024 37406 25059 37440
rect 25093 37406 25127 37440
rect 25161 37406 25195 37440
rect 25229 37406 25263 37440
rect 25297 37406 25331 37440
rect 25365 37406 25399 37440
rect 25433 37406 25467 37440
rect 25501 37406 25535 37440
rect 25569 37406 25603 37440
rect 25637 37406 25671 37440
rect 25705 37406 25739 37440
rect 25773 37406 25807 37440
rect 25841 37406 25875 37440
rect 25909 37406 25943 37440
rect 25977 37406 26011 37440
rect 26045 37406 26079 37440
rect 26113 37406 26147 37440
rect 26181 37406 26215 37440
rect 26249 37406 26283 37440
rect 26317 37406 26351 37440
rect 26385 37406 26419 37440
rect 26453 37406 26487 37440
rect 26521 37406 26555 37440
rect 26589 37406 26623 37440
rect 26657 37406 26691 37440
rect 26725 37406 26759 37440
rect 26793 37406 26827 37440
rect 26861 37406 26895 37440
rect 26929 37406 26963 37440
rect 26997 37406 27021 37440
rect 22823 37381 27021 37406
rect 22823 37347 22827 37381
rect 22861 37347 22897 37381
rect 22931 37347 22967 37381
rect 23001 37347 23037 37381
rect 23071 37347 23107 37381
rect 23141 37347 23177 37381
rect 23211 37347 23247 37381
rect 23281 37347 23317 37381
rect 23351 37347 23387 37381
rect 23421 37347 23457 37381
rect 23491 37347 23527 37381
rect 23561 37347 23597 37381
rect 23631 37368 27021 37381
rect 23631 37347 23711 37368
rect 22823 37334 23711 37347
rect 23745 37334 23794 37368
rect 23828 37334 23877 37368
rect 23911 37334 23959 37368
rect 23993 37362 27021 37368
rect 23993 37334 24093 37362
rect 22823 37328 24093 37334
rect 24127 37328 24162 37362
rect 24196 37328 24231 37362
rect 24265 37328 24300 37362
rect 24334 37328 24369 37362
rect 24403 37328 24438 37362
rect 24472 37328 24507 37362
rect 24541 37328 24576 37362
rect 24610 37328 24645 37362
rect 24679 37328 24714 37362
rect 24748 37328 24783 37362
rect 24817 37328 24852 37362
rect 24886 37328 24921 37362
rect 24955 37328 24990 37362
rect 25024 37328 25059 37362
rect 25093 37328 25127 37362
rect 25161 37328 25195 37362
rect 25229 37328 25263 37362
rect 25297 37328 25331 37362
rect 25365 37328 25399 37362
rect 25433 37328 25467 37362
rect 25501 37328 25535 37362
rect 25569 37328 25603 37362
rect 25637 37328 25671 37362
rect 25705 37328 25739 37362
rect 25773 37328 25807 37362
rect 25841 37328 25875 37362
rect 25909 37328 25943 37362
rect 25977 37328 26011 37362
rect 26045 37328 26079 37362
rect 26113 37328 26147 37362
rect 26181 37328 26215 37362
rect 26249 37328 26283 37362
rect 26317 37328 26351 37362
rect 26385 37328 26419 37362
rect 26453 37328 26487 37362
rect 26521 37328 26555 37362
rect 26589 37328 26623 37362
rect 26657 37328 26691 37362
rect 26725 37328 26759 37362
rect 26793 37328 26827 37362
rect 26861 37328 26895 37362
rect 26929 37328 26963 37362
rect 26997 37328 27021 37362
rect 22823 37313 27021 37328
rect 22823 37279 22827 37313
rect 22861 37279 22897 37313
rect 22931 37279 22967 37313
rect 23001 37279 23037 37313
rect 23071 37279 23107 37313
rect 23141 37279 23177 37313
rect 23211 37279 23247 37313
rect 23281 37279 23317 37313
rect 23351 37279 23387 37313
rect 23421 37279 23457 37313
rect 23491 37279 23527 37313
rect 23561 37279 23597 37313
rect 23631 37284 27021 37313
rect 23631 37282 24093 37284
rect 23631 37279 23711 37282
rect 22823 37248 23711 37279
rect 23745 37248 23794 37282
rect 23828 37248 23877 37282
rect 23911 37248 23959 37282
rect 23993 37250 24093 37282
rect 24127 37250 24162 37284
rect 24196 37250 24231 37284
rect 24265 37250 24300 37284
rect 24334 37250 24369 37284
rect 24403 37250 24438 37284
rect 24472 37250 24507 37284
rect 24541 37250 24576 37284
rect 24610 37250 24645 37284
rect 24679 37250 24714 37284
rect 24748 37250 24783 37284
rect 24817 37250 24852 37284
rect 24886 37250 24921 37284
rect 24955 37250 24990 37284
rect 25024 37250 25059 37284
rect 25093 37250 25127 37284
rect 25161 37250 25195 37284
rect 25229 37250 25263 37284
rect 25297 37250 25331 37284
rect 25365 37250 25399 37284
rect 25433 37250 25467 37284
rect 25501 37250 25535 37284
rect 25569 37250 25603 37284
rect 25637 37250 25671 37284
rect 25705 37250 25739 37284
rect 25773 37250 25807 37284
rect 25841 37250 25875 37284
rect 25909 37250 25943 37284
rect 25977 37250 26011 37284
rect 26045 37250 26079 37284
rect 26113 37250 26147 37284
rect 26181 37250 26215 37284
rect 26249 37250 26283 37284
rect 26317 37250 26351 37284
rect 26385 37250 26419 37284
rect 26453 37250 26487 37284
rect 26521 37250 26555 37284
rect 26589 37250 26623 37284
rect 26657 37250 26691 37284
rect 26725 37250 26759 37284
rect 26793 37250 26827 37284
rect 26861 37250 26895 37284
rect 26929 37250 26963 37284
rect 26997 37250 27021 37284
rect 23993 37248 27021 37250
rect 22823 37247 27021 37248
rect 22823 37245 23635 37247
rect 22823 37211 22827 37245
rect 22861 37211 22897 37245
rect 22931 37211 22967 37245
rect 23001 37211 23037 37245
rect 23071 37211 23107 37245
rect 23141 37211 23177 37245
rect 23211 37211 23247 37245
rect 23281 37211 23317 37245
rect 23351 37211 23387 37245
rect 23421 37211 23457 37245
rect 23491 37211 23527 37245
rect 23561 37211 23597 37245
rect 23631 37211 23635 37245
rect 22823 37177 23635 37211
rect 22823 37143 22827 37177
rect 22861 37143 22897 37177
rect 22931 37143 22967 37177
rect 23001 37143 23037 37177
rect 23071 37143 23107 37177
rect 23141 37143 23177 37177
rect 23211 37143 23247 37177
rect 23281 37143 23317 37177
rect 23351 37143 23387 37177
rect 23421 37143 23457 37177
rect 23491 37143 23527 37177
rect 23561 37143 23597 37177
rect 23631 37143 23635 37177
rect 22823 37109 23635 37143
rect 22823 37075 22827 37109
rect 22861 37075 22897 37109
rect 22931 37075 22967 37109
rect 23001 37075 23037 37109
rect 23071 37075 23107 37109
rect 23141 37075 23177 37109
rect 23211 37075 23247 37109
rect 23281 37075 23317 37109
rect 23351 37075 23387 37109
rect 23421 37075 23457 37109
rect 23491 37075 23527 37109
rect 23561 37075 23597 37109
rect 23631 37075 23635 37109
rect 22823 37041 23635 37075
rect 22823 37007 22827 37041
rect 22861 37007 22897 37041
rect 22931 37007 22967 37041
rect 23001 37007 23037 37041
rect 23071 37007 23107 37041
rect 23141 37007 23177 37041
rect 23211 37007 23247 37041
rect 23281 37007 23317 37041
rect 23351 37007 23387 37041
rect 23421 37007 23457 37041
rect 23491 37007 23527 37041
rect 23561 37007 23597 37041
rect 23631 37007 23635 37041
rect 22823 36973 23635 37007
rect 22823 36939 22827 36973
rect 22861 36939 22897 36973
rect 22931 36939 22967 36973
rect 23001 36939 23037 36973
rect 23071 36939 23107 36973
rect 23141 36939 23177 36973
rect 23211 36939 23247 36973
rect 23281 36939 23317 36973
rect 23351 36939 23387 36973
rect 23421 36939 23457 36973
rect 23491 36939 23527 36973
rect 23561 36939 23597 36973
rect 23631 36939 23635 36973
rect 22823 36905 23635 36939
rect 22823 36871 22827 36905
rect 22861 36871 22897 36905
rect 22931 36871 22967 36905
rect 23001 36871 23037 36905
rect 23071 36871 23107 36905
rect 23141 36871 23177 36905
rect 23211 36871 23247 36905
rect 23281 36871 23317 36905
rect 23351 36871 23387 36905
rect 23421 36871 23457 36905
rect 23491 36871 23527 36905
rect 23561 36871 23597 36905
rect 23631 36871 23635 36905
rect 22823 36837 23635 36871
rect 22823 36803 22827 36837
rect 22861 36803 22897 36837
rect 22931 36803 22967 36837
rect 23001 36803 23037 36837
rect 23071 36803 23107 36837
rect 23141 36803 23177 36837
rect 23211 36803 23247 36837
rect 23281 36803 23317 36837
rect 23351 36803 23387 36837
rect 23421 36803 23457 36837
rect 23491 36803 23527 36837
rect 23561 36803 23597 36837
rect 23631 36803 23635 36837
rect 22823 36769 23635 36803
rect 22823 36735 22827 36769
rect 22861 36735 22897 36769
rect 22931 36735 22967 36769
rect 23001 36735 23037 36769
rect 23071 36735 23107 36769
rect 23141 36735 23177 36769
rect 23211 36735 23247 36769
rect 23281 36735 23317 36769
rect 23351 36735 23387 36769
rect 23421 36735 23457 36769
rect 23491 36735 23527 36769
rect 23561 36735 23597 36769
rect 23631 36735 23635 36769
rect 22823 36701 23635 36735
rect 22823 36667 22827 36701
rect 22861 36667 22897 36701
rect 22931 36667 22967 36701
rect 23001 36667 23037 36701
rect 23071 36667 23107 36701
rect 23141 36667 23177 36701
rect 23211 36667 23247 36701
rect 23281 36667 23317 36701
rect 23351 36667 23387 36701
rect 23421 36667 23457 36701
rect 23491 36667 23527 36701
rect 23561 36667 23597 36701
rect 23631 36667 23635 36701
rect 22823 36633 23635 36667
rect 22823 36599 22827 36633
rect 22861 36599 22897 36633
rect 22931 36599 22967 36633
rect 23001 36599 23037 36633
rect 23071 36599 23107 36633
rect 23141 36599 23177 36633
rect 23211 36599 23247 36633
rect 23281 36599 23317 36633
rect 23351 36599 23387 36633
rect 23421 36599 23457 36633
rect 23491 36599 23527 36633
rect 23561 36599 23597 36633
rect 23631 36599 23635 36633
rect 22823 36565 23635 36599
rect 22823 36531 22827 36565
rect 22861 36531 22897 36565
rect 22931 36531 22967 36565
rect 23001 36531 23037 36565
rect 23071 36531 23107 36565
rect 23141 36531 23177 36565
rect 23211 36531 23247 36565
rect 23281 36531 23317 36565
rect 23351 36531 23387 36565
rect 23421 36531 23457 36565
rect 23491 36531 23527 36565
rect 23561 36531 23597 36565
rect 23631 36531 23635 36565
rect 22823 36497 23635 36531
rect 22823 36463 22827 36497
rect 22861 36463 22897 36497
rect 22931 36463 22967 36497
rect 23001 36463 23037 36497
rect 23071 36463 23107 36497
rect 23141 36463 23177 36497
rect 23211 36463 23247 36497
rect 23281 36463 23317 36497
rect 23351 36463 23387 36497
rect 23421 36463 23457 36497
rect 23491 36463 23527 36497
rect 23561 36463 23597 36497
rect 23631 36463 23635 36497
rect 22823 36429 23635 36463
rect 22823 36395 22827 36429
rect 22861 36395 22897 36429
rect 22931 36395 22967 36429
rect 23001 36395 23037 36429
rect 23071 36395 23107 36429
rect 23141 36395 23177 36429
rect 23211 36395 23247 36429
rect 23281 36395 23317 36429
rect 23351 36395 23387 36429
rect 23421 36395 23457 36429
rect 23491 36395 23527 36429
rect 23561 36395 23597 36429
rect 23631 36395 23635 36429
rect 22823 36361 23635 36395
rect 22823 36327 22827 36361
rect 22861 36327 22897 36361
rect 22931 36327 22967 36361
rect 23001 36327 23037 36361
rect 23071 36327 23107 36361
rect 23141 36327 23177 36361
rect 23211 36327 23247 36361
rect 23281 36327 23317 36361
rect 23351 36327 23387 36361
rect 23421 36327 23457 36361
rect 23491 36327 23527 36361
rect 23561 36327 23597 36361
rect 23631 36327 23635 36361
rect 22823 36293 23635 36327
rect 22823 36259 22827 36293
rect 22861 36259 22897 36293
rect 22931 36259 22967 36293
rect 23001 36259 23037 36293
rect 23071 36259 23107 36293
rect 23141 36259 23177 36293
rect 23211 36259 23247 36293
rect 23281 36259 23317 36293
rect 23351 36259 23387 36293
rect 23421 36259 23457 36293
rect 23491 36259 23527 36293
rect 23561 36259 23597 36293
rect 23631 36259 23635 36293
rect 22823 36225 23635 36259
rect 22823 36191 22827 36225
rect 22861 36191 22897 36225
rect 22931 36191 22967 36225
rect 23001 36191 23037 36225
rect 23071 36191 23107 36225
rect 23141 36191 23177 36225
rect 23211 36191 23247 36225
rect 23281 36191 23317 36225
rect 23351 36191 23387 36225
rect 23421 36191 23457 36225
rect 23491 36191 23527 36225
rect 23561 36191 23597 36225
rect 23631 36191 23635 36225
rect 22823 36157 23635 36191
rect 22823 36123 22827 36157
rect 22861 36123 22897 36157
rect 22931 36123 22967 36157
rect 23001 36123 23037 36157
rect 23071 36123 23107 36157
rect 23141 36123 23177 36157
rect 23211 36123 23247 36157
rect 23281 36123 23317 36157
rect 23351 36123 23387 36157
rect 23421 36123 23457 36157
rect 23491 36123 23527 36157
rect 23561 36123 23597 36157
rect 23631 36123 23635 36157
rect 22823 36089 23635 36123
rect 22823 36055 22827 36089
rect 22861 36055 22897 36089
rect 22931 36055 22967 36089
rect 23001 36055 23037 36089
rect 23071 36055 23107 36089
rect 23141 36055 23177 36089
rect 23211 36055 23247 36089
rect 23281 36055 23317 36089
rect 23351 36055 23387 36089
rect 23421 36055 23457 36089
rect 23491 36055 23527 36089
rect 23561 36055 23597 36089
rect 23631 36055 23635 36089
rect 22823 36021 23635 36055
rect 22823 35987 22827 36021
rect 22861 35987 22897 36021
rect 22931 35987 22967 36021
rect 23001 35987 23037 36021
rect 23071 35987 23107 36021
rect 23141 35987 23177 36021
rect 23211 35987 23247 36021
rect 23281 35987 23317 36021
rect 23351 35987 23387 36021
rect 23421 35987 23457 36021
rect 23491 35987 23527 36021
rect 23561 35987 23597 36021
rect 23631 35987 23635 36021
rect 22823 35953 23635 35987
rect 22823 35919 22827 35953
rect 22861 35919 22897 35953
rect 22931 35919 22967 35953
rect 23001 35919 23037 35953
rect 23071 35919 23107 35953
rect 23141 35919 23177 35953
rect 23211 35919 23247 35953
rect 23281 35919 23317 35953
rect 23351 35919 23387 35953
rect 23421 35919 23457 35953
rect 23491 35919 23527 35953
rect 23561 35919 23597 35953
rect 23631 35919 23635 35953
rect 22823 35885 23635 35919
rect 22823 35851 22827 35885
rect 22861 35851 22897 35885
rect 22931 35851 22967 35885
rect 23001 35851 23037 35885
rect 23071 35851 23107 35885
rect 23141 35851 23177 35885
rect 23211 35851 23247 35885
rect 23281 35851 23317 35885
rect 23351 35851 23387 35885
rect 23421 35851 23457 35885
rect 23491 35851 23527 35885
rect 23561 35851 23597 35885
rect 23631 35851 23635 35885
rect 22823 35817 23635 35851
rect 22823 35783 22827 35817
rect 22861 35783 22897 35817
rect 22931 35783 22967 35817
rect 23001 35783 23037 35817
rect 23071 35783 23107 35817
rect 23141 35783 23177 35817
rect 23211 35783 23247 35817
rect 23281 35783 23317 35817
rect 23351 35783 23387 35817
rect 23421 35783 23457 35817
rect 23491 35783 23527 35817
rect 23561 35783 23597 35817
rect 23631 35783 23635 35817
rect 22823 35749 23635 35783
rect 22823 35715 22827 35749
rect 22861 35715 22897 35749
rect 22931 35715 22967 35749
rect 23001 35715 23037 35749
rect 23071 35715 23107 35749
rect 23141 35715 23177 35749
rect 23211 35715 23247 35749
rect 23281 35715 23317 35749
rect 23351 35715 23387 35749
rect 23421 35715 23457 35749
rect 23491 35715 23527 35749
rect 23561 35715 23597 35749
rect 23631 35715 23635 35749
rect 22823 35681 23635 35715
rect 22823 35647 22827 35681
rect 22861 35647 22897 35681
rect 22931 35647 22967 35681
rect 23001 35647 23037 35681
rect 23071 35647 23107 35681
rect 23141 35647 23177 35681
rect 23211 35647 23247 35681
rect 23281 35647 23317 35681
rect 23351 35647 23387 35681
rect 23421 35647 23457 35681
rect 23491 35647 23527 35681
rect 23561 35647 23597 35681
rect 23631 35647 23635 35681
rect 22823 35613 23635 35647
rect 22823 35579 22827 35613
rect 22861 35579 22897 35613
rect 22931 35579 22967 35613
rect 23001 35579 23037 35613
rect 23071 35579 23107 35613
rect 23141 35579 23177 35613
rect 23211 35579 23247 35613
rect 23281 35579 23317 35613
rect 23351 35579 23387 35613
rect 23421 35579 23457 35613
rect 23491 35579 23527 35613
rect 23561 35579 23597 35613
rect 23631 35579 23635 35613
rect 22823 35545 23635 35579
rect 22823 35511 22827 35545
rect 22861 35511 22897 35545
rect 22931 35511 22967 35545
rect 23001 35511 23037 35545
rect 23071 35511 23107 35545
rect 23141 35511 23177 35545
rect 23211 35511 23247 35545
rect 23281 35511 23317 35545
rect 23351 35511 23387 35545
rect 23421 35511 23457 35545
rect 23491 35511 23527 35545
rect 23561 35511 23597 35545
rect 23631 35511 23635 35545
rect 22823 35477 23635 35511
rect 22823 35443 22827 35477
rect 22861 35443 22897 35477
rect 22931 35443 22967 35477
rect 23001 35443 23037 35477
rect 23071 35443 23107 35477
rect 23141 35443 23177 35477
rect 23211 35443 23247 35477
rect 23281 35443 23317 35477
rect 23351 35443 23387 35477
rect 23421 35443 23457 35477
rect 23491 35443 23527 35477
rect 23561 35443 23597 35477
rect 23631 35443 23635 35477
rect 22823 35409 23635 35443
rect 22823 35375 22827 35409
rect 22861 35375 22897 35409
rect 22931 35375 22967 35409
rect 23001 35375 23037 35409
rect 23071 35375 23107 35409
rect 23141 35375 23177 35409
rect 23211 35375 23247 35409
rect 23281 35375 23317 35409
rect 23351 35375 23387 35409
rect 23421 35375 23457 35409
rect 23491 35375 23527 35409
rect 23561 35375 23597 35409
rect 23631 35375 23635 35409
rect 22823 35341 23635 35375
rect 22823 35307 22827 35341
rect 22861 35307 22897 35341
rect 22931 35307 22967 35341
rect 23001 35307 23037 35341
rect 23071 35307 23107 35341
rect 23141 35307 23177 35341
rect 23211 35307 23247 35341
rect 23281 35307 23317 35341
rect 23351 35307 23387 35341
rect 23421 35307 23457 35341
rect 23491 35307 23527 35341
rect 23561 35307 23597 35341
rect 23631 35307 23635 35341
rect 22823 35273 23635 35307
rect 22823 35239 22827 35273
rect 22861 35239 22897 35273
rect 22931 35239 22967 35273
rect 23001 35239 23037 35273
rect 23071 35239 23107 35273
rect 23141 35239 23177 35273
rect 23211 35239 23247 35273
rect 23281 35239 23317 35273
rect 23351 35239 23387 35273
rect 23421 35239 23457 35273
rect 23491 35239 23527 35273
rect 23561 35239 23597 35273
rect 23631 35239 23635 35273
rect 22823 35205 23635 35239
rect 22823 35171 22827 35205
rect 22861 35171 22897 35205
rect 22931 35171 22967 35205
rect 23001 35171 23037 35205
rect 23071 35171 23107 35205
rect 23141 35171 23177 35205
rect 23211 35171 23247 35205
rect 23281 35171 23317 35205
rect 23351 35171 23387 35205
rect 23421 35171 23457 35205
rect 23491 35171 23527 35205
rect 23561 35171 23597 35205
rect 23631 35171 23635 35205
rect 22823 35137 23635 35171
rect 22823 35103 22827 35137
rect 22861 35103 22897 35137
rect 22931 35103 22967 35137
rect 23001 35103 23037 35137
rect 23071 35103 23107 35137
rect 23141 35103 23177 35137
rect 23211 35103 23247 35137
rect 23281 35103 23317 35137
rect 23351 35103 23387 35137
rect 23421 35103 23457 35137
rect 23491 35103 23527 35137
rect 23561 35103 23597 35137
rect 23631 35103 23635 35137
rect 22823 35069 23635 35103
rect 22823 35035 22827 35069
rect 22861 35035 22897 35069
rect 22931 35035 22967 35069
rect 23001 35035 23037 35069
rect 23071 35035 23107 35069
rect 23141 35035 23177 35069
rect 23211 35035 23247 35069
rect 23281 35035 23317 35069
rect 23351 35035 23387 35069
rect 23421 35035 23457 35069
rect 23491 35035 23527 35069
rect 23561 35035 23597 35069
rect 23631 35035 23635 35069
rect 22823 35001 23635 35035
rect 22823 34967 22827 35001
rect 22861 34967 22897 35001
rect 22931 34967 22967 35001
rect 23001 34967 23037 35001
rect 23071 34967 23107 35001
rect 23141 34967 23177 35001
rect 23211 34967 23247 35001
rect 23281 34967 23317 35001
rect 23351 34967 23387 35001
rect 23421 34967 23457 35001
rect 23491 34967 23527 35001
rect 23561 34967 23597 35001
rect 23631 34967 23635 35001
rect 22823 34933 23635 34967
rect 22823 34899 22827 34933
rect 22861 34899 22897 34933
rect 22931 34899 22967 34933
rect 23001 34899 23037 34933
rect 23071 34899 23107 34933
rect 23141 34899 23177 34933
rect 23211 34899 23247 34933
rect 23281 34899 23317 34933
rect 23351 34899 23387 34933
rect 23421 34899 23457 34933
rect 23491 34899 23527 34933
rect 23561 34899 23597 34933
rect 23631 34899 23635 34933
rect 22823 34865 23635 34899
rect 22823 34831 22827 34865
rect 22861 34831 22897 34865
rect 22931 34831 22967 34865
rect 23001 34831 23037 34865
rect 23071 34831 23107 34865
rect 23141 34831 23177 34865
rect 23211 34831 23247 34865
rect 23281 34831 23317 34865
rect 23351 34831 23387 34865
rect 23421 34831 23457 34865
rect 23491 34831 23527 34865
rect 23561 34831 23597 34865
rect 23631 34831 23635 34865
rect 22823 34797 23635 34831
rect 22823 34763 22827 34797
rect 22861 34763 22897 34797
rect 22931 34763 22967 34797
rect 23001 34763 23037 34797
rect 23071 34763 23107 34797
rect 23141 34763 23177 34797
rect 23211 34763 23247 34797
rect 23281 34763 23317 34797
rect 23351 34763 23387 34797
rect 23421 34763 23457 34797
rect 23491 34763 23527 34797
rect 23561 34763 23597 34797
rect 23631 34763 23635 34797
rect 22823 34729 23635 34763
rect 22823 34695 22827 34729
rect 22861 34695 22897 34729
rect 22931 34695 22967 34729
rect 23001 34695 23037 34729
rect 23071 34695 23107 34729
rect 23141 34695 23177 34729
rect 23211 34695 23247 34729
rect 23281 34695 23317 34729
rect 23351 34695 23387 34729
rect 23421 34695 23457 34729
rect 23491 34695 23527 34729
rect 23561 34695 23597 34729
rect 23631 34695 23635 34729
rect 22823 34661 23635 34695
rect 22823 34627 22827 34661
rect 22861 34627 22897 34661
rect 22931 34627 22967 34661
rect 23001 34627 23037 34661
rect 23071 34627 23107 34661
rect 23141 34627 23177 34661
rect 23211 34627 23247 34661
rect 23281 34627 23317 34661
rect 23351 34627 23387 34661
rect 23421 34627 23457 34661
rect 23491 34627 23527 34661
rect 23561 34627 23597 34661
rect 23631 34627 23635 34661
rect 22823 34593 23635 34627
rect 22823 34559 22827 34593
rect 22861 34559 22897 34593
rect 22931 34559 22967 34593
rect 23001 34559 23037 34593
rect 23071 34559 23107 34593
rect 23141 34559 23177 34593
rect 23211 34559 23247 34593
rect 23281 34559 23317 34593
rect 23351 34559 23387 34593
rect 23421 34559 23457 34593
rect 23491 34559 23527 34593
rect 23561 34559 23597 34593
rect 23631 34559 23635 34593
rect 22823 34525 23635 34559
rect 22823 34491 22827 34525
rect 22861 34491 22897 34525
rect 22931 34491 22967 34525
rect 23001 34491 23037 34525
rect 23071 34491 23107 34525
rect 23141 34491 23177 34525
rect 23211 34491 23247 34525
rect 23281 34491 23317 34525
rect 23351 34491 23387 34525
rect 23421 34491 23457 34525
rect 23491 34491 23527 34525
rect 23561 34491 23597 34525
rect 23631 34491 23635 34525
rect 22823 34457 23635 34491
rect 22823 34423 22827 34457
rect 22861 34423 22897 34457
rect 22931 34423 22967 34457
rect 23001 34423 23037 34457
rect 23071 34423 23107 34457
rect 23141 34423 23177 34457
rect 23211 34423 23247 34457
rect 23281 34423 23317 34457
rect 23351 34423 23387 34457
rect 23421 34423 23457 34457
rect 23491 34423 23527 34457
rect 23561 34423 23597 34457
rect 23631 34423 23635 34457
rect 22823 34389 23635 34423
rect 22823 34355 22827 34389
rect 22861 34355 22897 34389
rect 22931 34355 22967 34389
rect 23001 34355 23037 34389
rect 23071 34355 23107 34389
rect 23141 34355 23177 34389
rect 23211 34355 23247 34389
rect 23281 34355 23317 34389
rect 23351 34355 23387 34389
rect 23421 34355 23457 34389
rect 23491 34355 23527 34389
rect 23561 34355 23597 34389
rect 23631 34355 23635 34389
rect 22823 34321 23635 34355
rect 22823 34287 22827 34321
rect 22861 34287 22897 34321
rect 22931 34287 22967 34321
rect 23001 34287 23037 34321
rect 23071 34287 23107 34321
rect 23141 34287 23177 34321
rect 23211 34287 23247 34321
rect 23281 34287 23317 34321
rect 23351 34287 23387 34321
rect 23421 34287 23457 34321
rect 23491 34287 23527 34321
rect 23561 34287 23597 34321
rect 23631 34287 23635 34321
rect 22823 34253 23635 34287
rect 22823 34219 22827 34253
rect 22861 34219 22897 34253
rect 22931 34219 22967 34253
rect 23001 34219 23037 34253
rect 23071 34219 23107 34253
rect 23141 34219 23177 34253
rect 23211 34219 23247 34253
rect 23281 34219 23317 34253
rect 23351 34219 23387 34253
rect 23421 34219 23457 34253
rect 23491 34219 23527 34253
rect 23561 34219 23597 34253
rect 23631 34219 23635 34253
rect 22823 34185 23635 34219
rect 22823 34151 22827 34185
rect 22861 34151 22897 34185
rect 22931 34151 22967 34185
rect 23001 34151 23037 34185
rect 23071 34151 23107 34185
rect 23141 34151 23177 34185
rect 23211 34151 23247 34185
rect 23281 34151 23317 34185
rect 23351 34151 23387 34185
rect 23421 34151 23457 34185
rect 23491 34151 23527 34185
rect 23561 34151 23597 34185
rect 23631 34151 23635 34185
rect 22823 34117 23635 34151
rect 22823 34083 22827 34117
rect 22861 34083 22897 34117
rect 22931 34083 22967 34117
rect 23001 34083 23037 34117
rect 23071 34083 23107 34117
rect 23141 34083 23177 34117
rect 23211 34083 23247 34117
rect 23281 34083 23317 34117
rect 23351 34083 23387 34117
rect 23421 34083 23457 34117
rect 23491 34083 23527 34117
rect 23561 34083 23597 34117
rect 23631 34083 23635 34117
rect 22823 34049 23635 34083
rect 22823 34015 22827 34049
rect 22861 34015 22897 34049
rect 22931 34015 22967 34049
rect 23001 34015 23037 34049
rect 23071 34015 23107 34049
rect 23141 34015 23177 34049
rect 23211 34015 23247 34049
rect 23281 34015 23317 34049
rect 23351 34015 23387 34049
rect 23421 34015 23457 34049
rect 23491 34015 23527 34049
rect 23561 34015 23597 34049
rect 23631 34015 23635 34049
rect 22823 33981 23635 34015
rect 22823 33947 22827 33981
rect 22861 33947 22897 33981
rect 22931 33947 22967 33981
rect 23001 33947 23037 33981
rect 23071 33947 23107 33981
rect 23141 33947 23177 33981
rect 23211 33947 23247 33981
rect 23281 33947 23317 33981
rect 23351 33947 23387 33981
rect 23421 33947 23457 33981
rect 23491 33947 23527 33981
rect 23561 33947 23597 33981
rect 23631 33947 23635 33981
rect 22823 33913 23635 33947
rect 22823 33879 22827 33913
rect 22861 33879 22897 33913
rect 22931 33879 22967 33913
rect 23001 33879 23037 33913
rect 23071 33879 23107 33913
rect 23141 33879 23177 33913
rect 23211 33879 23247 33913
rect 23281 33879 23317 33913
rect 23351 33879 23387 33913
rect 23421 33879 23457 33913
rect 23491 33879 23527 33913
rect 23561 33879 23597 33913
rect 23631 33879 23635 33913
rect 22823 33845 23635 33879
rect 22823 33811 22827 33845
rect 22861 33811 22897 33845
rect 22931 33811 22967 33845
rect 23001 33811 23037 33845
rect 23071 33811 23107 33845
rect 23141 33811 23177 33845
rect 23211 33811 23247 33845
rect 23281 33811 23317 33845
rect 23351 33811 23387 33845
rect 23421 33811 23457 33845
rect 23491 33811 23527 33845
rect 23561 33811 23597 33845
rect 23631 33811 23635 33845
rect 22823 33777 23635 33811
rect 22823 33743 22827 33777
rect 22861 33743 22897 33777
rect 22931 33743 22967 33777
rect 23001 33743 23037 33777
rect 23071 33743 23107 33777
rect 23141 33743 23177 33777
rect 23211 33743 23247 33777
rect 23281 33743 23317 33777
rect 23351 33743 23387 33777
rect 23421 33743 23457 33777
rect 23491 33743 23527 33777
rect 23561 33743 23597 33777
rect 23631 33743 23635 33777
rect 22823 33709 23635 33743
rect 22823 33675 22827 33709
rect 22861 33675 22897 33709
rect 22931 33675 22967 33709
rect 23001 33675 23037 33709
rect 23071 33675 23107 33709
rect 23141 33675 23177 33709
rect 23211 33675 23247 33709
rect 23281 33675 23317 33709
rect 23351 33675 23387 33709
rect 23421 33675 23457 33709
rect 23491 33675 23527 33709
rect 23561 33675 23597 33709
rect 23631 33675 23635 33709
rect 22823 33641 23635 33675
rect 22823 33607 22827 33641
rect 22861 33607 22897 33641
rect 22931 33607 22967 33641
rect 23001 33607 23037 33641
rect 23071 33607 23107 33641
rect 23141 33607 23177 33641
rect 23211 33607 23247 33641
rect 23281 33607 23317 33641
rect 23351 33607 23387 33641
rect 23421 33607 23457 33641
rect 23491 33607 23527 33641
rect 23561 33607 23597 33641
rect 23631 33607 23635 33641
rect 22823 33573 23635 33607
rect 22823 33539 22827 33573
rect 22861 33539 22897 33573
rect 22931 33539 22967 33573
rect 23001 33539 23037 33573
rect 23071 33539 23107 33573
rect 23141 33539 23177 33573
rect 23211 33539 23247 33573
rect 23281 33539 23317 33573
rect 23351 33539 23387 33573
rect 23421 33539 23457 33573
rect 23491 33539 23527 33573
rect 23561 33539 23597 33573
rect 23631 33539 23635 33573
rect 22823 33505 23635 33539
rect 22823 33471 22827 33505
rect 22861 33471 22897 33505
rect 22931 33471 22967 33505
rect 23001 33471 23037 33505
rect 23071 33471 23107 33505
rect 23141 33471 23177 33505
rect 23211 33471 23247 33505
rect 23281 33471 23317 33505
rect 23351 33471 23387 33505
rect 23421 33471 23457 33505
rect 23491 33471 23527 33505
rect 23561 33471 23597 33505
rect 23631 33471 23635 33505
rect 22823 33437 23635 33471
rect 22823 33403 22827 33437
rect 22861 33403 22897 33437
rect 22931 33403 22967 33437
rect 23001 33403 23037 33437
rect 23071 33403 23107 33437
rect 23141 33403 23177 33437
rect 23211 33403 23247 33437
rect 23281 33403 23317 33437
rect 23351 33403 23387 33437
rect 23421 33403 23457 33437
rect 23491 33403 23527 33437
rect 23561 33403 23597 33437
rect 23631 33403 23635 33437
rect 22823 33369 23635 33403
rect 22823 33335 22827 33369
rect 22861 33335 22897 33369
rect 22931 33335 22967 33369
rect 23001 33335 23037 33369
rect 23071 33335 23107 33369
rect 23141 33335 23177 33369
rect 23211 33335 23247 33369
rect 23281 33335 23317 33369
rect 23351 33335 23387 33369
rect 23421 33335 23457 33369
rect 23491 33335 23527 33369
rect 23561 33335 23597 33369
rect 23631 33335 23635 33369
rect 269 33281 339 33316
rect 269 33247 278 33281
rect 312 33247 339 33281
rect 269 33212 339 33247
rect 269 33178 278 33212
rect 312 33178 339 33212
rect 269 33143 339 33178
rect 269 33109 278 33143
rect 312 33109 339 33143
rect 269 33074 339 33109
rect 269 33040 278 33074
rect 312 33040 339 33074
rect 269 33005 339 33040
rect 269 32971 278 33005
rect 312 32971 339 33005
rect 269 32936 339 32971
rect 269 32902 278 32936
rect 312 32902 339 32936
rect 269 32867 339 32902
rect 269 32833 278 32867
rect 312 32833 339 32867
rect 269 32798 339 32833
rect 269 32764 278 32798
rect 312 32764 339 32798
rect 269 32729 339 32764
rect 269 32695 278 32729
rect 312 32695 339 32729
rect 269 32660 339 32695
rect 269 32626 278 32660
rect 312 32626 339 32660
rect 269 32591 339 32626
rect 269 32557 278 32591
rect 312 32557 339 32591
rect 269 32522 339 32557
rect 269 32488 278 32522
rect 312 32488 339 32522
rect 269 32453 339 32488
rect 269 32419 278 32453
rect 312 32419 339 32453
rect 269 32384 339 32419
rect 269 32350 278 32384
rect 312 32350 339 32384
rect 269 32316 339 32350
rect 18022 33307 18442 33331
rect 18022 33273 18025 33307
rect 18059 33273 18101 33307
rect 18135 33273 18177 33307
rect 18211 33273 18253 33307
rect 18287 33273 18329 33307
rect 18363 33273 18405 33307
rect 18439 33273 18442 33307
rect 18022 33239 18442 33273
rect 18022 33205 18025 33239
rect 18059 33205 18101 33239
rect 18135 33205 18177 33239
rect 18211 33205 18253 33239
rect 18287 33205 18329 33239
rect 18363 33205 18405 33239
rect 18439 33205 18442 33239
rect 18022 33171 18442 33205
rect 18022 33137 18025 33171
rect 18059 33137 18101 33171
rect 18135 33137 18177 33171
rect 18211 33137 18253 33171
rect 18287 33137 18329 33171
rect 18363 33137 18405 33171
rect 18439 33137 18442 33171
rect 18022 33103 18442 33137
rect 18022 33069 18025 33103
rect 18059 33069 18101 33103
rect 18135 33069 18177 33103
rect 18211 33069 18253 33103
rect 18287 33069 18329 33103
rect 18363 33069 18405 33103
rect 18439 33069 18442 33103
rect 18022 33035 18442 33069
rect 18022 33001 18025 33035
rect 18059 33001 18101 33035
rect 18135 33001 18177 33035
rect 18211 33001 18253 33035
rect 18287 33001 18329 33035
rect 18363 33001 18405 33035
rect 18439 33001 18442 33035
rect 18022 32967 18442 33001
rect 18022 32933 18025 32967
rect 18059 32933 18101 32967
rect 18135 32933 18177 32967
rect 18211 32933 18253 32967
rect 18287 32933 18329 32967
rect 18363 32933 18405 32967
rect 18439 32933 18442 32967
rect 18022 32899 18442 32933
rect 18022 32865 18025 32899
rect 18059 32865 18101 32899
rect 18135 32865 18177 32899
rect 18211 32865 18253 32899
rect 18287 32865 18329 32899
rect 18363 32865 18405 32899
rect 18439 32865 18442 32899
rect 18022 32831 18442 32865
rect 18022 32797 18025 32831
rect 18059 32797 18101 32831
rect 18135 32797 18177 32831
rect 18211 32797 18253 32831
rect 18287 32797 18329 32831
rect 18363 32797 18405 32831
rect 18439 32797 18442 32831
rect 18022 32763 18442 32797
rect 18022 32729 18025 32763
rect 18059 32729 18101 32763
rect 18135 32729 18177 32763
rect 18211 32729 18253 32763
rect 18287 32729 18329 32763
rect 18363 32729 18405 32763
rect 18439 32729 18442 32763
rect 18022 32695 18442 32729
rect 18022 32661 18025 32695
rect 18059 32661 18101 32695
rect 18135 32661 18177 32695
rect 18211 32661 18253 32695
rect 18287 32661 18329 32695
rect 18363 32661 18405 32695
rect 18439 32661 18442 32695
rect 18022 32627 18442 32661
rect 18022 32593 18025 32627
rect 18059 32593 18101 32627
rect 18135 32593 18177 32627
rect 18211 32593 18253 32627
rect 18287 32593 18329 32627
rect 18363 32593 18405 32627
rect 18439 32593 18442 32627
rect 18022 32559 18442 32593
rect 18022 32525 18025 32559
rect 18059 32525 18101 32559
rect 18135 32525 18177 32559
rect 18211 32525 18253 32559
rect 18287 32525 18329 32559
rect 18363 32525 18405 32559
rect 18439 32525 18442 32559
rect 18022 32491 18442 32525
rect 18022 32457 18025 32491
rect 18059 32457 18101 32491
rect 18135 32457 18177 32491
rect 18211 32457 18253 32491
rect 18287 32457 18329 32491
rect 18363 32457 18405 32491
rect 18439 32457 18442 32491
rect 18022 32423 18442 32457
rect 18022 32389 18025 32423
rect 18059 32389 18101 32423
rect 18135 32389 18177 32423
rect 18211 32389 18253 32423
rect 18287 32389 18329 32423
rect 18363 32389 18405 32423
rect 18439 32389 18442 32423
rect 18022 32355 18442 32389
rect 18022 32321 18025 32355
rect 18059 32321 18101 32355
rect 18135 32321 18177 32355
rect 18211 32321 18253 32355
rect 18287 32321 18329 32355
rect 18363 32321 18405 32355
rect 18439 32321 18442 32355
rect 269 32315 912 32316
rect 269 32281 278 32315
rect 312 32282 912 32315
rect 312 32281 368 32282
rect 269 32248 368 32281
rect 402 32248 440 32282
rect 474 32248 512 32282
rect 546 32248 584 32282
rect 618 32248 656 32282
rect 690 32248 728 32282
rect 762 32248 800 32282
rect 834 32248 872 32282
rect 906 32248 912 32282
rect 269 32246 912 32248
rect 269 32212 278 32246
rect 312 32212 912 32246
rect 269 32206 912 32212
rect 269 32177 368 32206
rect 269 32143 278 32177
rect 312 32172 368 32177
rect 402 32172 440 32206
rect 474 32172 512 32206
rect 546 32172 584 32206
rect 618 32172 656 32206
rect 690 32172 728 32206
rect 762 32172 800 32206
rect 834 32172 872 32206
rect 906 32172 912 32206
rect 312 32143 912 32172
rect 269 32130 912 32143
rect 269 32108 368 32130
rect 269 32074 278 32108
rect 312 32096 368 32108
rect 402 32096 440 32130
rect 474 32096 512 32130
rect 546 32096 584 32130
rect 618 32096 656 32130
rect 690 32096 728 32130
rect 762 32096 800 32130
rect 834 32096 872 32130
rect 906 32096 912 32130
rect 312 32074 912 32096
rect 269 32054 912 32074
rect 269 32039 368 32054
rect 269 32005 278 32039
rect 312 32020 368 32039
rect 402 32020 440 32054
rect 474 32020 512 32054
rect 546 32020 584 32054
rect 618 32020 656 32054
rect 690 32020 728 32054
rect 762 32020 800 32054
rect 834 32020 872 32054
rect 906 32020 912 32054
rect 312 32005 912 32020
rect 269 31978 912 32005
rect 269 31970 368 31978
rect 269 31936 278 31970
rect 312 31944 368 31970
rect 402 31944 440 31978
rect 474 31944 512 31978
rect 546 31944 584 31978
rect 618 31944 656 31978
rect 690 31944 728 31978
rect 762 31944 800 31978
rect 834 31944 872 31978
rect 906 31944 912 31978
rect 312 31936 912 31944
rect 269 31902 912 31936
rect 269 31901 368 31902
rect 269 31867 278 31901
rect 312 31868 368 31901
rect 402 31868 440 31902
rect 474 31868 512 31902
rect 546 31868 584 31902
rect 618 31868 656 31902
rect 690 31868 728 31902
rect 762 31868 800 31902
rect 834 31868 872 31902
rect 906 31868 912 31902
rect 312 31867 912 31868
rect 269 31832 912 31867
rect 269 31798 278 31832
rect 312 31825 912 31832
rect 312 31798 368 31825
rect 269 31791 368 31798
rect 402 31791 440 31825
rect 474 31791 512 31825
rect 546 31791 584 31825
rect 618 31791 656 31825
rect 690 31791 728 31825
rect 762 31791 800 31825
rect 834 31791 872 31825
rect 906 31791 912 31825
rect 269 31763 912 31791
rect 269 31729 278 31763
rect 312 31729 912 31763
rect 269 31705 912 31729
rect 18022 32287 18442 32321
rect 18022 32253 18025 32287
rect 18059 32253 18101 32287
rect 18135 32253 18177 32287
rect 18211 32253 18253 32287
rect 18287 32253 18329 32287
rect 18363 32253 18405 32287
rect 18439 32253 18442 32287
rect 18022 32219 18442 32253
rect 18022 32185 18025 32219
rect 18059 32185 18101 32219
rect 18135 32185 18177 32219
rect 18211 32185 18253 32219
rect 18287 32185 18329 32219
rect 18363 32185 18405 32219
rect 18439 32185 18442 32219
rect 18022 32151 18442 32185
rect 18022 32117 18025 32151
rect 18059 32117 18101 32151
rect 18135 32117 18177 32151
rect 18211 32117 18253 32151
rect 18287 32117 18329 32151
rect 18363 32117 18405 32151
rect 18439 32117 18442 32151
rect 18022 32083 18442 32117
rect 18022 32049 18025 32083
rect 18059 32049 18101 32083
rect 18135 32049 18177 32083
rect 18211 32049 18253 32083
rect 18287 32049 18329 32083
rect 18363 32049 18405 32083
rect 18439 32049 18442 32083
rect 18022 32015 18442 32049
rect 18022 31981 18025 32015
rect 18059 31981 18101 32015
rect 18135 31981 18177 32015
rect 18211 31981 18253 32015
rect 18287 31981 18329 32015
rect 18363 31981 18405 32015
rect 18439 31981 18442 32015
rect 18022 31947 18442 31981
rect 18022 31913 18025 31947
rect 18059 31913 18101 31947
rect 18135 31913 18177 31947
rect 18211 31913 18253 31947
rect 18287 31913 18329 31947
rect 18363 31913 18405 31947
rect 18439 31913 18442 31947
rect 18022 31879 18442 31913
rect 18022 31845 18025 31879
rect 18059 31845 18101 31879
rect 18135 31845 18177 31879
rect 18211 31845 18253 31879
rect 18287 31845 18329 31879
rect 18363 31845 18405 31879
rect 18439 31845 18442 31879
rect 18022 31811 18442 31845
rect 18022 31777 18025 31811
rect 18059 31777 18101 31811
rect 18135 31777 18177 31811
rect 18211 31777 18253 31811
rect 18287 31777 18329 31811
rect 18363 31777 18405 31811
rect 18439 31777 18442 31811
rect 18022 31743 18442 31777
rect 18022 31709 18025 31743
rect 18059 31709 18101 31743
rect 18135 31709 18177 31743
rect 18211 31709 18253 31743
rect 18287 31709 18329 31743
rect 18363 31709 18405 31743
rect 18439 31709 18442 31743
rect 279 31645 332 31705
rect 1025 31671 1313 31705
rect 1025 31645 1051 31671
rect 279 23829 306 31645
rect 280 23803 306 23829
rect 324 23829 332 31645
rect 999 31637 1051 31645
rect 1085 31637 1127 31671
rect 1161 31637 1203 31671
rect 1237 31637 1279 31671
rect 999 31603 1313 31637
rect 999 31569 1051 31603
rect 1085 31569 1127 31603
rect 1161 31569 1203 31603
rect 1237 31569 1279 31603
rect 999 31535 1313 31569
rect 999 31501 1051 31535
rect 1085 31501 1127 31535
rect 1161 31501 1203 31535
rect 1237 31501 1279 31535
rect 999 31467 1313 31501
rect 999 31433 1051 31467
rect 1085 31433 1127 31467
rect 1161 31433 1203 31467
rect 1237 31433 1279 31467
rect 999 31399 1313 31433
rect 999 31365 1051 31399
rect 1085 31365 1127 31399
rect 1161 31365 1203 31399
rect 1237 31365 1279 31399
rect 999 31331 1313 31365
rect 999 31297 1051 31331
rect 1085 31297 1127 31331
rect 1161 31297 1203 31331
rect 1237 31297 1279 31331
rect 999 31263 1313 31297
rect 999 31229 1051 31263
rect 1085 31229 1127 31263
rect 1161 31229 1203 31263
rect 1237 31229 1279 31263
rect 999 31195 1313 31229
rect 999 31161 1051 31195
rect 1085 31161 1127 31195
rect 1161 31161 1203 31195
rect 1237 31161 1279 31195
rect 999 31127 1313 31161
rect 999 31093 1051 31127
rect 1085 31093 1127 31127
rect 1161 31093 1203 31127
rect 1237 31093 1279 31127
rect 999 31059 1313 31093
rect 999 31025 1051 31059
rect 1085 31025 1127 31059
rect 1161 31025 1203 31059
rect 1237 31025 1279 31059
rect 999 30991 1313 31025
rect 999 30957 1051 30991
rect 1085 30957 1127 30991
rect 1161 30957 1203 30991
rect 1237 30957 1279 30991
rect 999 30923 1313 30957
rect 999 30889 1051 30923
rect 1085 30889 1127 30923
rect 1161 30889 1203 30923
rect 1237 30889 1279 30923
rect 999 30855 1313 30889
rect 999 30821 1051 30855
rect 1085 30821 1127 30855
rect 1161 30821 1203 30855
rect 1237 30821 1279 30855
rect 999 30787 1313 30821
rect 999 30753 1051 30787
rect 1085 30753 1127 30787
rect 1161 30753 1203 30787
rect 1237 30753 1279 30787
rect 999 30719 1313 30753
rect 999 30685 1051 30719
rect 1085 30685 1127 30719
rect 1161 30685 1203 30719
rect 1237 30685 1279 30719
rect 999 30651 1313 30685
rect 999 30617 1051 30651
rect 1085 30617 1127 30651
rect 1161 30617 1203 30651
rect 1237 30617 1279 30651
rect 999 30583 1313 30617
rect 999 30549 1051 30583
rect 1085 30549 1127 30583
rect 1161 30549 1203 30583
rect 1237 30549 1279 30583
rect 999 30515 1313 30549
rect 999 30481 1051 30515
rect 1085 30481 1127 30515
rect 1161 30481 1203 30515
rect 1237 30481 1279 30515
rect 999 30447 1313 30481
rect 999 30413 1051 30447
rect 1085 30413 1127 30447
rect 1161 30413 1203 30447
rect 1237 30413 1279 30447
rect 999 30379 1313 30413
rect 999 30345 1051 30379
rect 1085 30345 1127 30379
rect 1161 30345 1203 30379
rect 1237 30345 1279 30379
rect 999 30311 1313 30345
rect 999 30277 1051 30311
rect 1085 30277 1127 30311
rect 1161 30277 1203 30311
rect 1237 30277 1279 30311
rect 999 30243 1313 30277
rect 999 30209 1051 30243
rect 1085 30209 1127 30243
rect 1161 30209 1203 30243
rect 1237 30209 1279 30243
rect 999 30175 1313 30209
rect 999 30141 1051 30175
rect 1085 30141 1127 30175
rect 1161 30141 1203 30175
rect 1237 30141 1279 30175
rect 999 30107 1313 30141
rect 999 30073 1051 30107
rect 1085 30073 1127 30107
rect 1161 30073 1203 30107
rect 1237 30073 1279 30107
rect 999 30039 1313 30073
rect 999 30005 1051 30039
rect 1085 30005 1127 30039
rect 1161 30005 1203 30039
rect 1237 30005 1279 30039
rect 999 29971 1313 30005
rect 999 29937 1051 29971
rect 1085 29937 1127 29971
rect 1161 29937 1203 29971
rect 1237 29937 1279 29971
rect 999 29903 1313 29937
rect 999 29869 1051 29903
rect 1085 29869 1127 29903
rect 1161 29869 1203 29903
rect 1237 29869 1279 29903
rect 999 29835 1313 29869
rect 999 29801 1051 29835
rect 1085 29801 1127 29835
rect 1161 29801 1203 29835
rect 1237 29801 1279 29835
rect 999 29767 1313 29801
rect 999 29733 1051 29767
rect 1085 29733 1127 29767
rect 1161 29733 1203 29767
rect 1237 29733 1279 29767
rect 999 29699 1313 29733
rect 999 29665 1051 29699
rect 1085 29665 1127 29699
rect 1161 29665 1203 29699
rect 1237 29665 1279 29699
rect 999 29631 1313 29665
rect 999 29597 1051 29631
rect 1085 29597 1127 29631
rect 1161 29597 1203 29631
rect 1237 29597 1279 29631
rect 999 29563 1313 29597
rect 999 29529 1051 29563
rect 1085 29529 1127 29563
rect 1161 29529 1203 29563
rect 1237 29529 1279 29563
rect 999 29495 1313 29529
rect 999 29461 1051 29495
rect 1085 29461 1127 29495
rect 1161 29461 1203 29495
rect 1237 29461 1279 29495
rect 999 29427 1313 29461
rect 999 29393 1051 29427
rect 1085 29393 1127 29427
rect 1161 29393 1203 29427
rect 1237 29393 1279 29427
rect 999 29359 1313 29393
rect 999 29325 1051 29359
rect 1085 29325 1127 29359
rect 1161 29325 1203 29359
rect 1237 29325 1279 29359
rect 999 29291 1313 29325
rect 999 29257 1051 29291
rect 1085 29257 1127 29291
rect 1161 29257 1203 29291
rect 1237 29257 1279 29291
rect 999 29223 1313 29257
rect 999 29189 1051 29223
rect 1085 29189 1127 29223
rect 1161 29189 1203 29223
rect 1237 29189 1279 29223
rect 999 29155 1313 29189
rect 999 29121 1051 29155
rect 1085 29121 1127 29155
rect 1161 29121 1203 29155
rect 1237 29121 1279 29155
rect 999 29086 1313 29121
rect 999 29052 1051 29086
rect 1085 29052 1127 29086
rect 1161 29052 1203 29086
rect 1237 29052 1279 29086
rect 999 29017 1313 29052
rect 999 28983 1051 29017
rect 1085 28983 1127 29017
rect 1161 28983 1203 29017
rect 1237 28983 1279 29017
rect 999 28948 1313 28983
rect 999 28914 1051 28948
rect 1085 28914 1127 28948
rect 1161 28914 1203 28948
rect 1237 28914 1279 28948
rect 999 28879 1313 28914
rect 999 28845 1051 28879
rect 1085 28845 1127 28879
rect 1161 28845 1203 28879
rect 1237 28845 1279 28879
rect 999 28810 1313 28845
rect 999 28776 1051 28810
rect 1085 28776 1127 28810
rect 1161 28776 1203 28810
rect 1237 28776 1279 28810
rect 999 28741 1313 28776
rect 999 28707 1051 28741
rect 1085 28707 1127 28741
rect 1161 28707 1203 28741
rect 1237 28707 1279 28741
rect 999 28672 1313 28707
rect 999 28638 1051 28672
rect 1085 28638 1127 28672
rect 1161 28638 1203 28672
rect 1237 28638 1279 28672
rect 999 28603 1313 28638
rect 999 28569 1051 28603
rect 1085 28569 1127 28603
rect 1161 28569 1203 28603
rect 1237 28569 1279 28603
rect 999 28534 1313 28569
rect 999 28500 1051 28534
rect 1085 28500 1127 28534
rect 1161 28500 1203 28534
rect 1237 28500 1279 28534
rect 999 28465 1313 28500
rect 999 28431 1051 28465
rect 1085 28431 1127 28465
rect 1161 28431 1203 28465
rect 1237 28431 1279 28465
rect 999 28396 1313 28431
rect 999 28362 1051 28396
rect 1085 28362 1127 28396
rect 1161 28362 1203 28396
rect 1237 28362 1279 28396
rect 999 28327 1313 28362
rect 999 28293 1051 28327
rect 1085 28293 1127 28327
rect 1161 28293 1203 28327
rect 1237 28293 1279 28327
rect 999 28258 1313 28293
rect 999 28224 1051 28258
rect 1085 28224 1127 28258
rect 1161 28224 1203 28258
rect 1237 28224 1279 28258
rect 999 28189 1313 28224
rect 999 28155 1051 28189
rect 1085 28155 1127 28189
rect 1161 28155 1203 28189
rect 1237 28155 1279 28189
rect 999 28120 1313 28155
rect 999 28086 1051 28120
rect 1085 28086 1127 28120
rect 1161 28086 1203 28120
rect 1237 28086 1279 28120
rect 999 28051 1313 28086
rect 999 28017 1051 28051
rect 1085 28017 1127 28051
rect 1161 28017 1203 28051
rect 1237 28017 1279 28051
rect 999 27982 1313 28017
rect 999 27948 1051 27982
rect 1085 27948 1127 27982
rect 1161 27948 1203 27982
rect 1237 27948 1279 27982
rect 999 27913 1313 27948
rect 999 27879 1051 27913
rect 1085 27879 1127 27913
rect 1161 27879 1203 27913
rect 1237 27879 1279 27913
rect 999 27844 1313 27879
rect 999 27810 1051 27844
rect 1085 27810 1127 27844
rect 1161 27810 1203 27844
rect 1237 27810 1279 27844
rect 999 27775 1313 27810
rect 999 27741 1051 27775
rect 1085 27741 1127 27775
rect 1161 27741 1203 27775
rect 1237 27741 1279 27775
rect 999 27706 1313 27741
rect 999 27672 1051 27706
rect 1085 27672 1127 27706
rect 1161 27672 1203 27706
rect 1237 27672 1279 27706
rect 999 27637 1313 27672
rect 999 27603 1051 27637
rect 1085 27603 1127 27637
rect 1161 27603 1203 27637
rect 1237 27603 1279 27637
rect 999 27568 1313 27603
rect 999 27534 1051 27568
rect 1085 27534 1127 27568
rect 1161 27534 1203 27568
rect 1237 27534 1279 27568
rect 999 27499 1313 27534
rect 999 27465 1051 27499
rect 1085 27465 1127 27499
rect 1161 27465 1203 27499
rect 1237 27465 1279 27499
rect 999 27430 1313 27465
rect 999 27396 1051 27430
rect 1085 27396 1127 27430
rect 1161 27396 1203 27430
rect 1237 27396 1279 27430
rect 999 27361 1313 27396
rect 999 27327 1051 27361
rect 1085 27327 1127 27361
rect 1161 27327 1203 27361
rect 1237 27327 1279 27361
rect 999 27292 1313 27327
rect 999 27258 1051 27292
rect 1085 27258 1127 27292
rect 1161 27258 1203 27292
rect 1237 27258 1279 27292
rect 999 27223 1313 27258
rect 999 27189 1051 27223
rect 1085 27189 1127 27223
rect 1161 27189 1203 27223
rect 1237 27189 1279 27223
rect 999 27103 1313 27189
rect 18022 31675 18442 31709
rect 18022 31641 18025 31675
rect 18059 31641 18101 31675
rect 18135 31641 18177 31675
rect 18211 31641 18253 31675
rect 18287 31641 18329 31675
rect 18363 31641 18405 31675
rect 18439 31641 18442 31675
rect 18022 31607 18442 31641
rect 18022 31573 18025 31607
rect 18059 31573 18101 31607
rect 18135 31573 18177 31607
rect 18211 31573 18253 31607
rect 18287 31573 18329 31607
rect 18363 31573 18405 31607
rect 18439 31573 18442 31607
rect 18022 31539 18442 31573
rect 18022 31505 18025 31539
rect 18059 31505 18101 31539
rect 18135 31505 18177 31539
rect 18211 31505 18253 31539
rect 18287 31505 18329 31539
rect 18363 31505 18405 31539
rect 18439 31505 18442 31539
rect 18022 31471 18442 31505
rect 18022 31437 18025 31471
rect 18059 31437 18101 31471
rect 18135 31437 18177 31471
rect 18211 31437 18253 31471
rect 18287 31437 18329 31471
rect 18363 31437 18405 31471
rect 18439 31437 18442 31471
rect 18022 31403 18442 31437
rect 18022 31369 18025 31403
rect 18059 31369 18101 31403
rect 18135 31369 18177 31403
rect 18211 31369 18253 31403
rect 18287 31369 18329 31403
rect 18363 31369 18405 31403
rect 18439 31369 18442 31403
rect 18022 31335 18442 31369
rect 18022 31301 18025 31335
rect 18059 31301 18101 31335
rect 18135 31301 18177 31335
rect 18211 31301 18253 31335
rect 18287 31301 18329 31335
rect 18363 31301 18405 31335
rect 18439 31301 18442 31335
rect 18022 31267 18442 31301
rect 18022 31233 18025 31267
rect 18059 31233 18101 31267
rect 18135 31233 18177 31267
rect 18211 31233 18253 31267
rect 18287 31233 18329 31267
rect 18363 31233 18405 31267
rect 18439 31233 18442 31267
rect 18022 31199 18442 31233
rect 18022 31165 18025 31199
rect 18059 31165 18101 31199
rect 18135 31165 18177 31199
rect 18211 31165 18253 31199
rect 18287 31165 18329 31199
rect 18363 31165 18405 31199
rect 18439 31165 18442 31199
rect 18022 31131 18442 31165
rect 18022 31097 18025 31131
rect 18059 31097 18101 31131
rect 18135 31097 18177 31131
rect 18211 31097 18253 31131
rect 18287 31097 18329 31131
rect 18363 31097 18405 31131
rect 18439 31097 18442 31131
rect 18022 31063 18442 31097
rect 18022 31029 18025 31063
rect 18059 31029 18101 31063
rect 18135 31029 18177 31063
rect 18211 31029 18253 31063
rect 18287 31029 18329 31063
rect 18363 31029 18405 31063
rect 18439 31029 18442 31063
rect 18022 30995 18442 31029
rect 18022 30961 18025 30995
rect 18059 30961 18101 30995
rect 18135 30961 18177 30995
rect 18211 30961 18253 30995
rect 18287 30961 18329 30995
rect 18363 30961 18405 30995
rect 18439 30961 18442 30995
rect 18022 30927 18442 30961
rect 18022 30893 18025 30927
rect 18059 30893 18101 30927
rect 18135 30893 18177 30927
rect 18211 30893 18253 30927
rect 18287 30893 18329 30927
rect 18363 30893 18405 30927
rect 18439 30893 18442 30927
rect 18022 30859 18442 30893
rect 18022 30825 18025 30859
rect 18059 30825 18101 30859
rect 18135 30825 18177 30859
rect 18211 30825 18253 30859
rect 18287 30825 18329 30859
rect 18363 30825 18405 30859
rect 18439 30825 18442 30859
rect 18022 30791 18442 30825
rect 18022 30757 18025 30791
rect 18059 30757 18101 30791
rect 18135 30757 18177 30791
rect 18211 30757 18253 30791
rect 18287 30757 18329 30791
rect 18363 30757 18405 30791
rect 18439 30757 18442 30791
rect 18022 30723 18442 30757
rect 18022 30689 18025 30723
rect 18059 30689 18101 30723
rect 18135 30689 18177 30723
rect 18211 30689 18253 30723
rect 18287 30689 18329 30723
rect 18363 30689 18405 30723
rect 18439 30705 18442 30723
rect 22823 33301 23635 33335
rect 22823 33267 22827 33301
rect 22861 33267 22897 33301
rect 22931 33267 22967 33301
rect 23001 33267 23037 33301
rect 23071 33267 23107 33301
rect 23141 33267 23177 33301
rect 23211 33267 23247 33301
rect 23281 33267 23317 33301
rect 23351 33267 23387 33301
rect 23421 33267 23457 33301
rect 23491 33267 23527 33301
rect 23561 33267 23597 33301
rect 23631 33267 23635 33301
rect 22823 33233 23635 33267
rect 22823 33199 22827 33233
rect 22861 33199 22897 33233
rect 22931 33199 22967 33233
rect 23001 33199 23037 33233
rect 23071 33199 23107 33233
rect 23141 33199 23177 33233
rect 23211 33199 23247 33233
rect 23281 33199 23317 33233
rect 23351 33199 23387 33233
rect 23421 33199 23457 33233
rect 23491 33199 23527 33233
rect 23561 33199 23597 33233
rect 23631 33199 23635 33233
rect 22823 33165 23635 33199
rect 22823 33131 22827 33165
rect 22861 33131 22897 33165
rect 22931 33131 22967 33165
rect 23001 33131 23037 33165
rect 23071 33131 23107 33165
rect 23141 33131 23177 33165
rect 23211 33131 23247 33165
rect 23281 33131 23317 33165
rect 23351 33131 23387 33165
rect 23421 33131 23457 33165
rect 23491 33131 23527 33165
rect 23561 33131 23597 33165
rect 23631 33131 23635 33165
rect 22823 33097 23635 33131
rect 22823 33063 22827 33097
rect 22861 33063 22897 33097
rect 22931 33063 22967 33097
rect 23001 33063 23037 33097
rect 23071 33063 23107 33097
rect 23141 33063 23177 33097
rect 23211 33063 23247 33097
rect 23281 33063 23317 33097
rect 23351 33063 23387 33097
rect 23421 33063 23457 33097
rect 23491 33063 23527 33097
rect 23561 33063 23597 33097
rect 23631 33063 23635 33097
rect 22823 33029 23635 33063
rect 22823 32995 22827 33029
rect 22861 32995 22897 33029
rect 22931 32995 22967 33029
rect 23001 32995 23037 33029
rect 23071 32995 23107 33029
rect 23141 32995 23177 33029
rect 23211 32995 23247 33029
rect 23281 32995 23317 33029
rect 23351 32995 23387 33029
rect 23421 32995 23457 33029
rect 23491 32995 23527 33029
rect 23561 32995 23597 33029
rect 23631 32995 23635 33029
rect 22823 32961 23635 32995
rect 22823 32927 22827 32961
rect 22861 32927 22897 32961
rect 22931 32927 22967 32961
rect 23001 32927 23037 32961
rect 23071 32927 23107 32961
rect 23141 32927 23177 32961
rect 23211 32927 23247 32961
rect 23281 32927 23317 32961
rect 23351 32927 23387 32961
rect 23421 32927 23457 32961
rect 23491 32927 23527 32961
rect 23561 32927 23597 32961
rect 23631 32927 23635 32961
rect 22823 32893 23635 32927
rect 22823 32859 22827 32893
rect 22861 32859 22897 32893
rect 22931 32859 22967 32893
rect 23001 32859 23037 32893
rect 23071 32859 23107 32893
rect 23141 32859 23177 32893
rect 23211 32859 23247 32893
rect 23281 32859 23317 32893
rect 23351 32859 23387 32893
rect 23421 32859 23457 32893
rect 23491 32859 23527 32893
rect 23561 32859 23597 32893
rect 23631 32859 23635 32893
rect 22823 32825 23635 32859
rect 22823 32791 22827 32825
rect 22861 32791 22897 32825
rect 22931 32791 22967 32825
rect 23001 32791 23037 32825
rect 23071 32791 23107 32825
rect 23141 32791 23177 32825
rect 23211 32791 23247 32825
rect 23281 32791 23317 32825
rect 23351 32791 23387 32825
rect 23421 32791 23457 32825
rect 23491 32791 23527 32825
rect 23561 32791 23597 32825
rect 23631 32791 23635 32825
rect 22823 32757 23635 32791
rect 22823 32723 22827 32757
rect 22861 32723 22897 32757
rect 22931 32723 22967 32757
rect 23001 32723 23037 32757
rect 23071 32723 23107 32757
rect 23141 32723 23177 32757
rect 23211 32723 23247 32757
rect 23281 32723 23317 32757
rect 23351 32723 23387 32757
rect 23421 32723 23457 32757
rect 23491 32723 23527 32757
rect 23561 32723 23597 32757
rect 23631 32723 23635 32757
rect 22823 32689 23635 32723
rect 22823 32655 22827 32689
rect 22861 32655 22897 32689
rect 22931 32655 22967 32689
rect 23001 32655 23037 32689
rect 23071 32655 23107 32689
rect 23141 32655 23177 32689
rect 23211 32655 23247 32689
rect 23281 32655 23317 32689
rect 23351 32655 23387 32689
rect 23421 32655 23457 32689
rect 23491 32655 23527 32689
rect 23561 32655 23597 32689
rect 23631 32655 23635 32689
rect 22823 32621 23635 32655
rect 22823 32587 22827 32621
rect 22861 32587 22897 32621
rect 22931 32587 22967 32621
rect 23001 32587 23037 32621
rect 23071 32587 23107 32621
rect 23141 32587 23177 32621
rect 23211 32587 23247 32621
rect 23281 32587 23317 32621
rect 23351 32587 23387 32621
rect 23421 32587 23457 32621
rect 23491 32587 23527 32621
rect 23561 32587 23597 32621
rect 23631 32587 23635 32621
rect 22823 32553 23635 32587
rect 22823 32519 22827 32553
rect 22861 32519 22897 32553
rect 22931 32519 22967 32553
rect 23001 32519 23037 32553
rect 23071 32519 23107 32553
rect 23141 32519 23177 32553
rect 23211 32519 23247 32553
rect 23281 32519 23317 32553
rect 23351 32519 23387 32553
rect 23421 32519 23457 32553
rect 23491 32519 23527 32553
rect 23561 32519 23597 32553
rect 23631 32519 23635 32553
rect 22823 32485 23635 32519
rect 22823 32451 22827 32485
rect 22861 32451 22897 32485
rect 22931 32451 22967 32485
rect 23001 32451 23037 32485
rect 23071 32451 23107 32485
rect 23141 32451 23177 32485
rect 23211 32451 23247 32485
rect 23281 32451 23317 32485
rect 23351 32451 23387 32485
rect 23421 32451 23457 32485
rect 23491 32451 23527 32485
rect 23561 32451 23597 32485
rect 23631 32451 23635 32485
rect 22823 32417 23635 32451
rect 22823 32383 22827 32417
rect 22861 32383 22897 32417
rect 22931 32383 22967 32417
rect 23001 32383 23037 32417
rect 23071 32383 23107 32417
rect 23141 32383 23177 32417
rect 23211 32383 23247 32417
rect 23281 32383 23317 32417
rect 23351 32383 23387 32417
rect 23421 32383 23457 32417
rect 23491 32383 23527 32417
rect 23561 32383 23597 32417
rect 23631 32383 23635 32417
rect 22823 32349 23635 32383
rect 22823 32315 22827 32349
rect 22861 32315 22897 32349
rect 22931 32315 22967 32349
rect 23001 32315 23037 32349
rect 23071 32315 23107 32349
rect 23141 32315 23177 32349
rect 23211 32315 23247 32349
rect 23281 32315 23317 32349
rect 23351 32315 23387 32349
rect 23421 32315 23457 32349
rect 23491 32315 23527 32349
rect 23561 32315 23597 32349
rect 23631 32315 23635 32349
rect 22823 32281 23635 32315
rect 22823 32247 22827 32281
rect 22861 32247 22897 32281
rect 22931 32247 22967 32281
rect 23001 32247 23037 32281
rect 23071 32247 23107 32281
rect 23141 32247 23177 32281
rect 23211 32247 23247 32281
rect 23281 32247 23317 32281
rect 23351 32247 23387 32281
rect 23421 32247 23457 32281
rect 23491 32247 23527 32281
rect 23561 32247 23597 32281
rect 23631 32247 23635 32281
rect 22823 32213 23635 32247
rect 22823 32179 22827 32213
rect 22861 32179 22897 32213
rect 22931 32179 22967 32213
rect 23001 32179 23037 32213
rect 23071 32179 23107 32213
rect 23141 32179 23177 32213
rect 23211 32179 23247 32213
rect 23281 32179 23317 32213
rect 23351 32179 23387 32213
rect 23421 32179 23457 32213
rect 23491 32179 23527 32213
rect 23561 32179 23597 32213
rect 23631 32179 23635 32213
rect 22823 32145 23635 32179
rect 22823 32111 22827 32145
rect 22861 32111 22897 32145
rect 22931 32111 22967 32145
rect 23001 32111 23037 32145
rect 23071 32111 23107 32145
rect 23141 32111 23177 32145
rect 23211 32111 23247 32145
rect 23281 32111 23317 32145
rect 23351 32111 23387 32145
rect 23421 32111 23457 32145
rect 23491 32111 23527 32145
rect 23561 32111 23597 32145
rect 23631 32111 23635 32145
rect 22823 32077 23635 32111
rect 22823 32043 22827 32077
rect 22861 32043 22897 32077
rect 22931 32043 22967 32077
rect 23001 32043 23037 32077
rect 23071 32043 23107 32077
rect 23141 32043 23177 32077
rect 23211 32043 23247 32077
rect 23281 32043 23317 32077
rect 23351 32043 23387 32077
rect 23421 32043 23457 32077
rect 23491 32043 23527 32077
rect 23561 32043 23597 32077
rect 23631 32043 23635 32077
rect 22823 32009 23635 32043
rect 22823 31975 22827 32009
rect 22861 31975 22897 32009
rect 22931 31975 22967 32009
rect 23001 31975 23037 32009
rect 23071 31975 23107 32009
rect 23141 31975 23177 32009
rect 23211 31975 23247 32009
rect 23281 31975 23317 32009
rect 23351 31975 23387 32009
rect 23421 31975 23457 32009
rect 23491 31975 23527 32009
rect 23561 31975 23597 32009
rect 23631 31975 23635 32009
rect 22823 31941 23635 31975
rect 22823 31907 22827 31941
rect 22861 31907 22897 31941
rect 22931 31907 22967 31941
rect 23001 31907 23037 31941
rect 23071 31907 23107 31941
rect 23141 31907 23177 31941
rect 23211 31907 23247 31941
rect 23281 31907 23317 31941
rect 23351 31907 23387 31941
rect 23421 31907 23457 31941
rect 23491 31907 23527 31941
rect 23561 31907 23597 31941
rect 23631 31907 23635 31941
rect 22823 31873 23635 31907
rect 22823 31839 22827 31873
rect 22861 31839 22897 31873
rect 22931 31839 22967 31873
rect 23001 31839 23037 31873
rect 23071 31839 23107 31873
rect 23141 31839 23177 31873
rect 23211 31839 23247 31873
rect 23281 31839 23317 31873
rect 23351 31839 23387 31873
rect 23421 31839 23457 31873
rect 23491 31839 23527 31873
rect 23561 31839 23597 31873
rect 23631 31839 23635 31873
rect 22823 31805 23635 31839
rect 22823 31771 22827 31805
rect 22861 31771 22897 31805
rect 22931 31771 22967 31805
rect 23001 31771 23037 31805
rect 23071 31771 23107 31805
rect 23141 31771 23177 31805
rect 23211 31771 23247 31805
rect 23281 31771 23317 31805
rect 23351 31771 23387 31805
rect 23421 31771 23457 31805
rect 23491 31771 23527 31805
rect 23561 31771 23597 31805
rect 23631 31771 23635 31805
rect 22823 31737 23635 31771
rect 22823 31703 22827 31737
rect 22861 31703 22897 31737
rect 22931 31703 22967 31737
rect 23001 31703 23037 31737
rect 23071 31703 23107 31737
rect 23141 31703 23177 31737
rect 23211 31703 23247 31737
rect 23281 31703 23317 31737
rect 23351 31703 23387 31737
rect 23421 31703 23457 31737
rect 23491 31703 23527 31737
rect 23561 31703 23597 31737
rect 23631 31703 23635 31737
rect 22823 31669 23635 31703
rect 22823 31635 22827 31669
rect 22861 31635 22897 31669
rect 22931 31635 22967 31669
rect 23001 31635 23037 31669
rect 23071 31635 23107 31669
rect 23141 31635 23177 31669
rect 23211 31635 23247 31669
rect 23281 31635 23317 31669
rect 23351 31635 23387 31669
rect 23421 31635 23457 31669
rect 23491 31635 23527 31669
rect 23561 31635 23597 31669
rect 23631 31635 23635 31669
rect 22823 31601 23635 31635
rect 22823 31567 22827 31601
rect 22861 31567 22897 31601
rect 22931 31567 22967 31601
rect 23001 31567 23037 31601
rect 23071 31567 23107 31601
rect 23141 31567 23177 31601
rect 23211 31567 23247 31601
rect 23281 31567 23317 31601
rect 23351 31567 23387 31601
rect 23421 31567 23457 31601
rect 23491 31567 23527 31601
rect 23561 31567 23597 31601
rect 23631 31567 23635 31601
rect 22823 31533 23635 31567
rect 22823 31499 22827 31533
rect 22861 31499 22897 31533
rect 22931 31499 22967 31533
rect 23001 31499 23037 31533
rect 23071 31499 23107 31533
rect 23141 31499 23177 31533
rect 23211 31499 23247 31533
rect 23281 31499 23317 31533
rect 23351 31499 23387 31533
rect 23421 31499 23457 31533
rect 23491 31499 23527 31533
rect 23561 31499 23597 31533
rect 23631 31499 23635 31533
rect 22823 31465 23635 31499
rect 22823 31431 22827 31465
rect 22861 31431 22897 31465
rect 22931 31431 22967 31465
rect 23001 31431 23037 31465
rect 23071 31431 23107 31465
rect 23141 31431 23177 31465
rect 23211 31431 23247 31465
rect 23281 31431 23317 31465
rect 23351 31431 23387 31465
rect 23421 31431 23457 31465
rect 23491 31431 23527 31465
rect 23561 31431 23597 31465
rect 23631 31431 23635 31465
rect 22823 31397 23635 31431
rect 22823 31363 22827 31397
rect 22861 31363 22897 31397
rect 22931 31363 22967 31397
rect 23001 31363 23037 31397
rect 23071 31363 23107 31397
rect 23141 31363 23177 31397
rect 23211 31363 23247 31397
rect 23281 31363 23317 31397
rect 23351 31363 23387 31397
rect 23421 31363 23457 31397
rect 23491 31363 23527 31397
rect 23561 31363 23597 31397
rect 23631 31363 23635 31397
rect 22823 31329 23635 31363
rect 22823 31295 22827 31329
rect 22861 31295 22897 31329
rect 22931 31295 22967 31329
rect 23001 31295 23037 31329
rect 23071 31295 23107 31329
rect 23141 31295 23177 31329
rect 23211 31295 23247 31329
rect 23281 31295 23317 31329
rect 23351 31295 23387 31329
rect 23421 31295 23457 31329
rect 23491 31295 23527 31329
rect 23561 31295 23597 31329
rect 23631 31295 23635 31329
rect 22823 31261 23635 31295
rect 22823 31227 22827 31261
rect 22861 31227 22897 31261
rect 22931 31227 22967 31261
rect 23001 31227 23037 31261
rect 23071 31227 23107 31261
rect 23141 31227 23177 31261
rect 23211 31227 23247 31261
rect 23281 31227 23317 31261
rect 23351 31227 23387 31261
rect 23421 31227 23457 31261
rect 23491 31227 23527 31261
rect 23561 31227 23597 31261
rect 23631 31227 23635 31261
rect 22823 31193 23635 31227
rect 22823 31159 22827 31193
rect 22861 31159 22897 31193
rect 22931 31159 22967 31193
rect 23001 31159 23037 31193
rect 23071 31159 23107 31193
rect 23141 31159 23177 31193
rect 23211 31159 23247 31193
rect 23281 31159 23317 31193
rect 23351 31159 23387 31193
rect 23421 31159 23457 31193
rect 23491 31159 23527 31193
rect 23561 31159 23597 31193
rect 23631 31159 23635 31193
rect 22823 31125 23635 31159
rect 22823 31091 22827 31125
rect 22861 31091 22897 31125
rect 22931 31091 22967 31125
rect 23001 31091 23037 31125
rect 23071 31091 23107 31125
rect 23141 31091 23177 31125
rect 23211 31091 23247 31125
rect 23281 31091 23317 31125
rect 23351 31091 23387 31125
rect 23421 31091 23457 31125
rect 23491 31091 23527 31125
rect 23561 31091 23597 31125
rect 23631 31091 23635 31125
rect 22823 31057 23635 31091
rect 22823 31023 22827 31057
rect 22861 31023 22897 31057
rect 22931 31023 22967 31057
rect 23001 31023 23037 31057
rect 23071 31023 23107 31057
rect 23141 31023 23177 31057
rect 23211 31023 23247 31057
rect 23281 31023 23317 31057
rect 23351 31023 23387 31057
rect 23421 31023 23457 31057
rect 23491 31023 23527 31057
rect 23561 31023 23597 31057
rect 23631 31023 23635 31057
rect 22823 30989 23635 31023
rect 22823 30955 22827 30989
rect 22861 30955 22897 30989
rect 22931 30955 22967 30989
rect 23001 30955 23037 30989
rect 23071 30955 23107 30989
rect 23141 30955 23177 30989
rect 23211 30955 23247 30989
rect 23281 30955 23317 30989
rect 23351 30955 23387 30989
rect 23421 30955 23457 30989
rect 23491 30955 23527 30989
rect 23561 30955 23597 30989
rect 23631 30955 23635 30989
rect 22823 30921 23635 30955
rect 22823 30887 22827 30921
rect 22861 30887 22897 30921
rect 22931 30887 22967 30921
rect 23001 30887 23037 30921
rect 23071 30887 23107 30921
rect 23141 30887 23177 30921
rect 23211 30887 23247 30921
rect 23281 30887 23317 30921
rect 23351 30887 23387 30921
rect 23421 30887 23457 30921
rect 23491 30887 23527 30921
rect 23561 30887 23597 30921
rect 23631 30887 23635 30921
rect 22823 30853 23635 30887
rect 22823 30819 22827 30853
rect 22861 30819 22897 30853
rect 22931 30819 22967 30853
rect 23001 30819 23037 30853
rect 23071 30819 23107 30853
rect 23141 30819 23177 30853
rect 23211 30819 23247 30853
rect 23281 30819 23317 30853
rect 23351 30819 23387 30853
rect 23421 30819 23457 30853
rect 23491 30819 23527 30853
rect 23561 30819 23597 30853
rect 23631 30819 23635 30853
rect 22823 30785 23635 30819
rect 22823 30751 22827 30785
rect 22861 30751 22897 30785
rect 22931 30751 22967 30785
rect 23001 30751 23037 30785
rect 23071 30751 23107 30785
rect 23141 30751 23177 30785
rect 23211 30751 23247 30785
rect 23281 30751 23317 30785
rect 23351 30751 23387 30785
rect 23421 30751 23457 30785
rect 23491 30751 23527 30785
rect 23561 30751 23597 30785
rect 23631 30751 23635 30785
rect 22823 30717 23635 30751
rect 18439 30689 19012 30705
rect 18022 30671 19012 30689
rect 18022 30655 18486 30671
rect 18022 30621 18025 30655
rect 18059 30621 18101 30655
rect 18135 30621 18177 30655
rect 18211 30621 18253 30655
rect 18287 30621 18329 30655
rect 18363 30621 18405 30655
rect 18439 30637 18486 30655
rect 18520 30637 18556 30671
rect 18590 30637 18626 30671
rect 18660 30637 18696 30671
rect 18730 30637 18766 30671
rect 18800 30637 18836 30671
rect 18870 30637 18906 30671
rect 18940 30637 18976 30671
rect 19010 30637 19012 30671
rect 18439 30621 19012 30637
rect 18022 30603 19012 30621
rect 18022 30587 18486 30603
rect 18022 30553 18025 30587
rect 18059 30553 18101 30587
rect 18135 30553 18177 30587
rect 18211 30553 18253 30587
rect 18287 30553 18329 30587
rect 18363 30553 18405 30587
rect 18439 30569 18486 30587
rect 18520 30569 18556 30603
rect 18590 30569 18626 30603
rect 18660 30569 18696 30603
rect 18730 30569 18766 30603
rect 18800 30569 18836 30603
rect 18870 30569 18906 30603
rect 18940 30569 18976 30603
rect 19010 30569 19012 30603
rect 18439 30553 19012 30569
rect 18022 30535 19012 30553
rect 18022 30519 18486 30535
rect 18022 30485 18025 30519
rect 18059 30485 18101 30519
rect 18135 30485 18177 30519
rect 18211 30485 18253 30519
rect 18287 30485 18329 30519
rect 18363 30485 18405 30519
rect 18439 30501 18486 30519
rect 18520 30501 18556 30535
rect 18590 30501 18626 30535
rect 18660 30501 18696 30535
rect 18730 30501 18766 30535
rect 18800 30501 18836 30535
rect 18870 30501 18906 30535
rect 18940 30501 18976 30535
rect 19010 30501 19012 30535
rect 18439 30485 19012 30501
rect 18022 30467 19012 30485
rect 18022 30451 18486 30467
rect 18022 30417 18025 30451
rect 18059 30417 18101 30451
rect 18135 30417 18177 30451
rect 18211 30417 18253 30451
rect 18287 30417 18329 30451
rect 18363 30417 18405 30451
rect 18439 30433 18486 30451
rect 18520 30433 18556 30467
rect 18590 30433 18626 30467
rect 18660 30433 18696 30467
rect 18730 30433 18766 30467
rect 18800 30433 18836 30467
rect 18870 30433 18906 30467
rect 18940 30433 18976 30467
rect 19010 30433 19012 30467
rect 18439 30417 19012 30433
rect 18022 30399 19012 30417
rect 18022 30383 18486 30399
rect 18022 30349 18025 30383
rect 18059 30349 18101 30383
rect 18135 30349 18177 30383
rect 18211 30349 18253 30383
rect 18287 30349 18329 30383
rect 18363 30349 18405 30383
rect 18439 30365 18486 30383
rect 18520 30365 18556 30399
rect 18590 30365 18626 30399
rect 18660 30365 18696 30399
rect 18730 30365 18766 30399
rect 18800 30365 18836 30399
rect 18870 30365 18906 30399
rect 18940 30365 18976 30399
rect 19010 30365 19012 30399
rect 18439 30349 19012 30365
rect 18022 30331 19012 30349
rect 18022 30315 18486 30331
rect 18022 30281 18025 30315
rect 18059 30281 18101 30315
rect 18135 30281 18177 30315
rect 18211 30281 18253 30315
rect 18287 30281 18329 30315
rect 18363 30281 18405 30315
rect 18439 30297 18486 30315
rect 18520 30297 18556 30331
rect 18590 30297 18626 30331
rect 18660 30297 18696 30331
rect 18730 30297 18766 30331
rect 18800 30297 18836 30331
rect 18870 30297 18906 30331
rect 18940 30297 18976 30331
rect 19010 30297 19012 30331
rect 18439 30281 19012 30297
rect 18022 30263 19012 30281
rect 18022 30247 18486 30263
rect 18022 30213 18025 30247
rect 18059 30213 18101 30247
rect 18135 30213 18177 30247
rect 18211 30213 18253 30247
rect 18287 30213 18329 30247
rect 18363 30213 18405 30247
rect 18439 30229 18486 30247
rect 18520 30229 18556 30263
rect 18590 30229 18626 30263
rect 18660 30229 18696 30263
rect 18730 30229 18766 30263
rect 18800 30229 18836 30263
rect 18870 30229 18906 30263
rect 18940 30229 18976 30263
rect 19010 30229 19012 30263
rect 18439 30213 19012 30229
rect 18022 30195 19012 30213
rect 18022 30179 18486 30195
rect 18022 30145 18025 30179
rect 18059 30145 18101 30179
rect 18135 30145 18177 30179
rect 18211 30145 18253 30179
rect 18287 30145 18329 30179
rect 18363 30145 18405 30179
rect 18439 30161 18486 30179
rect 18520 30161 18556 30195
rect 18590 30161 18626 30195
rect 18660 30161 18696 30195
rect 18730 30161 18766 30195
rect 18800 30161 18836 30195
rect 18870 30161 18906 30195
rect 18940 30161 18976 30195
rect 19010 30161 19012 30195
rect 18439 30145 19012 30161
rect 18022 30127 19012 30145
rect 18022 30111 18486 30127
rect 18022 30077 18025 30111
rect 18059 30077 18101 30111
rect 18135 30077 18177 30111
rect 18211 30077 18253 30111
rect 18287 30077 18329 30111
rect 18363 30077 18405 30111
rect 18439 30093 18486 30111
rect 18520 30093 18556 30127
rect 18590 30093 18626 30127
rect 18660 30093 18696 30127
rect 18730 30093 18766 30127
rect 18800 30093 18836 30127
rect 18870 30093 18906 30127
rect 18940 30093 18976 30127
rect 19010 30093 19012 30127
rect 18439 30077 19012 30093
rect 18022 30059 19012 30077
rect 18022 30043 18486 30059
rect 18022 30009 18025 30043
rect 18059 30009 18101 30043
rect 18135 30009 18177 30043
rect 18211 30009 18253 30043
rect 18287 30009 18329 30043
rect 18363 30009 18405 30043
rect 18439 30025 18486 30043
rect 18520 30025 18556 30059
rect 18590 30025 18626 30059
rect 18660 30025 18696 30059
rect 18730 30025 18766 30059
rect 18800 30025 18836 30059
rect 18870 30025 18906 30059
rect 18940 30025 18976 30059
rect 19010 30025 19012 30059
rect 18439 30009 19012 30025
rect 18022 29991 19012 30009
rect 18022 29975 18486 29991
rect 18022 29941 18025 29975
rect 18059 29941 18101 29975
rect 18135 29941 18177 29975
rect 18211 29941 18253 29975
rect 18287 29941 18329 29975
rect 18363 29941 18405 29975
rect 18439 29957 18486 29975
rect 18520 29957 18556 29991
rect 18590 29957 18626 29991
rect 18660 29957 18696 29991
rect 18730 29957 18766 29991
rect 18800 29957 18836 29991
rect 18870 29957 18906 29991
rect 18940 29957 18976 29991
rect 19010 29957 19012 29991
rect 18439 29941 19012 29957
rect 18022 29923 19012 29941
rect 18022 29907 18486 29923
rect 18022 29873 18025 29907
rect 18059 29873 18101 29907
rect 18135 29873 18177 29907
rect 18211 29873 18253 29907
rect 18287 29873 18329 29907
rect 18363 29873 18405 29907
rect 18439 29889 18486 29907
rect 18520 29889 18556 29923
rect 18590 29889 18626 29923
rect 18660 29889 18696 29923
rect 18730 29889 18766 29923
rect 18800 29889 18836 29923
rect 18870 29889 18906 29923
rect 18940 29889 18976 29923
rect 19010 29889 19012 29923
rect 18439 29873 19012 29889
rect 18022 29855 19012 29873
rect 18022 29839 18486 29855
rect 18022 29805 18025 29839
rect 18059 29805 18101 29839
rect 18135 29805 18177 29839
rect 18211 29805 18253 29839
rect 18287 29805 18329 29839
rect 18363 29805 18405 29839
rect 18439 29821 18486 29839
rect 18520 29821 18556 29855
rect 18590 29821 18626 29855
rect 18660 29821 18696 29855
rect 18730 29821 18766 29855
rect 18800 29821 18836 29855
rect 18870 29821 18906 29855
rect 18940 29821 18976 29855
rect 19010 29821 19012 29855
rect 18439 29805 19012 29821
rect 18022 29787 19012 29805
rect 18022 29771 18486 29787
rect 18022 29737 18025 29771
rect 18059 29737 18101 29771
rect 18135 29737 18177 29771
rect 18211 29737 18253 29771
rect 18287 29737 18329 29771
rect 18363 29737 18405 29771
rect 18439 29753 18486 29771
rect 18520 29753 18556 29787
rect 18590 29753 18626 29787
rect 18660 29753 18696 29787
rect 18730 29753 18766 29787
rect 18800 29753 18836 29787
rect 18870 29753 18906 29787
rect 18940 29753 18976 29787
rect 19010 29753 19012 29787
rect 18439 29737 19012 29753
rect 18022 29719 19012 29737
rect 18022 29703 18486 29719
rect 18022 29669 18025 29703
rect 18059 29669 18101 29703
rect 18135 29669 18177 29703
rect 18211 29669 18253 29703
rect 18287 29669 18329 29703
rect 18363 29669 18405 29703
rect 18439 29685 18486 29703
rect 18520 29685 18556 29719
rect 18590 29685 18626 29719
rect 18660 29685 18696 29719
rect 18730 29685 18766 29719
rect 18800 29685 18836 29719
rect 18870 29685 18906 29719
rect 18940 29685 18976 29719
rect 19010 29685 19012 29719
rect 18439 29669 19012 29685
rect 18022 29651 19012 29669
rect 18022 29635 18486 29651
rect 18022 29601 18025 29635
rect 18059 29601 18101 29635
rect 18135 29601 18177 29635
rect 18211 29601 18253 29635
rect 18287 29601 18329 29635
rect 18363 29601 18405 29635
rect 18439 29617 18486 29635
rect 18520 29617 18556 29651
rect 18590 29617 18626 29651
rect 18660 29617 18696 29651
rect 18730 29617 18766 29651
rect 18800 29617 18836 29651
rect 18870 29617 18906 29651
rect 18940 29617 18976 29651
rect 19010 29617 19012 29651
rect 18439 29601 19012 29617
rect 18022 29583 19012 29601
rect 18022 29567 18486 29583
rect 18022 29533 18025 29567
rect 18059 29533 18101 29567
rect 18135 29533 18177 29567
rect 18211 29533 18253 29567
rect 18287 29533 18329 29567
rect 18363 29533 18405 29567
rect 18439 29549 18486 29567
rect 18520 29549 18556 29583
rect 18590 29549 18626 29583
rect 18660 29549 18696 29583
rect 18730 29549 18766 29583
rect 18800 29549 18836 29583
rect 18870 29549 18906 29583
rect 18940 29549 18976 29583
rect 19010 29549 19012 29583
rect 18439 29533 19012 29549
rect 18022 29515 19012 29533
rect 18022 29499 18486 29515
rect 18022 29465 18025 29499
rect 18059 29465 18101 29499
rect 18135 29465 18177 29499
rect 18211 29465 18253 29499
rect 18287 29465 18329 29499
rect 18363 29465 18405 29499
rect 18439 29481 18486 29499
rect 18520 29481 18556 29515
rect 18590 29481 18626 29515
rect 18660 29481 18696 29515
rect 18730 29481 18766 29515
rect 18800 29481 18836 29515
rect 18870 29481 18906 29515
rect 18940 29481 18976 29515
rect 19010 29481 19012 29515
rect 18439 29465 19012 29481
rect 18022 29447 19012 29465
rect 18022 29431 18486 29447
rect 18022 29397 18025 29431
rect 18059 29397 18101 29431
rect 18135 29397 18177 29431
rect 18211 29397 18253 29431
rect 18287 29397 18329 29431
rect 18363 29397 18405 29431
rect 18439 29413 18486 29431
rect 18520 29413 18556 29447
rect 18590 29413 18626 29447
rect 18660 29413 18696 29447
rect 18730 29413 18766 29447
rect 18800 29413 18836 29447
rect 18870 29413 18906 29447
rect 18940 29413 18976 29447
rect 19010 29413 19012 29447
rect 18439 29397 19012 29413
rect 18022 29379 19012 29397
rect 18022 29363 18486 29379
rect 18022 29329 18025 29363
rect 18059 29329 18101 29363
rect 18135 29329 18177 29363
rect 18211 29329 18253 29363
rect 18287 29329 18329 29363
rect 18363 29329 18405 29363
rect 18439 29345 18486 29363
rect 18520 29345 18556 29379
rect 18590 29345 18626 29379
rect 18660 29345 18696 29379
rect 18730 29345 18766 29379
rect 18800 29345 18836 29379
rect 18870 29345 18906 29379
rect 18940 29345 18976 29379
rect 19010 29345 19012 29379
rect 18439 29329 19012 29345
rect 18022 29311 19012 29329
rect 18022 29295 18486 29311
rect 18022 29261 18025 29295
rect 18059 29261 18101 29295
rect 18135 29261 18177 29295
rect 18211 29261 18253 29295
rect 18287 29261 18329 29295
rect 18363 29261 18405 29295
rect 18439 29277 18486 29295
rect 18520 29277 18556 29311
rect 18590 29277 18626 29311
rect 18660 29277 18696 29311
rect 18730 29277 18766 29311
rect 18800 29277 18836 29311
rect 18870 29277 18906 29311
rect 18940 29277 18976 29311
rect 19010 29277 19012 29311
rect 18439 29261 19012 29277
rect 18022 29243 19012 29261
rect 18022 29227 18486 29243
rect 18022 29193 18025 29227
rect 18059 29193 18101 29227
rect 18135 29193 18177 29227
rect 18211 29193 18253 29227
rect 18287 29193 18329 29227
rect 18363 29193 18405 29227
rect 18439 29209 18486 29227
rect 18520 29209 18556 29243
rect 18590 29209 18626 29243
rect 18660 29209 18696 29243
rect 18730 29209 18766 29243
rect 18800 29209 18836 29243
rect 18870 29209 18906 29243
rect 18940 29209 18976 29243
rect 19010 29209 19012 29243
rect 18439 29193 19012 29209
rect 18022 29175 19012 29193
rect 18022 29159 18486 29175
rect 18022 29125 18025 29159
rect 18059 29125 18101 29159
rect 18135 29125 18177 29159
rect 18211 29125 18253 29159
rect 18287 29125 18329 29159
rect 18363 29125 18405 29159
rect 18439 29141 18486 29159
rect 18520 29141 18556 29175
rect 18590 29141 18626 29175
rect 18660 29141 18696 29175
rect 18730 29141 18766 29175
rect 18800 29141 18836 29175
rect 18870 29141 18906 29175
rect 18940 29141 18976 29175
rect 19010 29141 19012 29175
rect 18439 29125 19012 29141
rect 18022 29107 19012 29125
rect 18022 29091 18486 29107
rect 18022 29057 18025 29091
rect 18059 29057 18101 29091
rect 18135 29057 18177 29091
rect 18211 29057 18253 29091
rect 18287 29057 18329 29091
rect 18363 29057 18405 29091
rect 18439 29073 18486 29091
rect 18520 29073 18556 29107
rect 18590 29073 18626 29107
rect 18660 29073 18696 29107
rect 18730 29073 18766 29107
rect 18800 29073 18836 29107
rect 18870 29073 18906 29107
rect 18940 29073 18976 29107
rect 19010 29073 19012 29107
rect 18439 29057 19012 29073
rect 18022 29039 19012 29057
rect 18022 29023 18486 29039
rect 18022 28989 18025 29023
rect 18059 28989 18101 29023
rect 18135 28989 18177 29023
rect 18211 28989 18253 29023
rect 18287 28989 18329 29023
rect 18363 28989 18405 29023
rect 18439 29005 18486 29023
rect 18520 29005 18556 29039
rect 18590 29005 18626 29039
rect 18660 29005 18696 29039
rect 18730 29005 18766 29039
rect 18800 29005 18836 29039
rect 18870 29005 18906 29039
rect 18940 29005 18976 29039
rect 19010 29005 19012 29039
rect 18439 28989 19012 29005
rect 18022 28971 19012 28989
rect 18022 28955 18486 28971
rect 18022 28921 18025 28955
rect 18059 28921 18101 28955
rect 18135 28921 18177 28955
rect 18211 28921 18253 28955
rect 18287 28921 18329 28955
rect 18363 28921 18405 28955
rect 18439 28937 18486 28955
rect 18520 28937 18556 28971
rect 18590 28937 18626 28971
rect 18660 28937 18696 28971
rect 18730 28937 18766 28971
rect 18800 28937 18836 28971
rect 18870 28937 18906 28971
rect 18940 28937 18976 28971
rect 19010 28937 19012 28971
rect 18439 28921 19012 28937
rect 18022 28903 19012 28921
rect 18022 28887 18486 28903
rect 18022 28853 18025 28887
rect 18059 28853 18101 28887
rect 18135 28853 18177 28887
rect 18211 28853 18253 28887
rect 18287 28853 18329 28887
rect 18363 28853 18405 28887
rect 18439 28869 18486 28887
rect 18520 28869 18556 28903
rect 18590 28869 18626 28903
rect 18660 28869 18696 28903
rect 18730 28869 18766 28903
rect 18800 28869 18836 28903
rect 18870 28869 18906 28903
rect 18940 28869 18976 28903
rect 19010 28869 19012 28903
rect 18439 28853 19012 28869
rect 18022 28835 19012 28853
rect 18022 28819 18486 28835
rect 18022 28785 18025 28819
rect 18059 28785 18101 28819
rect 18135 28785 18177 28819
rect 18211 28785 18253 28819
rect 18287 28785 18329 28819
rect 18363 28785 18405 28819
rect 18439 28801 18486 28819
rect 18520 28801 18556 28835
rect 18590 28801 18626 28835
rect 18660 28801 18696 28835
rect 18730 28801 18766 28835
rect 18800 28801 18836 28835
rect 18870 28801 18906 28835
rect 18940 28801 18976 28835
rect 19010 28801 19012 28835
rect 18439 28785 19012 28801
rect 18022 28767 19012 28785
rect 18022 28751 18486 28767
rect 18022 28717 18025 28751
rect 18059 28717 18101 28751
rect 18135 28717 18177 28751
rect 18211 28717 18253 28751
rect 18287 28717 18329 28751
rect 18363 28717 18405 28751
rect 18439 28733 18486 28751
rect 18520 28733 18556 28767
rect 18590 28733 18626 28767
rect 18660 28733 18696 28767
rect 18730 28733 18766 28767
rect 18800 28733 18836 28767
rect 18870 28733 18906 28767
rect 18940 28733 18976 28767
rect 19010 28733 19012 28767
rect 18439 28717 19012 28733
rect 18022 28699 19012 28717
rect 18022 28683 18486 28699
rect 18022 28649 18025 28683
rect 18059 28649 18101 28683
rect 18135 28649 18177 28683
rect 18211 28649 18253 28683
rect 18287 28649 18329 28683
rect 18363 28649 18405 28683
rect 18439 28665 18486 28683
rect 18520 28665 18556 28699
rect 18590 28665 18626 28699
rect 18660 28665 18696 28699
rect 18730 28665 18766 28699
rect 18800 28665 18836 28699
rect 18870 28665 18906 28699
rect 18940 28665 18976 28699
rect 19010 28665 19012 28699
rect 18439 28649 19012 28665
rect 18022 28631 19012 28649
rect 18022 28615 18486 28631
rect 18022 28581 18025 28615
rect 18059 28581 18101 28615
rect 18135 28581 18177 28615
rect 18211 28581 18253 28615
rect 18287 28581 18329 28615
rect 18363 28581 18405 28615
rect 18439 28597 18486 28615
rect 18520 28597 18556 28631
rect 18590 28597 18626 28631
rect 18660 28597 18696 28631
rect 18730 28597 18766 28631
rect 18800 28597 18836 28631
rect 18870 28597 18906 28631
rect 18940 28597 18976 28631
rect 19010 28597 19012 28631
rect 18439 28581 19012 28597
rect 18022 28563 19012 28581
rect 18022 28547 18486 28563
rect 18022 28513 18025 28547
rect 18059 28513 18101 28547
rect 18135 28513 18177 28547
rect 18211 28513 18253 28547
rect 18287 28513 18329 28547
rect 18363 28513 18405 28547
rect 18439 28529 18486 28547
rect 18520 28529 18556 28563
rect 18590 28529 18626 28563
rect 18660 28529 18696 28563
rect 18730 28529 18766 28563
rect 18800 28529 18836 28563
rect 18870 28529 18906 28563
rect 18940 28529 18976 28563
rect 19010 28529 19012 28563
rect 18439 28513 19012 28529
rect 18022 28495 19012 28513
rect 18022 28479 18486 28495
rect 18022 28445 18025 28479
rect 18059 28445 18101 28479
rect 18135 28445 18177 28479
rect 18211 28445 18253 28479
rect 18287 28445 18329 28479
rect 18363 28445 18405 28479
rect 18439 28461 18486 28479
rect 18520 28461 18556 28495
rect 18590 28461 18626 28495
rect 18660 28461 18696 28495
rect 18730 28461 18766 28495
rect 18800 28461 18836 28495
rect 18870 28461 18906 28495
rect 18940 28461 18976 28495
rect 19010 28461 19012 28495
rect 18439 28445 19012 28461
rect 18022 28427 19012 28445
rect 18022 28411 18486 28427
rect 18022 28377 18025 28411
rect 18059 28377 18101 28411
rect 18135 28377 18177 28411
rect 18211 28377 18253 28411
rect 18287 28377 18329 28411
rect 18363 28377 18405 28411
rect 18439 28393 18486 28411
rect 18520 28393 18556 28427
rect 18590 28393 18626 28427
rect 18660 28393 18696 28427
rect 18730 28393 18766 28427
rect 18800 28393 18836 28427
rect 18870 28393 18906 28427
rect 18940 28393 18976 28427
rect 19010 28393 19012 28427
rect 18439 28377 19012 28393
rect 18022 28359 19012 28377
rect 18022 28343 18486 28359
rect 18022 28309 18025 28343
rect 18059 28309 18101 28343
rect 18135 28309 18177 28343
rect 18211 28309 18253 28343
rect 18287 28309 18329 28343
rect 18363 28309 18405 28343
rect 18439 28325 18486 28343
rect 18520 28325 18556 28359
rect 18590 28325 18626 28359
rect 18660 28325 18696 28359
rect 18730 28325 18766 28359
rect 18800 28325 18836 28359
rect 18870 28325 18906 28359
rect 18940 28325 18976 28359
rect 19010 28325 19012 28359
rect 18439 28309 19012 28325
rect 18022 28291 19012 28309
rect 18022 28275 18486 28291
rect 18022 28241 18025 28275
rect 18059 28241 18101 28275
rect 18135 28241 18177 28275
rect 18211 28241 18253 28275
rect 18287 28241 18329 28275
rect 18363 28241 18405 28275
rect 18439 28257 18486 28275
rect 18520 28257 18556 28291
rect 18590 28257 18626 28291
rect 18660 28257 18696 28291
rect 18730 28257 18766 28291
rect 18800 28257 18836 28291
rect 18870 28257 18906 28291
rect 18940 28257 18976 28291
rect 19010 28257 19012 28291
rect 18439 28241 19012 28257
rect 18022 28223 19012 28241
rect 18022 28207 18486 28223
rect 18022 28173 18025 28207
rect 18059 28173 18101 28207
rect 18135 28173 18177 28207
rect 18211 28173 18253 28207
rect 18287 28173 18329 28207
rect 18363 28173 18405 28207
rect 18439 28189 18486 28207
rect 18520 28189 18556 28223
rect 18590 28189 18626 28223
rect 18660 28189 18696 28223
rect 18730 28189 18766 28223
rect 18800 28189 18836 28223
rect 18870 28189 18906 28223
rect 18940 28189 18976 28223
rect 19010 28189 19012 28223
rect 18439 28173 19012 28189
rect 18022 28155 19012 28173
rect 18022 28139 18486 28155
rect 18022 28105 18025 28139
rect 18059 28105 18101 28139
rect 18135 28105 18177 28139
rect 18211 28105 18253 28139
rect 18287 28105 18329 28139
rect 18363 28105 18405 28139
rect 18439 28121 18486 28139
rect 18520 28121 18556 28155
rect 18590 28121 18626 28155
rect 18660 28121 18696 28155
rect 18730 28121 18766 28155
rect 18800 28121 18836 28155
rect 18870 28121 18906 28155
rect 18940 28121 18976 28155
rect 19010 28121 19012 28155
rect 18439 28105 19012 28121
rect 18022 28087 19012 28105
rect 18022 28071 18486 28087
rect 18022 28037 18025 28071
rect 18059 28037 18101 28071
rect 18135 28037 18177 28071
rect 18211 28037 18253 28071
rect 18287 28037 18329 28071
rect 18363 28037 18405 28071
rect 18439 28053 18486 28071
rect 18520 28053 18556 28087
rect 18590 28053 18626 28087
rect 18660 28053 18696 28087
rect 18730 28053 18766 28087
rect 18800 28053 18836 28087
rect 18870 28053 18906 28087
rect 18940 28053 18976 28087
rect 19010 28053 19012 28087
rect 18439 28037 19012 28053
rect 18022 28019 19012 28037
rect 18022 28003 18486 28019
rect 18022 27969 18025 28003
rect 18059 27969 18101 28003
rect 18135 27969 18177 28003
rect 18211 27969 18253 28003
rect 18287 27969 18329 28003
rect 18363 27969 18405 28003
rect 18439 27985 18486 28003
rect 18520 27985 18556 28019
rect 18590 27985 18626 28019
rect 18660 27985 18696 28019
rect 18730 27985 18766 28019
rect 18800 27985 18836 28019
rect 18870 27985 18906 28019
rect 18940 27985 18976 28019
rect 19010 27985 19012 28019
rect 18439 27969 19012 27985
rect 18022 27951 19012 27969
rect 18022 27935 18486 27951
rect 18022 27901 18025 27935
rect 18059 27901 18101 27935
rect 18135 27901 18177 27935
rect 18211 27901 18253 27935
rect 18287 27901 18329 27935
rect 18363 27901 18405 27935
rect 18439 27917 18486 27935
rect 18520 27917 18556 27951
rect 18590 27917 18626 27951
rect 18660 27917 18696 27951
rect 18730 27917 18766 27951
rect 18800 27917 18836 27951
rect 18870 27917 18906 27951
rect 18940 27917 18976 27951
rect 19010 27917 19012 27951
rect 18439 27901 19012 27917
rect 18022 27883 19012 27901
rect 18022 27867 18486 27883
rect 18022 27833 18025 27867
rect 18059 27833 18101 27867
rect 18135 27833 18177 27867
rect 18211 27833 18253 27867
rect 18287 27833 18329 27867
rect 18363 27833 18405 27867
rect 18439 27849 18486 27867
rect 18520 27849 18556 27883
rect 18590 27849 18626 27883
rect 18660 27849 18696 27883
rect 18730 27849 18766 27883
rect 18800 27849 18836 27883
rect 18870 27849 18906 27883
rect 18940 27849 18976 27883
rect 19010 27849 19012 27883
rect 18439 27833 19012 27849
rect 18022 27815 19012 27833
rect 18022 27799 18486 27815
rect 18022 27765 18025 27799
rect 18059 27765 18101 27799
rect 18135 27765 18177 27799
rect 18211 27765 18253 27799
rect 18287 27765 18329 27799
rect 18363 27765 18405 27799
rect 18439 27781 18486 27799
rect 18520 27781 18556 27815
rect 18590 27781 18626 27815
rect 18660 27781 18696 27815
rect 18730 27781 18766 27815
rect 18800 27781 18836 27815
rect 18870 27781 18906 27815
rect 18940 27781 18976 27815
rect 19010 27781 19012 27815
rect 18439 27765 19012 27781
rect 18022 27747 19012 27765
rect 18022 27731 18486 27747
rect 18022 27697 18025 27731
rect 18059 27697 18101 27731
rect 18135 27697 18177 27731
rect 18211 27697 18253 27731
rect 18287 27697 18329 27731
rect 18363 27697 18405 27731
rect 18439 27713 18486 27731
rect 18520 27713 18556 27747
rect 18590 27713 18626 27747
rect 18660 27713 18696 27747
rect 18730 27713 18766 27747
rect 18800 27713 18836 27747
rect 18870 27713 18906 27747
rect 18940 27713 18976 27747
rect 19010 27713 19012 27747
rect 18439 27697 19012 27713
rect 18022 27679 19012 27697
rect 18022 27663 18486 27679
rect 18022 27629 18025 27663
rect 18059 27629 18101 27663
rect 18135 27629 18177 27663
rect 18211 27629 18253 27663
rect 18287 27629 18329 27663
rect 18363 27629 18405 27663
rect 18439 27645 18486 27663
rect 18520 27645 18556 27679
rect 18590 27645 18626 27679
rect 18660 27645 18696 27679
rect 18730 27645 18766 27679
rect 18800 27645 18836 27679
rect 18870 27645 18906 27679
rect 18940 27645 18976 27679
rect 19010 27645 19012 27679
rect 18439 27629 19012 27645
rect 18022 27611 19012 27629
rect 18022 27595 18486 27611
rect 18022 27561 18025 27595
rect 18059 27561 18101 27595
rect 18135 27561 18177 27595
rect 18211 27561 18253 27595
rect 18287 27561 18329 27595
rect 18363 27561 18405 27595
rect 18439 27577 18486 27595
rect 18520 27577 18556 27611
rect 18590 27577 18626 27611
rect 18660 27577 18696 27611
rect 18730 27577 18766 27611
rect 18800 27577 18836 27611
rect 18870 27577 18906 27611
rect 18940 27577 18976 27611
rect 19010 27577 19012 27611
rect 18439 27561 19012 27577
rect 18022 27543 19012 27561
rect 18022 27527 18486 27543
rect 18022 27493 18025 27527
rect 18059 27493 18101 27527
rect 18135 27493 18177 27527
rect 18211 27493 18253 27527
rect 18287 27493 18329 27527
rect 18363 27493 18405 27527
rect 18439 27509 18486 27527
rect 18520 27509 18556 27543
rect 18590 27509 18626 27543
rect 18660 27509 18696 27543
rect 18730 27509 18766 27543
rect 18800 27509 18836 27543
rect 18870 27509 18906 27543
rect 18940 27509 18976 27543
rect 19010 27509 19012 27543
rect 18439 27493 19012 27509
rect 18022 27475 19012 27493
rect 18022 27459 18486 27475
rect 18022 27425 18025 27459
rect 18059 27425 18101 27459
rect 18135 27425 18177 27459
rect 18211 27425 18253 27459
rect 18287 27425 18329 27459
rect 18363 27425 18405 27459
rect 18439 27441 18486 27459
rect 18520 27441 18556 27475
rect 18590 27441 18626 27475
rect 18660 27441 18696 27475
rect 18730 27441 18766 27475
rect 18800 27441 18836 27475
rect 18870 27441 18906 27475
rect 18940 27441 18976 27475
rect 19010 27441 19012 27475
rect 18439 27425 19012 27441
rect 18022 27407 19012 27425
rect 18022 27391 18486 27407
rect 18022 27357 18025 27391
rect 18059 27357 18101 27391
rect 18135 27357 18177 27391
rect 18211 27357 18253 27391
rect 18287 27357 18329 27391
rect 18363 27357 18405 27391
rect 18439 27373 18486 27391
rect 18520 27373 18556 27407
rect 18590 27373 18626 27407
rect 18660 27373 18696 27407
rect 18730 27373 18766 27407
rect 18800 27373 18836 27407
rect 18870 27373 18906 27407
rect 18940 27373 18976 27407
rect 19010 27373 19012 27407
rect 18439 27357 19012 27373
rect 18022 27339 19012 27357
rect 18022 27323 18486 27339
rect 18022 27289 18025 27323
rect 18059 27289 18101 27323
rect 18135 27289 18177 27323
rect 18211 27289 18253 27323
rect 18287 27289 18329 27323
rect 18363 27289 18405 27323
rect 18439 27305 18486 27323
rect 18520 27305 18556 27339
rect 18590 27305 18626 27339
rect 18660 27305 18696 27339
rect 18730 27305 18766 27339
rect 18800 27305 18836 27339
rect 18870 27305 18906 27339
rect 18940 27305 18976 27339
rect 19010 27305 19012 27339
rect 18439 27289 19012 27305
rect 18022 27271 19012 27289
rect 18022 27255 18486 27271
rect 18022 27221 18025 27255
rect 18059 27221 18101 27255
rect 18135 27221 18177 27255
rect 18211 27221 18253 27255
rect 18287 27221 18329 27255
rect 18363 27221 18405 27255
rect 18439 27237 18486 27255
rect 18520 27237 18556 27271
rect 18590 27237 18626 27271
rect 18660 27237 18696 27271
rect 18730 27237 18766 27271
rect 18800 27237 18836 27271
rect 18870 27237 18906 27271
rect 18940 27237 18976 27271
rect 19010 27237 19012 27271
rect 18439 27221 19012 27237
rect 18022 27203 19012 27221
rect 18022 27187 18486 27203
rect 18022 27153 18025 27187
rect 18059 27153 18101 27187
rect 18135 27153 18177 27187
rect 18211 27153 18253 27187
rect 18287 27153 18329 27187
rect 18363 27153 18405 27187
rect 18439 27169 18486 27187
rect 18520 27169 18556 27203
rect 18590 27169 18626 27203
rect 18660 27169 18696 27203
rect 18730 27169 18766 27203
rect 18800 27169 18836 27203
rect 18870 27169 18906 27203
rect 18940 27169 18976 27203
rect 19010 27169 19012 27203
rect 18439 27153 19012 27169
rect 18022 27135 19012 27153
rect 18022 27119 18486 27135
rect 999 27079 1732 27103
rect 999 27045 1057 27079
rect 1091 27045 1125 27079
rect 1159 27045 1193 27079
rect 1227 27045 1261 27079
rect 1295 27045 1329 27079
rect 1363 27045 1397 27079
rect 1431 27045 1465 27079
rect 1499 27045 1533 27079
rect 1567 27045 1601 27079
rect 1635 27045 1669 27079
rect 1703 27045 1732 27079
rect 999 27010 1732 27045
rect 999 26976 1057 27010
rect 1091 26976 1125 27010
rect 1159 26976 1193 27010
rect 1227 26976 1261 27010
rect 1295 26976 1329 27010
rect 1363 26976 1397 27010
rect 1431 26976 1465 27010
rect 1499 26976 1533 27010
rect 1567 26976 1601 27010
rect 1635 26976 1669 27010
rect 1703 26976 1732 27010
rect 999 26941 1732 26976
rect 999 26907 1057 26941
rect 1091 26907 1125 26941
rect 1159 26907 1193 26941
rect 1227 26907 1261 26941
rect 1295 26907 1329 26941
rect 1363 26907 1397 26941
rect 1431 26907 1465 26941
rect 1499 26907 1533 26941
rect 1567 26907 1601 26941
rect 1635 26907 1669 26941
rect 1703 26907 1732 26941
rect 999 26872 1732 26907
rect 999 26838 1057 26872
rect 1091 26838 1125 26872
rect 1159 26838 1193 26872
rect 1227 26838 1261 26872
rect 1295 26838 1329 26872
rect 1363 26838 1397 26872
rect 1431 26838 1465 26872
rect 1499 26838 1533 26872
rect 1567 26838 1601 26872
rect 1635 26838 1669 26872
rect 1703 26838 1732 26872
rect 999 26803 1732 26838
rect 999 26769 1057 26803
rect 1091 26769 1125 26803
rect 1159 26769 1193 26803
rect 1227 26769 1261 26803
rect 1295 26769 1329 26803
rect 1363 26769 1397 26803
rect 1431 26769 1465 26803
rect 1499 26769 1533 26803
rect 1567 26769 1601 26803
rect 1635 26769 1669 26803
rect 1703 26769 1732 26803
rect 999 26734 1732 26769
rect 999 26700 1057 26734
rect 1091 26700 1125 26734
rect 1159 26700 1193 26734
rect 1227 26700 1261 26734
rect 1295 26700 1329 26734
rect 1363 26700 1397 26734
rect 1431 26700 1465 26734
rect 1499 26700 1533 26734
rect 1567 26700 1601 26734
rect 1635 26700 1669 26734
rect 1703 26700 1732 26734
rect 999 26665 1732 26700
rect 999 26631 1057 26665
rect 1091 26631 1125 26665
rect 1159 26631 1193 26665
rect 1227 26631 1261 26665
rect 1295 26631 1329 26665
rect 1363 26631 1397 26665
rect 1431 26631 1465 26665
rect 1499 26631 1533 26665
rect 1567 26631 1601 26665
rect 1635 26631 1669 26665
rect 1703 26631 1732 26665
rect 999 26596 1732 26631
rect 999 26562 1057 26596
rect 1091 26562 1125 26596
rect 1159 26562 1193 26596
rect 1227 26562 1261 26596
rect 1295 26562 1329 26596
rect 1363 26562 1397 26596
rect 1431 26562 1465 26596
rect 1499 26562 1533 26596
rect 1567 26562 1601 26596
rect 1635 26562 1669 26596
rect 1703 26562 1732 26596
rect 999 26527 1732 26562
rect 999 26493 1057 26527
rect 1091 26493 1125 26527
rect 1159 26493 1193 26527
rect 1227 26493 1261 26527
rect 1295 26493 1329 26527
rect 1363 26493 1397 26527
rect 1431 26493 1465 26527
rect 1499 26493 1533 26527
rect 1567 26493 1601 26527
rect 1635 26493 1669 26527
rect 1703 26493 1732 26527
rect 999 26458 1732 26493
rect 999 26424 1057 26458
rect 1091 26424 1125 26458
rect 1159 26424 1193 26458
rect 1227 26424 1261 26458
rect 1295 26424 1329 26458
rect 1363 26424 1397 26458
rect 1431 26424 1465 26458
rect 1499 26424 1533 26458
rect 1567 26424 1601 26458
rect 1635 26424 1669 26458
rect 1703 26424 1732 26458
rect 999 26389 1732 26424
rect 999 26355 1057 26389
rect 1091 26355 1125 26389
rect 1159 26355 1193 26389
rect 1227 26355 1261 26389
rect 1295 26355 1329 26389
rect 1363 26355 1397 26389
rect 1431 26355 1465 26389
rect 1499 26355 1533 26389
rect 1567 26355 1601 26389
rect 1635 26355 1669 26389
rect 1703 26355 1732 26389
rect 999 26320 1732 26355
rect 999 26286 1057 26320
rect 1091 26286 1125 26320
rect 1159 26286 1193 26320
rect 1227 26286 1261 26320
rect 1295 26286 1329 26320
rect 1363 26286 1397 26320
rect 1431 26286 1465 26320
rect 1499 26286 1533 26320
rect 1567 26286 1601 26320
rect 1635 26286 1669 26320
rect 1703 26286 1732 26320
rect 999 26251 1732 26286
rect 999 26217 1057 26251
rect 1091 26217 1125 26251
rect 1159 26217 1193 26251
rect 1227 26217 1261 26251
rect 1295 26217 1329 26251
rect 1363 26217 1397 26251
rect 1431 26217 1465 26251
rect 1499 26217 1533 26251
rect 1567 26217 1601 26251
rect 1635 26217 1669 26251
rect 1703 26217 1732 26251
rect 999 26182 1732 26217
rect 999 26148 1057 26182
rect 1091 26148 1125 26182
rect 1159 26148 1193 26182
rect 1227 26148 1261 26182
rect 1295 26148 1329 26182
rect 1363 26148 1397 26182
rect 1431 26148 1465 26182
rect 1499 26148 1533 26182
rect 1567 26148 1601 26182
rect 1635 26148 1669 26182
rect 1703 26148 1732 26182
rect 999 26113 1732 26148
rect 999 26079 1057 26113
rect 1091 26079 1125 26113
rect 1159 26079 1193 26113
rect 1227 26079 1261 26113
rect 1295 26079 1329 26113
rect 1363 26079 1397 26113
rect 1431 26079 1465 26113
rect 1499 26079 1533 26113
rect 1567 26079 1601 26113
rect 1635 26079 1669 26113
rect 1703 26079 1732 26113
rect 999 26044 1732 26079
rect 999 26010 1057 26044
rect 1091 26010 1125 26044
rect 1159 26010 1193 26044
rect 1227 26010 1261 26044
rect 1295 26010 1329 26044
rect 1363 26010 1397 26044
rect 1431 26010 1465 26044
rect 1499 26010 1533 26044
rect 1567 26010 1601 26044
rect 1635 26010 1669 26044
rect 1703 26010 1732 26044
rect 999 25975 1732 26010
rect 999 25941 1057 25975
rect 1091 25941 1125 25975
rect 1159 25941 1193 25975
rect 1227 25941 1261 25975
rect 1295 25941 1329 25975
rect 1363 25941 1397 25975
rect 1431 25941 1465 25975
rect 1499 25941 1533 25975
rect 1567 25941 1601 25975
rect 1635 25941 1669 25975
rect 1703 25941 1732 25975
rect 999 25906 1732 25941
rect 999 25872 1057 25906
rect 1091 25872 1125 25906
rect 1159 25872 1193 25906
rect 1227 25872 1261 25906
rect 1295 25872 1329 25906
rect 1363 25872 1397 25906
rect 1431 25872 1465 25906
rect 1499 25872 1533 25906
rect 1567 25872 1601 25906
rect 1635 25872 1669 25906
rect 1703 25872 1732 25906
rect 999 25837 1732 25872
rect 999 25803 1057 25837
rect 1091 25803 1125 25837
rect 1159 25803 1193 25837
rect 1227 25803 1261 25837
rect 1295 25803 1329 25837
rect 1363 25803 1397 25837
rect 1431 25803 1465 25837
rect 1499 25803 1533 25837
rect 1567 25803 1601 25837
rect 1635 25803 1669 25837
rect 1703 25803 1732 25837
rect 999 25768 1732 25803
rect 999 25734 1057 25768
rect 1091 25734 1125 25768
rect 1159 25734 1193 25768
rect 1227 25734 1261 25768
rect 1295 25734 1329 25768
rect 1363 25734 1397 25768
rect 1431 25734 1465 25768
rect 1499 25734 1533 25768
rect 1567 25734 1601 25768
rect 1635 25734 1669 25768
rect 1703 25734 1732 25768
rect 999 25699 1732 25734
rect 999 25665 1057 25699
rect 1091 25665 1125 25699
rect 1159 25665 1193 25699
rect 1227 25665 1261 25699
rect 1295 25665 1329 25699
rect 1363 25665 1397 25699
rect 1431 25665 1465 25699
rect 1499 25665 1533 25699
rect 1567 25665 1601 25699
rect 1635 25665 1669 25699
rect 1703 25665 1732 25699
rect 999 25630 1732 25665
rect 999 25596 1057 25630
rect 1091 25596 1125 25630
rect 1159 25596 1193 25630
rect 1227 25596 1261 25630
rect 1295 25596 1329 25630
rect 1363 25596 1397 25630
rect 1431 25596 1465 25630
rect 1499 25596 1533 25630
rect 1567 25596 1601 25630
rect 1635 25596 1669 25630
rect 1703 25596 1732 25630
rect 999 25561 1732 25596
rect 999 25527 1057 25561
rect 1091 25527 1125 25561
rect 1159 25527 1193 25561
rect 1227 25527 1261 25561
rect 1295 25527 1329 25561
rect 1363 25527 1397 25561
rect 1431 25527 1465 25561
rect 1499 25527 1533 25561
rect 1567 25527 1601 25561
rect 1635 25527 1669 25561
rect 1703 25527 1732 25561
rect 999 25492 1732 25527
rect 999 25458 1057 25492
rect 1091 25458 1125 25492
rect 1159 25458 1193 25492
rect 1227 25458 1261 25492
rect 1295 25458 1329 25492
rect 1363 25458 1397 25492
rect 1431 25458 1465 25492
rect 1499 25458 1533 25492
rect 1567 25458 1601 25492
rect 1635 25458 1669 25492
rect 1703 25458 1732 25492
rect 999 25423 1732 25458
rect 999 25389 1057 25423
rect 1091 25389 1125 25423
rect 1159 25389 1193 25423
rect 1227 25389 1261 25423
rect 1295 25389 1329 25423
rect 1363 25389 1397 25423
rect 1431 25389 1465 25423
rect 1499 25389 1533 25423
rect 1567 25389 1601 25423
rect 1635 25389 1669 25423
rect 1703 25389 1732 25423
rect 999 25354 1732 25389
rect 999 25320 1057 25354
rect 1091 25320 1125 25354
rect 1159 25320 1193 25354
rect 1227 25320 1261 25354
rect 1295 25320 1329 25354
rect 1363 25320 1397 25354
rect 1431 25320 1465 25354
rect 1499 25320 1533 25354
rect 1567 25320 1601 25354
rect 1635 25320 1669 25354
rect 1703 25320 1732 25354
rect 999 25285 1732 25320
rect 999 25251 1057 25285
rect 1091 25251 1125 25285
rect 1159 25251 1193 25285
rect 1227 25251 1261 25285
rect 1295 25251 1329 25285
rect 1363 25251 1397 25285
rect 1431 25251 1465 25285
rect 1499 25251 1533 25285
rect 1567 25251 1601 25285
rect 1635 25251 1669 25285
rect 1703 25251 1732 25285
rect 999 25216 1732 25251
rect 999 25182 1057 25216
rect 1091 25182 1125 25216
rect 1159 25182 1193 25216
rect 1227 25182 1261 25216
rect 1295 25182 1329 25216
rect 1363 25182 1397 25216
rect 1431 25182 1465 25216
rect 1499 25182 1533 25216
rect 1567 25182 1601 25216
rect 1635 25182 1669 25216
rect 1703 25182 1732 25216
rect 999 25147 1732 25182
rect 999 25113 1057 25147
rect 1091 25113 1125 25147
rect 1159 25113 1193 25147
rect 1227 25113 1261 25147
rect 1295 25113 1329 25147
rect 1363 25113 1397 25147
rect 1431 25113 1465 25147
rect 1499 25113 1533 25147
rect 1567 25113 1601 25147
rect 1635 25113 1669 25147
rect 1703 25113 1732 25147
rect 999 25077 1732 25113
rect 999 25043 1057 25077
rect 1091 25043 1125 25077
rect 1159 25043 1193 25077
rect 1227 25043 1261 25077
rect 1295 25043 1329 25077
rect 1363 25043 1397 25077
rect 1431 25043 1465 25077
rect 1499 25043 1533 25077
rect 1567 25043 1601 25077
rect 1635 25043 1669 25077
rect 1703 25043 1732 25077
rect 999 25007 1732 25043
rect 999 24973 1057 25007
rect 1091 24973 1125 25007
rect 1159 24973 1193 25007
rect 1227 24973 1261 25007
rect 1295 24973 1329 25007
rect 1363 24973 1397 25007
rect 1431 24973 1465 25007
rect 1499 24973 1533 25007
rect 1567 24973 1601 25007
rect 1635 24973 1669 25007
rect 1703 24973 1732 25007
rect 999 24937 1732 24973
rect 999 24903 1057 24937
rect 1091 24903 1125 24937
rect 1159 24903 1193 24937
rect 1227 24903 1261 24937
rect 1295 24903 1329 24937
rect 1363 24903 1397 24937
rect 1431 24903 1465 24937
rect 1499 24903 1533 24937
rect 1567 24903 1601 24937
rect 1635 24903 1669 24937
rect 1703 24903 1732 24937
rect 999 24867 1732 24903
rect 999 24833 1057 24867
rect 1091 24833 1125 24867
rect 1159 24833 1193 24867
rect 1227 24833 1261 24867
rect 1295 24833 1329 24867
rect 1363 24833 1397 24867
rect 1431 24833 1465 24867
rect 1499 24833 1533 24867
rect 1567 24833 1601 24867
rect 1635 24833 1669 24867
rect 1703 24833 1732 24867
rect 999 24797 1732 24833
rect 999 24763 1057 24797
rect 1091 24763 1125 24797
rect 1159 24763 1193 24797
rect 1227 24763 1261 24797
rect 1295 24763 1329 24797
rect 1363 24763 1397 24797
rect 1431 24763 1465 24797
rect 1499 24763 1533 24797
rect 1567 24763 1601 24797
rect 1635 24763 1669 24797
rect 1703 24763 1732 24797
rect 999 24727 1732 24763
rect 999 24693 1057 24727
rect 1091 24693 1125 24727
rect 1159 24693 1193 24727
rect 1227 24693 1261 24727
rect 1295 24693 1329 24727
rect 1363 24693 1397 24727
rect 1431 24693 1465 24727
rect 1499 24693 1533 24727
rect 1567 24693 1601 24727
rect 1635 24693 1669 24727
rect 1703 24693 1732 24727
rect 999 24657 1732 24693
rect 999 24623 1057 24657
rect 1091 24623 1125 24657
rect 1159 24623 1193 24657
rect 1227 24623 1261 24657
rect 1295 24623 1329 24657
rect 1363 24623 1397 24657
rect 1431 24623 1465 24657
rect 1499 24623 1533 24657
rect 1567 24623 1601 24657
rect 1635 24623 1669 24657
rect 1703 24623 1732 24657
rect 999 24587 1732 24623
rect 999 24553 1057 24587
rect 1091 24553 1125 24587
rect 1159 24553 1193 24587
rect 1227 24553 1261 24587
rect 1295 24553 1329 24587
rect 1363 24553 1397 24587
rect 1431 24553 1465 24587
rect 1499 24553 1533 24587
rect 1567 24553 1601 24587
rect 1635 24553 1669 24587
rect 1703 24553 1732 24587
rect 999 24517 1732 24553
rect 999 24483 1057 24517
rect 1091 24483 1125 24517
rect 1159 24483 1193 24517
rect 1227 24483 1261 24517
rect 1295 24483 1329 24517
rect 1363 24483 1397 24517
rect 1431 24483 1465 24517
rect 1499 24483 1533 24517
rect 1567 24483 1601 24517
rect 1635 24483 1669 24517
rect 1703 24483 1732 24517
rect 999 24447 1732 24483
rect 999 24413 1057 24447
rect 1091 24413 1125 24447
rect 1159 24413 1193 24447
rect 1227 24413 1261 24447
rect 1295 24413 1329 24447
rect 1363 24413 1397 24447
rect 1431 24413 1465 24447
rect 1499 24413 1533 24447
rect 1567 24413 1601 24447
rect 1635 24413 1669 24447
rect 1703 24413 1732 24447
rect 999 24377 1732 24413
rect 999 24343 1057 24377
rect 1091 24343 1125 24377
rect 1159 24343 1193 24377
rect 1227 24343 1261 24377
rect 1295 24343 1329 24377
rect 1363 24343 1397 24377
rect 1431 24343 1465 24377
rect 1499 24343 1533 24377
rect 1567 24343 1601 24377
rect 1635 24343 1669 24377
rect 1703 24343 1732 24377
rect 999 24307 1732 24343
rect 999 24273 1057 24307
rect 1091 24273 1125 24307
rect 1159 24273 1193 24307
rect 1227 24273 1261 24307
rect 1295 24273 1329 24307
rect 1363 24273 1397 24307
rect 1431 24273 1465 24307
rect 1499 24273 1533 24307
rect 1567 24273 1601 24307
rect 1635 24273 1669 24307
rect 1703 24273 1732 24307
rect 999 24237 1732 24273
rect 999 24203 1057 24237
rect 1091 24203 1125 24237
rect 1159 24203 1193 24237
rect 1227 24203 1261 24237
rect 1295 24203 1329 24237
rect 1363 24203 1397 24237
rect 1431 24203 1465 24237
rect 1499 24203 1533 24237
rect 1567 24203 1601 24237
rect 1635 24203 1669 24237
rect 1703 24203 1732 24237
rect 999 24167 1732 24203
rect 999 24133 1057 24167
rect 1091 24133 1125 24167
rect 1159 24133 1193 24167
rect 1227 24133 1261 24167
rect 1295 24133 1329 24167
rect 1363 24133 1397 24167
rect 1431 24133 1465 24167
rect 1499 24133 1533 24167
rect 1567 24133 1601 24167
rect 1635 24133 1669 24167
rect 1703 24133 1732 24167
rect 999 24097 1732 24133
rect 999 24063 1057 24097
rect 1091 24063 1125 24097
rect 1159 24063 1193 24097
rect 1227 24063 1261 24097
rect 1295 24063 1329 24097
rect 1363 24063 1397 24097
rect 1431 24063 1465 24097
rect 1499 24063 1533 24097
rect 1567 24063 1601 24097
rect 1635 24063 1669 24097
rect 1703 24063 1732 24097
rect 999 24027 1732 24063
rect 999 23993 1057 24027
rect 1091 23993 1125 24027
rect 1159 23993 1193 24027
rect 1227 23993 1261 24027
rect 1295 23993 1329 24027
rect 1363 23993 1397 24027
rect 1431 23993 1465 24027
rect 1499 23993 1533 24027
rect 1567 23993 1601 24027
rect 1635 23993 1669 24027
rect 1703 23993 1732 24027
rect 999 23957 1732 23993
rect 999 23923 1057 23957
rect 1091 23923 1125 23957
rect 1159 23923 1193 23957
rect 1227 23923 1261 23957
rect 1295 23923 1329 23957
rect 1363 23923 1397 23957
rect 1431 23923 1465 23957
rect 1499 23923 1533 23957
rect 1567 23923 1601 23957
rect 1635 23923 1669 23957
rect 1703 23923 1732 23957
rect 999 23887 1732 23923
rect 999 23853 1057 23887
rect 1091 23853 1125 23887
rect 1159 23853 1193 23887
rect 1227 23853 1261 23887
rect 1295 23853 1329 23887
rect 1363 23853 1397 23887
rect 1431 23853 1465 23887
rect 1499 23853 1533 23887
rect 1567 23853 1601 23887
rect 1635 23853 1669 23887
rect 1703 23853 1732 23887
rect 999 23829 1732 23853
rect 324 23803 1732 23829
rect 18022 27085 18025 27119
rect 18059 27085 18101 27119
rect 18135 27085 18177 27119
rect 18211 27085 18253 27119
rect 18287 27085 18329 27119
rect 18363 27085 18405 27119
rect 18439 27101 18486 27119
rect 18520 27101 18556 27135
rect 18590 27101 18626 27135
rect 18660 27101 18696 27135
rect 18730 27101 18766 27135
rect 18800 27101 18836 27135
rect 18870 27101 18906 27135
rect 18940 27101 18976 27135
rect 19010 27101 19012 27135
rect 18439 27085 19012 27101
rect 18022 27067 19012 27085
rect 18022 27051 18486 27067
rect 18022 27017 18025 27051
rect 18059 27017 18101 27051
rect 18135 27017 18177 27051
rect 18211 27017 18253 27051
rect 18287 27017 18329 27051
rect 18363 27017 18405 27051
rect 18439 27033 18486 27051
rect 18520 27033 18556 27067
rect 18590 27033 18626 27067
rect 18660 27033 18696 27067
rect 18730 27033 18766 27067
rect 18800 27033 18836 27067
rect 18870 27033 18906 27067
rect 18940 27033 18976 27067
rect 19010 27033 19012 27067
rect 18439 27017 19012 27033
rect 18022 26999 19012 27017
rect 18022 26983 18486 26999
rect 18022 26949 18025 26983
rect 18059 26949 18101 26983
rect 18135 26949 18177 26983
rect 18211 26949 18253 26983
rect 18287 26949 18329 26983
rect 18363 26949 18405 26983
rect 18439 26965 18486 26983
rect 18520 26965 18556 26999
rect 18590 26965 18626 26999
rect 18660 26965 18696 26999
rect 18730 26965 18766 26999
rect 18800 26965 18836 26999
rect 18870 26965 18906 26999
rect 18940 26965 18976 26999
rect 19010 26965 19012 26999
rect 18439 26949 19012 26965
rect 18022 26931 19012 26949
rect 18022 26915 18486 26931
rect 18022 26881 18025 26915
rect 18059 26881 18101 26915
rect 18135 26881 18177 26915
rect 18211 26881 18253 26915
rect 18287 26881 18329 26915
rect 18363 26881 18405 26915
rect 18439 26897 18486 26915
rect 18520 26897 18556 26931
rect 18590 26897 18626 26931
rect 18660 26897 18696 26931
rect 18730 26897 18766 26931
rect 18800 26897 18836 26931
rect 18870 26897 18906 26931
rect 18940 26897 18976 26931
rect 19010 26897 19012 26931
rect 18439 26881 19012 26897
rect 18022 26863 19012 26881
rect 18022 26847 18486 26863
rect 18022 26813 18025 26847
rect 18059 26813 18101 26847
rect 18135 26813 18177 26847
rect 18211 26813 18253 26847
rect 18287 26813 18329 26847
rect 18363 26813 18405 26847
rect 18439 26829 18486 26847
rect 18520 26829 18556 26863
rect 18590 26829 18626 26863
rect 18660 26829 18696 26863
rect 18730 26829 18766 26863
rect 18800 26829 18836 26863
rect 18870 26829 18906 26863
rect 18940 26829 18976 26863
rect 19010 26829 19012 26863
rect 18439 26813 19012 26829
rect 18022 26795 19012 26813
rect 18022 26779 18486 26795
rect 18022 26745 18025 26779
rect 18059 26745 18101 26779
rect 18135 26745 18177 26779
rect 18211 26745 18253 26779
rect 18287 26745 18329 26779
rect 18363 26745 18405 26779
rect 18439 26761 18486 26779
rect 18520 26761 18556 26795
rect 18590 26761 18626 26795
rect 18660 26761 18696 26795
rect 18730 26761 18766 26795
rect 18800 26761 18836 26795
rect 18870 26761 18906 26795
rect 18940 26761 18976 26795
rect 19010 26761 19012 26795
rect 18439 26745 19012 26761
rect 18022 26727 19012 26745
rect 18022 26711 18486 26727
rect 18022 26677 18025 26711
rect 18059 26677 18101 26711
rect 18135 26677 18177 26711
rect 18211 26677 18253 26711
rect 18287 26677 18329 26711
rect 18363 26677 18405 26711
rect 18439 26693 18486 26711
rect 18520 26693 18556 26727
rect 18590 26693 18626 26727
rect 18660 26693 18696 26727
rect 18730 26693 18766 26727
rect 18800 26693 18836 26727
rect 18870 26693 18906 26727
rect 18940 26693 18976 26727
rect 19010 26693 19012 26727
rect 18439 26677 19012 26693
rect 18022 26659 19012 26677
rect 18022 26643 18486 26659
rect 18022 26609 18025 26643
rect 18059 26609 18101 26643
rect 18135 26609 18177 26643
rect 18211 26609 18253 26643
rect 18287 26609 18329 26643
rect 18363 26609 18405 26643
rect 18439 26625 18486 26643
rect 18520 26625 18556 26659
rect 18590 26625 18626 26659
rect 18660 26625 18696 26659
rect 18730 26625 18766 26659
rect 18800 26625 18836 26659
rect 18870 26625 18906 26659
rect 18940 26625 18976 26659
rect 19010 26625 19012 26659
rect 18439 26609 19012 26625
rect 18022 26591 19012 26609
rect 18022 26575 18486 26591
rect 18022 26541 18025 26575
rect 18059 26541 18101 26575
rect 18135 26541 18177 26575
rect 18211 26541 18253 26575
rect 18287 26541 18329 26575
rect 18363 26541 18405 26575
rect 18439 26557 18486 26575
rect 18520 26557 18556 26591
rect 18590 26557 18626 26591
rect 18660 26557 18696 26591
rect 18730 26557 18766 26591
rect 18800 26557 18836 26591
rect 18870 26557 18906 26591
rect 18940 26557 18976 26591
rect 19010 26557 19012 26591
rect 18439 26541 19012 26557
rect 18022 26523 19012 26541
rect 18022 26507 18486 26523
rect 18022 26473 18025 26507
rect 18059 26473 18101 26507
rect 18135 26473 18177 26507
rect 18211 26473 18253 26507
rect 18287 26473 18329 26507
rect 18363 26473 18405 26507
rect 18439 26489 18486 26507
rect 18520 26489 18556 26523
rect 18590 26489 18626 26523
rect 18660 26489 18696 26523
rect 18730 26489 18766 26523
rect 18800 26489 18836 26523
rect 18870 26489 18906 26523
rect 18940 26489 18976 26523
rect 19010 26489 19012 26523
rect 18439 26473 19012 26489
rect 18022 26455 19012 26473
rect 18022 26439 18486 26455
rect 18022 26405 18025 26439
rect 18059 26405 18101 26439
rect 18135 26405 18177 26439
rect 18211 26405 18253 26439
rect 18287 26405 18329 26439
rect 18363 26405 18405 26439
rect 18439 26421 18486 26439
rect 18520 26421 18556 26455
rect 18590 26421 18626 26455
rect 18660 26421 18696 26455
rect 18730 26421 18766 26455
rect 18800 26421 18836 26455
rect 18870 26421 18906 26455
rect 18940 26421 18976 26455
rect 19010 26421 19012 26455
rect 18439 26405 19012 26421
rect 18022 26387 19012 26405
rect 18022 26371 18486 26387
rect 18022 26337 18025 26371
rect 18059 26337 18101 26371
rect 18135 26337 18177 26371
rect 18211 26337 18253 26371
rect 18287 26337 18329 26371
rect 18363 26337 18405 26371
rect 18439 26353 18486 26371
rect 18520 26353 18556 26387
rect 18590 26353 18626 26387
rect 18660 26353 18696 26387
rect 18730 26353 18766 26387
rect 18800 26353 18836 26387
rect 18870 26353 18906 26387
rect 18940 26353 18976 26387
rect 19010 26353 19012 26387
rect 18439 26337 19012 26353
rect 18022 26319 19012 26337
rect 18022 26303 18486 26319
rect 18022 26269 18025 26303
rect 18059 26269 18101 26303
rect 18135 26269 18177 26303
rect 18211 26269 18253 26303
rect 18287 26269 18329 26303
rect 18363 26269 18405 26303
rect 18439 26285 18486 26303
rect 18520 26285 18556 26319
rect 18590 26285 18626 26319
rect 18660 26285 18696 26319
rect 18730 26285 18766 26319
rect 18800 26285 18836 26319
rect 18870 26285 18906 26319
rect 18940 26285 18976 26319
rect 19010 26285 19012 26319
rect 18439 26269 19012 26285
rect 18022 26251 19012 26269
rect 18022 26235 18486 26251
rect 18022 26201 18025 26235
rect 18059 26201 18101 26235
rect 18135 26201 18177 26235
rect 18211 26201 18253 26235
rect 18287 26201 18329 26235
rect 18363 26201 18405 26235
rect 18439 26217 18486 26235
rect 18520 26217 18556 26251
rect 18590 26217 18626 26251
rect 18660 26217 18696 26251
rect 18730 26217 18766 26251
rect 18800 26217 18836 26251
rect 18870 26217 18906 26251
rect 18940 26217 18976 26251
rect 19010 26217 19012 26251
rect 18439 26201 19012 26217
rect 18022 26183 19012 26201
rect 18022 26167 18486 26183
rect 18022 26133 18025 26167
rect 18059 26133 18101 26167
rect 18135 26133 18177 26167
rect 18211 26133 18253 26167
rect 18287 26133 18329 26167
rect 18363 26133 18405 26167
rect 18439 26149 18486 26167
rect 18520 26149 18556 26183
rect 18590 26149 18626 26183
rect 18660 26149 18696 26183
rect 18730 26149 18766 26183
rect 18800 26149 18836 26183
rect 18870 26149 18906 26183
rect 18940 26149 18976 26183
rect 19010 26149 19012 26183
rect 18439 26133 19012 26149
rect 18022 26115 19012 26133
rect 18022 26099 18486 26115
rect 18022 26065 18025 26099
rect 18059 26065 18101 26099
rect 18135 26065 18177 26099
rect 18211 26065 18253 26099
rect 18287 26065 18329 26099
rect 18363 26065 18405 26099
rect 18439 26081 18486 26099
rect 18520 26081 18556 26115
rect 18590 26081 18626 26115
rect 18660 26081 18696 26115
rect 18730 26081 18766 26115
rect 18800 26081 18836 26115
rect 18870 26081 18906 26115
rect 18940 26081 18976 26115
rect 19010 26081 19012 26115
rect 18439 26065 19012 26081
rect 18022 26047 19012 26065
rect 18022 26031 18486 26047
rect 18022 25997 18025 26031
rect 18059 25997 18101 26031
rect 18135 25997 18177 26031
rect 18211 25997 18253 26031
rect 18287 25997 18329 26031
rect 18363 25997 18405 26031
rect 18439 26013 18486 26031
rect 18520 26013 18556 26047
rect 18590 26013 18626 26047
rect 18660 26013 18696 26047
rect 18730 26013 18766 26047
rect 18800 26013 18836 26047
rect 18870 26013 18906 26047
rect 18940 26013 18976 26047
rect 19010 26013 19012 26047
rect 18439 25997 19012 26013
rect 18022 25979 19012 25997
rect 18022 25963 18486 25979
rect 18022 25929 18025 25963
rect 18059 25929 18101 25963
rect 18135 25929 18177 25963
rect 18211 25929 18253 25963
rect 18287 25929 18329 25963
rect 18363 25929 18405 25963
rect 18439 25945 18486 25963
rect 18520 25945 18556 25979
rect 18590 25945 18626 25979
rect 18660 25945 18696 25979
rect 18730 25945 18766 25979
rect 18800 25945 18836 25979
rect 18870 25945 18906 25979
rect 18940 25945 18976 25979
rect 19010 25945 19012 25979
rect 18439 25929 19012 25945
rect 18022 25911 19012 25929
rect 18022 25895 18486 25911
rect 18022 25861 18025 25895
rect 18059 25861 18101 25895
rect 18135 25861 18177 25895
rect 18211 25861 18253 25895
rect 18287 25861 18329 25895
rect 18363 25861 18405 25895
rect 18439 25877 18486 25895
rect 18520 25877 18556 25911
rect 18590 25877 18626 25911
rect 18660 25877 18696 25911
rect 18730 25877 18766 25911
rect 18800 25877 18836 25911
rect 18870 25877 18906 25911
rect 18940 25877 18976 25911
rect 19010 25877 19012 25911
rect 18439 25861 19012 25877
rect 18022 25843 19012 25861
rect 18022 25827 18486 25843
rect 18022 25793 18025 25827
rect 18059 25793 18101 25827
rect 18135 25793 18177 25827
rect 18211 25793 18253 25827
rect 18287 25793 18329 25827
rect 18363 25793 18405 25827
rect 18439 25809 18486 25827
rect 18520 25809 18556 25843
rect 18590 25809 18626 25843
rect 18660 25809 18696 25843
rect 18730 25809 18766 25843
rect 18800 25809 18836 25843
rect 18870 25809 18906 25843
rect 18940 25809 18976 25843
rect 19010 25809 19012 25843
rect 18439 25793 19012 25809
rect 18022 25775 19012 25793
rect 18022 25759 18486 25775
rect 18022 25725 18025 25759
rect 18059 25725 18101 25759
rect 18135 25725 18177 25759
rect 18211 25725 18253 25759
rect 18287 25725 18329 25759
rect 18363 25725 18405 25759
rect 18439 25741 18486 25759
rect 18520 25741 18556 25775
rect 18590 25741 18626 25775
rect 18660 25741 18696 25775
rect 18730 25741 18766 25775
rect 18800 25741 18836 25775
rect 18870 25741 18906 25775
rect 18940 25741 18976 25775
rect 19010 25741 19012 25775
rect 18439 25725 19012 25741
rect 18022 25707 19012 25725
rect 18022 25691 18486 25707
rect 18022 25657 18025 25691
rect 18059 25657 18101 25691
rect 18135 25657 18177 25691
rect 18211 25657 18253 25691
rect 18287 25657 18329 25691
rect 18363 25657 18405 25691
rect 18439 25673 18486 25691
rect 18520 25673 18556 25707
rect 18590 25673 18626 25707
rect 18660 25673 18696 25707
rect 18730 25673 18766 25707
rect 18800 25673 18836 25707
rect 18870 25673 18906 25707
rect 18940 25673 18976 25707
rect 19010 25673 19012 25707
rect 18439 25657 19012 25673
rect 18022 25638 19012 25657
rect 18022 25623 18486 25638
rect 18022 25589 18025 25623
rect 18059 25589 18101 25623
rect 18135 25589 18177 25623
rect 18211 25589 18253 25623
rect 18287 25589 18329 25623
rect 18363 25589 18405 25623
rect 18439 25604 18486 25623
rect 18520 25604 18556 25638
rect 18590 25604 18626 25638
rect 18660 25604 18696 25638
rect 18730 25604 18766 25638
rect 18800 25604 18836 25638
rect 18870 25604 18906 25638
rect 18940 25604 18976 25638
rect 19010 25604 19012 25638
rect 18439 25589 19012 25604
rect 18022 25569 19012 25589
rect 18022 25555 18486 25569
rect 18022 25521 18025 25555
rect 18059 25521 18101 25555
rect 18135 25521 18177 25555
rect 18211 25521 18253 25555
rect 18287 25521 18329 25555
rect 18363 25521 18405 25555
rect 18439 25535 18486 25555
rect 18520 25535 18556 25569
rect 18590 25535 18626 25569
rect 18660 25535 18696 25569
rect 18730 25535 18766 25569
rect 18800 25535 18836 25569
rect 18870 25535 18906 25569
rect 18940 25535 18976 25569
rect 19010 25535 19012 25569
rect 18439 25521 19012 25535
rect 18022 25500 19012 25521
rect 18022 25487 18486 25500
rect 18022 25453 18025 25487
rect 18059 25453 18101 25487
rect 18135 25453 18177 25487
rect 18211 25453 18253 25487
rect 18287 25453 18329 25487
rect 18363 25453 18405 25487
rect 18439 25466 18486 25487
rect 18520 25466 18556 25500
rect 18590 25466 18626 25500
rect 18660 25466 18696 25500
rect 18730 25466 18766 25500
rect 18800 25466 18836 25500
rect 18870 25466 18906 25500
rect 18940 25466 18976 25500
rect 19010 25466 19012 25500
rect 18439 25453 19012 25466
rect 18022 25431 19012 25453
rect 18022 25419 18486 25431
rect 18022 25385 18025 25419
rect 18059 25385 18101 25419
rect 18135 25385 18177 25419
rect 18211 25385 18253 25419
rect 18287 25385 18329 25419
rect 18363 25385 18405 25419
rect 18439 25397 18486 25419
rect 18520 25397 18556 25431
rect 18590 25397 18626 25431
rect 18660 25397 18696 25431
rect 18730 25397 18766 25431
rect 18800 25397 18836 25431
rect 18870 25397 18906 25431
rect 18940 25397 18976 25431
rect 19010 25397 19012 25431
rect 18439 25385 19012 25397
rect 18022 25362 19012 25385
rect 18022 25351 18486 25362
rect 18022 25317 18025 25351
rect 18059 25317 18101 25351
rect 18135 25317 18177 25351
rect 18211 25317 18253 25351
rect 18287 25317 18329 25351
rect 18363 25317 18405 25351
rect 18439 25328 18486 25351
rect 18520 25328 18556 25362
rect 18590 25328 18626 25362
rect 18660 25328 18696 25362
rect 18730 25328 18766 25362
rect 18800 25328 18836 25362
rect 18870 25328 18906 25362
rect 18940 25328 18976 25362
rect 19010 25328 19012 25362
rect 18439 25317 19012 25328
rect 18022 25293 19012 25317
rect 18022 25283 18486 25293
rect 18022 25249 18025 25283
rect 18059 25249 18101 25283
rect 18135 25249 18177 25283
rect 18211 25249 18253 25283
rect 18287 25249 18329 25283
rect 18363 25249 18405 25283
rect 18439 25259 18486 25283
rect 18520 25259 18556 25293
rect 18590 25259 18626 25293
rect 18660 25259 18696 25293
rect 18730 25259 18766 25293
rect 18800 25259 18836 25293
rect 18870 25259 18906 25293
rect 18940 25259 18976 25293
rect 19010 25259 19012 25293
rect 18439 25249 19012 25259
rect 18022 25224 19012 25249
rect 18022 25214 18486 25224
rect 18022 25180 18025 25214
rect 18059 25180 18101 25214
rect 18135 25180 18177 25214
rect 18211 25180 18253 25214
rect 18287 25180 18329 25214
rect 18363 25180 18405 25214
rect 18439 25190 18486 25214
rect 18520 25190 18556 25224
rect 18590 25190 18626 25224
rect 18660 25190 18696 25224
rect 18730 25190 18766 25224
rect 18800 25190 18836 25224
rect 18870 25190 18906 25224
rect 18940 25190 18976 25224
rect 19010 25190 19012 25224
rect 18439 25180 19012 25190
rect 18022 25155 19012 25180
rect 18022 25145 18486 25155
rect 18022 25111 18025 25145
rect 18059 25111 18101 25145
rect 18135 25111 18177 25145
rect 18211 25111 18253 25145
rect 18287 25111 18329 25145
rect 18363 25111 18405 25145
rect 18439 25121 18486 25145
rect 18520 25121 18556 25155
rect 18590 25121 18626 25155
rect 18660 25121 18696 25155
rect 18730 25121 18766 25155
rect 18800 25121 18836 25155
rect 18870 25121 18906 25155
rect 18940 25121 18976 25155
rect 19010 25121 19012 25155
rect 18439 25111 19012 25121
rect 18022 25086 19012 25111
rect 18022 25076 18486 25086
rect 18022 25042 18025 25076
rect 18059 25042 18101 25076
rect 18135 25042 18177 25076
rect 18211 25042 18253 25076
rect 18287 25042 18329 25076
rect 18363 25042 18405 25076
rect 18439 25052 18486 25076
rect 18520 25052 18556 25086
rect 18590 25052 18626 25086
rect 18660 25052 18696 25086
rect 18730 25052 18766 25086
rect 18800 25052 18836 25086
rect 18870 25052 18906 25086
rect 18940 25052 18976 25086
rect 19010 25052 19012 25086
rect 18439 25042 19012 25052
rect 18022 25017 19012 25042
rect 18022 25007 18486 25017
rect 18022 24973 18025 25007
rect 18059 24973 18101 25007
rect 18135 24973 18177 25007
rect 18211 24973 18253 25007
rect 18287 24973 18329 25007
rect 18363 24973 18405 25007
rect 18439 24983 18486 25007
rect 18520 24983 18556 25017
rect 18590 24983 18626 25017
rect 18660 24983 18696 25017
rect 18730 24983 18766 25017
rect 18800 24983 18836 25017
rect 18870 24983 18906 25017
rect 18940 24983 18976 25017
rect 19010 24983 19012 25017
rect 18439 24973 19012 24983
rect 18022 24948 19012 24973
rect 18022 24938 18486 24948
rect 18022 24904 18025 24938
rect 18059 24904 18101 24938
rect 18135 24904 18177 24938
rect 18211 24904 18253 24938
rect 18287 24904 18329 24938
rect 18363 24904 18405 24938
rect 18439 24914 18486 24938
rect 18520 24914 18556 24948
rect 18590 24914 18626 24948
rect 18660 24914 18696 24948
rect 18730 24914 18766 24948
rect 18800 24914 18836 24948
rect 18870 24914 18906 24948
rect 18940 24914 18976 24948
rect 19010 24914 19012 24948
rect 18439 24904 19012 24914
rect 18022 24879 19012 24904
rect 18022 24869 18486 24879
rect 18022 24835 18025 24869
rect 18059 24835 18101 24869
rect 18135 24835 18177 24869
rect 18211 24835 18253 24869
rect 18287 24835 18329 24869
rect 18363 24835 18405 24869
rect 18439 24845 18486 24869
rect 18520 24845 18556 24879
rect 18590 24845 18626 24879
rect 18660 24845 18696 24879
rect 18730 24845 18766 24879
rect 18800 24845 18836 24879
rect 18870 24845 18906 24879
rect 18940 24845 18976 24879
rect 19010 24845 19012 24879
rect 18439 24835 19012 24845
rect 18022 24810 19012 24835
rect 18022 24800 18486 24810
rect 18022 24766 18025 24800
rect 18059 24766 18101 24800
rect 18135 24766 18177 24800
rect 18211 24766 18253 24800
rect 18287 24766 18329 24800
rect 18363 24766 18405 24800
rect 18439 24776 18486 24800
rect 18520 24776 18556 24810
rect 18590 24776 18626 24810
rect 18660 24776 18696 24810
rect 18730 24776 18766 24810
rect 18800 24776 18836 24810
rect 18870 24776 18906 24810
rect 18940 24776 18976 24810
rect 19010 24776 19012 24810
rect 18439 24766 19012 24776
rect 18022 24741 19012 24766
rect 18022 24731 18486 24741
rect 18022 24697 18025 24731
rect 18059 24697 18101 24731
rect 18135 24697 18177 24731
rect 18211 24697 18253 24731
rect 18287 24697 18329 24731
rect 18363 24697 18405 24731
rect 18439 24707 18486 24731
rect 18520 24707 18556 24741
rect 18590 24707 18626 24741
rect 18660 24707 18696 24741
rect 18730 24707 18766 24741
rect 18800 24707 18836 24741
rect 18870 24707 18906 24741
rect 18940 24707 18976 24741
rect 19010 24707 19012 24741
rect 18439 24697 19012 24707
rect 18022 24672 19012 24697
rect 18022 24662 18486 24672
rect 18022 24628 18025 24662
rect 18059 24628 18101 24662
rect 18135 24628 18177 24662
rect 18211 24628 18253 24662
rect 18287 24628 18329 24662
rect 18363 24628 18405 24662
rect 18439 24638 18486 24662
rect 18520 24638 18556 24672
rect 18590 24638 18626 24672
rect 18660 24638 18696 24672
rect 18730 24638 18766 24672
rect 18800 24638 18836 24672
rect 18870 24638 18906 24672
rect 18940 24638 18976 24672
rect 19010 24638 19012 24672
rect 18439 24628 19012 24638
rect 18022 24603 19012 24628
rect 18022 24593 18486 24603
rect 18022 24559 18025 24593
rect 18059 24559 18101 24593
rect 18135 24559 18177 24593
rect 18211 24559 18253 24593
rect 18287 24559 18329 24593
rect 18363 24559 18405 24593
rect 18439 24569 18486 24593
rect 18520 24569 18556 24603
rect 18590 24569 18626 24603
rect 18660 24569 18696 24603
rect 18730 24569 18766 24603
rect 18800 24569 18836 24603
rect 18870 24569 18906 24603
rect 18940 24569 18976 24603
rect 19010 24569 19012 24603
rect 18439 24559 19012 24569
rect 18022 24534 19012 24559
rect 18022 24524 18486 24534
rect 18022 24490 18025 24524
rect 18059 24490 18101 24524
rect 18135 24490 18177 24524
rect 18211 24490 18253 24524
rect 18287 24490 18329 24524
rect 18363 24490 18405 24524
rect 18439 24500 18486 24524
rect 18520 24500 18556 24534
rect 18590 24500 18626 24534
rect 18660 24500 18696 24534
rect 18730 24500 18766 24534
rect 18800 24500 18836 24534
rect 18870 24500 18906 24534
rect 18940 24500 18976 24534
rect 19010 24500 19012 24534
rect 18439 24490 19012 24500
rect 18022 24465 19012 24490
rect 18022 24455 18486 24465
rect 18022 24421 18025 24455
rect 18059 24421 18101 24455
rect 18135 24421 18177 24455
rect 18211 24421 18253 24455
rect 18287 24421 18329 24455
rect 18363 24421 18405 24455
rect 18439 24431 18486 24455
rect 18520 24431 18556 24465
rect 18590 24431 18626 24465
rect 18660 24431 18696 24465
rect 18730 24431 18766 24465
rect 18800 24431 18836 24465
rect 18870 24431 18906 24465
rect 18940 24431 18976 24465
rect 19010 24431 19012 24465
rect 18439 24421 19012 24431
rect 18022 24396 19012 24421
rect 18022 24386 18486 24396
rect 18022 24352 18025 24386
rect 18059 24352 18101 24386
rect 18135 24352 18177 24386
rect 18211 24352 18253 24386
rect 18287 24352 18329 24386
rect 18363 24352 18405 24386
rect 18439 24362 18486 24386
rect 18520 24362 18556 24396
rect 18590 24362 18626 24396
rect 18660 24362 18696 24396
rect 18730 24362 18766 24396
rect 18800 24362 18836 24396
rect 18870 24362 18906 24396
rect 18940 24362 18976 24396
rect 19010 24362 19012 24396
rect 18439 24352 19012 24362
rect 18022 24327 19012 24352
rect 18022 24317 18486 24327
rect 18022 24283 18025 24317
rect 18059 24283 18101 24317
rect 18135 24283 18177 24317
rect 18211 24283 18253 24317
rect 18287 24283 18329 24317
rect 18363 24283 18405 24317
rect 18439 24293 18486 24317
rect 18520 24293 18556 24327
rect 18590 24293 18626 24327
rect 18660 24293 18696 24327
rect 18730 24293 18766 24327
rect 18800 24293 18836 24327
rect 18870 24293 18906 24327
rect 18940 24293 18976 24327
rect 19010 24293 19012 24327
rect 18439 24283 19012 24293
rect 18022 24258 19012 24283
rect 18022 24248 18486 24258
rect 18022 24214 18025 24248
rect 18059 24214 18101 24248
rect 18135 24214 18177 24248
rect 18211 24214 18253 24248
rect 18287 24214 18329 24248
rect 18363 24214 18405 24248
rect 18439 24224 18486 24248
rect 18520 24224 18556 24258
rect 18590 24224 18626 24258
rect 18660 24224 18696 24258
rect 18730 24224 18766 24258
rect 18800 24224 18836 24258
rect 18870 24224 18906 24258
rect 18940 24224 18976 24258
rect 19010 24224 19012 24258
rect 18439 24214 19012 24224
rect 18022 24189 19012 24214
rect 18022 24179 18486 24189
rect 18022 24145 18025 24179
rect 18059 24145 18101 24179
rect 18135 24145 18177 24179
rect 18211 24145 18253 24179
rect 18287 24145 18329 24179
rect 18363 24145 18405 24179
rect 18439 24155 18486 24179
rect 18520 24155 18556 24189
rect 18590 24155 18626 24189
rect 18660 24155 18696 24189
rect 18730 24155 18766 24189
rect 18800 24155 18836 24189
rect 18870 24155 18906 24189
rect 18940 24155 18976 24189
rect 19010 24155 19012 24189
rect 18439 24145 19012 24155
rect 18022 24120 19012 24145
rect 18022 24110 18486 24120
rect 18022 24076 18025 24110
rect 18059 24076 18101 24110
rect 18135 24076 18177 24110
rect 18211 24076 18253 24110
rect 18287 24076 18329 24110
rect 18363 24076 18405 24110
rect 18439 24086 18486 24110
rect 18520 24086 18556 24120
rect 18590 24086 18626 24120
rect 18660 24086 18696 24120
rect 18730 24086 18766 24120
rect 18800 24086 18836 24120
rect 18870 24086 18906 24120
rect 18940 24086 18976 24120
rect 19010 24086 19012 24120
rect 18439 24076 19012 24086
rect 18022 24051 19012 24076
rect 18022 24041 18486 24051
rect 18022 24007 18025 24041
rect 18059 24007 18101 24041
rect 18135 24007 18177 24041
rect 18211 24007 18253 24041
rect 18287 24007 18329 24041
rect 18363 24007 18405 24041
rect 18439 24017 18486 24041
rect 18520 24017 18556 24051
rect 18590 24017 18626 24051
rect 18660 24017 18696 24051
rect 18730 24017 18766 24051
rect 18800 24017 18836 24051
rect 18870 24017 18906 24051
rect 18940 24017 18976 24051
rect 19010 24017 19012 24051
rect 18439 24007 19012 24017
rect 18022 23982 19012 24007
rect 18022 23972 18486 23982
rect 18022 23938 18025 23972
rect 18059 23938 18101 23972
rect 18135 23938 18177 23972
rect 18211 23938 18253 23972
rect 18287 23938 18329 23972
rect 18363 23938 18405 23972
rect 18439 23948 18486 23972
rect 18520 23948 18556 23982
rect 18590 23948 18626 23982
rect 18660 23948 18696 23982
rect 18730 23948 18766 23982
rect 18800 23948 18836 23982
rect 18870 23948 18906 23982
rect 18940 23948 18976 23982
rect 19010 23948 19012 23982
rect 18439 23938 19012 23948
rect 18022 23913 19012 23938
rect 18022 23903 18486 23913
rect 18022 23869 18025 23903
rect 18059 23869 18101 23903
rect 18135 23869 18177 23903
rect 18211 23869 18253 23903
rect 18287 23869 18329 23903
rect 18363 23869 18405 23903
rect 18439 23879 18486 23903
rect 18520 23879 18556 23913
rect 18590 23879 18626 23913
rect 18660 23879 18696 23913
rect 18730 23879 18766 23913
rect 18800 23879 18836 23913
rect 18870 23879 18906 23913
rect 18940 23879 18976 23913
rect 19010 23879 19012 23913
rect 18439 23869 19012 23879
rect 18022 23844 19012 23869
rect 18022 23834 18486 23844
rect 280 23753 1741 23803
rect 280 23719 314 23753
rect 348 23719 384 23753
rect 418 23719 454 23753
rect 488 23719 524 23753
rect 558 23719 594 23753
rect 628 23719 664 23753
rect 698 23719 734 23753
rect 768 23719 804 23753
rect 838 23719 874 23753
rect 908 23719 944 23753
rect 978 23719 1014 23753
rect 1048 23719 1084 23753
rect 1118 23719 1154 23753
rect 1188 23719 1224 23753
rect 1258 23719 1294 23753
rect 1328 23719 1364 23753
rect 1398 23719 1434 23753
rect 1468 23719 1545 23753
rect 1579 23719 1613 23753
rect 1647 23719 1681 23753
rect 1715 23719 1741 23753
rect 280 23683 1741 23719
rect 280 23649 314 23683
rect 348 23649 384 23683
rect 418 23649 454 23683
rect 488 23649 524 23683
rect 558 23649 594 23683
rect 628 23649 664 23683
rect 698 23649 734 23683
rect 768 23649 804 23683
rect 838 23649 874 23683
rect 908 23649 944 23683
rect 978 23649 1014 23683
rect 1048 23649 1084 23683
rect 1118 23649 1154 23683
rect 1188 23649 1224 23683
rect 1258 23649 1294 23683
rect 1328 23649 1364 23683
rect 1398 23649 1434 23683
rect 1468 23650 1741 23683
rect 1468 23649 1545 23650
rect 280 23616 1545 23649
rect 1579 23616 1613 23650
rect 1647 23616 1681 23650
rect 1715 23616 1741 23650
rect 280 23613 1741 23616
rect 280 23579 314 23613
rect 348 23579 384 23613
rect 418 23579 454 23613
rect 488 23579 524 23613
rect 558 23579 594 23613
rect 628 23579 664 23613
rect 698 23579 734 23613
rect 768 23579 804 23613
rect 838 23579 874 23613
rect 908 23579 944 23613
rect 978 23579 1014 23613
rect 1048 23579 1084 23613
rect 1118 23579 1154 23613
rect 1188 23579 1224 23613
rect 1258 23579 1294 23613
rect 1328 23579 1364 23613
rect 1398 23579 1434 23613
rect 1468 23592 1741 23613
rect 18022 23800 18025 23834
rect 18059 23800 18101 23834
rect 18135 23800 18177 23834
rect 18211 23800 18253 23834
rect 18287 23800 18329 23834
rect 18363 23800 18405 23834
rect 18439 23810 18486 23834
rect 18520 23810 18556 23844
rect 18590 23810 18626 23844
rect 18660 23810 18696 23844
rect 18730 23810 18766 23844
rect 18800 23810 18836 23844
rect 18870 23810 18906 23844
rect 18940 23810 18976 23844
rect 19010 23810 19012 23844
rect 18439 23800 19012 23810
rect 18022 23775 19012 23800
rect 18022 23765 18486 23775
rect 18022 23731 18025 23765
rect 18059 23731 18101 23765
rect 18135 23731 18177 23765
rect 18211 23731 18253 23765
rect 18287 23731 18329 23765
rect 18363 23731 18405 23765
rect 18439 23741 18486 23765
rect 18520 23741 18556 23775
rect 18590 23741 18626 23775
rect 18660 23741 18696 23775
rect 18730 23741 18766 23775
rect 18800 23741 18836 23775
rect 18870 23741 18906 23775
rect 18940 23741 18976 23775
rect 19010 23741 19012 23775
rect 18439 23731 19012 23741
rect 18022 23706 19012 23731
rect 18022 23696 18486 23706
rect 18022 23662 18025 23696
rect 18059 23662 18101 23696
rect 18135 23662 18177 23696
rect 18211 23662 18253 23696
rect 18287 23662 18329 23696
rect 18363 23662 18405 23696
rect 18439 23672 18486 23696
rect 18520 23672 18556 23706
rect 18590 23672 18626 23706
rect 18660 23672 18696 23706
rect 18730 23672 18766 23706
rect 18800 23672 18836 23706
rect 18870 23672 18906 23706
rect 18940 23672 18976 23706
rect 19010 23672 19012 23706
rect 18439 23662 19012 23672
rect 18022 23637 19012 23662
rect 18022 23627 18486 23637
rect 18022 23593 18025 23627
rect 18059 23593 18101 23627
rect 18135 23593 18177 23627
rect 18211 23593 18253 23627
rect 18287 23593 18329 23627
rect 18363 23593 18405 23627
rect 18439 23603 18486 23627
rect 18520 23603 18556 23637
rect 18590 23603 18626 23637
rect 18660 23603 18696 23637
rect 18730 23603 18766 23637
rect 18800 23603 18836 23637
rect 18870 23603 18906 23637
rect 18940 23603 18976 23637
rect 19010 23603 19012 23637
rect 18439 23593 19012 23603
rect 1468 23579 1502 23592
rect 280 23543 1502 23579
rect 280 23509 314 23543
rect 348 23509 384 23543
rect 418 23509 454 23543
rect 488 23509 524 23543
rect 558 23509 594 23543
rect 628 23509 664 23543
rect 698 23509 734 23543
rect 768 23509 804 23543
rect 838 23509 874 23543
rect 908 23509 944 23543
rect 978 23509 1014 23543
rect 1048 23509 1084 23543
rect 1118 23509 1154 23543
rect 1188 23509 1224 23543
rect 1258 23509 1294 23543
rect 1328 23509 1364 23543
rect 1398 23509 1434 23543
rect 1468 23509 1502 23543
rect 280 23473 1502 23509
rect 18022 23568 19012 23593
rect 18022 23558 18486 23568
rect 18022 23524 18025 23558
rect 18059 23524 18101 23558
rect 18135 23524 18177 23558
rect 18211 23524 18253 23558
rect 18287 23524 18329 23558
rect 18363 23524 18405 23558
rect 18439 23534 18486 23558
rect 18520 23534 18556 23568
rect 18590 23534 18626 23568
rect 18660 23534 18696 23568
rect 18730 23534 18766 23568
rect 18800 23534 18836 23568
rect 18870 23534 18906 23568
rect 18940 23534 18976 23568
rect 19010 23534 19012 23568
rect 18439 23524 19012 23534
rect 18022 23500 19012 23524
rect 22823 30683 22827 30717
rect 22861 30683 22897 30717
rect 22931 30683 22967 30717
rect 23001 30683 23037 30717
rect 23071 30683 23107 30717
rect 23141 30683 23177 30717
rect 23211 30683 23247 30717
rect 23281 30683 23317 30717
rect 23351 30683 23387 30717
rect 23421 30683 23457 30717
rect 23491 30683 23527 30717
rect 23561 30683 23597 30717
rect 23631 30683 23635 30717
rect 22823 30649 23635 30683
rect 22823 30615 22827 30649
rect 22861 30615 22897 30649
rect 22931 30615 22967 30649
rect 23001 30615 23037 30649
rect 23071 30615 23107 30649
rect 23141 30615 23177 30649
rect 23211 30615 23247 30649
rect 23281 30615 23317 30649
rect 23351 30615 23387 30649
rect 23421 30615 23457 30649
rect 23491 30615 23527 30649
rect 23561 30615 23597 30649
rect 23631 30615 23635 30649
rect 22823 30581 23635 30615
rect 22823 30547 22827 30581
rect 22861 30547 22897 30581
rect 22931 30547 22967 30581
rect 23001 30547 23037 30581
rect 23071 30547 23107 30581
rect 23141 30547 23177 30581
rect 23211 30547 23247 30581
rect 23281 30547 23317 30581
rect 23351 30547 23387 30581
rect 23421 30547 23457 30581
rect 23491 30547 23527 30581
rect 23561 30547 23597 30581
rect 23631 30547 23635 30581
rect 22823 30513 23635 30547
rect 22823 30479 22827 30513
rect 22861 30479 22897 30513
rect 22931 30479 22967 30513
rect 23001 30479 23037 30513
rect 23071 30479 23107 30513
rect 23141 30479 23177 30513
rect 23211 30479 23247 30513
rect 23281 30479 23317 30513
rect 23351 30479 23387 30513
rect 23421 30479 23457 30513
rect 23491 30479 23527 30513
rect 23561 30479 23597 30513
rect 23631 30479 23635 30513
rect 22823 30445 23635 30479
rect 22823 30411 22827 30445
rect 22861 30411 22897 30445
rect 22931 30411 22967 30445
rect 23001 30411 23037 30445
rect 23071 30411 23107 30445
rect 23141 30411 23177 30445
rect 23211 30411 23247 30445
rect 23281 30411 23317 30445
rect 23351 30411 23387 30445
rect 23421 30411 23457 30445
rect 23491 30411 23527 30445
rect 23561 30411 23597 30445
rect 23631 30411 23635 30445
rect 22823 30377 23635 30411
rect 22823 30343 22827 30377
rect 22861 30343 22897 30377
rect 22931 30343 22967 30377
rect 23001 30343 23037 30377
rect 23071 30343 23107 30377
rect 23141 30343 23177 30377
rect 23211 30343 23247 30377
rect 23281 30343 23317 30377
rect 23351 30343 23387 30377
rect 23421 30343 23457 30377
rect 23491 30343 23527 30377
rect 23561 30343 23597 30377
rect 23631 30343 23635 30377
rect 22823 30309 23635 30343
rect 22823 30275 22827 30309
rect 22861 30275 22897 30309
rect 22931 30275 22967 30309
rect 23001 30275 23037 30309
rect 23071 30275 23107 30309
rect 23141 30275 23177 30309
rect 23211 30275 23247 30309
rect 23281 30275 23317 30309
rect 23351 30275 23387 30309
rect 23421 30275 23457 30309
rect 23491 30275 23527 30309
rect 23561 30275 23597 30309
rect 23631 30275 23635 30309
rect 22823 30241 23635 30275
rect 22823 30207 22827 30241
rect 22861 30207 22897 30241
rect 22931 30207 22967 30241
rect 23001 30207 23037 30241
rect 23071 30207 23107 30241
rect 23141 30207 23177 30241
rect 23211 30207 23247 30241
rect 23281 30207 23317 30241
rect 23351 30207 23387 30241
rect 23421 30207 23457 30241
rect 23491 30207 23527 30241
rect 23561 30207 23597 30241
rect 23631 30207 23635 30241
rect 22823 30173 23635 30207
rect 22823 30139 22827 30173
rect 22861 30139 22897 30173
rect 22931 30139 22967 30173
rect 23001 30139 23037 30173
rect 23071 30139 23107 30173
rect 23141 30139 23177 30173
rect 23211 30139 23247 30173
rect 23281 30139 23317 30173
rect 23351 30139 23387 30173
rect 23421 30139 23457 30173
rect 23491 30139 23527 30173
rect 23561 30139 23597 30173
rect 23631 30139 23635 30173
rect 22823 30105 23635 30139
rect 22823 30071 22827 30105
rect 22861 30071 22897 30105
rect 22931 30071 22967 30105
rect 23001 30071 23037 30105
rect 23071 30071 23107 30105
rect 23141 30071 23177 30105
rect 23211 30071 23247 30105
rect 23281 30071 23317 30105
rect 23351 30071 23387 30105
rect 23421 30071 23457 30105
rect 23491 30071 23527 30105
rect 23561 30071 23597 30105
rect 23631 30071 23635 30105
rect 22823 30037 23635 30071
rect 22823 30003 22827 30037
rect 22861 30003 22897 30037
rect 22931 30003 22967 30037
rect 23001 30003 23037 30037
rect 23071 30003 23107 30037
rect 23141 30003 23177 30037
rect 23211 30003 23247 30037
rect 23281 30003 23317 30037
rect 23351 30003 23387 30037
rect 23421 30003 23457 30037
rect 23491 30003 23527 30037
rect 23561 30003 23597 30037
rect 23631 30003 23635 30037
rect 22823 29969 23635 30003
rect 22823 29935 22827 29969
rect 22861 29935 22897 29969
rect 22931 29935 22967 29969
rect 23001 29935 23037 29969
rect 23071 29935 23107 29969
rect 23141 29935 23177 29969
rect 23211 29935 23247 29969
rect 23281 29935 23317 29969
rect 23351 29935 23387 29969
rect 23421 29935 23457 29969
rect 23491 29935 23527 29969
rect 23561 29935 23597 29969
rect 23631 29935 23635 29969
rect 22823 29901 23635 29935
rect 22823 29867 22827 29901
rect 22861 29867 22897 29901
rect 22931 29867 22967 29901
rect 23001 29867 23037 29901
rect 23071 29867 23107 29901
rect 23141 29867 23177 29901
rect 23211 29867 23247 29901
rect 23281 29867 23317 29901
rect 23351 29867 23387 29901
rect 23421 29867 23457 29901
rect 23491 29867 23527 29901
rect 23561 29867 23597 29901
rect 23631 29867 23635 29901
rect 22823 29833 23635 29867
rect 22823 29799 22827 29833
rect 22861 29799 22897 29833
rect 22931 29799 22967 29833
rect 23001 29799 23037 29833
rect 23071 29799 23107 29833
rect 23141 29799 23177 29833
rect 23211 29799 23247 29833
rect 23281 29799 23317 29833
rect 23351 29799 23387 29833
rect 23421 29799 23457 29833
rect 23491 29799 23527 29833
rect 23561 29799 23597 29833
rect 23631 29799 23635 29833
rect 22823 29765 23635 29799
rect 22823 29731 22827 29765
rect 22861 29731 22897 29765
rect 22931 29731 22967 29765
rect 23001 29731 23037 29765
rect 23071 29731 23107 29765
rect 23141 29731 23177 29765
rect 23211 29731 23247 29765
rect 23281 29731 23317 29765
rect 23351 29731 23387 29765
rect 23421 29731 23457 29765
rect 23491 29731 23527 29765
rect 23561 29731 23597 29765
rect 23631 29731 23635 29765
rect 22823 29697 23635 29731
rect 22823 29663 22827 29697
rect 22861 29663 22897 29697
rect 22931 29663 22967 29697
rect 23001 29663 23037 29697
rect 23071 29663 23107 29697
rect 23141 29663 23177 29697
rect 23211 29663 23247 29697
rect 23281 29663 23317 29697
rect 23351 29663 23387 29697
rect 23421 29663 23457 29697
rect 23491 29663 23527 29697
rect 23561 29663 23597 29697
rect 23631 29663 23635 29697
rect 22823 29629 23635 29663
rect 22823 29595 22827 29629
rect 22861 29595 22897 29629
rect 22931 29595 22967 29629
rect 23001 29595 23037 29629
rect 23071 29595 23107 29629
rect 23141 29595 23177 29629
rect 23211 29595 23247 29629
rect 23281 29595 23317 29629
rect 23351 29595 23387 29629
rect 23421 29595 23457 29629
rect 23491 29595 23527 29629
rect 23561 29595 23597 29629
rect 23631 29595 23635 29629
rect 22823 29561 23635 29595
rect 22823 29527 22827 29561
rect 22861 29527 22897 29561
rect 22931 29527 22967 29561
rect 23001 29527 23037 29561
rect 23071 29527 23107 29561
rect 23141 29527 23177 29561
rect 23211 29527 23247 29561
rect 23281 29527 23317 29561
rect 23351 29527 23387 29561
rect 23421 29527 23457 29561
rect 23491 29527 23527 29561
rect 23561 29527 23597 29561
rect 23631 29527 23635 29561
rect 22823 29493 23635 29527
rect 22823 29459 22827 29493
rect 22861 29459 22897 29493
rect 22931 29459 22967 29493
rect 23001 29459 23037 29493
rect 23071 29459 23107 29493
rect 23141 29459 23177 29493
rect 23211 29459 23247 29493
rect 23281 29459 23317 29493
rect 23351 29459 23387 29493
rect 23421 29459 23457 29493
rect 23491 29459 23527 29493
rect 23561 29459 23597 29493
rect 23631 29459 23635 29493
rect 22823 29425 23635 29459
rect 22823 29391 22827 29425
rect 22861 29391 22897 29425
rect 22931 29391 22967 29425
rect 23001 29391 23037 29425
rect 23071 29391 23107 29425
rect 23141 29391 23177 29425
rect 23211 29391 23247 29425
rect 23281 29391 23317 29425
rect 23351 29391 23387 29425
rect 23421 29391 23457 29425
rect 23491 29391 23527 29425
rect 23561 29391 23597 29425
rect 23631 29391 23635 29425
rect 22823 29357 23635 29391
rect 22823 29323 22827 29357
rect 22861 29323 22897 29357
rect 22931 29323 22967 29357
rect 23001 29323 23037 29357
rect 23071 29323 23107 29357
rect 23141 29323 23177 29357
rect 23211 29323 23247 29357
rect 23281 29323 23317 29357
rect 23351 29323 23387 29357
rect 23421 29323 23457 29357
rect 23491 29323 23527 29357
rect 23561 29323 23597 29357
rect 23631 29323 23635 29357
rect 22823 29289 23635 29323
rect 22823 29255 22827 29289
rect 22861 29255 22897 29289
rect 22931 29255 22967 29289
rect 23001 29255 23037 29289
rect 23071 29255 23107 29289
rect 23141 29255 23177 29289
rect 23211 29255 23247 29289
rect 23281 29255 23317 29289
rect 23351 29255 23387 29289
rect 23421 29255 23457 29289
rect 23491 29255 23527 29289
rect 23561 29255 23597 29289
rect 23631 29255 23635 29289
rect 22823 29221 23635 29255
rect 22823 29187 22827 29221
rect 22861 29187 22897 29221
rect 22931 29187 22967 29221
rect 23001 29187 23037 29221
rect 23071 29187 23107 29221
rect 23141 29187 23177 29221
rect 23211 29187 23247 29221
rect 23281 29187 23317 29221
rect 23351 29187 23387 29221
rect 23421 29187 23457 29221
rect 23491 29187 23527 29221
rect 23561 29187 23597 29221
rect 23631 29187 23635 29221
rect 22823 29153 23635 29187
rect 22823 29119 22827 29153
rect 22861 29119 22897 29153
rect 22931 29119 22967 29153
rect 23001 29119 23037 29153
rect 23071 29119 23107 29153
rect 23141 29119 23177 29153
rect 23211 29119 23247 29153
rect 23281 29119 23317 29153
rect 23351 29119 23387 29153
rect 23421 29119 23457 29153
rect 23491 29119 23527 29153
rect 23561 29119 23597 29153
rect 23631 29119 23635 29153
rect 22823 29085 23635 29119
rect 22823 29051 22827 29085
rect 22861 29051 22897 29085
rect 22931 29051 22967 29085
rect 23001 29051 23037 29085
rect 23071 29051 23107 29085
rect 23141 29051 23177 29085
rect 23211 29051 23247 29085
rect 23281 29051 23317 29085
rect 23351 29051 23387 29085
rect 23421 29051 23457 29085
rect 23491 29051 23527 29085
rect 23561 29051 23597 29085
rect 23631 29051 23635 29085
rect 22823 29017 23635 29051
rect 22823 28983 22827 29017
rect 22861 28983 22897 29017
rect 22931 28983 22967 29017
rect 23001 28983 23037 29017
rect 23071 28983 23107 29017
rect 23141 28983 23177 29017
rect 23211 28983 23247 29017
rect 23281 28983 23317 29017
rect 23351 28983 23387 29017
rect 23421 28983 23457 29017
rect 23491 28983 23527 29017
rect 23561 28983 23597 29017
rect 23631 28983 23635 29017
rect 22823 28949 23635 28983
rect 22823 28915 22827 28949
rect 22861 28915 22897 28949
rect 22931 28915 22967 28949
rect 23001 28915 23037 28949
rect 23071 28915 23107 28949
rect 23141 28915 23177 28949
rect 23211 28915 23247 28949
rect 23281 28915 23317 28949
rect 23351 28915 23387 28949
rect 23421 28915 23457 28949
rect 23491 28915 23527 28949
rect 23561 28915 23597 28949
rect 23631 28915 23635 28949
rect 22823 28881 23635 28915
rect 22823 28847 22827 28881
rect 22861 28847 22897 28881
rect 22931 28847 22967 28881
rect 23001 28847 23037 28881
rect 23071 28847 23107 28881
rect 23141 28847 23177 28881
rect 23211 28847 23247 28881
rect 23281 28847 23317 28881
rect 23351 28847 23387 28881
rect 23421 28847 23457 28881
rect 23491 28847 23527 28881
rect 23561 28847 23597 28881
rect 23631 28847 23635 28881
rect 22823 28813 23635 28847
rect 22823 28779 22827 28813
rect 22861 28779 22897 28813
rect 22931 28779 22967 28813
rect 23001 28779 23037 28813
rect 23071 28779 23107 28813
rect 23141 28779 23177 28813
rect 23211 28779 23247 28813
rect 23281 28779 23317 28813
rect 23351 28779 23387 28813
rect 23421 28779 23457 28813
rect 23491 28779 23527 28813
rect 23561 28779 23597 28813
rect 23631 28779 23635 28813
rect 22823 28745 23635 28779
rect 22823 28711 22827 28745
rect 22861 28711 22897 28745
rect 22931 28711 22967 28745
rect 23001 28711 23037 28745
rect 23071 28711 23107 28745
rect 23141 28711 23177 28745
rect 23211 28711 23247 28745
rect 23281 28711 23317 28745
rect 23351 28711 23387 28745
rect 23421 28711 23457 28745
rect 23491 28711 23527 28745
rect 23561 28711 23597 28745
rect 23631 28711 23635 28745
rect 22823 28677 23635 28711
rect 22823 28643 22827 28677
rect 22861 28643 22897 28677
rect 22931 28643 22967 28677
rect 23001 28643 23037 28677
rect 23071 28643 23107 28677
rect 23141 28643 23177 28677
rect 23211 28643 23247 28677
rect 23281 28643 23317 28677
rect 23351 28643 23387 28677
rect 23421 28643 23457 28677
rect 23491 28643 23527 28677
rect 23561 28643 23597 28677
rect 23631 28643 23635 28677
rect 22823 28609 23635 28643
rect 22823 28575 22827 28609
rect 22861 28575 22897 28609
rect 22931 28575 22967 28609
rect 23001 28575 23037 28609
rect 23071 28575 23107 28609
rect 23141 28575 23177 28609
rect 23211 28575 23247 28609
rect 23281 28575 23317 28609
rect 23351 28575 23387 28609
rect 23421 28575 23457 28609
rect 23491 28575 23527 28609
rect 23561 28575 23597 28609
rect 23631 28575 23635 28609
rect 22823 28541 23635 28575
rect 22823 28507 22827 28541
rect 22861 28507 22897 28541
rect 22931 28507 22967 28541
rect 23001 28507 23037 28541
rect 23071 28507 23107 28541
rect 23141 28507 23177 28541
rect 23211 28507 23247 28541
rect 23281 28507 23317 28541
rect 23351 28507 23387 28541
rect 23421 28507 23457 28541
rect 23491 28507 23527 28541
rect 23561 28507 23597 28541
rect 23631 28507 23635 28541
rect 22823 28473 23635 28507
rect 22823 28439 22827 28473
rect 22861 28439 22897 28473
rect 22931 28439 22967 28473
rect 23001 28439 23037 28473
rect 23071 28439 23107 28473
rect 23141 28439 23177 28473
rect 23211 28439 23247 28473
rect 23281 28439 23317 28473
rect 23351 28439 23387 28473
rect 23421 28439 23457 28473
rect 23491 28439 23527 28473
rect 23561 28439 23597 28473
rect 23631 28439 23635 28473
rect 22823 28405 23635 28439
rect 22823 28371 22827 28405
rect 22861 28371 22897 28405
rect 22931 28371 22967 28405
rect 23001 28371 23037 28405
rect 23071 28371 23107 28405
rect 23141 28371 23177 28405
rect 23211 28371 23247 28405
rect 23281 28371 23317 28405
rect 23351 28371 23387 28405
rect 23421 28371 23457 28405
rect 23491 28371 23527 28405
rect 23561 28371 23597 28405
rect 23631 28371 23635 28405
rect 22823 28337 23635 28371
rect 22823 28303 22827 28337
rect 22861 28303 22897 28337
rect 22931 28303 22967 28337
rect 23001 28303 23037 28337
rect 23071 28303 23107 28337
rect 23141 28303 23177 28337
rect 23211 28303 23247 28337
rect 23281 28303 23317 28337
rect 23351 28303 23387 28337
rect 23421 28303 23457 28337
rect 23491 28303 23527 28337
rect 23561 28303 23597 28337
rect 23631 28303 23635 28337
rect 22823 28269 23635 28303
rect 22823 28235 22827 28269
rect 22861 28235 22897 28269
rect 22931 28235 22967 28269
rect 23001 28235 23037 28269
rect 23071 28235 23107 28269
rect 23141 28235 23177 28269
rect 23211 28235 23247 28269
rect 23281 28235 23317 28269
rect 23351 28235 23387 28269
rect 23421 28235 23457 28269
rect 23491 28235 23527 28269
rect 23561 28235 23597 28269
rect 23631 28235 23635 28269
rect 22823 28201 23635 28235
rect 22823 28167 22827 28201
rect 22861 28167 22897 28201
rect 22931 28167 22967 28201
rect 23001 28167 23037 28201
rect 23071 28167 23107 28201
rect 23141 28167 23177 28201
rect 23211 28167 23247 28201
rect 23281 28167 23317 28201
rect 23351 28167 23387 28201
rect 23421 28167 23457 28201
rect 23491 28167 23527 28201
rect 23561 28167 23597 28201
rect 23631 28167 23635 28201
rect 22823 28133 23635 28167
rect 22823 28099 22827 28133
rect 22861 28099 22897 28133
rect 22931 28099 22967 28133
rect 23001 28099 23037 28133
rect 23071 28099 23107 28133
rect 23141 28099 23177 28133
rect 23211 28099 23247 28133
rect 23281 28099 23317 28133
rect 23351 28099 23387 28133
rect 23421 28099 23457 28133
rect 23491 28099 23527 28133
rect 23561 28099 23597 28133
rect 23631 28099 23635 28133
rect 22823 28065 23635 28099
rect 22823 28031 22827 28065
rect 22861 28031 22897 28065
rect 22931 28031 22967 28065
rect 23001 28031 23037 28065
rect 23071 28031 23107 28065
rect 23141 28031 23177 28065
rect 23211 28031 23247 28065
rect 23281 28031 23317 28065
rect 23351 28031 23387 28065
rect 23421 28031 23457 28065
rect 23491 28031 23527 28065
rect 23561 28031 23597 28065
rect 23631 28031 23635 28065
rect 22823 27997 23635 28031
rect 22823 27963 22827 27997
rect 22861 27963 22897 27997
rect 22931 27963 22967 27997
rect 23001 27963 23037 27997
rect 23071 27963 23107 27997
rect 23141 27963 23177 27997
rect 23211 27963 23247 27997
rect 23281 27963 23317 27997
rect 23351 27963 23387 27997
rect 23421 27963 23457 27997
rect 23491 27963 23527 27997
rect 23561 27963 23597 27997
rect 23631 27963 23635 27997
rect 22823 27929 23635 27963
rect 22823 27895 22827 27929
rect 22861 27895 22897 27929
rect 22931 27895 22967 27929
rect 23001 27895 23037 27929
rect 23071 27895 23107 27929
rect 23141 27895 23177 27929
rect 23211 27895 23247 27929
rect 23281 27895 23317 27929
rect 23351 27895 23387 27929
rect 23421 27895 23457 27929
rect 23491 27895 23527 27929
rect 23561 27895 23597 27929
rect 23631 27895 23635 27929
rect 22823 27861 23635 27895
rect 22823 27827 22827 27861
rect 22861 27827 22897 27861
rect 22931 27827 22967 27861
rect 23001 27827 23037 27861
rect 23071 27827 23107 27861
rect 23141 27827 23177 27861
rect 23211 27827 23247 27861
rect 23281 27827 23317 27861
rect 23351 27827 23387 27861
rect 23421 27827 23457 27861
rect 23491 27827 23527 27861
rect 23561 27827 23597 27861
rect 23631 27827 23635 27861
rect 22823 27793 23635 27827
rect 22823 27759 22827 27793
rect 22861 27759 22897 27793
rect 22931 27759 22967 27793
rect 23001 27759 23037 27793
rect 23071 27759 23107 27793
rect 23141 27759 23177 27793
rect 23211 27759 23247 27793
rect 23281 27759 23317 27793
rect 23351 27759 23387 27793
rect 23421 27759 23457 27793
rect 23491 27759 23527 27793
rect 23561 27759 23597 27793
rect 23631 27759 23635 27793
rect 22823 27725 23635 27759
rect 22823 27691 22827 27725
rect 22861 27691 22897 27725
rect 22931 27691 22967 27725
rect 23001 27691 23037 27725
rect 23071 27691 23107 27725
rect 23141 27691 23177 27725
rect 23211 27691 23247 27725
rect 23281 27691 23317 27725
rect 23351 27691 23387 27725
rect 23421 27691 23457 27725
rect 23491 27691 23527 27725
rect 23561 27691 23597 27725
rect 23631 27691 23635 27725
rect 22823 27657 23635 27691
rect 22823 27623 22827 27657
rect 22861 27623 22897 27657
rect 22931 27623 22967 27657
rect 23001 27623 23037 27657
rect 23071 27623 23107 27657
rect 23141 27623 23177 27657
rect 23211 27623 23247 27657
rect 23281 27623 23317 27657
rect 23351 27623 23387 27657
rect 23421 27623 23457 27657
rect 23491 27623 23527 27657
rect 23561 27623 23597 27657
rect 23631 27623 23635 27657
rect 22823 27589 23635 27623
rect 22823 27555 22827 27589
rect 22861 27555 22897 27589
rect 22931 27555 22967 27589
rect 23001 27555 23037 27589
rect 23071 27555 23107 27589
rect 23141 27555 23177 27589
rect 23211 27555 23247 27589
rect 23281 27555 23317 27589
rect 23351 27555 23387 27589
rect 23421 27555 23457 27589
rect 23491 27555 23527 27589
rect 23561 27555 23597 27589
rect 23631 27555 23635 27589
rect 22823 27521 23635 27555
rect 22823 27487 22827 27521
rect 22861 27487 22897 27521
rect 22931 27487 22967 27521
rect 23001 27487 23037 27521
rect 23071 27487 23107 27521
rect 23141 27487 23177 27521
rect 23211 27487 23247 27521
rect 23281 27487 23317 27521
rect 23351 27487 23387 27521
rect 23421 27487 23457 27521
rect 23491 27487 23527 27521
rect 23561 27487 23597 27521
rect 23631 27487 23635 27521
rect 22823 27453 23635 27487
rect 22823 27419 22827 27453
rect 22861 27419 22897 27453
rect 22931 27419 22967 27453
rect 23001 27419 23037 27453
rect 23071 27419 23107 27453
rect 23141 27419 23177 27453
rect 23211 27419 23247 27453
rect 23281 27419 23317 27453
rect 23351 27419 23387 27453
rect 23421 27419 23457 27453
rect 23491 27419 23527 27453
rect 23561 27419 23597 27453
rect 23631 27419 23635 27453
rect 22823 27385 23635 27419
rect 22823 27351 22827 27385
rect 22861 27351 22897 27385
rect 22931 27351 22967 27385
rect 23001 27351 23037 27385
rect 23071 27351 23107 27385
rect 23141 27351 23177 27385
rect 23211 27351 23247 27385
rect 23281 27351 23317 27385
rect 23351 27351 23387 27385
rect 23421 27351 23457 27385
rect 23491 27351 23527 27385
rect 23561 27351 23597 27385
rect 23631 27351 23635 27385
rect 22823 27317 23635 27351
rect 22823 27283 22827 27317
rect 22861 27283 22897 27317
rect 22931 27283 22967 27317
rect 23001 27283 23037 27317
rect 23071 27283 23107 27317
rect 23141 27283 23177 27317
rect 23211 27283 23247 27317
rect 23281 27283 23317 27317
rect 23351 27283 23387 27317
rect 23421 27283 23457 27317
rect 23491 27283 23527 27317
rect 23561 27283 23597 27317
rect 23631 27283 23635 27317
rect 22823 27249 23635 27283
rect 22823 27215 22827 27249
rect 22861 27215 22897 27249
rect 22931 27215 22967 27249
rect 23001 27215 23037 27249
rect 23071 27215 23107 27249
rect 23141 27215 23177 27249
rect 23211 27215 23247 27249
rect 23281 27215 23317 27249
rect 23351 27215 23387 27249
rect 23421 27215 23457 27249
rect 23491 27215 23527 27249
rect 23561 27215 23597 27249
rect 23631 27215 23635 27249
rect 22823 27181 23635 27215
rect 22823 27147 22827 27181
rect 22861 27147 22897 27181
rect 22931 27147 22967 27181
rect 23001 27147 23037 27181
rect 23071 27147 23107 27181
rect 23141 27147 23177 27181
rect 23211 27147 23247 27181
rect 23281 27147 23317 27181
rect 23351 27147 23387 27181
rect 23421 27147 23457 27181
rect 23491 27147 23527 27181
rect 23561 27147 23597 27181
rect 23631 27147 23635 27181
rect 22823 27113 23635 27147
rect 22823 27079 22827 27113
rect 22861 27079 22897 27113
rect 22931 27079 22967 27113
rect 23001 27079 23037 27113
rect 23071 27079 23107 27113
rect 23141 27079 23177 27113
rect 23211 27079 23247 27113
rect 23281 27079 23317 27113
rect 23351 27079 23387 27113
rect 23421 27079 23457 27113
rect 23491 27079 23527 27113
rect 23561 27079 23597 27113
rect 23631 27079 23635 27113
rect 22823 27045 23635 27079
rect 22823 27011 22827 27045
rect 22861 27011 22897 27045
rect 22931 27011 22967 27045
rect 23001 27011 23037 27045
rect 23071 27011 23107 27045
rect 23141 27011 23177 27045
rect 23211 27011 23247 27045
rect 23281 27011 23317 27045
rect 23351 27011 23387 27045
rect 23421 27011 23457 27045
rect 23491 27011 23527 27045
rect 23561 27011 23597 27045
rect 23631 27011 23635 27045
rect 22823 26977 23635 27011
rect 22823 26943 22827 26977
rect 22861 26943 22897 26977
rect 22931 26943 22967 26977
rect 23001 26943 23037 26977
rect 23071 26943 23107 26977
rect 23141 26943 23177 26977
rect 23211 26943 23247 26977
rect 23281 26943 23317 26977
rect 23351 26943 23387 26977
rect 23421 26943 23457 26977
rect 23491 26943 23527 26977
rect 23561 26943 23597 26977
rect 23631 26943 23635 26977
rect 22823 26909 23635 26943
rect 22823 26875 22827 26909
rect 22861 26875 22897 26909
rect 22931 26875 22967 26909
rect 23001 26875 23037 26909
rect 23071 26875 23107 26909
rect 23141 26875 23177 26909
rect 23211 26875 23247 26909
rect 23281 26875 23317 26909
rect 23351 26875 23387 26909
rect 23421 26875 23457 26909
rect 23491 26875 23527 26909
rect 23561 26875 23597 26909
rect 23631 26875 23635 26909
rect 22823 26841 23635 26875
rect 22823 26807 22827 26841
rect 22861 26807 22897 26841
rect 22931 26807 22967 26841
rect 23001 26807 23037 26841
rect 23071 26807 23107 26841
rect 23141 26807 23177 26841
rect 23211 26807 23247 26841
rect 23281 26807 23317 26841
rect 23351 26807 23387 26841
rect 23421 26807 23457 26841
rect 23491 26807 23527 26841
rect 23561 26807 23597 26841
rect 23631 26807 23635 26841
rect 22823 26773 23635 26807
rect 22823 26739 22827 26773
rect 22861 26739 22897 26773
rect 22931 26739 22967 26773
rect 23001 26739 23037 26773
rect 23071 26739 23107 26773
rect 23141 26739 23177 26773
rect 23211 26739 23247 26773
rect 23281 26739 23317 26773
rect 23351 26739 23387 26773
rect 23421 26739 23457 26773
rect 23491 26739 23527 26773
rect 23561 26739 23597 26773
rect 23631 26739 23635 26773
rect 22823 26705 23635 26739
rect 22823 26671 22827 26705
rect 22861 26671 22897 26705
rect 22931 26671 22967 26705
rect 23001 26671 23037 26705
rect 23071 26671 23107 26705
rect 23141 26671 23177 26705
rect 23211 26671 23247 26705
rect 23281 26671 23317 26705
rect 23351 26671 23387 26705
rect 23421 26671 23457 26705
rect 23491 26671 23527 26705
rect 23561 26671 23597 26705
rect 23631 26671 23635 26705
rect 22823 26637 23635 26671
rect 22823 26603 22827 26637
rect 22861 26603 22897 26637
rect 22931 26603 22967 26637
rect 23001 26603 23037 26637
rect 23071 26603 23107 26637
rect 23141 26603 23177 26637
rect 23211 26603 23247 26637
rect 23281 26603 23317 26637
rect 23351 26603 23387 26637
rect 23421 26603 23457 26637
rect 23491 26603 23527 26637
rect 23561 26603 23597 26637
rect 23631 26603 23635 26637
rect 22823 26569 23635 26603
rect 22823 26535 22827 26569
rect 22861 26535 22897 26569
rect 22931 26535 22967 26569
rect 23001 26535 23037 26569
rect 23071 26535 23107 26569
rect 23141 26535 23177 26569
rect 23211 26535 23247 26569
rect 23281 26535 23317 26569
rect 23351 26535 23387 26569
rect 23421 26535 23457 26569
rect 23491 26535 23527 26569
rect 23561 26535 23597 26569
rect 23631 26535 23635 26569
rect 22823 26501 23635 26535
rect 22823 26467 22827 26501
rect 22861 26467 22897 26501
rect 22931 26467 22967 26501
rect 23001 26467 23037 26501
rect 23071 26467 23107 26501
rect 23141 26467 23177 26501
rect 23211 26467 23247 26501
rect 23281 26467 23317 26501
rect 23351 26467 23387 26501
rect 23421 26467 23457 26501
rect 23491 26467 23527 26501
rect 23561 26467 23597 26501
rect 23631 26467 23635 26501
rect 22823 26433 23635 26467
rect 22823 26399 22827 26433
rect 22861 26399 22897 26433
rect 22931 26399 22967 26433
rect 23001 26399 23037 26433
rect 23071 26399 23107 26433
rect 23141 26399 23177 26433
rect 23211 26399 23247 26433
rect 23281 26399 23317 26433
rect 23351 26399 23387 26433
rect 23421 26399 23457 26433
rect 23491 26399 23527 26433
rect 23561 26399 23597 26433
rect 23631 26399 23635 26433
rect 22823 26365 23635 26399
rect 22823 26331 22827 26365
rect 22861 26331 22897 26365
rect 22931 26331 22967 26365
rect 23001 26331 23037 26365
rect 23071 26331 23107 26365
rect 23141 26331 23177 26365
rect 23211 26331 23247 26365
rect 23281 26331 23317 26365
rect 23351 26331 23387 26365
rect 23421 26331 23457 26365
rect 23491 26331 23527 26365
rect 23561 26331 23597 26365
rect 23631 26331 23635 26365
rect 22823 26297 23635 26331
rect 22823 26263 22827 26297
rect 22861 26263 22897 26297
rect 22931 26263 22967 26297
rect 23001 26263 23037 26297
rect 23071 26263 23107 26297
rect 23141 26263 23177 26297
rect 23211 26263 23247 26297
rect 23281 26263 23317 26297
rect 23351 26263 23387 26297
rect 23421 26263 23457 26297
rect 23491 26263 23527 26297
rect 23561 26263 23597 26297
rect 23631 26263 23635 26297
rect 22823 26229 23635 26263
rect 22823 26195 22827 26229
rect 22861 26195 22897 26229
rect 22931 26195 22967 26229
rect 23001 26195 23037 26229
rect 23071 26195 23107 26229
rect 23141 26195 23177 26229
rect 23211 26195 23247 26229
rect 23281 26195 23317 26229
rect 23351 26195 23387 26229
rect 23421 26195 23457 26229
rect 23491 26195 23527 26229
rect 23561 26195 23597 26229
rect 23631 26195 23635 26229
rect 22823 26161 23635 26195
rect 22823 26127 22827 26161
rect 22861 26127 22897 26161
rect 22931 26127 22967 26161
rect 23001 26127 23037 26161
rect 23071 26127 23107 26161
rect 23141 26127 23177 26161
rect 23211 26127 23247 26161
rect 23281 26127 23317 26161
rect 23351 26127 23387 26161
rect 23421 26127 23457 26161
rect 23491 26127 23527 26161
rect 23561 26127 23597 26161
rect 23631 26127 23635 26161
rect 22823 26093 23635 26127
rect 22823 26059 22827 26093
rect 22861 26059 22897 26093
rect 22931 26059 22967 26093
rect 23001 26059 23037 26093
rect 23071 26059 23107 26093
rect 23141 26059 23177 26093
rect 23211 26059 23247 26093
rect 23281 26059 23317 26093
rect 23351 26059 23387 26093
rect 23421 26059 23457 26093
rect 23491 26059 23527 26093
rect 23561 26059 23597 26093
rect 23631 26059 23635 26093
rect 22823 26025 23635 26059
rect 22823 25991 22827 26025
rect 22861 25991 22897 26025
rect 22931 25991 22967 26025
rect 23001 25991 23037 26025
rect 23071 25991 23107 26025
rect 23141 25991 23177 26025
rect 23211 25991 23247 26025
rect 23281 25991 23317 26025
rect 23351 25991 23387 26025
rect 23421 25991 23457 26025
rect 23491 25991 23527 26025
rect 23561 25991 23597 26025
rect 23631 25991 23635 26025
rect 22823 25957 23635 25991
rect 22823 25923 22827 25957
rect 22861 25923 22897 25957
rect 22931 25923 22967 25957
rect 23001 25923 23037 25957
rect 23071 25923 23107 25957
rect 23141 25923 23177 25957
rect 23211 25923 23247 25957
rect 23281 25923 23317 25957
rect 23351 25923 23387 25957
rect 23421 25923 23457 25957
rect 23491 25923 23527 25957
rect 23561 25923 23597 25957
rect 23631 25923 23635 25957
rect 22823 25889 23635 25923
rect 22823 25855 22827 25889
rect 22861 25855 22897 25889
rect 22931 25855 22967 25889
rect 23001 25855 23037 25889
rect 23071 25855 23107 25889
rect 23141 25855 23177 25889
rect 23211 25855 23247 25889
rect 23281 25855 23317 25889
rect 23351 25855 23387 25889
rect 23421 25855 23457 25889
rect 23491 25855 23527 25889
rect 23561 25855 23597 25889
rect 23631 25855 23635 25889
rect 22823 25821 23635 25855
rect 22823 25787 22827 25821
rect 22861 25787 22897 25821
rect 22931 25787 22967 25821
rect 23001 25787 23037 25821
rect 23071 25787 23107 25821
rect 23141 25787 23177 25821
rect 23211 25787 23247 25821
rect 23281 25787 23317 25821
rect 23351 25787 23387 25821
rect 23421 25787 23457 25821
rect 23491 25787 23527 25821
rect 23561 25787 23597 25821
rect 23631 25787 23635 25821
rect 22823 25753 23635 25787
rect 22823 25719 22827 25753
rect 22861 25719 22897 25753
rect 22931 25719 22967 25753
rect 23001 25719 23037 25753
rect 23071 25719 23107 25753
rect 23141 25719 23177 25753
rect 23211 25719 23247 25753
rect 23281 25719 23317 25753
rect 23351 25719 23387 25753
rect 23421 25719 23457 25753
rect 23491 25719 23527 25753
rect 23561 25719 23597 25753
rect 23631 25719 23635 25753
rect 22823 25685 23635 25719
rect 22823 25651 22827 25685
rect 22861 25651 22897 25685
rect 22931 25651 22967 25685
rect 23001 25651 23037 25685
rect 23071 25651 23107 25685
rect 23141 25651 23177 25685
rect 23211 25651 23247 25685
rect 23281 25651 23317 25685
rect 23351 25651 23387 25685
rect 23421 25651 23457 25685
rect 23491 25651 23527 25685
rect 23561 25651 23597 25685
rect 23631 25651 23635 25685
rect 22823 25617 23635 25651
rect 22823 25583 22827 25617
rect 22861 25583 22897 25617
rect 22931 25583 22967 25617
rect 23001 25583 23037 25617
rect 23071 25583 23107 25617
rect 23141 25583 23177 25617
rect 23211 25583 23247 25617
rect 23281 25583 23317 25617
rect 23351 25583 23387 25617
rect 23421 25583 23457 25617
rect 23491 25583 23527 25617
rect 23561 25583 23597 25617
rect 23631 25583 23635 25617
rect 22823 25549 23635 25583
rect 22823 25515 22827 25549
rect 22861 25515 22897 25549
rect 22931 25515 22967 25549
rect 23001 25515 23037 25549
rect 23071 25515 23107 25549
rect 23141 25515 23177 25549
rect 23211 25515 23247 25549
rect 23281 25515 23317 25549
rect 23351 25515 23387 25549
rect 23421 25515 23457 25549
rect 23491 25515 23527 25549
rect 23561 25515 23597 25549
rect 23631 25515 23635 25549
rect 22823 25481 23635 25515
rect 22823 25447 22827 25481
rect 22861 25447 22897 25481
rect 22931 25447 22967 25481
rect 23001 25447 23037 25481
rect 23071 25447 23107 25481
rect 23141 25447 23177 25481
rect 23211 25447 23247 25481
rect 23281 25447 23317 25481
rect 23351 25447 23387 25481
rect 23421 25447 23457 25481
rect 23491 25447 23527 25481
rect 23561 25447 23597 25481
rect 23631 25447 23635 25481
rect 22823 25413 23635 25447
rect 22823 25379 22827 25413
rect 22861 25379 22897 25413
rect 22931 25379 22967 25413
rect 23001 25379 23037 25413
rect 23071 25379 23107 25413
rect 23141 25379 23177 25413
rect 23211 25379 23247 25413
rect 23281 25379 23317 25413
rect 23351 25379 23387 25413
rect 23421 25379 23457 25413
rect 23491 25379 23527 25413
rect 23561 25379 23597 25413
rect 23631 25379 23635 25413
rect 22823 25345 23635 25379
rect 22823 25311 22827 25345
rect 22861 25311 22897 25345
rect 22931 25311 22967 25345
rect 23001 25311 23037 25345
rect 23071 25311 23107 25345
rect 23141 25311 23177 25345
rect 23211 25311 23247 25345
rect 23281 25311 23317 25345
rect 23351 25311 23387 25345
rect 23421 25311 23457 25345
rect 23491 25311 23527 25345
rect 23561 25311 23597 25345
rect 23631 25311 23635 25345
rect 22823 25277 23635 25311
rect 22823 25243 22827 25277
rect 22861 25243 22897 25277
rect 22931 25243 22967 25277
rect 23001 25243 23037 25277
rect 23071 25243 23107 25277
rect 23141 25243 23177 25277
rect 23211 25243 23247 25277
rect 23281 25243 23317 25277
rect 23351 25243 23387 25277
rect 23421 25243 23457 25277
rect 23491 25243 23527 25277
rect 23561 25243 23597 25277
rect 23631 25243 23635 25277
rect 22823 25209 23635 25243
rect 22823 25175 22827 25209
rect 22861 25175 22897 25209
rect 22931 25175 22967 25209
rect 23001 25175 23037 25209
rect 23071 25175 23107 25209
rect 23141 25175 23177 25209
rect 23211 25175 23247 25209
rect 23281 25175 23317 25209
rect 23351 25175 23387 25209
rect 23421 25175 23457 25209
rect 23491 25175 23527 25209
rect 23561 25175 23597 25209
rect 23631 25175 23635 25209
rect 22823 25140 23635 25175
rect 22823 25106 22827 25140
rect 22861 25106 22897 25140
rect 22931 25106 22967 25140
rect 23001 25106 23037 25140
rect 23071 25106 23107 25140
rect 23141 25106 23177 25140
rect 23211 25106 23247 25140
rect 23281 25106 23317 25140
rect 23351 25106 23387 25140
rect 23421 25106 23457 25140
rect 23491 25106 23527 25140
rect 23561 25106 23597 25140
rect 23631 25106 23635 25140
rect 22823 25071 23635 25106
rect 22823 25037 22827 25071
rect 22861 25037 22897 25071
rect 22931 25037 22967 25071
rect 23001 25037 23037 25071
rect 23071 25037 23107 25071
rect 23141 25037 23177 25071
rect 23211 25037 23247 25071
rect 23281 25037 23317 25071
rect 23351 25037 23387 25071
rect 23421 25037 23457 25071
rect 23491 25037 23527 25071
rect 23561 25037 23597 25071
rect 23631 25037 23635 25071
rect 22823 25002 23635 25037
rect 22823 24968 22827 25002
rect 22861 24968 22897 25002
rect 22931 24968 22967 25002
rect 23001 24968 23037 25002
rect 23071 24968 23107 25002
rect 23141 24968 23177 25002
rect 23211 24968 23247 25002
rect 23281 24968 23317 25002
rect 23351 24968 23387 25002
rect 23421 24968 23457 25002
rect 23491 24968 23527 25002
rect 23561 24968 23597 25002
rect 23631 24968 23635 25002
rect 22823 24933 23635 24968
rect 22823 24899 22827 24933
rect 22861 24899 22897 24933
rect 22931 24899 22967 24933
rect 23001 24899 23037 24933
rect 23071 24899 23107 24933
rect 23141 24899 23177 24933
rect 23211 24899 23247 24933
rect 23281 24899 23317 24933
rect 23351 24899 23387 24933
rect 23421 24899 23457 24933
rect 23491 24899 23527 24933
rect 23561 24899 23597 24933
rect 23631 24899 23635 24933
rect 22823 24864 23635 24899
rect 22823 24830 22827 24864
rect 22861 24830 22897 24864
rect 22931 24830 22967 24864
rect 23001 24830 23037 24864
rect 23071 24830 23107 24864
rect 23141 24830 23177 24864
rect 23211 24830 23247 24864
rect 23281 24830 23317 24864
rect 23351 24830 23387 24864
rect 23421 24830 23457 24864
rect 23491 24830 23527 24864
rect 23561 24830 23597 24864
rect 23631 24830 23635 24864
rect 22823 24795 23635 24830
rect 22823 24761 22827 24795
rect 22861 24761 22897 24795
rect 22931 24761 22967 24795
rect 23001 24761 23037 24795
rect 23071 24761 23107 24795
rect 23141 24761 23177 24795
rect 23211 24761 23247 24795
rect 23281 24761 23317 24795
rect 23351 24761 23387 24795
rect 23421 24761 23457 24795
rect 23491 24761 23527 24795
rect 23561 24761 23597 24795
rect 23631 24761 23635 24795
rect 22823 24726 23635 24761
rect 22823 24692 22827 24726
rect 22861 24692 22897 24726
rect 22931 24692 22967 24726
rect 23001 24692 23037 24726
rect 23071 24692 23107 24726
rect 23141 24692 23177 24726
rect 23211 24692 23247 24726
rect 23281 24692 23317 24726
rect 23351 24692 23387 24726
rect 23421 24692 23457 24726
rect 23491 24692 23527 24726
rect 23561 24692 23597 24726
rect 23631 24692 23635 24726
rect 22823 24657 23635 24692
rect 22823 24623 22827 24657
rect 22861 24623 22897 24657
rect 22931 24623 22967 24657
rect 23001 24623 23037 24657
rect 23071 24623 23107 24657
rect 23141 24623 23177 24657
rect 23211 24623 23247 24657
rect 23281 24623 23317 24657
rect 23351 24623 23387 24657
rect 23421 24623 23457 24657
rect 23491 24623 23527 24657
rect 23561 24623 23597 24657
rect 23631 24623 23635 24657
rect 22823 24588 23635 24623
rect 22823 24554 22827 24588
rect 22861 24554 22897 24588
rect 22931 24554 22967 24588
rect 23001 24554 23037 24588
rect 23071 24554 23107 24588
rect 23141 24554 23177 24588
rect 23211 24554 23247 24588
rect 23281 24554 23317 24588
rect 23351 24554 23387 24588
rect 23421 24554 23457 24588
rect 23491 24554 23527 24588
rect 23561 24554 23597 24588
rect 23631 24554 23635 24588
rect 22823 24519 23635 24554
rect 22823 24485 22827 24519
rect 22861 24485 22897 24519
rect 22931 24485 22967 24519
rect 23001 24485 23037 24519
rect 23071 24485 23107 24519
rect 23141 24485 23177 24519
rect 23211 24485 23247 24519
rect 23281 24485 23317 24519
rect 23351 24485 23387 24519
rect 23421 24485 23457 24519
rect 23491 24485 23527 24519
rect 23561 24485 23597 24519
rect 23631 24485 23635 24519
rect 22823 24450 23635 24485
rect 22823 24416 22827 24450
rect 22861 24416 22897 24450
rect 22931 24416 22967 24450
rect 23001 24416 23037 24450
rect 23071 24416 23107 24450
rect 23141 24416 23177 24450
rect 23211 24416 23247 24450
rect 23281 24416 23317 24450
rect 23351 24416 23387 24450
rect 23421 24416 23457 24450
rect 23491 24416 23527 24450
rect 23561 24416 23597 24450
rect 23631 24416 23635 24450
rect 22823 24381 23635 24416
rect 22823 24347 22827 24381
rect 22861 24347 22897 24381
rect 22931 24347 22967 24381
rect 23001 24347 23037 24381
rect 23071 24347 23107 24381
rect 23141 24347 23177 24381
rect 23211 24347 23247 24381
rect 23281 24347 23317 24381
rect 23351 24347 23387 24381
rect 23421 24347 23457 24381
rect 23491 24347 23527 24381
rect 23561 24347 23597 24381
rect 23631 24347 23635 24381
rect 22823 24312 23635 24347
rect 22823 24278 22827 24312
rect 22861 24278 22897 24312
rect 22931 24278 22967 24312
rect 23001 24278 23037 24312
rect 23071 24278 23107 24312
rect 23141 24278 23177 24312
rect 23211 24278 23247 24312
rect 23281 24278 23317 24312
rect 23351 24278 23387 24312
rect 23421 24278 23457 24312
rect 23491 24278 23527 24312
rect 23561 24278 23597 24312
rect 23631 24278 23635 24312
rect 22823 24243 23635 24278
rect 22823 24209 22827 24243
rect 22861 24209 22897 24243
rect 22931 24209 22967 24243
rect 23001 24209 23037 24243
rect 23071 24209 23107 24243
rect 23141 24209 23177 24243
rect 23211 24209 23247 24243
rect 23281 24209 23317 24243
rect 23351 24209 23387 24243
rect 23421 24209 23457 24243
rect 23491 24209 23527 24243
rect 23561 24209 23597 24243
rect 23631 24209 23635 24243
rect 22823 24174 23635 24209
rect 22823 24140 22827 24174
rect 22861 24140 22897 24174
rect 22931 24140 22967 24174
rect 23001 24140 23037 24174
rect 23071 24140 23107 24174
rect 23141 24140 23177 24174
rect 23211 24140 23247 24174
rect 23281 24140 23317 24174
rect 23351 24140 23387 24174
rect 23421 24140 23457 24174
rect 23491 24140 23527 24174
rect 23561 24140 23597 24174
rect 23631 24140 23635 24174
rect 22823 24105 23635 24140
rect 22823 24071 22827 24105
rect 22861 24071 22897 24105
rect 22931 24071 22967 24105
rect 23001 24071 23037 24105
rect 23071 24071 23107 24105
rect 23141 24071 23177 24105
rect 23211 24071 23247 24105
rect 23281 24071 23317 24105
rect 23351 24071 23387 24105
rect 23421 24071 23457 24105
rect 23491 24071 23527 24105
rect 23561 24071 23597 24105
rect 23631 24071 23635 24105
rect 22823 24036 23635 24071
rect 22823 24002 22827 24036
rect 22861 24002 22897 24036
rect 22931 24002 22967 24036
rect 23001 24002 23037 24036
rect 23071 24002 23107 24036
rect 23141 24002 23177 24036
rect 23211 24002 23247 24036
rect 23281 24002 23317 24036
rect 23351 24002 23387 24036
rect 23421 24002 23457 24036
rect 23491 24002 23527 24036
rect 23561 24002 23597 24036
rect 23631 24002 23635 24036
rect 22823 23967 23635 24002
rect 22823 23933 22827 23967
rect 22861 23933 22897 23967
rect 22931 23933 22967 23967
rect 23001 23933 23037 23967
rect 23071 23933 23107 23967
rect 23141 23933 23177 23967
rect 23211 23933 23247 23967
rect 23281 23933 23317 23967
rect 23351 23933 23387 23967
rect 23421 23933 23457 23967
rect 23491 23933 23527 23967
rect 23561 23933 23597 23967
rect 23631 23933 23635 23967
rect 22823 23898 23635 23933
rect 22823 23864 22827 23898
rect 22861 23864 22897 23898
rect 22931 23864 22967 23898
rect 23001 23864 23037 23898
rect 23071 23864 23107 23898
rect 23141 23864 23177 23898
rect 23211 23864 23247 23898
rect 23281 23864 23317 23898
rect 23351 23864 23387 23898
rect 23421 23864 23457 23898
rect 23491 23864 23527 23898
rect 23561 23864 23597 23898
rect 23631 23864 23635 23898
rect 22823 23829 23635 23864
rect 22823 23795 22827 23829
rect 22861 23795 22897 23829
rect 22931 23795 22967 23829
rect 23001 23795 23037 23829
rect 23071 23795 23107 23829
rect 23141 23795 23177 23829
rect 23211 23795 23247 23829
rect 23281 23795 23317 23829
rect 23351 23795 23387 23829
rect 23421 23795 23457 23829
rect 23491 23795 23527 23829
rect 23561 23795 23597 23829
rect 23631 23795 23635 23829
rect 22823 23760 23635 23795
rect 22823 23726 22827 23760
rect 22861 23726 22897 23760
rect 22931 23726 22967 23760
rect 23001 23726 23037 23760
rect 23071 23726 23107 23760
rect 23141 23726 23177 23760
rect 23211 23726 23247 23760
rect 23281 23726 23317 23760
rect 23351 23726 23387 23760
rect 23421 23726 23457 23760
rect 23491 23726 23527 23760
rect 23561 23726 23597 23760
rect 23631 23726 23635 23760
rect 22823 23691 23635 23726
rect 22823 23657 22827 23691
rect 22861 23657 22897 23691
rect 22931 23657 22967 23691
rect 23001 23657 23037 23691
rect 23071 23657 23107 23691
rect 23141 23657 23177 23691
rect 23211 23657 23247 23691
rect 23281 23657 23317 23691
rect 23351 23657 23387 23691
rect 23421 23657 23457 23691
rect 23491 23657 23527 23691
rect 23561 23657 23597 23691
rect 23631 23657 23635 23691
rect 22823 23622 23635 23657
rect 22823 23588 22827 23622
rect 22861 23588 22897 23622
rect 22931 23588 22967 23622
rect 23001 23588 23037 23622
rect 23071 23588 23107 23622
rect 23141 23588 23177 23622
rect 23211 23588 23247 23622
rect 23281 23588 23317 23622
rect 23351 23588 23387 23622
rect 23421 23588 23457 23622
rect 23491 23588 23527 23622
rect 23561 23588 23597 23622
rect 23631 23588 23635 23622
rect 22823 23553 23635 23588
rect 22823 23519 22827 23553
rect 22861 23519 22897 23553
rect 22931 23519 22967 23553
rect 23001 23519 23037 23553
rect 23071 23519 23107 23553
rect 23141 23519 23177 23553
rect 23211 23519 23247 23553
rect 23281 23519 23317 23553
rect 23351 23519 23387 23553
rect 23421 23519 23457 23553
rect 23491 23519 23527 23553
rect 23561 23519 23597 23553
rect 23631 23519 23635 23553
rect 280 23439 314 23473
rect 348 23439 384 23473
rect 418 23439 454 23473
rect 488 23439 524 23473
rect 558 23439 594 23473
rect 628 23439 664 23473
rect 698 23439 734 23473
rect 768 23439 804 23473
rect 838 23439 874 23473
rect 908 23439 944 23473
rect 978 23439 1014 23473
rect 1048 23439 1084 23473
rect 1118 23439 1154 23473
rect 1188 23439 1224 23473
rect 1258 23439 1294 23473
rect 1328 23439 1364 23473
rect 1398 23439 1434 23473
rect 1468 23439 1502 23473
rect 280 23403 1502 23439
rect 280 23369 314 23403
rect 348 23369 384 23403
rect 418 23369 454 23403
rect 488 23369 524 23403
rect 558 23369 594 23403
rect 628 23369 664 23403
rect 698 23369 734 23403
rect 768 23369 804 23403
rect 838 23369 874 23403
rect 908 23369 944 23403
rect 978 23369 1014 23403
rect 1048 23369 1084 23403
rect 1118 23369 1154 23403
rect 1188 23369 1224 23403
rect 1258 23369 1294 23403
rect 1328 23369 1364 23403
rect 1398 23369 1434 23403
rect 1468 23369 1502 23403
rect 280 23333 1502 23369
rect 280 23299 314 23333
rect 348 23299 384 23333
rect 418 23299 454 23333
rect 488 23299 524 23333
rect 558 23299 594 23333
rect 628 23299 664 23333
rect 698 23299 734 23333
rect 768 23299 804 23333
rect 838 23299 874 23333
rect 908 23299 944 23333
rect 978 23299 1014 23333
rect 1048 23299 1084 23333
rect 1118 23299 1154 23333
rect 1188 23299 1224 23333
rect 1258 23299 1294 23333
rect 1328 23299 1364 23333
rect 1398 23299 1434 23333
rect 1468 23299 1502 23333
rect 280 23263 1502 23299
rect 280 23229 314 23263
rect 348 23229 384 23263
rect 418 23229 454 23263
rect 488 23229 524 23263
rect 558 23229 594 23263
rect 628 23229 664 23263
rect 698 23229 734 23263
rect 768 23229 804 23263
rect 838 23229 874 23263
rect 908 23229 944 23263
rect 978 23229 1014 23263
rect 1048 23229 1084 23263
rect 1118 23229 1154 23263
rect 1188 23229 1224 23263
rect 1258 23229 1294 23263
rect 1328 23229 1364 23263
rect 1398 23229 1434 23263
rect 1468 23229 1502 23263
rect 280 23193 1502 23229
rect 280 23159 314 23193
rect 348 23159 384 23193
rect 418 23159 454 23193
rect 488 23159 524 23193
rect 558 23159 594 23193
rect 628 23159 664 23193
rect 698 23159 734 23193
rect 768 23159 804 23193
rect 838 23159 874 23193
rect 908 23159 944 23193
rect 978 23159 1014 23193
rect 1048 23159 1084 23193
rect 1118 23159 1154 23193
rect 1188 23159 1224 23193
rect 1258 23159 1294 23193
rect 1328 23159 1364 23193
rect 1398 23159 1434 23193
rect 1468 23159 1502 23193
rect 280 23123 1502 23159
rect 280 23089 314 23123
rect 348 23089 384 23123
rect 418 23089 454 23123
rect 488 23089 524 23123
rect 558 23089 594 23123
rect 628 23089 664 23123
rect 698 23089 734 23123
rect 768 23089 804 23123
rect 838 23089 874 23123
rect 908 23089 944 23123
rect 978 23089 1014 23123
rect 1048 23089 1084 23123
rect 1118 23089 1154 23123
rect 1188 23089 1224 23123
rect 1258 23089 1294 23123
rect 1328 23089 1364 23123
rect 1398 23089 1434 23123
rect 1468 23089 1502 23123
rect 280 23053 1502 23089
rect 280 23019 314 23053
rect 348 23019 384 23053
rect 418 23019 454 23053
rect 488 23019 524 23053
rect 558 23019 594 23053
rect 628 23019 664 23053
rect 698 23019 734 23053
rect 768 23019 804 23053
rect 838 23019 874 23053
rect 908 23019 944 23053
rect 978 23019 1014 23053
rect 1048 23019 1084 23053
rect 1118 23019 1154 23053
rect 1188 23019 1224 23053
rect 1258 23019 1294 23053
rect 1328 23019 1364 23053
rect 1398 23019 1434 23053
rect 1468 23019 1502 23053
rect 280 22983 1502 23019
rect 280 22949 314 22983
rect 348 22949 384 22983
rect 418 22949 454 22983
rect 488 22949 524 22983
rect 558 22949 594 22983
rect 628 22949 664 22983
rect 698 22949 734 22983
rect 768 22949 804 22983
rect 838 22949 874 22983
rect 908 22949 944 22983
rect 978 22949 1014 22983
rect 1048 22949 1084 22983
rect 1118 22949 1154 22983
rect 1188 22949 1224 22983
rect 1258 22949 1294 22983
rect 1328 22949 1364 22983
rect 1398 22949 1434 22983
rect 1468 22949 1502 22983
rect 280 22913 1502 22949
rect 280 22879 314 22913
rect 348 22879 384 22913
rect 418 22879 454 22913
rect 488 22879 524 22913
rect 558 22879 594 22913
rect 628 22879 664 22913
rect 698 22879 734 22913
rect 768 22879 804 22913
rect 838 22879 874 22913
rect 908 22879 944 22913
rect 978 22879 1014 22913
rect 1048 22879 1084 22913
rect 1118 22879 1154 22913
rect 1188 22879 1224 22913
rect 1258 22879 1294 22913
rect 1328 22879 1364 22913
rect 1398 22879 1434 22913
rect 1468 22879 1502 22913
rect 280 22843 1502 22879
rect 280 22809 314 22843
rect 348 22809 384 22843
rect 418 22809 454 22843
rect 488 22809 524 22843
rect 558 22809 594 22843
rect 628 22809 664 22843
rect 698 22809 734 22843
rect 768 22809 804 22843
rect 838 22809 874 22843
rect 908 22809 944 22843
rect 978 22809 1014 22843
rect 1048 22809 1084 22843
rect 1118 22809 1154 22843
rect 1188 22809 1224 22843
rect 1258 22809 1294 22843
rect 1328 22809 1364 22843
rect 1398 22809 1434 22843
rect 1468 22809 1502 22843
rect 280 22773 1502 22809
rect 280 22739 314 22773
rect 348 22739 384 22773
rect 418 22739 454 22773
rect 488 22739 524 22773
rect 558 22739 594 22773
rect 628 22739 664 22773
rect 698 22739 734 22773
rect 768 22739 804 22773
rect 838 22739 874 22773
rect 908 22739 944 22773
rect 978 22739 1014 22773
rect 1048 22739 1084 22773
rect 1118 22739 1154 22773
rect 1188 22739 1224 22773
rect 1258 22739 1294 22773
rect 1328 22739 1364 22773
rect 1398 22739 1434 22773
rect 1468 22739 1502 22773
rect 280 22702 1502 22739
rect 280 22668 314 22702
rect 348 22668 384 22702
rect 418 22668 454 22702
rect 488 22668 524 22702
rect 558 22668 594 22702
rect 628 22668 664 22702
rect 698 22668 734 22702
rect 768 22668 804 22702
rect 838 22668 874 22702
rect 908 22668 944 22702
rect 978 22668 1014 22702
rect 1048 22668 1084 22702
rect 1118 22668 1154 22702
rect 1188 22668 1224 22702
rect 1258 22668 1294 22702
rect 1328 22668 1364 22702
rect 1398 22668 1434 22702
rect 1468 22668 1502 22702
rect 280 22631 1502 22668
rect 280 22597 314 22631
rect 348 22597 384 22631
rect 418 22597 454 22631
rect 488 22597 524 22631
rect 558 22597 594 22631
rect 628 22597 664 22631
rect 698 22597 734 22631
rect 768 22597 804 22631
rect 838 22597 874 22631
rect 908 22597 944 22631
rect 978 22597 1014 22631
rect 1048 22597 1084 22631
rect 1118 22597 1154 22631
rect 1188 22597 1224 22631
rect 1258 22597 1294 22631
rect 1328 22597 1364 22631
rect 1398 22597 1434 22631
rect 1468 22597 1502 22631
rect 280 22560 1502 22597
rect 280 22526 314 22560
rect 348 22526 384 22560
rect 418 22526 454 22560
rect 488 22526 524 22560
rect 558 22526 594 22560
rect 628 22526 664 22560
rect 698 22526 734 22560
rect 768 22526 804 22560
rect 838 22526 874 22560
rect 908 22526 944 22560
rect 978 22526 1014 22560
rect 1048 22526 1084 22560
rect 1118 22526 1154 22560
rect 1188 22526 1224 22560
rect 1258 22526 1294 22560
rect 1328 22526 1364 22560
rect 1398 22526 1434 22560
rect 1468 22526 1502 22560
rect 280 22489 1502 22526
rect 280 22455 314 22489
rect 348 22455 384 22489
rect 418 22455 454 22489
rect 488 22455 524 22489
rect 558 22455 594 22489
rect 628 22455 664 22489
rect 698 22455 734 22489
rect 768 22455 804 22489
rect 838 22455 874 22489
rect 908 22455 944 22489
rect 978 22455 1014 22489
rect 1048 22455 1084 22489
rect 1118 22455 1154 22489
rect 1188 22455 1224 22489
rect 1258 22455 1294 22489
rect 1328 22455 1364 22489
rect 1398 22455 1434 22489
rect 1468 22455 1502 22489
rect 280 22418 1502 22455
rect 280 22384 314 22418
rect 348 22384 384 22418
rect 418 22384 454 22418
rect 488 22384 524 22418
rect 558 22384 594 22418
rect 628 22384 664 22418
rect 698 22384 734 22418
rect 768 22384 804 22418
rect 838 22384 874 22418
rect 908 22384 944 22418
rect 978 22384 1014 22418
rect 1048 22384 1084 22418
rect 1118 22384 1154 22418
rect 1188 22384 1224 22418
rect 1258 22384 1294 22418
rect 1328 22384 1364 22418
rect 1398 22384 1434 22418
rect 1468 22384 1502 22418
rect 280 22347 1502 22384
rect 280 22313 314 22347
rect 348 22313 384 22347
rect 418 22313 454 22347
rect 488 22313 524 22347
rect 558 22313 594 22347
rect 628 22313 664 22347
rect 698 22313 734 22347
rect 768 22313 804 22347
rect 838 22313 874 22347
rect 908 22313 944 22347
rect 978 22313 1014 22347
rect 1048 22313 1084 22347
rect 1118 22313 1154 22347
rect 1188 22313 1224 22347
rect 1258 22313 1294 22347
rect 1328 22313 1364 22347
rect 1398 22313 1434 22347
rect 1468 22313 1502 22347
rect 280 22289 1502 22313
rect 22823 23484 23635 23519
rect 22823 23450 22827 23484
rect 22861 23450 22897 23484
rect 22931 23450 22967 23484
rect 23001 23450 23037 23484
rect 23071 23450 23107 23484
rect 23141 23450 23177 23484
rect 23211 23450 23247 23484
rect 23281 23450 23317 23484
rect 23351 23450 23387 23484
rect 23421 23450 23457 23484
rect 23491 23450 23527 23484
rect 23561 23450 23597 23484
rect 23631 23450 23635 23484
rect 22823 23415 23635 23450
rect 22823 23381 22827 23415
rect 22861 23381 22897 23415
rect 22931 23381 22967 23415
rect 23001 23381 23037 23415
rect 23071 23381 23107 23415
rect 23141 23381 23177 23415
rect 23211 23381 23247 23415
rect 23281 23381 23317 23415
rect 23351 23381 23387 23415
rect 23421 23381 23457 23415
rect 23491 23381 23527 23415
rect 23561 23381 23597 23415
rect 23631 23381 23635 23415
rect 22823 23346 23635 23381
rect 22823 23312 22827 23346
rect 22861 23312 22897 23346
rect 22931 23312 22967 23346
rect 23001 23312 23037 23346
rect 23071 23312 23107 23346
rect 23141 23312 23177 23346
rect 23211 23312 23247 23346
rect 23281 23312 23317 23346
rect 23351 23312 23387 23346
rect 23421 23312 23457 23346
rect 23491 23312 23527 23346
rect 23561 23312 23597 23346
rect 23631 23312 23635 23346
rect 22823 23277 23635 23312
rect 22823 23243 22827 23277
rect 22861 23243 22897 23277
rect 22931 23243 22967 23277
rect 23001 23243 23037 23277
rect 23071 23243 23107 23277
rect 23141 23243 23177 23277
rect 23211 23243 23247 23277
rect 23281 23243 23317 23277
rect 23351 23243 23387 23277
rect 23421 23243 23457 23277
rect 23491 23243 23527 23277
rect 23561 23243 23597 23277
rect 23631 23243 23635 23277
rect 22823 23208 23635 23243
rect 22823 23174 22827 23208
rect 22861 23174 22897 23208
rect 22931 23174 22967 23208
rect 23001 23174 23037 23208
rect 23071 23174 23107 23208
rect 23141 23174 23177 23208
rect 23211 23174 23247 23208
rect 23281 23174 23317 23208
rect 23351 23174 23387 23208
rect 23421 23174 23457 23208
rect 23491 23174 23527 23208
rect 23561 23174 23597 23208
rect 23631 23174 23635 23208
rect 22823 23139 23635 23174
rect 22823 23105 22827 23139
rect 22861 23105 22897 23139
rect 22931 23105 22967 23139
rect 23001 23105 23037 23139
rect 23071 23105 23107 23139
rect 23141 23105 23177 23139
rect 23211 23105 23247 23139
rect 23281 23105 23317 23139
rect 23351 23105 23387 23139
rect 23421 23105 23457 23139
rect 23491 23105 23527 23139
rect 23561 23105 23597 23139
rect 23631 23105 23635 23139
rect 22823 23070 23635 23105
rect 22823 23036 22827 23070
rect 22861 23036 22897 23070
rect 22931 23036 22967 23070
rect 23001 23036 23037 23070
rect 23071 23036 23107 23070
rect 23141 23036 23177 23070
rect 23211 23036 23247 23070
rect 23281 23036 23317 23070
rect 23351 23036 23387 23070
rect 23421 23036 23457 23070
rect 23491 23036 23527 23070
rect 23561 23036 23597 23070
rect 23631 23036 23635 23070
rect 22823 23001 23635 23036
rect 22823 22967 22827 23001
rect 22861 22967 22897 23001
rect 22931 22967 22967 23001
rect 23001 22967 23037 23001
rect 23071 22967 23107 23001
rect 23141 22967 23177 23001
rect 23211 22967 23247 23001
rect 23281 22967 23317 23001
rect 23351 22967 23387 23001
rect 23421 22967 23457 23001
rect 23491 22967 23527 23001
rect 23561 22967 23597 23001
rect 23631 22967 23635 23001
rect 22823 22932 23635 22967
rect 22823 22898 22827 22932
rect 22861 22898 22897 22932
rect 22931 22898 22967 22932
rect 23001 22898 23037 22932
rect 23071 22898 23107 22932
rect 23141 22898 23177 22932
rect 23211 22898 23247 22932
rect 23281 22898 23317 22932
rect 23351 22898 23387 22932
rect 23421 22898 23457 22932
rect 23491 22898 23527 22932
rect 23561 22898 23597 22932
rect 23631 22898 23635 22932
rect 22823 22863 23635 22898
rect 22823 22829 22827 22863
rect 22861 22829 22897 22863
rect 22931 22829 22967 22863
rect 23001 22829 23037 22863
rect 23071 22829 23107 22863
rect 23141 22829 23177 22863
rect 23211 22829 23247 22863
rect 23281 22829 23317 22863
rect 23351 22829 23387 22863
rect 23421 22829 23457 22863
rect 23491 22829 23527 22863
rect 23561 22829 23597 22863
rect 23631 22829 23635 22863
rect 22823 22794 23635 22829
rect 22823 22760 22827 22794
rect 22861 22760 22897 22794
rect 22931 22760 22967 22794
rect 23001 22760 23037 22794
rect 23071 22760 23107 22794
rect 23141 22760 23177 22794
rect 23211 22760 23247 22794
rect 23281 22760 23317 22794
rect 23351 22760 23387 22794
rect 23421 22760 23457 22794
rect 23491 22760 23527 22794
rect 23561 22760 23597 22794
rect 23631 22760 23635 22794
rect 22823 22725 23635 22760
rect 22823 22691 22827 22725
rect 22861 22691 22897 22725
rect 22931 22691 22967 22725
rect 23001 22691 23037 22725
rect 23071 22691 23107 22725
rect 23141 22691 23177 22725
rect 23211 22691 23247 22725
rect 23281 22691 23317 22725
rect 23351 22691 23387 22725
rect 23421 22691 23457 22725
rect 23491 22691 23527 22725
rect 23561 22691 23597 22725
rect 23631 22691 23635 22725
rect 22823 22656 23635 22691
rect 22823 22622 22827 22656
rect 22861 22622 22897 22656
rect 22931 22622 22967 22656
rect 23001 22622 23037 22656
rect 23071 22622 23107 22656
rect 23141 22622 23177 22656
rect 23211 22622 23247 22656
rect 23281 22622 23317 22656
rect 23351 22622 23387 22656
rect 23421 22622 23457 22656
rect 23491 22622 23527 22656
rect 23561 22622 23597 22656
rect 23631 22622 23635 22656
rect 22823 22587 23635 22622
rect 22823 22553 22827 22587
rect 22861 22553 22897 22587
rect 22931 22553 22967 22587
rect 23001 22553 23037 22587
rect 23071 22553 23107 22587
rect 23141 22553 23177 22587
rect 23211 22553 23247 22587
rect 23281 22553 23317 22587
rect 23351 22553 23387 22587
rect 23421 22553 23457 22587
rect 23491 22553 23527 22587
rect 23561 22553 23597 22587
rect 23631 22553 23635 22587
rect 22823 22518 23635 22553
rect 22823 22484 22827 22518
rect 22861 22484 22897 22518
rect 22931 22484 22967 22518
rect 23001 22484 23037 22518
rect 23071 22484 23107 22518
rect 23141 22484 23177 22518
rect 23211 22484 23247 22518
rect 23281 22484 23317 22518
rect 23351 22484 23387 22518
rect 23421 22484 23457 22518
rect 23491 22484 23527 22518
rect 23561 22484 23597 22518
rect 23631 22484 23635 22518
rect 22823 22449 23635 22484
rect 22823 22415 22827 22449
rect 22861 22415 22897 22449
rect 22931 22415 22967 22449
rect 23001 22415 23037 22449
rect 23071 22415 23107 22449
rect 23141 22415 23177 22449
rect 23211 22415 23247 22449
rect 23281 22415 23317 22449
rect 23351 22415 23387 22449
rect 23421 22415 23457 22449
rect 23491 22415 23527 22449
rect 23561 22415 23597 22449
rect 23631 22415 23635 22449
rect 22823 22380 23635 22415
rect 22823 22346 22827 22380
rect 22861 22346 22897 22380
rect 22931 22346 22967 22380
rect 23001 22346 23037 22380
rect 23071 22346 23107 22380
rect 23141 22346 23177 22380
rect 23211 22346 23247 22380
rect 23281 22346 23317 22380
rect 23351 22346 23387 22380
rect 23421 22346 23457 22380
rect 23491 22346 23527 22380
rect 23561 22346 23597 22380
rect 23631 22346 23635 22380
rect 22823 22311 23635 22346
rect 714 22213 1020 22289
rect 22823 22277 22827 22311
rect 22861 22277 22897 22311
rect 22931 22277 22967 22311
rect 23001 22277 23037 22311
rect 23071 22277 23107 22311
rect 23141 22277 23177 22311
rect 23211 22277 23247 22311
rect 23281 22277 23317 22311
rect 23351 22277 23387 22311
rect 23421 22277 23457 22311
rect 23491 22277 23527 22311
rect 23561 22277 23597 22311
rect 23631 22277 23635 22311
rect 22823 22242 23635 22277
rect 22823 22208 22827 22242
rect 22861 22208 22897 22242
rect 22931 22208 22967 22242
rect 23001 22208 23037 22242
rect 23071 22208 23107 22242
rect 23141 22208 23177 22242
rect 23211 22208 23247 22242
rect 23281 22208 23317 22242
rect 23351 22208 23387 22242
rect 23421 22208 23457 22242
rect 23491 22208 23527 22242
rect 23561 22208 23597 22242
rect 23631 22208 23635 22242
rect 22823 22173 23635 22208
rect 22823 22139 22827 22173
rect 22861 22139 22897 22173
rect 22931 22139 22967 22173
rect 23001 22139 23037 22173
rect 23071 22139 23107 22173
rect 23141 22139 23177 22173
rect 23211 22139 23247 22173
rect 23281 22139 23317 22173
rect 23351 22139 23387 22173
rect 23421 22139 23457 22173
rect 23491 22139 23527 22173
rect 23561 22139 23597 22173
rect 23631 22139 23635 22173
rect 22823 22115 23635 22139
rect 714 17384 1020 17419
rect 748 17350 782 17384
rect 816 17350 850 17384
rect 884 17350 918 17384
rect 952 17350 986 17384
rect 714 17315 1020 17350
rect 748 17281 782 17315
rect 816 17281 850 17315
rect 884 17281 918 17315
rect 952 17281 986 17315
rect 714 17246 1020 17281
rect 748 17212 782 17246
rect 816 17212 850 17246
rect 884 17212 918 17246
rect 952 17212 986 17246
rect 714 17177 1020 17212
rect 748 17143 782 17177
rect 816 17143 850 17177
rect 884 17143 918 17177
rect 952 17143 986 17177
rect 714 17108 1020 17143
rect 748 17074 782 17108
rect 816 17074 850 17108
rect 884 17074 918 17108
rect 952 17074 986 17108
rect 714 17039 1020 17074
rect 748 17005 782 17039
rect 816 17005 850 17039
rect 884 17005 918 17039
rect 952 17005 986 17039
rect 714 16970 1020 17005
rect 748 16936 782 16970
rect 816 16936 850 16970
rect 884 16936 918 16970
rect 952 16936 986 16970
rect 714 16901 1020 16936
rect 748 16867 782 16901
rect 816 16867 850 16901
rect 884 16867 918 16901
rect 952 16867 986 16901
rect 714 16832 1020 16867
rect 748 16798 782 16832
rect 816 16798 850 16832
rect 884 16798 918 16832
rect 952 16798 986 16832
rect 714 16763 1020 16798
rect 748 16729 782 16763
rect 816 16729 850 16763
rect 884 16729 918 16763
rect 952 16729 986 16763
rect 714 16694 1020 16729
rect 748 16660 782 16694
rect 816 16660 850 16694
rect 884 16660 918 16694
rect 952 16660 986 16694
rect 714 16625 1020 16660
rect 748 16591 782 16625
rect 816 16591 850 16625
rect 884 16591 918 16625
rect 952 16591 986 16625
rect 714 16556 1020 16591
rect 748 16522 782 16556
rect 816 16522 850 16556
rect 884 16522 918 16556
rect 952 16522 986 16556
rect 714 16487 1020 16522
rect 748 16453 782 16487
rect 816 16453 850 16487
rect 884 16453 918 16487
rect 952 16453 986 16487
rect 714 16418 1020 16453
rect 748 16384 782 16418
rect 816 16384 850 16418
rect 884 16384 918 16418
rect 952 16384 986 16418
rect 714 16349 1020 16384
rect 748 16315 782 16349
rect 816 16315 850 16349
rect 884 16315 918 16349
rect 952 16315 986 16349
rect 714 16280 1020 16315
rect 748 16246 782 16280
rect 816 16246 850 16280
rect 884 16246 918 16280
rect 952 16246 986 16280
rect 714 16222 1020 16246
rect 19676 11622 19797 11629
rect 6746 11618 16309 11622
rect 6746 11584 6770 11618
rect 6804 11584 6839 11618
rect 6873 11584 6908 11618
rect 6942 11584 6977 11618
rect 7011 11584 7046 11618
rect 7080 11584 7115 11618
rect 7149 11584 7184 11618
rect 7218 11584 7253 11618
rect 7287 11584 7322 11618
rect 7356 11584 7391 11618
rect 7425 11584 7460 11618
rect 7494 11584 7529 11618
rect 7563 11584 7598 11618
rect 7632 11584 7667 11618
rect 7701 11584 7736 11618
rect 7770 11584 7805 11618
rect 7839 11584 7874 11618
rect 7908 11584 7943 11618
rect 7977 11584 8012 11618
rect 8046 11584 8081 11618
rect 8115 11584 8150 11618
rect 8184 11584 8219 11618
rect 8253 11584 8288 11618
rect 8322 11584 8357 11618
rect 8391 11584 8426 11618
rect 8460 11584 8495 11618
rect 8529 11584 8564 11618
rect 8598 11584 8633 11618
rect 8667 11584 8702 11618
rect 8736 11584 8771 11618
rect 8805 11584 8840 11618
rect 8874 11584 8909 11618
rect 8943 11584 8978 11618
rect 9012 11584 9046 11618
rect 9080 11584 9114 11618
rect 9148 11584 9182 11618
rect 9216 11584 9250 11618
rect 9284 11584 9318 11618
rect 9352 11584 9386 11618
rect 9420 11584 9454 11618
rect 9488 11584 9522 11618
rect 9556 11584 9590 11618
rect 9624 11584 9658 11618
rect 9692 11584 9726 11618
rect 9760 11584 9794 11618
rect 9828 11584 9862 11618
rect 9896 11584 9930 11618
rect 9964 11584 9998 11618
rect 10032 11584 10066 11618
rect 10100 11584 10134 11618
rect 10168 11584 10202 11618
rect 10236 11584 10270 11618
rect 10304 11588 16309 11618
rect 16343 11588 16379 11622
rect 16413 11588 16449 11622
rect 16483 11588 16519 11622
rect 16553 11588 16589 11622
rect 16623 11588 16658 11622
rect 16692 11588 16727 11622
rect 16761 11588 16796 11622
rect 16830 11588 16865 11622
rect 16899 11588 16934 11622
rect 16968 11588 17003 11622
rect 17037 11588 17072 11622
rect 17106 11588 17141 11622
rect 17175 11588 17210 11622
rect 17244 11588 17279 11622
rect 17313 11588 17348 11622
rect 17382 11588 17417 11622
rect 17451 11588 17486 11622
rect 17520 11588 17555 11622
rect 17589 11588 17624 11622
rect 17658 11588 17693 11622
rect 17727 11588 17762 11622
rect 17796 11588 17831 11622
rect 17865 11588 17900 11622
rect 17934 11588 17969 11622
rect 18003 11588 18038 11622
rect 18072 11588 18107 11622
rect 18141 11588 18176 11622
rect 18210 11588 18245 11622
rect 18279 11588 18314 11622
rect 18348 11588 18383 11622
rect 18417 11588 18452 11622
rect 18486 11588 18521 11622
rect 18555 11588 18590 11622
rect 18624 11588 18659 11622
rect 18693 11588 18728 11622
rect 18762 11588 18797 11622
rect 18831 11588 18866 11622
rect 18900 11588 18935 11622
rect 18969 11588 19004 11622
rect 19038 11588 19073 11622
rect 19107 11588 19142 11622
rect 19176 11588 19211 11622
rect 19245 11588 19280 11622
rect 19314 11588 19349 11622
rect 19383 11588 19418 11622
rect 19452 11588 19487 11622
rect 19521 11588 19556 11622
rect 19590 11588 19625 11622
rect 19659 11595 19797 11622
rect 19831 11595 19866 11629
rect 19900 11595 19935 11629
rect 19969 11595 20004 11629
rect 20038 11595 20073 11629
rect 20107 11595 20142 11629
rect 20176 11595 20211 11629
rect 20245 11595 20280 11629
rect 20314 11595 20349 11629
rect 20383 11595 20418 11629
rect 20452 11595 20487 11629
rect 20521 11595 20556 11629
rect 20590 11595 20625 11629
rect 20659 11595 20694 11629
rect 20728 11595 20763 11629
rect 20797 11595 20832 11629
rect 20866 11595 20901 11629
rect 20935 11595 20970 11629
rect 21004 11595 21039 11629
rect 21073 11595 21108 11629
rect 21142 11595 21177 11629
rect 21211 11595 21246 11629
rect 21280 11595 21315 11629
rect 21349 11595 21384 11629
rect 21418 11595 21453 11629
rect 21487 11595 21522 11629
rect 21556 11595 21591 11629
rect 21625 11595 21660 11629
rect 21694 11595 21729 11629
rect 21763 11595 21798 11629
rect 21832 11595 21866 11629
rect 21900 11595 21934 11629
rect 21968 11595 22002 11629
rect 22036 11595 22070 11629
rect 22104 11595 22138 11629
rect 22172 11595 22206 11629
rect 22240 11595 22274 11629
rect 22308 11595 22342 11629
rect 22376 11595 22410 11629
rect 22444 11595 22478 11629
rect 22512 11595 22546 11629
rect 22580 11595 22614 11629
rect 22648 11595 22682 11629
rect 22716 11595 22750 11629
rect 22784 11595 22818 11629
rect 22852 11595 22886 11629
rect 22920 11595 22954 11629
rect 22988 11595 23022 11629
rect 23056 11595 23090 11629
rect 23124 11595 23158 11629
rect 23192 11595 23226 11629
rect 23260 11595 23294 11629
rect 23328 11595 23362 11629
rect 23396 11595 23430 11629
rect 23464 11595 23498 11629
rect 23532 11595 23566 11629
rect 23600 11595 23634 11629
rect 23668 11595 23702 11629
rect 23736 11595 23770 11629
rect 23804 11595 23838 11629
rect 23872 11595 23906 11629
rect 23940 11595 23974 11629
rect 24008 11595 24042 11629
rect 24076 11595 24110 11629
rect 24144 11595 24178 11629
rect 24212 11595 24246 11629
rect 24280 11595 24314 11629
rect 24348 11595 24382 11629
rect 24416 11595 24450 11629
rect 24484 11595 24518 11629
rect 24552 11595 24586 11629
rect 24620 11595 24654 11629
rect 24688 11595 24722 11629
rect 24756 11595 24790 11629
rect 24824 11595 24858 11629
rect 24892 11595 24926 11629
rect 24960 11595 24994 11629
rect 25028 11595 25062 11629
rect 25096 11595 25130 11629
rect 25164 11595 25198 11629
rect 25232 11595 25266 11629
rect 25300 11595 25334 11629
rect 25368 11595 25402 11629
rect 25436 11595 25470 11629
rect 25504 11595 25528 11629
rect 19659 11588 25528 11595
rect 10304 11584 25528 11588
rect 6746 11577 25528 11584
rect 6746 11546 10404 11577
rect 6746 11512 6770 11546
rect 6804 11512 6839 11546
rect 6873 11512 6908 11546
rect 6942 11512 6977 11546
rect 7011 11512 7046 11546
rect 7080 11512 7115 11546
rect 7149 11512 7184 11546
rect 7218 11512 7253 11546
rect 7287 11512 7322 11546
rect 7356 11512 7391 11546
rect 7425 11512 7460 11546
rect 7494 11512 7529 11546
rect 7563 11512 7598 11546
rect 7632 11512 7667 11546
rect 7701 11512 7736 11546
rect 7770 11512 7805 11546
rect 7839 11512 7874 11546
rect 7908 11512 7943 11546
rect 7977 11512 8012 11546
rect 8046 11512 8081 11546
rect 8115 11512 8150 11546
rect 8184 11512 8219 11546
rect 8253 11512 8288 11546
rect 8322 11512 8357 11546
rect 8391 11512 8426 11546
rect 8460 11512 8495 11546
rect 8529 11512 8564 11546
rect 8598 11512 8633 11546
rect 8667 11512 8702 11546
rect 8736 11512 8771 11546
rect 8805 11512 8840 11546
rect 8874 11512 8909 11546
rect 8943 11512 8978 11546
rect 9012 11512 9046 11546
rect 9080 11512 9114 11546
rect 9148 11512 9182 11546
rect 9216 11512 9250 11546
rect 9284 11512 9318 11546
rect 9352 11512 9386 11546
rect 9420 11512 9454 11546
rect 9488 11512 9522 11546
rect 9556 11512 9590 11546
rect 9624 11512 9658 11546
rect 9692 11512 9726 11546
rect 9760 11512 9794 11546
rect 9828 11512 9862 11546
rect 9896 11512 9930 11546
rect 9964 11512 9998 11546
rect 10032 11512 10066 11546
rect 10100 11512 10134 11546
rect 10168 11512 10202 11546
rect 10236 11512 10270 11546
rect 10304 11543 10404 11546
rect 10438 11543 10473 11577
rect 10507 11543 10542 11577
rect 10576 11543 10611 11577
rect 10645 11543 10680 11577
rect 10714 11543 10749 11577
rect 10783 11543 10818 11577
rect 10852 11543 10887 11577
rect 10921 11543 10956 11577
rect 10990 11543 11025 11577
rect 11059 11543 11094 11577
rect 11128 11543 11163 11577
rect 11197 11543 11232 11577
rect 11266 11543 11301 11577
rect 11335 11543 11370 11577
rect 11404 11543 11439 11577
rect 11473 11543 11508 11577
rect 11542 11543 11577 11577
rect 11611 11543 11646 11577
rect 11680 11543 11715 11577
rect 11749 11543 11784 11577
rect 11818 11543 11853 11577
rect 11887 11543 11922 11577
rect 11956 11543 11991 11577
rect 12025 11543 12060 11577
rect 12094 11543 12129 11577
rect 12163 11543 12198 11577
rect 12232 11543 12267 11577
rect 12301 11543 12336 11577
rect 12370 11543 12405 11577
rect 12439 11543 12474 11577
rect 12508 11543 12543 11577
rect 12577 11543 12612 11577
rect 12646 11543 12681 11577
rect 12715 11543 12750 11577
rect 12784 11543 12819 11577
rect 12853 11543 12888 11577
rect 12922 11543 12957 11577
rect 12991 11543 13026 11577
rect 13060 11543 13095 11577
rect 13129 11543 13164 11577
rect 13198 11543 13233 11577
rect 13267 11543 13302 11577
rect 13336 11543 13371 11577
rect 10304 11512 13371 11543
rect 6746 11509 13371 11512
rect 6746 11475 10404 11509
rect 10438 11475 10473 11509
rect 10507 11475 10542 11509
rect 10576 11475 10611 11509
rect 10645 11475 10680 11509
rect 10714 11475 10749 11509
rect 10783 11475 10818 11509
rect 10852 11475 10887 11509
rect 10921 11475 10956 11509
rect 10990 11475 11025 11509
rect 11059 11475 11094 11509
rect 11128 11475 11163 11509
rect 11197 11475 11232 11509
rect 11266 11475 11301 11509
rect 11335 11475 11370 11509
rect 11404 11475 11439 11509
rect 11473 11475 11508 11509
rect 11542 11475 11577 11509
rect 11611 11475 11646 11509
rect 11680 11475 11715 11509
rect 11749 11475 11784 11509
rect 11818 11475 11853 11509
rect 11887 11475 11922 11509
rect 11956 11475 11991 11509
rect 12025 11475 12060 11509
rect 12094 11475 12129 11509
rect 12163 11475 12198 11509
rect 12232 11475 12267 11509
rect 12301 11475 12336 11509
rect 12370 11475 12405 11509
rect 12439 11475 12474 11509
rect 12508 11475 12543 11509
rect 12577 11475 12612 11509
rect 12646 11475 12681 11509
rect 12715 11475 12750 11509
rect 12784 11475 12819 11509
rect 12853 11475 12888 11509
rect 12922 11475 12957 11509
rect 12991 11475 13026 11509
rect 13060 11475 13095 11509
rect 13129 11475 13164 11509
rect 13198 11475 13233 11509
rect 13267 11475 13302 11509
rect 13336 11475 13371 11509
rect 6746 11474 13371 11475
rect 6746 11440 6770 11474
rect 6804 11440 6839 11474
rect 6873 11440 6908 11474
rect 6942 11440 6977 11474
rect 7011 11440 7046 11474
rect 7080 11440 7115 11474
rect 7149 11440 7184 11474
rect 7218 11440 7253 11474
rect 7287 11440 7322 11474
rect 7356 11440 7391 11474
rect 7425 11440 7460 11474
rect 7494 11440 7529 11474
rect 7563 11440 7598 11474
rect 7632 11440 7667 11474
rect 7701 11440 7736 11474
rect 7770 11440 7805 11474
rect 7839 11440 7874 11474
rect 7908 11440 7943 11474
rect 7977 11440 8012 11474
rect 8046 11440 8081 11474
rect 8115 11440 8150 11474
rect 8184 11440 8219 11474
rect 8253 11440 8288 11474
rect 8322 11440 8357 11474
rect 8391 11440 8426 11474
rect 8460 11440 8495 11474
rect 8529 11440 8564 11474
rect 8598 11440 8633 11474
rect 8667 11440 8702 11474
rect 8736 11440 8771 11474
rect 8805 11440 8840 11474
rect 8874 11440 8909 11474
rect 8943 11440 8978 11474
rect 9012 11440 9046 11474
rect 9080 11440 9114 11474
rect 9148 11440 9182 11474
rect 9216 11440 9250 11474
rect 9284 11440 9318 11474
rect 9352 11440 9386 11474
rect 9420 11440 9454 11474
rect 9488 11440 9522 11474
rect 9556 11440 9590 11474
rect 9624 11440 9658 11474
rect 9692 11440 9726 11474
rect 9760 11440 9794 11474
rect 9828 11440 9862 11474
rect 9896 11440 9930 11474
rect 9964 11440 9998 11474
rect 10032 11440 10066 11474
rect 10100 11440 10134 11474
rect 10168 11440 10202 11474
rect 10236 11440 10270 11474
rect 10304 11441 13371 11474
rect 10304 11440 10404 11441
rect 6746 11407 10404 11440
rect 10438 11407 10473 11441
rect 10507 11407 10542 11441
rect 10576 11407 10611 11441
rect 10645 11407 10680 11441
rect 10714 11407 10749 11441
rect 10783 11407 10818 11441
rect 10852 11407 10887 11441
rect 10921 11407 10956 11441
rect 10990 11407 11025 11441
rect 11059 11407 11094 11441
rect 11128 11407 11163 11441
rect 11197 11407 11232 11441
rect 11266 11407 11301 11441
rect 11335 11407 11370 11441
rect 11404 11407 11439 11441
rect 11473 11407 11508 11441
rect 11542 11407 11577 11441
rect 11611 11407 11646 11441
rect 11680 11407 11715 11441
rect 11749 11407 11784 11441
rect 11818 11407 11853 11441
rect 11887 11407 11922 11441
rect 11956 11407 11991 11441
rect 12025 11407 12060 11441
rect 12094 11407 12129 11441
rect 12163 11407 12198 11441
rect 12232 11407 12267 11441
rect 12301 11407 12336 11441
rect 12370 11407 12405 11441
rect 12439 11407 12474 11441
rect 12508 11407 12543 11441
rect 12577 11407 12612 11441
rect 12646 11407 12681 11441
rect 12715 11407 12750 11441
rect 12784 11407 12819 11441
rect 12853 11407 12888 11441
rect 12922 11407 12957 11441
rect 12991 11407 13026 11441
rect 13060 11407 13095 11441
rect 13129 11407 13164 11441
rect 13198 11407 13233 11441
rect 13267 11407 13302 11441
rect 13336 11407 13371 11441
rect 16261 11554 25528 11577
rect 16261 11520 16309 11554
rect 16343 11520 16379 11554
rect 16413 11520 16449 11554
rect 16483 11520 16519 11554
rect 16553 11520 16589 11554
rect 16623 11520 16658 11554
rect 16692 11520 16727 11554
rect 16761 11520 16796 11554
rect 16830 11520 16865 11554
rect 16899 11520 16934 11554
rect 16968 11520 17003 11554
rect 17037 11520 17072 11554
rect 17106 11520 17141 11554
rect 17175 11520 17210 11554
rect 17244 11520 17279 11554
rect 17313 11520 17348 11554
rect 17382 11520 17417 11554
rect 17451 11520 17486 11554
rect 17520 11520 17555 11554
rect 17589 11520 17624 11554
rect 17658 11520 17693 11554
rect 17727 11520 17762 11554
rect 17796 11520 17831 11554
rect 17865 11520 17900 11554
rect 17934 11520 17969 11554
rect 18003 11520 18038 11554
rect 18072 11520 18107 11554
rect 18141 11520 18176 11554
rect 18210 11520 18245 11554
rect 18279 11520 18314 11554
rect 18348 11520 18383 11554
rect 18417 11520 18452 11554
rect 18486 11520 18521 11554
rect 18555 11520 18590 11554
rect 18624 11520 18659 11554
rect 18693 11520 18728 11554
rect 18762 11520 18797 11554
rect 18831 11520 18866 11554
rect 18900 11520 18935 11554
rect 18969 11520 19004 11554
rect 19038 11520 19073 11554
rect 19107 11520 19142 11554
rect 19176 11520 19211 11554
rect 19245 11520 19280 11554
rect 19314 11520 19349 11554
rect 19383 11520 19418 11554
rect 19452 11520 19487 11554
rect 19521 11520 19556 11554
rect 19590 11520 19625 11554
rect 19659 11527 25528 11554
rect 19659 11520 19683 11527
rect 16261 11486 19683 11520
rect 16261 11452 16309 11486
rect 16343 11452 16379 11486
rect 16413 11452 16449 11486
rect 16483 11452 16519 11486
rect 16553 11452 16589 11486
rect 16623 11452 16658 11486
rect 16692 11452 16727 11486
rect 16761 11452 16796 11486
rect 16830 11452 16865 11486
rect 16899 11452 16934 11486
rect 16968 11452 17003 11486
rect 17037 11452 17072 11486
rect 17106 11452 17141 11486
rect 17175 11452 17210 11486
rect 17244 11452 17279 11486
rect 17313 11452 17348 11486
rect 17382 11452 17417 11486
rect 17451 11452 17486 11486
rect 17520 11452 17555 11486
rect 17589 11452 17624 11486
rect 17658 11452 17693 11486
rect 17727 11452 17762 11486
rect 17796 11452 17831 11486
rect 17865 11452 17900 11486
rect 17934 11452 17969 11486
rect 18003 11452 18038 11486
rect 18072 11452 18107 11486
rect 18141 11452 18176 11486
rect 18210 11452 18245 11486
rect 18279 11452 18314 11486
rect 18348 11452 18383 11486
rect 18417 11452 18452 11486
rect 18486 11452 18521 11486
rect 18555 11452 18590 11486
rect 18624 11452 18659 11486
rect 18693 11452 18728 11486
rect 18762 11452 18797 11486
rect 18831 11452 18866 11486
rect 18900 11452 18935 11486
rect 18969 11452 19004 11486
rect 19038 11452 19073 11486
rect 19107 11452 19142 11486
rect 19176 11452 19211 11486
rect 19245 11452 19280 11486
rect 19314 11452 19349 11486
rect 19383 11452 19418 11486
rect 19452 11452 19487 11486
rect 19521 11452 19556 11486
rect 19590 11452 19625 11486
rect 19659 11452 19683 11486
rect 16261 11418 19683 11452
rect 16261 11407 16309 11418
rect 6746 11402 16309 11407
rect 6746 11368 6770 11402
rect 6804 11368 6839 11402
rect 6873 11368 6908 11402
rect 6942 11368 6977 11402
rect 7011 11368 7046 11402
rect 7080 11368 7115 11402
rect 7149 11368 7184 11402
rect 7218 11368 7253 11402
rect 7287 11368 7322 11402
rect 7356 11368 7391 11402
rect 7425 11368 7460 11402
rect 7494 11368 7529 11402
rect 7563 11368 7598 11402
rect 7632 11368 7667 11402
rect 7701 11368 7736 11402
rect 7770 11368 7805 11402
rect 7839 11368 7874 11402
rect 7908 11368 7943 11402
rect 7977 11368 8012 11402
rect 8046 11368 8081 11402
rect 8115 11368 8150 11402
rect 8184 11368 8219 11402
rect 8253 11368 8288 11402
rect 8322 11368 8357 11402
rect 8391 11368 8426 11402
rect 8460 11368 8495 11402
rect 8529 11368 8564 11402
rect 8598 11368 8633 11402
rect 8667 11368 8702 11402
rect 8736 11368 8771 11402
rect 8805 11368 8840 11402
rect 8874 11368 8909 11402
rect 8943 11368 8978 11402
rect 9012 11368 9046 11402
rect 9080 11368 9114 11402
rect 9148 11368 9182 11402
rect 9216 11368 9250 11402
rect 9284 11368 9318 11402
rect 9352 11368 9386 11402
rect 9420 11368 9454 11402
rect 9488 11368 9522 11402
rect 9556 11368 9590 11402
rect 9624 11368 9658 11402
rect 9692 11368 9726 11402
rect 9760 11368 9794 11402
rect 9828 11368 9862 11402
rect 9896 11368 9930 11402
rect 9964 11368 9998 11402
rect 10032 11368 10066 11402
rect 10100 11368 10134 11402
rect 10168 11368 10202 11402
rect 10236 11368 10270 11402
rect 10304 11384 16309 11402
rect 16343 11384 16379 11418
rect 16413 11384 16449 11418
rect 16483 11384 16519 11418
rect 16553 11384 16589 11418
rect 16623 11384 16658 11418
rect 16692 11384 16727 11418
rect 16761 11384 16796 11418
rect 16830 11384 16865 11418
rect 16899 11384 16934 11418
rect 16968 11384 17003 11418
rect 17037 11384 17072 11418
rect 17106 11384 17141 11418
rect 17175 11384 17210 11418
rect 17244 11384 17279 11418
rect 17313 11384 17348 11418
rect 17382 11384 17417 11418
rect 17451 11384 17486 11418
rect 17520 11384 17555 11418
rect 17589 11384 17624 11418
rect 17658 11384 17693 11418
rect 17727 11384 17762 11418
rect 17796 11384 17831 11418
rect 17865 11384 17900 11418
rect 17934 11384 17969 11418
rect 18003 11384 18038 11418
rect 18072 11384 18107 11418
rect 18141 11384 18176 11418
rect 18210 11384 18245 11418
rect 18279 11384 18314 11418
rect 18348 11384 18383 11418
rect 18417 11384 18452 11418
rect 18486 11384 18521 11418
rect 18555 11384 18590 11418
rect 18624 11384 18659 11418
rect 18693 11384 18728 11418
rect 18762 11384 18797 11418
rect 18831 11384 18866 11418
rect 18900 11384 18935 11418
rect 18969 11384 19004 11418
rect 19038 11384 19073 11418
rect 19107 11384 19142 11418
rect 19176 11384 19211 11418
rect 19245 11384 19280 11418
rect 19314 11384 19349 11418
rect 19383 11384 19418 11418
rect 19452 11384 19487 11418
rect 19521 11384 19556 11418
rect 19590 11384 19625 11418
rect 19659 11384 19683 11418
rect 10304 11368 19382 11384
rect 6746 11350 19382 11368
rect 25101 11355 25528 11527
rect 6746 11346 16319 11350
rect 6746 11330 10328 11346
rect 6746 11296 6770 11330
rect 6804 11296 6839 11330
rect 6873 11296 6908 11330
rect 6942 11296 6977 11330
rect 7011 11296 7046 11330
rect 7080 11296 7115 11330
rect 7149 11296 7184 11330
rect 7218 11296 7253 11330
rect 7287 11296 7322 11330
rect 7356 11296 7391 11330
rect 7425 11296 7460 11330
rect 7494 11296 7529 11330
rect 7563 11296 7598 11330
rect 7632 11296 7667 11330
rect 7701 11296 7736 11330
rect 7770 11296 7805 11330
rect 7839 11296 7874 11330
rect 7908 11296 7943 11330
rect 7977 11296 8012 11330
rect 8046 11296 8081 11330
rect 8115 11296 8150 11330
rect 8184 11296 8219 11330
rect 8253 11296 8288 11330
rect 8322 11296 8357 11330
rect 8391 11296 8426 11330
rect 8460 11296 8495 11330
rect 8529 11296 8564 11330
rect 8598 11296 8633 11330
rect 8667 11296 8702 11330
rect 8736 11296 8771 11330
rect 8805 11296 8840 11330
rect 8874 11296 8909 11330
rect 8943 11296 8978 11330
rect 9012 11296 9046 11330
rect 9080 11296 9114 11330
rect 9148 11296 9182 11330
rect 9216 11296 9250 11330
rect 9284 11296 9318 11330
rect 9352 11296 9386 11330
rect 9420 11296 9454 11330
rect 9488 11296 9522 11330
rect 9556 11296 9590 11330
rect 9624 11296 9658 11330
rect 9692 11296 9726 11330
rect 9760 11296 9794 11330
rect 9828 11296 9862 11330
rect 9896 11296 9930 11330
rect 9964 11296 9998 11330
rect 10032 11296 10066 11330
rect 10100 11296 10134 11330
rect 10168 11296 10202 11330
rect 10236 11296 10270 11330
rect 10304 11296 10328 11330
rect 14066 11316 16319 11346
rect 16353 11316 16388 11350
rect 16422 11316 16457 11350
rect 16491 11316 16526 11350
rect 16560 11316 16594 11350
rect 16628 11316 16662 11350
rect 16696 11316 16730 11350
rect 16764 11316 16798 11350
rect 16832 11316 16866 11350
rect 16900 11316 16934 11350
rect 16968 11316 17002 11350
rect 17036 11316 17070 11350
rect 17104 11316 17138 11350
rect 17172 11316 17206 11350
rect 17240 11316 17274 11350
rect 17308 11316 17342 11350
rect 17376 11316 17410 11350
rect 17444 11316 17478 11350
rect 17512 11316 17546 11350
rect 17580 11316 17614 11350
rect 17648 11316 17682 11350
rect 17716 11316 17750 11350
rect 17784 11316 17818 11350
rect 17852 11316 17886 11350
rect 17920 11316 17954 11350
rect 17988 11316 18022 11350
rect 18056 11316 18090 11350
rect 18124 11316 18158 11350
rect 18192 11316 18226 11350
rect 18260 11316 18294 11350
rect 18328 11316 18362 11350
rect 18396 11316 18430 11350
rect 18464 11316 18498 11350
rect 18532 11316 18566 11350
rect 18600 11316 18634 11350
rect 18668 11316 18702 11350
rect 18736 11316 18770 11350
rect 18804 11316 18838 11350
rect 18872 11316 18906 11350
rect 18940 11316 18974 11350
rect 19008 11316 19042 11350
rect 19076 11316 19110 11350
rect 19144 11316 19178 11350
rect 19212 11316 19246 11350
rect 19280 11316 19314 11350
rect 19348 11316 19382 11350
rect 6746 11258 10328 11296
rect 6746 11224 6770 11258
rect 6804 11224 6839 11258
rect 6873 11224 6908 11258
rect 6942 11224 6977 11258
rect 7011 11224 7046 11258
rect 7080 11224 7115 11258
rect 7149 11224 7184 11258
rect 7218 11224 7253 11258
rect 7287 11224 7322 11258
rect 7356 11224 7391 11258
rect 7425 11224 7460 11258
rect 7494 11224 7529 11258
rect 7563 11224 7598 11258
rect 7632 11224 7667 11258
rect 7701 11224 7736 11258
rect 7770 11224 7805 11258
rect 7839 11224 7874 11258
rect 7908 11224 7943 11258
rect 7977 11224 8012 11258
rect 8046 11224 8081 11258
rect 8115 11224 8150 11258
rect 8184 11224 8219 11258
rect 8253 11224 8288 11258
rect 8322 11224 8357 11258
rect 8391 11224 8426 11258
rect 8460 11224 8495 11258
rect 8529 11224 8564 11258
rect 8598 11224 8633 11258
rect 8667 11224 8702 11258
rect 8736 11224 8771 11258
rect 8805 11224 8840 11258
rect 8874 11224 8909 11258
rect 8943 11224 8978 11258
rect 9012 11224 9046 11258
rect 9080 11224 9114 11258
rect 9148 11224 9182 11258
rect 9216 11224 9250 11258
rect 9284 11224 9318 11258
rect 9352 11224 9386 11258
rect 9420 11224 9454 11258
rect 9488 11224 9522 11258
rect 9556 11224 9590 11258
rect 9624 11224 9658 11258
rect 9692 11224 9726 11258
rect 9760 11224 9794 11258
rect 9828 11224 9862 11258
rect 9896 11224 9930 11258
rect 9964 11224 9998 11258
rect 10032 11224 10066 11258
rect 10100 11224 10134 11258
rect 10168 11224 10202 11258
rect 10236 11224 10270 11258
rect 10304 11224 10328 11258
rect 6746 11186 10328 11224
rect 6746 11152 6770 11186
rect 6804 11152 6839 11186
rect 6873 11152 6908 11186
rect 6942 11152 6977 11186
rect 7011 11152 7046 11186
rect 7080 11152 7115 11186
rect 7149 11152 7184 11186
rect 7218 11152 7253 11186
rect 7287 11152 7322 11186
rect 7356 11152 7391 11186
rect 7425 11152 7460 11186
rect 7494 11152 7529 11186
rect 7563 11152 7598 11186
rect 7632 11152 7667 11186
rect 7701 11152 7736 11186
rect 7770 11152 7805 11186
rect 7839 11152 7874 11186
rect 7908 11152 7943 11186
rect 7977 11152 8012 11186
rect 8046 11152 8081 11186
rect 8115 11152 8150 11186
rect 8184 11152 8219 11186
rect 8253 11152 8288 11186
rect 8322 11152 8357 11186
rect 8391 11152 8426 11186
rect 8460 11152 8495 11186
rect 8529 11152 8564 11186
rect 8598 11152 8633 11186
rect 8667 11152 8702 11186
rect 8736 11152 8771 11186
rect 8805 11152 8840 11186
rect 8874 11152 8909 11186
rect 8943 11152 8978 11186
rect 9012 11152 9046 11186
rect 9080 11152 9114 11186
rect 9148 11152 9182 11186
rect 9216 11152 9250 11186
rect 9284 11152 9318 11186
rect 9352 11152 9386 11186
rect 9420 11152 9454 11186
rect 9488 11152 9522 11186
rect 9556 11152 9590 11186
rect 9624 11152 9658 11186
rect 9692 11152 9726 11186
rect 9760 11152 9794 11186
rect 9828 11152 9862 11186
rect 9896 11152 9930 11186
rect 9964 11152 9998 11186
rect 10032 11152 10066 11186
rect 10100 11152 10134 11186
rect 10168 11152 10202 11186
rect 10236 11152 10270 11186
rect 10304 11152 10328 11186
rect 6746 11148 10328 11152
rect 16285 11278 19382 11316
rect 16285 11244 16319 11278
rect 16353 11244 16388 11278
rect 16422 11244 16457 11278
rect 16491 11244 16526 11278
rect 16560 11244 16594 11278
rect 16628 11244 16662 11278
rect 16696 11244 16730 11278
rect 16764 11244 16798 11278
rect 16832 11244 16866 11278
rect 16900 11244 16934 11278
rect 16968 11244 17002 11278
rect 17036 11244 17070 11278
rect 17104 11244 17138 11278
rect 17172 11244 17206 11278
rect 17240 11244 17274 11278
rect 17308 11244 17342 11278
rect 17376 11244 17410 11278
rect 17444 11244 17478 11278
rect 17512 11244 17546 11278
rect 17580 11244 17614 11278
rect 17648 11244 17682 11278
rect 17716 11244 17750 11278
rect 17784 11244 17818 11278
rect 17852 11244 17886 11278
rect 17920 11244 17954 11278
rect 17988 11244 18022 11278
rect 18056 11244 18090 11278
rect 18124 11244 18158 11278
rect 18192 11244 18226 11278
rect 18260 11244 18294 11278
rect 18328 11244 18362 11278
rect 18396 11244 18430 11278
rect 18464 11244 18498 11278
rect 18532 11244 18566 11278
rect 18600 11244 18634 11278
rect 18668 11244 18702 11278
rect 18736 11244 18770 11278
rect 18804 11244 18838 11278
rect 18872 11244 18906 11278
rect 18940 11244 18974 11278
rect 19008 11244 19042 11278
rect 19076 11244 19110 11278
rect 19144 11244 19178 11278
rect 19212 11244 19246 11278
rect 19280 11244 19314 11278
rect 19348 11244 19382 11278
rect 25100 11321 25124 11355
rect 25158 11321 25196 11355
rect 25230 11321 25268 11355
rect 25302 11321 25340 11355
rect 25374 11321 25412 11355
rect 25446 11321 25484 11355
rect 25518 11321 25556 11355
rect 25590 11321 25627 11355
rect 25661 11321 25698 11355
rect 25732 11321 25769 11355
rect 25803 11321 25840 11355
rect 25874 11321 25911 11355
rect 25945 11321 25982 11355
rect 26016 11321 26053 11355
rect 26087 11321 26124 11355
rect 26158 11321 26195 11355
rect 26229 11321 26283 11355
rect 25100 11287 26283 11321
rect 25100 11253 25124 11287
rect 25158 11253 25196 11287
rect 25230 11253 25268 11287
rect 25302 11253 25340 11287
rect 25374 11253 25412 11287
rect 25446 11253 25484 11287
rect 25518 11253 25556 11287
rect 25590 11253 25627 11287
rect 25661 11253 25698 11287
rect 25732 11253 25769 11287
rect 25803 11253 25840 11287
rect 25874 11253 25911 11287
rect 25945 11253 25982 11287
rect 26016 11253 26053 11287
rect 26087 11253 26124 11287
rect 26158 11253 26195 11287
rect 26229 11253 26283 11287
rect 16285 11206 19382 11244
rect 16285 11172 16319 11206
rect 16353 11172 16388 11206
rect 16422 11172 16457 11206
rect 16491 11172 16526 11206
rect 16560 11172 16594 11206
rect 16628 11172 16662 11206
rect 16696 11172 16730 11206
rect 16764 11172 16798 11206
rect 16832 11172 16866 11206
rect 16900 11172 16934 11206
rect 16968 11172 17002 11206
rect 17036 11172 17070 11206
rect 17104 11172 17138 11206
rect 17172 11172 17206 11206
rect 17240 11172 17274 11206
rect 17308 11172 17342 11206
rect 17376 11172 17410 11206
rect 17444 11172 17478 11206
rect 17512 11172 17546 11206
rect 17580 11172 17614 11206
rect 17648 11172 17682 11206
rect 17716 11172 17750 11206
rect 17784 11172 17818 11206
rect 17852 11172 17886 11206
rect 17920 11172 17954 11206
rect 17988 11172 18022 11206
rect 18056 11172 18090 11206
rect 18124 11172 18158 11206
rect 18192 11172 18226 11206
rect 18260 11172 18294 11206
rect 18328 11172 18362 11206
rect 18396 11172 18430 11206
rect 18464 11172 18498 11206
rect 18532 11172 18566 11206
rect 18600 11172 18634 11206
rect 18668 11172 18702 11206
rect 18736 11172 18770 11206
rect 18804 11172 18838 11206
rect 18872 11172 18906 11206
rect 18940 11172 18974 11206
rect 19008 11172 19042 11206
rect 19076 11172 19110 11206
rect 19144 11172 19178 11206
rect 19212 11172 19246 11206
rect 19280 11172 19314 11206
rect 19348 11172 19382 11206
rect 6746 11072 7246 11148
rect 6746 11038 6751 11072
rect 6785 11038 6827 11072
rect 6861 11038 6903 11072
rect 6937 11038 6979 11072
rect 7013 11038 7055 11072
rect 7089 11038 7131 11072
rect 7165 11038 7207 11072
rect 7241 11038 7246 11072
rect 6746 11004 7246 11038
rect 6746 10970 6751 11004
rect 6785 10970 6827 11004
rect 6861 10970 6903 11004
rect 6937 10970 6979 11004
rect 7013 10970 7055 11004
rect 7089 10970 7131 11004
rect 7165 10970 7207 11004
rect 7241 10970 7246 11004
rect 6746 10936 7246 10970
rect 6746 10902 6751 10936
rect 6785 10902 6827 10936
rect 6861 10902 6903 10936
rect 6937 10902 6979 10936
rect 7013 10902 7055 10936
rect 7089 10902 7131 10936
rect 7165 10902 7207 10936
rect 7241 10902 7246 10936
rect 6746 10868 7246 10902
rect 6746 10834 6751 10868
rect 6785 10834 6827 10868
rect 6861 10834 6903 10868
rect 6937 10834 6979 10868
rect 7013 10834 7055 10868
rect 7089 10834 7131 10868
rect 7165 10834 7207 10868
rect 7241 10834 7246 10868
rect 6746 10800 7246 10834
rect 6746 10766 6751 10800
rect 6785 10766 6827 10800
rect 6861 10766 6903 10800
rect 6937 10766 6979 10800
rect 7013 10766 7055 10800
rect 7089 10766 7131 10800
rect 7165 10766 7207 10800
rect 7241 10766 7246 10800
rect 6746 10732 7246 10766
rect 6746 10698 6751 10732
rect 6785 10698 6827 10732
rect 6861 10698 6903 10732
rect 6937 10698 6979 10732
rect 7013 10698 7055 10732
rect 7089 10698 7131 10732
rect 7165 10698 7207 10732
rect 7241 10698 7246 10732
rect 6746 10664 7246 10698
rect 6746 10630 6751 10664
rect 6785 10630 6827 10664
rect 6861 10630 6903 10664
rect 6937 10630 6979 10664
rect 7013 10630 7055 10664
rect 7089 10630 7131 10664
rect 7165 10630 7207 10664
rect 7241 10630 7246 10664
rect 6746 10596 7246 10630
rect 6746 10562 6751 10596
rect 6785 10562 6827 10596
rect 6861 10562 6903 10596
rect 6937 10562 6979 10596
rect 7013 10562 7055 10596
rect 7089 10562 7131 10596
rect 7165 10562 7207 10596
rect 7241 10562 7246 10596
rect 6746 10528 7246 10562
rect 6746 10494 6751 10528
rect 6785 10494 6827 10528
rect 6861 10494 6903 10528
rect 6937 10494 6979 10528
rect 7013 10494 7055 10528
rect 7089 10494 7131 10528
rect 7165 10494 7207 10528
rect 7241 10494 7246 10528
rect 6746 10460 7246 10494
rect 6746 10426 6751 10460
rect 6785 10426 6827 10460
rect 6861 10426 6903 10460
rect 6937 10426 6979 10460
rect 7013 10426 7055 10460
rect 7089 10426 7131 10460
rect 7165 10426 7207 10460
rect 7241 10426 7246 10460
rect 6746 10392 7246 10426
rect 6746 10358 6751 10392
rect 6785 10358 6827 10392
rect 6861 10358 6903 10392
rect 6937 10358 6979 10392
rect 7013 10358 7055 10392
rect 7089 10358 7131 10392
rect 7165 10358 7207 10392
rect 7241 10358 7246 10392
rect 6746 10324 7246 10358
rect 6746 10290 6751 10324
rect 6785 10290 6827 10324
rect 6861 10290 6903 10324
rect 6937 10290 6979 10324
rect 7013 10290 7055 10324
rect 7089 10290 7131 10324
rect 7165 10290 7207 10324
rect 7241 10290 7246 10324
rect 6746 10256 7246 10290
rect 6746 10222 6751 10256
rect 6785 10222 6827 10256
rect 6861 10222 6903 10256
rect 6937 10222 6979 10256
rect 7013 10222 7055 10256
rect 7089 10222 7131 10256
rect 7165 10222 7207 10256
rect 7241 10222 7246 10256
rect 6746 10188 7246 10222
rect 6746 10154 6751 10188
rect 6785 10154 6827 10188
rect 6861 10154 6903 10188
rect 6937 10154 6979 10188
rect 7013 10154 7055 10188
rect 7089 10154 7131 10188
rect 7165 10154 7207 10188
rect 7241 10154 7246 10188
rect 6746 10120 7246 10154
rect 6746 10086 6751 10120
rect 6785 10086 6827 10120
rect 6861 10086 6903 10120
rect 6937 10086 6979 10120
rect 7013 10086 7055 10120
rect 7089 10086 7131 10120
rect 7165 10086 7207 10120
rect 7241 10086 7246 10120
rect 6746 10052 7246 10086
rect 6746 10018 6751 10052
rect 6785 10018 6827 10052
rect 6861 10018 6903 10052
rect 6937 10018 6979 10052
rect 7013 10018 7055 10052
rect 7089 10018 7131 10052
rect 7165 10018 7207 10052
rect 7241 10018 7246 10052
rect 6746 9984 7246 10018
rect 6746 9950 6751 9984
rect 6785 9950 6827 9984
rect 6861 9950 6903 9984
rect 6937 9950 6979 9984
rect 7013 9950 7055 9984
rect 7089 9950 7131 9984
rect 7165 9950 7207 9984
rect 7241 9950 7246 9984
rect 6746 9916 7246 9950
rect 6746 9882 6751 9916
rect 6785 9882 6827 9916
rect 6861 9882 6903 9916
rect 6937 9882 6979 9916
rect 7013 9882 7055 9916
rect 7089 9882 7131 9916
rect 7165 9882 7207 9916
rect 7241 9882 7246 9916
rect 6746 9848 7246 9882
rect 6746 9814 6751 9848
rect 6785 9814 6827 9848
rect 6861 9814 6903 9848
rect 6937 9814 6979 9848
rect 7013 9814 7055 9848
rect 7089 9814 7131 9848
rect 7165 9814 7207 9848
rect 7241 9814 7246 9848
rect 6746 9780 7246 9814
rect 6746 9746 6751 9780
rect 6785 9746 6827 9780
rect 6861 9746 6903 9780
rect 6937 9746 6979 9780
rect 7013 9746 7055 9780
rect 7089 9746 7131 9780
rect 7165 9746 7207 9780
rect 7241 9746 7246 9780
rect 6746 9712 7246 9746
rect 6746 9678 6751 9712
rect 6785 9678 6827 9712
rect 6861 9678 6903 9712
rect 6937 9678 6979 9712
rect 7013 9678 7055 9712
rect 7089 9678 7131 9712
rect 7165 9678 7207 9712
rect 7241 9678 7246 9712
rect 6746 9644 7246 9678
rect 6746 9610 6751 9644
rect 6785 9610 6827 9644
rect 6861 9610 6903 9644
rect 6937 9610 6979 9644
rect 7013 9610 7055 9644
rect 7089 9610 7131 9644
rect 7165 9610 7207 9644
rect 7241 9610 7246 9644
rect 6746 9589 7246 9610
rect 10049 11072 10219 11148
rect 16285 11134 19382 11172
rect 16285 11100 16319 11134
rect 16353 11100 16388 11134
rect 16422 11100 16457 11134
rect 16491 11100 16526 11134
rect 16560 11100 16594 11134
rect 16628 11100 16662 11134
rect 16696 11100 16730 11134
rect 16764 11100 16798 11134
rect 16832 11100 16866 11134
rect 16900 11100 16934 11134
rect 16968 11100 17002 11134
rect 17036 11100 17070 11134
rect 17104 11100 17138 11134
rect 17172 11100 17206 11134
rect 17240 11100 17274 11134
rect 17308 11100 17342 11134
rect 17376 11100 17410 11134
rect 17444 11100 17478 11134
rect 17512 11100 17546 11134
rect 17580 11100 17614 11134
rect 17648 11100 17682 11134
rect 17716 11100 17750 11134
rect 17784 11100 17818 11134
rect 17852 11100 17886 11134
rect 17920 11100 17954 11134
rect 17988 11100 18022 11134
rect 18056 11100 18090 11134
rect 18124 11100 18158 11134
rect 18192 11100 18226 11134
rect 18260 11100 18294 11134
rect 18328 11100 18362 11134
rect 18396 11100 18430 11134
rect 18464 11100 18498 11134
rect 18532 11100 18566 11134
rect 18600 11100 18634 11134
rect 18668 11100 18702 11134
rect 18736 11100 18770 11134
rect 18804 11100 18838 11134
rect 18872 11100 18906 11134
rect 18940 11100 18974 11134
rect 19008 11100 19042 11134
rect 19076 11100 19110 11134
rect 19144 11100 19178 11134
rect 19212 11100 19246 11134
rect 19280 11100 19314 11134
rect 19348 11100 19382 11134
rect 16285 11076 19382 11100
rect 10049 10255 10219 10290
rect 10083 10221 10117 10255
rect 10151 10221 10185 10255
rect 10049 10186 10219 10221
rect 10083 10152 10117 10186
rect 10151 10152 10185 10186
rect 10049 10117 10219 10152
rect 10083 10083 10117 10117
rect 10151 10083 10185 10117
rect 10049 10048 10219 10083
rect 10083 10014 10117 10048
rect 10151 10014 10185 10048
rect 10049 9979 10219 10014
rect 10083 9945 10117 9979
rect 10151 9945 10185 9979
rect 10049 9910 10219 9945
rect 10083 9876 10117 9910
rect 10151 9876 10185 9910
rect 10049 9841 10219 9876
rect 10083 9807 10117 9841
rect 10151 9807 10185 9841
rect 10049 9772 10219 9807
rect 10083 9738 10117 9772
rect 10151 9738 10185 9772
rect 10049 9703 10219 9738
rect 10083 9669 10117 9703
rect 10151 9669 10185 9703
rect 10049 9634 10219 9669
rect 10083 9600 10117 9634
rect 10151 9600 10185 9634
rect 10049 9589 10219 9600
rect 6746 9588 10219 9589
rect 6746 9576 7332 9588
rect 6746 9542 6751 9576
rect 6785 9542 6827 9576
rect 6861 9542 6903 9576
rect 6937 9542 6979 9576
rect 7013 9542 7055 9576
rect 7089 9542 7131 9576
rect 7165 9542 7207 9576
rect 7241 9554 7332 9576
rect 7366 9554 7401 9588
rect 7435 9554 7470 9588
rect 7504 9554 7539 9588
rect 7573 9554 7608 9588
rect 7642 9554 7677 9588
rect 7711 9554 7746 9588
rect 7780 9554 7815 9588
rect 7849 9554 7884 9588
rect 7918 9554 7953 9588
rect 7987 9554 8022 9588
rect 8056 9554 8091 9588
rect 8125 9554 8160 9588
rect 8194 9554 8229 9588
rect 8263 9554 8297 9588
rect 8331 9554 8365 9588
rect 8399 9554 8433 9588
rect 8467 9554 8501 9588
rect 8535 9554 8569 9588
rect 8603 9554 8637 9588
rect 8671 9554 8705 9588
rect 8739 9554 8773 9588
rect 8807 9554 8841 9588
rect 8875 9554 8909 9588
rect 8943 9554 8977 9588
rect 9011 9554 9045 9588
rect 9079 9554 9113 9588
rect 9147 9554 9181 9588
rect 9215 9554 9249 9588
rect 9283 9554 9317 9588
rect 9351 9554 9385 9588
rect 9419 9554 9453 9588
rect 9487 9554 9521 9588
rect 9555 9554 9589 9588
rect 9623 9554 9657 9588
rect 9691 9554 9725 9588
rect 9759 9554 9793 9588
rect 9827 9554 9861 9588
rect 9895 9554 9929 9588
rect 9963 9565 10219 9588
rect 9963 9554 10049 9565
rect 7241 9542 10049 9554
rect 6746 9531 10049 9542
rect 10083 9531 10117 9565
rect 10151 9531 10185 9565
rect 26249 10370 26283 11253
rect 26249 10336 26277 10370
rect 26311 10336 26348 10370
rect 26382 10336 26419 10370
rect 26453 10336 26490 10370
rect 26524 10336 26561 10370
rect 26595 10336 26632 10370
rect 26666 10336 26703 10370
rect 26737 10336 26774 10370
rect 26808 10336 26845 10370
rect 26879 10336 26916 10370
rect 26950 10336 26986 10370
rect 27020 10336 27056 10370
rect 27090 10336 27126 10370
rect 27160 10336 27196 10370
rect 27230 10336 27266 10370
rect 27300 10336 27336 10370
rect 27370 10336 27406 10370
rect 27440 10346 27853 10370
rect 27440 10336 27547 10346
rect 26249 10312 27547 10336
rect 27581 10312 27615 10346
rect 27649 10312 27683 10346
rect 27717 10312 27751 10346
rect 27785 10312 27819 10346
rect 26249 10302 27853 10312
rect 26249 10268 26277 10302
rect 26311 10268 26348 10302
rect 26382 10268 26419 10302
rect 26453 10268 26490 10302
rect 26524 10268 26561 10302
rect 26595 10268 26632 10302
rect 26666 10268 26703 10302
rect 26737 10268 26774 10302
rect 26808 10268 26845 10302
rect 26879 10268 26916 10302
rect 26950 10268 26986 10302
rect 27020 10268 27056 10302
rect 27090 10268 27126 10302
rect 27160 10268 27196 10302
rect 27230 10268 27266 10302
rect 27300 10268 27336 10302
rect 27370 10268 27406 10302
rect 27440 10277 27853 10302
rect 27440 10268 27547 10277
rect 26249 10243 27547 10268
rect 27581 10243 27615 10277
rect 27649 10243 27683 10277
rect 27717 10243 27751 10277
rect 27785 10243 27819 10277
rect 26249 10234 27853 10243
rect 26249 10200 26277 10234
rect 26311 10200 26348 10234
rect 26382 10200 26419 10234
rect 26453 10200 26490 10234
rect 26524 10200 26561 10234
rect 26595 10200 26632 10234
rect 26666 10200 26703 10234
rect 26737 10200 26774 10234
rect 26808 10200 26845 10234
rect 26879 10200 26916 10234
rect 26950 10200 26986 10234
rect 27020 10200 27056 10234
rect 27090 10200 27126 10234
rect 27160 10200 27196 10234
rect 27230 10200 27266 10234
rect 27300 10200 27336 10234
rect 27370 10200 27406 10234
rect 27440 10208 27853 10234
rect 27440 10200 27547 10208
rect 26249 10174 27547 10200
rect 27581 10174 27615 10208
rect 27649 10174 27683 10208
rect 27717 10174 27751 10208
rect 27785 10174 27819 10208
rect 26249 10166 27853 10174
rect 26249 10132 26277 10166
rect 26311 10132 26348 10166
rect 26382 10132 26419 10166
rect 26453 10132 26490 10166
rect 26524 10132 26561 10166
rect 26595 10132 26632 10166
rect 26666 10132 26703 10166
rect 26737 10132 26774 10166
rect 26808 10132 26845 10166
rect 26879 10132 26916 10166
rect 26950 10132 26986 10166
rect 27020 10132 27056 10166
rect 27090 10132 27126 10166
rect 27160 10132 27196 10166
rect 27230 10132 27266 10166
rect 27300 10132 27336 10166
rect 27370 10132 27406 10166
rect 27440 10139 27853 10166
rect 27440 10132 27547 10139
rect 26249 10105 27547 10132
rect 27581 10105 27615 10139
rect 27649 10105 27683 10139
rect 27717 10105 27751 10139
rect 27785 10105 27819 10139
rect 26249 10098 27853 10105
rect 26249 10064 26277 10098
rect 26311 10064 26348 10098
rect 26382 10064 26419 10098
rect 26453 10064 26490 10098
rect 26524 10064 26561 10098
rect 26595 10064 26632 10098
rect 26666 10064 26703 10098
rect 26737 10064 26774 10098
rect 26808 10064 26845 10098
rect 26879 10064 26916 10098
rect 26950 10064 26986 10098
rect 27020 10064 27056 10098
rect 27090 10064 27126 10098
rect 27160 10064 27196 10098
rect 27230 10064 27266 10098
rect 27300 10064 27336 10098
rect 27370 10064 27406 10098
rect 27440 10070 27853 10098
rect 27440 10064 27547 10070
rect 26249 10036 27547 10064
rect 27581 10036 27615 10070
rect 27649 10036 27683 10070
rect 27717 10036 27751 10070
rect 27785 10036 27819 10070
rect 26249 10030 27853 10036
rect 26249 9996 26277 10030
rect 26311 9996 26348 10030
rect 26382 9996 26419 10030
rect 26453 9996 26490 10030
rect 26524 9996 26561 10030
rect 26595 9996 26632 10030
rect 26666 9996 26703 10030
rect 26737 9996 26774 10030
rect 26808 9996 26845 10030
rect 26879 9996 26916 10030
rect 26950 9996 26986 10030
rect 27020 9996 27056 10030
rect 27090 9996 27126 10030
rect 27160 9996 27196 10030
rect 27230 9996 27266 10030
rect 27300 9996 27336 10030
rect 27370 9996 27406 10030
rect 27440 10001 27853 10030
rect 27440 9996 27547 10001
rect 26249 9967 27547 9996
rect 27581 9967 27615 10001
rect 27649 9967 27683 10001
rect 27717 9967 27751 10001
rect 27785 9967 27819 10001
rect 26249 9962 27853 9967
rect 26249 9928 26277 9962
rect 26311 9928 26348 9962
rect 26382 9928 26419 9962
rect 26453 9928 26490 9962
rect 26524 9928 26561 9962
rect 26595 9928 26632 9962
rect 26666 9928 26703 9962
rect 26737 9928 26774 9962
rect 26808 9928 26845 9962
rect 26879 9928 26916 9962
rect 26950 9928 26986 9962
rect 27020 9928 27056 9962
rect 27090 9928 27126 9962
rect 27160 9928 27196 9962
rect 27230 9928 27266 9962
rect 27300 9928 27336 9962
rect 27370 9928 27406 9962
rect 27440 9932 27853 9962
rect 27440 9928 27547 9932
rect 26249 9898 27547 9928
rect 27581 9898 27615 9932
rect 27649 9898 27683 9932
rect 27717 9898 27751 9932
rect 27785 9898 27819 9932
rect 26249 9894 27853 9898
rect 26249 9860 26277 9894
rect 26311 9860 26348 9894
rect 26382 9860 26419 9894
rect 26453 9860 26490 9894
rect 26524 9860 26561 9894
rect 26595 9860 26632 9894
rect 26666 9860 26703 9894
rect 26737 9860 26774 9894
rect 26808 9860 26845 9894
rect 26879 9860 26916 9894
rect 26950 9860 26986 9894
rect 27020 9860 27056 9894
rect 27090 9860 27126 9894
rect 27160 9860 27196 9894
rect 27230 9860 27266 9894
rect 27300 9860 27336 9894
rect 27370 9860 27406 9894
rect 27440 9863 27853 9894
rect 27440 9860 27547 9863
rect 27581 9829 27615 9863
rect 27649 9829 27683 9863
rect 27717 9829 27751 9863
rect 27785 9829 27819 9863
rect 27547 9794 27853 9829
rect 27581 9760 27615 9794
rect 27649 9760 27683 9794
rect 27717 9760 27751 9794
rect 27785 9760 27819 9794
rect 27547 9724 27853 9760
rect 27581 9690 27615 9724
rect 27649 9690 27683 9724
rect 27717 9690 27751 9724
rect 27785 9690 27819 9724
rect 27547 9654 27853 9690
rect 27581 9620 27615 9654
rect 27649 9620 27683 9654
rect 27717 9620 27751 9654
rect 27785 9620 27819 9654
rect 27547 9584 27853 9620
rect 27581 9550 27615 9584
rect 27649 9550 27683 9584
rect 27717 9550 27751 9584
rect 27785 9550 27819 9584
rect 6746 9527 10219 9531
rect 6746 9508 10305 9527
rect 6746 9474 6751 9508
rect 6785 9474 6827 9508
rect 6861 9474 6903 9508
rect 6937 9474 6979 9508
rect 7013 9474 7055 9508
rect 7089 9474 7131 9508
rect 7165 9474 7207 9508
rect 7241 9496 10305 9508
rect 7241 9474 7332 9496
rect 6746 9462 7332 9474
rect 7366 9462 7401 9496
rect 7435 9462 7470 9496
rect 7504 9462 7539 9496
rect 7573 9462 7608 9496
rect 7642 9462 7677 9496
rect 7711 9462 7746 9496
rect 7780 9462 7815 9496
rect 7849 9462 7884 9496
rect 7918 9462 7953 9496
rect 7987 9462 8022 9496
rect 8056 9462 8091 9496
rect 8125 9462 8160 9496
rect 8194 9462 8229 9496
rect 8263 9462 8297 9496
rect 8331 9462 8365 9496
rect 8399 9462 8433 9496
rect 8467 9462 8501 9496
rect 8535 9462 8569 9496
rect 8603 9462 8637 9496
rect 8671 9462 8705 9496
rect 8739 9462 8773 9496
rect 8807 9462 8841 9496
rect 8875 9462 8909 9496
rect 8943 9462 8977 9496
rect 9011 9462 9045 9496
rect 9079 9462 9113 9496
rect 9147 9462 9181 9496
rect 9215 9462 9249 9496
rect 9283 9462 9317 9496
rect 9351 9462 9385 9496
rect 9419 9462 9453 9496
rect 9487 9462 9521 9496
rect 9555 9462 9589 9496
rect 9623 9462 9657 9496
rect 9691 9462 9725 9496
rect 9759 9462 9793 9496
rect 9827 9462 9861 9496
rect 9895 9462 9929 9496
rect 9963 9462 10049 9496
rect 10083 9462 10117 9496
rect 10151 9462 10185 9496
rect 10219 9493 10305 9496
rect 10339 9493 10405 9527
rect 10439 9493 10505 9527
rect 10539 9493 10607 9527
rect 10219 9462 10607 9493
rect 6746 9455 10607 9462
rect 6746 9440 10573 9455
rect 6746 9406 6751 9440
rect 6785 9406 6827 9440
rect 6861 9406 6903 9440
rect 6937 9406 6979 9440
rect 7013 9406 7055 9440
rect 7089 9406 7131 9440
rect 7165 9406 7207 9440
rect 7241 9427 10573 9440
rect 7241 9406 10049 9427
rect 6746 9404 10049 9406
rect 6746 9372 7332 9404
rect 6746 9338 6751 9372
rect 6785 9338 6827 9372
rect 6861 9338 6903 9372
rect 6937 9338 6979 9372
rect 7013 9338 7055 9372
rect 7089 9338 7131 9372
rect 7165 9338 7207 9372
rect 7241 9370 7332 9372
rect 7366 9370 7401 9404
rect 7435 9370 7470 9404
rect 7504 9370 7539 9404
rect 7573 9370 7608 9404
rect 7642 9370 7677 9404
rect 7711 9370 7746 9404
rect 7780 9370 7815 9404
rect 7849 9370 7884 9404
rect 7918 9370 7953 9404
rect 7987 9370 8022 9404
rect 8056 9370 8091 9404
rect 8125 9370 8160 9404
rect 8194 9370 8229 9404
rect 8263 9370 8297 9404
rect 8331 9370 8365 9404
rect 8399 9370 8433 9404
rect 8467 9370 8501 9404
rect 8535 9370 8569 9404
rect 8603 9370 8637 9404
rect 8671 9370 8705 9404
rect 8739 9370 8773 9404
rect 8807 9370 8841 9404
rect 8875 9370 8909 9404
rect 8943 9370 8977 9404
rect 9011 9370 9045 9404
rect 9079 9370 9113 9404
rect 9147 9370 9181 9404
rect 9215 9370 9249 9404
rect 9283 9370 9317 9404
rect 9351 9370 9385 9404
rect 9419 9370 9453 9404
rect 9487 9370 9521 9404
rect 9555 9370 9589 9404
rect 9623 9370 9657 9404
rect 9691 9370 9725 9404
rect 9759 9370 9793 9404
rect 9827 9370 9861 9404
rect 9895 9370 9929 9404
rect 9963 9393 10049 9404
rect 10083 9393 10117 9427
rect 10151 9393 10185 9427
rect 10219 9421 10573 9427
rect 27547 9514 27853 9550
rect 27581 9480 27615 9514
rect 27649 9480 27683 9514
rect 27717 9480 27751 9514
rect 27785 9480 27819 9514
rect 27547 9444 27853 9480
rect 10219 9403 10607 9421
rect 10219 9393 10305 9403
rect 9963 9370 10305 9393
rect 7241 9369 10305 9370
rect 10339 9369 10377 9403
rect 10411 9369 10449 9403
rect 10483 9383 10607 9403
rect 10483 9369 10573 9383
rect 7241 9338 7246 9369
rect 6746 9304 7246 9338
rect 6746 9270 6751 9304
rect 6785 9270 6827 9304
rect 6861 9270 6903 9304
rect 6937 9270 6979 9304
rect 7013 9270 7055 9304
rect 7089 9270 7131 9304
rect 7165 9270 7207 9304
rect 7241 9270 7246 9304
rect 6746 9236 7246 9270
rect 6746 9202 6751 9236
rect 6785 9202 6827 9236
rect 6861 9202 6903 9236
rect 6937 9202 6979 9236
rect 7013 9202 7055 9236
rect 7089 9202 7131 9236
rect 7165 9202 7207 9236
rect 7241 9202 7246 9236
rect 6746 9168 7246 9202
rect 6746 9134 6751 9168
rect 6785 9134 6827 9168
rect 6861 9134 6903 9168
rect 6937 9134 6979 9168
rect 7013 9134 7055 9168
rect 7089 9134 7131 9168
rect 7165 9134 7207 9168
rect 7241 9134 7246 9168
rect 6746 9100 7246 9134
rect 6746 9066 6751 9100
rect 6785 9066 6827 9100
rect 6861 9066 6903 9100
rect 6937 9066 6979 9100
rect 7013 9066 7055 9100
rect 7089 9066 7131 9100
rect 7165 9066 7207 9100
rect 7241 9066 7246 9100
rect 6746 9032 7246 9066
rect 6746 8998 6751 9032
rect 6785 8998 6827 9032
rect 6861 8998 6903 9032
rect 6937 8998 6979 9032
rect 7013 8998 7055 9032
rect 7089 8998 7131 9032
rect 7165 8998 7207 9032
rect 7241 8998 7246 9032
rect 6746 8964 7246 8998
rect 6746 8930 6751 8964
rect 6785 8930 6827 8964
rect 6861 8930 6903 8964
rect 6937 8930 6979 8964
rect 7013 8930 7055 8964
rect 7089 8930 7131 8964
rect 7165 8930 7207 8964
rect 7241 8930 7246 8964
rect 6746 8896 7246 8930
rect 6746 8862 6751 8896
rect 6785 8862 6827 8896
rect 6861 8862 6903 8896
rect 6937 8862 6979 8896
rect 7013 8862 7055 8896
rect 7089 8862 7131 8896
rect 7165 8862 7207 8896
rect 7241 8862 7246 8896
rect 168 8856 1846 8861
rect 168 8822 192 8856
rect 226 8822 262 8856
rect 296 8822 332 8856
rect 366 8822 402 8856
rect 436 8822 472 8856
rect 506 8822 542 8856
rect 576 8822 612 8856
rect 646 8822 682 8856
rect 716 8822 752 8856
rect 786 8822 822 8856
rect 856 8822 891 8856
rect 925 8822 960 8856
rect 994 8822 1029 8856
rect 1063 8822 1098 8856
rect 1132 8822 1167 8856
rect 1201 8822 1236 8856
rect 1270 8822 1305 8856
rect 1339 8822 1374 8856
rect 1408 8822 1443 8856
rect 1477 8822 1512 8856
rect 1546 8822 1581 8856
rect 1615 8822 1650 8856
rect 1684 8822 1719 8856
rect 1753 8822 1788 8856
rect 1822 8822 1846 8856
rect 168 8782 1846 8822
rect 168 8748 192 8782
rect 226 8748 262 8782
rect 296 8748 332 8782
rect 366 8748 402 8782
rect 436 8748 472 8782
rect 506 8748 542 8782
rect 576 8748 612 8782
rect 646 8748 682 8782
rect 716 8748 752 8782
rect 786 8748 822 8782
rect 856 8748 891 8782
rect 925 8748 960 8782
rect 994 8748 1029 8782
rect 1063 8748 1098 8782
rect 1132 8748 1167 8782
rect 1201 8748 1236 8782
rect 1270 8748 1305 8782
rect 1339 8748 1374 8782
rect 1408 8748 1443 8782
rect 1477 8748 1512 8782
rect 1546 8748 1581 8782
rect 1615 8748 1650 8782
rect 1684 8748 1719 8782
rect 1753 8748 1788 8782
rect 1822 8748 1846 8782
rect 168 8708 1846 8748
rect 168 8674 192 8708
rect 226 8674 262 8708
rect 296 8674 332 8708
rect 366 8674 402 8708
rect 436 8674 472 8708
rect 506 8674 542 8708
rect 576 8674 612 8708
rect 646 8674 682 8708
rect 716 8674 752 8708
rect 786 8674 822 8708
rect 856 8674 891 8708
rect 925 8674 960 8708
rect 994 8674 1029 8708
rect 1063 8674 1098 8708
rect 1132 8674 1167 8708
rect 1201 8674 1236 8708
rect 1270 8674 1305 8708
rect 1339 8674 1374 8708
rect 1408 8674 1443 8708
rect 1477 8674 1512 8708
rect 1546 8674 1581 8708
rect 1615 8674 1650 8708
rect 1684 8674 1719 8708
rect 1753 8674 1788 8708
rect 1822 8674 1846 8708
rect 168 8634 1846 8674
rect 168 8600 192 8634
rect 226 8600 262 8634
rect 296 8600 332 8634
rect 366 8600 402 8634
rect 436 8600 472 8634
rect 506 8600 542 8634
rect 576 8600 612 8634
rect 646 8600 682 8634
rect 716 8600 752 8634
rect 786 8600 822 8634
rect 856 8600 891 8634
rect 925 8600 960 8634
rect 994 8600 1029 8634
rect 1063 8600 1098 8634
rect 1132 8600 1167 8634
rect 1201 8600 1236 8634
rect 1270 8600 1305 8634
rect 1339 8600 1374 8634
rect 1408 8600 1443 8634
rect 1477 8600 1512 8634
rect 1546 8600 1581 8634
rect 1615 8600 1650 8634
rect 1684 8600 1719 8634
rect 1753 8600 1788 8634
rect 1822 8600 1846 8634
rect 168 8560 1846 8600
rect 168 8526 192 8560
rect 226 8526 262 8560
rect 296 8526 332 8560
rect 366 8526 402 8560
rect 436 8526 472 8560
rect 506 8526 542 8560
rect 576 8526 612 8560
rect 646 8526 682 8560
rect 716 8526 752 8560
rect 786 8526 822 8560
rect 856 8526 891 8560
rect 925 8526 960 8560
rect 994 8526 1029 8560
rect 1063 8526 1098 8560
rect 1132 8526 1167 8560
rect 1201 8526 1236 8560
rect 1270 8526 1305 8560
rect 1339 8526 1374 8560
rect 1408 8526 1443 8560
rect 1477 8526 1512 8560
rect 1546 8526 1581 8560
rect 1615 8526 1650 8560
rect 1684 8526 1719 8560
rect 1753 8526 1788 8560
rect 1822 8526 1846 8560
rect 168 8486 1846 8526
rect 6746 8828 7246 8862
rect 6746 8794 6751 8828
rect 6785 8794 6827 8828
rect 6861 8794 6903 8828
rect 6937 8794 6979 8828
rect 7013 8794 7055 8828
rect 7089 8794 7131 8828
rect 7165 8794 7207 8828
rect 7241 8794 7246 8828
rect 6746 8760 7246 8794
rect 6746 8726 6751 8760
rect 6785 8726 6827 8760
rect 6861 8726 6903 8760
rect 6937 8726 6979 8760
rect 7013 8726 7055 8760
rect 7089 8726 7131 8760
rect 7165 8726 7207 8760
rect 7241 8726 7246 8760
rect 6746 8692 7246 8726
rect 6746 8658 6751 8692
rect 6785 8658 6827 8692
rect 6861 8658 6903 8692
rect 6937 8658 6979 8692
rect 7013 8658 7055 8692
rect 7089 8658 7131 8692
rect 7165 8658 7207 8692
rect 7241 8658 7246 8692
rect 6746 8624 7246 8658
rect 6746 8590 6751 8624
rect 6785 8590 6827 8624
rect 6861 8590 6903 8624
rect 6937 8590 6979 8624
rect 7013 8590 7055 8624
rect 7089 8590 7131 8624
rect 7165 8590 7207 8624
rect 7241 8590 7246 8624
rect 6746 8555 7246 8590
rect 6746 8521 6751 8555
rect 6785 8521 6827 8555
rect 6861 8521 6903 8555
rect 6937 8521 6979 8555
rect 7013 8521 7055 8555
rect 7089 8521 7131 8555
rect 7165 8521 7207 8555
rect 7241 8521 7246 8555
rect 6746 8497 7246 8521
rect 10449 9349 10573 9369
rect 10449 9335 10607 9349
rect 10483 9311 10607 9335
rect 10483 9301 10573 9311
rect 10449 9277 10573 9301
rect 10449 9267 10607 9277
rect 10483 9239 10607 9267
rect 10483 9233 10573 9239
rect 10449 9205 10573 9233
rect 10449 9199 10607 9205
rect 10483 9167 10607 9199
rect 10483 9165 10573 9167
rect 10449 9133 10573 9165
rect 10449 9131 10607 9133
rect 10483 9097 10607 9131
rect 10449 9095 10607 9097
rect 10449 9063 10573 9095
rect 10483 9061 10573 9063
rect 10483 9029 10607 9061
rect 10449 9023 10607 9029
rect 10449 8995 10573 9023
rect 10483 8989 10573 8995
rect 23855 9431 24068 9434
rect 23855 9397 23879 9431
rect 23913 9397 24010 9431
rect 24044 9397 24068 9431
rect 23855 9351 24068 9397
rect 23855 9317 23879 9351
rect 23913 9317 24010 9351
rect 24044 9317 24068 9351
rect 23855 9271 24068 9317
rect 23855 9237 23879 9271
rect 23913 9237 24010 9271
rect 24044 9237 24068 9271
rect 23855 9191 24068 9237
rect 23855 9157 23879 9191
rect 23913 9157 24010 9191
rect 24044 9157 24068 9191
rect 23855 9111 24068 9157
rect 23855 9077 23879 9111
rect 23913 9077 24010 9111
rect 24044 9077 24068 9111
rect 23855 9031 24068 9077
rect 23855 9006 23879 9031
rect 10483 8961 10607 8989
rect 23654 8972 23659 9006
rect 23693 8972 23728 9006
rect 23762 8972 23797 9006
rect 23831 8997 23879 9006
rect 23913 8997 24010 9031
rect 24044 8997 24068 9031
rect 23831 8972 24068 8997
rect 10449 8950 10607 8961
rect 10449 8927 10573 8950
rect 10483 8916 10573 8927
rect 21694 8942 22862 8948
rect 10483 8893 10607 8916
rect 10449 8877 10607 8893
rect 10449 8859 10573 8877
rect 10483 8843 10573 8859
rect 10483 8825 10607 8843
rect 10449 8804 10607 8825
rect 10449 8791 10573 8804
rect 10483 8770 10573 8791
rect 10483 8757 10607 8770
rect 10449 8731 10607 8757
rect 10449 8723 10573 8731
rect 10483 8697 10573 8723
rect 10483 8689 10607 8697
rect 10449 8658 10607 8689
rect 10449 8654 10573 8658
rect 10483 8624 10573 8654
rect 10483 8620 10607 8624
rect 10449 8585 10607 8620
rect 10483 8551 10573 8585
rect 20784 8939 22862 8942
rect 20784 8905 20808 8939
rect 20842 8905 20883 8939
rect 20917 8905 20958 8939
rect 20992 8905 21033 8939
rect 21067 8905 21108 8939
rect 21142 8905 21183 8939
rect 21217 8905 21258 8939
rect 21292 8905 21332 8939
rect 21366 8905 21406 8939
rect 21440 8905 21480 8939
rect 21514 8908 22862 8939
rect 23846 8942 24068 8972
rect 23846 8908 23870 8942
rect 23904 8908 23940 8942
rect 23974 8908 24010 8942
rect 24044 8908 24068 8942
rect 27581 9410 27615 9444
rect 27649 9410 27683 9444
rect 27717 9410 27751 9444
rect 27785 9410 27819 9444
rect 27547 9374 27853 9410
rect 27581 9340 27615 9374
rect 27649 9340 27683 9374
rect 27717 9340 27751 9374
rect 27785 9340 27819 9374
rect 27547 9304 27853 9340
rect 27581 9270 27615 9304
rect 27649 9270 27683 9304
rect 27717 9270 27751 9304
rect 27785 9270 27819 9304
rect 27547 9234 27853 9270
rect 27581 9200 27615 9234
rect 27649 9200 27683 9234
rect 27717 9200 27751 9234
rect 27785 9200 27819 9234
rect 27547 9164 27853 9200
rect 27581 9130 27615 9164
rect 27649 9130 27683 9164
rect 27717 9130 27751 9164
rect 27785 9130 27819 9164
rect 27547 9094 27853 9130
rect 27581 9060 27615 9094
rect 27649 9060 27683 9094
rect 27717 9060 27751 9094
rect 27785 9060 27819 9094
rect 27547 9024 27853 9060
rect 27581 8990 27615 9024
rect 27649 8990 27683 9024
rect 27717 8990 27751 9024
rect 27785 8990 27819 9024
rect 27547 8954 27853 8990
rect 27581 8920 27615 8954
rect 27649 8920 27683 8954
rect 27717 8920 27751 8954
rect 27785 8920 27819 8954
rect 21514 8905 21572 8908
rect 20784 8874 21572 8905
rect 21606 8874 21648 8908
rect 21682 8874 21724 8908
rect 21758 8874 21800 8908
rect 21834 8874 21876 8908
rect 21910 8874 21952 8908
rect 21986 8874 22027 8908
rect 22061 8874 22102 8908
rect 22136 8890 22862 8908
rect 22136 8874 22194 8890
rect 20784 8871 22194 8874
rect 20784 8837 20808 8871
rect 20842 8837 20883 8871
rect 20917 8837 20958 8871
rect 20992 8837 21033 8871
rect 21067 8837 21108 8871
rect 21142 8837 21183 8871
rect 21217 8837 21258 8871
rect 21292 8837 21332 8871
rect 21366 8837 21406 8871
rect 21440 8837 21480 8871
rect 21514 8856 22194 8871
rect 22228 8856 22269 8890
rect 22303 8856 22344 8890
rect 22378 8856 22419 8890
rect 22453 8856 22494 8890
rect 22528 8856 22569 8890
rect 22603 8856 22643 8890
rect 22677 8856 22717 8890
rect 22751 8856 22791 8890
rect 22825 8856 22865 8890
rect 22899 8856 22923 8890
rect 21514 8840 22923 8856
rect 21514 8837 21572 8840
rect 20784 8806 21572 8837
rect 21606 8806 21648 8840
rect 21682 8806 21724 8840
rect 21758 8806 21800 8840
rect 21834 8806 21876 8840
rect 21910 8806 21952 8840
rect 21986 8806 22027 8840
rect 22061 8806 22102 8840
rect 22136 8822 22923 8840
rect 22136 8806 22194 8822
rect 20784 8803 21538 8806
rect 20784 8769 20808 8803
rect 20842 8769 20883 8803
rect 20917 8769 20958 8803
rect 20992 8769 21033 8803
rect 21067 8769 21108 8803
rect 21142 8769 21183 8803
rect 21217 8769 21258 8803
rect 21292 8769 21332 8803
rect 21366 8769 21406 8803
rect 21440 8769 21480 8803
rect 21514 8769 21538 8803
rect 20784 8735 21538 8769
rect 20784 8701 20808 8735
rect 20842 8701 20883 8735
rect 20917 8701 20958 8735
rect 20992 8701 21033 8735
rect 21067 8701 21108 8735
rect 21142 8701 21183 8735
rect 21217 8701 21258 8735
rect 21292 8701 21332 8735
rect 21366 8701 21406 8735
rect 21440 8701 21480 8735
rect 21514 8701 21538 8735
rect 20784 8667 21538 8701
rect 20784 8633 20808 8667
rect 20842 8633 20883 8667
rect 20917 8633 20958 8667
rect 20992 8633 21033 8667
rect 21067 8633 21108 8667
rect 21142 8633 21183 8667
rect 21217 8633 21258 8667
rect 21292 8633 21332 8667
rect 21366 8633 21406 8667
rect 21440 8633 21480 8667
rect 21514 8633 21538 8667
rect 20784 8599 21538 8633
rect 20784 8565 20808 8599
rect 20842 8565 20883 8599
rect 20917 8565 20958 8599
rect 20992 8565 21033 8599
rect 21067 8565 21108 8599
rect 21142 8565 21183 8599
rect 21217 8565 21258 8599
rect 21292 8565 21332 8599
rect 21366 8565 21406 8599
rect 21440 8565 21480 8599
rect 21514 8565 21538 8599
rect 22170 8788 22194 8806
rect 22228 8788 22269 8822
rect 22303 8788 22344 8822
rect 22378 8788 22419 8822
rect 22453 8788 22494 8822
rect 22528 8788 22569 8822
rect 22603 8788 22643 8822
rect 22677 8788 22717 8822
rect 22751 8788 22791 8822
rect 22825 8788 22865 8822
rect 22899 8788 22923 8822
rect 22170 8754 22923 8788
rect 22170 8720 22194 8754
rect 22228 8720 22269 8754
rect 22303 8720 22344 8754
rect 22378 8720 22419 8754
rect 22453 8720 22494 8754
rect 22528 8720 22569 8754
rect 22603 8720 22643 8754
rect 22677 8720 22717 8754
rect 22751 8720 22791 8754
rect 22825 8720 22865 8754
rect 22899 8720 22923 8754
rect 22170 8686 22923 8720
rect 22170 8652 22194 8686
rect 22228 8652 22269 8686
rect 22303 8652 22344 8686
rect 22378 8652 22419 8686
rect 22453 8652 22494 8686
rect 22528 8652 22569 8686
rect 22603 8652 22643 8686
rect 22677 8652 22717 8686
rect 22751 8652 22791 8686
rect 22825 8652 22865 8686
rect 22899 8652 22923 8686
rect 22170 8618 22923 8652
rect 22170 8584 22194 8618
rect 22228 8584 22269 8618
rect 22303 8584 22344 8618
rect 22378 8584 22419 8618
rect 22453 8584 22494 8618
rect 22528 8584 22569 8618
rect 22603 8584 22643 8618
rect 22677 8584 22717 8618
rect 22751 8584 22791 8618
rect 22825 8584 22865 8618
rect 22899 8584 22923 8618
rect 27547 8884 27853 8920
rect 27581 8850 27615 8884
rect 27649 8850 27683 8884
rect 27717 8850 27751 8884
rect 27785 8850 27819 8884
rect 27547 8814 27853 8850
rect 27581 8780 27615 8814
rect 27649 8780 27683 8814
rect 27717 8780 27751 8814
rect 27785 8780 27819 8814
rect 27547 8744 27853 8780
rect 27581 8710 27615 8744
rect 27649 8710 27683 8744
rect 27717 8710 27751 8744
rect 27785 8710 27819 8744
rect 27547 8674 27853 8710
rect 27581 8640 27615 8674
rect 27649 8640 27683 8674
rect 27717 8640 27751 8674
rect 27785 8640 27819 8674
rect 27547 8604 27853 8640
rect 20784 8562 21538 8565
rect 27581 8570 27615 8604
rect 27649 8570 27683 8604
rect 27717 8570 27751 8604
rect 27785 8570 27819 8604
rect 10449 8517 10607 8551
rect 27547 8534 27853 8570
rect 168 8452 192 8486
rect 226 8452 262 8486
rect 296 8452 332 8486
rect 366 8452 402 8486
rect 436 8452 472 8486
rect 506 8452 542 8486
rect 576 8452 612 8486
rect 646 8452 682 8486
rect 716 8452 752 8486
rect 786 8452 822 8486
rect 856 8452 891 8486
rect 925 8452 960 8486
rect 994 8452 1029 8486
rect 1063 8452 1098 8486
rect 1132 8452 1167 8486
rect 1201 8452 1236 8486
rect 1270 8452 1305 8486
rect 1339 8452 1374 8486
rect 1408 8452 1443 8486
rect 1477 8452 1512 8486
rect 1546 8452 1581 8486
rect 1615 8452 1650 8486
rect 1684 8452 1719 8486
rect 1753 8452 1788 8486
rect 1822 8452 1846 8486
rect 168 8412 1846 8452
rect 168 8378 192 8412
rect 226 8378 262 8412
rect 296 8378 332 8412
rect 366 8378 402 8412
rect 436 8378 472 8412
rect 506 8378 542 8412
rect 576 8378 612 8412
rect 646 8378 682 8412
rect 716 8378 752 8412
rect 786 8378 822 8412
rect 856 8378 891 8412
rect 925 8378 960 8412
rect 994 8378 1029 8412
rect 1063 8378 1098 8412
rect 1132 8378 1167 8412
rect 1201 8378 1236 8412
rect 1270 8378 1305 8412
rect 1339 8378 1374 8412
rect 1408 8378 1443 8412
rect 1477 8378 1512 8412
rect 1546 8378 1581 8412
rect 1615 8378 1650 8412
rect 1684 8378 1719 8412
rect 1753 8378 1788 8412
rect 1822 8378 1846 8412
rect 168 8338 1846 8378
rect 168 8304 192 8338
rect 226 8304 262 8338
rect 296 8304 332 8338
rect 366 8304 402 8338
rect 436 8304 472 8338
rect 506 8304 542 8338
rect 576 8304 612 8338
rect 646 8304 682 8338
rect 716 8304 752 8338
rect 786 8304 822 8338
rect 856 8304 891 8338
rect 925 8304 960 8338
rect 994 8304 1029 8338
rect 1063 8304 1098 8338
rect 1132 8304 1167 8338
rect 1201 8304 1236 8338
rect 1270 8304 1305 8338
rect 1339 8304 1374 8338
rect 1408 8304 1443 8338
rect 1477 8304 1512 8338
rect 1546 8304 1581 8338
rect 1615 8304 1650 8338
rect 1684 8304 1719 8338
rect 1753 8304 1788 8338
rect 1822 8304 1846 8338
rect 168 8256 1846 8304
rect 168 8222 175 8256
rect 209 8222 245 8256
rect 279 8222 315 8256
rect 349 8222 385 8256
rect 419 8222 455 8256
rect 489 8222 525 8256
rect 559 8222 595 8256
rect 629 8222 665 8256
rect 699 8222 735 8256
rect 769 8222 805 8256
rect 839 8235 1846 8256
rect 7088 8463 7246 8497
rect 7122 8429 7212 8463
rect 7088 8394 7246 8429
rect 7122 8360 7212 8394
rect 27581 8500 27615 8534
rect 27649 8500 27683 8534
rect 27717 8500 27751 8534
rect 27785 8500 27819 8534
rect 27547 8464 27853 8500
rect 27581 8430 27615 8464
rect 27649 8430 27683 8464
rect 27717 8430 27751 8464
rect 27785 8430 27819 8464
rect 27547 8378 27853 8430
rect 7088 8325 7246 8360
rect 7122 8291 7212 8325
rect 7088 8256 7246 8291
rect 839 8222 846 8235
rect 168 8188 846 8222
rect 168 8154 175 8188
rect 209 8154 245 8188
rect 279 8154 315 8188
rect 349 8154 385 8188
rect 419 8154 455 8188
rect 489 8154 525 8188
rect 559 8154 595 8188
rect 629 8154 665 8188
rect 699 8154 735 8188
rect 769 8154 805 8188
rect 839 8154 846 8188
rect 168 8120 846 8154
rect 168 8086 175 8120
rect 209 8086 245 8120
rect 279 8086 315 8120
rect 349 8086 385 8120
rect 419 8086 455 8120
rect 489 8086 525 8120
rect 559 8086 595 8120
rect 629 8086 665 8120
rect 699 8086 735 8120
rect 769 8086 805 8120
rect 839 8086 846 8120
rect 168 8052 846 8086
rect 168 8018 175 8052
rect 209 8018 245 8052
rect 279 8018 315 8052
rect 349 8018 385 8052
rect 419 8018 455 8052
rect 489 8018 525 8052
rect 559 8018 595 8052
rect 629 8018 665 8052
rect 699 8018 735 8052
rect 769 8018 805 8052
rect 839 8018 846 8052
rect 168 7984 846 8018
rect 168 7950 175 7984
rect 209 7950 245 7984
rect 279 7950 315 7984
rect 349 7950 385 7984
rect 419 7950 455 7984
rect 489 7950 525 7984
rect 559 7950 595 7984
rect 629 7950 665 7984
rect 699 7950 735 7984
rect 769 7950 805 7984
rect 839 7950 846 7984
rect 168 7915 846 7950
rect 168 7881 175 7915
rect 209 7881 245 7915
rect 279 7881 315 7915
rect 349 7881 385 7915
rect 419 7881 455 7915
rect 489 7881 525 7915
rect 559 7881 595 7915
rect 629 7881 665 7915
rect 699 7881 735 7915
rect 769 7881 805 7915
rect 839 7881 846 7915
rect 168 7846 846 7881
rect 168 7812 175 7846
rect 209 7812 245 7846
rect 279 7812 315 7846
rect 349 7812 385 7846
rect 419 7812 455 7846
rect 489 7812 525 7846
rect 559 7812 595 7846
rect 629 7812 665 7846
rect 699 7812 735 7846
rect 769 7812 805 7846
rect 839 7812 846 7846
rect 168 7777 846 7812
rect 168 7743 175 7777
rect 209 7743 245 7777
rect 279 7743 315 7777
rect 349 7743 385 7777
rect 419 7743 455 7777
rect 489 7743 525 7777
rect 559 7743 595 7777
rect 629 7743 665 7777
rect 699 7743 735 7777
rect 769 7743 805 7777
rect 839 7743 846 7777
rect 168 7708 846 7743
rect 168 7674 175 7708
rect 209 7674 245 7708
rect 279 7674 315 7708
rect 349 7674 385 7708
rect 419 7674 455 7708
rect 489 7674 525 7708
rect 559 7674 595 7708
rect 629 7674 665 7708
rect 699 7674 735 7708
rect 769 7674 805 7708
rect 839 7674 846 7708
rect 168 7639 846 7674
rect 168 7605 175 7639
rect 209 7605 245 7639
rect 279 7605 315 7639
rect 349 7605 385 7639
rect 419 7605 455 7639
rect 489 7605 525 7639
rect 559 7605 595 7639
rect 629 7605 665 7639
rect 699 7605 735 7639
rect 769 7605 805 7639
rect 839 7605 846 7639
rect 168 7570 846 7605
rect 168 7536 175 7570
rect 209 7536 245 7570
rect 279 7536 315 7570
rect 349 7536 385 7570
rect 419 7536 455 7570
rect 489 7536 525 7570
rect 559 7536 595 7570
rect 629 7536 665 7570
rect 699 7536 735 7570
rect 769 7536 805 7570
rect 839 7536 846 7570
rect 168 7501 846 7536
rect 168 7467 175 7501
rect 209 7467 245 7501
rect 279 7467 315 7501
rect 349 7467 385 7501
rect 419 7467 455 7501
rect 489 7467 525 7501
rect 559 7467 595 7501
rect 629 7467 665 7501
rect 699 7467 735 7501
rect 769 7467 805 7501
rect 839 7467 846 7501
rect 168 7432 846 7467
rect 168 7398 175 7432
rect 209 7398 245 7432
rect 279 7398 315 7432
rect 349 7398 385 7432
rect 419 7398 455 7432
rect 489 7398 525 7432
rect 559 7398 595 7432
rect 629 7398 665 7432
rect 699 7398 735 7432
rect 769 7398 805 7432
rect 839 7398 846 7432
rect 168 7363 846 7398
rect 168 7329 175 7363
rect 209 7329 245 7363
rect 279 7329 315 7363
rect 349 7329 385 7363
rect 419 7329 455 7363
rect 489 7329 525 7363
rect 559 7329 595 7363
rect 629 7329 665 7363
rect 699 7329 735 7363
rect 769 7329 805 7363
rect 839 7329 846 7363
rect 168 7294 846 7329
rect 168 7260 175 7294
rect 209 7260 245 7294
rect 279 7260 315 7294
rect 349 7260 385 7294
rect 419 7260 455 7294
rect 489 7260 525 7294
rect 559 7260 595 7294
rect 629 7260 665 7294
rect 699 7260 735 7294
rect 769 7260 805 7294
rect 839 7260 846 7294
rect 7122 8222 7212 8256
rect 7088 8187 7246 8222
rect 7122 8153 7212 8187
rect 7088 8118 7246 8153
rect 7122 8084 7212 8118
rect 7088 8048 7246 8084
rect 7122 8014 7212 8048
rect 7088 7978 7246 8014
rect 7122 7944 7212 7978
rect 7088 7908 7246 7944
rect 7122 7874 7212 7908
rect 7088 7838 7246 7874
rect 7122 7804 7212 7838
rect 7088 7768 7246 7804
rect 7122 7734 7212 7768
rect 7088 7698 7246 7734
rect 7122 7664 7212 7698
rect 7088 7628 7246 7664
rect 27270 8354 27853 8378
rect 27304 8320 27338 8354
rect 27372 8320 27406 8354
rect 27440 8320 27474 8354
rect 27508 8320 27542 8354
rect 27576 8320 27610 8354
rect 27644 8320 27678 8354
rect 27712 8320 27746 8354
rect 27780 8320 27814 8354
rect 27848 8320 27853 8354
rect 27270 8283 27853 8320
rect 27304 8249 27338 8283
rect 27372 8249 27406 8283
rect 27440 8249 27474 8283
rect 27508 8249 27542 8283
rect 27576 8249 27610 8283
rect 27644 8249 27678 8283
rect 27712 8249 27746 8283
rect 27780 8249 27814 8283
rect 27848 8249 27853 8283
rect 27270 8212 27853 8249
rect 27304 8178 27338 8212
rect 27372 8178 27406 8212
rect 27440 8178 27474 8212
rect 27508 8178 27542 8212
rect 27576 8178 27610 8212
rect 27644 8178 27678 8212
rect 27712 8178 27746 8212
rect 27780 8178 27814 8212
rect 27848 8178 27853 8212
rect 27270 8141 27853 8178
rect 27304 8107 27338 8141
rect 27372 8107 27406 8141
rect 27440 8107 27474 8141
rect 27508 8107 27542 8141
rect 27576 8107 27610 8141
rect 27644 8107 27678 8141
rect 27712 8107 27746 8141
rect 27780 8107 27814 8141
rect 27848 8107 27853 8141
rect 27270 8070 27853 8107
rect 27304 8036 27338 8070
rect 27372 8036 27406 8070
rect 27440 8036 27474 8070
rect 27508 8036 27542 8070
rect 27576 8036 27610 8070
rect 27644 8036 27678 8070
rect 27712 8036 27746 8070
rect 27780 8036 27814 8070
rect 27848 8036 27853 8070
rect 27270 7999 27853 8036
rect 27304 7965 27338 7999
rect 27372 7965 27406 7999
rect 27440 7965 27474 7999
rect 27508 7965 27542 7999
rect 27576 7965 27610 7999
rect 27644 7965 27678 7999
rect 27712 7965 27746 7999
rect 27780 7965 27814 7999
rect 27848 7965 27853 7999
rect 27270 7928 27853 7965
rect 27304 7894 27338 7928
rect 27372 7894 27406 7928
rect 27440 7894 27474 7928
rect 27508 7894 27542 7928
rect 27576 7894 27610 7928
rect 27644 7894 27678 7928
rect 27712 7894 27746 7928
rect 27780 7894 27814 7928
rect 27848 7894 27853 7928
rect 27270 7857 27853 7894
rect 27304 7823 27338 7857
rect 27372 7823 27406 7857
rect 27440 7823 27474 7857
rect 27508 7823 27542 7857
rect 27576 7823 27610 7857
rect 27644 7823 27678 7857
rect 27712 7823 27746 7857
rect 27780 7823 27814 7857
rect 27848 7823 27853 7857
rect 27270 7786 27853 7823
rect 27304 7752 27338 7786
rect 27372 7752 27406 7786
rect 27440 7752 27474 7786
rect 27508 7752 27542 7786
rect 27576 7752 27610 7786
rect 27644 7752 27678 7786
rect 27712 7752 27746 7786
rect 27780 7752 27814 7786
rect 27848 7752 27853 7786
rect 27270 7714 27853 7752
rect 27304 7680 27338 7714
rect 27372 7680 27406 7714
rect 27440 7680 27474 7714
rect 27508 7680 27542 7714
rect 27576 7680 27610 7714
rect 27644 7680 27678 7714
rect 27712 7680 27746 7714
rect 27780 7680 27814 7714
rect 27848 7680 27853 7714
rect 27270 7656 27853 7680
rect 7122 7594 7212 7628
rect 7088 7558 7246 7594
rect 7122 7524 7212 7558
rect 7088 7488 7246 7524
rect 7122 7454 7212 7488
rect 7088 7418 7246 7454
rect 7122 7384 7212 7418
rect 7088 7348 7246 7384
rect 7122 7314 7212 7348
rect 7088 7280 7246 7314
rect 168 7225 846 7260
rect 168 7191 175 7225
rect 209 7191 245 7225
rect 279 7191 315 7225
rect 349 7191 385 7225
rect 419 7191 455 7225
rect 489 7191 525 7225
rect 559 7191 595 7225
rect 629 7191 665 7225
rect 699 7191 735 7225
rect 769 7191 805 7225
rect 839 7191 846 7225
rect 168 7156 846 7191
rect 168 7122 175 7156
rect 209 7122 245 7156
rect 279 7122 315 7156
rect 349 7122 385 7156
rect 419 7122 455 7156
rect 489 7122 525 7156
rect 559 7122 595 7156
rect 629 7122 665 7156
rect 699 7122 735 7156
rect 769 7122 805 7156
rect 839 7122 846 7156
rect 168 7087 846 7122
rect 168 7053 175 7087
rect 209 7053 245 7087
rect 279 7053 315 7087
rect 349 7053 385 7087
rect 419 7053 455 7087
rect 489 7053 525 7087
rect 559 7053 595 7087
rect 629 7053 665 7087
rect 699 7053 735 7087
rect 769 7053 805 7087
rect 839 7053 846 7087
rect 168 7018 846 7053
rect 168 6984 175 7018
rect 209 6984 245 7018
rect 279 6984 315 7018
rect 349 6984 385 7018
rect 419 6984 455 7018
rect 489 6984 525 7018
rect 559 6984 595 7018
rect 629 6984 665 7018
rect 699 6984 735 7018
rect 769 6984 805 7018
rect 839 6984 846 7018
rect 168 6949 846 6984
rect 168 6915 175 6949
rect 209 6915 245 6949
rect 279 6915 315 6949
rect 349 6915 385 6949
rect 419 6915 455 6949
rect 489 6915 525 6949
rect 559 6915 595 6949
rect 629 6915 665 6949
rect 699 6915 735 6949
rect 769 6915 805 6949
rect 839 6915 846 6949
rect 14257 7013 15093 7037
rect 14257 6979 14262 7013
rect 14296 6979 14334 7013
rect 14368 6979 14406 7013
rect 14440 6979 14478 7013
rect 14512 6979 14550 7013
rect 14584 6979 14622 7013
rect 14656 6979 14694 7013
rect 14728 6979 14766 7013
rect 14800 6979 14838 7013
rect 14872 6979 14910 7013
rect 14944 6979 14982 7013
rect 15016 6979 15054 7013
rect 15088 6979 15093 7013
rect 14257 6940 15093 6979
rect 14257 6930 14262 6940
rect 168 6880 846 6915
rect 168 6846 175 6880
rect 209 6846 245 6880
rect 279 6846 315 6880
rect 349 6846 385 6880
rect 419 6846 455 6880
rect 489 6846 525 6880
rect 559 6846 595 6880
rect 629 6846 665 6880
rect 699 6846 735 6880
rect 769 6846 805 6880
rect 839 6846 846 6880
rect 168 6811 846 6846
rect 168 6777 175 6811
rect 209 6777 245 6811
rect 279 6777 315 6811
rect 349 6777 385 6811
rect 419 6777 455 6811
rect 489 6777 525 6811
rect 559 6777 595 6811
rect 629 6777 665 6811
rect 699 6777 735 6811
rect 769 6777 805 6811
rect 839 6777 846 6811
rect 168 6742 846 6777
rect 168 6708 175 6742
rect 209 6708 245 6742
rect 279 6708 315 6742
rect 349 6708 385 6742
rect 419 6708 455 6742
rect 489 6708 525 6742
rect 559 6708 595 6742
rect 629 6708 665 6742
rect 699 6708 735 6742
rect 769 6708 805 6742
rect 839 6708 846 6742
rect 168 6673 846 6708
rect 168 6639 175 6673
rect 209 6639 245 6673
rect 279 6639 315 6673
rect 349 6639 385 6673
rect 419 6639 455 6673
rect 489 6639 525 6673
rect 559 6639 595 6673
rect 629 6639 665 6673
rect 699 6639 735 6673
rect 769 6639 805 6673
rect 839 6639 846 6673
rect 168 6604 846 6639
rect 168 6570 175 6604
rect 209 6570 245 6604
rect 279 6570 315 6604
rect 349 6570 385 6604
rect 419 6570 455 6604
rect 489 6570 525 6604
rect 559 6570 595 6604
rect 629 6570 665 6604
rect 699 6570 735 6604
rect 769 6570 805 6604
rect 839 6570 846 6604
rect 168 6535 846 6570
rect 168 6501 175 6535
rect 209 6501 245 6535
rect 279 6501 315 6535
rect 349 6501 385 6535
rect 419 6501 455 6535
rect 489 6501 525 6535
rect 559 6501 595 6535
rect 629 6501 665 6535
rect 699 6501 735 6535
rect 769 6501 805 6535
rect 839 6501 846 6535
rect 168 6466 846 6501
rect 168 6432 175 6466
rect 209 6432 245 6466
rect 279 6432 315 6466
rect 349 6432 385 6466
rect 419 6432 455 6466
rect 489 6432 525 6466
rect 559 6432 595 6466
rect 629 6432 665 6466
rect 699 6432 735 6466
rect 769 6432 805 6466
rect 839 6432 846 6466
rect 168 6397 846 6432
rect 168 6363 175 6397
rect 209 6363 245 6397
rect 279 6363 315 6397
rect 349 6363 385 6397
rect 419 6363 455 6397
rect 489 6363 525 6397
rect 559 6363 595 6397
rect 629 6363 665 6397
rect 699 6363 735 6397
rect 769 6363 805 6397
rect 839 6363 846 6397
rect 168 6328 846 6363
rect 168 6294 175 6328
rect 209 6294 245 6328
rect 279 6294 315 6328
rect 349 6294 385 6328
rect 419 6294 455 6328
rect 489 6294 525 6328
rect 559 6294 595 6328
rect 629 6294 665 6328
rect 699 6294 735 6328
rect 769 6294 805 6328
rect 839 6294 846 6328
rect 168 6259 846 6294
rect 13030 6923 14262 6930
rect 13030 6889 13054 6923
rect 13088 6889 13123 6923
rect 13157 6889 13192 6923
rect 13226 6889 13261 6923
rect 13295 6889 13330 6923
rect 13364 6889 13399 6923
rect 13433 6889 13467 6923
rect 13501 6889 13535 6923
rect 13569 6889 13603 6923
rect 13637 6889 13671 6923
rect 13705 6889 13739 6923
rect 13773 6889 13807 6923
rect 13841 6889 13875 6923
rect 13909 6889 13943 6923
rect 13977 6889 14011 6923
rect 14045 6889 14079 6923
rect 14113 6889 14147 6923
rect 14181 6906 14262 6923
rect 14296 6906 14334 6940
rect 14368 6906 14406 6940
rect 14440 6906 14478 6940
rect 14512 6906 14550 6940
rect 14584 6906 14622 6940
rect 14656 6906 14694 6940
rect 14728 6906 14766 6940
rect 14800 6906 14838 6940
rect 14872 6906 14910 6940
rect 14944 6906 14982 6940
rect 15016 6906 15054 6940
rect 15088 6906 15093 6940
rect 14181 6889 15093 6906
rect 13030 6866 15093 6889
rect 13030 6849 14262 6866
rect 13030 6815 13054 6849
rect 13088 6815 13123 6849
rect 13157 6815 13192 6849
rect 13226 6815 13261 6849
rect 13295 6815 13330 6849
rect 13364 6815 13399 6849
rect 13433 6815 13467 6849
rect 13501 6815 13535 6849
rect 13569 6815 13603 6849
rect 13637 6815 13671 6849
rect 13705 6815 13739 6849
rect 13773 6815 13807 6849
rect 13841 6815 13875 6849
rect 13909 6815 13943 6849
rect 13977 6815 14011 6849
rect 14045 6815 14079 6849
rect 14113 6815 14147 6849
rect 14181 6832 14262 6849
rect 14296 6832 14334 6866
rect 14368 6832 14406 6866
rect 14440 6832 14478 6866
rect 14512 6832 14550 6866
rect 14584 6832 14622 6866
rect 14656 6832 14694 6866
rect 14728 6832 14766 6866
rect 14800 6832 14838 6866
rect 14872 6832 14910 6866
rect 14944 6832 14982 6866
rect 15016 6832 15054 6866
rect 15088 6832 15093 6866
rect 14181 6815 15093 6832
rect 13030 6792 15093 6815
rect 13030 6775 14262 6792
rect 13030 6741 13054 6775
rect 13088 6741 13123 6775
rect 13157 6741 13192 6775
rect 13226 6741 13261 6775
rect 13295 6741 13330 6775
rect 13364 6741 13399 6775
rect 13433 6741 13467 6775
rect 13501 6741 13535 6775
rect 13569 6741 13603 6775
rect 13637 6741 13671 6775
rect 13705 6741 13739 6775
rect 13773 6741 13807 6775
rect 13841 6741 13875 6775
rect 13909 6741 13943 6775
rect 13977 6741 14011 6775
rect 14045 6741 14079 6775
rect 14113 6741 14147 6775
rect 14181 6758 14262 6775
rect 14296 6758 14334 6792
rect 14368 6758 14406 6792
rect 14440 6758 14478 6792
rect 14512 6758 14550 6792
rect 14584 6758 14622 6792
rect 14656 6758 14694 6792
rect 14728 6758 14766 6792
rect 14800 6758 14838 6792
rect 14872 6758 14910 6792
rect 14944 6758 14982 6792
rect 15016 6758 15054 6792
rect 15088 6758 15093 6792
rect 14181 6741 15093 6758
rect 13030 6718 15093 6741
rect 13030 6701 14262 6718
rect 13030 6667 13054 6701
rect 13088 6667 13123 6701
rect 13157 6667 13192 6701
rect 13226 6667 13261 6701
rect 13295 6667 13330 6701
rect 13364 6667 13399 6701
rect 13433 6667 13467 6701
rect 13501 6667 13535 6701
rect 13569 6667 13603 6701
rect 13637 6667 13671 6701
rect 13705 6667 13739 6701
rect 13773 6667 13807 6701
rect 13841 6667 13875 6701
rect 13909 6667 13943 6701
rect 13977 6667 14011 6701
rect 14045 6667 14079 6701
rect 14113 6667 14147 6701
rect 14181 6684 14262 6701
rect 14296 6684 14334 6718
rect 14368 6684 14406 6718
rect 14440 6684 14478 6718
rect 14512 6684 14550 6718
rect 14584 6684 14622 6718
rect 14656 6684 14694 6718
rect 14728 6684 14766 6718
rect 14800 6684 14838 6718
rect 14872 6684 14910 6718
rect 14944 6684 14982 6718
rect 15016 6684 15054 6718
rect 15088 6684 15093 6718
rect 14181 6667 15093 6684
rect 13030 6644 15093 6667
rect 13030 6627 14262 6644
rect 13030 6593 13054 6627
rect 13088 6593 13123 6627
rect 13157 6593 13192 6627
rect 13226 6593 13261 6627
rect 13295 6593 13330 6627
rect 13364 6593 13399 6627
rect 13433 6593 13467 6627
rect 13501 6593 13535 6627
rect 13569 6593 13603 6627
rect 13637 6593 13671 6627
rect 13705 6593 13739 6627
rect 13773 6593 13807 6627
rect 13841 6593 13875 6627
rect 13909 6593 13943 6627
rect 13977 6593 14011 6627
rect 14045 6593 14079 6627
rect 14113 6593 14147 6627
rect 14181 6610 14262 6627
rect 14296 6610 14334 6644
rect 14368 6610 14406 6644
rect 14440 6610 14478 6644
rect 14512 6610 14550 6644
rect 14584 6610 14622 6644
rect 14656 6610 14694 6644
rect 14728 6610 14766 6644
rect 14800 6610 14838 6644
rect 14872 6610 14910 6644
rect 14944 6610 14982 6644
rect 15016 6610 15054 6644
rect 15088 6610 15093 6644
rect 14181 6593 15093 6610
rect 13030 6570 15093 6593
rect 13030 6553 14262 6570
rect 13030 6519 13054 6553
rect 13088 6519 13123 6553
rect 13157 6519 13192 6553
rect 13226 6519 13261 6553
rect 13295 6519 13330 6553
rect 13364 6519 13399 6553
rect 13433 6519 13467 6553
rect 13501 6519 13535 6553
rect 13569 6519 13603 6553
rect 13637 6519 13671 6553
rect 13705 6519 13739 6553
rect 13773 6519 13807 6553
rect 13841 6519 13875 6553
rect 13909 6519 13943 6553
rect 13977 6519 14011 6553
rect 14045 6519 14079 6553
rect 14113 6519 14147 6553
rect 14181 6536 14262 6553
rect 14296 6536 14334 6570
rect 14368 6536 14406 6570
rect 14440 6536 14478 6570
rect 14512 6536 14550 6570
rect 14584 6536 14622 6570
rect 14656 6536 14694 6570
rect 14728 6536 14766 6570
rect 14800 6536 14838 6570
rect 14872 6536 14910 6570
rect 14944 6536 14982 6570
rect 15016 6536 15054 6570
rect 15088 6536 15093 6570
rect 14181 6519 15093 6536
rect 13030 6496 15093 6519
rect 13030 6479 14262 6496
rect 13030 6445 13054 6479
rect 13088 6445 13123 6479
rect 13157 6445 13192 6479
rect 13226 6445 13261 6479
rect 13295 6445 13330 6479
rect 13364 6445 13399 6479
rect 13433 6445 13467 6479
rect 13501 6445 13535 6479
rect 13569 6445 13603 6479
rect 13637 6445 13671 6479
rect 13705 6445 13739 6479
rect 13773 6445 13807 6479
rect 13841 6445 13875 6479
rect 13909 6445 13943 6479
rect 13977 6445 14011 6479
rect 14045 6445 14079 6479
rect 14113 6445 14147 6479
rect 14181 6462 14262 6479
rect 14296 6462 14334 6496
rect 14368 6462 14406 6496
rect 14440 6462 14478 6496
rect 14512 6462 14550 6496
rect 14584 6462 14622 6496
rect 14656 6462 14694 6496
rect 14728 6462 14766 6496
rect 14800 6462 14838 6496
rect 14872 6462 14910 6496
rect 14944 6462 14982 6496
rect 15016 6462 15054 6496
rect 15088 6462 15093 6496
rect 14181 6445 15093 6462
rect 13030 6422 15093 6445
rect 13030 6405 14262 6422
rect 13030 6371 13054 6405
rect 13088 6371 13123 6405
rect 13157 6371 13192 6405
rect 13226 6371 13261 6405
rect 13295 6371 13330 6405
rect 13364 6371 13399 6405
rect 13433 6371 13467 6405
rect 13501 6371 13535 6405
rect 13569 6371 13603 6405
rect 13637 6371 13671 6405
rect 13705 6371 13739 6405
rect 13773 6371 13807 6405
rect 13841 6371 13875 6405
rect 13909 6371 13943 6405
rect 13977 6371 14011 6405
rect 14045 6371 14079 6405
rect 14113 6371 14147 6405
rect 14181 6388 14262 6405
rect 14296 6388 14334 6422
rect 14368 6388 14406 6422
rect 14440 6388 14478 6422
rect 14512 6388 14550 6422
rect 14584 6388 14622 6422
rect 14656 6388 14694 6422
rect 14728 6388 14766 6422
rect 14800 6388 14838 6422
rect 14872 6388 14910 6422
rect 14944 6388 14982 6422
rect 15016 6388 15054 6422
rect 15088 6388 15093 6422
rect 14181 6371 15093 6388
rect 13030 6348 15093 6371
rect 13030 6331 14262 6348
rect 13030 6297 13054 6331
rect 13088 6297 13123 6331
rect 13157 6297 13192 6331
rect 13226 6297 13261 6331
rect 13295 6297 13330 6331
rect 13364 6297 13399 6331
rect 13433 6297 13467 6331
rect 13501 6297 13535 6331
rect 13569 6297 13603 6331
rect 13637 6297 13671 6331
rect 13705 6297 13739 6331
rect 13773 6297 13807 6331
rect 13841 6297 13875 6331
rect 13909 6297 13943 6331
rect 13977 6297 14011 6331
rect 14045 6297 14079 6331
rect 14113 6297 14147 6331
rect 14181 6314 14262 6331
rect 14296 6314 14334 6348
rect 14368 6314 14406 6348
rect 14440 6314 14478 6348
rect 14512 6314 14550 6348
rect 14584 6314 14622 6348
rect 14656 6314 14694 6348
rect 14728 6314 14766 6348
rect 14800 6314 14838 6348
rect 14872 6314 14910 6348
rect 14944 6314 14982 6348
rect 15016 6314 15054 6348
rect 15088 6314 15093 6348
rect 14181 6297 15093 6314
rect 13030 6290 15093 6297
rect 168 6225 175 6259
rect 209 6225 245 6259
rect 279 6225 315 6259
rect 349 6225 385 6259
rect 419 6225 455 6259
rect 489 6225 525 6259
rect 559 6225 595 6259
rect 629 6225 665 6259
rect 699 6225 735 6259
rect 769 6225 805 6259
rect 839 6225 846 6259
rect 168 6201 846 6225
rect 168 6125 356 6201
rect 168 6091 169 6125
rect 203 6091 245 6125
rect 279 6091 321 6125
rect 355 6091 356 6125
rect 168 6056 356 6091
rect 168 6022 169 6056
rect 203 6022 245 6056
rect 279 6022 321 6056
rect 355 6022 356 6056
rect 168 5987 356 6022
rect 168 5953 169 5987
rect 203 5953 245 5987
rect 279 5953 321 5987
rect 355 5953 356 5987
rect 168 5918 356 5953
rect 168 5884 169 5918
rect 203 5884 245 5918
rect 279 5884 321 5918
rect 355 5884 356 5918
rect 168 5849 356 5884
rect 168 5815 169 5849
rect 203 5815 245 5849
rect 279 5815 321 5849
rect 355 5815 356 5849
rect 168 5780 356 5815
rect 168 5746 169 5780
rect 203 5746 245 5780
rect 279 5746 321 5780
rect 355 5746 356 5780
rect 168 5711 356 5746
rect 168 5677 169 5711
rect 203 5677 245 5711
rect 279 5677 321 5711
rect 355 5677 356 5711
rect 168 5642 356 5677
rect 168 5608 169 5642
rect 203 5608 245 5642
rect 279 5608 321 5642
rect 355 5608 356 5642
rect 168 5573 356 5608
rect 168 5539 169 5573
rect 203 5539 245 5573
rect 279 5539 321 5573
rect 355 5539 356 5573
rect 168 5504 356 5539
rect 168 5470 169 5504
rect 203 5470 245 5504
rect 279 5470 321 5504
rect 355 5470 356 5504
rect 168 5435 356 5470
rect 168 5401 169 5435
rect 203 5401 245 5435
rect 279 5401 321 5435
rect 355 5401 356 5435
rect 168 5366 356 5401
rect 168 5332 169 5366
rect 203 5332 245 5366
rect 279 5332 321 5366
rect 355 5332 356 5366
rect 168 5297 356 5332
rect 168 5263 169 5297
rect 203 5263 245 5297
rect 279 5263 321 5297
rect 355 5263 356 5297
rect 168 5228 356 5263
rect 168 5194 169 5228
rect 203 5194 245 5228
rect 279 5194 321 5228
rect 355 5194 356 5228
rect 168 5159 356 5194
rect 168 5125 169 5159
rect 203 5125 245 5159
rect 279 5125 321 5159
rect 355 5125 356 5159
rect 168 5090 356 5125
rect 168 5056 169 5090
rect 203 5056 245 5090
rect 279 5056 321 5090
rect 355 5056 356 5090
rect 168 5021 356 5056
rect 168 4987 169 5021
rect 203 4987 245 5021
rect 279 4987 321 5021
rect 355 4987 356 5021
rect 168 4952 356 4987
rect 168 4918 169 4952
rect 203 4918 245 4952
rect 279 4918 321 4952
rect 355 4918 408 4952
rect 168 4883 408 4918
rect 168 4849 169 4883
rect 203 4849 245 4883
rect 279 4849 321 4883
rect 355 4849 408 4883
rect 168 4814 408 4849
rect 168 4780 169 4814
rect 203 4780 245 4814
rect 279 4780 321 4814
rect 355 4780 408 4814
rect 168 4745 408 4780
rect 168 4711 169 4745
rect 203 4711 245 4745
rect 279 4711 321 4745
rect 355 4711 408 4745
rect 168 4676 408 4711
rect 168 4642 169 4676
rect 203 4642 245 4676
rect 279 4642 321 4676
rect 355 4642 408 4676
rect 168 4607 408 4642
rect 168 4573 169 4607
rect 203 4573 245 4607
rect 279 4573 321 4607
rect 355 4573 408 4607
rect 168 4538 408 4573
rect 168 4504 169 4538
rect 203 4504 245 4538
rect 279 4504 321 4538
rect 355 4504 408 4538
rect 168 4469 408 4504
rect 168 4435 169 4469
rect 203 4435 245 4469
rect 279 4435 321 4469
rect 355 4435 408 4469
rect 168 4400 408 4435
rect 168 4366 169 4400
rect 203 4366 245 4400
rect 279 4366 321 4400
rect 355 4366 408 4400
rect 168 4331 408 4366
rect 168 4297 169 4331
rect 203 4297 245 4331
rect 279 4297 321 4331
rect 355 4297 408 4331
rect 168 4262 408 4297
rect 168 4228 169 4262
rect 203 4228 245 4262
rect 279 4228 321 4262
rect 355 4228 408 4262
rect 168 4193 408 4228
rect 168 4159 169 4193
rect 203 4159 245 4193
rect 279 4159 321 4193
rect 355 4159 408 4193
rect 168 4156 408 4159
rect 168 4125 1048 4156
rect 168 4124 1074 4125
rect 168 4090 169 4124
rect 203 4090 245 4124
rect 279 4090 321 4124
rect 355 4107 1074 4124
rect 355 4090 2120 4107
rect 168 4081 2120 4090
rect 168 4055 442 4081
rect 168 4021 169 4055
rect 203 4021 245 4055
rect 279 4021 321 4055
rect 355 4047 442 4055
rect 476 4047 512 4081
rect 546 4047 582 4081
rect 616 4047 652 4081
rect 686 4047 722 4081
rect 756 4047 792 4081
rect 826 4047 862 4081
rect 896 4047 932 4081
rect 966 4047 1002 4081
rect 1036 4047 1072 4081
rect 1106 4047 1142 4081
rect 1176 4047 1212 4081
rect 1246 4047 1282 4081
rect 1316 4047 1352 4081
rect 1386 4047 1422 4081
rect 1456 4047 1492 4081
rect 1526 4047 1562 4081
rect 1596 4047 1632 4081
rect 1666 4047 1702 4081
rect 1736 4047 1772 4081
rect 1806 4047 1842 4081
rect 1876 4047 1912 4081
rect 1946 4047 1982 4081
rect 2016 4047 2052 4081
rect 2086 4047 2120 4081
rect 355 4021 2120 4047
rect 168 3986 2120 4021
rect 168 3952 169 3986
rect 203 3952 245 3986
rect 279 3952 321 3986
rect 355 3955 2120 3986
rect 355 3952 442 3955
rect 168 3921 442 3952
rect 476 3921 512 3955
rect 546 3921 582 3955
rect 616 3921 652 3955
rect 686 3921 722 3955
rect 756 3921 792 3955
rect 826 3921 862 3955
rect 896 3921 932 3955
rect 966 3921 1002 3955
rect 1036 3921 1072 3955
rect 1106 3921 1142 3955
rect 1176 3921 1212 3955
rect 1246 3921 1282 3955
rect 1316 3921 1352 3955
rect 1386 3921 1422 3955
rect 1456 3921 1492 3955
rect 1526 3921 1562 3955
rect 1596 3921 1632 3955
rect 1666 3921 1702 3955
rect 1736 3921 1772 3955
rect 1806 3921 1842 3955
rect 1876 3921 1912 3955
rect 1946 3921 1982 3955
rect 2016 3921 2052 3955
rect 2086 3921 2120 3955
rect 168 3917 668 3921
rect 168 3883 169 3917
rect 203 3883 245 3917
rect 279 3883 321 3917
rect 355 3883 668 3917
rect 168 3848 668 3883
rect 168 3814 169 3848
rect 203 3814 245 3848
rect 279 3814 321 3848
rect 355 3845 668 3848
rect 355 3814 410 3845
rect 168 3811 410 3814
rect 444 3811 484 3845
rect 518 3811 558 3845
rect 592 3811 632 3845
rect 666 3811 668 3845
rect 168 3779 668 3811
rect 168 3745 169 3779
rect 203 3745 245 3779
rect 279 3745 321 3779
rect 355 3774 668 3779
rect 355 3745 410 3774
rect 168 3740 410 3745
rect 444 3740 484 3774
rect 518 3740 558 3774
rect 592 3740 632 3774
rect 666 3740 668 3774
rect 168 3710 668 3740
rect 168 3676 169 3710
rect 203 3676 245 3710
rect 279 3676 321 3710
rect 355 3702 668 3710
rect 355 3676 410 3702
rect 168 3668 410 3676
rect 444 3668 484 3702
rect 518 3668 558 3702
rect 592 3668 632 3702
rect 666 3668 668 3702
rect 168 3641 668 3668
rect 168 3607 169 3641
rect 203 3607 245 3641
rect 279 3607 321 3641
rect 355 3630 668 3641
rect 355 3607 410 3630
rect 168 3596 410 3607
rect 444 3596 484 3630
rect 518 3596 558 3630
rect 592 3596 632 3630
rect 666 3596 668 3630
rect 168 3571 668 3596
rect 168 3537 169 3571
rect 203 3537 245 3571
rect 279 3537 321 3571
rect 355 3558 668 3571
rect 355 3537 410 3558
rect 168 3524 410 3537
rect 444 3524 484 3558
rect 518 3524 558 3558
rect 592 3524 632 3558
rect 666 3524 668 3558
rect 168 3501 668 3524
rect 168 3467 169 3501
rect 203 3467 245 3501
rect 279 3467 321 3501
rect 355 3486 668 3501
rect 355 3467 410 3486
rect 168 3452 410 3467
rect 444 3452 484 3486
rect 518 3452 558 3486
rect 592 3452 632 3486
rect 666 3452 668 3486
rect 168 3431 668 3452
rect 168 3397 169 3431
rect 203 3397 245 3431
rect 279 3397 321 3431
rect 355 3414 668 3431
rect 355 3397 410 3414
rect 168 3380 410 3397
rect 444 3380 484 3414
rect 518 3380 558 3414
rect 592 3380 632 3414
rect 666 3380 668 3414
rect 168 3361 668 3380
rect 168 3327 169 3361
rect 203 3327 245 3361
rect 279 3327 321 3361
rect 355 3342 668 3361
rect 355 3327 410 3342
rect 168 3308 410 3327
rect 444 3308 484 3342
rect 518 3308 558 3342
rect 592 3308 632 3342
rect 666 3308 668 3342
rect 168 3291 668 3308
rect 168 3257 169 3291
rect 203 3257 245 3291
rect 279 3257 321 3291
rect 355 3270 668 3291
rect 355 3257 410 3270
rect 168 3236 410 3257
rect 444 3236 484 3270
rect 518 3236 558 3270
rect 592 3236 632 3270
rect 666 3236 668 3270
rect 168 3221 668 3236
rect 168 3187 169 3221
rect 203 3187 245 3221
rect 279 3187 321 3221
rect 355 3198 668 3221
rect 355 3187 410 3198
rect 168 3164 410 3187
rect 444 3164 484 3198
rect 518 3164 558 3198
rect 592 3164 632 3198
rect 666 3164 668 3198
rect 168 3151 668 3164
rect 168 3117 169 3151
rect 203 3117 245 3151
rect 279 3117 321 3151
rect 355 3117 668 3151
rect 168 3089 668 3117
rect 1339 3841 2120 3921
rect 1339 3807 1373 3841
rect 1407 3807 1449 3841
rect 1483 3807 1525 3841
rect 1559 3807 1601 3841
rect 1635 3807 1677 3841
rect 1711 3807 1752 3841
rect 1786 3807 1827 3841
rect 1861 3807 1902 3841
rect 1936 3807 1977 3841
rect 2011 3807 2052 3841
rect 2086 3807 2120 3841
rect 1339 3761 2120 3807
rect 1339 3727 1373 3761
rect 1407 3727 1449 3761
rect 1483 3727 1525 3761
rect 1559 3727 1601 3761
rect 1635 3727 1677 3761
rect 1711 3727 1752 3761
rect 1786 3727 1827 3761
rect 1861 3727 1902 3761
rect 1936 3727 1977 3761
rect 2011 3727 2052 3761
rect 2086 3727 2120 3761
rect 1339 3681 2120 3727
rect 1339 3647 1373 3681
rect 1407 3647 1449 3681
rect 1483 3647 1525 3681
rect 1559 3647 1601 3681
rect 1635 3647 1677 3681
rect 1711 3647 1752 3681
rect 1786 3647 1827 3681
rect 1861 3647 1902 3681
rect 1936 3647 1977 3681
rect 2011 3647 2052 3681
rect 2086 3647 2120 3681
rect 1339 3601 2120 3647
rect 1339 3567 1373 3601
rect 1407 3567 1449 3601
rect 1483 3567 1525 3601
rect 1559 3567 1601 3601
rect 1635 3567 1677 3601
rect 1711 3567 1752 3601
rect 1786 3567 1827 3601
rect 1861 3567 1902 3601
rect 1936 3567 1977 3601
rect 2011 3567 2052 3601
rect 2086 3567 2120 3601
rect 1339 3521 2120 3567
rect 1339 3487 1373 3521
rect 1407 3487 1449 3521
rect 1483 3487 1525 3521
rect 1559 3487 1601 3521
rect 1635 3487 1677 3521
rect 1711 3487 1752 3521
rect 1786 3487 1827 3521
rect 1861 3487 1902 3521
rect 1936 3487 1977 3521
rect 2011 3487 2052 3521
rect 2086 3487 2120 3521
rect 1339 3441 2120 3487
rect 1339 3407 1373 3441
rect 1407 3407 1449 3441
rect 1483 3407 1525 3441
rect 1559 3407 1601 3441
rect 1635 3407 1677 3441
rect 1711 3407 1752 3441
rect 1786 3407 1827 3441
rect 1861 3407 1902 3441
rect 1936 3407 1977 3441
rect 2011 3407 2052 3441
rect 2086 3407 2120 3441
rect 1339 3371 2120 3407
rect 1339 3337 1389 3371
rect 1423 3337 1464 3371
rect 1498 3337 1539 3371
rect 1573 3337 1614 3371
rect 1648 3337 1689 3371
rect 1723 3337 1764 3371
rect 1798 3337 1839 3371
rect 1873 3337 1914 3371
rect 1948 3337 1988 3371
rect 2022 3337 2062 3371
rect 2096 3337 2120 3371
rect 1339 3303 2120 3337
rect 1339 3269 1389 3303
rect 1423 3269 1464 3303
rect 1498 3269 1539 3303
rect 1573 3269 1614 3303
rect 1648 3269 1689 3303
rect 1723 3269 1764 3303
rect 1798 3269 1839 3303
rect 1873 3269 1914 3303
rect 1948 3269 1988 3303
rect 2022 3269 2062 3303
rect 2096 3269 2120 3303
rect 1339 3233 2120 3269
rect 1339 3199 1363 3233
rect 1397 3199 1432 3233
rect 1466 3199 1501 3233
rect 1535 3199 1570 3233
rect 1604 3199 1639 3233
rect 1673 3199 1708 3233
rect 1742 3199 1777 3233
rect 1811 3199 1846 3233
rect 1880 3199 1915 3233
rect 1949 3199 1984 3233
rect 2018 3199 2053 3233
rect 2087 3199 2122 3233
rect 2156 3199 2191 3233
rect 2225 3199 2259 3233
rect 2293 3199 2327 3233
rect 2361 3199 2395 3233
rect 2429 3199 2463 3233
rect 2497 3199 2531 3233
rect 2565 3199 2599 3233
rect 2633 3199 2667 3233
rect 2701 3199 2735 3233
rect 2769 3199 2803 3233
rect 2837 3199 2871 3233
rect 2905 3199 2939 3233
rect 2973 3199 3007 3233
rect 3041 3199 3075 3233
rect 3109 3199 3133 3233
rect 1339 3159 3133 3199
rect 1339 3125 1363 3159
rect 1397 3125 1432 3159
rect 1466 3125 1501 3159
rect 1535 3125 1570 3159
rect 1604 3125 1639 3159
rect 1673 3125 1708 3159
rect 1742 3125 1777 3159
rect 1811 3125 1846 3159
rect 1880 3125 1915 3159
rect 1949 3125 1984 3159
rect 2018 3125 2053 3159
rect 2087 3125 2122 3159
rect 2156 3125 2191 3159
rect 2225 3125 2259 3159
rect 2293 3125 2327 3159
rect 2361 3125 2395 3159
rect 2429 3125 2463 3159
rect 2497 3125 2531 3159
rect 2565 3125 2599 3159
rect 2633 3125 2667 3159
rect 2701 3125 2735 3159
rect 2769 3125 2803 3159
rect 2837 3125 2871 3159
rect 2905 3125 2939 3159
rect 2973 3125 3007 3159
rect 3041 3125 3075 3159
rect 3109 3125 3133 3159
rect 1339 3089 3133 3125
rect 168 3087 3133 3089
rect 168 3081 410 3087
rect 168 3047 169 3081
rect 203 3047 245 3081
rect 279 3047 321 3081
rect 355 3053 410 3081
rect 444 3053 481 3087
rect 515 3053 552 3087
rect 586 3053 623 3087
rect 657 3053 694 3087
rect 728 3053 765 3087
rect 799 3053 835 3087
rect 869 3053 905 3087
rect 939 3053 975 3087
rect 1009 3053 1045 3087
rect 1079 3053 1115 3087
rect 1149 3053 1185 3087
rect 1219 3053 1255 3087
rect 1289 3085 3133 3087
rect 1289 3053 1363 3085
rect 355 3051 1363 3053
rect 1397 3051 1432 3085
rect 1466 3051 1501 3085
rect 1535 3051 1570 3085
rect 1604 3051 1639 3085
rect 1673 3051 1708 3085
rect 1742 3051 1777 3085
rect 1811 3051 1846 3085
rect 1880 3051 1915 3085
rect 1949 3051 1984 3085
rect 2018 3051 2053 3085
rect 2087 3051 2122 3085
rect 2156 3051 2191 3085
rect 2225 3051 2259 3085
rect 2293 3051 2327 3085
rect 2361 3051 2395 3085
rect 2429 3051 2463 3085
rect 2497 3051 2531 3085
rect 2565 3051 2599 3085
rect 2633 3051 2667 3085
rect 2701 3051 2735 3085
rect 2769 3051 2803 3085
rect 2837 3051 2871 3085
rect 2905 3051 2939 3085
rect 2973 3051 3007 3085
rect 3041 3051 3075 3085
rect 3109 3051 3133 3085
rect 355 3047 3133 3051
rect 168 3013 3133 3047
rect 168 3011 410 3013
rect 168 2977 169 3011
rect 203 2977 245 3011
rect 279 2977 321 3011
rect 355 2979 410 3011
rect 444 2979 481 3013
rect 515 2979 552 3013
rect 586 2979 623 3013
rect 657 2979 694 3013
rect 728 2979 765 3013
rect 799 2979 835 3013
rect 869 2979 905 3013
rect 939 2979 975 3013
rect 1009 2979 1045 3013
rect 1079 2979 1115 3013
rect 1149 2979 1185 3013
rect 1219 2979 1255 3013
rect 1289 3011 3133 3013
rect 1289 2979 1363 3011
rect 355 2977 1363 2979
rect 1397 2977 1432 3011
rect 1466 2977 1501 3011
rect 1535 2977 1570 3011
rect 1604 2977 1639 3011
rect 1673 2977 1708 3011
rect 1742 2977 1777 3011
rect 1811 2977 1846 3011
rect 1880 2977 1915 3011
rect 1949 2977 1984 3011
rect 2018 2977 2053 3011
rect 2087 2977 2122 3011
rect 2156 2977 2191 3011
rect 2225 2977 2259 3011
rect 2293 2977 2327 3011
rect 2361 2977 2395 3011
rect 2429 2977 2463 3011
rect 2497 2977 2531 3011
rect 2565 2977 2599 3011
rect 2633 2977 2667 3011
rect 2701 2977 2735 3011
rect 2769 2977 2803 3011
rect 2837 2977 2871 3011
rect 2905 2977 2939 3011
rect 2973 2977 3007 3011
rect 3041 2977 3075 3011
rect 3109 2977 3133 3011
rect 168 2941 3133 2977
rect 168 2907 169 2941
rect 203 2907 245 2941
rect 279 2907 321 2941
rect 355 2939 3133 2941
rect 355 2907 410 2939
rect 168 2905 410 2907
rect 444 2905 481 2939
rect 515 2905 552 2939
rect 586 2905 623 2939
rect 657 2905 694 2939
rect 728 2905 765 2939
rect 799 2905 835 2939
rect 869 2905 905 2939
rect 939 2905 975 2939
rect 1009 2905 1045 2939
rect 1079 2905 1115 2939
rect 1149 2905 1185 2939
rect 1219 2905 1255 2939
rect 1289 2937 3133 2939
rect 1289 2905 1363 2937
rect 168 2903 1363 2905
rect 1397 2903 1432 2937
rect 1466 2903 1501 2937
rect 1535 2903 1570 2937
rect 1604 2903 1639 2937
rect 1673 2903 1708 2937
rect 1742 2903 1777 2937
rect 1811 2903 1846 2937
rect 1880 2903 1915 2937
rect 1949 2903 1984 2937
rect 2018 2903 2053 2937
rect 2087 2903 2122 2937
rect 2156 2903 2191 2937
rect 2225 2903 2259 2937
rect 2293 2903 2327 2937
rect 2361 2903 2395 2937
rect 2429 2903 2463 2937
rect 2497 2903 2531 2937
rect 2565 2903 2599 2937
rect 2633 2903 2667 2937
rect 2701 2903 2735 2937
rect 2769 2903 2803 2937
rect 2837 2903 2871 2937
rect 2905 2903 2939 2937
rect 2973 2903 3007 2937
rect 3041 2903 3075 2937
rect 3109 2903 3133 2937
rect 168 2871 3133 2903
rect 168 2837 169 2871
rect 203 2837 245 2871
rect 279 2837 321 2871
rect 355 2865 3133 2871
rect 355 2837 410 2865
rect 168 2831 410 2837
rect 444 2831 481 2865
rect 515 2831 552 2865
rect 586 2831 623 2865
rect 657 2831 694 2865
rect 728 2831 765 2865
rect 799 2831 835 2865
rect 869 2831 905 2865
rect 939 2831 975 2865
rect 1009 2831 1045 2865
rect 1079 2831 1115 2865
rect 1149 2831 1185 2865
rect 1219 2831 1255 2865
rect 1289 2863 3133 2865
rect 1289 2831 1363 2863
rect 168 2829 1363 2831
rect 1397 2829 1432 2863
rect 1466 2829 1501 2863
rect 1535 2829 1570 2863
rect 1604 2829 1639 2863
rect 1673 2829 1708 2863
rect 1742 2829 1777 2863
rect 1811 2829 1846 2863
rect 1880 2829 1915 2863
rect 1949 2829 1984 2863
rect 2018 2829 2053 2863
rect 2087 2829 2122 2863
rect 2156 2829 2191 2863
rect 2225 2829 2259 2863
rect 2293 2829 2327 2863
rect 2361 2829 2395 2863
rect 2429 2829 2463 2863
rect 2497 2829 2531 2863
rect 2565 2829 2599 2863
rect 2633 2829 2667 2863
rect 2701 2829 2735 2863
rect 2769 2829 2803 2863
rect 2837 2829 2871 2863
rect 2905 2829 2939 2863
rect 2973 2829 3007 2863
rect 3041 2829 3075 2863
rect 3109 2829 3133 2863
rect 168 2801 3133 2829
rect 168 2767 169 2801
rect 203 2767 245 2801
rect 279 2767 321 2801
rect 355 2791 3133 2801
rect 355 2767 410 2791
rect 168 2757 410 2767
rect 444 2757 481 2791
rect 515 2757 552 2791
rect 586 2757 623 2791
rect 657 2757 694 2791
rect 728 2757 765 2791
rect 799 2757 835 2791
rect 869 2757 905 2791
rect 939 2757 975 2791
rect 1009 2757 1045 2791
rect 1079 2757 1115 2791
rect 1149 2757 1185 2791
rect 1219 2757 1255 2791
rect 1289 2789 3133 2791
rect 1289 2757 1363 2789
rect 168 2755 1363 2757
rect 1397 2755 1432 2789
rect 1466 2755 1501 2789
rect 1535 2755 1570 2789
rect 1604 2755 1639 2789
rect 1673 2755 1708 2789
rect 1742 2755 1777 2789
rect 1811 2755 1846 2789
rect 1880 2755 1915 2789
rect 1949 2755 1984 2789
rect 2018 2755 2053 2789
rect 2087 2755 2122 2789
rect 2156 2755 2191 2789
rect 2225 2755 2259 2789
rect 2293 2755 2327 2789
rect 2361 2755 2395 2789
rect 2429 2755 2463 2789
rect 2497 2755 2531 2789
rect 2565 2755 2599 2789
rect 2633 2755 2667 2789
rect 2701 2755 2735 2789
rect 2769 2755 2803 2789
rect 2837 2755 2871 2789
rect 2905 2755 2939 2789
rect 2973 2755 3007 2789
rect 3041 2755 3075 2789
rect 3109 2755 3133 2789
rect 168 2731 3133 2755
rect 168 2697 169 2731
rect 203 2697 245 2731
rect 279 2697 321 2731
rect 355 2717 3133 2731
rect 355 2697 410 2717
rect 168 2683 410 2697
rect 444 2683 481 2717
rect 515 2683 552 2717
rect 586 2683 623 2717
rect 657 2683 694 2717
rect 728 2683 765 2717
rect 799 2683 835 2717
rect 869 2683 905 2717
rect 939 2683 975 2717
rect 1009 2683 1045 2717
rect 1079 2683 1115 2717
rect 1149 2683 1185 2717
rect 1219 2683 1255 2717
rect 1289 2715 3133 2717
rect 1289 2683 1363 2715
rect 168 2681 1363 2683
rect 1397 2681 1432 2715
rect 1466 2681 1501 2715
rect 1535 2681 1570 2715
rect 1604 2681 1639 2715
rect 1673 2681 1708 2715
rect 1742 2681 1777 2715
rect 1811 2681 1846 2715
rect 1880 2681 1915 2715
rect 1949 2681 1984 2715
rect 2018 2681 2053 2715
rect 2087 2681 2122 2715
rect 2156 2681 2191 2715
rect 2225 2681 2259 2715
rect 2293 2681 2327 2715
rect 2361 2681 2395 2715
rect 2429 2681 2463 2715
rect 2497 2681 2531 2715
rect 2565 2681 2599 2715
rect 2633 2681 2667 2715
rect 2701 2681 2735 2715
rect 2769 2681 2803 2715
rect 2837 2681 2871 2715
rect 2905 2681 2939 2715
rect 2973 2681 3007 2715
rect 3041 2681 3075 2715
rect 3109 2681 3133 2715
rect 168 2661 3133 2681
rect 168 2627 169 2661
rect 203 2627 245 2661
rect 279 2627 321 2661
rect 355 2643 3133 2661
rect 355 2627 410 2643
rect 168 2609 410 2627
rect 444 2609 481 2643
rect 515 2609 552 2643
rect 586 2609 623 2643
rect 657 2609 694 2643
rect 728 2609 765 2643
rect 799 2609 835 2643
rect 869 2609 905 2643
rect 939 2609 975 2643
rect 1009 2609 1045 2643
rect 1079 2609 1115 2643
rect 1149 2609 1185 2643
rect 1219 2609 1255 2643
rect 1289 2641 3133 2643
rect 1289 2609 1363 2641
rect 168 2607 1363 2609
rect 1397 2607 1432 2641
rect 1466 2607 1501 2641
rect 1535 2607 1570 2641
rect 1604 2607 1639 2641
rect 1673 2607 1708 2641
rect 1742 2607 1777 2641
rect 1811 2607 1846 2641
rect 1880 2607 1915 2641
rect 1949 2607 1984 2641
rect 2018 2607 2053 2641
rect 2087 2607 2122 2641
rect 2156 2607 2191 2641
rect 2225 2607 2259 2641
rect 2293 2607 2327 2641
rect 2361 2607 2395 2641
rect 2429 2607 2463 2641
rect 2497 2607 2531 2641
rect 2565 2607 2599 2641
rect 2633 2607 2667 2641
rect 2701 2607 2735 2641
rect 2769 2607 2803 2641
rect 2837 2607 2871 2641
rect 2905 2607 2939 2641
rect 2973 2607 3007 2641
rect 3041 2607 3075 2641
rect 3109 2607 3133 2641
rect 168 2591 3133 2607
rect 168 2557 169 2591
rect 203 2557 245 2591
rect 279 2557 321 2591
rect 355 2569 3133 2591
rect 355 2557 410 2569
rect 168 2535 410 2557
rect 444 2535 481 2569
rect 515 2535 552 2569
rect 586 2535 623 2569
rect 657 2535 694 2569
rect 728 2535 765 2569
rect 799 2535 835 2569
rect 869 2535 905 2569
rect 939 2535 975 2569
rect 1009 2535 1045 2569
rect 1079 2535 1115 2569
rect 1149 2535 1185 2569
rect 1219 2535 1255 2569
rect 1289 2567 3133 2569
rect 1289 2535 1363 2567
rect 168 2533 1363 2535
rect 1397 2533 1432 2567
rect 1466 2533 1501 2567
rect 1535 2533 1570 2567
rect 1604 2533 1639 2567
rect 1673 2533 1708 2567
rect 1742 2533 1777 2567
rect 1811 2533 1846 2567
rect 1880 2533 1915 2567
rect 1949 2533 1984 2567
rect 2018 2533 2053 2567
rect 2087 2533 2122 2567
rect 2156 2533 2191 2567
rect 2225 2533 2259 2567
rect 2293 2533 2327 2567
rect 2361 2533 2395 2567
rect 2429 2533 2463 2567
rect 2497 2533 2531 2567
rect 2565 2533 2599 2567
rect 2633 2533 2667 2567
rect 2701 2533 2735 2567
rect 2769 2533 2803 2567
rect 2837 2533 2871 2567
rect 2905 2533 2939 2567
rect 2973 2533 3007 2567
rect 3041 2533 3075 2567
rect 3109 2533 3133 2567
rect 25812 2033 27880 2034
rect 25812 1999 25846 2033
rect 25880 1999 25917 2033
rect 25951 1999 25988 2033
rect 26022 1999 26059 2033
rect 26093 1999 26130 2033
rect 26164 1999 26201 2033
rect 26235 1999 26272 2033
rect 26306 1999 26342 2033
rect 26376 1999 26412 2033
rect 26446 1999 26482 2033
rect 26516 1999 26552 2033
rect 26586 1999 26622 2033
rect 26656 1999 26692 2033
rect 26726 1999 26762 2033
rect 26796 1999 26832 2033
rect 26866 1999 26902 2033
rect 26936 1999 26972 2033
rect 27006 1999 27042 2033
rect 27076 1999 27112 2033
rect 27146 1999 27182 2033
rect 27216 1999 27252 2033
rect 27286 1999 27322 2033
rect 27356 1999 27392 2033
rect 27426 1999 27462 2033
rect 27496 1999 27532 2033
rect 27566 1999 27602 2033
rect 27636 1999 27672 2033
rect 27706 1999 27742 2033
rect 27776 1999 27812 2033
rect 27846 1999 27880 2033
rect 25812 1947 27880 1999
rect 25812 1913 25846 1947
rect 25880 1913 25917 1947
rect 25951 1913 25988 1947
rect 26022 1913 26059 1947
rect 26093 1913 26130 1947
rect 26164 1913 26201 1947
rect 26235 1913 26272 1947
rect 26306 1913 26342 1947
rect 26376 1913 26412 1947
rect 26446 1913 26482 1947
rect 26516 1913 26552 1947
rect 26586 1913 26622 1947
rect 26656 1913 26692 1947
rect 26726 1913 26762 1947
rect 26796 1913 26832 1947
rect 26866 1913 26902 1947
rect 26936 1913 26972 1947
rect 27006 1913 27042 1947
rect 27076 1913 27112 1947
rect 27146 1913 27182 1947
rect 27216 1913 27252 1947
rect 27286 1913 27322 1947
rect 27356 1913 27392 1947
rect 27426 1913 27462 1947
rect 27496 1913 27532 1947
rect 27566 1913 27602 1947
rect 27636 1913 27672 1947
rect 27706 1913 27742 1947
rect 27776 1913 27812 1947
rect 27846 1913 27880 1947
rect 25812 1861 27880 1913
rect 25812 1827 25846 1861
rect 25880 1827 25917 1861
rect 25951 1827 25988 1861
rect 26022 1827 26059 1861
rect 26093 1827 26130 1861
rect 26164 1827 26201 1861
rect 26235 1827 26272 1861
rect 26306 1827 26342 1861
rect 26376 1827 26412 1861
rect 26446 1827 26482 1861
rect 26516 1827 26552 1861
rect 26586 1827 26622 1861
rect 26656 1827 26692 1861
rect 26726 1827 26762 1861
rect 26796 1827 26832 1861
rect 26866 1827 26902 1861
rect 26936 1827 26972 1861
rect 27006 1827 27042 1861
rect 27076 1827 27112 1861
rect 27146 1827 27182 1861
rect 27216 1827 27252 1861
rect 27286 1827 27322 1861
rect 27356 1827 27392 1861
rect 27426 1827 27462 1861
rect 27496 1827 27532 1861
rect 27566 1827 27602 1861
rect 27636 1827 27672 1861
rect 27706 1827 27742 1861
rect 27776 1827 27812 1861
rect 27846 1827 27880 1861
rect 25812 1775 27880 1827
rect 25812 1741 25846 1775
rect 25880 1741 25917 1775
rect 25951 1741 25988 1775
rect 26022 1741 26059 1775
rect 26093 1741 26130 1775
rect 26164 1741 26201 1775
rect 26235 1741 26272 1775
rect 26306 1741 26342 1775
rect 26376 1741 26412 1775
rect 26446 1741 26482 1775
rect 26516 1741 26552 1775
rect 26586 1741 26622 1775
rect 26656 1741 26692 1775
rect 26726 1741 26762 1775
rect 26796 1741 26832 1775
rect 26866 1741 26902 1775
rect 26936 1741 26972 1775
rect 27006 1741 27042 1775
rect 27076 1741 27112 1775
rect 27146 1741 27182 1775
rect 27216 1741 27252 1775
rect 27286 1741 27322 1775
rect 27356 1741 27392 1775
rect 27426 1741 27462 1775
rect 27496 1741 27532 1775
rect 27566 1741 27602 1775
rect 27636 1741 27672 1775
rect 27706 1741 27742 1775
rect 27776 1741 27812 1775
rect 27846 1741 27880 1775
rect 25812 1740 27880 1741
<< mvnsubdiff >>
rect 2335 20750 3196 20804
rect 2335 20716 2401 20750
rect 2435 20716 2474 20750
rect 2508 20716 2547 20750
rect 2581 20716 2620 20750
rect 2654 20716 2693 20750
rect 2727 20716 2766 20750
rect 2800 20716 2839 20750
rect 2873 20716 2912 20750
rect 2946 20716 2984 20750
rect 3018 20716 3056 20750
rect 3090 20716 3128 20750
rect 3162 20716 3196 20750
rect 2335 20672 3196 20716
rect 2335 20638 2401 20672
rect 2435 20638 2474 20672
rect 2508 20638 2547 20672
rect 2581 20638 2620 20672
rect 2654 20638 2693 20672
rect 2727 20638 2766 20672
rect 2800 20638 2839 20672
rect 2873 20638 2912 20672
rect 2946 20638 2984 20672
rect 3018 20638 3056 20672
rect 3090 20638 3128 20672
rect 3162 20638 3196 20672
rect 2335 20594 3196 20638
rect 2335 20560 2401 20594
rect 2435 20560 2474 20594
rect 2508 20560 2547 20594
rect 2581 20560 2620 20594
rect 2654 20560 2693 20594
rect 2727 20560 2766 20594
rect 2800 20560 2839 20594
rect 2873 20560 2912 20594
rect 2946 20560 2984 20594
rect 3018 20560 3056 20594
rect 3090 20560 3128 20594
rect 3162 20560 3196 20594
rect 2335 20516 3196 20560
rect 2335 20482 2401 20516
rect 2435 20482 2474 20516
rect 2508 20482 2547 20516
rect 2581 20482 2620 20516
rect 2654 20482 2693 20516
rect 2727 20482 2766 20516
rect 2800 20482 2839 20516
rect 2873 20482 2912 20516
rect 2946 20482 2984 20516
rect 3018 20482 3056 20516
rect 3090 20482 3128 20516
rect 3162 20482 3196 20516
rect 2335 20438 3196 20482
rect 2335 20404 2401 20438
rect 2435 20404 2474 20438
rect 2508 20404 2547 20438
rect 2581 20404 2620 20438
rect 2654 20404 2693 20438
rect 2727 20404 2766 20438
rect 2800 20404 2839 20438
rect 2873 20404 2912 20438
rect 2946 20404 2984 20438
rect 3018 20404 3056 20438
rect 3090 20404 3128 20438
rect 3162 20404 3196 20438
rect 26366 20718 26952 20804
rect 26366 20684 26371 20718
rect 26405 20684 26441 20718
rect 26475 20684 26511 20718
rect 26545 20684 26581 20718
rect 26615 20684 26651 20718
rect 26685 20684 26721 20718
rect 26755 20684 26791 20718
rect 26825 20684 26861 20718
rect 26895 20684 26952 20718
rect 26366 20647 26952 20684
rect 26366 20613 26371 20647
rect 26405 20613 26441 20647
rect 26475 20613 26511 20647
rect 26545 20613 26581 20647
rect 26615 20613 26651 20647
rect 26685 20613 26721 20647
rect 26755 20613 26791 20647
rect 26825 20613 26861 20647
rect 26895 20613 26952 20647
rect 26366 20576 26952 20613
rect 26366 20542 26371 20576
rect 26405 20542 26441 20576
rect 26475 20542 26511 20576
rect 26545 20542 26581 20576
rect 26615 20542 26651 20576
rect 26685 20542 26721 20576
rect 26755 20542 26791 20576
rect 26825 20542 26861 20576
rect 26895 20542 26952 20576
rect 26366 20505 26952 20542
rect 26366 20471 26371 20505
rect 26405 20471 26441 20505
rect 26475 20471 26511 20505
rect 26545 20471 26581 20505
rect 26615 20471 26651 20505
rect 26685 20471 26721 20505
rect 26755 20471 26791 20505
rect 26825 20471 26861 20505
rect 26895 20471 26952 20505
rect 26366 20434 26952 20471
rect 26366 20400 26371 20434
rect 26405 20400 26441 20434
rect 26475 20400 26511 20434
rect 26545 20400 26581 20434
rect 26615 20400 26651 20434
rect 26685 20400 26721 20434
rect 26755 20400 26791 20434
rect 26825 20400 26861 20434
rect 26895 20400 26952 20434
rect 26366 20363 26952 20400
rect 26366 20329 26371 20363
rect 26405 20329 26441 20363
rect 26475 20329 26511 20363
rect 26545 20329 26581 20363
rect 26615 20329 26651 20363
rect 26685 20329 26721 20363
rect 26755 20329 26791 20363
rect 26825 20329 26861 20363
rect 26895 20329 26952 20363
rect 26366 20292 26952 20329
rect 26366 20258 26371 20292
rect 26405 20258 26441 20292
rect 26475 20258 26511 20292
rect 26545 20258 26581 20292
rect 26615 20258 26651 20292
rect 26685 20258 26721 20292
rect 26755 20258 26791 20292
rect 26825 20258 26861 20292
rect 26895 20258 26952 20292
rect 26366 20221 26952 20258
rect 26366 20187 26371 20221
rect 26405 20187 26441 20221
rect 26475 20187 26511 20221
rect 26545 20187 26581 20221
rect 26615 20187 26651 20221
rect 26685 20187 26721 20221
rect 26755 20187 26791 20221
rect 26825 20187 26861 20221
rect 26895 20187 26952 20221
rect 26366 20150 26952 20187
rect 26366 20116 26371 20150
rect 26405 20116 26441 20150
rect 26475 20116 26511 20150
rect 26545 20116 26581 20150
rect 26615 20116 26651 20150
rect 26685 20116 26721 20150
rect 26755 20116 26791 20150
rect 26825 20116 26861 20150
rect 26895 20116 26952 20150
rect 26366 20078 26952 20116
rect 26366 20044 26371 20078
rect 26405 20044 26441 20078
rect 26475 20044 26511 20078
rect 26545 20044 26581 20078
rect 26615 20044 26651 20078
rect 26685 20044 26721 20078
rect 26755 20044 26791 20078
rect 26825 20044 26861 20078
rect 26895 20044 26952 20078
rect 26366 20010 26952 20044
rect 3484 19551 4095 19585
rect 3484 19517 3485 19551
rect 3519 19517 3561 19551
rect 3595 19517 3637 19551
rect 3671 19517 3713 19551
rect 3747 19517 3789 19551
rect 3823 19517 3865 19551
rect 3899 19517 3941 19551
rect 3975 19517 4017 19551
rect 4051 19517 4095 19551
rect 3484 19483 4095 19517
rect 3484 19449 3485 19483
rect 3519 19449 3561 19483
rect 3595 19449 3637 19483
rect 3671 19449 3713 19483
rect 3747 19449 3789 19483
rect 3823 19449 3865 19483
rect 3899 19449 3941 19483
rect 3975 19449 4017 19483
rect 4051 19449 4095 19483
rect 3484 19415 4095 19449
rect 3484 19381 3485 19415
rect 3519 19381 3561 19415
rect 3595 19381 3637 19415
rect 3671 19381 3713 19415
rect 3747 19381 3789 19415
rect 3823 19381 3865 19415
rect 3899 19381 3941 19415
rect 3975 19381 4017 19415
rect 4051 19381 4095 19415
rect 3484 19347 4095 19381
rect 3484 19313 3485 19347
rect 3519 19313 3561 19347
rect 3595 19313 3637 19347
rect 3671 19313 3713 19347
rect 3747 19313 3789 19347
rect 3823 19313 3865 19347
rect 3899 19313 3941 19347
rect 3975 19313 4017 19347
rect 4051 19313 4095 19347
rect 3484 19279 4095 19313
rect 3484 19245 3485 19279
rect 3519 19245 3561 19279
rect 3595 19245 3637 19279
rect 3671 19245 3713 19279
rect 3747 19245 3789 19279
rect 3823 19245 3865 19279
rect 3899 19245 3941 19279
rect 3975 19245 4017 19279
rect 4051 19245 4095 19279
rect 3484 19210 4095 19245
rect 3484 19176 3485 19210
rect 3519 19176 3561 19210
rect 3595 19176 3637 19210
rect 3671 19176 3713 19210
rect 3747 19176 3789 19210
rect 3823 19176 3865 19210
rect 3899 19176 3941 19210
rect 3975 19176 4017 19210
rect 4051 19176 4095 19210
rect 3484 19141 4095 19176
rect 3484 19107 3485 19141
rect 3519 19107 3561 19141
rect 3595 19107 3637 19141
rect 3671 19107 3713 19141
rect 3747 19107 3789 19141
rect 3823 19107 3865 19141
rect 3899 19107 3941 19141
rect 3975 19107 4017 19141
rect 4051 19107 4095 19141
rect 3484 19072 4095 19107
rect 3484 19038 3485 19072
rect 3519 19038 3561 19072
rect 3595 19038 3637 19072
rect 3671 19038 3713 19072
rect 3747 19038 3789 19072
rect 3823 19038 3865 19072
rect 3899 19038 3941 19072
rect 3975 19038 4017 19072
rect 4051 19038 4095 19072
rect 3484 19003 4095 19038
rect 3484 18969 3485 19003
rect 3519 18969 3561 19003
rect 3595 18969 3637 19003
rect 3671 18969 3713 19003
rect 3747 18969 3789 19003
rect 3823 18969 3865 19003
rect 3899 18969 3941 19003
rect 3975 18969 4017 19003
rect 4051 18969 4095 19003
rect 3484 18934 4095 18969
rect 3484 18900 3485 18934
rect 3519 18900 3561 18934
rect 3595 18900 3637 18934
rect 3671 18900 3713 18934
rect 3747 18900 3789 18934
rect 3823 18900 3865 18934
rect 3899 18900 3941 18934
rect 3975 18900 4017 18934
rect 4051 18900 4095 18934
rect 3484 18865 4095 18900
rect 3484 18831 3485 18865
rect 3519 18831 3561 18865
rect 3595 18831 3637 18865
rect 3671 18831 3713 18865
rect 3747 18831 3789 18865
rect 3823 18831 3865 18865
rect 3899 18831 3941 18865
rect 3975 18831 4017 18865
rect 4051 18831 4095 18865
rect 3484 18796 4095 18831
rect 3484 18762 3485 18796
rect 3519 18762 3561 18796
rect 3595 18762 3637 18796
rect 3671 18762 3713 18796
rect 3747 18762 3789 18796
rect 3823 18762 3865 18796
rect 3899 18762 3941 18796
rect 3975 18762 4017 18796
rect 4051 18762 4095 18796
rect 3484 18727 4095 18762
rect 3484 18693 3485 18727
rect 3519 18693 3561 18727
rect 3595 18693 3637 18727
rect 3671 18693 3713 18727
rect 3747 18693 3789 18727
rect 3823 18693 3865 18727
rect 3899 18693 3941 18727
rect 3975 18693 4017 18727
rect 4051 18693 4095 18727
rect 3484 18658 4095 18693
rect 3484 18624 3485 18658
rect 3519 18624 3561 18658
rect 3595 18624 3637 18658
rect 3671 18624 3713 18658
rect 3747 18624 3789 18658
rect 3823 18624 3865 18658
rect 3899 18624 3941 18658
rect 3975 18624 4017 18658
rect 4051 18624 4095 18658
rect 3484 18589 4095 18624
rect 3484 18555 3485 18589
rect 3519 18555 3561 18589
rect 3595 18555 3637 18589
rect 3671 18555 3713 18589
rect 3747 18555 3789 18589
rect 3823 18555 3865 18589
rect 3899 18555 3941 18589
rect 3975 18555 4017 18589
rect 4051 18555 4095 18589
rect 3484 18520 4095 18555
rect 3484 18486 3485 18520
rect 3519 18486 3561 18520
rect 3595 18486 3637 18520
rect 3671 18486 3713 18520
rect 3747 18486 3789 18520
rect 3823 18486 3865 18520
rect 3899 18486 3941 18520
rect 3975 18486 4017 18520
rect 4051 18486 4095 18520
rect 3484 18451 4095 18486
rect 3484 18417 3485 18451
rect 3519 18417 3561 18451
rect 3595 18417 3637 18451
rect 3671 18417 3713 18451
rect 3747 18417 3789 18451
rect 3823 18417 3865 18451
rect 3899 18417 3941 18451
rect 3975 18417 4017 18451
rect 4051 18417 4095 18451
rect 3484 18382 4095 18417
rect 3484 18348 3485 18382
rect 3519 18348 3561 18382
rect 3595 18348 3637 18382
rect 3671 18348 3713 18382
rect 3747 18348 3789 18382
rect 3823 18348 3865 18382
rect 3899 18348 3941 18382
rect 3975 18348 4017 18382
rect 4051 18348 4095 18382
rect 3484 18313 4095 18348
rect 3484 18279 3485 18313
rect 3519 18279 3561 18313
rect 3595 18279 3637 18313
rect 3671 18279 3713 18313
rect 3747 18279 3789 18313
rect 3823 18279 3865 18313
rect 3899 18279 3941 18313
rect 3975 18279 4017 18313
rect 4051 18279 4095 18313
rect 3484 18244 4095 18279
rect 3484 18210 3485 18244
rect 3519 18210 3561 18244
rect 3595 18210 3637 18244
rect 3671 18210 3713 18244
rect 3747 18210 3789 18244
rect 3823 18210 3865 18244
rect 3899 18210 3941 18244
rect 3975 18210 4017 18244
rect 4051 18210 4095 18244
rect 3484 18175 4095 18210
rect 3484 18141 3485 18175
rect 3519 18141 3561 18175
rect 3595 18141 3637 18175
rect 3671 18141 3713 18175
rect 3747 18141 3789 18175
rect 3823 18141 3865 18175
rect 3899 18141 3941 18175
rect 3975 18141 4017 18175
rect 4051 18141 4095 18175
rect 3484 18106 4095 18141
rect 3484 18072 3485 18106
rect 3519 18072 3561 18106
rect 3595 18072 3637 18106
rect 3671 18072 3713 18106
rect 3747 18072 3789 18106
rect 3823 18072 3865 18106
rect 3899 18072 3941 18106
rect 3975 18072 4017 18106
rect 4051 18072 4095 18106
rect 3484 18037 4095 18072
rect 3484 18003 3485 18037
rect 3519 18003 3561 18037
rect 3595 18003 3637 18037
rect 3671 18003 3713 18037
rect 3747 18003 3789 18037
rect 3823 18003 3865 18037
rect 3899 18003 3941 18037
rect 3975 18003 4017 18037
rect 4051 18003 4095 18037
rect 3484 17968 4095 18003
rect 3484 17934 3485 17968
rect 3519 17934 3561 17968
rect 3595 17934 3637 17968
rect 3671 17934 3713 17968
rect 3747 17934 3789 17968
rect 3823 17934 3865 17968
rect 3899 17934 3941 17968
rect 3975 17934 4017 17968
rect 4051 17934 4095 17968
rect 3484 17899 4095 17934
rect 3484 17865 3485 17899
rect 3519 17865 3561 17899
rect 3595 17865 3637 17899
rect 3671 17865 3713 17899
rect 3747 17865 3789 17899
rect 3823 17865 3865 17899
rect 3899 17865 3941 17899
rect 3975 17865 4017 17899
rect 4051 17865 4095 17899
rect 3484 17830 4095 17865
rect 3484 17796 3485 17830
rect 3519 17796 3561 17830
rect 3595 17796 3637 17830
rect 3671 17796 3713 17830
rect 3747 17796 3789 17830
rect 3823 17796 3865 17830
rect 3899 17796 3941 17830
rect 3975 17796 4017 17830
rect 4051 17796 4095 17830
rect 3484 17761 4095 17796
rect 3484 17727 3485 17761
rect 3519 17727 3561 17761
rect 3595 17727 3637 17761
rect 3671 17727 3713 17761
rect 3747 17727 3789 17761
rect 3823 17727 3865 17761
rect 3899 17727 3941 17761
rect 3975 17727 4017 17761
rect 4051 17727 4095 17761
rect 3484 17692 4095 17727
rect 3484 17658 3485 17692
rect 3519 17658 3561 17692
rect 3595 17658 3637 17692
rect 3671 17658 3713 17692
rect 3747 17658 3789 17692
rect 3823 17658 3865 17692
rect 3899 17658 3941 17692
rect 3975 17658 4017 17692
rect 4051 17658 4095 17692
rect 3484 17623 4095 17658
rect 3484 17589 3485 17623
rect 3519 17589 3561 17623
rect 3595 17589 3637 17623
rect 3671 17589 3713 17623
rect 3747 17589 3789 17623
rect 3823 17589 3865 17623
rect 3899 17589 3941 17623
rect 3975 17589 4017 17623
rect 4051 17589 4095 17623
rect 3484 17554 4095 17589
rect 3484 17520 3485 17554
rect 3519 17520 3561 17554
rect 3595 17520 3637 17554
rect 3671 17520 3713 17554
rect 3747 17520 3789 17554
rect 3823 17520 3865 17554
rect 3899 17520 3941 17554
rect 3975 17520 4017 17554
rect 4051 17520 4095 17554
rect 3484 17485 4095 17520
rect 3484 17451 3485 17485
rect 3519 17451 3561 17485
rect 3595 17451 3637 17485
rect 3671 17451 3713 17485
rect 3747 17451 3789 17485
rect 3823 17451 3865 17485
rect 3899 17451 3941 17485
rect 3975 17451 4017 17485
rect 4051 17451 4095 17485
rect 3484 17416 4095 17451
rect 3484 17382 3485 17416
rect 3519 17382 3561 17416
rect 3595 17382 3637 17416
rect 3671 17382 3713 17416
rect 3747 17382 3789 17416
rect 3823 17382 3865 17416
rect 3899 17382 3941 17416
rect 3975 17382 4017 17416
rect 4051 17382 4095 17416
rect 3484 17347 4095 17382
rect 3484 17313 3485 17347
rect 3519 17313 3561 17347
rect 3595 17313 3637 17347
rect 3671 17313 3713 17347
rect 3747 17313 3789 17347
rect 3823 17313 3865 17347
rect 3899 17313 3941 17347
rect 3975 17313 4017 17347
rect 4051 17313 4095 17347
rect 3484 17278 4095 17313
rect 3484 17244 3485 17278
rect 3519 17244 3561 17278
rect 3595 17244 3637 17278
rect 3671 17244 3713 17278
rect 3747 17244 3789 17278
rect 3823 17244 3865 17278
rect 3899 17244 3941 17278
rect 3975 17244 4017 17278
rect 4051 17244 4095 17278
rect 3484 17209 4095 17244
rect 3484 17175 3485 17209
rect 3519 17175 3561 17209
rect 3595 17175 3637 17209
rect 3671 17175 3713 17209
rect 3747 17175 3789 17209
rect 3823 17175 3865 17209
rect 3899 17175 3941 17209
rect 3975 17175 4017 17209
rect 4051 17175 4095 17209
rect 3484 17140 4095 17175
rect 3484 17106 3485 17140
rect 3519 17106 3561 17140
rect 3595 17106 3637 17140
rect 3671 17106 3713 17140
rect 3747 17106 3789 17140
rect 3823 17106 3865 17140
rect 3899 17106 3941 17140
rect 3975 17106 4017 17140
rect 4051 17106 4095 17140
rect 3484 17047 4095 17106
rect 3484 17013 3767 17047
rect 3801 17013 3835 17047
rect 3869 17013 3903 17047
rect 3937 17013 3971 17047
rect 4005 17013 4039 17047
rect 4073 17013 4095 17047
rect 3484 17006 4095 17013
rect 3701 16973 4095 17006
rect 3701 16939 3767 16973
rect 3801 16939 3835 16973
rect 3869 16939 3903 16973
rect 3937 16939 3971 16973
rect 4005 16939 4039 16973
rect 4073 16939 4095 16973
rect 3701 16899 4095 16939
rect 3701 16865 3767 16899
rect 3801 16865 3835 16899
rect 3869 16865 3903 16899
rect 3937 16865 3971 16899
rect 4005 16865 4039 16899
rect 4073 16865 4095 16899
rect 3701 16825 4095 16865
rect 3701 16791 3767 16825
rect 3801 16791 3835 16825
rect 3869 16791 3903 16825
rect 3937 16791 3971 16825
rect 4005 16791 4039 16825
rect 4073 16791 4095 16825
rect 3701 16751 4095 16791
rect 3701 16717 3767 16751
rect 3801 16717 3835 16751
rect 3869 16717 3903 16751
rect 3937 16717 3971 16751
rect 4005 16717 4039 16751
rect 4073 16717 4095 16751
rect 3701 16677 4095 16717
rect 3701 16643 3767 16677
rect 3801 16643 3835 16677
rect 3869 16643 3903 16677
rect 3937 16643 3971 16677
rect 4005 16643 4039 16677
rect 4073 16643 4095 16677
rect 3701 16603 4095 16643
rect 3701 16569 3767 16603
rect 3801 16569 3835 16603
rect 3869 16569 3903 16603
rect 3937 16569 3971 16603
rect 4005 16569 4039 16603
rect 4073 16569 4095 16603
rect 3701 16529 4095 16569
rect 3701 16495 3767 16529
rect 3801 16495 3835 16529
rect 3869 16495 3903 16529
rect 3937 16495 3971 16529
rect 4005 16495 4039 16529
rect 4073 16495 4095 16529
rect 3701 16455 4095 16495
rect 3701 16421 3767 16455
rect 3801 16421 3835 16455
rect 3869 16421 3903 16455
rect 3937 16421 3971 16455
rect 4005 16421 4039 16455
rect 4073 16421 4095 16455
rect 3701 16380 4095 16421
rect 3701 16360 3767 16380
rect 3484 16346 3767 16360
rect 3801 16346 3835 16380
rect 3869 16346 3903 16380
rect 3937 16346 3971 16380
rect 4005 16346 4039 16380
rect 4073 16346 4095 16380
rect 3484 16312 4095 16346
rect 3484 16294 3732 16312
rect 2950 16260 3732 16294
rect 2984 16226 3018 16260
rect 3052 16226 3086 16260
rect 3120 16226 3154 16260
rect 3188 16226 3222 16260
rect 3256 16226 3290 16260
rect 3324 16226 3358 16260
rect 3392 16226 3426 16260
rect 3460 16226 3494 16260
rect 3528 16226 3562 16260
rect 3596 16226 3630 16260
rect 3664 16226 3698 16260
rect 2950 16188 3732 16226
rect 2984 16154 3018 16188
rect 3052 16154 3086 16188
rect 3120 16154 3154 16188
rect 3188 16154 3222 16188
rect 3256 16154 3290 16188
rect 3324 16154 3358 16188
rect 3392 16154 3426 16188
rect 3460 16154 3494 16188
rect 3528 16154 3562 16188
rect 3596 16154 3630 16188
rect 3664 16154 3698 16188
rect 2950 16116 3732 16154
rect 2984 16082 3018 16116
rect 3052 16082 3086 16116
rect 3120 16082 3154 16116
rect 3188 16082 3222 16116
rect 3256 16082 3290 16116
rect 3324 16082 3358 16116
rect 3392 16082 3426 16116
rect 3460 16082 3494 16116
rect 3528 16082 3562 16116
rect 3596 16082 3630 16116
rect 3664 16082 3698 16116
rect 2950 16044 3732 16082
rect 2984 16010 3018 16044
rect 3052 16010 3086 16044
rect 3120 16010 3154 16044
rect 3188 16010 3222 16044
rect 3256 16010 3290 16044
rect 3324 16010 3358 16044
rect 3392 16010 3426 16044
rect 3460 16010 3494 16044
rect 3528 16010 3562 16044
rect 3596 16010 3630 16044
rect 3664 16010 3698 16044
rect 2950 15972 3732 16010
rect 2984 15938 3018 15972
rect 3052 15938 3086 15972
rect 3120 15938 3154 15972
rect 3188 15938 3222 15972
rect 3256 15938 3290 15972
rect 3324 15938 3358 15972
rect 3392 15938 3426 15972
rect 3460 15938 3494 15972
rect 3528 15938 3562 15972
rect 3596 15938 3630 15972
rect 3664 15938 3698 15972
rect 2950 15900 3732 15938
rect 2984 15866 3018 15900
rect 3052 15866 3086 15900
rect 3120 15866 3154 15900
rect 3188 15866 3222 15900
rect 3256 15866 3290 15900
rect 3324 15866 3358 15900
rect 3392 15866 3426 15900
rect 3460 15866 3494 15900
rect 3528 15866 3562 15900
rect 3596 15866 3630 15900
rect 3664 15866 3698 15900
rect 2950 15828 3732 15866
rect 2984 15794 3018 15828
rect 3052 15794 3086 15828
rect 3120 15794 3154 15828
rect 3188 15794 3222 15828
rect 3256 15794 3290 15828
rect 3324 15794 3358 15828
rect 3392 15794 3426 15828
rect 3460 15794 3494 15828
rect 3528 15794 3562 15828
rect 3596 15794 3630 15828
rect 3664 15794 3698 15828
rect 2950 15756 3732 15794
rect 2984 15722 3018 15756
rect 3052 15722 3086 15756
rect 3120 15722 3154 15756
rect 3188 15722 3222 15756
rect 3256 15722 3290 15756
rect 3324 15722 3358 15756
rect 3392 15722 3426 15756
rect 3460 15722 3494 15756
rect 3528 15722 3562 15756
rect 3596 15722 3630 15756
rect 3664 15722 3698 15756
rect 2950 15684 3732 15722
rect 2984 15650 3018 15684
rect 3052 15650 3086 15684
rect 3120 15650 3154 15684
rect 3188 15650 3222 15684
rect 3256 15650 3290 15684
rect 3324 15650 3358 15684
rect 3392 15650 3426 15684
rect 3460 15650 3494 15684
rect 3528 15650 3562 15684
rect 3596 15650 3630 15684
rect 3664 15650 3698 15684
rect 2950 15612 3732 15650
rect 2984 15578 3018 15612
rect 3052 15578 3086 15612
rect 3120 15578 3154 15612
rect 3188 15578 3222 15612
rect 3256 15578 3290 15612
rect 3324 15578 3358 15612
rect 3392 15578 3426 15612
rect 3460 15578 3494 15612
rect 3528 15578 3562 15612
rect 3596 15578 3630 15612
rect 3664 15578 3698 15612
rect 2950 15540 3732 15578
rect 2984 15506 3018 15540
rect 3052 15506 3086 15540
rect 3120 15506 3154 15540
rect 3188 15506 3222 15540
rect 3256 15506 3290 15540
rect 3324 15506 3358 15540
rect 3392 15506 3426 15540
rect 3460 15506 3494 15540
rect 3528 15506 3562 15540
rect 3596 15506 3630 15540
rect 3664 15506 3698 15540
rect 2950 15468 3732 15506
rect 2984 15434 3018 15468
rect 3052 15434 3086 15468
rect 3120 15434 3154 15468
rect 3188 15434 3222 15468
rect 3256 15434 3290 15468
rect 3324 15434 3358 15468
rect 3392 15434 3426 15468
rect 3460 15434 3494 15468
rect 3528 15434 3562 15468
rect 3596 15434 3630 15468
rect 3664 15434 3698 15468
rect 2950 15400 3732 15434
rect 7855 16278 8275 16312
rect 7855 16244 7858 16278
rect 7892 16244 7934 16278
rect 7968 16244 8010 16278
rect 8044 16244 8086 16278
rect 8120 16244 8162 16278
rect 8196 16244 8238 16278
rect 8272 16244 8275 16278
rect 7855 16209 8275 16244
rect 7855 16175 7858 16209
rect 7892 16175 7934 16209
rect 7968 16175 8010 16209
rect 8044 16175 8086 16209
rect 8120 16175 8162 16209
rect 8196 16175 8238 16209
rect 8272 16175 8275 16209
rect 7855 16140 8275 16175
rect 7855 16106 7858 16140
rect 7892 16106 7934 16140
rect 7968 16106 8010 16140
rect 8044 16106 8086 16140
rect 8120 16106 8162 16140
rect 8196 16106 8238 16140
rect 8272 16106 8275 16140
rect 7855 16071 8275 16106
rect 7855 16037 7858 16071
rect 7892 16037 7934 16071
rect 7968 16037 8010 16071
rect 8044 16037 8086 16071
rect 8120 16037 8162 16071
rect 8196 16037 8238 16071
rect 8272 16037 8275 16071
rect 7855 16002 8275 16037
rect 7855 15968 7858 16002
rect 7892 15968 7934 16002
rect 7968 15968 8010 16002
rect 8044 15968 8086 16002
rect 8120 15968 8162 16002
rect 8196 15968 8238 16002
rect 8272 15968 8275 16002
rect 7855 15933 8275 15968
rect 7855 15899 7858 15933
rect 7892 15899 7934 15933
rect 7968 15899 8010 15933
rect 8044 15899 8086 15933
rect 8120 15899 8162 15933
rect 8196 15899 8238 15933
rect 8272 15899 8275 15933
rect 7855 15864 8275 15899
rect 7855 15830 7858 15864
rect 7892 15830 7934 15864
rect 7968 15830 8010 15864
rect 8044 15830 8086 15864
rect 8120 15830 8162 15864
rect 8196 15830 8238 15864
rect 8272 15830 8275 15864
rect 7855 15795 8275 15830
rect 7855 15761 7858 15795
rect 7892 15761 7934 15795
rect 7968 15761 8010 15795
rect 8044 15761 8086 15795
rect 8120 15761 8162 15795
rect 8196 15761 8238 15795
rect 8272 15761 8275 15795
rect 7855 15726 8275 15761
rect 7855 15692 7858 15726
rect 7892 15692 7934 15726
rect 7968 15692 8010 15726
rect 8044 15692 8086 15726
rect 8120 15692 8162 15726
rect 8196 15692 8238 15726
rect 8272 15692 8275 15726
rect 7855 15657 8275 15692
rect 7855 15623 7858 15657
rect 7892 15623 7934 15657
rect 7968 15623 8010 15657
rect 8044 15623 8086 15657
rect 8120 15623 8162 15657
rect 8196 15623 8238 15657
rect 8272 15623 8275 15657
rect 7855 15588 8275 15623
rect 7855 15554 7858 15588
rect 7892 15554 7934 15588
rect 7968 15554 8010 15588
rect 8044 15554 8086 15588
rect 8120 15554 8162 15588
rect 8196 15554 8238 15588
rect 8272 15554 8275 15588
rect 7855 15519 8275 15554
rect 7855 15485 7858 15519
rect 7892 15485 7934 15519
rect 7968 15485 8010 15519
rect 8044 15485 8086 15519
rect 8120 15485 8162 15519
rect 8196 15485 8238 15519
rect 8272 15485 8275 15519
rect 7855 15449 8275 15485
rect 7855 15415 7858 15449
rect 7892 15415 7934 15449
rect 7968 15415 8010 15449
rect 8044 15415 8086 15449
rect 8120 15415 8162 15449
rect 8196 15415 8238 15449
rect 8272 15415 8275 15449
rect 7855 15381 8275 15415
<< psubdiffcont >>
rect 76 39866 110 39900
rect 198 39866 232 39900
rect 76 39797 110 39831
rect 198 39797 232 39831
rect 76 39728 110 39762
rect 198 39728 232 39762
rect 76 39659 110 39693
rect 198 39659 232 39693
rect 76 39590 110 39624
rect 198 39590 232 39624
rect 76 39521 110 39555
rect 198 39521 232 39555
rect 76 39452 110 39486
rect 198 39452 232 39486
rect 76 39383 110 39417
rect 198 39383 232 39417
rect 76 39314 110 39348
rect 198 39314 232 39348
rect 76 39245 110 39279
rect 198 39245 232 39279
rect 76 39175 110 39209
rect 198 39175 232 39209
rect 76 39105 110 39139
rect 198 39105 232 39139
rect 76 39035 110 39069
rect 198 39035 232 39069
rect 76 38965 110 38999
rect 198 38965 232 38999
rect 76 38895 110 38929
rect 198 38895 232 38929
rect 76 38825 110 38859
rect 198 38825 232 38859
rect 76 38755 110 38789
rect 198 38755 232 38789
rect 76 38685 110 38719
rect 198 38685 232 38719
rect 76 38615 110 38649
rect 198 38615 232 38649
rect 76 38545 110 38579
rect 198 38545 232 38579
rect 76 38475 110 38509
rect 198 38475 232 38509
rect 76 38405 110 38439
rect 198 38405 232 38439
rect 76 38335 110 38369
rect 198 38335 232 38369
rect 76 38265 110 38299
rect 198 38265 232 38299
rect 76 38195 110 38229
rect 198 38195 232 38229
rect 76 38125 110 38159
rect 198 38125 232 38159
rect 76 38055 110 38089
rect 198 38055 232 38089
rect 233 12914 267 12948
rect 301 12914 335 12948
rect 369 12914 403 12948
rect 437 12914 471 12948
rect 505 12914 539 12948
rect 573 12914 607 12948
rect 641 12914 675 12948
rect 709 12914 743 12948
rect 777 12914 811 12948
rect 845 12914 879 12948
rect 913 12914 947 12948
rect 981 12914 1015 12948
rect 1049 12914 1083 12948
rect 1117 12914 1151 12948
rect 1185 12914 1219 12948
rect 233 12843 267 12877
rect 301 12843 335 12877
rect 369 12843 403 12877
rect 437 12843 471 12877
rect 505 12843 539 12877
rect 573 12843 607 12877
rect 641 12843 675 12877
rect 709 12843 743 12877
rect 777 12843 811 12877
rect 845 12843 879 12877
rect 913 12843 947 12877
rect 981 12843 1015 12877
rect 1049 12843 1083 12877
rect 1117 12843 1151 12877
rect 1185 12843 1219 12877
rect 233 12772 267 12806
rect 301 12772 335 12806
rect 369 12772 403 12806
rect 437 12772 471 12806
rect 505 12772 539 12806
rect 573 12772 607 12806
rect 641 12772 675 12806
rect 709 12772 743 12806
rect 777 12772 811 12806
rect 845 12772 879 12806
rect 913 12772 947 12806
rect 981 12772 1015 12806
rect 1049 12772 1083 12806
rect 1117 12772 1151 12806
rect 1185 12772 1219 12806
rect 233 12701 267 12735
rect 301 12701 335 12735
rect 369 12701 403 12735
rect 437 12701 471 12735
rect 505 12701 539 12735
rect 573 12701 607 12735
rect 641 12701 675 12735
rect 709 12701 743 12735
rect 777 12701 811 12735
rect 845 12701 879 12735
rect 913 12701 947 12735
rect 981 12701 1015 12735
rect 1049 12701 1083 12735
rect 1117 12701 1151 12735
rect 1185 12701 1219 12735
rect 233 12630 267 12664
rect 301 12630 335 12664
rect 369 12630 403 12664
rect 437 12630 471 12664
rect 505 12630 539 12664
rect 573 12630 607 12664
rect 641 12630 675 12664
rect 709 12630 743 12664
rect 777 12630 811 12664
rect 845 12630 879 12664
rect 913 12630 947 12664
rect 981 12630 1015 12664
rect 1049 12630 1083 12664
rect 1117 12630 1151 12664
rect 1185 12630 1219 12664
rect 233 12559 267 12593
rect 301 12559 335 12593
rect 369 12559 403 12593
rect 437 12559 471 12593
rect 505 12559 539 12593
rect 573 12559 607 12593
rect 641 12559 675 12593
rect 709 12559 743 12593
rect 777 12559 811 12593
rect 845 12559 879 12593
rect 913 12559 947 12593
rect 981 12559 1015 12593
rect 1049 12559 1083 12593
rect 1117 12559 1151 12593
rect 1185 12559 1219 12593
rect 233 12488 267 12522
rect 301 12488 335 12522
rect 369 12488 403 12522
rect 437 12488 471 12522
rect 505 12488 539 12522
rect 573 12488 607 12522
rect 641 12488 675 12522
rect 709 12488 743 12522
rect 777 12488 811 12522
rect 845 12488 879 12522
rect 913 12488 947 12522
rect 981 12488 1015 12522
rect 1049 12488 1083 12522
rect 1117 12488 1151 12522
rect 1185 12488 1219 12522
rect 233 12417 267 12451
rect 301 12417 335 12451
rect 369 12417 403 12451
rect 437 12417 471 12451
rect 505 12417 539 12451
rect 573 12417 607 12451
rect 641 12417 675 12451
rect 709 12417 743 12451
rect 777 12417 811 12451
rect 845 12417 879 12451
rect 913 12417 947 12451
rect 981 12417 1015 12451
rect 1049 12417 1083 12451
rect 1117 12417 1151 12451
rect 1185 12417 1219 12451
rect 233 12346 267 12380
rect 301 12346 335 12380
rect 369 12346 403 12380
rect 437 12346 471 12380
rect 505 12346 539 12380
rect 573 12346 607 12380
rect 641 12346 675 12380
rect 709 12346 743 12380
rect 777 12346 811 12380
rect 845 12346 879 12380
rect 913 12346 947 12380
rect 981 12346 1015 12380
rect 1049 12346 1083 12380
rect 1117 12346 1151 12380
rect 1185 12346 1219 12380
rect 233 12275 267 12309
rect 301 12275 335 12309
rect 369 12275 403 12309
rect 437 12275 471 12309
rect 505 12275 539 12309
rect 573 12275 607 12309
rect 641 12275 675 12309
rect 709 12275 743 12309
rect 777 12275 811 12309
rect 845 12275 879 12309
rect 913 12275 947 12309
rect 981 12275 1015 12309
rect 1049 12275 1083 12309
rect 1117 12275 1151 12309
rect 1185 12275 1219 12309
rect 233 12204 267 12238
rect 301 12204 335 12238
rect 369 12204 403 12238
rect 437 12204 471 12238
rect 505 12204 539 12238
rect 573 12204 607 12238
rect 641 12204 675 12238
rect 709 12204 743 12238
rect 777 12204 811 12238
rect 845 12204 879 12238
rect 913 12204 947 12238
rect 981 12204 1015 12238
rect 1049 12204 1083 12238
rect 1117 12204 1151 12238
rect 1185 12204 1219 12238
rect 233 12133 267 12167
rect 301 12133 335 12167
rect 369 12133 403 12167
rect 437 12133 471 12167
rect 505 12133 539 12167
rect 573 12133 607 12167
rect 641 12133 675 12167
rect 709 12133 743 12167
rect 777 12133 811 12167
rect 845 12133 879 12167
rect 913 12133 947 12167
rect 981 12133 1015 12167
rect 1049 12133 1083 12167
rect 1117 12133 1151 12167
rect 1185 12133 1219 12167
rect 233 12062 267 12096
rect 301 12062 335 12096
rect 369 12062 403 12096
rect 437 12062 471 12096
rect 505 12062 539 12096
rect 573 12062 607 12096
rect 641 12062 675 12096
rect 709 12062 743 12096
rect 777 12062 811 12096
rect 845 12062 879 12096
rect 913 12062 947 12096
rect 981 12062 1015 12096
rect 1049 12062 1083 12096
rect 1117 12062 1151 12096
rect 1185 12062 1219 12096
rect 233 11991 267 12025
rect 301 11991 335 12025
rect 369 11991 403 12025
rect 437 11991 471 12025
rect 505 11991 539 12025
rect 573 11991 607 12025
rect 641 11991 675 12025
rect 709 11991 743 12025
rect 777 11991 811 12025
rect 845 11991 879 12025
rect 913 11991 947 12025
rect 981 11991 1015 12025
rect 1049 11991 1083 12025
rect 1117 11991 1151 12025
rect 1185 11991 1219 12025
rect 233 11920 267 11954
rect 301 11920 335 11954
rect 369 11920 403 11954
rect 437 11920 471 11954
rect 505 11920 539 11954
rect 573 11920 607 11954
rect 641 11920 675 11954
rect 709 11920 743 11954
rect 777 11920 811 11954
rect 845 11920 879 11954
rect 913 11920 947 11954
rect 981 11920 1015 11954
rect 1049 11920 1083 11954
rect 1117 11920 1151 11954
rect 1185 11920 1219 11954
rect 233 11849 267 11883
rect 301 11849 335 11883
rect 369 11849 403 11883
rect 437 11849 471 11883
rect 505 11849 539 11883
rect 573 11849 607 11883
rect 641 11849 675 11883
rect 709 11849 743 11883
rect 777 11849 811 11883
rect 845 11849 879 11883
rect 913 11849 947 11883
rect 981 11849 1015 11883
rect 1049 11849 1083 11883
rect 1117 11849 1151 11883
rect 1185 11849 1219 11883
rect 233 11778 267 11812
rect 301 11778 335 11812
rect 369 11778 403 11812
rect 437 11778 471 11812
rect 505 11778 539 11812
rect 573 11778 607 11812
rect 641 11778 675 11812
rect 709 11778 743 11812
rect 777 11778 811 11812
rect 845 11778 879 11812
rect 913 11778 947 11812
rect 981 11778 1015 11812
rect 1049 11778 1083 11812
rect 1117 11778 1151 11812
rect 1185 11778 1219 11812
rect 233 11707 267 11741
rect 301 11707 335 11741
rect 369 11707 403 11741
rect 437 11707 471 11741
rect 505 11707 539 11741
rect 573 11707 607 11741
rect 641 11707 675 11741
rect 709 11707 743 11741
rect 777 11707 811 11741
rect 845 11707 879 11741
rect 913 11707 947 11741
rect 981 11707 1015 11741
rect 1049 11707 1083 11741
rect 1117 11707 1151 11741
rect 1185 11707 1219 11741
rect 233 11636 267 11670
rect 301 11636 335 11670
rect 369 11636 403 11670
rect 437 11636 471 11670
rect 505 11636 539 11670
rect 573 11636 607 11670
rect 641 11636 675 11670
rect 709 11636 743 11670
rect 777 11636 811 11670
rect 845 11636 879 11670
rect 913 11636 947 11670
rect 981 11636 1015 11670
rect 1049 11636 1083 11670
rect 1117 11636 1151 11670
rect 1185 11636 1219 11670
rect 233 11564 267 11598
rect 301 11564 335 11598
rect 369 11564 403 11598
rect 437 11564 471 11598
rect 505 11564 539 11598
rect 573 11564 607 11598
rect 641 11564 675 11598
rect 709 11564 743 11598
rect 777 11564 811 11598
rect 845 11564 879 11598
rect 913 11564 947 11598
rect 981 11564 1015 11598
rect 1049 11564 1083 11598
rect 1117 11564 1151 11598
rect 1185 11564 1219 11598
rect 233 11492 267 11526
rect 301 11492 335 11526
rect 369 11492 403 11526
rect 437 11492 471 11526
rect 505 11492 539 11526
rect 573 11492 607 11526
rect 641 11492 675 11526
rect 709 11492 743 11526
rect 777 11492 811 11526
rect 845 11492 879 11526
rect 913 11492 947 11526
rect 981 11492 1015 11526
rect 1049 11492 1083 11526
rect 1117 11492 1151 11526
rect 1185 11492 1219 11526
rect 16319 11028 16353 11062
rect 16388 11028 16422 11062
rect 16457 11028 16491 11062
rect 16526 11028 16560 11062
rect 16594 11028 16628 11062
rect 16662 11028 16696 11062
rect 16730 11028 16764 11062
rect 16798 11028 16832 11062
rect 16866 11028 16900 11062
rect 16934 11028 16968 11062
rect 17002 11028 17036 11062
rect 17070 11028 17104 11062
rect 17138 11028 17172 11062
rect 17206 11028 17240 11062
rect 17274 11028 17308 11062
rect 17342 11028 17376 11062
rect 17410 11028 17444 11062
rect 17478 11028 17512 11062
rect 17546 11028 17580 11062
rect 17614 11028 17648 11062
rect 17682 11028 17716 11062
rect 17750 11028 17784 11062
rect 17818 11028 17852 11062
rect 17886 11028 17920 11062
rect 17954 11028 17988 11062
rect 18022 11028 18056 11062
rect 18090 11028 18124 11062
rect 18158 11028 18192 11062
rect 18226 11028 18260 11062
rect 18294 11028 18328 11062
rect 18362 11028 18396 11062
rect 18430 11028 18464 11062
rect 18498 11028 18532 11062
rect 18566 11028 18600 11062
rect 18634 11028 18668 11062
rect 18702 11028 18736 11062
rect 18770 11028 18804 11062
rect 18838 11028 18872 11062
rect 18906 11028 18940 11062
rect 18974 11028 19008 11062
rect 19042 11028 19076 11062
rect 19110 11028 19144 11062
rect 19178 11028 19212 11062
rect 19246 11028 19280 11062
rect 19314 11028 19348 11062
rect 19548 11002 19582 11036
rect 19616 11002 19650 11036
rect 19548 10899 19582 10933
rect 19616 10899 19650 10933
rect 19548 10796 19582 10830
rect 19616 10796 19650 10830
rect 19548 10693 19582 10727
rect 19616 10693 19650 10727
rect 19548 10589 19582 10623
rect 19616 10589 19650 10623
rect 19548 10485 19582 10519
rect 19616 10485 19650 10519
rect 19548 10381 19582 10415
rect 19616 10381 19650 10415
rect 16563 10221 16597 10255
rect 16631 10221 16665 10255
rect 16699 10221 16733 10255
rect 16767 10221 16801 10255
rect 16563 10148 16597 10182
rect 16631 10148 16665 10182
rect 16699 10148 16733 10182
rect 16767 10148 16801 10182
rect 16563 10075 16597 10109
rect 16631 10075 16665 10109
rect 16699 10075 16733 10109
rect 16767 10075 16801 10109
rect 16563 10002 16597 10036
rect 16631 10002 16665 10036
rect 16699 10002 16733 10036
rect 16767 10002 16801 10036
rect 16563 9928 16597 9962
rect 16631 9928 16665 9962
rect 16699 9928 16733 9962
rect 16767 9928 16801 9962
rect 16563 9854 16597 9888
rect 16631 9854 16665 9888
rect 16699 9854 16733 9888
rect 16767 9854 16801 9888
rect 19548 10277 19582 10311
rect 19616 10277 19650 10311
rect 19548 10173 19582 10207
rect 19616 10173 19650 10207
rect 19548 10069 19582 10103
rect 19616 10069 19650 10103
rect 19548 9965 19582 9999
rect 19616 9965 19650 9999
rect 19548 9861 19582 9895
rect 19616 9861 19650 9895
rect 16563 9780 16597 9814
rect 16631 9780 16665 9814
rect 16699 9780 16733 9814
rect 16767 9780 16801 9814
rect 16563 9706 16597 9740
rect 16631 9706 16665 9740
rect 16699 9706 16733 9740
rect 16767 9706 16801 9740
rect 16563 9632 16597 9666
rect 16631 9632 16665 9666
rect 16699 9632 16733 9666
rect 16767 9632 16801 9666
rect 16563 9558 16597 9592
rect 16631 9558 16665 9592
rect 16699 9558 16733 9592
rect 16767 9558 16801 9592
rect 23590 8972 23624 9006
<< mvpsubdiffcont >>
rect 24093 37640 24127 37674
rect 24162 37640 24196 37674
rect 24231 37640 24265 37674
rect 24300 37640 24334 37674
rect 24369 37640 24403 37674
rect 24438 37640 24472 37674
rect 24507 37640 24541 37674
rect 24576 37640 24610 37674
rect 24645 37640 24679 37674
rect 24714 37640 24748 37674
rect 24783 37640 24817 37674
rect 24852 37640 24886 37674
rect 24921 37640 24955 37674
rect 24990 37640 25024 37674
rect 25059 37640 25093 37674
rect 25127 37640 25161 37674
rect 25195 37640 25229 37674
rect 25263 37640 25297 37674
rect 25331 37640 25365 37674
rect 25399 37640 25433 37674
rect 25467 37640 25501 37674
rect 25535 37640 25569 37674
rect 25603 37640 25637 37674
rect 25671 37640 25705 37674
rect 25739 37640 25773 37674
rect 25807 37640 25841 37674
rect 25875 37640 25909 37674
rect 25943 37640 25977 37674
rect 26011 37640 26045 37674
rect 26079 37640 26113 37674
rect 26147 37640 26181 37674
rect 26215 37640 26249 37674
rect 26283 37640 26317 37674
rect 26351 37640 26385 37674
rect 26419 37640 26453 37674
rect 26487 37640 26521 37674
rect 26555 37640 26589 37674
rect 26623 37640 26657 37674
rect 26691 37640 26725 37674
rect 26759 37640 26793 37674
rect 26827 37640 26861 37674
rect 26895 37640 26929 37674
rect 26963 37640 26997 37674
rect 24093 37562 24127 37596
rect 24162 37562 24196 37596
rect 24231 37562 24265 37596
rect 24300 37562 24334 37596
rect 24369 37562 24403 37596
rect 24438 37562 24472 37596
rect 24507 37562 24541 37596
rect 24576 37562 24610 37596
rect 24645 37562 24679 37596
rect 24714 37562 24748 37596
rect 24783 37562 24817 37596
rect 24852 37562 24886 37596
rect 24921 37562 24955 37596
rect 24990 37562 25024 37596
rect 25059 37562 25093 37596
rect 25127 37562 25161 37596
rect 25195 37562 25229 37596
rect 25263 37562 25297 37596
rect 25331 37562 25365 37596
rect 25399 37562 25433 37596
rect 25467 37562 25501 37596
rect 25535 37562 25569 37596
rect 25603 37562 25637 37596
rect 25671 37562 25705 37596
rect 25739 37562 25773 37596
rect 25807 37562 25841 37596
rect 25875 37562 25909 37596
rect 25943 37562 25977 37596
rect 26011 37562 26045 37596
rect 26079 37562 26113 37596
rect 26147 37562 26181 37596
rect 26215 37562 26249 37596
rect 26283 37562 26317 37596
rect 26351 37562 26385 37596
rect 26419 37562 26453 37596
rect 26487 37562 26521 37596
rect 26555 37562 26589 37596
rect 26623 37562 26657 37596
rect 26691 37562 26725 37596
rect 26759 37562 26793 37596
rect 26827 37562 26861 37596
rect 26895 37562 26929 37596
rect 26963 37562 26997 37596
rect 219 37450 253 37484
rect 305 37450 339 37484
rect 219 37381 253 37415
rect 305 37381 339 37415
rect 219 37312 253 37346
rect 305 37312 339 37346
rect 219 37243 253 37277
rect 305 37243 339 37277
rect 219 37174 253 37208
rect 305 37174 339 37208
rect 219 37105 253 37139
rect 305 37105 339 37139
rect 219 37036 253 37070
rect 305 37036 339 37070
rect 219 36967 253 37001
rect 305 36967 339 37001
rect 219 36898 253 36932
rect 305 36898 339 36932
rect 219 36829 253 36863
rect 305 36829 339 36863
rect 219 36760 253 36794
rect 305 36760 339 36794
rect 219 36691 253 36725
rect 305 36691 339 36725
rect 219 36621 253 36655
rect 305 36621 339 36655
rect 219 36551 253 36585
rect 305 36551 339 36585
rect 219 36481 253 36515
rect 305 36481 339 36515
rect 219 36411 253 36445
rect 305 36411 339 36445
rect 219 36341 253 36375
rect 305 36341 339 36375
rect 219 36271 253 36305
rect 305 36271 339 36305
rect 219 36201 253 36235
rect 305 36201 339 36235
rect 219 36131 253 36165
rect 305 36131 339 36165
rect 219 36061 253 36095
rect 305 36061 339 36095
rect 219 35991 253 36025
rect 305 35991 339 36025
rect 278 35857 312 35891
rect 278 35789 312 35823
rect 278 35721 312 35755
rect 278 35653 312 35687
rect 278 35585 312 35619
rect 278 35517 312 35551
rect 278 35449 312 35483
rect 278 35381 312 35415
rect 278 35313 312 35347
rect 278 35245 312 35279
rect 278 35177 312 35211
rect 278 35109 312 35143
rect 278 35041 312 35075
rect 278 34972 312 35006
rect 278 34903 312 34937
rect 278 34834 312 34868
rect 278 34765 312 34799
rect 278 34696 312 34730
rect 278 34627 312 34661
rect 278 34558 312 34592
rect 278 34489 312 34523
rect 278 34420 312 34454
rect 278 34351 312 34385
rect 278 34282 312 34316
rect 278 34213 312 34247
rect 278 34144 312 34178
rect 278 34075 312 34109
rect 278 34006 312 34040
rect 278 33937 312 33971
rect 278 33868 312 33902
rect 278 33799 312 33833
rect 278 33730 312 33764
rect 278 33661 312 33695
rect 278 33592 312 33626
rect 278 33523 312 33557
rect 278 33454 312 33488
rect 278 33385 312 33419
rect 278 33316 312 33350
rect 22827 37483 22861 37517
rect 22897 37483 22931 37517
rect 22967 37483 23001 37517
rect 23037 37483 23071 37517
rect 23107 37483 23141 37517
rect 23177 37483 23211 37517
rect 23247 37483 23281 37517
rect 23317 37483 23351 37517
rect 23387 37483 23421 37517
rect 23457 37483 23491 37517
rect 23527 37483 23561 37517
rect 23597 37483 23631 37517
rect 23711 37506 23745 37540
rect 23794 37506 23828 37540
rect 23877 37506 23911 37540
rect 23959 37506 23993 37540
rect 24093 37484 24127 37518
rect 24162 37484 24196 37518
rect 24231 37484 24265 37518
rect 24300 37484 24334 37518
rect 24369 37484 24403 37518
rect 24438 37484 24472 37518
rect 24507 37484 24541 37518
rect 24576 37484 24610 37518
rect 24645 37484 24679 37518
rect 24714 37484 24748 37518
rect 24783 37484 24817 37518
rect 24852 37484 24886 37518
rect 24921 37484 24955 37518
rect 24990 37484 25024 37518
rect 25059 37484 25093 37518
rect 25127 37484 25161 37518
rect 25195 37484 25229 37518
rect 25263 37484 25297 37518
rect 25331 37484 25365 37518
rect 25399 37484 25433 37518
rect 25467 37484 25501 37518
rect 25535 37484 25569 37518
rect 25603 37484 25637 37518
rect 25671 37484 25705 37518
rect 25739 37484 25773 37518
rect 25807 37484 25841 37518
rect 25875 37484 25909 37518
rect 25943 37484 25977 37518
rect 26011 37484 26045 37518
rect 26079 37484 26113 37518
rect 26147 37484 26181 37518
rect 26215 37484 26249 37518
rect 26283 37484 26317 37518
rect 26351 37484 26385 37518
rect 26419 37484 26453 37518
rect 26487 37484 26521 37518
rect 26555 37484 26589 37518
rect 26623 37484 26657 37518
rect 26691 37484 26725 37518
rect 26759 37484 26793 37518
rect 26827 37484 26861 37518
rect 26895 37484 26929 37518
rect 26963 37484 26997 37518
rect 22827 37415 22861 37449
rect 22897 37415 22931 37449
rect 22967 37415 23001 37449
rect 23037 37415 23071 37449
rect 23107 37415 23141 37449
rect 23177 37415 23211 37449
rect 23247 37415 23281 37449
rect 23317 37415 23351 37449
rect 23387 37415 23421 37449
rect 23457 37415 23491 37449
rect 23527 37415 23561 37449
rect 23597 37415 23631 37449
rect 23711 37420 23745 37454
rect 23794 37420 23828 37454
rect 23877 37420 23911 37454
rect 23959 37420 23993 37454
rect 24093 37406 24127 37440
rect 24162 37406 24196 37440
rect 24231 37406 24265 37440
rect 24300 37406 24334 37440
rect 24369 37406 24403 37440
rect 24438 37406 24472 37440
rect 24507 37406 24541 37440
rect 24576 37406 24610 37440
rect 24645 37406 24679 37440
rect 24714 37406 24748 37440
rect 24783 37406 24817 37440
rect 24852 37406 24886 37440
rect 24921 37406 24955 37440
rect 24990 37406 25024 37440
rect 25059 37406 25093 37440
rect 25127 37406 25161 37440
rect 25195 37406 25229 37440
rect 25263 37406 25297 37440
rect 25331 37406 25365 37440
rect 25399 37406 25433 37440
rect 25467 37406 25501 37440
rect 25535 37406 25569 37440
rect 25603 37406 25637 37440
rect 25671 37406 25705 37440
rect 25739 37406 25773 37440
rect 25807 37406 25841 37440
rect 25875 37406 25909 37440
rect 25943 37406 25977 37440
rect 26011 37406 26045 37440
rect 26079 37406 26113 37440
rect 26147 37406 26181 37440
rect 26215 37406 26249 37440
rect 26283 37406 26317 37440
rect 26351 37406 26385 37440
rect 26419 37406 26453 37440
rect 26487 37406 26521 37440
rect 26555 37406 26589 37440
rect 26623 37406 26657 37440
rect 26691 37406 26725 37440
rect 26759 37406 26793 37440
rect 26827 37406 26861 37440
rect 26895 37406 26929 37440
rect 26963 37406 26997 37440
rect 22827 37347 22861 37381
rect 22897 37347 22931 37381
rect 22967 37347 23001 37381
rect 23037 37347 23071 37381
rect 23107 37347 23141 37381
rect 23177 37347 23211 37381
rect 23247 37347 23281 37381
rect 23317 37347 23351 37381
rect 23387 37347 23421 37381
rect 23457 37347 23491 37381
rect 23527 37347 23561 37381
rect 23597 37347 23631 37381
rect 23711 37334 23745 37368
rect 23794 37334 23828 37368
rect 23877 37334 23911 37368
rect 23959 37334 23993 37368
rect 24093 37328 24127 37362
rect 24162 37328 24196 37362
rect 24231 37328 24265 37362
rect 24300 37328 24334 37362
rect 24369 37328 24403 37362
rect 24438 37328 24472 37362
rect 24507 37328 24541 37362
rect 24576 37328 24610 37362
rect 24645 37328 24679 37362
rect 24714 37328 24748 37362
rect 24783 37328 24817 37362
rect 24852 37328 24886 37362
rect 24921 37328 24955 37362
rect 24990 37328 25024 37362
rect 25059 37328 25093 37362
rect 25127 37328 25161 37362
rect 25195 37328 25229 37362
rect 25263 37328 25297 37362
rect 25331 37328 25365 37362
rect 25399 37328 25433 37362
rect 25467 37328 25501 37362
rect 25535 37328 25569 37362
rect 25603 37328 25637 37362
rect 25671 37328 25705 37362
rect 25739 37328 25773 37362
rect 25807 37328 25841 37362
rect 25875 37328 25909 37362
rect 25943 37328 25977 37362
rect 26011 37328 26045 37362
rect 26079 37328 26113 37362
rect 26147 37328 26181 37362
rect 26215 37328 26249 37362
rect 26283 37328 26317 37362
rect 26351 37328 26385 37362
rect 26419 37328 26453 37362
rect 26487 37328 26521 37362
rect 26555 37328 26589 37362
rect 26623 37328 26657 37362
rect 26691 37328 26725 37362
rect 26759 37328 26793 37362
rect 26827 37328 26861 37362
rect 26895 37328 26929 37362
rect 26963 37328 26997 37362
rect 22827 37279 22861 37313
rect 22897 37279 22931 37313
rect 22967 37279 23001 37313
rect 23037 37279 23071 37313
rect 23107 37279 23141 37313
rect 23177 37279 23211 37313
rect 23247 37279 23281 37313
rect 23317 37279 23351 37313
rect 23387 37279 23421 37313
rect 23457 37279 23491 37313
rect 23527 37279 23561 37313
rect 23597 37279 23631 37313
rect 23711 37248 23745 37282
rect 23794 37248 23828 37282
rect 23877 37248 23911 37282
rect 23959 37248 23993 37282
rect 24093 37250 24127 37284
rect 24162 37250 24196 37284
rect 24231 37250 24265 37284
rect 24300 37250 24334 37284
rect 24369 37250 24403 37284
rect 24438 37250 24472 37284
rect 24507 37250 24541 37284
rect 24576 37250 24610 37284
rect 24645 37250 24679 37284
rect 24714 37250 24748 37284
rect 24783 37250 24817 37284
rect 24852 37250 24886 37284
rect 24921 37250 24955 37284
rect 24990 37250 25024 37284
rect 25059 37250 25093 37284
rect 25127 37250 25161 37284
rect 25195 37250 25229 37284
rect 25263 37250 25297 37284
rect 25331 37250 25365 37284
rect 25399 37250 25433 37284
rect 25467 37250 25501 37284
rect 25535 37250 25569 37284
rect 25603 37250 25637 37284
rect 25671 37250 25705 37284
rect 25739 37250 25773 37284
rect 25807 37250 25841 37284
rect 25875 37250 25909 37284
rect 25943 37250 25977 37284
rect 26011 37250 26045 37284
rect 26079 37250 26113 37284
rect 26147 37250 26181 37284
rect 26215 37250 26249 37284
rect 26283 37250 26317 37284
rect 26351 37250 26385 37284
rect 26419 37250 26453 37284
rect 26487 37250 26521 37284
rect 26555 37250 26589 37284
rect 26623 37250 26657 37284
rect 26691 37250 26725 37284
rect 26759 37250 26793 37284
rect 26827 37250 26861 37284
rect 26895 37250 26929 37284
rect 26963 37250 26997 37284
rect 22827 37211 22861 37245
rect 22897 37211 22931 37245
rect 22967 37211 23001 37245
rect 23037 37211 23071 37245
rect 23107 37211 23141 37245
rect 23177 37211 23211 37245
rect 23247 37211 23281 37245
rect 23317 37211 23351 37245
rect 23387 37211 23421 37245
rect 23457 37211 23491 37245
rect 23527 37211 23561 37245
rect 23597 37211 23631 37245
rect 22827 37143 22861 37177
rect 22897 37143 22931 37177
rect 22967 37143 23001 37177
rect 23037 37143 23071 37177
rect 23107 37143 23141 37177
rect 23177 37143 23211 37177
rect 23247 37143 23281 37177
rect 23317 37143 23351 37177
rect 23387 37143 23421 37177
rect 23457 37143 23491 37177
rect 23527 37143 23561 37177
rect 23597 37143 23631 37177
rect 22827 37075 22861 37109
rect 22897 37075 22931 37109
rect 22967 37075 23001 37109
rect 23037 37075 23071 37109
rect 23107 37075 23141 37109
rect 23177 37075 23211 37109
rect 23247 37075 23281 37109
rect 23317 37075 23351 37109
rect 23387 37075 23421 37109
rect 23457 37075 23491 37109
rect 23527 37075 23561 37109
rect 23597 37075 23631 37109
rect 22827 37007 22861 37041
rect 22897 37007 22931 37041
rect 22967 37007 23001 37041
rect 23037 37007 23071 37041
rect 23107 37007 23141 37041
rect 23177 37007 23211 37041
rect 23247 37007 23281 37041
rect 23317 37007 23351 37041
rect 23387 37007 23421 37041
rect 23457 37007 23491 37041
rect 23527 37007 23561 37041
rect 23597 37007 23631 37041
rect 22827 36939 22861 36973
rect 22897 36939 22931 36973
rect 22967 36939 23001 36973
rect 23037 36939 23071 36973
rect 23107 36939 23141 36973
rect 23177 36939 23211 36973
rect 23247 36939 23281 36973
rect 23317 36939 23351 36973
rect 23387 36939 23421 36973
rect 23457 36939 23491 36973
rect 23527 36939 23561 36973
rect 23597 36939 23631 36973
rect 22827 36871 22861 36905
rect 22897 36871 22931 36905
rect 22967 36871 23001 36905
rect 23037 36871 23071 36905
rect 23107 36871 23141 36905
rect 23177 36871 23211 36905
rect 23247 36871 23281 36905
rect 23317 36871 23351 36905
rect 23387 36871 23421 36905
rect 23457 36871 23491 36905
rect 23527 36871 23561 36905
rect 23597 36871 23631 36905
rect 22827 36803 22861 36837
rect 22897 36803 22931 36837
rect 22967 36803 23001 36837
rect 23037 36803 23071 36837
rect 23107 36803 23141 36837
rect 23177 36803 23211 36837
rect 23247 36803 23281 36837
rect 23317 36803 23351 36837
rect 23387 36803 23421 36837
rect 23457 36803 23491 36837
rect 23527 36803 23561 36837
rect 23597 36803 23631 36837
rect 22827 36735 22861 36769
rect 22897 36735 22931 36769
rect 22967 36735 23001 36769
rect 23037 36735 23071 36769
rect 23107 36735 23141 36769
rect 23177 36735 23211 36769
rect 23247 36735 23281 36769
rect 23317 36735 23351 36769
rect 23387 36735 23421 36769
rect 23457 36735 23491 36769
rect 23527 36735 23561 36769
rect 23597 36735 23631 36769
rect 22827 36667 22861 36701
rect 22897 36667 22931 36701
rect 22967 36667 23001 36701
rect 23037 36667 23071 36701
rect 23107 36667 23141 36701
rect 23177 36667 23211 36701
rect 23247 36667 23281 36701
rect 23317 36667 23351 36701
rect 23387 36667 23421 36701
rect 23457 36667 23491 36701
rect 23527 36667 23561 36701
rect 23597 36667 23631 36701
rect 22827 36599 22861 36633
rect 22897 36599 22931 36633
rect 22967 36599 23001 36633
rect 23037 36599 23071 36633
rect 23107 36599 23141 36633
rect 23177 36599 23211 36633
rect 23247 36599 23281 36633
rect 23317 36599 23351 36633
rect 23387 36599 23421 36633
rect 23457 36599 23491 36633
rect 23527 36599 23561 36633
rect 23597 36599 23631 36633
rect 22827 36531 22861 36565
rect 22897 36531 22931 36565
rect 22967 36531 23001 36565
rect 23037 36531 23071 36565
rect 23107 36531 23141 36565
rect 23177 36531 23211 36565
rect 23247 36531 23281 36565
rect 23317 36531 23351 36565
rect 23387 36531 23421 36565
rect 23457 36531 23491 36565
rect 23527 36531 23561 36565
rect 23597 36531 23631 36565
rect 22827 36463 22861 36497
rect 22897 36463 22931 36497
rect 22967 36463 23001 36497
rect 23037 36463 23071 36497
rect 23107 36463 23141 36497
rect 23177 36463 23211 36497
rect 23247 36463 23281 36497
rect 23317 36463 23351 36497
rect 23387 36463 23421 36497
rect 23457 36463 23491 36497
rect 23527 36463 23561 36497
rect 23597 36463 23631 36497
rect 22827 36395 22861 36429
rect 22897 36395 22931 36429
rect 22967 36395 23001 36429
rect 23037 36395 23071 36429
rect 23107 36395 23141 36429
rect 23177 36395 23211 36429
rect 23247 36395 23281 36429
rect 23317 36395 23351 36429
rect 23387 36395 23421 36429
rect 23457 36395 23491 36429
rect 23527 36395 23561 36429
rect 23597 36395 23631 36429
rect 22827 36327 22861 36361
rect 22897 36327 22931 36361
rect 22967 36327 23001 36361
rect 23037 36327 23071 36361
rect 23107 36327 23141 36361
rect 23177 36327 23211 36361
rect 23247 36327 23281 36361
rect 23317 36327 23351 36361
rect 23387 36327 23421 36361
rect 23457 36327 23491 36361
rect 23527 36327 23561 36361
rect 23597 36327 23631 36361
rect 22827 36259 22861 36293
rect 22897 36259 22931 36293
rect 22967 36259 23001 36293
rect 23037 36259 23071 36293
rect 23107 36259 23141 36293
rect 23177 36259 23211 36293
rect 23247 36259 23281 36293
rect 23317 36259 23351 36293
rect 23387 36259 23421 36293
rect 23457 36259 23491 36293
rect 23527 36259 23561 36293
rect 23597 36259 23631 36293
rect 22827 36191 22861 36225
rect 22897 36191 22931 36225
rect 22967 36191 23001 36225
rect 23037 36191 23071 36225
rect 23107 36191 23141 36225
rect 23177 36191 23211 36225
rect 23247 36191 23281 36225
rect 23317 36191 23351 36225
rect 23387 36191 23421 36225
rect 23457 36191 23491 36225
rect 23527 36191 23561 36225
rect 23597 36191 23631 36225
rect 22827 36123 22861 36157
rect 22897 36123 22931 36157
rect 22967 36123 23001 36157
rect 23037 36123 23071 36157
rect 23107 36123 23141 36157
rect 23177 36123 23211 36157
rect 23247 36123 23281 36157
rect 23317 36123 23351 36157
rect 23387 36123 23421 36157
rect 23457 36123 23491 36157
rect 23527 36123 23561 36157
rect 23597 36123 23631 36157
rect 22827 36055 22861 36089
rect 22897 36055 22931 36089
rect 22967 36055 23001 36089
rect 23037 36055 23071 36089
rect 23107 36055 23141 36089
rect 23177 36055 23211 36089
rect 23247 36055 23281 36089
rect 23317 36055 23351 36089
rect 23387 36055 23421 36089
rect 23457 36055 23491 36089
rect 23527 36055 23561 36089
rect 23597 36055 23631 36089
rect 22827 35987 22861 36021
rect 22897 35987 22931 36021
rect 22967 35987 23001 36021
rect 23037 35987 23071 36021
rect 23107 35987 23141 36021
rect 23177 35987 23211 36021
rect 23247 35987 23281 36021
rect 23317 35987 23351 36021
rect 23387 35987 23421 36021
rect 23457 35987 23491 36021
rect 23527 35987 23561 36021
rect 23597 35987 23631 36021
rect 22827 35919 22861 35953
rect 22897 35919 22931 35953
rect 22967 35919 23001 35953
rect 23037 35919 23071 35953
rect 23107 35919 23141 35953
rect 23177 35919 23211 35953
rect 23247 35919 23281 35953
rect 23317 35919 23351 35953
rect 23387 35919 23421 35953
rect 23457 35919 23491 35953
rect 23527 35919 23561 35953
rect 23597 35919 23631 35953
rect 22827 35851 22861 35885
rect 22897 35851 22931 35885
rect 22967 35851 23001 35885
rect 23037 35851 23071 35885
rect 23107 35851 23141 35885
rect 23177 35851 23211 35885
rect 23247 35851 23281 35885
rect 23317 35851 23351 35885
rect 23387 35851 23421 35885
rect 23457 35851 23491 35885
rect 23527 35851 23561 35885
rect 23597 35851 23631 35885
rect 22827 35783 22861 35817
rect 22897 35783 22931 35817
rect 22967 35783 23001 35817
rect 23037 35783 23071 35817
rect 23107 35783 23141 35817
rect 23177 35783 23211 35817
rect 23247 35783 23281 35817
rect 23317 35783 23351 35817
rect 23387 35783 23421 35817
rect 23457 35783 23491 35817
rect 23527 35783 23561 35817
rect 23597 35783 23631 35817
rect 22827 35715 22861 35749
rect 22897 35715 22931 35749
rect 22967 35715 23001 35749
rect 23037 35715 23071 35749
rect 23107 35715 23141 35749
rect 23177 35715 23211 35749
rect 23247 35715 23281 35749
rect 23317 35715 23351 35749
rect 23387 35715 23421 35749
rect 23457 35715 23491 35749
rect 23527 35715 23561 35749
rect 23597 35715 23631 35749
rect 22827 35647 22861 35681
rect 22897 35647 22931 35681
rect 22967 35647 23001 35681
rect 23037 35647 23071 35681
rect 23107 35647 23141 35681
rect 23177 35647 23211 35681
rect 23247 35647 23281 35681
rect 23317 35647 23351 35681
rect 23387 35647 23421 35681
rect 23457 35647 23491 35681
rect 23527 35647 23561 35681
rect 23597 35647 23631 35681
rect 22827 35579 22861 35613
rect 22897 35579 22931 35613
rect 22967 35579 23001 35613
rect 23037 35579 23071 35613
rect 23107 35579 23141 35613
rect 23177 35579 23211 35613
rect 23247 35579 23281 35613
rect 23317 35579 23351 35613
rect 23387 35579 23421 35613
rect 23457 35579 23491 35613
rect 23527 35579 23561 35613
rect 23597 35579 23631 35613
rect 22827 35511 22861 35545
rect 22897 35511 22931 35545
rect 22967 35511 23001 35545
rect 23037 35511 23071 35545
rect 23107 35511 23141 35545
rect 23177 35511 23211 35545
rect 23247 35511 23281 35545
rect 23317 35511 23351 35545
rect 23387 35511 23421 35545
rect 23457 35511 23491 35545
rect 23527 35511 23561 35545
rect 23597 35511 23631 35545
rect 22827 35443 22861 35477
rect 22897 35443 22931 35477
rect 22967 35443 23001 35477
rect 23037 35443 23071 35477
rect 23107 35443 23141 35477
rect 23177 35443 23211 35477
rect 23247 35443 23281 35477
rect 23317 35443 23351 35477
rect 23387 35443 23421 35477
rect 23457 35443 23491 35477
rect 23527 35443 23561 35477
rect 23597 35443 23631 35477
rect 22827 35375 22861 35409
rect 22897 35375 22931 35409
rect 22967 35375 23001 35409
rect 23037 35375 23071 35409
rect 23107 35375 23141 35409
rect 23177 35375 23211 35409
rect 23247 35375 23281 35409
rect 23317 35375 23351 35409
rect 23387 35375 23421 35409
rect 23457 35375 23491 35409
rect 23527 35375 23561 35409
rect 23597 35375 23631 35409
rect 22827 35307 22861 35341
rect 22897 35307 22931 35341
rect 22967 35307 23001 35341
rect 23037 35307 23071 35341
rect 23107 35307 23141 35341
rect 23177 35307 23211 35341
rect 23247 35307 23281 35341
rect 23317 35307 23351 35341
rect 23387 35307 23421 35341
rect 23457 35307 23491 35341
rect 23527 35307 23561 35341
rect 23597 35307 23631 35341
rect 22827 35239 22861 35273
rect 22897 35239 22931 35273
rect 22967 35239 23001 35273
rect 23037 35239 23071 35273
rect 23107 35239 23141 35273
rect 23177 35239 23211 35273
rect 23247 35239 23281 35273
rect 23317 35239 23351 35273
rect 23387 35239 23421 35273
rect 23457 35239 23491 35273
rect 23527 35239 23561 35273
rect 23597 35239 23631 35273
rect 22827 35171 22861 35205
rect 22897 35171 22931 35205
rect 22967 35171 23001 35205
rect 23037 35171 23071 35205
rect 23107 35171 23141 35205
rect 23177 35171 23211 35205
rect 23247 35171 23281 35205
rect 23317 35171 23351 35205
rect 23387 35171 23421 35205
rect 23457 35171 23491 35205
rect 23527 35171 23561 35205
rect 23597 35171 23631 35205
rect 22827 35103 22861 35137
rect 22897 35103 22931 35137
rect 22967 35103 23001 35137
rect 23037 35103 23071 35137
rect 23107 35103 23141 35137
rect 23177 35103 23211 35137
rect 23247 35103 23281 35137
rect 23317 35103 23351 35137
rect 23387 35103 23421 35137
rect 23457 35103 23491 35137
rect 23527 35103 23561 35137
rect 23597 35103 23631 35137
rect 22827 35035 22861 35069
rect 22897 35035 22931 35069
rect 22967 35035 23001 35069
rect 23037 35035 23071 35069
rect 23107 35035 23141 35069
rect 23177 35035 23211 35069
rect 23247 35035 23281 35069
rect 23317 35035 23351 35069
rect 23387 35035 23421 35069
rect 23457 35035 23491 35069
rect 23527 35035 23561 35069
rect 23597 35035 23631 35069
rect 22827 34967 22861 35001
rect 22897 34967 22931 35001
rect 22967 34967 23001 35001
rect 23037 34967 23071 35001
rect 23107 34967 23141 35001
rect 23177 34967 23211 35001
rect 23247 34967 23281 35001
rect 23317 34967 23351 35001
rect 23387 34967 23421 35001
rect 23457 34967 23491 35001
rect 23527 34967 23561 35001
rect 23597 34967 23631 35001
rect 22827 34899 22861 34933
rect 22897 34899 22931 34933
rect 22967 34899 23001 34933
rect 23037 34899 23071 34933
rect 23107 34899 23141 34933
rect 23177 34899 23211 34933
rect 23247 34899 23281 34933
rect 23317 34899 23351 34933
rect 23387 34899 23421 34933
rect 23457 34899 23491 34933
rect 23527 34899 23561 34933
rect 23597 34899 23631 34933
rect 22827 34831 22861 34865
rect 22897 34831 22931 34865
rect 22967 34831 23001 34865
rect 23037 34831 23071 34865
rect 23107 34831 23141 34865
rect 23177 34831 23211 34865
rect 23247 34831 23281 34865
rect 23317 34831 23351 34865
rect 23387 34831 23421 34865
rect 23457 34831 23491 34865
rect 23527 34831 23561 34865
rect 23597 34831 23631 34865
rect 22827 34763 22861 34797
rect 22897 34763 22931 34797
rect 22967 34763 23001 34797
rect 23037 34763 23071 34797
rect 23107 34763 23141 34797
rect 23177 34763 23211 34797
rect 23247 34763 23281 34797
rect 23317 34763 23351 34797
rect 23387 34763 23421 34797
rect 23457 34763 23491 34797
rect 23527 34763 23561 34797
rect 23597 34763 23631 34797
rect 22827 34695 22861 34729
rect 22897 34695 22931 34729
rect 22967 34695 23001 34729
rect 23037 34695 23071 34729
rect 23107 34695 23141 34729
rect 23177 34695 23211 34729
rect 23247 34695 23281 34729
rect 23317 34695 23351 34729
rect 23387 34695 23421 34729
rect 23457 34695 23491 34729
rect 23527 34695 23561 34729
rect 23597 34695 23631 34729
rect 22827 34627 22861 34661
rect 22897 34627 22931 34661
rect 22967 34627 23001 34661
rect 23037 34627 23071 34661
rect 23107 34627 23141 34661
rect 23177 34627 23211 34661
rect 23247 34627 23281 34661
rect 23317 34627 23351 34661
rect 23387 34627 23421 34661
rect 23457 34627 23491 34661
rect 23527 34627 23561 34661
rect 23597 34627 23631 34661
rect 22827 34559 22861 34593
rect 22897 34559 22931 34593
rect 22967 34559 23001 34593
rect 23037 34559 23071 34593
rect 23107 34559 23141 34593
rect 23177 34559 23211 34593
rect 23247 34559 23281 34593
rect 23317 34559 23351 34593
rect 23387 34559 23421 34593
rect 23457 34559 23491 34593
rect 23527 34559 23561 34593
rect 23597 34559 23631 34593
rect 22827 34491 22861 34525
rect 22897 34491 22931 34525
rect 22967 34491 23001 34525
rect 23037 34491 23071 34525
rect 23107 34491 23141 34525
rect 23177 34491 23211 34525
rect 23247 34491 23281 34525
rect 23317 34491 23351 34525
rect 23387 34491 23421 34525
rect 23457 34491 23491 34525
rect 23527 34491 23561 34525
rect 23597 34491 23631 34525
rect 22827 34423 22861 34457
rect 22897 34423 22931 34457
rect 22967 34423 23001 34457
rect 23037 34423 23071 34457
rect 23107 34423 23141 34457
rect 23177 34423 23211 34457
rect 23247 34423 23281 34457
rect 23317 34423 23351 34457
rect 23387 34423 23421 34457
rect 23457 34423 23491 34457
rect 23527 34423 23561 34457
rect 23597 34423 23631 34457
rect 22827 34355 22861 34389
rect 22897 34355 22931 34389
rect 22967 34355 23001 34389
rect 23037 34355 23071 34389
rect 23107 34355 23141 34389
rect 23177 34355 23211 34389
rect 23247 34355 23281 34389
rect 23317 34355 23351 34389
rect 23387 34355 23421 34389
rect 23457 34355 23491 34389
rect 23527 34355 23561 34389
rect 23597 34355 23631 34389
rect 22827 34287 22861 34321
rect 22897 34287 22931 34321
rect 22967 34287 23001 34321
rect 23037 34287 23071 34321
rect 23107 34287 23141 34321
rect 23177 34287 23211 34321
rect 23247 34287 23281 34321
rect 23317 34287 23351 34321
rect 23387 34287 23421 34321
rect 23457 34287 23491 34321
rect 23527 34287 23561 34321
rect 23597 34287 23631 34321
rect 22827 34219 22861 34253
rect 22897 34219 22931 34253
rect 22967 34219 23001 34253
rect 23037 34219 23071 34253
rect 23107 34219 23141 34253
rect 23177 34219 23211 34253
rect 23247 34219 23281 34253
rect 23317 34219 23351 34253
rect 23387 34219 23421 34253
rect 23457 34219 23491 34253
rect 23527 34219 23561 34253
rect 23597 34219 23631 34253
rect 22827 34151 22861 34185
rect 22897 34151 22931 34185
rect 22967 34151 23001 34185
rect 23037 34151 23071 34185
rect 23107 34151 23141 34185
rect 23177 34151 23211 34185
rect 23247 34151 23281 34185
rect 23317 34151 23351 34185
rect 23387 34151 23421 34185
rect 23457 34151 23491 34185
rect 23527 34151 23561 34185
rect 23597 34151 23631 34185
rect 22827 34083 22861 34117
rect 22897 34083 22931 34117
rect 22967 34083 23001 34117
rect 23037 34083 23071 34117
rect 23107 34083 23141 34117
rect 23177 34083 23211 34117
rect 23247 34083 23281 34117
rect 23317 34083 23351 34117
rect 23387 34083 23421 34117
rect 23457 34083 23491 34117
rect 23527 34083 23561 34117
rect 23597 34083 23631 34117
rect 22827 34015 22861 34049
rect 22897 34015 22931 34049
rect 22967 34015 23001 34049
rect 23037 34015 23071 34049
rect 23107 34015 23141 34049
rect 23177 34015 23211 34049
rect 23247 34015 23281 34049
rect 23317 34015 23351 34049
rect 23387 34015 23421 34049
rect 23457 34015 23491 34049
rect 23527 34015 23561 34049
rect 23597 34015 23631 34049
rect 22827 33947 22861 33981
rect 22897 33947 22931 33981
rect 22967 33947 23001 33981
rect 23037 33947 23071 33981
rect 23107 33947 23141 33981
rect 23177 33947 23211 33981
rect 23247 33947 23281 33981
rect 23317 33947 23351 33981
rect 23387 33947 23421 33981
rect 23457 33947 23491 33981
rect 23527 33947 23561 33981
rect 23597 33947 23631 33981
rect 22827 33879 22861 33913
rect 22897 33879 22931 33913
rect 22967 33879 23001 33913
rect 23037 33879 23071 33913
rect 23107 33879 23141 33913
rect 23177 33879 23211 33913
rect 23247 33879 23281 33913
rect 23317 33879 23351 33913
rect 23387 33879 23421 33913
rect 23457 33879 23491 33913
rect 23527 33879 23561 33913
rect 23597 33879 23631 33913
rect 22827 33811 22861 33845
rect 22897 33811 22931 33845
rect 22967 33811 23001 33845
rect 23037 33811 23071 33845
rect 23107 33811 23141 33845
rect 23177 33811 23211 33845
rect 23247 33811 23281 33845
rect 23317 33811 23351 33845
rect 23387 33811 23421 33845
rect 23457 33811 23491 33845
rect 23527 33811 23561 33845
rect 23597 33811 23631 33845
rect 22827 33743 22861 33777
rect 22897 33743 22931 33777
rect 22967 33743 23001 33777
rect 23037 33743 23071 33777
rect 23107 33743 23141 33777
rect 23177 33743 23211 33777
rect 23247 33743 23281 33777
rect 23317 33743 23351 33777
rect 23387 33743 23421 33777
rect 23457 33743 23491 33777
rect 23527 33743 23561 33777
rect 23597 33743 23631 33777
rect 22827 33675 22861 33709
rect 22897 33675 22931 33709
rect 22967 33675 23001 33709
rect 23037 33675 23071 33709
rect 23107 33675 23141 33709
rect 23177 33675 23211 33709
rect 23247 33675 23281 33709
rect 23317 33675 23351 33709
rect 23387 33675 23421 33709
rect 23457 33675 23491 33709
rect 23527 33675 23561 33709
rect 23597 33675 23631 33709
rect 22827 33607 22861 33641
rect 22897 33607 22931 33641
rect 22967 33607 23001 33641
rect 23037 33607 23071 33641
rect 23107 33607 23141 33641
rect 23177 33607 23211 33641
rect 23247 33607 23281 33641
rect 23317 33607 23351 33641
rect 23387 33607 23421 33641
rect 23457 33607 23491 33641
rect 23527 33607 23561 33641
rect 23597 33607 23631 33641
rect 22827 33539 22861 33573
rect 22897 33539 22931 33573
rect 22967 33539 23001 33573
rect 23037 33539 23071 33573
rect 23107 33539 23141 33573
rect 23177 33539 23211 33573
rect 23247 33539 23281 33573
rect 23317 33539 23351 33573
rect 23387 33539 23421 33573
rect 23457 33539 23491 33573
rect 23527 33539 23561 33573
rect 23597 33539 23631 33573
rect 22827 33471 22861 33505
rect 22897 33471 22931 33505
rect 22967 33471 23001 33505
rect 23037 33471 23071 33505
rect 23107 33471 23141 33505
rect 23177 33471 23211 33505
rect 23247 33471 23281 33505
rect 23317 33471 23351 33505
rect 23387 33471 23421 33505
rect 23457 33471 23491 33505
rect 23527 33471 23561 33505
rect 23597 33471 23631 33505
rect 22827 33403 22861 33437
rect 22897 33403 22931 33437
rect 22967 33403 23001 33437
rect 23037 33403 23071 33437
rect 23107 33403 23141 33437
rect 23177 33403 23211 33437
rect 23247 33403 23281 33437
rect 23317 33403 23351 33437
rect 23387 33403 23421 33437
rect 23457 33403 23491 33437
rect 23527 33403 23561 33437
rect 23597 33403 23631 33437
rect 22827 33335 22861 33369
rect 22897 33335 22931 33369
rect 22967 33335 23001 33369
rect 23037 33335 23071 33369
rect 23107 33335 23141 33369
rect 23177 33335 23211 33369
rect 23247 33335 23281 33369
rect 23317 33335 23351 33369
rect 23387 33335 23421 33369
rect 23457 33335 23491 33369
rect 23527 33335 23561 33369
rect 23597 33335 23631 33369
rect 278 33247 312 33281
rect 278 33178 312 33212
rect 278 33109 312 33143
rect 278 33040 312 33074
rect 278 32971 312 33005
rect 278 32902 312 32936
rect 278 32833 312 32867
rect 278 32764 312 32798
rect 278 32695 312 32729
rect 278 32626 312 32660
rect 278 32557 312 32591
rect 278 32488 312 32522
rect 278 32419 312 32453
rect 278 32350 312 32384
rect 18025 33273 18059 33307
rect 18101 33273 18135 33307
rect 18177 33273 18211 33307
rect 18253 33273 18287 33307
rect 18329 33273 18363 33307
rect 18405 33273 18439 33307
rect 18025 33205 18059 33239
rect 18101 33205 18135 33239
rect 18177 33205 18211 33239
rect 18253 33205 18287 33239
rect 18329 33205 18363 33239
rect 18405 33205 18439 33239
rect 18025 33137 18059 33171
rect 18101 33137 18135 33171
rect 18177 33137 18211 33171
rect 18253 33137 18287 33171
rect 18329 33137 18363 33171
rect 18405 33137 18439 33171
rect 18025 33069 18059 33103
rect 18101 33069 18135 33103
rect 18177 33069 18211 33103
rect 18253 33069 18287 33103
rect 18329 33069 18363 33103
rect 18405 33069 18439 33103
rect 18025 33001 18059 33035
rect 18101 33001 18135 33035
rect 18177 33001 18211 33035
rect 18253 33001 18287 33035
rect 18329 33001 18363 33035
rect 18405 33001 18439 33035
rect 18025 32933 18059 32967
rect 18101 32933 18135 32967
rect 18177 32933 18211 32967
rect 18253 32933 18287 32967
rect 18329 32933 18363 32967
rect 18405 32933 18439 32967
rect 18025 32865 18059 32899
rect 18101 32865 18135 32899
rect 18177 32865 18211 32899
rect 18253 32865 18287 32899
rect 18329 32865 18363 32899
rect 18405 32865 18439 32899
rect 18025 32797 18059 32831
rect 18101 32797 18135 32831
rect 18177 32797 18211 32831
rect 18253 32797 18287 32831
rect 18329 32797 18363 32831
rect 18405 32797 18439 32831
rect 18025 32729 18059 32763
rect 18101 32729 18135 32763
rect 18177 32729 18211 32763
rect 18253 32729 18287 32763
rect 18329 32729 18363 32763
rect 18405 32729 18439 32763
rect 18025 32661 18059 32695
rect 18101 32661 18135 32695
rect 18177 32661 18211 32695
rect 18253 32661 18287 32695
rect 18329 32661 18363 32695
rect 18405 32661 18439 32695
rect 18025 32593 18059 32627
rect 18101 32593 18135 32627
rect 18177 32593 18211 32627
rect 18253 32593 18287 32627
rect 18329 32593 18363 32627
rect 18405 32593 18439 32627
rect 18025 32525 18059 32559
rect 18101 32525 18135 32559
rect 18177 32525 18211 32559
rect 18253 32525 18287 32559
rect 18329 32525 18363 32559
rect 18405 32525 18439 32559
rect 18025 32457 18059 32491
rect 18101 32457 18135 32491
rect 18177 32457 18211 32491
rect 18253 32457 18287 32491
rect 18329 32457 18363 32491
rect 18405 32457 18439 32491
rect 18025 32389 18059 32423
rect 18101 32389 18135 32423
rect 18177 32389 18211 32423
rect 18253 32389 18287 32423
rect 18329 32389 18363 32423
rect 18405 32389 18439 32423
rect 18025 32321 18059 32355
rect 18101 32321 18135 32355
rect 18177 32321 18211 32355
rect 18253 32321 18287 32355
rect 18329 32321 18363 32355
rect 18405 32321 18439 32355
rect 278 32281 312 32315
rect 368 32248 402 32282
rect 440 32248 474 32282
rect 512 32248 546 32282
rect 584 32248 618 32282
rect 656 32248 690 32282
rect 728 32248 762 32282
rect 800 32248 834 32282
rect 872 32248 906 32282
rect 278 32212 312 32246
rect 278 32143 312 32177
rect 368 32172 402 32206
rect 440 32172 474 32206
rect 512 32172 546 32206
rect 584 32172 618 32206
rect 656 32172 690 32206
rect 728 32172 762 32206
rect 800 32172 834 32206
rect 872 32172 906 32206
rect 278 32074 312 32108
rect 368 32096 402 32130
rect 440 32096 474 32130
rect 512 32096 546 32130
rect 584 32096 618 32130
rect 656 32096 690 32130
rect 728 32096 762 32130
rect 800 32096 834 32130
rect 872 32096 906 32130
rect 278 32005 312 32039
rect 368 32020 402 32054
rect 440 32020 474 32054
rect 512 32020 546 32054
rect 584 32020 618 32054
rect 656 32020 690 32054
rect 728 32020 762 32054
rect 800 32020 834 32054
rect 872 32020 906 32054
rect 278 31936 312 31970
rect 368 31944 402 31978
rect 440 31944 474 31978
rect 512 31944 546 31978
rect 584 31944 618 31978
rect 656 31944 690 31978
rect 728 31944 762 31978
rect 800 31944 834 31978
rect 872 31944 906 31978
rect 278 31867 312 31901
rect 368 31868 402 31902
rect 440 31868 474 31902
rect 512 31868 546 31902
rect 584 31868 618 31902
rect 656 31868 690 31902
rect 728 31868 762 31902
rect 800 31868 834 31902
rect 872 31868 906 31902
rect 278 31798 312 31832
rect 368 31791 402 31825
rect 440 31791 474 31825
rect 512 31791 546 31825
rect 584 31791 618 31825
rect 656 31791 690 31825
rect 728 31791 762 31825
rect 800 31791 834 31825
rect 872 31791 906 31825
rect 278 31729 312 31763
rect 18025 32253 18059 32287
rect 18101 32253 18135 32287
rect 18177 32253 18211 32287
rect 18253 32253 18287 32287
rect 18329 32253 18363 32287
rect 18405 32253 18439 32287
rect 18025 32185 18059 32219
rect 18101 32185 18135 32219
rect 18177 32185 18211 32219
rect 18253 32185 18287 32219
rect 18329 32185 18363 32219
rect 18405 32185 18439 32219
rect 18025 32117 18059 32151
rect 18101 32117 18135 32151
rect 18177 32117 18211 32151
rect 18253 32117 18287 32151
rect 18329 32117 18363 32151
rect 18405 32117 18439 32151
rect 18025 32049 18059 32083
rect 18101 32049 18135 32083
rect 18177 32049 18211 32083
rect 18253 32049 18287 32083
rect 18329 32049 18363 32083
rect 18405 32049 18439 32083
rect 18025 31981 18059 32015
rect 18101 31981 18135 32015
rect 18177 31981 18211 32015
rect 18253 31981 18287 32015
rect 18329 31981 18363 32015
rect 18405 31981 18439 32015
rect 18025 31913 18059 31947
rect 18101 31913 18135 31947
rect 18177 31913 18211 31947
rect 18253 31913 18287 31947
rect 18329 31913 18363 31947
rect 18405 31913 18439 31947
rect 18025 31845 18059 31879
rect 18101 31845 18135 31879
rect 18177 31845 18211 31879
rect 18253 31845 18287 31879
rect 18329 31845 18363 31879
rect 18405 31845 18439 31879
rect 18025 31777 18059 31811
rect 18101 31777 18135 31811
rect 18177 31777 18211 31811
rect 18253 31777 18287 31811
rect 18329 31777 18363 31811
rect 18405 31777 18439 31811
rect 18025 31709 18059 31743
rect 18101 31709 18135 31743
rect 18177 31709 18211 31743
rect 18253 31709 18287 31743
rect 18329 31709 18363 31743
rect 18405 31709 18439 31743
rect 1051 31637 1085 31671
rect 1127 31637 1161 31671
rect 1203 31637 1237 31671
rect 1279 31637 1313 31671
rect 1051 31569 1085 31603
rect 1127 31569 1161 31603
rect 1203 31569 1237 31603
rect 1279 31569 1313 31603
rect 1051 31501 1085 31535
rect 1127 31501 1161 31535
rect 1203 31501 1237 31535
rect 1279 31501 1313 31535
rect 1051 31433 1085 31467
rect 1127 31433 1161 31467
rect 1203 31433 1237 31467
rect 1279 31433 1313 31467
rect 1051 31365 1085 31399
rect 1127 31365 1161 31399
rect 1203 31365 1237 31399
rect 1279 31365 1313 31399
rect 1051 31297 1085 31331
rect 1127 31297 1161 31331
rect 1203 31297 1237 31331
rect 1279 31297 1313 31331
rect 1051 31229 1085 31263
rect 1127 31229 1161 31263
rect 1203 31229 1237 31263
rect 1279 31229 1313 31263
rect 1051 31161 1085 31195
rect 1127 31161 1161 31195
rect 1203 31161 1237 31195
rect 1279 31161 1313 31195
rect 1051 31093 1085 31127
rect 1127 31093 1161 31127
rect 1203 31093 1237 31127
rect 1279 31093 1313 31127
rect 1051 31025 1085 31059
rect 1127 31025 1161 31059
rect 1203 31025 1237 31059
rect 1279 31025 1313 31059
rect 1051 30957 1085 30991
rect 1127 30957 1161 30991
rect 1203 30957 1237 30991
rect 1279 30957 1313 30991
rect 1051 30889 1085 30923
rect 1127 30889 1161 30923
rect 1203 30889 1237 30923
rect 1279 30889 1313 30923
rect 1051 30821 1085 30855
rect 1127 30821 1161 30855
rect 1203 30821 1237 30855
rect 1279 30821 1313 30855
rect 1051 30753 1085 30787
rect 1127 30753 1161 30787
rect 1203 30753 1237 30787
rect 1279 30753 1313 30787
rect 1051 30685 1085 30719
rect 1127 30685 1161 30719
rect 1203 30685 1237 30719
rect 1279 30685 1313 30719
rect 1051 30617 1085 30651
rect 1127 30617 1161 30651
rect 1203 30617 1237 30651
rect 1279 30617 1313 30651
rect 1051 30549 1085 30583
rect 1127 30549 1161 30583
rect 1203 30549 1237 30583
rect 1279 30549 1313 30583
rect 1051 30481 1085 30515
rect 1127 30481 1161 30515
rect 1203 30481 1237 30515
rect 1279 30481 1313 30515
rect 1051 30413 1085 30447
rect 1127 30413 1161 30447
rect 1203 30413 1237 30447
rect 1279 30413 1313 30447
rect 1051 30345 1085 30379
rect 1127 30345 1161 30379
rect 1203 30345 1237 30379
rect 1279 30345 1313 30379
rect 1051 30277 1085 30311
rect 1127 30277 1161 30311
rect 1203 30277 1237 30311
rect 1279 30277 1313 30311
rect 1051 30209 1085 30243
rect 1127 30209 1161 30243
rect 1203 30209 1237 30243
rect 1279 30209 1313 30243
rect 1051 30141 1085 30175
rect 1127 30141 1161 30175
rect 1203 30141 1237 30175
rect 1279 30141 1313 30175
rect 1051 30073 1085 30107
rect 1127 30073 1161 30107
rect 1203 30073 1237 30107
rect 1279 30073 1313 30107
rect 1051 30005 1085 30039
rect 1127 30005 1161 30039
rect 1203 30005 1237 30039
rect 1279 30005 1313 30039
rect 1051 29937 1085 29971
rect 1127 29937 1161 29971
rect 1203 29937 1237 29971
rect 1279 29937 1313 29971
rect 1051 29869 1085 29903
rect 1127 29869 1161 29903
rect 1203 29869 1237 29903
rect 1279 29869 1313 29903
rect 1051 29801 1085 29835
rect 1127 29801 1161 29835
rect 1203 29801 1237 29835
rect 1279 29801 1313 29835
rect 1051 29733 1085 29767
rect 1127 29733 1161 29767
rect 1203 29733 1237 29767
rect 1279 29733 1313 29767
rect 1051 29665 1085 29699
rect 1127 29665 1161 29699
rect 1203 29665 1237 29699
rect 1279 29665 1313 29699
rect 1051 29597 1085 29631
rect 1127 29597 1161 29631
rect 1203 29597 1237 29631
rect 1279 29597 1313 29631
rect 1051 29529 1085 29563
rect 1127 29529 1161 29563
rect 1203 29529 1237 29563
rect 1279 29529 1313 29563
rect 1051 29461 1085 29495
rect 1127 29461 1161 29495
rect 1203 29461 1237 29495
rect 1279 29461 1313 29495
rect 1051 29393 1085 29427
rect 1127 29393 1161 29427
rect 1203 29393 1237 29427
rect 1279 29393 1313 29427
rect 1051 29325 1085 29359
rect 1127 29325 1161 29359
rect 1203 29325 1237 29359
rect 1279 29325 1313 29359
rect 1051 29257 1085 29291
rect 1127 29257 1161 29291
rect 1203 29257 1237 29291
rect 1279 29257 1313 29291
rect 1051 29189 1085 29223
rect 1127 29189 1161 29223
rect 1203 29189 1237 29223
rect 1279 29189 1313 29223
rect 1051 29121 1085 29155
rect 1127 29121 1161 29155
rect 1203 29121 1237 29155
rect 1279 29121 1313 29155
rect 1051 29052 1085 29086
rect 1127 29052 1161 29086
rect 1203 29052 1237 29086
rect 1279 29052 1313 29086
rect 1051 28983 1085 29017
rect 1127 28983 1161 29017
rect 1203 28983 1237 29017
rect 1279 28983 1313 29017
rect 1051 28914 1085 28948
rect 1127 28914 1161 28948
rect 1203 28914 1237 28948
rect 1279 28914 1313 28948
rect 1051 28845 1085 28879
rect 1127 28845 1161 28879
rect 1203 28845 1237 28879
rect 1279 28845 1313 28879
rect 1051 28776 1085 28810
rect 1127 28776 1161 28810
rect 1203 28776 1237 28810
rect 1279 28776 1313 28810
rect 1051 28707 1085 28741
rect 1127 28707 1161 28741
rect 1203 28707 1237 28741
rect 1279 28707 1313 28741
rect 1051 28638 1085 28672
rect 1127 28638 1161 28672
rect 1203 28638 1237 28672
rect 1279 28638 1313 28672
rect 1051 28569 1085 28603
rect 1127 28569 1161 28603
rect 1203 28569 1237 28603
rect 1279 28569 1313 28603
rect 1051 28500 1085 28534
rect 1127 28500 1161 28534
rect 1203 28500 1237 28534
rect 1279 28500 1313 28534
rect 1051 28431 1085 28465
rect 1127 28431 1161 28465
rect 1203 28431 1237 28465
rect 1279 28431 1313 28465
rect 1051 28362 1085 28396
rect 1127 28362 1161 28396
rect 1203 28362 1237 28396
rect 1279 28362 1313 28396
rect 1051 28293 1085 28327
rect 1127 28293 1161 28327
rect 1203 28293 1237 28327
rect 1279 28293 1313 28327
rect 1051 28224 1085 28258
rect 1127 28224 1161 28258
rect 1203 28224 1237 28258
rect 1279 28224 1313 28258
rect 1051 28155 1085 28189
rect 1127 28155 1161 28189
rect 1203 28155 1237 28189
rect 1279 28155 1313 28189
rect 1051 28086 1085 28120
rect 1127 28086 1161 28120
rect 1203 28086 1237 28120
rect 1279 28086 1313 28120
rect 1051 28017 1085 28051
rect 1127 28017 1161 28051
rect 1203 28017 1237 28051
rect 1279 28017 1313 28051
rect 1051 27948 1085 27982
rect 1127 27948 1161 27982
rect 1203 27948 1237 27982
rect 1279 27948 1313 27982
rect 1051 27879 1085 27913
rect 1127 27879 1161 27913
rect 1203 27879 1237 27913
rect 1279 27879 1313 27913
rect 1051 27810 1085 27844
rect 1127 27810 1161 27844
rect 1203 27810 1237 27844
rect 1279 27810 1313 27844
rect 1051 27741 1085 27775
rect 1127 27741 1161 27775
rect 1203 27741 1237 27775
rect 1279 27741 1313 27775
rect 1051 27672 1085 27706
rect 1127 27672 1161 27706
rect 1203 27672 1237 27706
rect 1279 27672 1313 27706
rect 1051 27603 1085 27637
rect 1127 27603 1161 27637
rect 1203 27603 1237 27637
rect 1279 27603 1313 27637
rect 1051 27534 1085 27568
rect 1127 27534 1161 27568
rect 1203 27534 1237 27568
rect 1279 27534 1313 27568
rect 1051 27465 1085 27499
rect 1127 27465 1161 27499
rect 1203 27465 1237 27499
rect 1279 27465 1313 27499
rect 1051 27396 1085 27430
rect 1127 27396 1161 27430
rect 1203 27396 1237 27430
rect 1279 27396 1313 27430
rect 1051 27327 1085 27361
rect 1127 27327 1161 27361
rect 1203 27327 1237 27361
rect 1279 27327 1313 27361
rect 1051 27258 1085 27292
rect 1127 27258 1161 27292
rect 1203 27258 1237 27292
rect 1279 27258 1313 27292
rect 1051 27189 1085 27223
rect 1127 27189 1161 27223
rect 1203 27189 1237 27223
rect 1279 27189 1313 27223
rect 18025 31641 18059 31675
rect 18101 31641 18135 31675
rect 18177 31641 18211 31675
rect 18253 31641 18287 31675
rect 18329 31641 18363 31675
rect 18405 31641 18439 31675
rect 18025 31573 18059 31607
rect 18101 31573 18135 31607
rect 18177 31573 18211 31607
rect 18253 31573 18287 31607
rect 18329 31573 18363 31607
rect 18405 31573 18439 31607
rect 18025 31505 18059 31539
rect 18101 31505 18135 31539
rect 18177 31505 18211 31539
rect 18253 31505 18287 31539
rect 18329 31505 18363 31539
rect 18405 31505 18439 31539
rect 18025 31437 18059 31471
rect 18101 31437 18135 31471
rect 18177 31437 18211 31471
rect 18253 31437 18287 31471
rect 18329 31437 18363 31471
rect 18405 31437 18439 31471
rect 18025 31369 18059 31403
rect 18101 31369 18135 31403
rect 18177 31369 18211 31403
rect 18253 31369 18287 31403
rect 18329 31369 18363 31403
rect 18405 31369 18439 31403
rect 18025 31301 18059 31335
rect 18101 31301 18135 31335
rect 18177 31301 18211 31335
rect 18253 31301 18287 31335
rect 18329 31301 18363 31335
rect 18405 31301 18439 31335
rect 18025 31233 18059 31267
rect 18101 31233 18135 31267
rect 18177 31233 18211 31267
rect 18253 31233 18287 31267
rect 18329 31233 18363 31267
rect 18405 31233 18439 31267
rect 18025 31165 18059 31199
rect 18101 31165 18135 31199
rect 18177 31165 18211 31199
rect 18253 31165 18287 31199
rect 18329 31165 18363 31199
rect 18405 31165 18439 31199
rect 18025 31097 18059 31131
rect 18101 31097 18135 31131
rect 18177 31097 18211 31131
rect 18253 31097 18287 31131
rect 18329 31097 18363 31131
rect 18405 31097 18439 31131
rect 18025 31029 18059 31063
rect 18101 31029 18135 31063
rect 18177 31029 18211 31063
rect 18253 31029 18287 31063
rect 18329 31029 18363 31063
rect 18405 31029 18439 31063
rect 18025 30961 18059 30995
rect 18101 30961 18135 30995
rect 18177 30961 18211 30995
rect 18253 30961 18287 30995
rect 18329 30961 18363 30995
rect 18405 30961 18439 30995
rect 18025 30893 18059 30927
rect 18101 30893 18135 30927
rect 18177 30893 18211 30927
rect 18253 30893 18287 30927
rect 18329 30893 18363 30927
rect 18405 30893 18439 30927
rect 18025 30825 18059 30859
rect 18101 30825 18135 30859
rect 18177 30825 18211 30859
rect 18253 30825 18287 30859
rect 18329 30825 18363 30859
rect 18405 30825 18439 30859
rect 18025 30757 18059 30791
rect 18101 30757 18135 30791
rect 18177 30757 18211 30791
rect 18253 30757 18287 30791
rect 18329 30757 18363 30791
rect 18405 30757 18439 30791
rect 18025 30689 18059 30723
rect 18101 30689 18135 30723
rect 18177 30689 18211 30723
rect 18253 30689 18287 30723
rect 18329 30689 18363 30723
rect 18405 30689 18439 30723
rect 22827 33267 22861 33301
rect 22897 33267 22931 33301
rect 22967 33267 23001 33301
rect 23037 33267 23071 33301
rect 23107 33267 23141 33301
rect 23177 33267 23211 33301
rect 23247 33267 23281 33301
rect 23317 33267 23351 33301
rect 23387 33267 23421 33301
rect 23457 33267 23491 33301
rect 23527 33267 23561 33301
rect 23597 33267 23631 33301
rect 22827 33199 22861 33233
rect 22897 33199 22931 33233
rect 22967 33199 23001 33233
rect 23037 33199 23071 33233
rect 23107 33199 23141 33233
rect 23177 33199 23211 33233
rect 23247 33199 23281 33233
rect 23317 33199 23351 33233
rect 23387 33199 23421 33233
rect 23457 33199 23491 33233
rect 23527 33199 23561 33233
rect 23597 33199 23631 33233
rect 22827 33131 22861 33165
rect 22897 33131 22931 33165
rect 22967 33131 23001 33165
rect 23037 33131 23071 33165
rect 23107 33131 23141 33165
rect 23177 33131 23211 33165
rect 23247 33131 23281 33165
rect 23317 33131 23351 33165
rect 23387 33131 23421 33165
rect 23457 33131 23491 33165
rect 23527 33131 23561 33165
rect 23597 33131 23631 33165
rect 22827 33063 22861 33097
rect 22897 33063 22931 33097
rect 22967 33063 23001 33097
rect 23037 33063 23071 33097
rect 23107 33063 23141 33097
rect 23177 33063 23211 33097
rect 23247 33063 23281 33097
rect 23317 33063 23351 33097
rect 23387 33063 23421 33097
rect 23457 33063 23491 33097
rect 23527 33063 23561 33097
rect 23597 33063 23631 33097
rect 22827 32995 22861 33029
rect 22897 32995 22931 33029
rect 22967 32995 23001 33029
rect 23037 32995 23071 33029
rect 23107 32995 23141 33029
rect 23177 32995 23211 33029
rect 23247 32995 23281 33029
rect 23317 32995 23351 33029
rect 23387 32995 23421 33029
rect 23457 32995 23491 33029
rect 23527 32995 23561 33029
rect 23597 32995 23631 33029
rect 22827 32927 22861 32961
rect 22897 32927 22931 32961
rect 22967 32927 23001 32961
rect 23037 32927 23071 32961
rect 23107 32927 23141 32961
rect 23177 32927 23211 32961
rect 23247 32927 23281 32961
rect 23317 32927 23351 32961
rect 23387 32927 23421 32961
rect 23457 32927 23491 32961
rect 23527 32927 23561 32961
rect 23597 32927 23631 32961
rect 22827 32859 22861 32893
rect 22897 32859 22931 32893
rect 22967 32859 23001 32893
rect 23037 32859 23071 32893
rect 23107 32859 23141 32893
rect 23177 32859 23211 32893
rect 23247 32859 23281 32893
rect 23317 32859 23351 32893
rect 23387 32859 23421 32893
rect 23457 32859 23491 32893
rect 23527 32859 23561 32893
rect 23597 32859 23631 32893
rect 22827 32791 22861 32825
rect 22897 32791 22931 32825
rect 22967 32791 23001 32825
rect 23037 32791 23071 32825
rect 23107 32791 23141 32825
rect 23177 32791 23211 32825
rect 23247 32791 23281 32825
rect 23317 32791 23351 32825
rect 23387 32791 23421 32825
rect 23457 32791 23491 32825
rect 23527 32791 23561 32825
rect 23597 32791 23631 32825
rect 22827 32723 22861 32757
rect 22897 32723 22931 32757
rect 22967 32723 23001 32757
rect 23037 32723 23071 32757
rect 23107 32723 23141 32757
rect 23177 32723 23211 32757
rect 23247 32723 23281 32757
rect 23317 32723 23351 32757
rect 23387 32723 23421 32757
rect 23457 32723 23491 32757
rect 23527 32723 23561 32757
rect 23597 32723 23631 32757
rect 22827 32655 22861 32689
rect 22897 32655 22931 32689
rect 22967 32655 23001 32689
rect 23037 32655 23071 32689
rect 23107 32655 23141 32689
rect 23177 32655 23211 32689
rect 23247 32655 23281 32689
rect 23317 32655 23351 32689
rect 23387 32655 23421 32689
rect 23457 32655 23491 32689
rect 23527 32655 23561 32689
rect 23597 32655 23631 32689
rect 22827 32587 22861 32621
rect 22897 32587 22931 32621
rect 22967 32587 23001 32621
rect 23037 32587 23071 32621
rect 23107 32587 23141 32621
rect 23177 32587 23211 32621
rect 23247 32587 23281 32621
rect 23317 32587 23351 32621
rect 23387 32587 23421 32621
rect 23457 32587 23491 32621
rect 23527 32587 23561 32621
rect 23597 32587 23631 32621
rect 22827 32519 22861 32553
rect 22897 32519 22931 32553
rect 22967 32519 23001 32553
rect 23037 32519 23071 32553
rect 23107 32519 23141 32553
rect 23177 32519 23211 32553
rect 23247 32519 23281 32553
rect 23317 32519 23351 32553
rect 23387 32519 23421 32553
rect 23457 32519 23491 32553
rect 23527 32519 23561 32553
rect 23597 32519 23631 32553
rect 22827 32451 22861 32485
rect 22897 32451 22931 32485
rect 22967 32451 23001 32485
rect 23037 32451 23071 32485
rect 23107 32451 23141 32485
rect 23177 32451 23211 32485
rect 23247 32451 23281 32485
rect 23317 32451 23351 32485
rect 23387 32451 23421 32485
rect 23457 32451 23491 32485
rect 23527 32451 23561 32485
rect 23597 32451 23631 32485
rect 22827 32383 22861 32417
rect 22897 32383 22931 32417
rect 22967 32383 23001 32417
rect 23037 32383 23071 32417
rect 23107 32383 23141 32417
rect 23177 32383 23211 32417
rect 23247 32383 23281 32417
rect 23317 32383 23351 32417
rect 23387 32383 23421 32417
rect 23457 32383 23491 32417
rect 23527 32383 23561 32417
rect 23597 32383 23631 32417
rect 22827 32315 22861 32349
rect 22897 32315 22931 32349
rect 22967 32315 23001 32349
rect 23037 32315 23071 32349
rect 23107 32315 23141 32349
rect 23177 32315 23211 32349
rect 23247 32315 23281 32349
rect 23317 32315 23351 32349
rect 23387 32315 23421 32349
rect 23457 32315 23491 32349
rect 23527 32315 23561 32349
rect 23597 32315 23631 32349
rect 22827 32247 22861 32281
rect 22897 32247 22931 32281
rect 22967 32247 23001 32281
rect 23037 32247 23071 32281
rect 23107 32247 23141 32281
rect 23177 32247 23211 32281
rect 23247 32247 23281 32281
rect 23317 32247 23351 32281
rect 23387 32247 23421 32281
rect 23457 32247 23491 32281
rect 23527 32247 23561 32281
rect 23597 32247 23631 32281
rect 22827 32179 22861 32213
rect 22897 32179 22931 32213
rect 22967 32179 23001 32213
rect 23037 32179 23071 32213
rect 23107 32179 23141 32213
rect 23177 32179 23211 32213
rect 23247 32179 23281 32213
rect 23317 32179 23351 32213
rect 23387 32179 23421 32213
rect 23457 32179 23491 32213
rect 23527 32179 23561 32213
rect 23597 32179 23631 32213
rect 22827 32111 22861 32145
rect 22897 32111 22931 32145
rect 22967 32111 23001 32145
rect 23037 32111 23071 32145
rect 23107 32111 23141 32145
rect 23177 32111 23211 32145
rect 23247 32111 23281 32145
rect 23317 32111 23351 32145
rect 23387 32111 23421 32145
rect 23457 32111 23491 32145
rect 23527 32111 23561 32145
rect 23597 32111 23631 32145
rect 22827 32043 22861 32077
rect 22897 32043 22931 32077
rect 22967 32043 23001 32077
rect 23037 32043 23071 32077
rect 23107 32043 23141 32077
rect 23177 32043 23211 32077
rect 23247 32043 23281 32077
rect 23317 32043 23351 32077
rect 23387 32043 23421 32077
rect 23457 32043 23491 32077
rect 23527 32043 23561 32077
rect 23597 32043 23631 32077
rect 22827 31975 22861 32009
rect 22897 31975 22931 32009
rect 22967 31975 23001 32009
rect 23037 31975 23071 32009
rect 23107 31975 23141 32009
rect 23177 31975 23211 32009
rect 23247 31975 23281 32009
rect 23317 31975 23351 32009
rect 23387 31975 23421 32009
rect 23457 31975 23491 32009
rect 23527 31975 23561 32009
rect 23597 31975 23631 32009
rect 22827 31907 22861 31941
rect 22897 31907 22931 31941
rect 22967 31907 23001 31941
rect 23037 31907 23071 31941
rect 23107 31907 23141 31941
rect 23177 31907 23211 31941
rect 23247 31907 23281 31941
rect 23317 31907 23351 31941
rect 23387 31907 23421 31941
rect 23457 31907 23491 31941
rect 23527 31907 23561 31941
rect 23597 31907 23631 31941
rect 22827 31839 22861 31873
rect 22897 31839 22931 31873
rect 22967 31839 23001 31873
rect 23037 31839 23071 31873
rect 23107 31839 23141 31873
rect 23177 31839 23211 31873
rect 23247 31839 23281 31873
rect 23317 31839 23351 31873
rect 23387 31839 23421 31873
rect 23457 31839 23491 31873
rect 23527 31839 23561 31873
rect 23597 31839 23631 31873
rect 22827 31771 22861 31805
rect 22897 31771 22931 31805
rect 22967 31771 23001 31805
rect 23037 31771 23071 31805
rect 23107 31771 23141 31805
rect 23177 31771 23211 31805
rect 23247 31771 23281 31805
rect 23317 31771 23351 31805
rect 23387 31771 23421 31805
rect 23457 31771 23491 31805
rect 23527 31771 23561 31805
rect 23597 31771 23631 31805
rect 22827 31703 22861 31737
rect 22897 31703 22931 31737
rect 22967 31703 23001 31737
rect 23037 31703 23071 31737
rect 23107 31703 23141 31737
rect 23177 31703 23211 31737
rect 23247 31703 23281 31737
rect 23317 31703 23351 31737
rect 23387 31703 23421 31737
rect 23457 31703 23491 31737
rect 23527 31703 23561 31737
rect 23597 31703 23631 31737
rect 22827 31635 22861 31669
rect 22897 31635 22931 31669
rect 22967 31635 23001 31669
rect 23037 31635 23071 31669
rect 23107 31635 23141 31669
rect 23177 31635 23211 31669
rect 23247 31635 23281 31669
rect 23317 31635 23351 31669
rect 23387 31635 23421 31669
rect 23457 31635 23491 31669
rect 23527 31635 23561 31669
rect 23597 31635 23631 31669
rect 22827 31567 22861 31601
rect 22897 31567 22931 31601
rect 22967 31567 23001 31601
rect 23037 31567 23071 31601
rect 23107 31567 23141 31601
rect 23177 31567 23211 31601
rect 23247 31567 23281 31601
rect 23317 31567 23351 31601
rect 23387 31567 23421 31601
rect 23457 31567 23491 31601
rect 23527 31567 23561 31601
rect 23597 31567 23631 31601
rect 22827 31499 22861 31533
rect 22897 31499 22931 31533
rect 22967 31499 23001 31533
rect 23037 31499 23071 31533
rect 23107 31499 23141 31533
rect 23177 31499 23211 31533
rect 23247 31499 23281 31533
rect 23317 31499 23351 31533
rect 23387 31499 23421 31533
rect 23457 31499 23491 31533
rect 23527 31499 23561 31533
rect 23597 31499 23631 31533
rect 22827 31431 22861 31465
rect 22897 31431 22931 31465
rect 22967 31431 23001 31465
rect 23037 31431 23071 31465
rect 23107 31431 23141 31465
rect 23177 31431 23211 31465
rect 23247 31431 23281 31465
rect 23317 31431 23351 31465
rect 23387 31431 23421 31465
rect 23457 31431 23491 31465
rect 23527 31431 23561 31465
rect 23597 31431 23631 31465
rect 22827 31363 22861 31397
rect 22897 31363 22931 31397
rect 22967 31363 23001 31397
rect 23037 31363 23071 31397
rect 23107 31363 23141 31397
rect 23177 31363 23211 31397
rect 23247 31363 23281 31397
rect 23317 31363 23351 31397
rect 23387 31363 23421 31397
rect 23457 31363 23491 31397
rect 23527 31363 23561 31397
rect 23597 31363 23631 31397
rect 22827 31295 22861 31329
rect 22897 31295 22931 31329
rect 22967 31295 23001 31329
rect 23037 31295 23071 31329
rect 23107 31295 23141 31329
rect 23177 31295 23211 31329
rect 23247 31295 23281 31329
rect 23317 31295 23351 31329
rect 23387 31295 23421 31329
rect 23457 31295 23491 31329
rect 23527 31295 23561 31329
rect 23597 31295 23631 31329
rect 22827 31227 22861 31261
rect 22897 31227 22931 31261
rect 22967 31227 23001 31261
rect 23037 31227 23071 31261
rect 23107 31227 23141 31261
rect 23177 31227 23211 31261
rect 23247 31227 23281 31261
rect 23317 31227 23351 31261
rect 23387 31227 23421 31261
rect 23457 31227 23491 31261
rect 23527 31227 23561 31261
rect 23597 31227 23631 31261
rect 22827 31159 22861 31193
rect 22897 31159 22931 31193
rect 22967 31159 23001 31193
rect 23037 31159 23071 31193
rect 23107 31159 23141 31193
rect 23177 31159 23211 31193
rect 23247 31159 23281 31193
rect 23317 31159 23351 31193
rect 23387 31159 23421 31193
rect 23457 31159 23491 31193
rect 23527 31159 23561 31193
rect 23597 31159 23631 31193
rect 22827 31091 22861 31125
rect 22897 31091 22931 31125
rect 22967 31091 23001 31125
rect 23037 31091 23071 31125
rect 23107 31091 23141 31125
rect 23177 31091 23211 31125
rect 23247 31091 23281 31125
rect 23317 31091 23351 31125
rect 23387 31091 23421 31125
rect 23457 31091 23491 31125
rect 23527 31091 23561 31125
rect 23597 31091 23631 31125
rect 22827 31023 22861 31057
rect 22897 31023 22931 31057
rect 22967 31023 23001 31057
rect 23037 31023 23071 31057
rect 23107 31023 23141 31057
rect 23177 31023 23211 31057
rect 23247 31023 23281 31057
rect 23317 31023 23351 31057
rect 23387 31023 23421 31057
rect 23457 31023 23491 31057
rect 23527 31023 23561 31057
rect 23597 31023 23631 31057
rect 22827 30955 22861 30989
rect 22897 30955 22931 30989
rect 22967 30955 23001 30989
rect 23037 30955 23071 30989
rect 23107 30955 23141 30989
rect 23177 30955 23211 30989
rect 23247 30955 23281 30989
rect 23317 30955 23351 30989
rect 23387 30955 23421 30989
rect 23457 30955 23491 30989
rect 23527 30955 23561 30989
rect 23597 30955 23631 30989
rect 22827 30887 22861 30921
rect 22897 30887 22931 30921
rect 22967 30887 23001 30921
rect 23037 30887 23071 30921
rect 23107 30887 23141 30921
rect 23177 30887 23211 30921
rect 23247 30887 23281 30921
rect 23317 30887 23351 30921
rect 23387 30887 23421 30921
rect 23457 30887 23491 30921
rect 23527 30887 23561 30921
rect 23597 30887 23631 30921
rect 22827 30819 22861 30853
rect 22897 30819 22931 30853
rect 22967 30819 23001 30853
rect 23037 30819 23071 30853
rect 23107 30819 23141 30853
rect 23177 30819 23211 30853
rect 23247 30819 23281 30853
rect 23317 30819 23351 30853
rect 23387 30819 23421 30853
rect 23457 30819 23491 30853
rect 23527 30819 23561 30853
rect 23597 30819 23631 30853
rect 22827 30751 22861 30785
rect 22897 30751 22931 30785
rect 22967 30751 23001 30785
rect 23037 30751 23071 30785
rect 23107 30751 23141 30785
rect 23177 30751 23211 30785
rect 23247 30751 23281 30785
rect 23317 30751 23351 30785
rect 23387 30751 23421 30785
rect 23457 30751 23491 30785
rect 23527 30751 23561 30785
rect 23597 30751 23631 30785
rect 18025 30621 18059 30655
rect 18101 30621 18135 30655
rect 18177 30621 18211 30655
rect 18253 30621 18287 30655
rect 18329 30621 18363 30655
rect 18405 30621 18439 30655
rect 18486 30637 18520 30671
rect 18556 30637 18590 30671
rect 18626 30637 18660 30671
rect 18696 30637 18730 30671
rect 18766 30637 18800 30671
rect 18836 30637 18870 30671
rect 18906 30637 18940 30671
rect 18976 30637 19010 30671
rect 18025 30553 18059 30587
rect 18101 30553 18135 30587
rect 18177 30553 18211 30587
rect 18253 30553 18287 30587
rect 18329 30553 18363 30587
rect 18405 30553 18439 30587
rect 18486 30569 18520 30603
rect 18556 30569 18590 30603
rect 18626 30569 18660 30603
rect 18696 30569 18730 30603
rect 18766 30569 18800 30603
rect 18836 30569 18870 30603
rect 18906 30569 18940 30603
rect 18976 30569 19010 30603
rect 18025 30485 18059 30519
rect 18101 30485 18135 30519
rect 18177 30485 18211 30519
rect 18253 30485 18287 30519
rect 18329 30485 18363 30519
rect 18405 30485 18439 30519
rect 18486 30501 18520 30535
rect 18556 30501 18590 30535
rect 18626 30501 18660 30535
rect 18696 30501 18730 30535
rect 18766 30501 18800 30535
rect 18836 30501 18870 30535
rect 18906 30501 18940 30535
rect 18976 30501 19010 30535
rect 18025 30417 18059 30451
rect 18101 30417 18135 30451
rect 18177 30417 18211 30451
rect 18253 30417 18287 30451
rect 18329 30417 18363 30451
rect 18405 30417 18439 30451
rect 18486 30433 18520 30467
rect 18556 30433 18590 30467
rect 18626 30433 18660 30467
rect 18696 30433 18730 30467
rect 18766 30433 18800 30467
rect 18836 30433 18870 30467
rect 18906 30433 18940 30467
rect 18976 30433 19010 30467
rect 18025 30349 18059 30383
rect 18101 30349 18135 30383
rect 18177 30349 18211 30383
rect 18253 30349 18287 30383
rect 18329 30349 18363 30383
rect 18405 30349 18439 30383
rect 18486 30365 18520 30399
rect 18556 30365 18590 30399
rect 18626 30365 18660 30399
rect 18696 30365 18730 30399
rect 18766 30365 18800 30399
rect 18836 30365 18870 30399
rect 18906 30365 18940 30399
rect 18976 30365 19010 30399
rect 18025 30281 18059 30315
rect 18101 30281 18135 30315
rect 18177 30281 18211 30315
rect 18253 30281 18287 30315
rect 18329 30281 18363 30315
rect 18405 30281 18439 30315
rect 18486 30297 18520 30331
rect 18556 30297 18590 30331
rect 18626 30297 18660 30331
rect 18696 30297 18730 30331
rect 18766 30297 18800 30331
rect 18836 30297 18870 30331
rect 18906 30297 18940 30331
rect 18976 30297 19010 30331
rect 18025 30213 18059 30247
rect 18101 30213 18135 30247
rect 18177 30213 18211 30247
rect 18253 30213 18287 30247
rect 18329 30213 18363 30247
rect 18405 30213 18439 30247
rect 18486 30229 18520 30263
rect 18556 30229 18590 30263
rect 18626 30229 18660 30263
rect 18696 30229 18730 30263
rect 18766 30229 18800 30263
rect 18836 30229 18870 30263
rect 18906 30229 18940 30263
rect 18976 30229 19010 30263
rect 18025 30145 18059 30179
rect 18101 30145 18135 30179
rect 18177 30145 18211 30179
rect 18253 30145 18287 30179
rect 18329 30145 18363 30179
rect 18405 30145 18439 30179
rect 18486 30161 18520 30195
rect 18556 30161 18590 30195
rect 18626 30161 18660 30195
rect 18696 30161 18730 30195
rect 18766 30161 18800 30195
rect 18836 30161 18870 30195
rect 18906 30161 18940 30195
rect 18976 30161 19010 30195
rect 18025 30077 18059 30111
rect 18101 30077 18135 30111
rect 18177 30077 18211 30111
rect 18253 30077 18287 30111
rect 18329 30077 18363 30111
rect 18405 30077 18439 30111
rect 18486 30093 18520 30127
rect 18556 30093 18590 30127
rect 18626 30093 18660 30127
rect 18696 30093 18730 30127
rect 18766 30093 18800 30127
rect 18836 30093 18870 30127
rect 18906 30093 18940 30127
rect 18976 30093 19010 30127
rect 18025 30009 18059 30043
rect 18101 30009 18135 30043
rect 18177 30009 18211 30043
rect 18253 30009 18287 30043
rect 18329 30009 18363 30043
rect 18405 30009 18439 30043
rect 18486 30025 18520 30059
rect 18556 30025 18590 30059
rect 18626 30025 18660 30059
rect 18696 30025 18730 30059
rect 18766 30025 18800 30059
rect 18836 30025 18870 30059
rect 18906 30025 18940 30059
rect 18976 30025 19010 30059
rect 18025 29941 18059 29975
rect 18101 29941 18135 29975
rect 18177 29941 18211 29975
rect 18253 29941 18287 29975
rect 18329 29941 18363 29975
rect 18405 29941 18439 29975
rect 18486 29957 18520 29991
rect 18556 29957 18590 29991
rect 18626 29957 18660 29991
rect 18696 29957 18730 29991
rect 18766 29957 18800 29991
rect 18836 29957 18870 29991
rect 18906 29957 18940 29991
rect 18976 29957 19010 29991
rect 18025 29873 18059 29907
rect 18101 29873 18135 29907
rect 18177 29873 18211 29907
rect 18253 29873 18287 29907
rect 18329 29873 18363 29907
rect 18405 29873 18439 29907
rect 18486 29889 18520 29923
rect 18556 29889 18590 29923
rect 18626 29889 18660 29923
rect 18696 29889 18730 29923
rect 18766 29889 18800 29923
rect 18836 29889 18870 29923
rect 18906 29889 18940 29923
rect 18976 29889 19010 29923
rect 18025 29805 18059 29839
rect 18101 29805 18135 29839
rect 18177 29805 18211 29839
rect 18253 29805 18287 29839
rect 18329 29805 18363 29839
rect 18405 29805 18439 29839
rect 18486 29821 18520 29855
rect 18556 29821 18590 29855
rect 18626 29821 18660 29855
rect 18696 29821 18730 29855
rect 18766 29821 18800 29855
rect 18836 29821 18870 29855
rect 18906 29821 18940 29855
rect 18976 29821 19010 29855
rect 18025 29737 18059 29771
rect 18101 29737 18135 29771
rect 18177 29737 18211 29771
rect 18253 29737 18287 29771
rect 18329 29737 18363 29771
rect 18405 29737 18439 29771
rect 18486 29753 18520 29787
rect 18556 29753 18590 29787
rect 18626 29753 18660 29787
rect 18696 29753 18730 29787
rect 18766 29753 18800 29787
rect 18836 29753 18870 29787
rect 18906 29753 18940 29787
rect 18976 29753 19010 29787
rect 18025 29669 18059 29703
rect 18101 29669 18135 29703
rect 18177 29669 18211 29703
rect 18253 29669 18287 29703
rect 18329 29669 18363 29703
rect 18405 29669 18439 29703
rect 18486 29685 18520 29719
rect 18556 29685 18590 29719
rect 18626 29685 18660 29719
rect 18696 29685 18730 29719
rect 18766 29685 18800 29719
rect 18836 29685 18870 29719
rect 18906 29685 18940 29719
rect 18976 29685 19010 29719
rect 18025 29601 18059 29635
rect 18101 29601 18135 29635
rect 18177 29601 18211 29635
rect 18253 29601 18287 29635
rect 18329 29601 18363 29635
rect 18405 29601 18439 29635
rect 18486 29617 18520 29651
rect 18556 29617 18590 29651
rect 18626 29617 18660 29651
rect 18696 29617 18730 29651
rect 18766 29617 18800 29651
rect 18836 29617 18870 29651
rect 18906 29617 18940 29651
rect 18976 29617 19010 29651
rect 18025 29533 18059 29567
rect 18101 29533 18135 29567
rect 18177 29533 18211 29567
rect 18253 29533 18287 29567
rect 18329 29533 18363 29567
rect 18405 29533 18439 29567
rect 18486 29549 18520 29583
rect 18556 29549 18590 29583
rect 18626 29549 18660 29583
rect 18696 29549 18730 29583
rect 18766 29549 18800 29583
rect 18836 29549 18870 29583
rect 18906 29549 18940 29583
rect 18976 29549 19010 29583
rect 18025 29465 18059 29499
rect 18101 29465 18135 29499
rect 18177 29465 18211 29499
rect 18253 29465 18287 29499
rect 18329 29465 18363 29499
rect 18405 29465 18439 29499
rect 18486 29481 18520 29515
rect 18556 29481 18590 29515
rect 18626 29481 18660 29515
rect 18696 29481 18730 29515
rect 18766 29481 18800 29515
rect 18836 29481 18870 29515
rect 18906 29481 18940 29515
rect 18976 29481 19010 29515
rect 18025 29397 18059 29431
rect 18101 29397 18135 29431
rect 18177 29397 18211 29431
rect 18253 29397 18287 29431
rect 18329 29397 18363 29431
rect 18405 29397 18439 29431
rect 18486 29413 18520 29447
rect 18556 29413 18590 29447
rect 18626 29413 18660 29447
rect 18696 29413 18730 29447
rect 18766 29413 18800 29447
rect 18836 29413 18870 29447
rect 18906 29413 18940 29447
rect 18976 29413 19010 29447
rect 18025 29329 18059 29363
rect 18101 29329 18135 29363
rect 18177 29329 18211 29363
rect 18253 29329 18287 29363
rect 18329 29329 18363 29363
rect 18405 29329 18439 29363
rect 18486 29345 18520 29379
rect 18556 29345 18590 29379
rect 18626 29345 18660 29379
rect 18696 29345 18730 29379
rect 18766 29345 18800 29379
rect 18836 29345 18870 29379
rect 18906 29345 18940 29379
rect 18976 29345 19010 29379
rect 18025 29261 18059 29295
rect 18101 29261 18135 29295
rect 18177 29261 18211 29295
rect 18253 29261 18287 29295
rect 18329 29261 18363 29295
rect 18405 29261 18439 29295
rect 18486 29277 18520 29311
rect 18556 29277 18590 29311
rect 18626 29277 18660 29311
rect 18696 29277 18730 29311
rect 18766 29277 18800 29311
rect 18836 29277 18870 29311
rect 18906 29277 18940 29311
rect 18976 29277 19010 29311
rect 18025 29193 18059 29227
rect 18101 29193 18135 29227
rect 18177 29193 18211 29227
rect 18253 29193 18287 29227
rect 18329 29193 18363 29227
rect 18405 29193 18439 29227
rect 18486 29209 18520 29243
rect 18556 29209 18590 29243
rect 18626 29209 18660 29243
rect 18696 29209 18730 29243
rect 18766 29209 18800 29243
rect 18836 29209 18870 29243
rect 18906 29209 18940 29243
rect 18976 29209 19010 29243
rect 18025 29125 18059 29159
rect 18101 29125 18135 29159
rect 18177 29125 18211 29159
rect 18253 29125 18287 29159
rect 18329 29125 18363 29159
rect 18405 29125 18439 29159
rect 18486 29141 18520 29175
rect 18556 29141 18590 29175
rect 18626 29141 18660 29175
rect 18696 29141 18730 29175
rect 18766 29141 18800 29175
rect 18836 29141 18870 29175
rect 18906 29141 18940 29175
rect 18976 29141 19010 29175
rect 18025 29057 18059 29091
rect 18101 29057 18135 29091
rect 18177 29057 18211 29091
rect 18253 29057 18287 29091
rect 18329 29057 18363 29091
rect 18405 29057 18439 29091
rect 18486 29073 18520 29107
rect 18556 29073 18590 29107
rect 18626 29073 18660 29107
rect 18696 29073 18730 29107
rect 18766 29073 18800 29107
rect 18836 29073 18870 29107
rect 18906 29073 18940 29107
rect 18976 29073 19010 29107
rect 18025 28989 18059 29023
rect 18101 28989 18135 29023
rect 18177 28989 18211 29023
rect 18253 28989 18287 29023
rect 18329 28989 18363 29023
rect 18405 28989 18439 29023
rect 18486 29005 18520 29039
rect 18556 29005 18590 29039
rect 18626 29005 18660 29039
rect 18696 29005 18730 29039
rect 18766 29005 18800 29039
rect 18836 29005 18870 29039
rect 18906 29005 18940 29039
rect 18976 29005 19010 29039
rect 18025 28921 18059 28955
rect 18101 28921 18135 28955
rect 18177 28921 18211 28955
rect 18253 28921 18287 28955
rect 18329 28921 18363 28955
rect 18405 28921 18439 28955
rect 18486 28937 18520 28971
rect 18556 28937 18590 28971
rect 18626 28937 18660 28971
rect 18696 28937 18730 28971
rect 18766 28937 18800 28971
rect 18836 28937 18870 28971
rect 18906 28937 18940 28971
rect 18976 28937 19010 28971
rect 18025 28853 18059 28887
rect 18101 28853 18135 28887
rect 18177 28853 18211 28887
rect 18253 28853 18287 28887
rect 18329 28853 18363 28887
rect 18405 28853 18439 28887
rect 18486 28869 18520 28903
rect 18556 28869 18590 28903
rect 18626 28869 18660 28903
rect 18696 28869 18730 28903
rect 18766 28869 18800 28903
rect 18836 28869 18870 28903
rect 18906 28869 18940 28903
rect 18976 28869 19010 28903
rect 18025 28785 18059 28819
rect 18101 28785 18135 28819
rect 18177 28785 18211 28819
rect 18253 28785 18287 28819
rect 18329 28785 18363 28819
rect 18405 28785 18439 28819
rect 18486 28801 18520 28835
rect 18556 28801 18590 28835
rect 18626 28801 18660 28835
rect 18696 28801 18730 28835
rect 18766 28801 18800 28835
rect 18836 28801 18870 28835
rect 18906 28801 18940 28835
rect 18976 28801 19010 28835
rect 18025 28717 18059 28751
rect 18101 28717 18135 28751
rect 18177 28717 18211 28751
rect 18253 28717 18287 28751
rect 18329 28717 18363 28751
rect 18405 28717 18439 28751
rect 18486 28733 18520 28767
rect 18556 28733 18590 28767
rect 18626 28733 18660 28767
rect 18696 28733 18730 28767
rect 18766 28733 18800 28767
rect 18836 28733 18870 28767
rect 18906 28733 18940 28767
rect 18976 28733 19010 28767
rect 18025 28649 18059 28683
rect 18101 28649 18135 28683
rect 18177 28649 18211 28683
rect 18253 28649 18287 28683
rect 18329 28649 18363 28683
rect 18405 28649 18439 28683
rect 18486 28665 18520 28699
rect 18556 28665 18590 28699
rect 18626 28665 18660 28699
rect 18696 28665 18730 28699
rect 18766 28665 18800 28699
rect 18836 28665 18870 28699
rect 18906 28665 18940 28699
rect 18976 28665 19010 28699
rect 18025 28581 18059 28615
rect 18101 28581 18135 28615
rect 18177 28581 18211 28615
rect 18253 28581 18287 28615
rect 18329 28581 18363 28615
rect 18405 28581 18439 28615
rect 18486 28597 18520 28631
rect 18556 28597 18590 28631
rect 18626 28597 18660 28631
rect 18696 28597 18730 28631
rect 18766 28597 18800 28631
rect 18836 28597 18870 28631
rect 18906 28597 18940 28631
rect 18976 28597 19010 28631
rect 18025 28513 18059 28547
rect 18101 28513 18135 28547
rect 18177 28513 18211 28547
rect 18253 28513 18287 28547
rect 18329 28513 18363 28547
rect 18405 28513 18439 28547
rect 18486 28529 18520 28563
rect 18556 28529 18590 28563
rect 18626 28529 18660 28563
rect 18696 28529 18730 28563
rect 18766 28529 18800 28563
rect 18836 28529 18870 28563
rect 18906 28529 18940 28563
rect 18976 28529 19010 28563
rect 18025 28445 18059 28479
rect 18101 28445 18135 28479
rect 18177 28445 18211 28479
rect 18253 28445 18287 28479
rect 18329 28445 18363 28479
rect 18405 28445 18439 28479
rect 18486 28461 18520 28495
rect 18556 28461 18590 28495
rect 18626 28461 18660 28495
rect 18696 28461 18730 28495
rect 18766 28461 18800 28495
rect 18836 28461 18870 28495
rect 18906 28461 18940 28495
rect 18976 28461 19010 28495
rect 18025 28377 18059 28411
rect 18101 28377 18135 28411
rect 18177 28377 18211 28411
rect 18253 28377 18287 28411
rect 18329 28377 18363 28411
rect 18405 28377 18439 28411
rect 18486 28393 18520 28427
rect 18556 28393 18590 28427
rect 18626 28393 18660 28427
rect 18696 28393 18730 28427
rect 18766 28393 18800 28427
rect 18836 28393 18870 28427
rect 18906 28393 18940 28427
rect 18976 28393 19010 28427
rect 18025 28309 18059 28343
rect 18101 28309 18135 28343
rect 18177 28309 18211 28343
rect 18253 28309 18287 28343
rect 18329 28309 18363 28343
rect 18405 28309 18439 28343
rect 18486 28325 18520 28359
rect 18556 28325 18590 28359
rect 18626 28325 18660 28359
rect 18696 28325 18730 28359
rect 18766 28325 18800 28359
rect 18836 28325 18870 28359
rect 18906 28325 18940 28359
rect 18976 28325 19010 28359
rect 18025 28241 18059 28275
rect 18101 28241 18135 28275
rect 18177 28241 18211 28275
rect 18253 28241 18287 28275
rect 18329 28241 18363 28275
rect 18405 28241 18439 28275
rect 18486 28257 18520 28291
rect 18556 28257 18590 28291
rect 18626 28257 18660 28291
rect 18696 28257 18730 28291
rect 18766 28257 18800 28291
rect 18836 28257 18870 28291
rect 18906 28257 18940 28291
rect 18976 28257 19010 28291
rect 18025 28173 18059 28207
rect 18101 28173 18135 28207
rect 18177 28173 18211 28207
rect 18253 28173 18287 28207
rect 18329 28173 18363 28207
rect 18405 28173 18439 28207
rect 18486 28189 18520 28223
rect 18556 28189 18590 28223
rect 18626 28189 18660 28223
rect 18696 28189 18730 28223
rect 18766 28189 18800 28223
rect 18836 28189 18870 28223
rect 18906 28189 18940 28223
rect 18976 28189 19010 28223
rect 18025 28105 18059 28139
rect 18101 28105 18135 28139
rect 18177 28105 18211 28139
rect 18253 28105 18287 28139
rect 18329 28105 18363 28139
rect 18405 28105 18439 28139
rect 18486 28121 18520 28155
rect 18556 28121 18590 28155
rect 18626 28121 18660 28155
rect 18696 28121 18730 28155
rect 18766 28121 18800 28155
rect 18836 28121 18870 28155
rect 18906 28121 18940 28155
rect 18976 28121 19010 28155
rect 18025 28037 18059 28071
rect 18101 28037 18135 28071
rect 18177 28037 18211 28071
rect 18253 28037 18287 28071
rect 18329 28037 18363 28071
rect 18405 28037 18439 28071
rect 18486 28053 18520 28087
rect 18556 28053 18590 28087
rect 18626 28053 18660 28087
rect 18696 28053 18730 28087
rect 18766 28053 18800 28087
rect 18836 28053 18870 28087
rect 18906 28053 18940 28087
rect 18976 28053 19010 28087
rect 18025 27969 18059 28003
rect 18101 27969 18135 28003
rect 18177 27969 18211 28003
rect 18253 27969 18287 28003
rect 18329 27969 18363 28003
rect 18405 27969 18439 28003
rect 18486 27985 18520 28019
rect 18556 27985 18590 28019
rect 18626 27985 18660 28019
rect 18696 27985 18730 28019
rect 18766 27985 18800 28019
rect 18836 27985 18870 28019
rect 18906 27985 18940 28019
rect 18976 27985 19010 28019
rect 18025 27901 18059 27935
rect 18101 27901 18135 27935
rect 18177 27901 18211 27935
rect 18253 27901 18287 27935
rect 18329 27901 18363 27935
rect 18405 27901 18439 27935
rect 18486 27917 18520 27951
rect 18556 27917 18590 27951
rect 18626 27917 18660 27951
rect 18696 27917 18730 27951
rect 18766 27917 18800 27951
rect 18836 27917 18870 27951
rect 18906 27917 18940 27951
rect 18976 27917 19010 27951
rect 18025 27833 18059 27867
rect 18101 27833 18135 27867
rect 18177 27833 18211 27867
rect 18253 27833 18287 27867
rect 18329 27833 18363 27867
rect 18405 27833 18439 27867
rect 18486 27849 18520 27883
rect 18556 27849 18590 27883
rect 18626 27849 18660 27883
rect 18696 27849 18730 27883
rect 18766 27849 18800 27883
rect 18836 27849 18870 27883
rect 18906 27849 18940 27883
rect 18976 27849 19010 27883
rect 18025 27765 18059 27799
rect 18101 27765 18135 27799
rect 18177 27765 18211 27799
rect 18253 27765 18287 27799
rect 18329 27765 18363 27799
rect 18405 27765 18439 27799
rect 18486 27781 18520 27815
rect 18556 27781 18590 27815
rect 18626 27781 18660 27815
rect 18696 27781 18730 27815
rect 18766 27781 18800 27815
rect 18836 27781 18870 27815
rect 18906 27781 18940 27815
rect 18976 27781 19010 27815
rect 18025 27697 18059 27731
rect 18101 27697 18135 27731
rect 18177 27697 18211 27731
rect 18253 27697 18287 27731
rect 18329 27697 18363 27731
rect 18405 27697 18439 27731
rect 18486 27713 18520 27747
rect 18556 27713 18590 27747
rect 18626 27713 18660 27747
rect 18696 27713 18730 27747
rect 18766 27713 18800 27747
rect 18836 27713 18870 27747
rect 18906 27713 18940 27747
rect 18976 27713 19010 27747
rect 18025 27629 18059 27663
rect 18101 27629 18135 27663
rect 18177 27629 18211 27663
rect 18253 27629 18287 27663
rect 18329 27629 18363 27663
rect 18405 27629 18439 27663
rect 18486 27645 18520 27679
rect 18556 27645 18590 27679
rect 18626 27645 18660 27679
rect 18696 27645 18730 27679
rect 18766 27645 18800 27679
rect 18836 27645 18870 27679
rect 18906 27645 18940 27679
rect 18976 27645 19010 27679
rect 18025 27561 18059 27595
rect 18101 27561 18135 27595
rect 18177 27561 18211 27595
rect 18253 27561 18287 27595
rect 18329 27561 18363 27595
rect 18405 27561 18439 27595
rect 18486 27577 18520 27611
rect 18556 27577 18590 27611
rect 18626 27577 18660 27611
rect 18696 27577 18730 27611
rect 18766 27577 18800 27611
rect 18836 27577 18870 27611
rect 18906 27577 18940 27611
rect 18976 27577 19010 27611
rect 18025 27493 18059 27527
rect 18101 27493 18135 27527
rect 18177 27493 18211 27527
rect 18253 27493 18287 27527
rect 18329 27493 18363 27527
rect 18405 27493 18439 27527
rect 18486 27509 18520 27543
rect 18556 27509 18590 27543
rect 18626 27509 18660 27543
rect 18696 27509 18730 27543
rect 18766 27509 18800 27543
rect 18836 27509 18870 27543
rect 18906 27509 18940 27543
rect 18976 27509 19010 27543
rect 18025 27425 18059 27459
rect 18101 27425 18135 27459
rect 18177 27425 18211 27459
rect 18253 27425 18287 27459
rect 18329 27425 18363 27459
rect 18405 27425 18439 27459
rect 18486 27441 18520 27475
rect 18556 27441 18590 27475
rect 18626 27441 18660 27475
rect 18696 27441 18730 27475
rect 18766 27441 18800 27475
rect 18836 27441 18870 27475
rect 18906 27441 18940 27475
rect 18976 27441 19010 27475
rect 18025 27357 18059 27391
rect 18101 27357 18135 27391
rect 18177 27357 18211 27391
rect 18253 27357 18287 27391
rect 18329 27357 18363 27391
rect 18405 27357 18439 27391
rect 18486 27373 18520 27407
rect 18556 27373 18590 27407
rect 18626 27373 18660 27407
rect 18696 27373 18730 27407
rect 18766 27373 18800 27407
rect 18836 27373 18870 27407
rect 18906 27373 18940 27407
rect 18976 27373 19010 27407
rect 18025 27289 18059 27323
rect 18101 27289 18135 27323
rect 18177 27289 18211 27323
rect 18253 27289 18287 27323
rect 18329 27289 18363 27323
rect 18405 27289 18439 27323
rect 18486 27305 18520 27339
rect 18556 27305 18590 27339
rect 18626 27305 18660 27339
rect 18696 27305 18730 27339
rect 18766 27305 18800 27339
rect 18836 27305 18870 27339
rect 18906 27305 18940 27339
rect 18976 27305 19010 27339
rect 18025 27221 18059 27255
rect 18101 27221 18135 27255
rect 18177 27221 18211 27255
rect 18253 27221 18287 27255
rect 18329 27221 18363 27255
rect 18405 27221 18439 27255
rect 18486 27237 18520 27271
rect 18556 27237 18590 27271
rect 18626 27237 18660 27271
rect 18696 27237 18730 27271
rect 18766 27237 18800 27271
rect 18836 27237 18870 27271
rect 18906 27237 18940 27271
rect 18976 27237 19010 27271
rect 18025 27153 18059 27187
rect 18101 27153 18135 27187
rect 18177 27153 18211 27187
rect 18253 27153 18287 27187
rect 18329 27153 18363 27187
rect 18405 27153 18439 27187
rect 18486 27169 18520 27203
rect 18556 27169 18590 27203
rect 18626 27169 18660 27203
rect 18696 27169 18730 27203
rect 18766 27169 18800 27203
rect 18836 27169 18870 27203
rect 18906 27169 18940 27203
rect 18976 27169 19010 27203
rect 1057 27045 1091 27079
rect 1125 27045 1159 27079
rect 1193 27045 1227 27079
rect 1261 27045 1295 27079
rect 1329 27045 1363 27079
rect 1397 27045 1431 27079
rect 1465 27045 1499 27079
rect 1533 27045 1567 27079
rect 1601 27045 1635 27079
rect 1669 27045 1703 27079
rect 1057 26976 1091 27010
rect 1125 26976 1159 27010
rect 1193 26976 1227 27010
rect 1261 26976 1295 27010
rect 1329 26976 1363 27010
rect 1397 26976 1431 27010
rect 1465 26976 1499 27010
rect 1533 26976 1567 27010
rect 1601 26976 1635 27010
rect 1669 26976 1703 27010
rect 1057 26907 1091 26941
rect 1125 26907 1159 26941
rect 1193 26907 1227 26941
rect 1261 26907 1295 26941
rect 1329 26907 1363 26941
rect 1397 26907 1431 26941
rect 1465 26907 1499 26941
rect 1533 26907 1567 26941
rect 1601 26907 1635 26941
rect 1669 26907 1703 26941
rect 1057 26838 1091 26872
rect 1125 26838 1159 26872
rect 1193 26838 1227 26872
rect 1261 26838 1295 26872
rect 1329 26838 1363 26872
rect 1397 26838 1431 26872
rect 1465 26838 1499 26872
rect 1533 26838 1567 26872
rect 1601 26838 1635 26872
rect 1669 26838 1703 26872
rect 1057 26769 1091 26803
rect 1125 26769 1159 26803
rect 1193 26769 1227 26803
rect 1261 26769 1295 26803
rect 1329 26769 1363 26803
rect 1397 26769 1431 26803
rect 1465 26769 1499 26803
rect 1533 26769 1567 26803
rect 1601 26769 1635 26803
rect 1669 26769 1703 26803
rect 1057 26700 1091 26734
rect 1125 26700 1159 26734
rect 1193 26700 1227 26734
rect 1261 26700 1295 26734
rect 1329 26700 1363 26734
rect 1397 26700 1431 26734
rect 1465 26700 1499 26734
rect 1533 26700 1567 26734
rect 1601 26700 1635 26734
rect 1669 26700 1703 26734
rect 1057 26631 1091 26665
rect 1125 26631 1159 26665
rect 1193 26631 1227 26665
rect 1261 26631 1295 26665
rect 1329 26631 1363 26665
rect 1397 26631 1431 26665
rect 1465 26631 1499 26665
rect 1533 26631 1567 26665
rect 1601 26631 1635 26665
rect 1669 26631 1703 26665
rect 1057 26562 1091 26596
rect 1125 26562 1159 26596
rect 1193 26562 1227 26596
rect 1261 26562 1295 26596
rect 1329 26562 1363 26596
rect 1397 26562 1431 26596
rect 1465 26562 1499 26596
rect 1533 26562 1567 26596
rect 1601 26562 1635 26596
rect 1669 26562 1703 26596
rect 1057 26493 1091 26527
rect 1125 26493 1159 26527
rect 1193 26493 1227 26527
rect 1261 26493 1295 26527
rect 1329 26493 1363 26527
rect 1397 26493 1431 26527
rect 1465 26493 1499 26527
rect 1533 26493 1567 26527
rect 1601 26493 1635 26527
rect 1669 26493 1703 26527
rect 1057 26424 1091 26458
rect 1125 26424 1159 26458
rect 1193 26424 1227 26458
rect 1261 26424 1295 26458
rect 1329 26424 1363 26458
rect 1397 26424 1431 26458
rect 1465 26424 1499 26458
rect 1533 26424 1567 26458
rect 1601 26424 1635 26458
rect 1669 26424 1703 26458
rect 1057 26355 1091 26389
rect 1125 26355 1159 26389
rect 1193 26355 1227 26389
rect 1261 26355 1295 26389
rect 1329 26355 1363 26389
rect 1397 26355 1431 26389
rect 1465 26355 1499 26389
rect 1533 26355 1567 26389
rect 1601 26355 1635 26389
rect 1669 26355 1703 26389
rect 1057 26286 1091 26320
rect 1125 26286 1159 26320
rect 1193 26286 1227 26320
rect 1261 26286 1295 26320
rect 1329 26286 1363 26320
rect 1397 26286 1431 26320
rect 1465 26286 1499 26320
rect 1533 26286 1567 26320
rect 1601 26286 1635 26320
rect 1669 26286 1703 26320
rect 1057 26217 1091 26251
rect 1125 26217 1159 26251
rect 1193 26217 1227 26251
rect 1261 26217 1295 26251
rect 1329 26217 1363 26251
rect 1397 26217 1431 26251
rect 1465 26217 1499 26251
rect 1533 26217 1567 26251
rect 1601 26217 1635 26251
rect 1669 26217 1703 26251
rect 1057 26148 1091 26182
rect 1125 26148 1159 26182
rect 1193 26148 1227 26182
rect 1261 26148 1295 26182
rect 1329 26148 1363 26182
rect 1397 26148 1431 26182
rect 1465 26148 1499 26182
rect 1533 26148 1567 26182
rect 1601 26148 1635 26182
rect 1669 26148 1703 26182
rect 1057 26079 1091 26113
rect 1125 26079 1159 26113
rect 1193 26079 1227 26113
rect 1261 26079 1295 26113
rect 1329 26079 1363 26113
rect 1397 26079 1431 26113
rect 1465 26079 1499 26113
rect 1533 26079 1567 26113
rect 1601 26079 1635 26113
rect 1669 26079 1703 26113
rect 1057 26010 1091 26044
rect 1125 26010 1159 26044
rect 1193 26010 1227 26044
rect 1261 26010 1295 26044
rect 1329 26010 1363 26044
rect 1397 26010 1431 26044
rect 1465 26010 1499 26044
rect 1533 26010 1567 26044
rect 1601 26010 1635 26044
rect 1669 26010 1703 26044
rect 1057 25941 1091 25975
rect 1125 25941 1159 25975
rect 1193 25941 1227 25975
rect 1261 25941 1295 25975
rect 1329 25941 1363 25975
rect 1397 25941 1431 25975
rect 1465 25941 1499 25975
rect 1533 25941 1567 25975
rect 1601 25941 1635 25975
rect 1669 25941 1703 25975
rect 1057 25872 1091 25906
rect 1125 25872 1159 25906
rect 1193 25872 1227 25906
rect 1261 25872 1295 25906
rect 1329 25872 1363 25906
rect 1397 25872 1431 25906
rect 1465 25872 1499 25906
rect 1533 25872 1567 25906
rect 1601 25872 1635 25906
rect 1669 25872 1703 25906
rect 1057 25803 1091 25837
rect 1125 25803 1159 25837
rect 1193 25803 1227 25837
rect 1261 25803 1295 25837
rect 1329 25803 1363 25837
rect 1397 25803 1431 25837
rect 1465 25803 1499 25837
rect 1533 25803 1567 25837
rect 1601 25803 1635 25837
rect 1669 25803 1703 25837
rect 1057 25734 1091 25768
rect 1125 25734 1159 25768
rect 1193 25734 1227 25768
rect 1261 25734 1295 25768
rect 1329 25734 1363 25768
rect 1397 25734 1431 25768
rect 1465 25734 1499 25768
rect 1533 25734 1567 25768
rect 1601 25734 1635 25768
rect 1669 25734 1703 25768
rect 1057 25665 1091 25699
rect 1125 25665 1159 25699
rect 1193 25665 1227 25699
rect 1261 25665 1295 25699
rect 1329 25665 1363 25699
rect 1397 25665 1431 25699
rect 1465 25665 1499 25699
rect 1533 25665 1567 25699
rect 1601 25665 1635 25699
rect 1669 25665 1703 25699
rect 1057 25596 1091 25630
rect 1125 25596 1159 25630
rect 1193 25596 1227 25630
rect 1261 25596 1295 25630
rect 1329 25596 1363 25630
rect 1397 25596 1431 25630
rect 1465 25596 1499 25630
rect 1533 25596 1567 25630
rect 1601 25596 1635 25630
rect 1669 25596 1703 25630
rect 1057 25527 1091 25561
rect 1125 25527 1159 25561
rect 1193 25527 1227 25561
rect 1261 25527 1295 25561
rect 1329 25527 1363 25561
rect 1397 25527 1431 25561
rect 1465 25527 1499 25561
rect 1533 25527 1567 25561
rect 1601 25527 1635 25561
rect 1669 25527 1703 25561
rect 1057 25458 1091 25492
rect 1125 25458 1159 25492
rect 1193 25458 1227 25492
rect 1261 25458 1295 25492
rect 1329 25458 1363 25492
rect 1397 25458 1431 25492
rect 1465 25458 1499 25492
rect 1533 25458 1567 25492
rect 1601 25458 1635 25492
rect 1669 25458 1703 25492
rect 1057 25389 1091 25423
rect 1125 25389 1159 25423
rect 1193 25389 1227 25423
rect 1261 25389 1295 25423
rect 1329 25389 1363 25423
rect 1397 25389 1431 25423
rect 1465 25389 1499 25423
rect 1533 25389 1567 25423
rect 1601 25389 1635 25423
rect 1669 25389 1703 25423
rect 1057 25320 1091 25354
rect 1125 25320 1159 25354
rect 1193 25320 1227 25354
rect 1261 25320 1295 25354
rect 1329 25320 1363 25354
rect 1397 25320 1431 25354
rect 1465 25320 1499 25354
rect 1533 25320 1567 25354
rect 1601 25320 1635 25354
rect 1669 25320 1703 25354
rect 1057 25251 1091 25285
rect 1125 25251 1159 25285
rect 1193 25251 1227 25285
rect 1261 25251 1295 25285
rect 1329 25251 1363 25285
rect 1397 25251 1431 25285
rect 1465 25251 1499 25285
rect 1533 25251 1567 25285
rect 1601 25251 1635 25285
rect 1669 25251 1703 25285
rect 1057 25182 1091 25216
rect 1125 25182 1159 25216
rect 1193 25182 1227 25216
rect 1261 25182 1295 25216
rect 1329 25182 1363 25216
rect 1397 25182 1431 25216
rect 1465 25182 1499 25216
rect 1533 25182 1567 25216
rect 1601 25182 1635 25216
rect 1669 25182 1703 25216
rect 1057 25113 1091 25147
rect 1125 25113 1159 25147
rect 1193 25113 1227 25147
rect 1261 25113 1295 25147
rect 1329 25113 1363 25147
rect 1397 25113 1431 25147
rect 1465 25113 1499 25147
rect 1533 25113 1567 25147
rect 1601 25113 1635 25147
rect 1669 25113 1703 25147
rect 1057 25043 1091 25077
rect 1125 25043 1159 25077
rect 1193 25043 1227 25077
rect 1261 25043 1295 25077
rect 1329 25043 1363 25077
rect 1397 25043 1431 25077
rect 1465 25043 1499 25077
rect 1533 25043 1567 25077
rect 1601 25043 1635 25077
rect 1669 25043 1703 25077
rect 1057 24973 1091 25007
rect 1125 24973 1159 25007
rect 1193 24973 1227 25007
rect 1261 24973 1295 25007
rect 1329 24973 1363 25007
rect 1397 24973 1431 25007
rect 1465 24973 1499 25007
rect 1533 24973 1567 25007
rect 1601 24973 1635 25007
rect 1669 24973 1703 25007
rect 1057 24903 1091 24937
rect 1125 24903 1159 24937
rect 1193 24903 1227 24937
rect 1261 24903 1295 24937
rect 1329 24903 1363 24937
rect 1397 24903 1431 24937
rect 1465 24903 1499 24937
rect 1533 24903 1567 24937
rect 1601 24903 1635 24937
rect 1669 24903 1703 24937
rect 1057 24833 1091 24867
rect 1125 24833 1159 24867
rect 1193 24833 1227 24867
rect 1261 24833 1295 24867
rect 1329 24833 1363 24867
rect 1397 24833 1431 24867
rect 1465 24833 1499 24867
rect 1533 24833 1567 24867
rect 1601 24833 1635 24867
rect 1669 24833 1703 24867
rect 1057 24763 1091 24797
rect 1125 24763 1159 24797
rect 1193 24763 1227 24797
rect 1261 24763 1295 24797
rect 1329 24763 1363 24797
rect 1397 24763 1431 24797
rect 1465 24763 1499 24797
rect 1533 24763 1567 24797
rect 1601 24763 1635 24797
rect 1669 24763 1703 24797
rect 1057 24693 1091 24727
rect 1125 24693 1159 24727
rect 1193 24693 1227 24727
rect 1261 24693 1295 24727
rect 1329 24693 1363 24727
rect 1397 24693 1431 24727
rect 1465 24693 1499 24727
rect 1533 24693 1567 24727
rect 1601 24693 1635 24727
rect 1669 24693 1703 24727
rect 1057 24623 1091 24657
rect 1125 24623 1159 24657
rect 1193 24623 1227 24657
rect 1261 24623 1295 24657
rect 1329 24623 1363 24657
rect 1397 24623 1431 24657
rect 1465 24623 1499 24657
rect 1533 24623 1567 24657
rect 1601 24623 1635 24657
rect 1669 24623 1703 24657
rect 1057 24553 1091 24587
rect 1125 24553 1159 24587
rect 1193 24553 1227 24587
rect 1261 24553 1295 24587
rect 1329 24553 1363 24587
rect 1397 24553 1431 24587
rect 1465 24553 1499 24587
rect 1533 24553 1567 24587
rect 1601 24553 1635 24587
rect 1669 24553 1703 24587
rect 1057 24483 1091 24517
rect 1125 24483 1159 24517
rect 1193 24483 1227 24517
rect 1261 24483 1295 24517
rect 1329 24483 1363 24517
rect 1397 24483 1431 24517
rect 1465 24483 1499 24517
rect 1533 24483 1567 24517
rect 1601 24483 1635 24517
rect 1669 24483 1703 24517
rect 1057 24413 1091 24447
rect 1125 24413 1159 24447
rect 1193 24413 1227 24447
rect 1261 24413 1295 24447
rect 1329 24413 1363 24447
rect 1397 24413 1431 24447
rect 1465 24413 1499 24447
rect 1533 24413 1567 24447
rect 1601 24413 1635 24447
rect 1669 24413 1703 24447
rect 1057 24343 1091 24377
rect 1125 24343 1159 24377
rect 1193 24343 1227 24377
rect 1261 24343 1295 24377
rect 1329 24343 1363 24377
rect 1397 24343 1431 24377
rect 1465 24343 1499 24377
rect 1533 24343 1567 24377
rect 1601 24343 1635 24377
rect 1669 24343 1703 24377
rect 1057 24273 1091 24307
rect 1125 24273 1159 24307
rect 1193 24273 1227 24307
rect 1261 24273 1295 24307
rect 1329 24273 1363 24307
rect 1397 24273 1431 24307
rect 1465 24273 1499 24307
rect 1533 24273 1567 24307
rect 1601 24273 1635 24307
rect 1669 24273 1703 24307
rect 1057 24203 1091 24237
rect 1125 24203 1159 24237
rect 1193 24203 1227 24237
rect 1261 24203 1295 24237
rect 1329 24203 1363 24237
rect 1397 24203 1431 24237
rect 1465 24203 1499 24237
rect 1533 24203 1567 24237
rect 1601 24203 1635 24237
rect 1669 24203 1703 24237
rect 1057 24133 1091 24167
rect 1125 24133 1159 24167
rect 1193 24133 1227 24167
rect 1261 24133 1295 24167
rect 1329 24133 1363 24167
rect 1397 24133 1431 24167
rect 1465 24133 1499 24167
rect 1533 24133 1567 24167
rect 1601 24133 1635 24167
rect 1669 24133 1703 24167
rect 1057 24063 1091 24097
rect 1125 24063 1159 24097
rect 1193 24063 1227 24097
rect 1261 24063 1295 24097
rect 1329 24063 1363 24097
rect 1397 24063 1431 24097
rect 1465 24063 1499 24097
rect 1533 24063 1567 24097
rect 1601 24063 1635 24097
rect 1669 24063 1703 24097
rect 1057 23993 1091 24027
rect 1125 23993 1159 24027
rect 1193 23993 1227 24027
rect 1261 23993 1295 24027
rect 1329 23993 1363 24027
rect 1397 23993 1431 24027
rect 1465 23993 1499 24027
rect 1533 23993 1567 24027
rect 1601 23993 1635 24027
rect 1669 23993 1703 24027
rect 1057 23923 1091 23957
rect 1125 23923 1159 23957
rect 1193 23923 1227 23957
rect 1261 23923 1295 23957
rect 1329 23923 1363 23957
rect 1397 23923 1431 23957
rect 1465 23923 1499 23957
rect 1533 23923 1567 23957
rect 1601 23923 1635 23957
rect 1669 23923 1703 23957
rect 1057 23853 1091 23887
rect 1125 23853 1159 23887
rect 1193 23853 1227 23887
rect 1261 23853 1295 23887
rect 1329 23853 1363 23887
rect 1397 23853 1431 23887
rect 1465 23853 1499 23887
rect 1533 23853 1567 23887
rect 1601 23853 1635 23887
rect 1669 23853 1703 23887
rect 18025 27085 18059 27119
rect 18101 27085 18135 27119
rect 18177 27085 18211 27119
rect 18253 27085 18287 27119
rect 18329 27085 18363 27119
rect 18405 27085 18439 27119
rect 18486 27101 18520 27135
rect 18556 27101 18590 27135
rect 18626 27101 18660 27135
rect 18696 27101 18730 27135
rect 18766 27101 18800 27135
rect 18836 27101 18870 27135
rect 18906 27101 18940 27135
rect 18976 27101 19010 27135
rect 18025 27017 18059 27051
rect 18101 27017 18135 27051
rect 18177 27017 18211 27051
rect 18253 27017 18287 27051
rect 18329 27017 18363 27051
rect 18405 27017 18439 27051
rect 18486 27033 18520 27067
rect 18556 27033 18590 27067
rect 18626 27033 18660 27067
rect 18696 27033 18730 27067
rect 18766 27033 18800 27067
rect 18836 27033 18870 27067
rect 18906 27033 18940 27067
rect 18976 27033 19010 27067
rect 18025 26949 18059 26983
rect 18101 26949 18135 26983
rect 18177 26949 18211 26983
rect 18253 26949 18287 26983
rect 18329 26949 18363 26983
rect 18405 26949 18439 26983
rect 18486 26965 18520 26999
rect 18556 26965 18590 26999
rect 18626 26965 18660 26999
rect 18696 26965 18730 26999
rect 18766 26965 18800 26999
rect 18836 26965 18870 26999
rect 18906 26965 18940 26999
rect 18976 26965 19010 26999
rect 18025 26881 18059 26915
rect 18101 26881 18135 26915
rect 18177 26881 18211 26915
rect 18253 26881 18287 26915
rect 18329 26881 18363 26915
rect 18405 26881 18439 26915
rect 18486 26897 18520 26931
rect 18556 26897 18590 26931
rect 18626 26897 18660 26931
rect 18696 26897 18730 26931
rect 18766 26897 18800 26931
rect 18836 26897 18870 26931
rect 18906 26897 18940 26931
rect 18976 26897 19010 26931
rect 18025 26813 18059 26847
rect 18101 26813 18135 26847
rect 18177 26813 18211 26847
rect 18253 26813 18287 26847
rect 18329 26813 18363 26847
rect 18405 26813 18439 26847
rect 18486 26829 18520 26863
rect 18556 26829 18590 26863
rect 18626 26829 18660 26863
rect 18696 26829 18730 26863
rect 18766 26829 18800 26863
rect 18836 26829 18870 26863
rect 18906 26829 18940 26863
rect 18976 26829 19010 26863
rect 18025 26745 18059 26779
rect 18101 26745 18135 26779
rect 18177 26745 18211 26779
rect 18253 26745 18287 26779
rect 18329 26745 18363 26779
rect 18405 26745 18439 26779
rect 18486 26761 18520 26795
rect 18556 26761 18590 26795
rect 18626 26761 18660 26795
rect 18696 26761 18730 26795
rect 18766 26761 18800 26795
rect 18836 26761 18870 26795
rect 18906 26761 18940 26795
rect 18976 26761 19010 26795
rect 18025 26677 18059 26711
rect 18101 26677 18135 26711
rect 18177 26677 18211 26711
rect 18253 26677 18287 26711
rect 18329 26677 18363 26711
rect 18405 26677 18439 26711
rect 18486 26693 18520 26727
rect 18556 26693 18590 26727
rect 18626 26693 18660 26727
rect 18696 26693 18730 26727
rect 18766 26693 18800 26727
rect 18836 26693 18870 26727
rect 18906 26693 18940 26727
rect 18976 26693 19010 26727
rect 18025 26609 18059 26643
rect 18101 26609 18135 26643
rect 18177 26609 18211 26643
rect 18253 26609 18287 26643
rect 18329 26609 18363 26643
rect 18405 26609 18439 26643
rect 18486 26625 18520 26659
rect 18556 26625 18590 26659
rect 18626 26625 18660 26659
rect 18696 26625 18730 26659
rect 18766 26625 18800 26659
rect 18836 26625 18870 26659
rect 18906 26625 18940 26659
rect 18976 26625 19010 26659
rect 18025 26541 18059 26575
rect 18101 26541 18135 26575
rect 18177 26541 18211 26575
rect 18253 26541 18287 26575
rect 18329 26541 18363 26575
rect 18405 26541 18439 26575
rect 18486 26557 18520 26591
rect 18556 26557 18590 26591
rect 18626 26557 18660 26591
rect 18696 26557 18730 26591
rect 18766 26557 18800 26591
rect 18836 26557 18870 26591
rect 18906 26557 18940 26591
rect 18976 26557 19010 26591
rect 18025 26473 18059 26507
rect 18101 26473 18135 26507
rect 18177 26473 18211 26507
rect 18253 26473 18287 26507
rect 18329 26473 18363 26507
rect 18405 26473 18439 26507
rect 18486 26489 18520 26523
rect 18556 26489 18590 26523
rect 18626 26489 18660 26523
rect 18696 26489 18730 26523
rect 18766 26489 18800 26523
rect 18836 26489 18870 26523
rect 18906 26489 18940 26523
rect 18976 26489 19010 26523
rect 18025 26405 18059 26439
rect 18101 26405 18135 26439
rect 18177 26405 18211 26439
rect 18253 26405 18287 26439
rect 18329 26405 18363 26439
rect 18405 26405 18439 26439
rect 18486 26421 18520 26455
rect 18556 26421 18590 26455
rect 18626 26421 18660 26455
rect 18696 26421 18730 26455
rect 18766 26421 18800 26455
rect 18836 26421 18870 26455
rect 18906 26421 18940 26455
rect 18976 26421 19010 26455
rect 18025 26337 18059 26371
rect 18101 26337 18135 26371
rect 18177 26337 18211 26371
rect 18253 26337 18287 26371
rect 18329 26337 18363 26371
rect 18405 26337 18439 26371
rect 18486 26353 18520 26387
rect 18556 26353 18590 26387
rect 18626 26353 18660 26387
rect 18696 26353 18730 26387
rect 18766 26353 18800 26387
rect 18836 26353 18870 26387
rect 18906 26353 18940 26387
rect 18976 26353 19010 26387
rect 18025 26269 18059 26303
rect 18101 26269 18135 26303
rect 18177 26269 18211 26303
rect 18253 26269 18287 26303
rect 18329 26269 18363 26303
rect 18405 26269 18439 26303
rect 18486 26285 18520 26319
rect 18556 26285 18590 26319
rect 18626 26285 18660 26319
rect 18696 26285 18730 26319
rect 18766 26285 18800 26319
rect 18836 26285 18870 26319
rect 18906 26285 18940 26319
rect 18976 26285 19010 26319
rect 18025 26201 18059 26235
rect 18101 26201 18135 26235
rect 18177 26201 18211 26235
rect 18253 26201 18287 26235
rect 18329 26201 18363 26235
rect 18405 26201 18439 26235
rect 18486 26217 18520 26251
rect 18556 26217 18590 26251
rect 18626 26217 18660 26251
rect 18696 26217 18730 26251
rect 18766 26217 18800 26251
rect 18836 26217 18870 26251
rect 18906 26217 18940 26251
rect 18976 26217 19010 26251
rect 18025 26133 18059 26167
rect 18101 26133 18135 26167
rect 18177 26133 18211 26167
rect 18253 26133 18287 26167
rect 18329 26133 18363 26167
rect 18405 26133 18439 26167
rect 18486 26149 18520 26183
rect 18556 26149 18590 26183
rect 18626 26149 18660 26183
rect 18696 26149 18730 26183
rect 18766 26149 18800 26183
rect 18836 26149 18870 26183
rect 18906 26149 18940 26183
rect 18976 26149 19010 26183
rect 18025 26065 18059 26099
rect 18101 26065 18135 26099
rect 18177 26065 18211 26099
rect 18253 26065 18287 26099
rect 18329 26065 18363 26099
rect 18405 26065 18439 26099
rect 18486 26081 18520 26115
rect 18556 26081 18590 26115
rect 18626 26081 18660 26115
rect 18696 26081 18730 26115
rect 18766 26081 18800 26115
rect 18836 26081 18870 26115
rect 18906 26081 18940 26115
rect 18976 26081 19010 26115
rect 18025 25997 18059 26031
rect 18101 25997 18135 26031
rect 18177 25997 18211 26031
rect 18253 25997 18287 26031
rect 18329 25997 18363 26031
rect 18405 25997 18439 26031
rect 18486 26013 18520 26047
rect 18556 26013 18590 26047
rect 18626 26013 18660 26047
rect 18696 26013 18730 26047
rect 18766 26013 18800 26047
rect 18836 26013 18870 26047
rect 18906 26013 18940 26047
rect 18976 26013 19010 26047
rect 18025 25929 18059 25963
rect 18101 25929 18135 25963
rect 18177 25929 18211 25963
rect 18253 25929 18287 25963
rect 18329 25929 18363 25963
rect 18405 25929 18439 25963
rect 18486 25945 18520 25979
rect 18556 25945 18590 25979
rect 18626 25945 18660 25979
rect 18696 25945 18730 25979
rect 18766 25945 18800 25979
rect 18836 25945 18870 25979
rect 18906 25945 18940 25979
rect 18976 25945 19010 25979
rect 18025 25861 18059 25895
rect 18101 25861 18135 25895
rect 18177 25861 18211 25895
rect 18253 25861 18287 25895
rect 18329 25861 18363 25895
rect 18405 25861 18439 25895
rect 18486 25877 18520 25911
rect 18556 25877 18590 25911
rect 18626 25877 18660 25911
rect 18696 25877 18730 25911
rect 18766 25877 18800 25911
rect 18836 25877 18870 25911
rect 18906 25877 18940 25911
rect 18976 25877 19010 25911
rect 18025 25793 18059 25827
rect 18101 25793 18135 25827
rect 18177 25793 18211 25827
rect 18253 25793 18287 25827
rect 18329 25793 18363 25827
rect 18405 25793 18439 25827
rect 18486 25809 18520 25843
rect 18556 25809 18590 25843
rect 18626 25809 18660 25843
rect 18696 25809 18730 25843
rect 18766 25809 18800 25843
rect 18836 25809 18870 25843
rect 18906 25809 18940 25843
rect 18976 25809 19010 25843
rect 18025 25725 18059 25759
rect 18101 25725 18135 25759
rect 18177 25725 18211 25759
rect 18253 25725 18287 25759
rect 18329 25725 18363 25759
rect 18405 25725 18439 25759
rect 18486 25741 18520 25775
rect 18556 25741 18590 25775
rect 18626 25741 18660 25775
rect 18696 25741 18730 25775
rect 18766 25741 18800 25775
rect 18836 25741 18870 25775
rect 18906 25741 18940 25775
rect 18976 25741 19010 25775
rect 18025 25657 18059 25691
rect 18101 25657 18135 25691
rect 18177 25657 18211 25691
rect 18253 25657 18287 25691
rect 18329 25657 18363 25691
rect 18405 25657 18439 25691
rect 18486 25673 18520 25707
rect 18556 25673 18590 25707
rect 18626 25673 18660 25707
rect 18696 25673 18730 25707
rect 18766 25673 18800 25707
rect 18836 25673 18870 25707
rect 18906 25673 18940 25707
rect 18976 25673 19010 25707
rect 18025 25589 18059 25623
rect 18101 25589 18135 25623
rect 18177 25589 18211 25623
rect 18253 25589 18287 25623
rect 18329 25589 18363 25623
rect 18405 25589 18439 25623
rect 18486 25604 18520 25638
rect 18556 25604 18590 25638
rect 18626 25604 18660 25638
rect 18696 25604 18730 25638
rect 18766 25604 18800 25638
rect 18836 25604 18870 25638
rect 18906 25604 18940 25638
rect 18976 25604 19010 25638
rect 18025 25521 18059 25555
rect 18101 25521 18135 25555
rect 18177 25521 18211 25555
rect 18253 25521 18287 25555
rect 18329 25521 18363 25555
rect 18405 25521 18439 25555
rect 18486 25535 18520 25569
rect 18556 25535 18590 25569
rect 18626 25535 18660 25569
rect 18696 25535 18730 25569
rect 18766 25535 18800 25569
rect 18836 25535 18870 25569
rect 18906 25535 18940 25569
rect 18976 25535 19010 25569
rect 18025 25453 18059 25487
rect 18101 25453 18135 25487
rect 18177 25453 18211 25487
rect 18253 25453 18287 25487
rect 18329 25453 18363 25487
rect 18405 25453 18439 25487
rect 18486 25466 18520 25500
rect 18556 25466 18590 25500
rect 18626 25466 18660 25500
rect 18696 25466 18730 25500
rect 18766 25466 18800 25500
rect 18836 25466 18870 25500
rect 18906 25466 18940 25500
rect 18976 25466 19010 25500
rect 18025 25385 18059 25419
rect 18101 25385 18135 25419
rect 18177 25385 18211 25419
rect 18253 25385 18287 25419
rect 18329 25385 18363 25419
rect 18405 25385 18439 25419
rect 18486 25397 18520 25431
rect 18556 25397 18590 25431
rect 18626 25397 18660 25431
rect 18696 25397 18730 25431
rect 18766 25397 18800 25431
rect 18836 25397 18870 25431
rect 18906 25397 18940 25431
rect 18976 25397 19010 25431
rect 18025 25317 18059 25351
rect 18101 25317 18135 25351
rect 18177 25317 18211 25351
rect 18253 25317 18287 25351
rect 18329 25317 18363 25351
rect 18405 25317 18439 25351
rect 18486 25328 18520 25362
rect 18556 25328 18590 25362
rect 18626 25328 18660 25362
rect 18696 25328 18730 25362
rect 18766 25328 18800 25362
rect 18836 25328 18870 25362
rect 18906 25328 18940 25362
rect 18976 25328 19010 25362
rect 18025 25249 18059 25283
rect 18101 25249 18135 25283
rect 18177 25249 18211 25283
rect 18253 25249 18287 25283
rect 18329 25249 18363 25283
rect 18405 25249 18439 25283
rect 18486 25259 18520 25293
rect 18556 25259 18590 25293
rect 18626 25259 18660 25293
rect 18696 25259 18730 25293
rect 18766 25259 18800 25293
rect 18836 25259 18870 25293
rect 18906 25259 18940 25293
rect 18976 25259 19010 25293
rect 18025 25180 18059 25214
rect 18101 25180 18135 25214
rect 18177 25180 18211 25214
rect 18253 25180 18287 25214
rect 18329 25180 18363 25214
rect 18405 25180 18439 25214
rect 18486 25190 18520 25224
rect 18556 25190 18590 25224
rect 18626 25190 18660 25224
rect 18696 25190 18730 25224
rect 18766 25190 18800 25224
rect 18836 25190 18870 25224
rect 18906 25190 18940 25224
rect 18976 25190 19010 25224
rect 18025 25111 18059 25145
rect 18101 25111 18135 25145
rect 18177 25111 18211 25145
rect 18253 25111 18287 25145
rect 18329 25111 18363 25145
rect 18405 25111 18439 25145
rect 18486 25121 18520 25155
rect 18556 25121 18590 25155
rect 18626 25121 18660 25155
rect 18696 25121 18730 25155
rect 18766 25121 18800 25155
rect 18836 25121 18870 25155
rect 18906 25121 18940 25155
rect 18976 25121 19010 25155
rect 18025 25042 18059 25076
rect 18101 25042 18135 25076
rect 18177 25042 18211 25076
rect 18253 25042 18287 25076
rect 18329 25042 18363 25076
rect 18405 25042 18439 25076
rect 18486 25052 18520 25086
rect 18556 25052 18590 25086
rect 18626 25052 18660 25086
rect 18696 25052 18730 25086
rect 18766 25052 18800 25086
rect 18836 25052 18870 25086
rect 18906 25052 18940 25086
rect 18976 25052 19010 25086
rect 18025 24973 18059 25007
rect 18101 24973 18135 25007
rect 18177 24973 18211 25007
rect 18253 24973 18287 25007
rect 18329 24973 18363 25007
rect 18405 24973 18439 25007
rect 18486 24983 18520 25017
rect 18556 24983 18590 25017
rect 18626 24983 18660 25017
rect 18696 24983 18730 25017
rect 18766 24983 18800 25017
rect 18836 24983 18870 25017
rect 18906 24983 18940 25017
rect 18976 24983 19010 25017
rect 18025 24904 18059 24938
rect 18101 24904 18135 24938
rect 18177 24904 18211 24938
rect 18253 24904 18287 24938
rect 18329 24904 18363 24938
rect 18405 24904 18439 24938
rect 18486 24914 18520 24948
rect 18556 24914 18590 24948
rect 18626 24914 18660 24948
rect 18696 24914 18730 24948
rect 18766 24914 18800 24948
rect 18836 24914 18870 24948
rect 18906 24914 18940 24948
rect 18976 24914 19010 24948
rect 18025 24835 18059 24869
rect 18101 24835 18135 24869
rect 18177 24835 18211 24869
rect 18253 24835 18287 24869
rect 18329 24835 18363 24869
rect 18405 24835 18439 24869
rect 18486 24845 18520 24879
rect 18556 24845 18590 24879
rect 18626 24845 18660 24879
rect 18696 24845 18730 24879
rect 18766 24845 18800 24879
rect 18836 24845 18870 24879
rect 18906 24845 18940 24879
rect 18976 24845 19010 24879
rect 18025 24766 18059 24800
rect 18101 24766 18135 24800
rect 18177 24766 18211 24800
rect 18253 24766 18287 24800
rect 18329 24766 18363 24800
rect 18405 24766 18439 24800
rect 18486 24776 18520 24810
rect 18556 24776 18590 24810
rect 18626 24776 18660 24810
rect 18696 24776 18730 24810
rect 18766 24776 18800 24810
rect 18836 24776 18870 24810
rect 18906 24776 18940 24810
rect 18976 24776 19010 24810
rect 18025 24697 18059 24731
rect 18101 24697 18135 24731
rect 18177 24697 18211 24731
rect 18253 24697 18287 24731
rect 18329 24697 18363 24731
rect 18405 24697 18439 24731
rect 18486 24707 18520 24741
rect 18556 24707 18590 24741
rect 18626 24707 18660 24741
rect 18696 24707 18730 24741
rect 18766 24707 18800 24741
rect 18836 24707 18870 24741
rect 18906 24707 18940 24741
rect 18976 24707 19010 24741
rect 18025 24628 18059 24662
rect 18101 24628 18135 24662
rect 18177 24628 18211 24662
rect 18253 24628 18287 24662
rect 18329 24628 18363 24662
rect 18405 24628 18439 24662
rect 18486 24638 18520 24672
rect 18556 24638 18590 24672
rect 18626 24638 18660 24672
rect 18696 24638 18730 24672
rect 18766 24638 18800 24672
rect 18836 24638 18870 24672
rect 18906 24638 18940 24672
rect 18976 24638 19010 24672
rect 18025 24559 18059 24593
rect 18101 24559 18135 24593
rect 18177 24559 18211 24593
rect 18253 24559 18287 24593
rect 18329 24559 18363 24593
rect 18405 24559 18439 24593
rect 18486 24569 18520 24603
rect 18556 24569 18590 24603
rect 18626 24569 18660 24603
rect 18696 24569 18730 24603
rect 18766 24569 18800 24603
rect 18836 24569 18870 24603
rect 18906 24569 18940 24603
rect 18976 24569 19010 24603
rect 18025 24490 18059 24524
rect 18101 24490 18135 24524
rect 18177 24490 18211 24524
rect 18253 24490 18287 24524
rect 18329 24490 18363 24524
rect 18405 24490 18439 24524
rect 18486 24500 18520 24534
rect 18556 24500 18590 24534
rect 18626 24500 18660 24534
rect 18696 24500 18730 24534
rect 18766 24500 18800 24534
rect 18836 24500 18870 24534
rect 18906 24500 18940 24534
rect 18976 24500 19010 24534
rect 18025 24421 18059 24455
rect 18101 24421 18135 24455
rect 18177 24421 18211 24455
rect 18253 24421 18287 24455
rect 18329 24421 18363 24455
rect 18405 24421 18439 24455
rect 18486 24431 18520 24465
rect 18556 24431 18590 24465
rect 18626 24431 18660 24465
rect 18696 24431 18730 24465
rect 18766 24431 18800 24465
rect 18836 24431 18870 24465
rect 18906 24431 18940 24465
rect 18976 24431 19010 24465
rect 18025 24352 18059 24386
rect 18101 24352 18135 24386
rect 18177 24352 18211 24386
rect 18253 24352 18287 24386
rect 18329 24352 18363 24386
rect 18405 24352 18439 24386
rect 18486 24362 18520 24396
rect 18556 24362 18590 24396
rect 18626 24362 18660 24396
rect 18696 24362 18730 24396
rect 18766 24362 18800 24396
rect 18836 24362 18870 24396
rect 18906 24362 18940 24396
rect 18976 24362 19010 24396
rect 18025 24283 18059 24317
rect 18101 24283 18135 24317
rect 18177 24283 18211 24317
rect 18253 24283 18287 24317
rect 18329 24283 18363 24317
rect 18405 24283 18439 24317
rect 18486 24293 18520 24327
rect 18556 24293 18590 24327
rect 18626 24293 18660 24327
rect 18696 24293 18730 24327
rect 18766 24293 18800 24327
rect 18836 24293 18870 24327
rect 18906 24293 18940 24327
rect 18976 24293 19010 24327
rect 18025 24214 18059 24248
rect 18101 24214 18135 24248
rect 18177 24214 18211 24248
rect 18253 24214 18287 24248
rect 18329 24214 18363 24248
rect 18405 24214 18439 24248
rect 18486 24224 18520 24258
rect 18556 24224 18590 24258
rect 18626 24224 18660 24258
rect 18696 24224 18730 24258
rect 18766 24224 18800 24258
rect 18836 24224 18870 24258
rect 18906 24224 18940 24258
rect 18976 24224 19010 24258
rect 18025 24145 18059 24179
rect 18101 24145 18135 24179
rect 18177 24145 18211 24179
rect 18253 24145 18287 24179
rect 18329 24145 18363 24179
rect 18405 24145 18439 24179
rect 18486 24155 18520 24189
rect 18556 24155 18590 24189
rect 18626 24155 18660 24189
rect 18696 24155 18730 24189
rect 18766 24155 18800 24189
rect 18836 24155 18870 24189
rect 18906 24155 18940 24189
rect 18976 24155 19010 24189
rect 18025 24076 18059 24110
rect 18101 24076 18135 24110
rect 18177 24076 18211 24110
rect 18253 24076 18287 24110
rect 18329 24076 18363 24110
rect 18405 24076 18439 24110
rect 18486 24086 18520 24120
rect 18556 24086 18590 24120
rect 18626 24086 18660 24120
rect 18696 24086 18730 24120
rect 18766 24086 18800 24120
rect 18836 24086 18870 24120
rect 18906 24086 18940 24120
rect 18976 24086 19010 24120
rect 18025 24007 18059 24041
rect 18101 24007 18135 24041
rect 18177 24007 18211 24041
rect 18253 24007 18287 24041
rect 18329 24007 18363 24041
rect 18405 24007 18439 24041
rect 18486 24017 18520 24051
rect 18556 24017 18590 24051
rect 18626 24017 18660 24051
rect 18696 24017 18730 24051
rect 18766 24017 18800 24051
rect 18836 24017 18870 24051
rect 18906 24017 18940 24051
rect 18976 24017 19010 24051
rect 18025 23938 18059 23972
rect 18101 23938 18135 23972
rect 18177 23938 18211 23972
rect 18253 23938 18287 23972
rect 18329 23938 18363 23972
rect 18405 23938 18439 23972
rect 18486 23948 18520 23982
rect 18556 23948 18590 23982
rect 18626 23948 18660 23982
rect 18696 23948 18730 23982
rect 18766 23948 18800 23982
rect 18836 23948 18870 23982
rect 18906 23948 18940 23982
rect 18976 23948 19010 23982
rect 18025 23869 18059 23903
rect 18101 23869 18135 23903
rect 18177 23869 18211 23903
rect 18253 23869 18287 23903
rect 18329 23869 18363 23903
rect 18405 23869 18439 23903
rect 18486 23879 18520 23913
rect 18556 23879 18590 23913
rect 18626 23879 18660 23913
rect 18696 23879 18730 23913
rect 18766 23879 18800 23913
rect 18836 23879 18870 23913
rect 18906 23879 18940 23913
rect 18976 23879 19010 23913
rect 314 23719 348 23753
rect 384 23719 418 23753
rect 454 23719 488 23753
rect 524 23719 558 23753
rect 594 23719 628 23753
rect 664 23719 698 23753
rect 734 23719 768 23753
rect 804 23719 838 23753
rect 874 23719 908 23753
rect 944 23719 978 23753
rect 1014 23719 1048 23753
rect 1084 23719 1118 23753
rect 1154 23719 1188 23753
rect 1224 23719 1258 23753
rect 1294 23719 1328 23753
rect 1364 23719 1398 23753
rect 1434 23719 1468 23753
rect 1545 23719 1579 23753
rect 1613 23719 1647 23753
rect 1681 23719 1715 23753
rect 314 23649 348 23683
rect 384 23649 418 23683
rect 454 23649 488 23683
rect 524 23649 558 23683
rect 594 23649 628 23683
rect 664 23649 698 23683
rect 734 23649 768 23683
rect 804 23649 838 23683
rect 874 23649 908 23683
rect 944 23649 978 23683
rect 1014 23649 1048 23683
rect 1084 23649 1118 23683
rect 1154 23649 1188 23683
rect 1224 23649 1258 23683
rect 1294 23649 1328 23683
rect 1364 23649 1398 23683
rect 1434 23649 1468 23683
rect 1545 23616 1579 23650
rect 1613 23616 1647 23650
rect 1681 23616 1715 23650
rect 314 23579 348 23613
rect 384 23579 418 23613
rect 454 23579 488 23613
rect 524 23579 558 23613
rect 594 23579 628 23613
rect 664 23579 698 23613
rect 734 23579 768 23613
rect 804 23579 838 23613
rect 874 23579 908 23613
rect 944 23579 978 23613
rect 1014 23579 1048 23613
rect 1084 23579 1118 23613
rect 1154 23579 1188 23613
rect 1224 23579 1258 23613
rect 1294 23579 1328 23613
rect 1364 23579 1398 23613
rect 1434 23579 1468 23613
rect 18025 23800 18059 23834
rect 18101 23800 18135 23834
rect 18177 23800 18211 23834
rect 18253 23800 18287 23834
rect 18329 23800 18363 23834
rect 18405 23800 18439 23834
rect 18486 23810 18520 23844
rect 18556 23810 18590 23844
rect 18626 23810 18660 23844
rect 18696 23810 18730 23844
rect 18766 23810 18800 23844
rect 18836 23810 18870 23844
rect 18906 23810 18940 23844
rect 18976 23810 19010 23844
rect 18025 23731 18059 23765
rect 18101 23731 18135 23765
rect 18177 23731 18211 23765
rect 18253 23731 18287 23765
rect 18329 23731 18363 23765
rect 18405 23731 18439 23765
rect 18486 23741 18520 23775
rect 18556 23741 18590 23775
rect 18626 23741 18660 23775
rect 18696 23741 18730 23775
rect 18766 23741 18800 23775
rect 18836 23741 18870 23775
rect 18906 23741 18940 23775
rect 18976 23741 19010 23775
rect 18025 23662 18059 23696
rect 18101 23662 18135 23696
rect 18177 23662 18211 23696
rect 18253 23662 18287 23696
rect 18329 23662 18363 23696
rect 18405 23662 18439 23696
rect 18486 23672 18520 23706
rect 18556 23672 18590 23706
rect 18626 23672 18660 23706
rect 18696 23672 18730 23706
rect 18766 23672 18800 23706
rect 18836 23672 18870 23706
rect 18906 23672 18940 23706
rect 18976 23672 19010 23706
rect 18025 23593 18059 23627
rect 18101 23593 18135 23627
rect 18177 23593 18211 23627
rect 18253 23593 18287 23627
rect 18329 23593 18363 23627
rect 18405 23593 18439 23627
rect 18486 23603 18520 23637
rect 18556 23603 18590 23637
rect 18626 23603 18660 23637
rect 18696 23603 18730 23637
rect 18766 23603 18800 23637
rect 18836 23603 18870 23637
rect 18906 23603 18940 23637
rect 18976 23603 19010 23637
rect 314 23509 348 23543
rect 384 23509 418 23543
rect 454 23509 488 23543
rect 524 23509 558 23543
rect 594 23509 628 23543
rect 664 23509 698 23543
rect 734 23509 768 23543
rect 804 23509 838 23543
rect 874 23509 908 23543
rect 944 23509 978 23543
rect 1014 23509 1048 23543
rect 1084 23509 1118 23543
rect 1154 23509 1188 23543
rect 1224 23509 1258 23543
rect 1294 23509 1328 23543
rect 1364 23509 1398 23543
rect 1434 23509 1468 23543
rect 18025 23524 18059 23558
rect 18101 23524 18135 23558
rect 18177 23524 18211 23558
rect 18253 23524 18287 23558
rect 18329 23524 18363 23558
rect 18405 23524 18439 23558
rect 18486 23534 18520 23568
rect 18556 23534 18590 23568
rect 18626 23534 18660 23568
rect 18696 23534 18730 23568
rect 18766 23534 18800 23568
rect 18836 23534 18870 23568
rect 18906 23534 18940 23568
rect 18976 23534 19010 23568
rect 22827 30683 22861 30717
rect 22897 30683 22931 30717
rect 22967 30683 23001 30717
rect 23037 30683 23071 30717
rect 23107 30683 23141 30717
rect 23177 30683 23211 30717
rect 23247 30683 23281 30717
rect 23317 30683 23351 30717
rect 23387 30683 23421 30717
rect 23457 30683 23491 30717
rect 23527 30683 23561 30717
rect 23597 30683 23631 30717
rect 22827 30615 22861 30649
rect 22897 30615 22931 30649
rect 22967 30615 23001 30649
rect 23037 30615 23071 30649
rect 23107 30615 23141 30649
rect 23177 30615 23211 30649
rect 23247 30615 23281 30649
rect 23317 30615 23351 30649
rect 23387 30615 23421 30649
rect 23457 30615 23491 30649
rect 23527 30615 23561 30649
rect 23597 30615 23631 30649
rect 22827 30547 22861 30581
rect 22897 30547 22931 30581
rect 22967 30547 23001 30581
rect 23037 30547 23071 30581
rect 23107 30547 23141 30581
rect 23177 30547 23211 30581
rect 23247 30547 23281 30581
rect 23317 30547 23351 30581
rect 23387 30547 23421 30581
rect 23457 30547 23491 30581
rect 23527 30547 23561 30581
rect 23597 30547 23631 30581
rect 22827 30479 22861 30513
rect 22897 30479 22931 30513
rect 22967 30479 23001 30513
rect 23037 30479 23071 30513
rect 23107 30479 23141 30513
rect 23177 30479 23211 30513
rect 23247 30479 23281 30513
rect 23317 30479 23351 30513
rect 23387 30479 23421 30513
rect 23457 30479 23491 30513
rect 23527 30479 23561 30513
rect 23597 30479 23631 30513
rect 22827 30411 22861 30445
rect 22897 30411 22931 30445
rect 22967 30411 23001 30445
rect 23037 30411 23071 30445
rect 23107 30411 23141 30445
rect 23177 30411 23211 30445
rect 23247 30411 23281 30445
rect 23317 30411 23351 30445
rect 23387 30411 23421 30445
rect 23457 30411 23491 30445
rect 23527 30411 23561 30445
rect 23597 30411 23631 30445
rect 22827 30343 22861 30377
rect 22897 30343 22931 30377
rect 22967 30343 23001 30377
rect 23037 30343 23071 30377
rect 23107 30343 23141 30377
rect 23177 30343 23211 30377
rect 23247 30343 23281 30377
rect 23317 30343 23351 30377
rect 23387 30343 23421 30377
rect 23457 30343 23491 30377
rect 23527 30343 23561 30377
rect 23597 30343 23631 30377
rect 22827 30275 22861 30309
rect 22897 30275 22931 30309
rect 22967 30275 23001 30309
rect 23037 30275 23071 30309
rect 23107 30275 23141 30309
rect 23177 30275 23211 30309
rect 23247 30275 23281 30309
rect 23317 30275 23351 30309
rect 23387 30275 23421 30309
rect 23457 30275 23491 30309
rect 23527 30275 23561 30309
rect 23597 30275 23631 30309
rect 22827 30207 22861 30241
rect 22897 30207 22931 30241
rect 22967 30207 23001 30241
rect 23037 30207 23071 30241
rect 23107 30207 23141 30241
rect 23177 30207 23211 30241
rect 23247 30207 23281 30241
rect 23317 30207 23351 30241
rect 23387 30207 23421 30241
rect 23457 30207 23491 30241
rect 23527 30207 23561 30241
rect 23597 30207 23631 30241
rect 22827 30139 22861 30173
rect 22897 30139 22931 30173
rect 22967 30139 23001 30173
rect 23037 30139 23071 30173
rect 23107 30139 23141 30173
rect 23177 30139 23211 30173
rect 23247 30139 23281 30173
rect 23317 30139 23351 30173
rect 23387 30139 23421 30173
rect 23457 30139 23491 30173
rect 23527 30139 23561 30173
rect 23597 30139 23631 30173
rect 22827 30071 22861 30105
rect 22897 30071 22931 30105
rect 22967 30071 23001 30105
rect 23037 30071 23071 30105
rect 23107 30071 23141 30105
rect 23177 30071 23211 30105
rect 23247 30071 23281 30105
rect 23317 30071 23351 30105
rect 23387 30071 23421 30105
rect 23457 30071 23491 30105
rect 23527 30071 23561 30105
rect 23597 30071 23631 30105
rect 22827 30003 22861 30037
rect 22897 30003 22931 30037
rect 22967 30003 23001 30037
rect 23037 30003 23071 30037
rect 23107 30003 23141 30037
rect 23177 30003 23211 30037
rect 23247 30003 23281 30037
rect 23317 30003 23351 30037
rect 23387 30003 23421 30037
rect 23457 30003 23491 30037
rect 23527 30003 23561 30037
rect 23597 30003 23631 30037
rect 22827 29935 22861 29969
rect 22897 29935 22931 29969
rect 22967 29935 23001 29969
rect 23037 29935 23071 29969
rect 23107 29935 23141 29969
rect 23177 29935 23211 29969
rect 23247 29935 23281 29969
rect 23317 29935 23351 29969
rect 23387 29935 23421 29969
rect 23457 29935 23491 29969
rect 23527 29935 23561 29969
rect 23597 29935 23631 29969
rect 22827 29867 22861 29901
rect 22897 29867 22931 29901
rect 22967 29867 23001 29901
rect 23037 29867 23071 29901
rect 23107 29867 23141 29901
rect 23177 29867 23211 29901
rect 23247 29867 23281 29901
rect 23317 29867 23351 29901
rect 23387 29867 23421 29901
rect 23457 29867 23491 29901
rect 23527 29867 23561 29901
rect 23597 29867 23631 29901
rect 22827 29799 22861 29833
rect 22897 29799 22931 29833
rect 22967 29799 23001 29833
rect 23037 29799 23071 29833
rect 23107 29799 23141 29833
rect 23177 29799 23211 29833
rect 23247 29799 23281 29833
rect 23317 29799 23351 29833
rect 23387 29799 23421 29833
rect 23457 29799 23491 29833
rect 23527 29799 23561 29833
rect 23597 29799 23631 29833
rect 22827 29731 22861 29765
rect 22897 29731 22931 29765
rect 22967 29731 23001 29765
rect 23037 29731 23071 29765
rect 23107 29731 23141 29765
rect 23177 29731 23211 29765
rect 23247 29731 23281 29765
rect 23317 29731 23351 29765
rect 23387 29731 23421 29765
rect 23457 29731 23491 29765
rect 23527 29731 23561 29765
rect 23597 29731 23631 29765
rect 22827 29663 22861 29697
rect 22897 29663 22931 29697
rect 22967 29663 23001 29697
rect 23037 29663 23071 29697
rect 23107 29663 23141 29697
rect 23177 29663 23211 29697
rect 23247 29663 23281 29697
rect 23317 29663 23351 29697
rect 23387 29663 23421 29697
rect 23457 29663 23491 29697
rect 23527 29663 23561 29697
rect 23597 29663 23631 29697
rect 22827 29595 22861 29629
rect 22897 29595 22931 29629
rect 22967 29595 23001 29629
rect 23037 29595 23071 29629
rect 23107 29595 23141 29629
rect 23177 29595 23211 29629
rect 23247 29595 23281 29629
rect 23317 29595 23351 29629
rect 23387 29595 23421 29629
rect 23457 29595 23491 29629
rect 23527 29595 23561 29629
rect 23597 29595 23631 29629
rect 22827 29527 22861 29561
rect 22897 29527 22931 29561
rect 22967 29527 23001 29561
rect 23037 29527 23071 29561
rect 23107 29527 23141 29561
rect 23177 29527 23211 29561
rect 23247 29527 23281 29561
rect 23317 29527 23351 29561
rect 23387 29527 23421 29561
rect 23457 29527 23491 29561
rect 23527 29527 23561 29561
rect 23597 29527 23631 29561
rect 22827 29459 22861 29493
rect 22897 29459 22931 29493
rect 22967 29459 23001 29493
rect 23037 29459 23071 29493
rect 23107 29459 23141 29493
rect 23177 29459 23211 29493
rect 23247 29459 23281 29493
rect 23317 29459 23351 29493
rect 23387 29459 23421 29493
rect 23457 29459 23491 29493
rect 23527 29459 23561 29493
rect 23597 29459 23631 29493
rect 22827 29391 22861 29425
rect 22897 29391 22931 29425
rect 22967 29391 23001 29425
rect 23037 29391 23071 29425
rect 23107 29391 23141 29425
rect 23177 29391 23211 29425
rect 23247 29391 23281 29425
rect 23317 29391 23351 29425
rect 23387 29391 23421 29425
rect 23457 29391 23491 29425
rect 23527 29391 23561 29425
rect 23597 29391 23631 29425
rect 22827 29323 22861 29357
rect 22897 29323 22931 29357
rect 22967 29323 23001 29357
rect 23037 29323 23071 29357
rect 23107 29323 23141 29357
rect 23177 29323 23211 29357
rect 23247 29323 23281 29357
rect 23317 29323 23351 29357
rect 23387 29323 23421 29357
rect 23457 29323 23491 29357
rect 23527 29323 23561 29357
rect 23597 29323 23631 29357
rect 22827 29255 22861 29289
rect 22897 29255 22931 29289
rect 22967 29255 23001 29289
rect 23037 29255 23071 29289
rect 23107 29255 23141 29289
rect 23177 29255 23211 29289
rect 23247 29255 23281 29289
rect 23317 29255 23351 29289
rect 23387 29255 23421 29289
rect 23457 29255 23491 29289
rect 23527 29255 23561 29289
rect 23597 29255 23631 29289
rect 22827 29187 22861 29221
rect 22897 29187 22931 29221
rect 22967 29187 23001 29221
rect 23037 29187 23071 29221
rect 23107 29187 23141 29221
rect 23177 29187 23211 29221
rect 23247 29187 23281 29221
rect 23317 29187 23351 29221
rect 23387 29187 23421 29221
rect 23457 29187 23491 29221
rect 23527 29187 23561 29221
rect 23597 29187 23631 29221
rect 22827 29119 22861 29153
rect 22897 29119 22931 29153
rect 22967 29119 23001 29153
rect 23037 29119 23071 29153
rect 23107 29119 23141 29153
rect 23177 29119 23211 29153
rect 23247 29119 23281 29153
rect 23317 29119 23351 29153
rect 23387 29119 23421 29153
rect 23457 29119 23491 29153
rect 23527 29119 23561 29153
rect 23597 29119 23631 29153
rect 22827 29051 22861 29085
rect 22897 29051 22931 29085
rect 22967 29051 23001 29085
rect 23037 29051 23071 29085
rect 23107 29051 23141 29085
rect 23177 29051 23211 29085
rect 23247 29051 23281 29085
rect 23317 29051 23351 29085
rect 23387 29051 23421 29085
rect 23457 29051 23491 29085
rect 23527 29051 23561 29085
rect 23597 29051 23631 29085
rect 22827 28983 22861 29017
rect 22897 28983 22931 29017
rect 22967 28983 23001 29017
rect 23037 28983 23071 29017
rect 23107 28983 23141 29017
rect 23177 28983 23211 29017
rect 23247 28983 23281 29017
rect 23317 28983 23351 29017
rect 23387 28983 23421 29017
rect 23457 28983 23491 29017
rect 23527 28983 23561 29017
rect 23597 28983 23631 29017
rect 22827 28915 22861 28949
rect 22897 28915 22931 28949
rect 22967 28915 23001 28949
rect 23037 28915 23071 28949
rect 23107 28915 23141 28949
rect 23177 28915 23211 28949
rect 23247 28915 23281 28949
rect 23317 28915 23351 28949
rect 23387 28915 23421 28949
rect 23457 28915 23491 28949
rect 23527 28915 23561 28949
rect 23597 28915 23631 28949
rect 22827 28847 22861 28881
rect 22897 28847 22931 28881
rect 22967 28847 23001 28881
rect 23037 28847 23071 28881
rect 23107 28847 23141 28881
rect 23177 28847 23211 28881
rect 23247 28847 23281 28881
rect 23317 28847 23351 28881
rect 23387 28847 23421 28881
rect 23457 28847 23491 28881
rect 23527 28847 23561 28881
rect 23597 28847 23631 28881
rect 22827 28779 22861 28813
rect 22897 28779 22931 28813
rect 22967 28779 23001 28813
rect 23037 28779 23071 28813
rect 23107 28779 23141 28813
rect 23177 28779 23211 28813
rect 23247 28779 23281 28813
rect 23317 28779 23351 28813
rect 23387 28779 23421 28813
rect 23457 28779 23491 28813
rect 23527 28779 23561 28813
rect 23597 28779 23631 28813
rect 22827 28711 22861 28745
rect 22897 28711 22931 28745
rect 22967 28711 23001 28745
rect 23037 28711 23071 28745
rect 23107 28711 23141 28745
rect 23177 28711 23211 28745
rect 23247 28711 23281 28745
rect 23317 28711 23351 28745
rect 23387 28711 23421 28745
rect 23457 28711 23491 28745
rect 23527 28711 23561 28745
rect 23597 28711 23631 28745
rect 22827 28643 22861 28677
rect 22897 28643 22931 28677
rect 22967 28643 23001 28677
rect 23037 28643 23071 28677
rect 23107 28643 23141 28677
rect 23177 28643 23211 28677
rect 23247 28643 23281 28677
rect 23317 28643 23351 28677
rect 23387 28643 23421 28677
rect 23457 28643 23491 28677
rect 23527 28643 23561 28677
rect 23597 28643 23631 28677
rect 22827 28575 22861 28609
rect 22897 28575 22931 28609
rect 22967 28575 23001 28609
rect 23037 28575 23071 28609
rect 23107 28575 23141 28609
rect 23177 28575 23211 28609
rect 23247 28575 23281 28609
rect 23317 28575 23351 28609
rect 23387 28575 23421 28609
rect 23457 28575 23491 28609
rect 23527 28575 23561 28609
rect 23597 28575 23631 28609
rect 22827 28507 22861 28541
rect 22897 28507 22931 28541
rect 22967 28507 23001 28541
rect 23037 28507 23071 28541
rect 23107 28507 23141 28541
rect 23177 28507 23211 28541
rect 23247 28507 23281 28541
rect 23317 28507 23351 28541
rect 23387 28507 23421 28541
rect 23457 28507 23491 28541
rect 23527 28507 23561 28541
rect 23597 28507 23631 28541
rect 22827 28439 22861 28473
rect 22897 28439 22931 28473
rect 22967 28439 23001 28473
rect 23037 28439 23071 28473
rect 23107 28439 23141 28473
rect 23177 28439 23211 28473
rect 23247 28439 23281 28473
rect 23317 28439 23351 28473
rect 23387 28439 23421 28473
rect 23457 28439 23491 28473
rect 23527 28439 23561 28473
rect 23597 28439 23631 28473
rect 22827 28371 22861 28405
rect 22897 28371 22931 28405
rect 22967 28371 23001 28405
rect 23037 28371 23071 28405
rect 23107 28371 23141 28405
rect 23177 28371 23211 28405
rect 23247 28371 23281 28405
rect 23317 28371 23351 28405
rect 23387 28371 23421 28405
rect 23457 28371 23491 28405
rect 23527 28371 23561 28405
rect 23597 28371 23631 28405
rect 22827 28303 22861 28337
rect 22897 28303 22931 28337
rect 22967 28303 23001 28337
rect 23037 28303 23071 28337
rect 23107 28303 23141 28337
rect 23177 28303 23211 28337
rect 23247 28303 23281 28337
rect 23317 28303 23351 28337
rect 23387 28303 23421 28337
rect 23457 28303 23491 28337
rect 23527 28303 23561 28337
rect 23597 28303 23631 28337
rect 22827 28235 22861 28269
rect 22897 28235 22931 28269
rect 22967 28235 23001 28269
rect 23037 28235 23071 28269
rect 23107 28235 23141 28269
rect 23177 28235 23211 28269
rect 23247 28235 23281 28269
rect 23317 28235 23351 28269
rect 23387 28235 23421 28269
rect 23457 28235 23491 28269
rect 23527 28235 23561 28269
rect 23597 28235 23631 28269
rect 22827 28167 22861 28201
rect 22897 28167 22931 28201
rect 22967 28167 23001 28201
rect 23037 28167 23071 28201
rect 23107 28167 23141 28201
rect 23177 28167 23211 28201
rect 23247 28167 23281 28201
rect 23317 28167 23351 28201
rect 23387 28167 23421 28201
rect 23457 28167 23491 28201
rect 23527 28167 23561 28201
rect 23597 28167 23631 28201
rect 22827 28099 22861 28133
rect 22897 28099 22931 28133
rect 22967 28099 23001 28133
rect 23037 28099 23071 28133
rect 23107 28099 23141 28133
rect 23177 28099 23211 28133
rect 23247 28099 23281 28133
rect 23317 28099 23351 28133
rect 23387 28099 23421 28133
rect 23457 28099 23491 28133
rect 23527 28099 23561 28133
rect 23597 28099 23631 28133
rect 22827 28031 22861 28065
rect 22897 28031 22931 28065
rect 22967 28031 23001 28065
rect 23037 28031 23071 28065
rect 23107 28031 23141 28065
rect 23177 28031 23211 28065
rect 23247 28031 23281 28065
rect 23317 28031 23351 28065
rect 23387 28031 23421 28065
rect 23457 28031 23491 28065
rect 23527 28031 23561 28065
rect 23597 28031 23631 28065
rect 22827 27963 22861 27997
rect 22897 27963 22931 27997
rect 22967 27963 23001 27997
rect 23037 27963 23071 27997
rect 23107 27963 23141 27997
rect 23177 27963 23211 27997
rect 23247 27963 23281 27997
rect 23317 27963 23351 27997
rect 23387 27963 23421 27997
rect 23457 27963 23491 27997
rect 23527 27963 23561 27997
rect 23597 27963 23631 27997
rect 22827 27895 22861 27929
rect 22897 27895 22931 27929
rect 22967 27895 23001 27929
rect 23037 27895 23071 27929
rect 23107 27895 23141 27929
rect 23177 27895 23211 27929
rect 23247 27895 23281 27929
rect 23317 27895 23351 27929
rect 23387 27895 23421 27929
rect 23457 27895 23491 27929
rect 23527 27895 23561 27929
rect 23597 27895 23631 27929
rect 22827 27827 22861 27861
rect 22897 27827 22931 27861
rect 22967 27827 23001 27861
rect 23037 27827 23071 27861
rect 23107 27827 23141 27861
rect 23177 27827 23211 27861
rect 23247 27827 23281 27861
rect 23317 27827 23351 27861
rect 23387 27827 23421 27861
rect 23457 27827 23491 27861
rect 23527 27827 23561 27861
rect 23597 27827 23631 27861
rect 22827 27759 22861 27793
rect 22897 27759 22931 27793
rect 22967 27759 23001 27793
rect 23037 27759 23071 27793
rect 23107 27759 23141 27793
rect 23177 27759 23211 27793
rect 23247 27759 23281 27793
rect 23317 27759 23351 27793
rect 23387 27759 23421 27793
rect 23457 27759 23491 27793
rect 23527 27759 23561 27793
rect 23597 27759 23631 27793
rect 22827 27691 22861 27725
rect 22897 27691 22931 27725
rect 22967 27691 23001 27725
rect 23037 27691 23071 27725
rect 23107 27691 23141 27725
rect 23177 27691 23211 27725
rect 23247 27691 23281 27725
rect 23317 27691 23351 27725
rect 23387 27691 23421 27725
rect 23457 27691 23491 27725
rect 23527 27691 23561 27725
rect 23597 27691 23631 27725
rect 22827 27623 22861 27657
rect 22897 27623 22931 27657
rect 22967 27623 23001 27657
rect 23037 27623 23071 27657
rect 23107 27623 23141 27657
rect 23177 27623 23211 27657
rect 23247 27623 23281 27657
rect 23317 27623 23351 27657
rect 23387 27623 23421 27657
rect 23457 27623 23491 27657
rect 23527 27623 23561 27657
rect 23597 27623 23631 27657
rect 22827 27555 22861 27589
rect 22897 27555 22931 27589
rect 22967 27555 23001 27589
rect 23037 27555 23071 27589
rect 23107 27555 23141 27589
rect 23177 27555 23211 27589
rect 23247 27555 23281 27589
rect 23317 27555 23351 27589
rect 23387 27555 23421 27589
rect 23457 27555 23491 27589
rect 23527 27555 23561 27589
rect 23597 27555 23631 27589
rect 22827 27487 22861 27521
rect 22897 27487 22931 27521
rect 22967 27487 23001 27521
rect 23037 27487 23071 27521
rect 23107 27487 23141 27521
rect 23177 27487 23211 27521
rect 23247 27487 23281 27521
rect 23317 27487 23351 27521
rect 23387 27487 23421 27521
rect 23457 27487 23491 27521
rect 23527 27487 23561 27521
rect 23597 27487 23631 27521
rect 22827 27419 22861 27453
rect 22897 27419 22931 27453
rect 22967 27419 23001 27453
rect 23037 27419 23071 27453
rect 23107 27419 23141 27453
rect 23177 27419 23211 27453
rect 23247 27419 23281 27453
rect 23317 27419 23351 27453
rect 23387 27419 23421 27453
rect 23457 27419 23491 27453
rect 23527 27419 23561 27453
rect 23597 27419 23631 27453
rect 22827 27351 22861 27385
rect 22897 27351 22931 27385
rect 22967 27351 23001 27385
rect 23037 27351 23071 27385
rect 23107 27351 23141 27385
rect 23177 27351 23211 27385
rect 23247 27351 23281 27385
rect 23317 27351 23351 27385
rect 23387 27351 23421 27385
rect 23457 27351 23491 27385
rect 23527 27351 23561 27385
rect 23597 27351 23631 27385
rect 22827 27283 22861 27317
rect 22897 27283 22931 27317
rect 22967 27283 23001 27317
rect 23037 27283 23071 27317
rect 23107 27283 23141 27317
rect 23177 27283 23211 27317
rect 23247 27283 23281 27317
rect 23317 27283 23351 27317
rect 23387 27283 23421 27317
rect 23457 27283 23491 27317
rect 23527 27283 23561 27317
rect 23597 27283 23631 27317
rect 22827 27215 22861 27249
rect 22897 27215 22931 27249
rect 22967 27215 23001 27249
rect 23037 27215 23071 27249
rect 23107 27215 23141 27249
rect 23177 27215 23211 27249
rect 23247 27215 23281 27249
rect 23317 27215 23351 27249
rect 23387 27215 23421 27249
rect 23457 27215 23491 27249
rect 23527 27215 23561 27249
rect 23597 27215 23631 27249
rect 22827 27147 22861 27181
rect 22897 27147 22931 27181
rect 22967 27147 23001 27181
rect 23037 27147 23071 27181
rect 23107 27147 23141 27181
rect 23177 27147 23211 27181
rect 23247 27147 23281 27181
rect 23317 27147 23351 27181
rect 23387 27147 23421 27181
rect 23457 27147 23491 27181
rect 23527 27147 23561 27181
rect 23597 27147 23631 27181
rect 22827 27079 22861 27113
rect 22897 27079 22931 27113
rect 22967 27079 23001 27113
rect 23037 27079 23071 27113
rect 23107 27079 23141 27113
rect 23177 27079 23211 27113
rect 23247 27079 23281 27113
rect 23317 27079 23351 27113
rect 23387 27079 23421 27113
rect 23457 27079 23491 27113
rect 23527 27079 23561 27113
rect 23597 27079 23631 27113
rect 22827 27011 22861 27045
rect 22897 27011 22931 27045
rect 22967 27011 23001 27045
rect 23037 27011 23071 27045
rect 23107 27011 23141 27045
rect 23177 27011 23211 27045
rect 23247 27011 23281 27045
rect 23317 27011 23351 27045
rect 23387 27011 23421 27045
rect 23457 27011 23491 27045
rect 23527 27011 23561 27045
rect 23597 27011 23631 27045
rect 22827 26943 22861 26977
rect 22897 26943 22931 26977
rect 22967 26943 23001 26977
rect 23037 26943 23071 26977
rect 23107 26943 23141 26977
rect 23177 26943 23211 26977
rect 23247 26943 23281 26977
rect 23317 26943 23351 26977
rect 23387 26943 23421 26977
rect 23457 26943 23491 26977
rect 23527 26943 23561 26977
rect 23597 26943 23631 26977
rect 22827 26875 22861 26909
rect 22897 26875 22931 26909
rect 22967 26875 23001 26909
rect 23037 26875 23071 26909
rect 23107 26875 23141 26909
rect 23177 26875 23211 26909
rect 23247 26875 23281 26909
rect 23317 26875 23351 26909
rect 23387 26875 23421 26909
rect 23457 26875 23491 26909
rect 23527 26875 23561 26909
rect 23597 26875 23631 26909
rect 22827 26807 22861 26841
rect 22897 26807 22931 26841
rect 22967 26807 23001 26841
rect 23037 26807 23071 26841
rect 23107 26807 23141 26841
rect 23177 26807 23211 26841
rect 23247 26807 23281 26841
rect 23317 26807 23351 26841
rect 23387 26807 23421 26841
rect 23457 26807 23491 26841
rect 23527 26807 23561 26841
rect 23597 26807 23631 26841
rect 22827 26739 22861 26773
rect 22897 26739 22931 26773
rect 22967 26739 23001 26773
rect 23037 26739 23071 26773
rect 23107 26739 23141 26773
rect 23177 26739 23211 26773
rect 23247 26739 23281 26773
rect 23317 26739 23351 26773
rect 23387 26739 23421 26773
rect 23457 26739 23491 26773
rect 23527 26739 23561 26773
rect 23597 26739 23631 26773
rect 22827 26671 22861 26705
rect 22897 26671 22931 26705
rect 22967 26671 23001 26705
rect 23037 26671 23071 26705
rect 23107 26671 23141 26705
rect 23177 26671 23211 26705
rect 23247 26671 23281 26705
rect 23317 26671 23351 26705
rect 23387 26671 23421 26705
rect 23457 26671 23491 26705
rect 23527 26671 23561 26705
rect 23597 26671 23631 26705
rect 22827 26603 22861 26637
rect 22897 26603 22931 26637
rect 22967 26603 23001 26637
rect 23037 26603 23071 26637
rect 23107 26603 23141 26637
rect 23177 26603 23211 26637
rect 23247 26603 23281 26637
rect 23317 26603 23351 26637
rect 23387 26603 23421 26637
rect 23457 26603 23491 26637
rect 23527 26603 23561 26637
rect 23597 26603 23631 26637
rect 22827 26535 22861 26569
rect 22897 26535 22931 26569
rect 22967 26535 23001 26569
rect 23037 26535 23071 26569
rect 23107 26535 23141 26569
rect 23177 26535 23211 26569
rect 23247 26535 23281 26569
rect 23317 26535 23351 26569
rect 23387 26535 23421 26569
rect 23457 26535 23491 26569
rect 23527 26535 23561 26569
rect 23597 26535 23631 26569
rect 22827 26467 22861 26501
rect 22897 26467 22931 26501
rect 22967 26467 23001 26501
rect 23037 26467 23071 26501
rect 23107 26467 23141 26501
rect 23177 26467 23211 26501
rect 23247 26467 23281 26501
rect 23317 26467 23351 26501
rect 23387 26467 23421 26501
rect 23457 26467 23491 26501
rect 23527 26467 23561 26501
rect 23597 26467 23631 26501
rect 22827 26399 22861 26433
rect 22897 26399 22931 26433
rect 22967 26399 23001 26433
rect 23037 26399 23071 26433
rect 23107 26399 23141 26433
rect 23177 26399 23211 26433
rect 23247 26399 23281 26433
rect 23317 26399 23351 26433
rect 23387 26399 23421 26433
rect 23457 26399 23491 26433
rect 23527 26399 23561 26433
rect 23597 26399 23631 26433
rect 22827 26331 22861 26365
rect 22897 26331 22931 26365
rect 22967 26331 23001 26365
rect 23037 26331 23071 26365
rect 23107 26331 23141 26365
rect 23177 26331 23211 26365
rect 23247 26331 23281 26365
rect 23317 26331 23351 26365
rect 23387 26331 23421 26365
rect 23457 26331 23491 26365
rect 23527 26331 23561 26365
rect 23597 26331 23631 26365
rect 22827 26263 22861 26297
rect 22897 26263 22931 26297
rect 22967 26263 23001 26297
rect 23037 26263 23071 26297
rect 23107 26263 23141 26297
rect 23177 26263 23211 26297
rect 23247 26263 23281 26297
rect 23317 26263 23351 26297
rect 23387 26263 23421 26297
rect 23457 26263 23491 26297
rect 23527 26263 23561 26297
rect 23597 26263 23631 26297
rect 22827 26195 22861 26229
rect 22897 26195 22931 26229
rect 22967 26195 23001 26229
rect 23037 26195 23071 26229
rect 23107 26195 23141 26229
rect 23177 26195 23211 26229
rect 23247 26195 23281 26229
rect 23317 26195 23351 26229
rect 23387 26195 23421 26229
rect 23457 26195 23491 26229
rect 23527 26195 23561 26229
rect 23597 26195 23631 26229
rect 22827 26127 22861 26161
rect 22897 26127 22931 26161
rect 22967 26127 23001 26161
rect 23037 26127 23071 26161
rect 23107 26127 23141 26161
rect 23177 26127 23211 26161
rect 23247 26127 23281 26161
rect 23317 26127 23351 26161
rect 23387 26127 23421 26161
rect 23457 26127 23491 26161
rect 23527 26127 23561 26161
rect 23597 26127 23631 26161
rect 22827 26059 22861 26093
rect 22897 26059 22931 26093
rect 22967 26059 23001 26093
rect 23037 26059 23071 26093
rect 23107 26059 23141 26093
rect 23177 26059 23211 26093
rect 23247 26059 23281 26093
rect 23317 26059 23351 26093
rect 23387 26059 23421 26093
rect 23457 26059 23491 26093
rect 23527 26059 23561 26093
rect 23597 26059 23631 26093
rect 22827 25991 22861 26025
rect 22897 25991 22931 26025
rect 22967 25991 23001 26025
rect 23037 25991 23071 26025
rect 23107 25991 23141 26025
rect 23177 25991 23211 26025
rect 23247 25991 23281 26025
rect 23317 25991 23351 26025
rect 23387 25991 23421 26025
rect 23457 25991 23491 26025
rect 23527 25991 23561 26025
rect 23597 25991 23631 26025
rect 22827 25923 22861 25957
rect 22897 25923 22931 25957
rect 22967 25923 23001 25957
rect 23037 25923 23071 25957
rect 23107 25923 23141 25957
rect 23177 25923 23211 25957
rect 23247 25923 23281 25957
rect 23317 25923 23351 25957
rect 23387 25923 23421 25957
rect 23457 25923 23491 25957
rect 23527 25923 23561 25957
rect 23597 25923 23631 25957
rect 22827 25855 22861 25889
rect 22897 25855 22931 25889
rect 22967 25855 23001 25889
rect 23037 25855 23071 25889
rect 23107 25855 23141 25889
rect 23177 25855 23211 25889
rect 23247 25855 23281 25889
rect 23317 25855 23351 25889
rect 23387 25855 23421 25889
rect 23457 25855 23491 25889
rect 23527 25855 23561 25889
rect 23597 25855 23631 25889
rect 22827 25787 22861 25821
rect 22897 25787 22931 25821
rect 22967 25787 23001 25821
rect 23037 25787 23071 25821
rect 23107 25787 23141 25821
rect 23177 25787 23211 25821
rect 23247 25787 23281 25821
rect 23317 25787 23351 25821
rect 23387 25787 23421 25821
rect 23457 25787 23491 25821
rect 23527 25787 23561 25821
rect 23597 25787 23631 25821
rect 22827 25719 22861 25753
rect 22897 25719 22931 25753
rect 22967 25719 23001 25753
rect 23037 25719 23071 25753
rect 23107 25719 23141 25753
rect 23177 25719 23211 25753
rect 23247 25719 23281 25753
rect 23317 25719 23351 25753
rect 23387 25719 23421 25753
rect 23457 25719 23491 25753
rect 23527 25719 23561 25753
rect 23597 25719 23631 25753
rect 22827 25651 22861 25685
rect 22897 25651 22931 25685
rect 22967 25651 23001 25685
rect 23037 25651 23071 25685
rect 23107 25651 23141 25685
rect 23177 25651 23211 25685
rect 23247 25651 23281 25685
rect 23317 25651 23351 25685
rect 23387 25651 23421 25685
rect 23457 25651 23491 25685
rect 23527 25651 23561 25685
rect 23597 25651 23631 25685
rect 22827 25583 22861 25617
rect 22897 25583 22931 25617
rect 22967 25583 23001 25617
rect 23037 25583 23071 25617
rect 23107 25583 23141 25617
rect 23177 25583 23211 25617
rect 23247 25583 23281 25617
rect 23317 25583 23351 25617
rect 23387 25583 23421 25617
rect 23457 25583 23491 25617
rect 23527 25583 23561 25617
rect 23597 25583 23631 25617
rect 22827 25515 22861 25549
rect 22897 25515 22931 25549
rect 22967 25515 23001 25549
rect 23037 25515 23071 25549
rect 23107 25515 23141 25549
rect 23177 25515 23211 25549
rect 23247 25515 23281 25549
rect 23317 25515 23351 25549
rect 23387 25515 23421 25549
rect 23457 25515 23491 25549
rect 23527 25515 23561 25549
rect 23597 25515 23631 25549
rect 22827 25447 22861 25481
rect 22897 25447 22931 25481
rect 22967 25447 23001 25481
rect 23037 25447 23071 25481
rect 23107 25447 23141 25481
rect 23177 25447 23211 25481
rect 23247 25447 23281 25481
rect 23317 25447 23351 25481
rect 23387 25447 23421 25481
rect 23457 25447 23491 25481
rect 23527 25447 23561 25481
rect 23597 25447 23631 25481
rect 22827 25379 22861 25413
rect 22897 25379 22931 25413
rect 22967 25379 23001 25413
rect 23037 25379 23071 25413
rect 23107 25379 23141 25413
rect 23177 25379 23211 25413
rect 23247 25379 23281 25413
rect 23317 25379 23351 25413
rect 23387 25379 23421 25413
rect 23457 25379 23491 25413
rect 23527 25379 23561 25413
rect 23597 25379 23631 25413
rect 22827 25311 22861 25345
rect 22897 25311 22931 25345
rect 22967 25311 23001 25345
rect 23037 25311 23071 25345
rect 23107 25311 23141 25345
rect 23177 25311 23211 25345
rect 23247 25311 23281 25345
rect 23317 25311 23351 25345
rect 23387 25311 23421 25345
rect 23457 25311 23491 25345
rect 23527 25311 23561 25345
rect 23597 25311 23631 25345
rect 22827 25243 22861 25277
rect 22897 25243 22931 25277
rect 22967 25243 23001 25277
rect 23037 25243 23071 25277
rect 23107 25243 23141 25277
rect 23177 25243 23211 25277
rect 23247 25243 23281 25277
rect 23317 25243 23351 25277
rect 23387 25243 23421 25277
rect 23457 25243 23491 25277
rect 23527 25243 23561 25277
rect 23597 25243 23631 25277
rect 22827 25175 22861 25209
rect 22897 25175 22931 25209
rect 22967 25175 23001 25209
rect 23037 25175 23071 25209
rect 23107 25175 23141 25209
rect 23177 25175 23211 25209
rect 23247 25175 23281 25209
rect 23317 25175 23351 25209
rect 23387 25175 23421 25209
rect 23457 25175 23491 25209
rect 23527 25175 23561 25209
rect 23597 25175 23631 25209
rect 22827 25106 22861 25140
rect 22897 25106 22931 25140
rect 22967 25106 23001 25140
rect 23037 25106 23071 25140
rect 23107 25106 23141 25140
rect 23177 25106 23211 25140
rect 23247 25106 23281 25140
rect 23317 25106 23351 25140
rect 23387 25106 23421 25140
rect 23457 25106 23491 25140
rect 23527 25106 23561 25140
rect 23597 25106 23631 25140
rect 22827 25037 22861 25071
rect 22897 25037 22931 25071
rect 22967 25037 23001 25071
rect 23037 25037 23071 25071
rect 23107 25037 23141 25071
rect 23177 25037 23211 25071
rect 23247 25037 23281 25071
rect 23317 25037 23351 25071
rect 23387 25037 23421 25071
rect 23457 25037 23491 25071
rect 23527 25037 23561 25071
rect 23597 25037 23631 25071
rect 22827 24968 22861 25002
rect 22897 24968 22931 25002
rect 22967 24968 23001 25002
rect 23037 24968 23071 25002
rect 23107 24968 23141 25002
rect 23177 24968 23211 25002
rect 23247 24968 23281 25002
rect 23317 24968 23351 25002
rect 23387 24968 23421 25002
rect 23457 24968 23491 25002
rect 23527 24968 23561 25002
rect 23597 24968 23631 25002
rect 22827 24899 22861 24933
rect 22897 24899 22931 24933
rect 22967 24899 23001 24933
rect 23037 24899 23071 24933
rect 23107 24899 23141 24933
rect 23177 24899 23211 24933
rect 23247 24899 23281 24933
rect 23317 24899 23351 24933
rect 23387 24899 23421 24933
rect 23457 24899 23491 24933
rect 23527 24899 23561 24933
rect 23597 24899 23631 24933
rect 22827 24830 22861 24864
rect 22897 24830 22931 24864
rect 22967 24830 23001 24864
rect 23037 24830 23071 24864
rect 23107 24830 23141 24864
rect 23177 24830 23211 24864
rect 23247 24830 23281 24864
rect 23317 24830 23351 24864
rect 23387 24830 23421 24864
rect 23457 24830 23491 24864
rect 23527 24830 23561 24864
rect 23597 24830 23631 24864
rect 22827 24761 22861 24795
rect 22897 24761 22931 24795
rect 22967 24761 23001 24795
rect 23037 24761 23071 24795
rect 23107 24761 23141 24795
rect 23177 24761 23211 24795
rect 23247 24761 23281 24795
rect 23317 24761 23351 24795
rect 23387 24761 23421 24795
rect 23457 24761 23491 24795
rect 23527 24761 23561 24795
rect 23597 24761 23631 24795
rect 22827 24692 22861 24726
rect 22897 24692 22931 24726
rect 22967 24692 23001 24726
rect 23037 24692 23071 24726
rect 23107 24692 23141 24726
rect 23177 24692 23211 24726
rect 23247 24692 23281 24726
rect 23317 24692 23351 24726
rect 23387 24692 23421 24726
rect 23457 24692 23491 24726
rect 23527 24692 23561 24726
rect 23597 24692 23631 24726
rect 22827 24623 22861 24657
rect 22897 24623 22931 24657
rect 22967 24623 23001 24657
rect 23037 24623 23071 24657
rect 23107 24623 23141 24657
rect 23177 24623 23211 24657
rect 23247 24623 23281 24657
rect 23317 24623 23351 24657
rect 23387 24623 23421 24657
rect 23457 24623 23491 24657
rect 23527 24623 23561 24657
rect 23597 24623 23631 24657
rect 22827 24554 22861 24588
rect 22897 24554 22931 24588
rect 22967 24554 23001 24588
rect 23037 24554 23071 24588
rect 23107 24554 23141 24588
rect 23177 24554 23211 24588
rect 23247 24554 23281 24588
rect 23317 24554 23351 24588
rect 23387 24554 23421 24588
rect 23457 24554 23491 24588
rect 23527 24554 23561 24588
rect 23597 24554 23631 24588
rect 22827 24485 22861 24519
rect 22897 24485 22931 24519
rect 22967 24485 23001 24519
rect 23037 24485 23071 24519
rect 23107 24485 23141 24519
rect 23177 24485 23211 24519
rect 23247 24485 23281 24519
rect 23317 24485 23351 24519
rect 23387 24485 23421 24519
rect 23457 24485 23491 24519
rect 23527 24485 23561 24519
rect 23597 24485 23631 24519
rect 22827 24416 22861 24450
rect 22897 24416 22931 24450
rect 22967 24416 23001 24450
rect 23037 24416 23071 24450
rect 23107 24416 23141 24450
rect 23177 24416 23211 24450
rect 23247 24416 23281 24450
rect 23317 24416 23351 24450
rect 23387 24416 23421 24450
rect 23457 24416 23491 24450
rect 23527 24416 23561 24450
rect 23597 24416 23631 24450
rect 22827 24347 22861 24381
rect 22897 24347 22931 24381
rect 22967 24347 23001 24381
rect 23037 24347 23071 24381
rect 23107 24347 23141 24381
rect 23177 24347 23211 24381
rect 23247 24347 23281 24381
rect 23317 24347 23351 24381
rect 23387 24347 23421 24381
rect 23457 24347 23491 24381
rect 23527 24347 23561 24381
rect 23597 24347 23631 24381
rect 22827 24278 22861 24312
rect 22897 24278 22931 24312
rect 22967 24278 23001 24312
rect 23037 24278 23071 24312
rect 23107 24278 23141 24312
rect 23177 24278 23211 24312
rect 23247 24278 23281 24312
rect 23317 24278 23351 24312
rect 23387 24278 23421 24312
rect 23457 24278 23491 24312
rect 23527 24278 23561 24312
rect 23597 24278 23631 24312
rect 22827 24209 22861 24243
rect 22897 24209 22931 24243
rect 22967 24209 23001 24243
rect 23037 24209 23071 24243
rect 23107 24209 23141 24243
rect 23177 24209 23211 24243
rect 23247 24209 23281 24243
rect 23317 24209 23351 24243
rect 23387 24209 23421 24243
rect 23457 24209 23491 24243
rect 23527 24209 23561 24243
rect 23597 24209 23631 24243
rect 22827 24140 22861 24174
rect 22897 24140 22931 24174
rect 22967 24140 23001 24174
rect 23037 24140 23071 24174
rect 23107 24140 23141 24174
rect 23177 24140 23211 24174
rect 23247 24140 23281 24174
rect 23317 24140 23351 24174
rect 23387 24140 23421 24174
rect 23457 24140 23491 24174
rect 23527 24140 23561 24174
rect 23597 24140 23631 24174
rect 22827 24071 22861 24105
rect 22897 24071 22931 24105
rect 22967 24071 23001 24105
rect 23037 24071 23071 24105
rect 23107 24071 23141 24105
rect 23177 24071 23211 24105
rect 23247 24071 23281 24105
rect 23317 24071 23351 24105
rect 23387 24071 23421 24105
rect 23457 24071 23491 24105
rect 23527 24071 23561 24105
rect 23597 24071 23631 24105
rect 22827 24002 22861 24036
rect 22897 24002 22931 24036
rect 22967 24002 23001 24036
rect 23037 24002 23071 24036
rect 23107 24002 23141 24036
rect 23177 24002 23211 24036
rect 23247 24002 23281 24036
rect 23317 24002 23351 24036
rect 23387 24002 23421 24036
rect 23457 24002 23491 24036
rect 23527 24002 23561 24036
rect 23597 24002 23631 24036
rect 22827 23933 22861 23967
rect 22897 23933 22931 23967
rect 22967 23933 23001 23967
rect 23037 23933 23071 23967
rect 23107 23933 23141 23967
rect 23177 23933 23211 23967
rect 23247 23933 23281 23967
rect 23317 23933 23351 23967
rect 23387 23933 23421 23967
rect 23457 23933 23491 23967
rect 23527 23933 23561 23967
rect 23597 23933 23631 23967
rect 22827 23864 22861 23898
rect 22897 23864 22931 23898
rect 22967 23864 23001 23898
rect 23037 23864 23071 23898
rect 23107 23864 23141 23898
rect 23177 23864 23211 23898
rect 23247 23864 23281 23898
rect 23317 23864 23351 23898
rect 23387 23864 23421 23898
rect 23457 23864 23491 23898
rect 23527 23864 23561 23898
rect 23597 23864 23631 23898
rect 22827 23795 22861 23829
rect 22897 23795 22931 23829
rect 22967 23795 23001 23829
rect 23037 23795 23071 23829
rect 23107 23795 23141 23829
rect 23177 23795 23211 23829
rect 23247 23795 23281 23829
rect 23317 23795 23351 23829
rect 23387 23795 23421 23829
rect 23457 23795 23491 23829
rect 23527 23795 23561 23829
rect 23597 23795 23631 23829
rect 22827 23726 22861 23760
rect 22897 23726 22931 23760
rect 22967 23726 23001 23760
rect 23037 23726 23071 23760
rect 23107 23726 23141 23760
rect 23177 23726 23211 23760
rect 23247 23726 23281 23760
rect 23317 23726 23351 23760
rect 23387 23726 23421 23760
rect 23457 23726 23491 23760
rect 23527 23726 23561 23760
rect 23597 23726 23631 23760
rect 22827 23657 22861 23691
rect 22897 23657 22931 23691
rect 22967 23657 23001 23691
rect 23037 23657 23071 23691
rect 23107 23657 23141 23691
rect 23177 23657 23211 23691
rect 23247 23657 23281 23691
rect 23317 23657 23351 23691
rect 23387 23657 23421 23691
rect 23457 23657 23491 23691
rect 23527 23657 23561 23691
rect 23597 23657 23631 23691
rect 22827 23588 22861 23622
rect 22897 23588 22931 23622
rect 22967 23588 23001 23622
rect 23037 23588 23071 23622
rect 23107 23588 23141 23622
rect 23177 23588 23211 23622
rect 23247 23588 23281 23622
rect 23317 23588 23351 23622
rect 23387 23588 23421 23622
rect 23457 23588 23491 23622
rect 23527 23588 23561 23622
rect 23597 23588 23631 23622
rect 22827 23519 22861 23553
rect 22897 23519 22931 23553
rect 22967 23519 23001 23553
rect 23037 23519 23071 23553
rect 23107 23519 23141 23553
rect 23177 23519 23211 23553
rect 23247 23519 23281 23553
rect 23317 23519 23351 23553
rect 23387 23519 23421 23553
rect 23457 23519 23491 23553
rect 23527 23519 23561 23553
rect 23597 23519 23631 23553
rect 314 23439 348 23473
rect 384 23439 418 23473
rect 454 23439 488 23473
rect 524 23439 558 23473
rect 594 23439 628 23473
rect 664 23439 698 23473
rect 734 23439 768 23473
rect 804 23439 838 23473
rect 874 23439 908 23473
rect 944 23439 978 23473
rect 1014 23439 1048 23473
rect 1084 23439 1118 23473
rect 1154 23439 1188 23473
rect 1224 23439 1258 23473
rect 1294 23439 1328 23473
rect 1364 23439 1398 23473
rect 1434 23439 1468 23473
rect 314 23369 348 23403
rect 384 23369 418 23403
rect 454 23369 488 23403
rect 524 23369 558 23403
rect 594 23369 628 23403
rect 664 23369 698 23403
rect 734 23369 768 23403
rect 804 23369 838 23403
rect 874 23369 908 23403
rect 944 23369 978 23403
rect 1014 23369 1048 23403
rect 1084 23369 1118 23403
rect 1154 23369 1188 23403
rect 1224 23369 1258 23403
rect 1294 23369 1328 23403
rect 1364 23369 1398 23403
rect 1434 23369 1468 23403
rect 314 23299 348 23333
rect 384 23299 418 23333
rect 454 23299 488 23333
rect 524 23299 558 23333
rect 594 23299 628 23333
rect 664 23299 698 23333
rect 734 23299 768 23333
rect 804 23299 838 23333
rect 874 23299 908 23333
rect 944 23299 978 23333
rect 1014 23299 1048 23333
rect 1084 23299 1118 23333
rect 1154 23299 1188 23333
rect 1224 23299 1258 23333
rect 1294 23299 1328 23333
rect 1364 23299 1398 23333
rect 1434 23299 1468 23333
rect 314 23229 348 23263
rect 384 23229 418 23263
rect 454 23229 488 23263
rect 524 23229 558 23263
rect 594 23229 628 23263
rect 664 23229 698 23263
rect 734 23229 768 23263
rect 804 23229 838 23263
rect 874 23229 908 23263
rect 944 23229 978 23263
rect 1014 23229 1048 23263
rect 1084 23229 1118 23263
rect 1154 23229 1188 23263
rect 1224 23229 1258 23263
rect 1294 23229 1328 23263
rect 1364 23229 1398 23263
rect 1434 23229 1468 23263
rect 314 23159 348 23193
rect 384 23159 418 23193
rect 454 23159 488 23193
rect 524 23159 558 23193
rect 594 23159 628 23193
rect 664 23159 698 23193
rect 734 23159 768 23193
rect 804 23159 838 23193
rect 874 23159 908 23193
rect 944 23159 978 23193
rect 1014 23159 1048 23193
rect 1084 23159 1118 23193
rect 1154 23159 1188 23193
rect 1224 23159 1258 23193
rect 1294 23159 1328 23193
rect 1364 23159 1398 23193
rect 1434 23159 1468 23193
rect 314 23089 348 23123
rect 384 23089 418 23123
rect 454 23089 488 23123
rect 524 23089 558 23123
rect 594 23089 628 23123
rect 664 23089 698 23123
rect 734 23089 768 23123
rect 804 23089 838 23123
rect 874 23089 908 23123
rect 944 23089 978 23123
rect 1014 23089 1048 23123
rect 1084 23089 1118 23123
rect 1154 23089 1188 23123
rect 1224 23089 1258 23123
rect 1294 23089 1328 23123
rect 1364 23089 1398 23123
rect 1434 23089 1468 23123
rect 314 23019 348 23053
rect 384 23019 418 23053
rect 454 23019 488 23053
rect 524 23019 558 23053
rect 594 23019 628 23053
rect 664 23019 698 23053
rect 734 23019 768 23053
rect 804 23019 838 23053
rect 874 23019 908 23053
rect 944 23019 978 23053
rect 1014 23019 1048 23053
rect 1084 23019 1118 23053
rect 1154 23019 1188 23053
rect 1224 23019 1258 23053
rect 1294 23019 1328 23053
rect 1364 23019 1398 23053
rect 1434 23019 1468 23053
rect 314 22949 348 22983
rect 384 22949 418 22983
rect 454 22949 488 22983
rect 524 22949 558 22983
rect 594 22949 628 22983
rect 664 22949 698 22983
rect 734 22949 768 22983
rect 804 22949 838 22983
rect 874 22949 908 22983
rect 944 22949 978 22983
rect 1014 22949 1048 22983
rect 1084 22949 1118 22983
rect 1154 22949 1188 22983
rect 1224 22949 1258 22983
rect 1294 22949 1328 22983
rect 1364 22949 1398 22983
rect 1434 22949 1468 22983
rect 314 22879 348 22913
rect 384 22879 418 22913
rect 454 22879 488 22913
rect 524 22879 558 22913
rect 594 22879 628 22913
rect 664 22879 698 22913
rect 734 22879 768 22913
rect 804 22879 838 22913
rect 874 22879 908 22913
rect 944 22879 978 22913
rect 1014 22879 1048 22913
rect 1084 22879 1118 22913
rect 1154 22879 1188 22913
rect 1224 22879 1258 22913
rect 1294 22879 1328 22913
rect 1364 22879 1398 22913
rect 1434 22879 1468 22913
rect 314 22809 348 22843
rect 384 22809 418 22843
rect 454 22809 488 22843
rect 524 22809 558 22843
rect 594 22809 628 22843
rect 664 22809 698 22843
rect 734 22809 768 22843
rect 804 22809 838 22843
rect 874 22809 908 22843
rect 944 22809 978 22843
rect 1014 22809 1048 22843
rect 1084 22809 1118 22843
rect 1154 22809 1188 22843
rect 1224 22809 1258 22843
rect 1294 22809 1328 22843
rect 1364 22809 1398 22843
rect 1434 22809 1468 22843
rect 314 22739 348 22773
rect 384 22739 418 22773
rect 454 22739 488 22773
rect 524 22739 558 22773
rect 594 22739 628 22773
rect 664 22739 698 22773
rect 734 22739 768 22773
rect 804 22739 838 22773
rect 874 22739 908 22773
rect 944 22739 978 22773
rect 1014 22739 1048 22773
rect 1084 22739 1118 22773
rect 1154 22739 1188 22773
rect 1224 22739 1258 22773
rect 1294 22739 1328 22773
rect 1364 22739 1398 22773
rect 1434 22739 1468 22773
rect 314 22668 348 22702
rect 384 22668 418 22702
rect 454 22668 488 22702
rect 524 22668 558 22702
rect 594 22668 628 22702
rect 664 22668 698 22702
rect 734 22668 768 22702
rect 804 22668 838 22702
rect 874 22668 908 22702
rect 944 22668 978 22702
rect 1014 22668 1048 22702
rect 1084 22668 1118 22702
rect 1154 22668 1188 22702
rect 1224 22668 1258 22702
rect 1294 22668 1328 22702
rect 1364 22668 1398 22702
rect 1434 22668 1468 22702
rect 314 22597 348 22631
rect 384 22597 418 22631
rect 454 22597 488 22631
rect 524 22597 558 22631
rect 594 22597 628 22631
rect 664 22597 698 22631
rect 734 22597 768 22631
rect 804 22597 838 22631
rect 874 22597 908 22631
rect 944 22597 978 22631
rect 1014 22597 1048 22631
rect 1084 22597 1118 22631
rect 1154 22597 1188 22631
rect 1224 22597 1258 22631
rect 1294 22597 1328 22631
rect 1364 22597 1398 22631
rect 1434 22597 1468 22631
rect 314 22526 348 22560
rect 384 22526 418 22560
rect 454 22526 488 22560
rect 524 22526 558 22560
rect 594 22526 628 22560
rect 664 22526 698 22560
rect 734 22526 768 22560
rect 804 22526 838 22560
rect 874 22526 908 22560
rect 944 22526 978 22560
rect 1014 22526 1048 22560
rect 1084 22526 1118 22560
rect 1154 22526 1188 22560
rect 1224 22526 1258 22560
rect 1294 22526 1328 22560
rect 1364 22526 1398 22560
rect 1434 22526 1468 22560
rect 314 22455 348 22489
rect 384 22455 418 22489
rect 454 22455 488 22489
rect 524 22455 558 22489
rect 594 22455 628 22489
rect 664 22455 698 22489
rect 734 22455 768 22489
rect 804 22455 838 22489
rect 874 22455 908 22489
rect 944 22455 978 22489
rect 1014 22455 1048 22489
rect 1084 22455 1118 22489
rect 1154 22455 1188 22489
rect 1224 22455 1258 22489
rect 1294 22455 1328 22489
rect 1364 22455 1398 22489
rect 1434 22455 1468 22489
rect 314 22384 348 22418
rect 384 22384 418 22418
rect 454 22384 488 22418
rect 524 22384 558 22418
rect 594 22384 628 22418
rect 664 22384 698 22418
rect 734 22384 768 22418
rect 804 22384 838 22418
rect 874 22384 908 22418
rect 944 22384 978 22418
rect 1014 22384 1048 22418
rect 1084 22384 1118 22418
rect 1154 22384 1188 22418
rect 1224 22384 1258 22418
rect 1294 22384 1328 22418
rect 1364 22384 1398 22418
rect 1434 22384 1468 22418
rect 314 22313 348 22347
rect 384 22313 418 22347
rect 454 22313 488 22347
rect 524 22313 558 22347
rect 594 22313 628 22347
rect 664 22313 698 22347
rect 734 22313 768 22347
rect 804 22313 838 22347
rect 874 22313 908 22347
rect 944 22313 978 22347
rect 1014 22313 1048 22347
rect 1084 22313 1118 22347
rect 1154 22313 1188 22347
rect 1224 22313 1258 22347
rect 1294 22313 1328 22347
rect 1364 22313 1398 22347
rect 1434 22313 1468 22347
rect 22827 23450 22861 23484
rect 22897 23450 22931 23484
rect 22967 23450 23001 23484
rect 23037 23450 23071 23484
rect 23107 23450 23141 23484
rect 23177 23450 23211 23484
rect 23247 23450 23281 23484
rect 23317 23450 23351 23484
rect 23387 23450 23421 23484
rect 23457 23450 23491 23484
rect 23527 23450 23561 23484
rect 23597 23450 23631 23484
rect 22827 23381 22861 23415
rect 22897 23381 22931 23415
rect 22967 23381 23001 23415
rect 23037 23381 23071 23415
rect 23107 23381 23141 23415
rect 23177 23381 23211 23415
rect 23247 23381 23281 23415
rect 23317 23381 23351 23415
rect 23387 23381 23421 23415
rect 23457 23381 23491 23415
rect 23527 23381 23561 23415
rect 23597 23381 23631 23415
rect 22827 23312 22861 23346
rect 22897 23312 22931 23346
rect 22967 23312 23001 23346
rect 23037 23312 23071 23346
rect 23107 23312 23141 23346
rect 23177 23312 23211 23346
rect 23247 23312 23281 23346
rect 23317 23312 23351 23346
rect 23387 23312 23421 23346
rect 23457 23312 23491 23346
rect 23527 23312 23561 23346
rect 23597 23312 23631 23346
rect 22827 23243 22861 23277
rect 22897 23243 22931 23277
rect 22967 23243 23001 23277
rect 23037 23243 23071 23277
rect 23107 23243 23141 23277
rect 23177 23243 23211 23277
rect 23247 23243 23281 23277
rect 23317 23243 23351 23277
rect 23387 23243 23421 23277
rect 23457 23243 23491 23277
rect 23527 23243 23561 23277
rect 23597 23243 23631 23277
rect 22827 23174 22861 23208
rect 22897 23174 22931 23208
rect 22967 23174 23001 23208
rect 23037 23174 23071 23208
rect 23107 23174 23141 23208
rect 23177 23174 23211 23208
rect 23247 23174 23281 23208
rect 23317 23174 23351 23208
rect 23387 23174 23421 23208
rect 23457 23174 23491 23208
rect 23527 23174 23561 23208
rect 23597 23174 23631 23208
rect 22827 23105 22861 23139
rect 22897 23105 22931 23139
rect 22967 23105 23001 23139
rect 23037 23105 23071 23139
rect 23107 23105 23141 23139
rect 23177 23105 23211 23139
rect 23247 23105 23281 23139
rect 23317 23105 23351 23139
rect 23387 23105 23421 23139
rect 23457 23105 23491 23139
rect 23527 23105 23561 23139
rect 23597 23105 23631 23139
rect 22827 23036 22861 23070
rect 22897 23036 22931 23070
rect 22967 23036 23001 23070
rect 23037 23036 23071 23070
rect 23107 23036 23141 23070
rect 23177 23036 23211 23070
rect 23247 23036 23281 23070
rect 23317 23036 23351 23070
rect 23387 23036 23421 23070
rect 23457 23036 23491 23070
rect 23527 23036 23561 23070
rect 23597 23036 23631 23070
rect 22827 22967 22861 23001
rect 22897 22967 22931 23001
rect 22967 22967 23001 23001
rect 23037 22967 23071 23001
rect 23107 22967 23141 23001
rect 23177 22967 23211 23001
rect 23247 22967 23281 23001
rect 23317 22967 23351 23001
rect 23387 22967 23421 23001
rect 23457 22967 23491 23001
rect 23527 22967 23561 23001
rect 23597 22967 23631 23001
rect 22827 22898 22861 22932
rect 22897 22898 22931 22932
rect 22967 22898 23001 22932
rect 23037 22898 23071 22932
rect 23107 22898 23141 22932
rect 23177 22898 23211 22932
rect 23247 22898 23281 22932
rect 23317 22898 23351 22932
rect 23387 22898 23421 22932
rect 23457 22898 23491 22932
rect 23527 22898 23561 22932
rect 23597 22898 23631 22932
rect 22827 22829 22861 22863
rect 22897 22829 22931 22863
rect 22967 22829 23001 22863
rect 23037 22829 23071 22863
rect 23107 22829 23141 22863
rect 23177 22829 23211 22863
rect 23247 22829 23281 22863
rect 23317 22829 23351 22863
rect 23387 22829 23421 22863
rect 23457 22829 23491 22863
rect 23527 22829 23561 22863
rect 23597 22829 23631 22863
rect 22827 22760 22861 22794
rect 22897 22760 22931 22794
rect 22967 22760 23001 22794
rect 23037 22760 23071 22794
rect 23107 22760 23141 22794
rect 23177 22760 23211 22794
rect 23247 22760 23281 22794
rect 23317 22760 23351 22794
rect 23387 22760 23421 22794
rect 23457 22760 23491 22794
rect 23527 22760 23561 22794
rect 23597 22760 23631 22794
rect 22827 22691 22861 22725
rect 22897 22691 22931 22725
rect 22967 22691 23001 22725
rect 23037 22691 23071 22725
rect 23107 22691 23141 22725
rect 23177 22691 23211 22725
rect 23247 22691 23281 22725
rect 23317 22691 23351 22725
rect 23387 22691 23421 22725
rect 23457 22691 23491 22725
rect 23527 22691 23561 22725
rect 23597 22691 23631 22725
rect 22827 22622 22861 22656
rect 22897 22622 22931 22656
rect 22967 22622 23001 22656
rect 23037 22622 23071 22656
rect 23107 22622 23141 22656
rect 23177 22622 23211 22656
rect 23247 22622 23281 22656
rect 23317 22622 23351 22656
rect 23387 22622 23421 22656
rect 23457 22622 23491 22656
rect 23527 22622 23561 22656
rect 23597 22622 23631 22656
rect 22827 22553 22861 22587
rect 22897 22553 22931 22587
rect 22967 22553 23001 22587
rect 23037 22553 23071 22587
rect 23107 22553 23141 22587
rect 23177 22553 23211 22587
rect 23247 22553 23281 22587
rect 23317 22553 23351 22587
rect 23387 22553 23421 22587
rect 23457 22553 23491 22587
rect 23527 22553 23561 22587
rect 23597 22553 23631 22587
rect 22827 22484 22861 22518
rect 22897 22484 22931 22518
rect 22967 22484 23001 22518
rect 23037 22484 23071 22518
rect 23107 22484 23141 22518
rect 23177 22484 23211 22518
rect 23247 22484 23281 22518
rect 23317 22484 23351 22518
rect 23387 22484 23421 22518
rect 23457 22484 23491 22518
rect 23527 22484 23561 22518
rect 23597 22484 23631 22518
rect 22827 22415 22861 22449
rect 22897 22415 22931 22449
rect 22967 22415 23001 22449
rect 23037 22415 23071 22449
rect 23107 22415 23141 22449
rect 23177 22415 23211 22449
rect 23247 22415 23281 22449
rect 23317 22415 23351 22449
rect 23387 22415 23421 22449
rect 23457 22415 23491 22449
rect 23527 22415 23561 22449
rect 23597 22415 23631 22449
rect 22827 22346 22861 22380
rect 22897 22346 22931 22380
rect 22967 22346 23001 22380
rect 23037 22346 23071 22380
rect 23107 22346 23141 22380
rect 23177 22346 23211 22380
rect 23247 22346 23281 22380
rect 23317 22346 23351 22380
rect 23387 22346 23421 22380
rect 23457 22346 23491 22380
rect 23527 22346 23561 22380
rect 23597 22346 23631 22380
rect 714 17419 1020 22213
rect 22827 22277 22861 22311
rect 22897 22277 22931 22311
rect 22967 22277 23001 22311
rect 23037 22277 23071 22311
rect 23107 22277 23141 22311
rect 23177 22277 23211 22311
rect 23247 22277 23281 22311
rect 23317 22277 23351 22311
rect 23387 22277 23421 22311
rect 23457 22277 23491 22311
rect 23527 22277 23561 22311
rect 23597 22277 23631 22311
rect 22827 22208 22861 22242
rect 22897 22208 22931 22242
rect 22967 22208 23001 22242
rect 23037 22208 23071 22242
rect 23107 22208 23141 22242
rect 23177 22208 23211 22242
rect 23247 22208 23281 22242
rect 23317 22208 23351 22242
rect 23387 22208 23421 22242
rect 23457 22208 23491 22242
rect 23527 22208 23561 22242
rect 23597 22208 23631 22242
rect 22827 22139 22861 22173
rect 22897 22139 22931 22173
rect 22967 22139 23001 22173
rect 23037 22139 23071 22173
rect 23107 22139 23141 22173
rect 23177 22139 23211 22173
rect 23247 22139 23281 22173
rect 23317 22139 23351 22173
rect 23387 22139 23421 22173
rect 23457 22139 23491 22173
rect 23527 22139 23561 22173
rect 23597 22139 23631 22173
rect 714 17350 748 17384
rect 782 17350 816 17384
rect 850 17350 884 17384
rect 918 17350 952 17384
rect 986 17350 1020 17384
rect 714 17281 748 17315
rect 782 17281 816 17315
rect 850 17281 884 17315
rect 918 17281 952 17315
rect 986 17281 1020 17315
rect 714 17212 748 17246
rect 782 17212 816 17246
rect 850 17212 884 17246
rect 918 17212 952 17246
rect 986 17212 1020 17246
rect 714 17143 748 17177
rect 782 17143 816 17177
rect 850 17143 884 17177
rect 918 17143 952 17177
rect 986 17143 1020 17177
rect 714 17074 748 17108
rect 782 17074 816 17108
rect 850 17074 884 17108
rect 918 17074 952 17108
rect 986 17074 1020 17108
rect 714 17005 748 17039
rect 782 17005 816 17039
rect 850 17005 884 17039
rect 918 17005 952 17039
rect 986 17005 1020 17039
rect 714 16936 748 16970
rect 782 16936 816 16970
rect 850 16936 884 16970
rect 918 16936 952 16970
rect 986 16936 1020 16970
rect 714 16867 748 16901
rect 782 16867 816 16901
rect 850 16867 884 16901
rect 918 16867 952 16901
rect 986 16867 1020 16901
rect 714 16798 748 16832
rect 782 16798 816 16832
rect 850 16798 884 16832
rect 918 16798 952 16832
rect 986 16798 1020 16832
rect 714 16729 748 16763
rect 782 16729 816 16763
rect 850 16729 884 16763
rect 918 16729 952 16763
rect 986 16729 1020 16763
rect 714 16660 748 16694
rect 782 16660 816 16694
rect 850 16660 884 16694
rect 918 16660 952 16694
rect 986 16660 1020 16694
rect 714 16591 748 16625
rect 782 16591 816 16625
rect 850 16591 884 16625
rect 918 16591 952 16625
rect 986 16591 1020 16625
rect 714 16522 748 16556
rect 782 16522 816 16556
rect 850 16522 884 16556
rect 918 16522 952 16556
rect 986 16522 1020 16556
rect 714 16453 748 16487
rect 782 16453 816 16487
rect 850 16453 884 16487
rect 918 16453 952 16487
rect 986 16453 1020 16487
rect 714 16384 748 16418
rect 782 16384 816 16418
rect 850 16384 884 16418
rect 918 16384 952 16418
rect 986 16384 1020 16418
rect 714 16315 748 16349
rect 782 16315 816 16349
rect 850 16315 884 16349
rect 918 16315 952 16349
rect 986 16315 1020 16349
rect 714 16246 748 16280
rect 782 16246 816 16280
rect 850 16246 884 16280
rect 918 16246 952 16280
rect 986 16246 1020 16280
rect 6770 11584 6804 11618
rect 6839 11584 6873 11618
rect 6908 11584 6942 11618
rect 6977 11584 7011 11618
rect 7046 11584 7080 11618
rect 7115 11584 7149 11618
rect 7184 11584 7218 11618
rect 7253 11584 7287 11618
rect 7322 11584 7356 11618
rect 7391 11584 7425 11618
rect 7460 11584 7494 11618
rect 7529 11584 7563 11618
rect 7598 11584 7632 11618
rect 7667 11584 7701 11618
rect 7736 11584 7770 11618
rect 7805 11584 7839 11618
rect 7874 11584 7908 11618
rect 7943 11584 7977 11618
rect 8012 11584 8046 11618
rect 8081 11584 8115 11618
rect 8150 11584 8184 11618
rect 8219 11584 8253 11618
rect 8288 11584 8322 11618
rect 8357 11584 8391 11618
rect 8426 11584 8460 11618
rect 8495 11584 8529 11618
rect 8564 11584 8598 11618
rect 8633 11584 8667 11618
rect 8702 11584 8736 11618
rect 8771 11584 8805 11618
rect 8840 11584 8874 11618
rect 8909 11584 8943 11618
rect 8978 11584 9012 11618
rect 9046 11584 9080 11618
rect 9114 11584 9148 11618
rect 9182 11584 9216 11618
rect 9250 11584 9284 11618
rect 9318 11584 9352 11618
rect 9386 11584 9420 11618
rect 9454 11584 9488 11618
rect 9522 11584 9556 11618
rect 9590 11584 9624 11618
rect 9658 11584 9692 11618
rect 9726 11584 9760 11618
rect 9794 11584 9828 11618
rect 9862 11584 9896 11618
rect 9930 11584 9964 11618
rect 9998 11584 10032 11618
rect 10066 11584 10100 11618
rect 10134 11584 10168 11618
rect 10202 11584 10236 11618
rect 10270 11584 10304 11618
rect 16309 11588 16343 11622
rect 16379 11588 16413 11622
rect 16449 11588 16483 11622
rect 16519 11588 16553 11622
rect 16589 11588 16623 11622
rect 16658 11588 16692 11622
rect 16727 11588 16761 11622
rect 16796 11588 16830 11622
rect 16865 11588 16899 11622
rect 16934 11588 16968 11622
rect 17003 11588 17037 11622
rect 17072 11588 17106 11622
rect 17141 11588 17175 11622
rect 17210 11588 17244 11622
rect 17279 11588 17313 11622
rect 17348 11588 17382 11622
rect 17417 11588 17451 11622
rect 17486 11588 17520 11622
rect 17555 11588 17589 11622
rect 17624 11588 17658 11622
rect 17693 11588 17727 11622
rect 17762 11588 17796 11622
rect 17831 11588 17865 11622
rect 17900 11588 17934 11622
rect 17969 11588 18003 11622
rect 18038 11588 18072 11622
rect 18107 11588 18141 11622
rect 18176 11588 18210 11622
rect 18245 11588 18279 11622
rect 18314 11588 18348 11622
rect 18383 11588 18417 11622
rect 18452 11588 18486 11622
rect 18521 11588 18555 11622
rect 18590 11588 18624 11622
rect 18659 11588 18693 11622
rect 18728 11588 18762 11622
rect 18797 11588 18831 11622
rect 18866 11588 18900 11622
rect 18935 11588 18969 11622
rect 19004 11588 19038 11622
rect 19073 11588 19107 11622
rect 19142 11588 19176 11622
rect 19211 11588 19245 11622
rect 19280 11588 19314 11622
rect 19349 11588 19383 11622
rect 19418 11588 19452 11622
rect 19487 11588 19521 11622
rect 19556 11588 19590 11622
rect 19625 11588 19659 11622
rect 19797 11595 19831 11629
rect 19866 11595 19900 11629
rect 19935 11595 19969 11629
rect 20004 11595 20038 11629
rect 20073 11595 20107 11629
rect 20142 11595 20176 11629
rect 20211 11595 20245 11629
rect 20280 11595 20314 11629
rect 20349 11595 20383 11629
rect 20418 11595 20452 11629
rect 20487 11595 20521 11629
rect 20556 11595 20590 11629
rect 20625 11595 20659 11629
rect 20694 11595 20728 11629
rect 20763 11595 20797 11629
rect 20832 11595 20866 11629
rect 20901 11595 20935 11629
rect 20970 11595 21004 11629
rect 21039 11595 21073 11629
rect 21108 11595 21142 11629
rect 21177 11595 21211 11629
rect 21246 11595 21280 11629
rect 21315 11595 21349 11629
rect 21384 11595 21418 11629
rect 21453 11595 21487 11629
rect 21522 11595 21556 11629
rect 21591 11595 21625 11629
rect 21660 11595 21694 11629
rect 21729 11595 21763 11629
rect 21798 11595 21832 11629
rect 21866 11595 21900 11629
rect 21934 11595 21968 11629
rect 22002 11595 22036 11629
rect 22070 11595 22104 11629
rect 22138 11595 22172 11629
rect 22206 11595 22240 11629
rect 22274 11595 22308 11629
rect 22342 11595 22376 11629
rect 22410 11595 22444 11629
rect 22478 11595 22512 11629
rect 22546 11595 22580 11629
rect 22614 11595 22648 11629
rect 22682 11595 22716 11629
rect 22750 11595 22784 11629
rect 22818 11595 22852 11629
rect 22886 11595 22920 11629
rect 22954 11595 22988 11629
rect 23022 11595 23056 11629
rect 23090 11595 23124 11629
rect 23158 11595 23192 11629
rect 23226 11595 23260 11629
rect 23294 11595 23328 11629
rect 23362 11595 23396 11629
rect 23430 11595 23464 11629
rect 23498 11595 23532 11629
rect 23566 11595 23600 11629
rect 23634 11595 23668 11629
rect 23702 11595 23736 11629
rect 23770 11595 23804 11629
rect 23838 11595 23872 11629
rect 23906 11595 23940 11629
rect 23974 11595 24008 11629
rect 24042 11595 24076 11629
rect 24110 11595 24144 11629
rect 24178 11595 24212 11629
rect 24246 11595 24280 11629
rect 24314 11595 24348 11629
rect 24382 11595 24416 11629
rect 24450 11595 24484 11629
rect 24518 11595 24552 11629
rect 24586 11595 24620 11629
rect 24654 11595 24688 11629
rect 24722 11595 24756 11629
rect 24790 11595 24824 11629
rect 24858 11595 24892 11629
rect 24926 11595 24960 11629
rect 24994 11595 25028 11629
rect 25062 11595 25096 11629
rect 25130 11595 25164 11629
rect 25198 11595 25232 11629
rect 25266 11595 25300 11629
rect 25334 11595 25368 11629
rect 25402 11595 25436 11629
rect 25470 11595 25504 11629
rect 6770 11512 6804 11546
rect 6839 11512 6873 11546
rect 6908 11512 6942 11546
rect 6977 11512 7011 11546
rect 7046 11512 7080 11546
rect 7115 11512 7149 11546
rect 7184 11512 7218 11546
rect 7253 11512 7287 11546
rect 7322 11512 7356 11546
rect 7391 11512 7425 11546
rect 7460 11512 7494 11546
rect 7529 11512 7563 11546
rect 7598 11512 7632 11546
rect 7667 11512 7701 11546
rect 7736 11512 7770 11546
rect 7805 11512 7839 11546
rect 7874 11512 7908 11546
rect 7943 11512 7977 11546
rect 8012 11512 8046 11546
rect 8081 11512 8115 11546
rect 8150 11512 8184 11546
rect 8219 11512 8253 11546
rect 8288 11512 8322 11546
rect 8357 11512 8391 11546
rect 8426 11512 8460 11546
rect 8495 11512 8529 11546
rect 8564 11512 8598 11546
rect 8633 11512 8667 11546
rect 8702 11512 8736 11546
rect 8771 11512 8805 11546
rect 8840 11512 8874 11546
rect 8909 11512 8943 11546
rect 8978 11512 9012 11546
rect 9046 11512 9080 11546
rect 9114 11512 9148 11546
rect 9182 11512 9216 11546
rect 9250 11512 9284 11546
rect 9318 11512 9352 11546
rect 9386 11512 9420 11546
rect 9454 11512 9488 11546
rect 9522 11512 9556 11546
rect 9590 11512 9624 11546
rect 9658 11512 9692 11546
rect 9726 11512 9760 11546
rect 9794 11512 9828 11546
rect 9862 11512 9896 11546
rect 9930 11512 9964 11546
rect 9998 11512 10032 11546
rect 10066 11512 10100 11546
rect 10134 11512 10168 11546
rect 10202 11512 10236 11546
rect 10270 11512 10304 11546
rect 10404 11543 10438 11577
rect 10473 11543 10507 11577
rect 10542 11543 10576 11577
rect 10611 11543 10645 11577
rect 10680 11543 10714 11577
rect 10749 11543 10783 11577
rect 10818 11543 10852 11577
rect 10887 11543 10921 11577
rect 10956 11543 10990 11577
rect 11025 11543 11059 11577
rect 11094 11543 11128 11577
rect 11163 11543 11197 11577
rect 11232 11543 11266 11577
rect 11301 11543 11335 11577
rect 11370 11543 11404 11577
rect 11439 11543 11473 11577
rect 11508 11543 11542 11577
rect 11577 11543 11611 11577
rect 11646 11543 11680 11577
rect 11715 11543 11749 11577
rect 11784 11543 11818 11577
rect 11853 11543 11887 11577
rect 11922 11543 11956 11577
rect 11991 11543 12025 11577
rect 12060 11543 12094 11577
rect 12129 11543 12163 11577
rect 12198 11543 12232 11577
rect 12267 11543 12301 11577
rect 12336 11543 12370 11577
rect 12405 11543 12439 11577
rect 12474 11543 12508 11577
rect 12543 11543 12577 11577
rect 12612 11543 12646 11577
rect 12681 11543 12715 11577
rect 12750 11543 12784 11577
rect 12819 11543 12853 11577
rect 12888 11543 12922 11577
rect 12957 11543 12991 11577
rect 13026 11543 13060 11577
rect 13095 11543 13129 11577
rect 13164 11543 13198 11577
rect 13233 11543 13267 11577
rect 13302 11543 13336 11577
rect 10404 11475 10438 11509
rect 10473 11475 10507 11509
rect 10542 11475 10576 11509
rect 10611 11475 10645 11509
rect 10680 11475 10714 11509
rect 10749 11475 10783 11509
rect 10818 11475 10852 11509
rect 10887 11475 10921 11509
rect 10956 11475 10990 11509
rect 11025 11475 11059 11509
rect 11094 11475 11128 11509
rect 11163 11475 11197 11509
rect 11232 11475 11266 11509
rect 11301 11475 11335 11509
rect 11370 11475 11404 11509
rect 11439 11475 11473 11509
rect 11508 11475 11542 11509
rect 11577 11475 11611 11509
rect 11646 11475 11680 11509
rect 11715 11475 11749 11509
rect 11784 11475 11818 11509
rect 11853 11475 11887 11509
rect 11922 11475 11956 11509
rect 11991 11475 12025 11509
rect 12060 11475 12094 11509
rect 12129 11475 12163 11509
rect 12198 11475 12232 11509
rect 12267 11475 12301 11509
rect 12336 11475 12370 11509
rect 12405 11475 12439 11509
rect 12474 11475 12508 11509
rect 12543 11475 12577 11509
rect 12612 11475 12646 11509
rect 12681 11475 12715 11509
rect 12750 11475 12784 11509
rect 12819 11475 12853 11509
rect 12888 11475 12922 11509
rect 12957 11475 12991 11509
rect 13026 11475 13060 11509
rect 13095 11475 13129 11509
rect 13164 11475 13198 11509
rect 13233 11475 13267 11509
rect 13302 11475 13336 11509
rect 6770 11440 6804 11474
rect 6839 11440 6873 11474
rect 6908 11440 6942 11474
rect 6977 11440 7011 11474
rect 7046 11440 7080 11474
rect 7115 11440 7149 11474
rect 7184 11440 7218 11474
rect 7253 11440 7287 11474
rect 7322 11440 7356 11474
rect 7391 11440 7425 11474
rect 7460 11440 7494 11474
rect 7529 11440 7563 11474
rect 7598 11440 7632 11474
rect 7667 11440 7701 11474
rect 7736 11440 7770 11474
rect 7805 11440 7839 11474
rect 7874 11440 7908 11474
rect 7943 11440 7977 11474
rect 8012 11440 8046 11474
rect 8081 11440 8115 11474
rect 8150 11440 8184 11474
rect 8219 11440 8253 11474
rect 8288 11440 8322 11474
rect 8357 11440 8391 11474
rect 8426 11440 8460 11474
rect 8495 11440 8529 11474
rect 8564 11440 8598 11474
rect 8633 11440 8667 11474
rect 8702 11440 8736 11474
rect 8771 11440 8805 11474
rect 8840 11440 8874 11474
rect 8909 11440 8943 11474
rect 8978 11440 9012 11474
rect 9046 11440 9080 11474
rect 9114 11440 9148 11474
rect 9182 11440 9216 11474
rect 9250 11440 9284 11474
rect 9318 11440 9352 11474
rect 9386 11440 9420 11474
rect 9454 11440 9488 11474
rect 9522 11440 9556 11474
rect 9590 11440 9624 11474
rect 9658 11440 9692 11474
rect 9726 11440 9760 11474
rect 9794 11440 9828 11474
rect 9862 11440 9896 11474
rect 9930 11440 9964 11474
rect 9998 11440 10032 11474
rect 10066 11440 10100 11474
rect 10134 11440 10168 11474
rect 10202 11440 10236 11474
rect 10270 11440 10304 11474
rect 10404 11407 10438 11441
rect 10473 11407 10507 11441
rect 10542 11407 10576 11441
rect 10611 11407 10645 11441
rect 10680 11407 10714 11441
rect 10749 11407 10783 11441
rect 10818 11407 10852 11441
rect 10887 11407 10921 11441
rect 10956 11407 10990 11441
rect 11025 11407 11059 11441
rect 11094 11407 11128 11441
rect 11163 11407 11197 11441
rect 11232 11407 11266 11441
rect 11301 11407 11335 11441
rect 11370 11407 11404 11441
rect 11439 11407 11473 11441
rect 11508 11407 11542 11441
rect 11577 11407 11611 11441
rect 11646 11407 11680 11441
rect 11715 11407 11749 11441
rect 11784 11407 11818 11441
rect 11853 11407 11887 11441
rect 11922 11407 11956 11441
rect 11991 11407 12025 11441
rect 12060 11407 12094 11441
rect 12129 11407 12163 11441
rect 12198 11407 12232 11441
rect 12267 11407 12301 11441
rect 12336 11407 12370 11441
rect 12405 11407 12439 11441
rect 12474 11407 12508 11441
rect 12543 11407 12577 11441
rect 12612 11407 12646 11441
rect 12681 11407 12715 11441
rect 12750 11407 12784 11441
rect 12819 11407 12853 11441
rect 12888 11407 12922 11441
rect 12957 11407 12991 11441
rect 13026 11407 13060 11441
rect 13095 11407 13129 11441
rect 13164 11407 13198 11441
rect 13233 11407 13267 11441
rect 13302 11407 13336 11441
rect 13371 11407 16261 11577
rect 16309 11520 16343 11554
rect 16379 11520 16413 11554
rect 16449 11520 16483 11554
rect 16519 11520 16553 11554
rect 16589 11520 16623 11554
rect 16658 11520 16692 11554
rect 16727 11520 16761 11554
rect 16796 11520 16830 11554
rect 16865 11520 16899 11554
rect 16934 11520 16968 11554
rect 17003 11520 17037 11554
rect 17072 11520 17106 11554
rect 17141 11520 17175 11554
rect 17210 11520 17244 11554
rect 17279 11520 17313 11554
rect 17348 11520 17382 11554
rect 17417 11520 17451 11554
rect 17486 11520 17520 11554
rect 17555 11520 17589 11554
rect 17624 11520 17658 11554
rect 17693 11520 17727 11554
rect 17762 11520 17796 11554
rect 17831 11520 17865 11554
rect 17900 11520 17934 11554
rect 17969 11520 18003 11554
rect 18038 11520 18072 11554
rect 18107 11520 18141 11554
rect 18176 11520 18210 11554
rect 18245 11520 18279 11554
rect 18314 11520 18348 11554
rect 18383 11520 18417 11554
rect 18452 11520 18486 11554
rect 18521 11520 18555 11554
rect 18590 11520 18624 11554
rect 18659 11520 18693 11554
rect 18728 11520 18762 11554
rect 18797 11520 18831 11554
rect 18866 11520 18900 11554
rect 18935 11520 18969 11554
rect 19004 11520 19038 11554
rect 19073 11520 19107 11554
rect 19142 11520 19176 11554
rect 19211 11520 19245 11554
rect 19280 11520 19314 11554
rect 19349 11520 19383 11554
rect 19418 11520 19452 11554
rect 19487 11520 19521 11554
rect 19556 11520 19590 11554
rect 19625 11520 19659 11554
rect 16309 11452 16343 11486
rect 16379 11452 16413 11486
rect 16449 11452 16483 11486
rect 16519 11452 16553 11486
rect 16589 11452 16623 11486
rect 16658 11452 16692 11486
rect 16727 11452 16761 11486
rect 16796 11452 16830 11486
rect 16865 11452 16899 11486
rect 16934 11452 16968 11486
rect 17003 11452 17037 11486
rect 17072 11452 17106 11486
rect 17141 11452 17175 11486
rect 17210 11452 17244 11486
rect 17279 11452 17313 11486
rect 17348 11452 17382 11486
rect 17417 11452 17451 11486
rect 17486 11452 17520 11486
rect 17555 11452 17589 11486
rect 17624 11452 17658 11486
rect 17693 11452 17727 11486
rect 17762 11452 17796 11486
rect 17831 11452 17865 11486
rect 17900 11452 17934 11486
rect 17969 11452 18003 11486
rect 18038 11452 18072 11486
rect 18107 11452 18141 11486
rect 18176 11452 18210 11486
rect 18245 11452 18279 11486
rect 18314 11452 18348 11486
rect 18383 11452 18417 11486
rect 18452 11452 18486 11486
rect 18521 11452 18555 11486
rect 18590 11452 18624 11486
rect 18659 11452 18693 11486
rect 18728 11452 18762 11486
rect 18797 11452 18831 11486
rect 18866 11452 18900 11486
rect 18935 11452 18969 11486
rect 19004 11452 19038 11486
rect 19073 11452 19107 11486
rect 19142 11452 19176 11486
rect 19211 11452 19245 11486
rect 19280 11452 19314 11486
rect 19349 11452 19383 11486
rect 19418 11452 19452 11486
rect 19487 11452 19521 11486
rect 19556 11452 19590 11486
rect 19625 11452 19659 11486
rect 6770 11368 6804 11402
rect 6839 11368 6873 11402
rect 6908 11368 6942 11402
rect 6977 11368 7011 11402
rect 7046 11368 7080 11402
rect 7115 11368 7149 11402
rect 7184 11368 7218 11402
rect 7253 11368 7287 11402
rect 7322 11368 7356 11402
rect 7391 11368 7425 11402
rect 7460 11368 7494 11402
rect 7529 11368 7563 11402
rect 7598 11368 7632 11402
rect 7667 11368 7701 11402
rect 7736 11368 7770 11402
rect 7805 11368 7839 11402
rect 7874 11368 7908 11402
rect 7943 11368 7977 11402
rect 8012 11368 8046 11402
rect 8081 11368 8115 11402
rect 8150 11368 8184 11402
rect 8219 11368 8253 11402
rect 8288 11368 8322 11402
rect 8357 11368 8391 11402
rect 8426 11368 8460 11402
rect 8495 11368 8529 11402
rect 8564 11368 8598 11402
rect 8633 11368 8667 11402
rect 8702 11368 8736 11402
rect 8771 11368 8805 11402
rect 8840 11368 8874 11402
rect 8909 11368 8943 11402
rect 8978 11368 9012 11402
rect 9046 11368 9080 11402
rect 9114 11368 9148 11402
rect 9182 11368 9216 11402
rect 9250 11368 9284 11402
rect 9318 11368 9352 11402
rect 9386 11368 9420 11402
rect 9454 11368 9488 11402
rect 9522 11368 9556 11402
rect 9590 11368 9624 11402
rect 9658 11368 9692 11402
rect 9726 11368 9760 11402
rect 9794 11368 9828 11402
rect 9862 11368 9896 11402
rect 9930 11368 9964 11402
rect 9998 11368 10032 11402
rect 10066 11368 10100 11402
rect 10134 11368 10168 11402
rect 10202 11368 10236 11402
rect 10270 11368 10304 11402
rect 16309 11384 16343 11418
rect 16379 11384 16413 11418
rect 16449 11384 16483 11418
rect 16519 11384 16553 11418
rect 16589 11384 16623 11418
rect 16658 11384 16692 11418
rect 16727 11384 16761 11418
rect 16796 11384 16830 11418
rect 16865 11384 16899 11418
rect 16934 11384 16968 11418
rect 17003 11384 17037 11418
rect 17072 11384 17106 11418
rect 17141 11384 17175 11418
rect 17210 11384 17244 11418
rect 17279 11384 17313 11418
rect 17348 11384 17382 11418
rect 17417 11384 17451 11418
rect 17486 11384 17520 11418
rect 17555 11384 17589 11418
rect 17624 11384 17658 11418
rect 17693 11384 17727 11418
rect 17762 11384 17796 11418
rect 17831 11384 17865 11418
rect 17900 11384 17934 11418
rect 17969 11384 18003 11418
rect 18038 11384 18072 11418
rect 18107 11384 18141 11418
rect 18176 11384 18210 11418
rect 18245 11384 18279 11418
rect 18314 11384 18348 11418
rect 18383 11384 18417 11418
rect 18452 11384 18486 11418
rect 18521 11384 18555 11418
rect 18590 11384 18624 11418
rect 18659 11384 18693 11418
rect 18728 11384 18762 11418
rect 18797 11384 18831 11418
rect 18866 11384 18900 11418
rect 18935 11384 18969 11418
rect 19004 11384 19038 11418
rect 19073 11384 19107 11418
rect 19142 11384 19176 11418
rect 19211 11384 19245 11418
rect 19280 11384 19314 11418
rect 19349 11384 19383 11418
rect 19418 11384 19452 11418
rect 19487 11384 19521 11418
rect 19556 11384 19590 11418
rect 19625 11384 19659 11418
rect 6770 11296 6804 11330
rect 6839 11296 6873 11330
rect 6908 11296 6942 11330
rect 6977 11296 7011 11330
rect 7046 11296 7080 11330
rect 7115 11296 7149 11330
rect 7184 11296 7218 11330
rect 7253 11296 7287 11330
rect 7322 11296 7356 11330
rect 7391 11296 7425 11330
rect 7460 11296 7494 11330
rect 7529 11296 7563 11330
rect 7598 11296 7632 11330
rect 7667 11296 7701 11330
rect 7736 11296 7770 11330
rect 7805 11296 7839 11330
rect 7874 11296 7908 11330
rect 7943 11296 7977 11330
rect 8012 11296 8046 11330
rect 8081 11296 8115 11330
rect 8150 11296 8184 11330
rect 8219 11296 8253 11330
rect 8288 11296 8322 11330
rect 8357 11296 8391 11330
rect 8426 11296 8460 11330
rect 8495 11296 8529 11330
rect 8564 11296 8598 11330
rect 8633 11296 8667 11330
rect 8702 11296 8736 11330
rect 8771 11296 8805 11330
rect 8840 11296 8874 11330
rect 8909 11296 8943 11330
rect 8978 11296 9012 11330
rect 9046 11296 9080 11330
rect 9114 11296 9148 11330
rect 9182 11296 9216 11330
rect 9250 11296 9284 11330
rect 9318 11296 9352 11330
rect 9386 11296 9420 11330
rect 9454 11296 9488 11330
rect 9522 11296 9556 11330
rect 9590 11296 9624 11330
rect 9658 11296 9692 11330
rect 9726 11296 9760 11330
rect 9794 11296 9828 11330
rect 9862 11296 9896 11330
rect 9930 11296 9964 11330
rect 9998 11296 10032 11330
rect 10066 11296 10100 11330
rect 10134 11296 10168 11330
rect 10202 11296 10236 11330
rect 10270 11296 10304 11330
rect 16319 11316 16353 11350
rect 16388 11316 16422 11350
rect 16457 11316 16491 11350
rect 16526 11316 16560 11350
rect 16594 11316 16628 11350
rect 16662 11316 16696 11350
rect 16730 11316 16764 11350
rect 16798 11316 16832 11350
rect 16866 11316 16900 11350
rect 16934 11316 16968 11350
rect 17002 11316 17036 11350
rect 17070 11316 17104 11350
rect 17138 11316 17172 11350
rect 17206 11316 17240 11350
rect 17274 11316 17308 11350
rect 17342 11316 17376 11350
rect 17410 11316 17444 11350
rect 17478 11316 17512 11350
rect 17546 11316 17580 11350
rect 17614 11316 17648 11350
rect 17682 11316 17716 11350
rect 17750 11316 17784 11350
rect 17818 11316 17852 11350
rect 17886 11316 17920 11350
rect 17954 11316 17988 11350
rect 18022 11316 18056 11350
rect 18090 11316 18124 11350
rect 18158 11316 18192 11350
rect 18226 11316 18260 11350
rect 18294 11316 18328 11350
rect 18362 11316 18396 11350
rect 18430 11316 18464 11350
rect 18498 11316 18532 11350
rect 18566 11316 18600 11350
rect 18634 11316 18668 11350
rect 18702 11316 18736 11350
rect 18770 11316 18804 11350
rect 18838 11316 18872 11350
rect 18906 11316 18940 11350
rect 18974 11316 19008 11350
rect 19042 11316 19076 11350
rect 19110 11316 19144 11350
rect 19178 11316 19212 11350
rect 19246 11316 19280 11350
rect 19314 11316 19348 11350
rect 6770 11224 6804 11258
rect 6839 11224 6873 11258
rect 6908 11224 6942 11258
rect 6977 11224 7011 11258
rect 7046 11224 7080 11258
rect 7115 11224 7149 11258
rect 7184 11224 7218 11258
rect 7253 11224 7287 11258
rect 7322 11224 7356 11258
rect 7391 11224 7425 11258
rect 7460 11224 7494 11258
rect 7529 11224 7563 11258
rect 7598 11224 7632 11258
rect 7667 11224 7701 11258
rect 7736 11224 7770 11258
rect 7805 11224 7839 11258
rect 7874 11224 7908 11258
rect 7943 11224 7977 11258
rect 8012 11224 8046 11258
rect 8081 11224 8115 11258
rect 8150 11224 8184 11258
rect 8219 11224 8253 11258
rect 8288 11224 8322 11258
rect 8357 11224 8391 11258
rect 8426 11224 8460 11258
rect 8495 11224 8529 11258
rect 8564 11224 8598 11258
rect 8633 11224 8667 11258
rect 8702 11224 8736 11258
rect 8771 11224 8805 11258
rect 8840 11224 8874 11258
rect 8909 11224 8943 11258
rect 8978 11224 9012 11258
rect 9046 11224 9080 11258
rect 9114 11224 9148 11258
rect 9182 11224 9216 11258
rect 9250 11224 9284 11258
rect 9318 11224 9352 11258
rect 9386 11224 9420 11258
rect 9454 11224 9488 11258
rect 9522 11224 9556 11258
rect 9590 11224 9624 11258
rect 9658 11224 9692 11258
rect 9726 11224 9760 11258
rect 9794 11224 9828 11258
rect 9862 11224 9896 11258
rect 9930 11224 9964 11258
rect 9998 11224 10032 11258
rect 10066 11224 10100 11258
rect 10134 11224 10168 11258
rect 10202 11224 10236 11258
rect 10270 11224 10304 11258
rect 6770 11152 6804 11186
rect 6839 11152 6873 11186
rect 6908 11152 6942 11186
rect 6977 11152 7011 11186
rect 7046 11152 7080 11186
rect 7115 11152 7149 11186
rect 7184 11152 7218 11186
rect 7253 11152 7287 11186
rect 7322 11152 7356 11186
rect 7391 11152 7425 11186
rect 7460 11152 7494 11186
rect 7529 11152 7563 11186
rect 7598 11152 7632 11186
rect 7667 11152 7701 11186
rect 7736 11152 7770 11186
rect 7805 11152 7839 11186
rect 7874 11152 7908 11186
rect 7943 11152 7977 11186
rect 8012 11152 8046 11186
rect 8081 11152 8115 11186
rect 8150 11152 8184 11186
rect 8219 11152 8253 11186
rect 8288 11152 8322 11186
rect 8357 11152 8391 11186
rect 8426 11152 8460 11186
rect 8495 11152 8529 11186
rect 8564 11152 8598 11186
rect 8633 11152 8667 11186
rect 8702 11152 8736 11186
rect 8771 11152 8805 11186
rect 8840 11152 8874 11186
rect 8909 11152 8943 11186
rect 8978 11152 9012 11186
rect 9046 11152 9080 11186
rect 9114 11152 9148 11186
rect 9182 11152 9216 11186
rect 9250 11152 9284 11186
rect 9318 11152 9352 11186
rect 9386 11152 9420 11186
rect 9454 11152 9488 11186
rect 9522 11152 9556 11186
rect 9590 11152 9624 11186
rect 9658 11152 9692 11186
rect 9726 11152 9760 11186
rect 9794 11152 9828 11186
rect 9862 11152 9896 11186
rect 9930 11152 9964 11186
rect 9998 11152 10032 11186
rect 10066 11152 10100 11186
rect 10134 11152 10168 11186
rect 10202 11152 10236 11186
rect 10270 11152 10304 11186
rect 16319 11244 16353 11278
rect 16388 11244 16422 11278
rect 16457 11244 16491 11278
rect 16526 11244 16560 11278
rect 16594 11244 16628 11278
rect 16662 11244 16696 11278
rect 16730 11244 16764 11278
rect 16798 11244 16832 11278
rect 16866 11244 16900 11278
rect 16934 11244 16968 11278
rect 17002 11244 17036 11278
rect 17070 11244 17104 11278
rect 17138 11244 17172 11278
rect 17206 11244 17240 11278
rect 17274 11244 17308 11278
rect 17342 11244 17376 11278
rect 17410 11244 17444 11278
rect 17478 11244 17512 11278
rect 17546 11244 17580 11278
rect 17614 11244 17648 11278
rect 17682 11244 17716 11278
rect 17750 11244 17784 11278
rect 17818 11244 17852 11278
rect 17886 11244 17920 11278
rect 17954 11244 17988 11278
rect 18022 11244 18056 11278
rect 18090 11244 18124 11278
rect 18158 11244 18192 11278
rect 18226 11244 18260 11278
rect 18294 11244 18328 11278
rect 18362 11244 18396 11278
rect 18430 11244 18464 11278
rect 18498 11244 18532 11278
rect 18566 11244 18600 11278
rect 18634 11244 18668 11278
rect 18702 11244 18736 11278
rect 18770 11244 18804 11278
rect 18838 11244 18872 11278
rect 18906 11244 18940 11278
rect 18974 11244 19008 11278
rect 19042 11244 19076 11278
rect 19110 11244 19144 11278
rect 19178 11244 19212 11278
rect 19246 11244 19280 11278
rect 19314 11244 19348 11278
rect 25124 11321 25158 11355
rect 25196 11321 25230 11355
rect 25268 11321 25302 11355
rect 25340 11321 25374 11355
rect 25412 11321 25446 11355
rect 25484 11321 25518 11355
rect 25556 11321 25590 11355
rect 25627 11321 25661 11355
rect 25698 11321 25732 11355
rect 25769 11321 25803 11355
rect 25840 11321 25874 11355
rect 25911 11321 25945 11355
rect 25982 11321 26016 11355
rect 26053 11321 26087 11355
rect 26124 11321 26158 11355
rect 26195 11321 26229 11355
rect 25124 11253 25158 11287
rect 25196 11253 25230 11287
rect 25268 11253 25302 11287
rect 25340 11253 25374 11287
rect 25412 11253 25446 11287
rect 25484 11253 25518 11287
rect 25556 11253 25590 11287
rect 25627 11253 25661 11287
rect 25698 11253 25732 11287
rect 25769 11253 25803 11287
rect 25840 11253 25874 11287
rect 25911 11253 25945 11287
rect 25982 11253 26016 11287
rect 26053 11253 26087 11287
rect 26124 11253 26158 11287
rect 26195 11253 26229 11287
rect 16319 11172 16353 11206
rect 16388 11172 16422 11206
rect 16457 11172 16491 11206
rect 16526 11172 16560 11206
rect 16594 11172 16628 11206
rect 16662 11172 16696 11206
rect 16730 11172 16764 11206
rect 16798 11172 16832 11206
rect 16866 11172 16900 11206
rect 16934 11172 16968 11206
rect 17002 11172 17036 11206
rect 17070 11172 17104 11206
rect 17138 11172 17172 11206
rect 17206 11172 17240 11206
rect 17274 11172 17308 11206
rect 17342 11172 17376 11206
rect 17410 11172 17444 11206
rect 17478 11172 17512 11206
rect 17546 11172 17580 11206
rect 17614 11172 17648 11206
rect 17682 11172 17716 11206
rect 17750 11172 17784 11206
rect 17818 11172 17852 11206
rect 17886 11172 17920 11206
rect 17954 11172 17988 11206
rect 18022 11172 18056 11206
rect 18090 11172 18124 11206
rect 18158 11172 18192 11206
rect 18226 11172 18260 11206
rect 18294 11172 18328 11206
rect 18362 11172 18396 11206
rect 18430 11172 18464 11206
rect 18498 11172 18532 11206
rect 18566 11172 18600 11206
rect 18634 11172 18668 11206
rect 18702 11172 18736 11206
rect 18770 11172 18804 11206
rect 18838 11172 18872 11206
rect 18906 11172 18940 11206
rect 18974 11172 19008 11206
rect 19042 11172 19076 11206
rect 19110 11172 19144 11206
rect 19178 11172 19212 11206
rect 19246 11172 19280 11206
rect 19314 11172 19348 11206
rect 6751 11038 6785 11072
rect 6827 11038 6861 11072
rect 6903 11038 6937 11072
rect 6979 11038 7013 11072
rect 7055 11038 7089 11072
rect 7131 11038 7165 11072
rect 7207 11038 7241 11072
rect 6751 10970 6785 11004
rect 6827 10970 6861 11004
rect 6903 10970 6937 11004
rect 6979 10970 7013 11004
rect 7055 10970 7089 11004
rect 7131 10970 7165 11004
rect 7207 10970 7241 11004
rect 6751 10902 6785 10936
rect 6827 10902 6861 10936
rect 6903 10902 6937 10936
rect 6979 10902 7013 10936
rect 7055 10902 7089 10936
rect 7131 10902 7165 10936
rect 7207 10902 7241 10936
rect 6751 10834 6785 10868
rect 6827 10834 6861 10868
rect 6903 10834 6937 10868
rect 6979 10834 7013 10868
rect 7055 10834 7089 10868
rect 7131 10834 7165 10868
rect 7207 10834 7241 10868
rect 6751 10766 6785 10800
rect 6827 10766 6861 10800
rect 6903 10766 6937 10800
rect 6979 10766 7013 10800
rect 7055 10766 7089 10800
rect 7131 10766 7165 10800
rect 7207 10766 7241 10800
rect 6751 10698 6785 10732
rect 6827 10698 6861 10732
rect 6903 10698 6937 10732
rect 6979 10698 7013 10732
rect 7055 10698 7089 10732
rect 7131 10698 7165 10732
rect 7207 10698 7241 10732
rect 6751 10630 6785 10664
rect 6827 10630 6861 10664
rect 6903 10630 6937 10664
rect 6979 10630 7013 10664
rect 7055 10630 7089 10664
rect 7131 10630 7165 10664
rect 7207 10630 7241 10664
rect 6751 10562 6785 10596
rect 6827 10562 6861 10596
rect 6903 10562 6937 10596
rect 6979 10562 7013 10596
rect 7055 10562 7089 10596
rect 7131 10562 7165 10596
rect 7207 10562 7241 10596
rect 6751 10494 6785 10528
rect 6827 10494 6861 10528
rect 6903 10494 6937 10528
rect 6979 10494 7013 10528
rect 7055 10494 7089 10528
rect 7131 10494 7165 10528
rect 7207 10494 7241 10528
rect 6751 10426 6785 10460
rect 6827 10426 6861 10460
rect 6903 10426 6937 10460
rect 6979 10426 7013 10460
rect 7055 10426 7089 10460
rect 7131 10426 7165 10460
rect 7207 10426 7241 10460
rect 6751 10358 6785 10392
rect 6827 10358 6861 10392
rect 6903 10358 6937 10392
rect 6979 10358 7013 10392
rect 7055 10358 7089 10392
rect 7131 10358 7165 10392
rect 7207 10358 7241 10392
rect 6751 10290 6785 10324
rect 6827 10290 6861 10324
rect 6903 10290 6937 10324
rect 6979 10290 7013 10324
rect 7055 10290 7089 10324
rect 7131 10290 7165 10324
rect 7207 10290 7241 10324
rect 6751 10222 6785 10256
rect 6827 10222 6861 10256
rect 6903 10222 6937 10256
rect 6979 10222 7013 10256
rect 7055 10222 7089 10256
rect 7131 10222 7165 10256
rect 7207 10222 7241 10256
rect 6751 10154 6785 10188
rect 6827 10154 6861 10188
rect 6903 10154 6937 10188
rect 6979 10154 7013 10188
rect 7055 10154 7089 10188
rect 7131 10154 7165 10188
rect 7207 10154 7241 10188
rect 6751 10086 6785 10120
rect 6827 10086 6861 10120
rect 6903 10086 6937 10120
rect 6979 10086 7013 10120
rect 7055 10086 7089 10120
rect 7131 10086 7165 10120
rect 7207 10086 7241 10120
rect 6751 10018 6785 10052
rect 6827 10018 6861 10052
rect 6903 10018 6937 10052
rect 6979 10018 7013 10052
rect 7055 10018 7089 10052
rect 7131 10018 7165 10052
rect 7207 10018 7241 10052
rect 6751 9950 6785 9984
rect 6827 9950 6861 9984
rect 6903 9950 6937 9984
rect 6979 9950 7013 9984
rect 7055 9950 7089 9984
rect 7131 9950 7165 9984
rect 7207 9950 7241 9984
rect 6751 9882 6785 9916
rect 6827 9882 6861 9916
rect 6903 9882 6937 9916
rect 6979 9882 7013 9916
rect 7055 9882 7089 9916
rect 7131 9882 7165 9916
rect 7207 9882 7241 9916
rect 6751 9814 6785 9848
rect 6827 9814 6861 9848
rect 6903 9814 6937 9848
rect 6979 9814 7013 9848
rect 7055 9814 7089 9848
rect 7131 9814 7165 9848
rect 7207 9814 7241 9848
rect 6751 9746 6785 9780
rect 6827 9746 6861 9780
rect 6903 9746 6937 9780
rect 6979 9746 7013 9780
rect 7055 9746 7089 9780
rect 7131 9746 7165 9780
rect 7207 9746 7241 9780
rect 6751 9678 6785 9712
rect 6827 9678 6861 9712
rect 6903 9678 6937 9712
rect 6979 9678 7013 9712
rect 7055 9678 7089 9712
rect 7131 9678 7165 9712
rect 7207 9678 7241 9712
rect 6751 9610 6785 9644
rect 6827 9610 6861 9644
rect 6903 9610 6937 9644
rect 6979 9610 7013 9644
rect 7055 9610 7089 9644
rect 7131 9610 7165 9644
rect 7207 9610 7241 9644
rect 10049 10290 10219 11072
rect 16319 11100 16353 11134
rect 16388 11100 16422 11134
rect 16457 11100 16491 11134
rect 16526 11100 16560 11134
rect 16594 11100 16628 11134
rect 16662 11100 16696 11134
rect 16730 11100 16764 11134
rect 16798 11100 16832 11134
rect 16866 11100 16900 11134
rect 16934 11100 16968 11134
rect 17002 11100 17036 11134
rect 17070 11100 17104 11134
rect 17138 11100 17172 11134
rect 17206 11100 17240 11134
rect 17274 11100 17308 11134
rect 17342 11100 17376 11134
rect 17410 11100 17444 11134
rect 17478 11100 17512 11134
rect 17546 11100 17580 11134
rect 17614 11100 17648 11134
rect 17682 11100 17716 11134
rect 17750 11100 17784 11134
rect 17818 11100 17852 11134
rect 17886 11100 17920 11134
rect 17954 11100 17988 11134
rect 18022 11100 18056 11134
rect 18090 11100 18124 11134
rect 18158 11100 18192 11134
rect 18226 11100 18260 11134
rect 18294 11100 18328 11134
rect 18362 11100 18396 11134
rect 18430 11100 18464 11134
rect 18498 11100 18532 11134
rect 18566 11100 18600 11134
rect 18634 11100 18668 11134
rect 18702 11100 18736 11134
rect 18770 11100 18804 11134
rect 18838 11100 18872 11134
rect 18906 11100 18940 11134
rect 18974 11100 19008 11134
rect 19042 11100 19076 11134
rect 19110 11100 19144 11134
rect 19178 11100 19212 11134
rect 19246 11100 19280 11134
rect 19314 11100 19348 11134
rect 10049 10221 10083 10255
rect 10117 10221 10151 10255
rect 10185 10221 10219 10255
rect 10049 10152 10083 10186
rect 10117 10152 10151 10186
rect 10185 10152 10219 10186
rect 10049 10083 10083 10117
rect 10117 10083 10151 10117
rect 10185 10083 10219 10117
rect 10049 10014 10083 10048
rect 10117 10014 10151 10048
rect 10185 10014 10219 10048
rect 10049 9945 10083 9979
rect 10117 9945 10151 9979
rect 10185 9945 10219 9979
rect 10049 9876 10083 9910
rect 10117 9876 10151 9910
rect 10185 9876 10219 9910
rect 10049 9807 10083 9841
rect 10117 9807 10151 9841
rect 10185 9807 10219 9841
rect 10049 9738 10083 9772
rect 10117 9738 10151 9772
rect 10185 9738 10219 9772
rect 10049 9669 10083 9703
rect 10117 9669 10151 9703
rect 10185 9669 10219 9703
rect 10049 9600 10083 9634
rect 10117 9600 10151 9634
rect 10185 9600 10219 9634
rect 6751 9542 6785 9576
rect 6827 9542 6861 9576
rect 6903 9542 6937 9576
rect 6979 9542 7013 9576
rect 7055 9542 7089 9576
rect 7131 9542 7165 9576
rect 7207 9542 7241 9576
rect 7332 9554 7366 9588
rect 7401 9554 7435 9588
rect 7470 9554 7504 9588
rect 7539 9554 7573 9588
rect 7608 9554 7642 9588
rect 7677 9554 7711 9588
rect 7746 9554 7780 9588
rect 7815 9554 7849 9588
rect 7884 9554 7918 9588
rect 7953 9554 7987 9588
rect 8022 9554 8056 9588
rect 8091 9554 8125 9588
rect 8160 9554 8194 9588
rect 8229 9554 8263 9588
rect 8297 9554 8331 9588
rect 8365 9554 8399 9588
rect 8433 9554 8467 9588
rect 8501 9554 8535 9588
rect 8569 9554 8603 9588
rect 8637 9554 8671 9588
rect 8705 9554 8739 9588
rect 8773 9554 8807 9588
rect 8841 9554 8875 9588
rect 8909 9554 8943 9588
rect 8977 9554 9011 9588
rect 9045 9554 9079 9588
rect 9113 9554 9147 9588
rect 9181 9554 9215 9588
rect 9249 9554 9283 9588
rect 9317 9554 9351 9588
rect 9385 9554 9419 9588
rect 9453 9554 9487 9588
rect 9521 9554 9555 9588
rect 9589 9554 9623 9588
rect 9657 9554 9691 9588
rect 9725 9554 9759 9588
rect 9793 9554 9827 9588
rect 9861 9554 9895 9588
rect 9929 9554 9963 9588
rect 10049 9531 10083 9565
rect 10117 9531 10151 9565
rect 10185 9531 10219 9565
rect 26277 10336 26311 10370
rect 26348 10336 26382 10370
rect 26419 10336 26453 10370
rect 26490 10336 26524 10370
rect 26561 10336 26595 10370
rect 26632 10336 26666 10370
rect 26703 10336 26737 10370
rect 26774 10336 26808 10370
rect 26845 10336 26879 10370
rect 26916 10336 26950 10370
rect 26986 10336 27020 10370
rect 27056 10336 27090 10370
rect 27126 10336 27160 10370
rect 27196 10336 27230 10370
rect 27266 10336 27300 10370
rect 27336 10336 27370 10370
rect 27406 10336 27440 10370
rect 27547 10312 27581 10346
rect 27615 10312 27649 10346
rect 27683 10312 27717 10346
rect 27751 10312 27785 10346
rect 27819 10312 27853 10346
rect 26277 10268 26311 10302
rect 26348 10268 26382 10302
rect 26419 10268 26453 10302
rect 26490 10268 26524 10302
rect 26561 10268 26595 10302
rect 26632 10268 26666 10302
rect 26703 10268 26737 10302
rect 26774 10268 26808 10302
rect 26845 10268 26879 10302
rect 26916 10268 26950 10302
rect 26986 10268 27020 10302
rect 27056 10268 27090 10302
rect 27126 10268 27160 10302
rect 27196 10268 27230 10302
rect 27266 10268 27300 10302
rect 27336 10268 27370 10302
rect 27406 10268 27440 10302
rect 27547 10243 27581 10277
rect 27615 10243 27649 10277
rect 27683 10243 27717 10277
rect 27751 10243 27785 10277
rect 27819 10243 27853 10277
rect 26277 10200 26311 10234
rect 26348 10200 26382 10234
rect 26419 10200 26453 10234
rect 26490 10200 26524 10234
rect 26561 10200 26595 10234
rect 26632 10200 26666 10234
rect 26703 10200 26737 10234
rect 26774 10200 26808 10234
rect 26845 10200 26879 10234
rect 26916 10200 26950 10234
rect 26986 10200 27020 10234
rect 27056 10200 27090 10234
rect 27126 10200 27160 10234
rect 27196 10200 27230 10234
rect 27266 10200 27300 10234
rect 27336 10200 27370 10234
rect 27406 10200 27440 10234
rect 27547 10174 27581 10208
rect 27615 10174 27649 10208
rect 27683 10174 27717 10208
rect 27751 10174 27785 10208
rect 27819 10174 27853 10208
rect 26277 10132 26311 10166
rect 26348 10132 26382 10166
rect 26419 10132 26453 10166
rect 26490 10132 26524 10166
rect 26561 10132 26595 10166
rect 26632 10132 26666 10166
rect 26703 10132 26737 10166
rect 26774 10132 26808 10166
rect 26845 10132 26879 10166
rect 26916 10132 26950 10166
rect 26986 10132 27020 10166
rect 27056 10132 27090 10166
rect 27126 10132 27160 10166
rect 27196 10132 27230 10166
rect 27266 10132 27300 10166
rect 27336 10132 27370 10166
rect 27406 10132 27440 10166
rect 27547 10105 27581 10139
rect 27615 10105 27649 10139
rect 27683 10105 27717 10139
rect 27751 10105 27785 10139
rect 27819 10105 27853 10139
rect 26277 10064 26311 10098
rect 26348 10064 26382 10098
rect 26419 10064 26453 10098
rect 26490 10064 26524 10098
rect 26561 10064 26595 10098
rect 26632 10064 26666 10098
rect 26703 10064 26737 10098
rect 26774 10064 26808 10098
rect 26845 10064 26879 10098
rect 26916 10064 26950 10098
rect 26986 10064 27020 10098
rect 27056 10064 27090 10098
rect 27126 10064 27160 10098
rect 27196 10064 27230 10098
rect 27266 10064 27300 10098
rect 27336 10064 27370 10098
rect 27406 10064 27440 10098
rect 27547 10036 27581 10070
rect 27615 10036 27649 10070
rect 27683 10036 27717 10070
rect 27751 10036 27785 10070
rect 27819 10036 27853 10070
rect 26277 9996 26311 10030
rect 26348 9996 26382 10030
rect 26419 9996 26453 10030
rect 26490 9996 26524 10030
rect 26561 9996 26595 10030
rect 26632 9996 26666 10030
rect 26703 9996 26737 10030
rect 26774 9996 26808 10030
rect 26845 9996 26879 10030
rect 26916 9996 26950 10030
rect 26986 9996 27020 10030
rect 27056 9996 27090 10030
rect 27126 9996 27160 10030
rect 27196 9996 27230 10030
rect 27266 9996 27300 10030
rect 27336 9996 27370 10030
rect 27406 9996 27440 10030
rect 27547 9967 27581 10001
rect 27615 9967 27649 10001
rect 27683 9967 27717 10001
rect 27751 9967 27785 10001
rect 27819 9967 27853 10001
rect 26277 9928 26311 9962
rect 26348 9928 26382 9962
rect 26419 9928 26453 9962
rect 26490 9928 26524 9962
rect 26561 9928 26595 9962
rect 26632 9928 26666 9962
rect 26703 9928 26737 9962
rect 26774 9928 26808 9962
rect 26845 9928 26879 9962
rect 26916 9928 26950 9962
rect 26986 9928 27020 9962
rect 27056 9928 27090 9962
rect 27126 9928 27160 9962
rect 27196 9928 27230 9962
rect 27266 9928 27300 9962
rect 27336 9928 27370 9962
rect 27406 9928 27440 9962
rect 27547 9898 27581 9932
rect 27615 9898 27649 9932
rect 27683 9898 27717 9932
rect 27751 9898 27785 9932
rect 27819 9898 27853 9932
rect 26277 9860 26311 9894
rect 26348 9860 26382 9894
rect 26419 9860 26453 9894
rect 26490 9860 26524 9894
rect 26561 9860 26595 9894
rect 26632 9860 26666 9894
rect 26703 9860 26737 9894
rect 26774 9860 26808 9894
rect 26845 9860 26879 9894
rect 26916 9860 26950 9894
rect 26986 9860 27020 9894
rect 27056 9860 27090 9894
rect 27126 9860 27160 9894
rect 27196 9860 27230 9894
rect 27266 9860 27300 9894
rect 27336 9860 27370 9894
rect 27406 9860 27440 9894
rect 27547 9829 27581 9863
rect 27615 9829 27649 9863
rect 27683 9829 27717 9863
rect 27751 9829 27785 9863
rect 27819 9829 27853 9863
rect 27547 9760 27581 9794
rect 27615 9760 27649 9794
rect 27683 9760 27717 9794
rect 27751 9760 27785 9794
rect 27819 9760 27853 9794
rect 27547 9690 27581 9724
rect 27615 9690 27649 9724
rect 27683 9690 27717 9724
rect 27751 9690 27785 9724
rect 27819 9690 27853 9724
rect 27547 9620 27581 9654
rect 27615 9620 27649 9654
rect 27683 9620 27717 9654
rect 27751 9620 27785 9654
rect 27819 9620 27853 9654
rect 27547 9550 27581 9584
rect 27615 9550 27649 9584
rect 27683 9550 27717 9584
rect 27751 9550 27785 9584
rect 27819 9550 27853 9584
rect 6751 9474 6785 9508
rect 6827 9474 6861 9508
rect 6903 9474 6937 9508
rect 6979 9474 7013 9508
rect 7055 9474 7089 9508
rect 7131 9474 7165 9508
rect 7207 9474 7241 9508
rect 7332 9462 7366 9496
rect 7401 9462 7435 9496
rect 7470 9462 7504 9496
rect 7539 9462 7573 9496
rect 7608 9462 7642 9496
rect 7677 9462 7711 9496
rect 7746 9462 7780 9496
rect 7815 9462 7849 9496
rect 7884 9462 7918 9496
rect 7953 9462 7987 9496
rect 8022 9462 8056 9496
rect 8091 9462 8125 9496
rect 8160 9462 8194 9496
rect 8229 9462 8263 9496
rect 8297 9462 8331 9496
rect 8365 9462 8399 9496
rect 8433 9462 8467 9496
rect 8501 9462 8535 9496
rect 8569 9462 8603 9496
rect 8637 9462 8671 9496
rect 8705 9462 8739 9496
rect 8773 9462 8807 9496
rect 8841 9462 8875 9496
rect 8909 9462 8943 9496
rect 8977 9462 9011 9496
rect 9045 9462 9079 9496
rect 9113 9462 9147 9496
rect 9181 9462 9215 9496
rect 9249 9462 9283 9496
rect 9317 9462 9351 9496
rect 9385 9462 9419 9496
rect 9453 9462 9487 9496
rect 9521 9462 9555 9496
rect 9589 9462 9623 9496
rect 9657 9462 9691 9496
rect 9725 9462 9759 9496
rect 9793 9462 9827 9496
rect 9861 9462 9895 9496
rect 9929 9462 9963 9496
rect 10049 9462 10083 9496
rect 10117 9462 10151 9496
rect 10185 9462 10219 9496
rect 10305 9493 10339 9527
rect 10405 9493 10439 9527
rect 10505 9493 10539 9527
rect 6751 9406 6785 9440
rect 6827 9406 6861 9440
rect 6903 9406 6937 9440
rect 6979 9406 7013 9440
rect 7055 9406 7089 9440
rect 7131 9406 7165 9440
rect 7207 9406 7241 9440
rect 6751 9338 6785 9372
rect 6827 9338 6861 9372
rect 6903 9338 6937 9372
rect 6979 9338 7013 9372
rect 7055 9338 7089 9372
rect 7131 9338 7165 9372
rect 7207 9338 7241 9372
rect 7332 9370 7366 9404
rect 7401 9370 7435 9404
rect 7470 9370 7504 9404
rect 7539 9370 7573 9404
rect 7608 9370 7642 9404
rect 7677 9370 7711 9404
rect 7746 9370 7780 9404
rect 7815 9370 7849 9404
rect 7884 9370 7918 9404
rect 7953 9370 7987 9404
rect 8022 9370 8056 9404
rect 8091 9370 8125 9404
rect 8160 9370 8194 9404
rect 8229 9370 8263 9404
rect 8297 9370 8331 9404
rect 8365 9370 8399 9404
rect 8433 9370 8467 9404
rect 8501 9370 8535 9404
rect 8569 9370 8603 9404
rect 8637 9370 8671 9404
rect 8705 9370 8739 9404
rect 8773 9370 8807 9404
rect 8841 9370 8875 9404
rect 8909 9370 8943 9404
rect 8977 9370 9011 9404
rect 9045 9370 9079 9404
rect 9113 9370 9147 9404
rect 9181 9370 9215 9404
rect 9249 9370 9283 9404
rect 9317 9370 9351 9404
rect 9385 9370 9419 9404
rect 9453 9370 9487 9404
rect 9521 9370 9555 9404
rect 9589 9370 9623 9404
rect 9657 9370 9691 9404
rect 9725 9370 9759 9404
rect 9793 9370 9827 9404
rect 9861 9370 9895 9404
rect 9929 9370 9963 9404
rect 10049 9393 10083 9427
rect 10117 9393 10151 9427
rect 10185 9393 10219 9427
rect 10573 9421 10607 9455
rect 27547 9480 27581 9514
rect 27615 9480 27649 9514
rect 27683 9480 27717 9514
rect 27751 9480 27785 9514
rect 27819 9480 27853 9514
rect 10305 9369 10339 9403
rect 10377 9369 10411 9403
rect 10449 9369 10483 9403
rect 6751 9270 6785 9304
rect 6827 9270 6861 9304
rect 6903 9270 6937 9304
rect 6979 9270 7013 9304
rect 7055 9270 7089 9304
rect 7131 9270 7165 9304
rect 7207 9270 7241 9304
rect 6751 9202 6785 9236
rect 6827 9202 6861 9236
rect 6903 9202 6937 9236
rect 6979 9202 7013 9236
rect 7055 9202 7089 9236
rect 7131 9202 7165 9236
rect 7207 9202 7241 9236
rect 6751 9134 6785 9168
rect 6827 9134 6861 9168
rect 6903 9134 6937 9168
rect 6979 9134 7013 9168
rect 7055 9134 7089 9168
rect 7131 9134 7165 9168
rect 7207 9134 7241 9168
rect 6751 9066 6785 9100
rect 6827 9066 6861 9100
rect 6903 9066 6937 9100
rect 6979 9066 7013 9100
rect 7055 9066 7089 9100
rect 7131 9066 7165 9100
rect 7207 9066 7241 9100
rect 6751 8998 6785 9032
rect 6827 8998 6861 9032
rect 6903 8998 6937 9032
rect 6979 8998 7013 9032
rect 7055 8998 7089 9032
rect 7131 8998 7165 9032
rect 7207 8998 7241 9032
rect 6751 8930 6785 8964
rect 6827 8930 6861 8964
rect 6903 8930 6937 8964
rect 6979 8930 7013 8964
rect 7055 8930 7089 8964
rect 7131 8930 7165 8964
rect 7207 8930 7241 8964
rect 6751 8862 6785 8896
rect 6827 8862 6861 8896
rect 6903 8862 6937 8896
rect 6979 8862 7013 8896
rect 7055 8862 7089 8896
rect 7131 8862 7165 8896
rect 7207 8862 7241 8896
rect 192 8822 226 8856
rect 262 8822 296 8856
rect 332 8822 366 8856
rect 402 8822 436 8856
rect 472 8822 506 8856
rect 542 8822 576 8856
rect 612 8822 646 8856
rect 682 8822 716 8856
rect 752 8822 786 8856
rect 822 8822 856 8856
rect 891 8822 925 8856
rect 960 8822 994 8856
rect 1029 8822 1063 8856
rect 1098 8822 1132 8856
rect 1167 8822 1201 8856
rect 1236 8822 1270 8856
rect 1305 8822 1339 8856
rect 1374 8822 1408 8856
rect 1443 8822 1477 8856
rect 1512 8822 1546 8856
rect 1581 8822 1615 8856
rect 1650 8822 1684 8856
rect 1719 8822 1753 8856
rect 1788 8822 1822 8856
rect 192 8748 226 8782
rect 262 8748 296 8782
rect 332 8748 366 8782
rect 402 8748 436 8782
rect 472 8748 506 8782
rect 542 8748 576 8782
rect 612 8748 646 8782
rect 682 8748 716 8782
rect 752 8748 786 8782
rect 822 8748 856 8782
rect 891 8748 925 8782
rect 960 8748 994 8782
rect 1029 8748 1063 8782
rect 1098 8748 1132 8782
rect 1167 8748 1201 8782
rect 1236 8748 1270 8782
rect 1305 8748 1339 8782
rect 1374 8748 1408 8782
rect 1443 8748 1477 8782
rect 1512 8748 1546 8782
rect 1581 8748 1615 8782
rect 1650 8748 1684 8782
rect 1719 8748 1753 8782
rect 1788 8748 1822 8782
rect 192 8674 226 8708
rect 262 8674 296 8708
rect 332 8674 366 8708
rect 402 8674 436 8708
rect 472 8674 506 8708
rect 542 8674 576 8708
rect 612 8674 646 8708
rect 682 8674 716 8708
rect 752 8674 786 8708
rect 822 8674 856 8708
rect 891 8674 925 8708
rect 960 8674 994 8708
rect 1029 8674 1063 8708
rect 1098 8674 1132 8708
rect 1167 8674 1201 8708
rect 1236 8674 1270 8708
rect 1305 8674 1339 8708
rect 1374 8674 1408 8708
rect 1443 8674 1477 8708
rect 1512 8674 1546 8708
rect 1581 8674 1615 8708
rect 1650 8674 1684 8708
rect 1719 8674 1753 8708
rect 1788 8674 1822 8708
rect 192 8600 226 8634
rect 262 8600 296 8634
rect 332 8600 366 8634
rect 402 8600 436 8634
rect 472 8600 506 8634
rect 542 8600 576 8634
rect 612 8600 646 8634
rect 682 8600 716 8634
rect 752 8600 786 8634
rect 822 8600 856 8634
rect 891 8600 925 8634
rect 960 8600 994 8634
rect 1029 8600 1063 8634
rect 1098 8600 1132 8634
rect 1167 8600 1201 8634
rect 1236 8600 1270 8634
rect 1305 8600 1339 8634
rect 1374 8600 1408 8634
rect 1443 8600 1477 8634
rect 1512 8600 1546 8634
rect 1581 8600 1615 8634
rect 1650 8600 1684 8634
rect 1719 8600 1753 8634
rect 1788 8600 1822 8634
rect 192 8526 226 8560
rect 262 8526 296 8560
rect 332 8526 366 8560
rect 402 8526 436 8560
rect 472 8526 506 8560
rect 542 8526 576 8560
rect 612 8526 646 8560
rect 682 8526 716 8560
rect 752 8526 786 8560
rect 822 8526 856 8560
rect 891 8526 925 8560
rect 960 8526 994 8560
rect 1029 8526 1063 8560
rect 1098 8526 1132 8560
rect 1167 8526 1201 8560
rect 1236 8526 1270 8560
rect 1305 8526 1339 8560
rect 1374 8526 1408 8560
rect 1443 8526 1477 8560
rect 1512 8526 1546 8560
rect 1581 8526 1615 8560
rect 1650 8526 1684 8560
rect 1719 8526 1753 8560
rect 1788 8526 1822 8560
rect 6751 8794 6785 8828
rect 6827 8794 6861 8828
rect 6903 8794 6937 8828
rect 6979 8794 7013 8828
rect 7055 8794 7089 8828
rect 7131 8794 7165 8828
rect 7207 8794 7241 8828
rect 6751 8726 6785 8760
rect 6827 8726 6861 8760
rect 6903 8726 6937 8760
rect 6979 8726 7013 8760
rect 7055 8726 7089 8760
rect 7131 8726 7165 8760
rect 7207 8726 7241 8760
rect 6751 8658 6785 8692
rect 6827 8658 6861 8692
rect 6903 8658 6937 8692
rect 6979 8658 7013 8692
rect 7055 8658 7089 8692
rect 7131 8658 7165 8692
rect 7207 8658 7241 8692
rect 6751 8590 6785 8624
rect 6827 8590 6861 8624
rect 6903 8590 6937 8624
rect 6979 8590 7013 8624
rect 7055 8590 7089 8624
rect 7131 8590 7165 8624
rect 7207 8590 7241 8624
rect 6751 8521 6785 8555
rect 6827 8521 6861 8555
rect 6903 8521 6937 8555
rect 6979 8521 7013 8555
rect 7055 8521 7089 8555
rect 7131 8521 7165 8555
rect 7207 8521 7241 8555
rect 10573 9349 10607 9383
rect 10449 9301 10483 9335
rect 10573 9277 10607 9311
rect 10449 9233 10483 9267
rect 10573 9205 10607 9239
rect 10449 9165 10483 9199
rect 10573 9133 10607 9167
rect 10449 9097 10483 9131
rect 10449 9029 10483 9063
rect 10573 9061 10607 9095
rect 10449 8961 10483 8995
rect 10573 8989 10607 9023
rect 23879 9397 23913 9431
rect 24010 9397 24044 9431
rect 23879 9317 23913 9351
rect 24010 9317 24044 9351
rect 23879 9237 23913 9271
rect 24010 9237 24044 9271
rect 23879 9157 23913 9191
rect 24010 9157 24044 9191
rect 23879 9077 23913 9111
rect 24010 9077 24044 9111
rect 23659 8972 23693 9006
rect 23728 8972 23762 9006
rect 23797 8972 23831 9006
rect 23879 8997 23913 9031
rect 24010 8997 24044 9031
rect 10449 8893 10483 8927
rect 10573 8916 10607 8950
rect 10449 8825 10483 8859
rect 10573 8843 10607 8877
rect 10449 8757 10483 8791
rect 10573 8770 10607 8804
rect 10449 8689 10483 8723
rect 10573 8697 10607 8731
rect 10449 8620 10483 8654
rect 10573 8624 10607 8658
rect 10449 8551 10483 8585
rect 10573 8551 10607 8585
rect 20808 8905 20842 8939
rect 20883 8905 20917 8939
rect 20958 8905 20992 8939
rect 21033 8905 21067 8939
rect 21108 8905 21142 8939
rect 21183 8905 21217 8939
rect 21258 8905 21292 8939
rect 21332 8905 21366 8939
rect 21406 8905 21440 8939
rect 21480 8905 21514 8939
rect 23870 8908 23904 8942
rect 23940 8908 23974 8942
rect 24010 8908 24044 8942
rect 27547 9410 27581 9444
rect 27615 9410 27649 9444
rect 27683 9410 27717 9444
rect 27751 9410 27785 9444
rect 27819 9410 27853 9444
rect 27547 9340 27581 9374
rect 27615 9340 27649 9374
rect 27683 9340 27717 9374
rect 27751 9340 27785 9374
rect 27819 9340 27853 9374
rect 27547 9270 27581 9304
rect 27615 9270 27649 9304
rect 27683 9270 27717 9304
rect 27751 9270 27785 9304
rect 27819 9270 27853 9304
rect 27547 9200 27581 9234
rect 27615 9200 27649 9234
rect 27683 9200 27717 9234
rect 27751 9200 27785 9234
rect 27819 9200 27853 9234
rect 27547 9130 27581 9164
rect 27615 9130 27649 9164
rect 27683 9130 27717 9164
rect 27751 9130 27785 9164
rect 27819 9130 27853 9164
rect 27547 9060 27581 9094
rect 27615 9060 27649 9094
rect 27683 9060 27717 9094
rect 27751 9060 27785 9094
rect 27819 9060 27853 9094
rect 27547 8990 27581 9024
rect 27615 8990 27649 9024
rect 27683 8990 27717 9024
rect 27751 8990 27785 9024
rect 27819 8990 27853 9024
rect 27547 8920 27581 8954
rect 27615 8920 27649 8954
rect 27683 8920 27717 8954
rect 27751 8920 27785 8954
rect 27819 8920 27853 8954
rect 21572 8874 21606 8908
rect 21648 8874 21682 8908
rect 21724 8874 21758 8908
rect 21800 8874 21834 8908
rect 21876 8874 21910 8908
rect 21952 8874 21986 8908
rect 22027 8874 22061 8908
rect 22102 8874 22136 8908
rect 20808 8837 20842 8871
rect 20883 8837 20917 8871
rect 20958 8837 20992 8871
rect 21033 8837 21067 8871
rect 21108 8837 21142 8871
rect 21183 8837 21217 8871
rect 21258 8837 21292 8871
rect 21332 8837 21366 8871
rect 21406 8837 21440 8871
rect 21480 8837 21514 8871
rect 22194 8856 22228 8890
rect 22269 8856 22303 8890
rect 22344 8856 22378 8890
rect 22419 8856 22453 8890
rect 22494 8856 22528 8890
rect 22569 8856 22603 8890
rect 22643 8856 22677 8890
rect 22717 8856 22751 8890
rect 22791 8856 22825 8890
rect 22865 8856 22899 8890
rect 21572 8806 21606 8840
rect 21648 8806 21682 8840
rect 21724 8806 21758 8840
rect 21800 8806 21834 8840
rect 21876 8806 21910 8840
rect 21952 8806 21986 8840
rect 22027 8806 22061 8840
rect 22102 8806 22136 8840
rect 20808 8769 20842 8803
rect 20883 8769 20917 8803
rect 20958 8769 20992 8803
rect 21033 8769 21067 8803
rect 21108 8769 21142 8803
rect 21183 8769 21217 8803
rect 21258 8769 21292 8803
rect 21332 8769 21366 8803
rect 21406 8769 21440 8803
rect 21480 8769 21514 8803
rect 20808 8701 20842 8735
rect 20883 8701 20917 8735
rect 20958 8701 20992 8735
rect 21033 8701 21067 8735
rect 21108 8701 21142 8735
rect 21183 8701 21217 8735
rect 21258 8701 21292 8735
rect 21332 8701 21366 8735
rect 21406 8701 21440 8735
rect 21480 8701 21514 8735
rect 20808 8633 20842 8667
rect 20883 8633 20917 8667
rect 20958 8633 20992 8667
rect 21033 8633 21067 8667
rect 21108 8633 21142 8667
rect 21183 8633 21217 8667
rect 21258 8633 21292 8667
rect 21332 8633 21366 8667
rect 21406 8633 21440 8667
rect 21480 8633 21514 8667
rect 20808 8565 20842 8599
rect 20883 8565 20917 8599
rect 20958 8565 20992 8599
rect 21033 8565 21067 8599
rect 21108 8565 21142 8599
rect 21183 8565 21217 8599
rect 21258 8565 21292 8599
rect 21332 8565 21366 8599
rect 21406 8565 21440 8599
rect 21480 8565 21514 8599
rect 22194 8788 22228 8822
rect 22269 8788 22303 8822
rect 22344 8788 22378 8822
rect 22419 8788 22453 8822
rect 22494 8788 22528 8822
rect 22569 8788 22603 8822
rect 22643 8788 22677 8822
rect 22717 8788 22751 8822
rect 22791 8788 22825 8822
rect 22865 8788 22899 8822
rect 22194 8720 22228 8754
rect 22269 8720 22303 8754
rect 22344 8720 22378 8754
rect 22419 8720 22453 8754
rect 22494 8720 22528 8754
rect 22569 8720 22603 8754
rect 22643 8720 22677 8754
rect 22717 8720 22751 8754
rect 22791 8720 22825 8754
rect 22865 8720 22899 8754
rect 22194 8652 22228 8686
rect 22269 8652 22303 8686
rect 22344 8652 22378 8686
rect 22419 8652 22453 8686
rect 22494 8652 22528 8686
rect 22569 8652 22603 8686
rect 22643 8652 22677 8686
rect 22717 8652 22751 8686
rect 22791 8652 22825 8686
rect 22865 8652 22899 8686
rect 22194 8584 22228 8618
rect 22269 8584 22303 8618
rect 22344 8584 22378 8618
rect 22419 8584 22453 8618
rect 22494 8584 22528 8618
rect 22569 8584 22603 8618
rect 22643 8584 22677 8618
rect 22717 8584 22751 8618
rect 22791 8584 22825 8618
rect 22865 8584 22899 8618
rect 27547 8850 27581 8884
rect 27615 8850 27649 8884
rect 27683 8850 27717 8884
rect 27751 8850 27785 8884
rect 27819 8850 27853 8884
rect 27547 8780 27581 8814
rect 27615 8780 27649 8814
rect 27683 8780 27717 8814
rect 27751 8780 27785 8814
rect 27819 8780 27853 8814
rect 27547 8710 27581 8744
rect 27615 8710 27649 8744
rect 27683 8710 27717 8744
rect 27751 8710 27785 8744
rect 27819 8710 27853 8744
rect 27547 8640 27581 8674
rect 27615 8640 27649 8674
rect 27683 8640 27717 8674
rect 27751 8640 27785 8674
rect 27819 8640 27853 8674
rect 27547 8570 27581 8604
rect 27615 8570 27649 8604
rect 27683 8570 27717 8604
rect 27751 8570 27785 8604
rect 27819 8570 27853 8604
rect 192 8452 226 8486
rect 262 8452 296 8486
rect 332 8452 366 8486
rect 402 8452 436 8486
rect 472 8452 506 8486
rect 542 8452 576 8486
rect 612 8452 646 8486
rect 682 8452 716 8486
rect 752 8452 786 8486
rect 822 8452 856 8486
rect 891 8452 925 8486
rect 960 8452 994 8486
rect 1029 8452 1063 8486
rect 1098 8452 1132 8486
rect 1167 8452 1201 8486
rect 1236 8452 1270 8486
rect 1305 8452 1339 8486
rect 1374 8452 1408 8486
rect 1443 8452 1477 8486
rect 1512 8452 1546 8486
rect 1581 8452 1615 8486
rect 1650 8452 1684 8486
rect 1719 8452 1753 8486
rect 1788 8452 1822 8486
rect 192 8378 226 8412
rect 262 8378 296 8412
rect 332 8378 366 8412
rect 402 8378 436 8412
rect 472 8378 506 8412
rect 542 8378 576 8412
rect 612 8378 646 8412
rect 682 8378 716 8412
rect 752 8378 786 8412
rect 822 8378 856 8412
rect 891 8378 925 8412
rect 960 8378 994 8412
rect 1029 8378 1063 8412
rect 1098 8378 1132 8412
rect 1167 8378 1201 8412
rect 1236 8378 1270 8412
rect 1305 8378 1339 8412
rect 1374 8378 1408 8412
rect 1443 8378 1477 8412
rect 1512 8378 1546 8412
rect 1581 8378 1615 8412
rect 1650 8378 1684 8412
rect 1719 8378 1753 8412
rect 1788 8378 1822 8412
rect 192 8304 226 8338
rect 262 8304 296 8338
rect 332 8304 366 8338
rect 402 8304 436 8338
rect 472 8304 506 8338
rect 542 8304 576 8338
rect 612 8304 646 8338
rect 682 8304 716 8338
rect 752 8304 786 8338
rect 822 8304 856 8338
rect 891 8304 925 8338
rect 960 8304 994 8338
rect 1029 8304 1063 8338
rect 1098 8304 1132 8338
rect 1167 8304 1201 8338
rect 1236 8304 1270 8338
rect 1305 8304 1339 8338
rect 1374 8304 1408 8338
rect 1443 8304 1477 8338
rect 1512 8304 1546 8338
rect 1581 8304 1615 8338
rect 1650 8304 1684 8338
rect 1719 8304 1753 8338
rect 1788 8304 1822 8338
rect 175 8222 209 8256
rect 245 8222 279 8256
rect 315 8222 349 8256
rect 385 8222 419 8256
rect 455 8222 489 8256
rect 525 8222 559 8256
rect 595 8222 629 8256
rect 665 8222 699 8256
rect 735 8222 769 8256
rect 805 8222 839 8256
rect 7088 8429 7122 8463
rect 7212 8429 7246 8463
rect 7088 8360 7122 8394
rect 7212 8360 7246 8394
rect 27547 8500 27581 8534
rect 27615 8500 27649 8534
rect 27683 8500 27717 8534
rect 27751 8500 27785 8534
rect 27819 8500 27853 8534
rect 27547 8430 27581 8464
rect 27615 8430 27649 8464
rect 27683 8430 27717 8464
rect 27751 8430 27785 8464
rect 27819 8430 27853 8464
rect 7088 8291 7122 8325
rect 7212 8291 7246 8325
rect 175 8154 209 8188
rect 245 8154 279 8188
rect 315 8154 349 8188
rect 385 8154 419 8188
rect 455 8154 489 8188
rect 525 8154 559 8188
rect 595 8154 629 8188
rect 665 8154 699 8188
rect 735 8154 769 8188
rect 805 8154 839 8188
rect 175 8086 209 8120
rect 245 8086 279 8120
rect 315 8086 349 8120
rect 385 8086 419 8120
rect 455 8086 489 8120
rect 525 8086 559 8120
rect 595 8086 629 8120
rect 665 8086 699 8120
rect 735 8086 769 8120
rect 805 8086 839 8120
rect 175 8018 209 8052
rect 245 8018 279 8052
rect 315 8018 349 8052
rect 385 8018 419 8052
rect 455 8018 489 8052
rect 525 8018 559 8052
rect 595 8018 629 8052
rect 665 8018 699 8052
rect 735 8018 769 8052
rect 805 8018 839 8052
rect 175 7950 209 7984
rect 245 7950 279 7984
rect 315 7950 349 7984
rect 385 7950 419 7984
rect 455 7950 489 7984
rect 525 7950 559 7984
rect 595 7950 629 7984
rect 665 7950 699 7984
rect 735 7950 769 7984
rect 805 7950 839 7984
rect 175 7881 209 7915
rect 245 7881 279 7915
rect 315 7881 349 7915
rect 385 7881 419 7915
rect 455 7881 489 7915
rect 525 7881 559 7915
rect 595 7881 629 7915
rect 665 7881 699 7915
rect 735 7881 769 7915
rect 805 7881 839 7915
rect 175 7812 209 7846
rect 245 7812 279 7846
rect 315 7812 349 7846
rect 385 7812 419 7846
rect 455 7812 489 7846
rect 525 7812 559 7846
rect 595 7812 629 7846
rect 665 7812 699 7846
rect 735 7812 769 7846
rect 805 7812 839 7846
rect 175 7743 209 7777
rect 245 7743 279 7777
rect 315 7743 349 7777
rect 385 7743 419 7777
rect 455 7743 489 7777
rect 525 7743 559 7777
rect 595 7743 629 7777
rect 665 7743 699 7777
rect 735 7743 769 7777
rect 805 7743 839 7777
rect 175 7674 209 7708
rect 245 7674 279 7708
rect 315 7674 349 7708
rect 385 7674 419 7708
rect 455 7674 489 7708
rect 525 7674 559 7708
rect 595 7674 629 7708
rect 665 7674 699 7708
rect 735 7674 769 7708
rect 805 7674 839 7708
rect 175 7605 209 7639
rect 245 7605 279 7639
rect 315 7605 349 7639
rect 385 7605 419 7639
rect 455 7605 489 7639
rect 525 7605 559 7639
rect 595 7605 629 7639
rect 665 7605 699 7639
rect 735 7605 769 7639
rect 805 7605 839 7639
rect 175 7536 209 7570
rect 245 7536 279 7570
rect 315 7536 349 7570
rect 385 7536 419 7570
rect 455 7536 489 7570
rect 525 7536 559 7570
rect 595 7536 629 7570
rect 665 7536 699 7570
rect 735 7536 769 7570
rect 805 7536 839 7570
rect 175 7467 209 7501
rect 245 7467 279 7501
rect 315 7467 349 7501
rect 385 7467 419 7501
rect 455 7467 489 7501
rect 525 7467 559 7501
rect 595 7467 629 7501
rect 665 7467 699 7501
rect 735 7467 769 7501
rect 805 7467 839 7501
rect 175 7398 209 7432
rect 245 7398 279 7432
rect 315 7398 349 7432
rect 385 7398 419 7432
rect 455 7398 489 7432
rect 525 7398 559 7432
rect 595 7398 629 7432
rect 665 7398 699 7432
rect 735 7398 769 7432
rect 805 7398 839 7432
rect 175 7329 209 7363
rect 245 7329 279 7363
rect 315 7329 349 7363
rect 385 7329 419 7363
rect 455 7329 489 7363
rect 525 7329 559 7363
rect 595 7329 629 7363
rect 665 7329 699 7363
rect 735 7329 769 7363
rect 805 7329 839 7363
rect 175 7260 209 7294
rect 245 7260 279 7294
rect 315 7260 349 7294
rect 385 7260 419 7294
rect 455 7260 489 7294
rect 525 7260 559 7294
rect 595 7260 629 7294
rect 665 7260 699 7294
rect 735 7260 769 7294
rect 805 7260 839 7294
rect 7088 8222 7122 8256
rect 7212 8222 7246 8256
rect 7088 8153 7122 8187
rect 7212 8153 7246 8187
rect 7088 8084 7122 8118
rect 7212 8084 7246 8118
rect 7088 8014 7122 8048
rect 7212 8014 7246 8048
rect 7088 7944 7122 7978
rect 7212 7944 7246 7978
rect 7088 7874 7122 7908
rect 7212 7874 7246 7908
rect 7088 7804 7122 7838
rect 7212 7804 7246 7838
rect 7088 7734 7122 7768
rect 7212 7734 7246 7768
rect 7088 7664 7122 7698
rect 7212 7664 7246 7698
rect 27270 8320 27304 8354
rect 27338 8320 27372 8354
rect 27406 8320 27440 8354
rect 27474 8320 27508 8354
rect 27542 8320 27576 8354
rect 27610 8320 27644 8354
rect 27678 8320 27712 8354
rect 27746 8320 27780 8354
rect 27814 8320 27848 8354
rect 27270 8249 27304 8283
rect 27338 8249 27372 8283
rect 27406 8249 27440 8283
rect 27474 8249 27508 8283
rect 27542 8249 27576 8283
rect 27610 8249 27644 8283
rect 27678 8249 27712 8283
rect 27746 8249 27780 8283
rect 27814 8249 27848 8283
rect 27270 8178 27304 8212
rect 27338 8178 27372 8212
rect 27406 8178 27440 8212
rect 27474 8178 27508 8212
rect 27542 8178 27576 8212
rect 27610 8178 27644 8212
rect 27678 8178 27712 8212
rect 27746 8178 27780 8212
rect 27814 8178 27848 8212
rect 27270 8107 27304 8141
rect 27338 8107 27372 8141
rect 27406 8107 27440 8141
rect 27474 8107 27508 8141
rect 27542 8107 27576 8141
rect 27610 8107 27644 8141
rect 27678 8107 27712 8141
rect 27746 8107 27780 8141
rect 27814 8107 27848 8141
rect 27270 8036 27304 8070
rect 27338 8036 27372 8070
rect 27406 8036 27440 8070
rect 27474 8036 27508 8070
rect 27542 8036 27576 8070
rect 27610 8036 27644 8070
rect 27678 8036 27712 8070
rect 27746 8036 27780 8070
rect 27814 8036 27848 8070
rect 27270 7965 27304 7999
rect 27338 7965 27372 7999
rect 27406 7965 27440 7999
rect 27474 7965 27508 7999
rect 27542 7965 27576 7999
rect 27610 7965 27644 7999
rect 27678 7965 27712 7999
rect 27746 7965 27780 7999
rect 27814 7965 27848 7999
rect 27270 7894 27304 7928
rect 27338 7894 27372 7928
rect 27406 7894 27440 7928
rect 27474 7894 27508 7928
rect 27542 7894 27576 7928
rect 27610 7894 27644 7928
rect 27678 7894 27712 7928
rect 27746 7894 27780 7928
rect 27814 7894 27848 7928
rect 27270 7823 27304 7857
rect 27338 7823 27372 7857
rect 27406 7823 27440 7857
rect 27474 7823 27508 7857
rect 27542 7823 27576 7857
rect 27610 7823 27644 7857
rect 27678 7823 27712 7857
rect 27746 7823 27780 7857
rect 27814 7823 27848 7857
rect 27270 7752 27304 7786
rect 27338 7752 27372 7786
rect 27406 7752 27440 7786
rect 27474 7752 27508 7786
rect 27542 7752 27576 7786
rect 27610 7752 27644 7786
rect 27678 7752 27712 7786
rect 27746 7752 27780 7786
rect 27814 7752 27848 7786
rect 27270 7680 27304 7714
rect 27338 7680 27372 7714
rect 27406 7680 27440 7714
rect 27474 7680 27508 7714
rect 27542 7680 27576 7714
rect 27610 7680 27644 7714
rect 27678 7680 27712 7714
rect 27746 7680 27780 7714
rect 27814 7680 27848 7714
rect 7088 7594 7122 7628
rect 7212 7594 7246 7628
rect 7088 7524 7122 7558
rect 7212 7524 7246 7558
rect 7088 7454 7122 7488
rect 7212 7454 7246 7488
rect 7088 7384 7122 7418
rect 7212 7384 7246 7418
rect 7088 7314 7122 7348
rect 7212 7314 7246 7348
rect 175 7191 209 7225
rect 245 7191 279 7225
rect 315 7191 349 7225
rect 385 7191 419 7225
rect 455 7191 489 7225
rect 525 7191 559 7225
rect 595 7191 629 7225
rect 665 7191 699 7225
rect 735 7191 769 7225
rect 805 7191 839 7225
rect 175 7122 209 7156
rect 245 7122 279 7156
rect 315 7122 349 7156
rect 385 7122 419 7156
rect 455 7122 489 7156
rect 525 7122 559 7156
rect 595 7122 629 7156
rect 665 7122 699 7156
rect 735 7122 769 7156
rect 805 7122 839 7156
rect 175 7053 209 7087
rect 245 7053 279 7087
rect 315 7053 349 7087
rect 385 7053 419 7087
rect 455 7053 489 7087
rect 525 7053 559 7087
rect 595 7053 629 7087
rect 665 7053 699 7087
rect 735 7053 769 7087
rect 805 7053 839 7087
rect 175 6984 209 7018
rect 245 6984 279 7018
rect 315 6984 349 7018
rect 385 6984 419 7018
rect 455 6984 489 7018
rect 525 6984 559 7018
rect 595 6984 629 7018
rect 665 6984 699 7018
rect 735 6984 769 7018
rect 805 6984 839 7018
rect 175 6915 209 6949
rect 245 6915 279 6949
rect 315 6915 349 6949
rect 385 6915 419 6949
rect 455 6915 489 6949
rect 525 6915 559 6949
rect 595 6915 629 6949
rect 665 6915 699 6949
rect 735 6915 769 6949
rect 805 6915 839 6949
rect 14262 6979 14296 7013
rect 14334 6979 14368 7013
rect 14406 6979 14440 7013
rect 14478 6979 14512 7013
rect 14550 6979 14584 7013
rect 14622 6979 14656 7013
rect 14694 6979 14728 7013
rect 14766 6979 14800 7013
rect 14838 6979 14872 7013
rect 14910 6979 14944 7013
rect 14982 6979 15016 7013
rect 15054 6979 15088 7013
rect 175 6846 209 6880
rect 245 6846 279 6880
rect 315 6846 349 6880
rect 385 6846 419 6880
rect 455 6846 489 6880
rect 525 6846 559 6880
rect 595 6846 629 6880
rect 665 6846 699 6880
rect 735 6846 769 6880
rect 805 6846 839 6880
rect 175 6777 209 6811
rect 245 6777 279 6811
rect 315 6777 349 6811
rect 385 6777 419 6811
rect 455 6777 489 6811
rect 525 6777 559 6811
rect 595 6777 629 6811
rect 665 6777 699 6811
rect 735 6777 769 6811
rect 805 6777 839 6811
rect 175 6708 209 6742
rect 245 6708 279 6742
rect 315 6708 349 6742
rect 385 6708 419 6742
rect 455 6708 489 6742
rect 525 6708 559 6742
rect 595 6708 629 6742
rect 665 6708 699 6742
rect 735 6708 769 6742
rect 805 6708 839 6742
rect 175 6639 209 6673
rect 245 6639 279 6673
rect 315 6639 349 6673
rect 385 6639 419 6673
rect 455 6639 489 6673
rect 525 6639 559 6673
rect 595 6639 629 6673
rect 665 6639 699 6673
rect 735 6639 769 6673
rect 805 6639 839 6673
rect 175 6570 209 6604
rect 245 6570 279 6604
rect 315 6570 349 6604
rect 385 6570 419 6604
rect 455 6570 489 6604
rect 525 6570 559 6604
rect 595 6570 629 6604
rect 665 6570 699 6604
rect 735 6570 769 6604
rect 805 6570 839 6604
rect 175 6501 209 6535
rect 245 6501 279 6535
rect 315 6501 349 6535
rect 385 6501 419 6535
rect 455 6501 489 6535
rect 525 6501 559 6535
rect 595 6501 629 6535
rect 665 6501 699 6535
rect 735 6501 769 6535
rect 805 6501 839 6535
rect 175 6432 209 6466
rect 245 6432 279 6466
rect 315 6432 349 6466
rect 385 6432 419 6466
rect 455 6432 489 6466
rect 525 6432 559 6466
rect 595 6432 629 6466
rect 665 6432 699 6466
rect 735 6432 769 6466
rect 805 6432 839 6466
rect 175 6363 209 6397
rect 245 6363 279 6397
rect 315 6363 349 6397
rect 385 6363 419 6397
rect 455 6363 489 6397
rect 525 6363 559 6397
rect 595 6363 629 6397
rect 665 6363 699 6397
rect 735 6363 769 6397
rect 805 6363 839 6397
rect 175 6294 209 6328
rect 245 6294 279 6328
rect 315 6294 349 6328
rect 385 6294 419 6328
rect 455 6294 489 6328
rect 525 6294 559 6328
rect 595 6294 629 6328
rect 665 6294 699 6328
rect 735 6294 769 6328
rect 805 6294 839 6328
rect 13054 6889 13088 6923
rect 13123 6889 13157 6923
rect 13192 6889 13226 6923
rect 13261 6889 13295 6923
rect 13330 6889 13364 6923
rect 13399 6889 13433 6923
rect 13467 6889 13501 6923
rect 13535 6889 13569 6923
rect 13603 6889 13637 6923
rect 13671 6889 13705 6923
rect 13739 6889 13773 6923
rect 13807 6889 13841 6923
rect 13875 6889 13909 6923
rect 13943 6889 13977 6923
rect 14011 6889 14045 6923
rect 14079 6889 14113 6923
rect 14147 6889 14181 6923
rect 14262 6906 14296 6940
rect 14334 6906 14368 6940
rect 14406 6906 14440 6940
rect 14478 6906 14512 6940
rect 14550 6906 14584 6940
rect 14622 6906 14656 6940
rect 14694 6906 14728 6940
rect 14766 6906 14800 6940
rect 14838 6906 14872 6940
rect 14910 6906 14944 6940
rect 14982 6906 15016 6940
rect 15054 6906 15088 6940
rect 13054 6815 13088 6849
rect 13123 6815 13157 6849
rect 13192 6815 13226 6849
rect 13261 6815 13295 6849
rect 13330 6815 13364 6849
rect 13399 6815 13433 6849
rect 13467 6815 13501 6849
rect 13535 6815 13569 6849
rect 13603 6815 13637 6849
rect 13671 6815 13705 6849
rect 13739 6815 13773 6849
rect 13807 6815 13841 6849
rect 13875 6815 13909 6849
rect 13943 6815 13977 6849
rect 14011 6815 14045 6849
rect 14079 6815 14113 6849
rect 14147 6815 14181 6849
rect 14262 6832 14296 6866
rect 14334 6832 14368 6866
rect 14406 6832 14440 6866
rect 14478 6832 14512 6866
rect 14550 6832 14584 6866
rect 14622 6832 14656 6866
rect 14694 6832 14728 6866
rect 14766 6832 14800 6866
rect 14838 6832 14872 6866
rect 14910 6832 14944 6866
rect 14982 6832 15016 6866
rect 15054 6832 15088 6866
rect 13054 6741 13088 6775
rect 13123 6741 13157 6775
rect 13192 6741 13226 6775
rect 13261 6741 13295 6775
rect 13330 6741 13364 6775
rect 13399 6741 13433 6775
rect 13467 6741 13501 6775
rect 13535 6741 13569 6775
rect 13603 6741 13637 6775
rect 13671 6741 13705 6775
rect 13739 6741 13773 6775
rect 13807 6741 13841 6775
rect 13875 6741 13909 6775
rect 13943 6741 13977 6775
rect 14011 6741 14045 6775
rect 14079 6741 14113 6775
rect 14147 6741 14181 6775
rect 14262 6758 14296 6792
rect 14334 6758 14368 6792
rect 14406 6758 14440 6792
rect 14478 6758 14512 6792
rect 14550 6758 14584 6792
rect 14622 6758 14656 6792
rect 14694 6758 14728 6792
rect 14766 6758 14800 6792
rect 14838 6758 14872 6792
rect 14910 6758 14944 6792
rect 14982 6758 15016 6792
rect 15054 6758 15088 6792
rect 13054 6667 13088 6701
rect 13123 6667 13157 6701
rect 13192 6667 13226 6701
rect 13261 6667 13295 6701
rect 13330 6667 13364 6701
rect 13399 6667 13433 6701
rect 13467 6667 13501 6701
rect 13535 6667 13569 6701
rect 13603 6667 13637 6701
rect 13671 6667 13705 6701
rect 13739 6667 13773 6701
rect 13807 6667 13841 6701
rect 13875 6667 13909 6701
rect 13943 6667 13977 6701
rect 14011 6667 14045 6701
rect 14079 6667 14113 6701
rect 14147 6667 14181 6701
rect 14262 6684 14296 6718
rect 14334 6684 14368 6718
rect 14406 6684 14440 6718
rect 14478 6684 14512 6718
rect 14550 6684 14584 6718
rect 14622 6684 14656 6718
rect 14694 6684 14728 6718
rect 14766 6684 14800 6718
rect 14838 6684 14872 6718
rect 14910 6684 14944 6718
rect 14982 6684 15016 6718
rect 15054 6684 15088 6718
rect 13054 6593 13088 6627
rect 13123 6593 13157 6627
rect 13192 6593 13226 6627
rect 13261 6593 13295 6627
rect 13330 6593 13364 6627
rect 13399 6593 13433 6627
rect 13467 6593 13501 6627
rect 13535 6593 13569 6627
rect 13603 6593 13637 6627
rect 13671 6593 13705 6627
rect 13739 6593 13773 6627
rect 13807 6593 13841 6627
rect 13875 6593 13909 6627
rect 13943 6593 13977 6627
rect 14011 6593 14045 6627
rect 14079 6593 14113 6627
rect 14147 6593 14181 6627
rect 14262 6610 14296 6644
rect 14334 6610 14368 6644
rect 14406 6610 14440 6644
rect 14478 6610 14512 6644
rect 14550 6610 14584 6644
rect 14622 6610 14656 6644
rect 14694 6610 14728 6644
rect 14766 6610 14800 6644
rect 14838 6610 14872 6644
rect 14910 6610 14944 6644
rect 14982 6610 15016 6644
rect 15054 6610 15088 6644
rect 13054 6519 13088 6553
rect 13123 6519 13157 6553
rect 13192 6519 13226 6553
rect 13261 6519 13295 6553
rect 13330 6519 13364 6553
rect 13399 6519 13433 6553
rect 13467 6519 13501 6553
rect 13535 6519 13569 6553
rect 13603 6519 13637 6553
rect 13671 6519 13705 6553
rect 13739 6519 13773 6553
rect 13807 6519 13841 6553
rect 13875 6519 13909 6553
rect 13943 6519 13977 6553
rect 14011 6519 14045 6553
rect 14079 6519 14113 6553
rect 14147 6519 14181 6553
rect 14262 6536 14296 6570
rect 14334 6536 14368 6570
rect 14406 6536 14440 6570
rect 14478 6536 14512 6570
rect 14550 6536 14584 6570
rect 14622 6536 14656 6570
rect 14694 6536 14728 6570
rect 14766 6536 14800 6570
rect 14838 6536 14872 6570
rect 14910 6536 14944 6570
rect 14982 6536 15016 6570
rect 15054 6536 15088 6570
rect 13054 6445 13088 6479
rect 13123 6445 13157 6479
rect 13192 6445 13226 6479
rect 13261 6445 13295 6479
rect 13330 6445 13364 6479
rect 13399 6445 13433 6479
rect 13467 6445 13501 6479
rect 13535 6445 13569 6479
rect 13603 6445 13637 6479
rect 13671 6445 13705 6479
rect 13739 6445 13773 6479
rect 13807 6445 13841 6479
rect 13875 6445 13909 6479
rect 13943 6445 13977 6479
rect 14011 6445 14045 6479
rect 14079 6445 14113 6479
rect 14147 6445 14181 6479
rect 14262 6462 14296 6496
rect 14334 6462 14368 6496
rect 14406 6462 14440 6496
rect 14478 6462 14512 6496
rect 14550 6462 14584 6496
rect 14622 6462 14656 6496
rect 14694 6462 14728 6496
rect 14766 6462 14800 6496
rect 14838 6462 14872 6496
rect 14910 6462 14944 6496
rect 14982 6462 15016 6496
rect 15054 6462 15088 6496
rect 13054 6371 13088 6405
rect 13123 6371 13157 6405
rect 13192 6371 13226 6405
rect 13261 6371 13295 6405
rect 13330 6371 13364 6405
rect 13399 6371 13433 6405
rect 13467 6371 13501 6405
rect 13535 6371 13569 6405
rect 13603 6371 13637 6405
rect 13671 6371 13705 6405
rect 13739 6371 13773 6405
rect 13807 6371 13841 6405
rect 13875 6371 13909 6405
rect 13943 6371 13977 6405
rect 14011 6371 14045 6405
rect 14079 6371 14113 6405
rect 14147 6371 14181 6405
rect 14262 6388 14296 6422
rect 14334 6388 14368 6422
rect 14406 6388 14440 6422
rect 14478 6388 14512 6422
rect 14550 6388 14584 6422
rect 14622 6388 14656 6422
rect 14694 6388 14728 6422
rect 14766 6388 14800 6422
rect 14838 6388 14872 6422
rect 14910 6388 14944 6422
rect 14982 6388 15016 6422
rect 15054 6388 15088 6422
rect 13054 6297 13088 6331
rect 13123 6297 13157 6331
rect 13192 6297 13226 6331
rect 13261 6297 13295 6331
rect 13330 6297 13364 6331
rect 13399 6297 13433 6331
rect 13467 6297 13501 6331
rect 13535 6297 13569 6331
rect 13603 6297 13637 6331
rect 13671 6297 13705 6331
rect 13739 6297 13773 6331
rect 13807 6297 13841 6331
rect 13875 6297 13909 6331
rect 13943 6297 13977 6331
rect 14011 6297 14045 6331
rect 14079 6297 14113 6331
rect 14147 6297 14181 6331
rect 14262 6314 14296 6348
rect 14334 6314 14368 6348
rect 14406 6314 14440 6348
rect 14478 6314 14512 6348
rect 14550 6314 14584 6348
rect 14622 6314 14656 6348
rect 14694 6314 14728 6348
rect 14766 6314 14800 6348
rect 14838 6314 14872 6348
rect 14910 6314 14944 6348
rect 14982 6314 15016 6348
rect 15054 6314 15088 6348
rect 175 6225 209 6259
rect 245 6225 279 6259
rect 315 6225 349 6259
rect 385 6225 419 6259
rect 455 6225 489 6259
rect 525 6225 559 6259
rect 595 6225 629 6259
rect 665 6225 699 6259
rect 735 6225 769 6259
rect 805 6225 839 6259
rect 169 6091 203 6125
rect 245 6091 279 6125
rect 321 6091 355 6125
rect 169 6022 203 6056
rect 245 6022 279 6056
rect 321 6022 355 6056
rect 169 5953 203 5987
rect 245 5953 279 5987
rect 321 5953 355 5987
rect 169 5884 203 5918
rect 245 5884 279 5918
rect 321 5884 355 5918
rect 169 5815 203 5849
rect 245 5815 279 5849
rect 321 5815 355 5849
rect 169 5746 203 5780
rect 245 5746 279 5780
rect 321 5746 355 5780
rect 169 5677 203 5711
rect 245 5677 279 5711
rect 321 5677 355 5711
rect 169 5608 203 5642
rect 245 5608 279 5642
rect 321 5608 355 5642
rect 169 5539 203 5573
rect 245 5539 279 5573
rect 321 5539 355 5573
rect 169 5470 203 5504
rect 245 5470 279 5504
rect 321 5470 355 5504
rect 169 5401 203 5435
rect 245 5401 279 5435
rect 321 5401 355 5435
rect 169 5332 203 5366
rect 245 5332 279 5366
rect 321 5332 355 5366
rect 169 5263 203 5297
rect 245 5263 279 5297
rect 321 5263 355 5297
rect 169 5194 203 5228
rect 245 5194 279 5228
rect 321 5194 355 5228
rect 169 5125 203 5159
rect 245 5125 279 5159
rect 321 5125 355 5159
rect 169 5056 203 5090
rect 245 5056 279 5090
rect 321 5056 355 5090
rect 169 4987 203 5021
rect 245 4987 279 5021
rect 321 4987 355 5021
rect 169 4918 203 4952
rect 245 4918 279 4952
rect 321 4918 355 4952
rect 169 4849 203 4883
rect 245 4849 279 4883
rect 321 4849 355 4883
rect 169 4780 203 4814
rect 245 4780 279 4814
rect 321 4780 355 4814
rect 169 4711 203 4745
rect 245 4711 279 4745
rect 321 4711 355 4745
rect 169 4642 203 4676
rect 245 4642 279 4676
rect 321 4642 355 4676
rect 169 4573 203 4607
rect 245 4573 279 4607
rect 321 4573 355 4607
rect 169 4504 203 4538
rect 245 4504 279 4538
rect 321 4504 355 4538
rect 169 4435 203 4469
rect 245 4435 279 4469
rect 321 4435 355 4469
rect 169 4366 203 4400
rect 245 4366 279 4400
rect 321 4366 355 4400
rect 169 4297 203 4331
rect 245 4297 279 4331
rect 321 4297 355 4331
rect 169 4228 203 4262
rect 245 4228 279 4262
rect 321 4228 355 4262
rect 169 4159 203 4193
rect 245 4159 279 4193
rect 321 4159 355 4193
rect 169 4090 203 4124
rect 245 4090 279 4124
rect 321 4090 355 4124
rect 169 4021 203 4055
rect 245 4021 279 4055
rect 321 4021 355 4055
rect 442 4047 476 4081
rect 512 4047 546 4081
rect 582 4047 616 4081
rect 652 4047 686 4081
rect 722 4047 756 4081
rect 792 4047 826 4081
rect 862 4047 896 4081
rect 932 4047 966 4081
rect 1002 4047 1036 4081
rect 1072 4047 1106 4081
rect 1142 4047 1176 4081
rect 1212 4047 1246 4081
rect 1282 4047 1316 4081
rect 1352 4047 1386 4081
rect 1422 4047 1456 4081
rect 1492 4047 1526 4081
rect 1562 4047 1596 4081
rect 1632 4047 1666 4081
rect 1702 4047 1736 4081
rect 1772 4047 1806 4081
rect 1842 4047 1876 4081
rect 1912 4047 1946 4081
rect 1982 4047 2016 4081
rect 2052 4047 2086 4081
rect 169 3952 203 3986
rect 245 3952 279 3986
rect 321 3952 355 3986
rect 442 3921 476 3955
rect 512 3921 546 3955
rect 582 3921 616 3955
rect 652 3921 686 3955
rect 722 3921 756 3955
rect 792 3921 826 3955
rect 862 3921 896 3955
rect 932 3921 966 3955
rect 1002 3921 1036 3955
rect 1072 3921 1106 3955
rect 1142 3921 1176 3955
rect 1212 3921 1246 3955
rect 1282 3921 1316 3955
rect 1352 3921 1386 3955
rect 1422 3921 1456 3955
rect 1492 3921 1526 3955
rect 1562 3921 1596 3955
rect 1632 3921 1666 3955
rect 1702 3921 1736 3955
rect 1772 3921 1806 3955
rect 1842 3921 1876 3955
rect 1912 3921 1946 3955
rect 1982 3921 2016 3955
rect 2052 3921 2086 3955
rect 169 3883 203 3917
rect 245 3883 279 3917
rect 321 3883 355 3917
rect 169 3814 203 3848
rect 245 3814 279 3848
rect 321 3814 355 3848
rect 410 3811 444 3845
rect 484 3811 518 3845
rect 558 3811 592 3845
rect 632 3811 666 3845
rect 169 3745 203 3779
rect 245 3745 279 3779
rect 321 3745 355 3779
rect 410 3740 444 3774
rect 484 3740 518 3774
rect 558 3740 592 3774
rect 632 3740 666 3774
rect 169 3676 203 3710
rect 245 3676 279 3710
rect 321 3676 355 3710
rect 410 3668 444 3702
rect 484 3668 518 3702
rect 558 3668 592 3702
rect 632 3668 666 3702
rect 169 3607 203 3641
rect 245 3607 279 3641
rect 321 3607 355 3641
rect 410 3596 444 3630
rect 484 3596 518 3630
rect 558 3596 592 3630
rect 632 3596 666 3630
rect 169 3537 203 3571
rect 245 3537 279 3571
rect 321 3537 355 3571
rect 410 3524 444 3558
rect 484 3524 518 3558
rect 558 3524 592 3558
rect 632 3524 666 3558
rect 169 3467 203 3501
rect 245 3467 279 3501
rect 321 3467 355 3501
rect 410 3452 444 3486
rect 484 3452 518 3486
rect 558 3452 592 3486
rect 632 3452 666 3486
rect 169 3397 203 3431
rect 245 3397 279 3431
rect 321 3397 355 3431
rect 410 3380 444 3414
rect 484 3380 518 3414
rect 558 3380 592 3414
rect 632 3380 666 3414
rect 169 3327 203 3361
rect 245 3327 279 3361
rect 321 3327 355 3361
rect 410 3308 444 3342
rect 484 3308 518 3342
rect 558 3308 592 3342
rect 632 3308 666 3342
rect 169 3257 203 3291
rect 245 3257 279 3291
rect 321 3257 355 3291
rect 410 3236 444 3270
rect 484 3236 518 3270
rect 558 3236 592 3270
rect 632 3236 666 3270
rect 169 3187 203 3221
rect 245 3187 279 3221
rect 321 3187 355 3221
rect 410 3164 444 3198
rect 484 3164 518 3198
rect 558 3164 592 3198
rect 632 3164 666 3198
rect 169 3117 203 3151
rect 245 3117 279 3151
rect 321 3117 355 3151
rect 1373 3807 1407 3841
rect 1449 3807 1483 3841
rect 1525 3807 1559 3841
rect 1601 3807 1635 3841
rect 1677 3807 1711 3841
rect 1752 3807 1786 3841
rect 1827 3807 1861 3841
rect 1902 3807 1936 3841
rect 1977 3807 2011 3841
rect 2052 3807 2086 3841
rect 1373 3727 1407 3761
rect 1449 3727 1483 3761
rect 1525 3727 1559 3761
rect 1601 3727 1635 3761
rect 1677 3727 1711 3761
rect 1752 3727 1786 3761
rect 1827 3727 1861 3761
rect 1902 3727 1936 3761
rect 1977 3727 2011 3761
rect 2052 3727 2086 3761
rect 1373 3647 1407 3681
rect 1449 3647 1483 3681
rect 1525 3647 1559 3681
rect 1601 3647 1635 3681
rect 1677 3647 1711 3681
rect 1752 3647 1786 3681
rect 1827 3647 1861 3681
rect 1902 3647 1936 3681
rect 1977 3647 2011 3681
rect 2052 3647 2086 3681
rect 1373 3567 1407 3601
rect 1449 3567 1483 3601
rect 1525 3567 1559 3601
rect 1601 3567 1635 3601
rect 1677 3567 1711 3601
rect 1752 3567 1786 3601
rect 1827 3567 1861 3601
rect 1902 3567 1936 3601
rect 1977 3567 2011 3601
rect 2052 3567 2086 3601
rect 1373 3487 1407 3521
rect 1449 3487 1483 3521
rect 1525 3487 1559 3521
rect 1601 3487 1635 3521
rect 1677 3487 1711 3521
rect 1752 3487 1786 3521
rect 1827 3487 1861 3521
rect 1902 3487 1936 3521
rect 1977 3487 2011 3521
rect 2052 3487 2086 3521
rect 1373 3407 1407 3441
rect 1449 3407 1483 3441
rect 1525 3407 1559 3441
rect 1601 3407 1635 3441
rect 1677 3407 1711 3441
rect 1752 3407 1786 3441
rect 1827 3407 1861 3441
rect 1902 3407 1936 3441
rect 1977 3407 2011 3441
rect 2052 3407 2086 3441
rect 1389 3337 1423 3371
rect 1464 3337 1498 3371
rect 1539 3337 1573 3371
rect 1614 3337 1648 3371
rect 1689 3337 1723 3371
rect 1764 3337 1798 3371
rect 1839 3337 1873 3371
rect 1914 3337 1948 3371
rect 1988 3337 2022 3371
rect 2062 3337 2096 3371
rect 1389 3269 1423 3303
rect 1464 3269 1498 3303
rect 1539 3269 1573 3303
rect 1614 3269 1648 3303
rect 1689 3269 1723 3303
rect 1764 3269 1798 3303
rect 1839 3269 1873 3303
rect 1914 3269 1948 3303
rect 1988 3269 2022 3303
rect 2062 3269 2096 3303
rect 1363 3199 1397 3233
rect 1432 3199 1466 3233
rect 1501 3199 1535 3233
rect 1570 3199 1604 3233
rect 1639 3199 1673 3233
rect 1708 3199 1742 3233
rect 1777 3199 1811 3233
rect 1846 3199 1880 3233
rect 1915 3199 1949 3233
rect 1984 3199 2018 3233
rect 2053 3199 2087 3233
rect 2122 3199 2156 3233
rect 2191 3199 2225 3233
rect 2259 3199 2293 3233
rect 2327 3199 2361 3233
rect 2395 3199 2429 3233
rect 2463 3199 2497 3233
rect 2531 3199 2565 3233
rect 2599 3199 2633 3233
rect 2667 3199 2701 3233
rect 2735 3199 2769 3233
rect 2803 3199 2837 3233
rect 2871 3199 2905 3233
rect 2939 3199 2973 3233
rect 3007 3199 3041 3233
rect 3075 3199 3109 3233
rect 1363 3125 1397 3159
rect 1432 3125 1466 3159
rect 1501 3125 1535 3159
rect 1570 3125 1604 3159
rect 1639 3125 1673 3159
rect 1708 3125 1742 3159
rect 1777 3125 1811 3159
rect 1846 3125 1880 3159
rect 1915 3125 1949 3159
rect 1984 3125 2018 3159
rect 2053 3125 2087 3159
rect 2122 3125 2156 3159
rect 2191 3125 2225 3159
rect 2259 3125 2293 3159
rect 2327 3125 2361 3159
rect 2395 3125 2429 3159
rect 2463 3125 2497 3159
rect 2531 3125 2565 3159
rect 2599 3125 2633 3159
rect 2667 3125 2701 3159
rect 2735 3125 2769 3159
rect 2803 3125 2837 3159
rect 2871 3125 2905 3159
rect 2939 3125 2973 3159
rect 3007 3125 3041 3159
rect 3075 3125 3109 3159
rect 169 3047 203 3081
rect 245 3047 279 3081
rect 321 3047 355 3081
rect 410 3053 444 3087
rect 481 3053 515 3087
rect 552 3053 586 3087
rect 623 3053 657 3087
rect 694 3053 728 3087
rect 765 3053 799 3087
rect 835 3053 869 3087
rect 905 3053 939 3087
rect 975 3053 1009 3087
rect 1045 3053 1079 3087
rect 1115 3053 1149 3087
rect 1185 3053 1219 3087
rect 1255 3053 1289 3087
rect 1363 3051 1397 3085
rect 1432 3051 1466 3085
rect 1501 3051 1535 3085
rect 1570 3051 1604 3085
rect 1639 3051 1673 3085
rect 1708 3051 1742 3085
rect 1777 3051 1811 3085
rect 1846 3051 1880 3085
rect 1915 3051 1949 3085
rect 1984 3051 2018 3085
rect 2053 3051 2087 3085
rect 2122 3051 2156 3085
rect 2191 3051 2225 3085
rect 2259 3051 2293 3085
rect 2327 3051 2361 3085
rect 2395 3051 2429 3085
rect 2463 3051 2497 3085
rect 2531 3051 2565 3085
rect 2599 3051 2633 3085
rect 2667 3051 2701 3085
rect 2735 3051 2769 3085
rect 2803 3051 2837 3085
rect 2871 3051 2905 3085
rect 2939 3051 2973 3085
rect 3007 3051 3041 3085
rect 3075 3051 3109 3085
rect 169 2977 203 3011
rect 245 2977 279 3011
rect 321 2977 355 3011
rect 410 2979 444 3013
rect 481 2979 515 3013
rect 552 2979 586 3013
rect 623 2979 657 3013
rect 694 2979 728 3013
rect 765 2979 799 3013
rect 835 2979 869 3013
rect 905 2979 939 3013
rect 975 2979 1009 3013
rect 1045 2979 1079 3013
rect 1115 2979 1149 3013
rect 1185 2979 1219 3013
rect 1255 2979 1289 3013
rect 1363 2977 1397 3011
rect 1432 2977 1466 3011
rect 1501 2977 1535 3011
rect 1570 2977 1604 3011
rect 1639 2977 1673 3011
rect 1708 2977 1742 3011
rect 1777 2977 1811 3011
rect 1846 2977 1880 3011
rect 1915 2977 1949 3011
rect 1984 2977 2018 3011
rect 2053 2977 2087 3011
rect 2122 2977 2156 3011
rect 2191 2977 2225 3011
rect 2259 2977 2293 3011
rect 2327 2977 2361 3011
rect 2395 2977 2429 3011
rect 2463 2977 2497 3011
rect 2531 2977 2565 3011
rect 2599 2977 2633 3011
rect 2667 2977 2701 3011
rect 2735 2977 2769 3011
rect 2803 2977 2837 3011
rect 2871 2977 2905 3011
rect 2939 2977 2973 3011
rect 3007 2977 3041 3011
rect 3075 2977 3109 3011
rect 169 2907 203 2941
rect 245 2907 279 2941
rect 321 2907 355 2941
rect 410 2905 444 2939
rect 481 2905 515 2939
rect 552 2905 586 2939
rect 623 2905 657 2939
rect 694 2905 728 2939
rect 765 2905 799 2939
rect 835 2905 869 2939
rect 905 2905 939 2939
rect 975 2905 1009 2939
rect 1045 2905 1079 2939
rect 1115 2905 1149 2939
rect 1185 2905 1219 2939
rect 1255 2905 1289 2939
rect 1363 2903 1397 2937
rect 1432 2903 1466 2937
rect 1501 2903 1535 2937
rect 1570 2903 1604 2937
rect 1639 2903 1673 2937
rect 1708 2903 1742 2937
rect 1777 2903 1811 2937
rect 1846 2903 1880 2937
rect 1915 2903 1949 2937
rect 1984 2903 2018 2937
rect 2053 2903 2087 2937
rect 2122 2903 2156 2937
rect 2191 2903 2225 2937
rect 2259 2903 2293 2937
rect 2327 2903 2361 2937
rect 2395 2903 2429 2937
rect 2463 2903 2497 2937
rect 2531 2903 2565 2937
rect 2599 2903 2633 2937
rect 2667 2903 2701 2937
rect 2735 2903 2769 2937
rect 2803 2903 2837 2937
rect 2871 2903 2905 2937
rect 2939 2903 2973 2937
rect 3007 2903 3041 2937
rect 3075 2903 3109 2937
rect 169 2837 203 2871
rect 245 2837 279 2871
rect 321 2837 355 2871
rect 410 2831 444 2865
rect 481 2831 515 2865
rect 552 2831 586 2865
rect 623 2831 657 2865
rect 694 2831 728 2865
rect 765 2831 799 2865
rect 835 2831 869 2865
rect 905 2831 939 2865
rect 975 2831 1009 2865
rect 1045 2831 1079 2865
rect 1115 2831 1149 2865
rect 1185 2831 1219 2865
rect 1255 2831 1289 2865
rect 1363 2829 1397 2863
rect 1432 2829 1466 2863
rect 1501 2829 1535 2863
rect 1570 2829 1604 2863
rect 1639 2829 1673 2863
rect 1708 2829 1742 2863
rect 1777 2829 1811 2863
rect 1846 2829 1880 2863
rect 1915 2829 1949 2863
rect 1984 2829 2018 2863
rect 2053 2829 2087 2863
rect 2122 2829 2156 2863
rect 2191 2829 2225 2863
rect 2259 2829 2293 2863
rect 2327 2829 2361 2863
rect 2395 2829 2429 2863
rect 2463 2829 2497 2863
rect 2531 2829 2565 2863
rect 2599 2829 2633 2863
rect 2667 2829 2701 2863
rect 2735 2829 2769 2863
rect 2803 2829 2837 2863
rect 2871 2829 2905 2863
rect 2939 2829 2973 2863
rect 3007 2829 3041 2863
rect 3075 2829 3109 2863
rect 169 2767 203 2801
rect 245 2767 279 2801
rect 321 2767 355 2801
rect 410 2757 444 2791
rect 481 2757 515 2791
rect 552 2757 586 2791
rect 623 2757 657 2791
rect 694 2757 728 2791
rect 765 2757 799 2791
rect 835 2757 869 2791
rect 905 2757 939 2791
rect 975 2757 1009 2791
rect 1045 2757 1079 2791
rect 1115 2757 1149 2791
rect 1185 2757 1219 2791
rect 1255 2757 1289 2791
rect 1363 2755 1397 2789
rect 1432 2755 1466 2789
rect 1501 2755 1535 2789
rect 1570 2755 1604 2789
rect 1639 2755 1673 2789
rect 1708 2755 1742 2789
rect 1777 2755 1811 2789
rect 1846 2755 1880 2789
rect 1915 2755 1949 2789
rect 1984 2755 2018 2789
rect 2053 2755 2087 2789
rect 2122 2755 2156 2789
rect 2191 2755 2225 2789
rect 2259 2755 2293 2789
rect 2327 2755 2361 2789
rect 2395 2755 2429 2789
rect 2463 2755 2497 2789
rect 2531 2755 2565 2789
rect 2599 2755 2633 2789
rect 2667 2755 2701 2789
rect 2735 2755 2769 2789
rect 2803 2755 2837 2789
rect 2871 2755 2905 2789
rect 2939 2755 2973 2789
rect 3007 2755 3041 2789
rect 3075 2755 3109 2789
rect 169 2697 203 2731
rect 245 2697 279 2731
rect 321 2697 355 2731
rect 410 2683 444 2717
rect 481 2683 515 2717
rect 552 2683 586 2717
rect 623 2683 657 2717
rect 694 2683 728 2717
rect 765 2683 799 2717
rect 835 2683 869 2717
rect 905 2683 939 2717
rect 975 2683 1009 2717
rect 1045 2683 1079 2717
rect 1115 2683 1149 2717
rect 1185 2683 1219 2717
rect 1255 2683 1289 2717
rect 1363 2681 1397 2715
rect 1432 2681 1466 2715
rect 1501 2681 1535 2715
rect 1570 2681 1604 2715
rect 1639 2681 1673 2715
rect 1708 2681 1742 2715
rect 1777 2681 1811 2715
rect 1846 2681 1880 2715
rect 1915 2681 1949 2715
rect 1984 2681 2018 2715
rect 2053 2681 2087 2715
rect 2122 2681 2156 2715
rect 2191 2681 2225 2715
rect 2259 2681 2293 2715
rect 2327 2681 2361 2715
rect 2395 2681 2429 2715
rect 2463 2681 2497 2715
rect 2531 2681 2565 2715
rect 2599 2681 2633 2715
rect 2667 2681 2701 2715
rect 2735 2681 2769 2715
rect 2803 2681 2837 2715
rect 2871 2681 2905 2715
rect 2939 2681 2973 2715
rect 3007 2681 3041 2715
rect 3075 2681 3109 2715
rect 169 2627 203 2661
rect 245 2627 279 2661
rect 321 2627 355 2661
rect 410 2609 444 2643
rect 481 2609 515 2643
rect 552 2609 586 2643
rect 623 2609 657 2643
rect 694 2609 728 2643
rect 765 2609 799 2643
rect 835 2609 869 2643
rect 905 2609 939 2643
rect 975 2609 1009 2643
rect 1045 2609 1079 2643
rect 1115 2609 1149 2643
rect 1185 2609 1219 2643
rect 1255 2609 1289 2643
rect 1363 2607 1397 2641
rect 1432 2607 1466 2641
rect 1501 2607 1535 2641
rect 1570 2607 1604 2641
rect 1639 2607 1673 2641
rect 1708 2607 1742 2641
rect 1777 2607 1811 2641
rect 1846 2607 1880 2641
rect 1915 2607 1949 2641
rect 1984 2607 2018 2641
rect 2053 2607 2087 2641
rect 2122 2607 2156 2641
rect 2191 2607 2225 2641
rect 2259 2607 2293 2641
rect 2327 2607 2361 2641
rect 2395 2607 2429 2641
rect 2463 2607 2497 2641
rect 2531 2607 2565 2641
rect 2599 2607 2633 2641
rect 2667 2607 2701 2641
rect 2735 2607 2769 2641
rect 2803 2607 2837 2641
rect 2871 2607 2905 2641
rect 2939 2607 2973 2641
rect 3007 2607 3041 2641
rect 3075 2607 3109 2641
rect 169 2557 203 2591
rect 245 2557 279 2591
rect 321 2557 355 2591
rect 410 2535 444 2569
rect 481 2535 515 2569
rect 552 2535 586 2569
rect 623 2535 657 2569
rect 694 2535 728 2569
rect 765 2535 799 2569
rect 835 2535 869 2569
rect 905 2535 939 2569
rect 975 2535 1009 2569
rect 1045 2535 1079 2569
rect 1115 2535 1149 2569
rect 1185 2535 1219 2569
rect 1255 2535 1289 2569
rect 1363 2533 1397 2567
rect 1432 2533 1466 2567
rect 1501 2533 1535 2567
rect 1570 2533 1604 2567
rect 1639 2533 1673 2567
rect 1708 2533 1742 2567
rect 1777 2533 1811 2567
rect 1846 2533 1880 2567
rect 1915 2533 1949 2567
rect 1984 2533 2018 2567
rect 2053 2533 2087 2567
rect 2122 2533 2156 2567
rect 2191 2533 2225 2567
rect 2259 2533 2293 2567
rect 2327 2533 2361 2567
rect 2395 2533 2429 2567
rect 2463 2533 2497 2567
rect 2531 2533 2565 2567
rect 2599 2533 2633 2567
rect 2667 2533 2701 2567
rect 2735 2533 2769 2567
rect 2803 2533 2837 2567
rect 2871 2533 2905 2567
rect 2939 2533 2973 2567
rect 3007 2533 3041 2567
rect 3075 2533 3109 2567
rect 25846 1999 25880 2033
rect 25917 1999 25951 2033
rect 25988 1999 26022 2033
rect 26059 1999 26093 2033
rect 26130 1999 26164 2033
rect 26201 1999 26235 2033
rect 26272 1999 26306 2033
rect 26342 1999 26376 2033
rect 26412 1999 26446 2033
rect 26482 1999 26516 2033
rect 26552 1999 26586 2033
rect 26622 1999 26656 2033
rect 26692 1999 26726 2033
rect 26762 1999 26796 2033
rect 26832 1999 26866 2033
rect 26902 1999 26936 2033
rect 26972 1999 27006 2033
rect 27042 1999 27076 2033
rect 27112 1999 27146 2033
rect 27182 1999 27216 2033
rect 27252 1999 27286 2033
rect 27322 1999 27356 2033
rect 27392 1999 27426 2033
rect 27462 1999 27496 2033
rect 27532 1999 27566 2033
rect 27602 1999 27636 2033
rect 27672 1999 27706 2033
rect 27742 1999 27776 2033
rect 27812 1999 27846 2033
rect 25846 1913 25880 1947
rect 25917 1913 25951 1947
rect 25988 1913 26022 1947
rect 26059 1913 26093 1947
rect 26130 1913 26164 1947
rect 26201 1913 26235 1947
rect 26272 1913 26306 1947
rect 26342 1913 26376 1947
rect 26412 1913 26446 1947
rect 26482 1913 26516 1947
rect 26552 1913 26586 1947
rect 26622 1913 26656 1947
rect 26692 1913 26726 1947
rect 26762 1913 26796 1947
rect 26832 1913 26866 1947
rect 26902 1913 26936 1947
rect 26972 1913 27006 1947
rect 27042 1913 27076 1947
rect 27112 1913 27146 1947
rect 27182 1913 27216 1947
rect 27252 1913 27286 1947
rect 27322 1913 27356 1947
rect 27392 1913 27426 1947
rect 27462 1913 27496 1947
rect 27532 1913 27566 1947
rect 27602 1913 27636 1947
rect 27672 1913 27706 1947
rect 27742 1913 27776 1947
rect 27812 1913 27846 1947
rect 25846 1827 25880 1861
rect 25917 1827 25951 1861
rect 25988 1827 26022 1861
rect 26059 1827 26093 1861
rect 26130 1827 26164 1861
rect 26201 1827 26235 1861
rect 26272 1827 26306 1861
rect 26342 1827 26376 1861
rect 26412 1827 26446 1861
rect 26482 1827 26516 1861
rect 26552 1827 26586 1861
rect 26622 1827 26656 1861
rect 26692 1827 26726 1861
rect 26762 1827 26796 1861
rect 26832 1827 26866 1861
rect 26902 1827 26936 1861
rect 26972 1827 27006 1861
rect 27042 1827 27076 1861
rect 27112 1827 27146 1861
rect 27182 1827 27216 1861
rect 27252 1827 27286 1861
rect 27322 1827 27356 1861
rect 27392 1827 27426 1861
rect 27462 1827 27496 1861
rect 27532 1827 27566 1861
rect 27602 1827 27636 1861
rect 27672 1827 27706 1861
rect 27742 1827 27776 1861
rect 27812 1827 27846 1861
rect 25846 1741 25880 1775
rect 25917 1741 25951 1775
rect 25988 1741 26022 1775
rect 26059 1741 26093 1775
rect 26130 1741 26164 1775
rect 26201 1741 26235 1775
rect 26272 1741 26306 1775
rect 26342 1741 26376 1775
rect 26412 1741 26446 1775
rect 26482 1741 26516 1775
rect 26552 1741 26586 1775
rect 26622 1741 26656 1775
rect 26692 1741 26726 1775
rect 26762 1741 26796 1775
rect 26832 1741 26866 1775
rect 26902 1741 26936 1775
rect 26972 1741 27006 1775
rect 27042 1741 27076 1775
rect 27112 1741 27146 1775
rect 27182 1741 27216 1775
rect 27252 1741 27286 1775
rect 27322 1741 27356 1775
rect 27392 1741 27426 1775
rect 27462 1741 27496 1775
rect 27532 1741 27566 1775
rect 27602 1741 27636 1775
rect 27672 1741 27706 1775
rect 27742 1741 27776 1775
rect 27812 1741 27846 1775
<< mvnsubdiffcont >>
rect 2401 20716 2435 20750
rect 2474 20716 2508 20750
rect 2547 20716 2581 20750
rect 2620 20716 2654 20750
rect 2693 20716 2727 20750
rect 2766 20716 2800 20750
rect 2839 20716 2873 20750
rect 2912 20716 2946 20750
rect 2984 20716 3018 20750
rect 3056 20716 3090 20750
rect 3128 20716 3162 20750
rect 2401 20638 2435 20672
rect 2474 20638 2508 20672
rect 2547 20638 2581 20672
rect 2620 20638 2654 20672
rect 2693 20638 2727 20672
rect 2766 20638 2800 20672
rect 2839 20638 2873 20672
rect 2912 20638 2946 20672
rect 2984 20638 3018 20672
rect 3056 20638 3090 20672
rect 3128 20638 3162 20672
rect 2401 20560 2435 20594
rect 2474 20560 2508 20594
rect 2547 20560 2581 20594
rect 2620 20560 2654 20594
rect 2693 20560 2727 20594
rect 2766 20560 2800 20594
rect 2839 20560 2873 20594
rect 2912 20560 2946 20594
rect 2984 20560 3018 20594
rect 3056 20560 3090 20594
rect 3128 20560 3162 20594
rect 2401 20482 2435 20516
rect 2474 20482 2508 20516
rect 2547 20482 2581 20516
rect 2620 20482 2654 20516
rect 2693 20482 2727 20516
rect 2766 20482 2800 20516
rect 2839 20482 2873 20516
rect 2912 20482 2946 20516
rect 2984 20482 3018 20516
rect 3056 20482 3090 20516
rect 3128 20482 3162 20516
rect 2401 20404 2435 20438
rect 2474 20404 2508 20438
rect 2547 20404 2581 20438
rect 2620 20404 2654 20438
rect 2693 20404 2727 20438
rect 2766 20404 2800 20438
rect 2839 20404 2873 20438
rect 2912 20404 2946 20438
rect 2984 20404 3018 20438
rect 3056 20404 3090 20438
rect 3128 20404 3162 20438
rect 26371 20684 26405 20718
rect 26441 20684 26475 20718
rect 26511 20684 26545 20718
rect 26581 20684 26615 20718
rect 26651 20684 26685 20718
rect 26721 20684 26755 20718
rect 26791 20684 26825 20718
rect 26861 20684 26895 20718
rect 26371 20613 26405 20647
rect 26441 20613 26475 20647
rect 26511 20613 26545 20647
rect 26581 20613 26615 20647
rect 26651 20613 26685 20647
rect 26721 20613 26755 20647
rect 26791 20613 26825 20647
rect 26861 20613 26895 20647
rect 26371 20542 26405 20576
rect 26441 20542 26475 20576
rect 26511 20542 26545 20576
rect 26581 20542 26615 20576
rect 26651 20542 26685 20576
rect 26721 20542 26755 20576
rect 26791 20542 26825 20576
rect 26861 20542 26895 20576
rect 26371 20471 26405 20505
rect 26441 20471 26475 20505
rect 26511 20471 26545 20505
rect 26581 20471 26615 20505
rect 26651 20471 26685 20505
rect 26721 20471 26755 20505
rect 26791 20471 26825 20505
rect 26861 20471 26895 20505
rect 26371 20400 26405 20434
rect 26441 20400 26475 20434
rect 26511 20400 26545 20434
rect 26581 20400 26615 20434
rect 26651 20400 26685 20434
rect 26721 20400 26755 20434
rect 26791 20400 26825 20434
rect 26861 20400 26895 20434
rect 26371 20329 26405 20363
rect 26441 20329 26475 20363
rect 26511 20329 26545 20363
rect 26581 20329 26615 20363
rect 26651 20329 26685 20363
rect 26721 20329 26755 20363
rect 26791 20329 26825 20363
rect 26861 20329 26895 20363
rect 26371 20258 26405 20292
rect 26441 20258 26475 20292
rect 26511 20258 26545 20292
rect 26581 20258 26615 20292
rect 26651 20258 26685 20292
rect 26721 20258 26755 20292
rect 26791 20258 26825 20292
rect 26861 20258 26895 20292
rect 26371 20187 26405 20221
rect 26441 20187 26475 20221
rect 26511 20187 26545 20221
rect 26581 20187 26615 20221
rect 26651 20187 26685 20221
rect 26721 20187 26755 20221
rect 26791 20187 26825 20221
rect 26861 20187 26895 20221
rect 26371 20116 26405 20150
rect 26441 20116 26475 20150
rect 26511 20116 26545 20150
rect 26581 20116 26615 20150
rect 26651 20116 26685 20150
rect 26721 20116 26755 20150
rect 26791 20116 26825 20150
rect 26861 20116 26895 20150
rect 26371 20044 26405 20078
rect 26441 20044 26475 20078
rect 26511 20044 26545 20078
rect 26581 20044 26615 20078
rect 26651 20044 26685 20078
rect 26721 20044 26755 20078
rect 26791 20044 26825 20078
rect 26861 20044 26895 20078
rect 3485 19517 3519 19551
rect 3561 19517 3595 19551
rect 3637 19517 3671 19551
rect 3713 19517 3747 19551
rect 3789 19517 3823 19551
rect 3865 19517 3899 19551
rect 3941 19517 3975 19551
rect 4017 19517 4051 19551
rect 3485 19449 3519 19483
rect 3561 19449 3595 19483
rect 3637 19449 3671 19483
rect 3713 19449 3747 19483
rect 3789 19449 3823 19483
rect 3865 19449 3899 19483
rect 3941 19449 3975 19483
rect 4017 19449 4051 19483
rect 3485 19381 3519 19415
rect 3561 19381 3595 19415
rect 3637 19381 3671 19415
rect 3713 19381 3747 19415
rect 3789 19381 3823 19415
rect 3865 19381 3899 19415
rect 3941 19381 3975 19415
rect 4017 19381 4051 19415
rect 3485 19313 3519 19347
rect 3561 19313 3595 19347
rect 3637 19313 3671 19347
rect 3713 19313 3747 19347
rect 3789 19313 3823 19347
rect 3865 19313 3899 19347
rect 3941 19313 3975 19347
rect 4017 19313 4051 19347
rect 3485 19245 3519 19279
rect 3561 19245 3595 19279
rect 3637 19245 3671 19279
rect 3713 19245 3747 19279
rect 3789 19245 3823 19279
rect 3865 19245 3899 19279
rect 3941 19245 3975 19279
rect 4017 19245 4051 19279
rect 3485 19176 3519 19210
rect 3561 19176 3595 19210
rect 3637 19176 3671 19210
rect 3713 19176 3747 19210
rect 3789 19176 3823 19210
rect 3865 19176 3899 19210
rect 3941 19176 3975 19210
rect 4017 19176 4051 19210
rect 3485 19107 3519 19141
rect 3561 19107 3595 19141
rect 3637 19107 3671 19141
rect 3713 19107 3747 19141
rect 3789 19107 3823 19141
rect 3865 19107 3899 19141
rect 3941 19107 3975 19141
rect 4017 19107 4051 19141
rect 3485 19038 3519 19072
rect 3561 19038 3595 19072
rect 3637 19038 3671 19072
rect 3713 19038 3747 19072
rect 3789 19038 3823 19072
rect 3865 19038 3899 19072
rect 3941 19038 3975 19072
rect 4017 19038 4051 19072
rect 3485 18969 3519 19003
rect 3561 18969 3595 19003
rect 3637 18969 3671 19003
rect 3713 18969 3747 19003
rect 3789 18969 3823 19003
rect 3865 18969 3899 19003
rect 3941 18969 3975 19003
rect 4017 18969 4051 19003
rect 3485 18900 3519 18934
rect 3561 18900 3595 18934
rect 3637 18900 3671 18934
rect 3713 18900 3747 18934
rect 3789 18900 3823 18934
rect 3865 18900 3899 18934
rect 3941 18900 3975 18934
rect 4017 18900 4051 18934
rect 3485 18831 3519 18865
rect 3561 18831 3595 18865
rect 3637 18831 3671 18865
rect 3713 18831 3747 18865
rect 3789 18831 3823 18865
rect 3865 18831 3899 18865
rect 3941 18831 3975 18865
rect 4017 18831 4051 18865
rect 3485 18762 3519 18796
rect 3561 18762 3595 18796
rect 3637 18762 3671 18796
rect 3713 18762 3747 18796
rect 3789 18762 3823 18796
rect 3865 18762 3899 18796
rect 3941 18762 3975 18796
rect 4017 18762 4051 18796
rect 3485 18693 3519 18727
rect 3561 18693 3595 18727
rect 3637 18693 3671 18727
rect 3713 18693 3747 18727
rect 3789 18693 3823 18727
rect 3865 18693 3899 18727
rect 3941 18693 3975 18727
rect 4017 18693 4051 18727
rect 3485 18624 3519 18658
rect 3561 18624 3595 18658
rect 3637 18624 3671 18658
rect 3713 18624 3747 18658
rect 3789 18624 3823 18658
rect 3865 18624 3899 18658
rect 3941 18624 3975 18658
rect 4017 18624 4051 18658
rect 3485 18555 3519 18589
rect 3561 18555 3595 18589
rect 3637 18555 3671 18589
rect 3713 18555 3747 18589
rect 3789 18555 3823 18589
rect 3865 18555 3899 18589
rect 3941 18555 3975 18589
rect 4017 18555 4051 18589
rect 3485 18486 3519 18520
rect 3561 18486 3595 18520
rect 3637 18486 3671 18520
rect 3713 18486 3747 18520
rect 3789 18486 3823 18520
rect 3865 18486 3899 18520
rect 3941 18486 3975 18520
rect 4017 18486 4051 18520
rect 3485 18417 3519 18451
rect 3561 18417 3595 18451
rect 3637 18417 3671 18451
rect 3713 18417 3747 18451
rect 3789 18417 3823 18451
rect 3865 18417 3899 18451
rect 3941 18417 3975 18451
rect 4017 18417 4051 18451
rect 3485 18348 3519 18382
rect 3561 18348 3595 18382
rect 3637 18348 3671 18382
rect 3713 18348 3747 18382
rect 3789 18348 3823 18382
rect 3865 18348 3899 18382
rect 3941 18348 3975 18382
rect 4017 18348 4051 18382
rect 3485 18279 3519 18313
rect 3561 18279 3595 18313
rect 3637 18279 3671 18313
rect 3713 18279 3747 18313
rect 3789 18279 3823 18313
rect 3865 18279 3899 18313
rect 3941 18279 3975 18313
rect 4017 18279 4051 18313
rect 3485 18210 3519 18244
rect 3561 18210 3595 18244
rect 3637 18210 3671 18244
rect 3713 18210 3747 18244
rect 3789 18210 3823 18244
rect 3865 18210 3899 18244
rect 3941 18210 3975 18244
rect 4017 18210 4051 18244
rect 3485 18141 3519 18175
rect 3561 18141 3595 18175
rect 3637 18141 3671 18175
rect 3713 18141 3747 18175
rect 3789 18141 3823 18175
rect 3865 18141 3899 18175
rect 3941 18141 3975 18175
rect 4017 18141 4051 18175
rect 3485 18072 3519 18106
rect 3561 18072 3595 18106
rect 3637 18072 3671 18106
rect 3713 18072 3747 18106
rect 3789 18072 3823 18106
rect 3865 18072 3899 18106
rect 3941 18072 3975 18106
rect 4017 18072 4051 18106
rect 3485 18003 3519 18037
rect 3561 18003 3595 18037
rect 3637 18003 3671 18037
rect 3713 18003 3747 18037
rect 3789 18003 3823 18037
rect 3865 18003 3899 18037
rect 3941 18003 3975 18037
rect 4017 18003 4051 18037
rect 3485 17934 3519 17968
rect 3561 17934 3595 17968
rect 3637 17934 3671 17968
rect 3713 17934 3747 17968
rect 3789 17934 3823 17968
rect 3865 17934 3899 17968
rect 3941 17934 3975 17968
rect 4017 17934 4051 17968
rect 3485 17865 3519 17899
rect 3561 17865 3595 17899
rect 3637 17865 3671 17899
rect 3713 17865 3747 17899
rect 3789 17865 3823 17899
rect 3865 17865 3899 17899
rect 3941 17865 3975 17899
rect 4017 17865 4051 17899
rect 3485 17796 3519 17830
rect 3561 17796 3595 17830
rect 3637 17796 3671 17830
rect 3713 17796 3747 17830
rect 3789 17796 3823 17830
rect 3865 17796 3899 17830
rect 3941 17796 3975 17830
rect 4017 17796 4051 17830
rect 3485 17727 3519 17761
rect 3561 17727 3595 17761
rect 3637 17727 3671 17761
rect 3713 17727 3747 17761
rect 3789 17727 3823 17761
rect 3865 17727 3899 17761
rect 3941 17727 3975 17761
rect 4017 17727 4051 17761
rect 3485 17658 3519 17692
rect 3561 17658 3595 17692
rect 3637 17658 3671 17692
rect 3713 17658 3747 17692
rect 3789 17658 3823 17692
rect 3865 17658 3899 17692
rect 3941 17658 3975 17692
rect 4017 17658 4051 17692
rect 3485 17589 3519 17623
rect 3561 17589 3595 17623
rect 3637 17589 3671 17623
rect 3713 17589 3747 17623
rect 3789 17589 3823 17623
rect 3865 17589 3899 17623
rect 3941 17589 3975 17623
rect 4017 17589 4051 17623
rect 3485 17520 3519 17554
rect 3561 17520 3595 17554
rect 3637 17520 3671 17554
rect 3713 17520 3747 17554
rect 3789 17520 3823 17554
rect 3865 17520 3899 17554
rect 3941 17520 3975 17554
rect 4017 17520 4051 17554
rect 3485 17451 3519 17485
rect 3561 17451 3595 17485
rect 3637 17451 3671 17485
rect 3713 17451 3747 17485
rect 3789 17451 3823 17485
rect 3865 17451 3899 17485
rect 3941 17451 3975 17485
rect 4017 17451 4051 17485
rect 3485 17382 3519 17416
rect 3561 17382 3595 17416
rect 3637 17382 3671 17416
rect 3713 17382 3747 17416
rect 3789 17382 3823 17416
rect 3865 17382 3899 17416
rect 3941 17382 3975 17416
rect 4017 17382 4051 17416
rect 3485 17313 3519 17347
rect 3561 17313 3595 17347
rect 3637 17313 3671 17347
rect 3713 17313 3747 17347
rect 3789 17313 3823 17347
rect 3865 17313 3899 17347
rect 3941 17313 3975 17347
rect 4017 17313 4051 17347
rect 3485 17244 3519 17278
rect 3561 17244 3595 17278
rect 3637 17244 3671 17278
rect 3713 17244 3747 17278
rect 3789 17244 3823 17278
rect 3865 17244 3899 17278
rect 3941 17244 3975 17278
rect 4017 17244 4051 17278
rect 3485 17175 3519 17209
rect 3561 17175 3595 17209
rect 3637 17175 3671 17209
rect 3713 17175 3747 17209
rect 3789 17175 3823 17209
rect 3865 17175 3899 17209
rect 3941 17175 3975 17209
rect 4017 17175 4051 17209
rect 3485 17106 3519 17140
rect 3561 17106 3595 17140
rect 3637 17106 3671 17140
rect 3713 17106 3747 17140
rect 3789 17106 3823 17140
rect 3865 17106 3899 17140
rect 3941 17106 3975 17140
rect 4017 17106 4051 17140
rect 3767 17013 3801 17047
rect 3835 17013 3869 17047
rect 3903 17013 3937 17047
rect 3971 17013 4005 17047
rect 4039 17013 4073 17047
rect 3767 16939 3801 16973
rect 3835 16939 3869 16973
rect 3903 16939 3937 16973
rect 3971 16939 4005 16973
rect 4039 16939 4073 16973
rect 3767 16865 3801 16899
rect 3835 16865 3869 16899
rect 3903 16865 3937 16899
rect 3971 16865 4005 16899
rect 4039 16865 4073 16899
rect 3767 16791 3801 16825
rect 3835 16791 3869 16825
rect 3903 16791 3937 16825
rect 3971 16791 4005 16825
rect 4039 16791 4073 16825
rect 3767 16717 3801 16751
rect 3835 16717 3869 16751
rect 3903 16717 3937 16751
rect 3971 16717 4005 16751
rect 4039 16717 4073 16751
rect 3767 16643 3801 16677
rect 3835 16643 3869 16677
rect 3903 16643 3937 16677
rect 3971 16643 4005 16677
rect 4039 16643 4073 16677
rect 3767 16569 3801 16603
rect 3835 16569 3869 16603
rect 3903 16569 3937 16603
rect 3971 16569 4005 16603
rect 4039 16569 4073 16603
rect 3767 16495 3801 16529
rect 3835 16495 3869 16529
rect 3903 16495 3937 16529
rect 3971 16495 4005 16529
rect 4039 16495 4073 16529
rect 3767 16421 3801 16455
rect 3835 16421 3869 16455
rect 3903 16421 3937 16455
rect 3971 16421 4005 16455
rect 4039 16421 4073 16455
rect 3767 16346 3801 16380
rect 3835 16346 3869 16380
rect 3903 16346 3937 16380
rect 3971 16346 4005 16380
rect 4039 16346 4073 16380
rect 2950 16226 2984 16260
rect 3018 16226 3052 16260
rect 3086 16226 3120 16260
rect 3154 16226 3188 16260
rect 3222 16226 3256 16260
rect 3290 16226 3324 16260
rect 3358 16226 3392 16260
rect 3426 16226 3460 16260
rect 3494 16226 3528 16260
rect 3562 16226 3596 16260
rect 3630 16226 3664 16260
rect 3698 16226 3732 16260
rect 2950 16154 2984 16188
rect 3018 16154 3052 16188
rect 3086 16154 3120 16188
rect 3154 16154 3188 16188
rect 3222 16154 3256 16188
rect 3290 16154 3324 16188
rect 3358 16154 3392 16188
rect 3426 16154 3460 16188
rect 3494 16154 3528 16188
rect 3562 16154 3596 16188
rect 3630 16154 3664 16188
rect 3698 16154 3732 16188
rect 2950 16082 2984 16116
rect 3018 16082 3052 16116
rect 3086 16082 3120 16116
rect 3154 16082 3188 16116
rect 3222 16082 3256 16116
rect 3290 16082 3324 16116
rect 3358 16082 3392 16116
rect 3426 16082 3460 16116
rect 3494 16082 3528 16116
rect 3562 16082 3596 16116
rect 3630 16082 3664 16116
rect 3698 16082 3732 16116
rect 2950 16010 2984 16044
rect 3018 16010 3052 16044
rect 3086 16010 3120 16044
rect 3154 16010 3188 16044
rect 3222 16010 3256 16044
rect 3290 16010 3324 16044
rect 3358 16010 3392 16044
rect 3426 16010 3460 16044
rect 3494 16010 3528 16044
rect 3562 16010 3596 16044
rect 3630 16010 3664 16044
rect 3698 16010 3732 16044
rect 2950 15938 2984 15972
rect 3018 15938 3052 15972
rect 3086 15938 3120 15972
rect 3154 15938 3188 15972
rect 3222 15938 3256 15972
rect 3290 15938 3324 15972
rect 3358 15938 3392 15972
rect 3426 15938 3460 15972
rect 3494 15938 3528 15972
rect 3562 15938 3596 15972
rect 3630 15938 3664 15972
rect 3698 15938 3732 15972
rect 2950 15866 2984 15900
rect 3018 15866 3052 15900
rect 3086 15866 3120 15900
rect 3154 15866 3188 15900
rect 3222 15866 3256 15900
rect 3290 15866 3324 15900
rect 3358 15866 3392 15900
rect 3426 15866 3460 15900
rect 3494 15866 3528 15900
rect 3562 15866 3596 15900
rect 3630 15866 3664 15900
rect 3698 15866 3732 15900
rect 2950 15794 2984 15828
rect 3018 15794 3052 15828
rect 3086 15794 3120 15828
rect 3154 15794 3188 15828
rect 3222 15794 3256 15828
rect 3290 15794 3324 15828
rect 3358 15794 3392 15828
rect 3426 15794 3460 15828
rect 3494 15794 3528 15828
rect 3562 15794 3596 15828
rect 3630 15794 3664 15828
rect 3698 15794 3732 15828
rect 2950 15722 2984 15756
rect 3018 15722 3052 15756
rect 3086 15722 3120 15756
rect 3154 15722 3188 15756
rect 3222 15722 3256 15756
rect 3290 15722 3324 15756
rect 3358 15722 3392 15756
rect 3426 15722 3460 15756
rect 3494 15722 3528 15756
rect 3562 15722 3596 15756
rect 3630 15722 3664 15756
rect 3698 15722 3732 15756
rect 2950 15650 2984 15684
rect 3018 15650 3052 15684
rect 3086 15650 3120 15684
rect 3154 15650 3188 15684
rect 3222 15650 3256 15684
rect 3290 15650 3324 15684
rect 3358 15650 3392 15684
rect 3426 15650 3460 15684
rect 3494 15650 3528 15684
rect 3562 15650 3596 15684
rect 3630 15650 3664 15684
rect 3698 15650 3732 15684
rect 2950 15578 2984 15612
rect 3018 15578 3052 15612
rect 3086 15578 3120 15612
rect 3154 15578 3188 15612
rect 3222 15578 3256 15612
rect 3290 15578 3324 15612
rect 3358 15578 3392 15612
rect 3426 15578 3460 15612
rect 3494 15578 3528 15612
rect 3562 15578 3596 15612
rect 3630 15578 3664 15612
rect 3698 15578 3732 15612
rect 2950 15506 2984 15540
rect 3018 15506 3052 15540
rect 3086 15506 3120 15540
rect 3154 15506 3188 15540
rect 3222 15506 3256 15540
rect 3290 15506 3324 15540
rect 3358 15506 3392 15540
rect 3426 15506 3460 15540
rect 3494 15506 3528 15540
rect 3562 15506 3596 15540
rect 3630 15506 3664 15540
rect 3698 15506 3732 15540
rect 2950 15434 2984 15468
rect 3018 15434 3052 15468
rect 3086 15434 3120 15468
rect 3154 15434 3188 15468
rect 3222 15434 3256 15468
rect 3290 15434 3324 15468
rect 3358 15434 3392 15468
rect 3426 15434 3460 15468
rect 3494 15434 3528 15468
rect 3562 15434 3596 15468
rect 3630 15434 3664 15468
rect 3698 15434 3732 15468
rect 7858 16244 7892 16278
rect 7934 16244 7968 16278
rect 8010 16244 8044 16278
rect 8086 16244 8120 16278
rect 8162 16244 8196 16278
rect 8238 16244 8272 16278
rect 7858 16175 7892 16209
rect 7934 16175 7968 16209
rect 8010 16175 8044 16209
rect 8086 16175 8120 16209
rect 8162 16175 8196 16209
rect 8238 16175 8272 16209
rect 7858 16106 7892 16140
rect 7934 16106 7968 16140
rect 8010 16106 8044 16140
rect 8086 16106 8120 16140
rect 8162 16106 8196 16140
rect 8238 16106 8272 16140
rect 7858 16037 7892 16071
rect 7934 16037 7968 16071
rect 8010 16037 8044 16071
rect 8086 16037 8120 16071
rect 8162 16037 8196 16071
rect 8238 16037 8272 16071
rect 7858 15968 7892 16002
rect 7934 15968 7968 16002
rect 8010 15968 8044 16002
rect 8086 15968 8120 16002
rect 8162 15968 8196 16002
rect 8238 15968 8272 16002
rect 7858 15899 7892 15933
rect 7934 15899 7968 15933
rect 8010 15899 8044 15933
rect 8086 15899 8120 15933
rect 8162 15899 8196 15933
rect 8238 15899 8272 15933
rect 7858 15830 7892 15864
rect 7934 15830 7968 15864
rect 8010 15830 8044 15864
rect 8086 15830 8120 15864
rect 8162 15830 8196 15864
rect 8238 15830 8272 15864
rect 7858 15761 7892 15795
rect 7934 15761 7968 15795
rect 8010 15761 8044 15795
rect 8086 15761 8120 15795
rect 8162 15761 8196 15795
rect 8238 15761 8272 15795
rect 7858 15692 7892 15726
rect 7934 15692 7968 15726
rect 8010 15692 8044 15726
rect 8086 15692 8120 15726
rect 8162 15692 8196 15726
rect 8238 15692 8272 15726
rect 7858 15623 7892 15657
rect 7934 15623 7968 15657
rect 8010 15623 8044 15657
rect 8086 15623 8120 15657
rect 8162 15623 8196 15657
rect 8238 15623 8272 15657
rect 7858 15554 7892 15588
rect 7934 15554 7968 15588
rect 8010 15554 8044 15588
rect 8086 15554 8120 15588
rect 8162 15554 8196 15588
rect 8238 15554 8272 15588
rect 7858 15485 7892 15519
rect 7934 15485 7968 15519
rect 8010 15485 8044 15519
rect 8086 15485 8120 15519
rect 8162 15485 8196 15519
rect 8238 15485 8272 15519
rect 7858 15415 7892 15449
rect 7934 15415 7968 15449
rect 8010 15415 8044 15449
rect 8086 15415 8120 15449
rect 8162 15415 8196 15449
rect 8238 15415 8272 15449
<< locali >>
rect 76 39912 232 39924
rect 76 39900 92 39912
rect 126 39878 174 39912
rect 208 39900 232 39912
rect 110 39866 198 39878
rect 76 39840 232 39866
rect 76 39831 92 39840
rect 126 39806 174 39840
rect 208 39831 232 39840
rect 110 39797 198 39806
rect 76 39768 232 39797
rect 76 39762 92 39768
rect 126 39734 174 39768
rect 208 39762 232 39768
rect 110 39728 198 39734
rect 76 39696 232 39728
rect 76 39693 92 39696
rect 126 39662 174 39696
rect 208 39693 232 39696
rect 110 39659 198 39662
rect 76 39624 232 39659
rect 126 39590 174 39624
rect 76 39555 232 39590
rect 110 39552 198 39555
rect 76 39518 92 39521
rect 126 39518 174 39552
rect 208 39518 232 39521
rect 76 39486 232 39518
rect 110 39480 198 39486
rect 76 39446 92 39452
rect 126 39446 174 39480
rect 208 39446 232 39452
rect 76 39417 232 39446
rect 110 39408 198 39417
rect 76 39374 92 39383
rect 126 39374 174 39408
rect 208 39374 232 39383
rect 76 39348 232 39374
rect 110 39336 198 39348
rect 76 39302 92 39314
rect 126 39302 174 39336
rect 208 39302 232 39314
rect 76 39279 232 39302
rect 110 39264 198 39279
rect 76 39230 92 39245
rect 126 39230 174 39264
rect 208 39230 232 39245
rect 76 39209 232 39230
rect 110 39192 198 39209
rect 76 39158 92 39175
rect 126 39158 174 39192
rect 208 39158 232 39175
rect 76 39139 232 39158
rect 110 39120 198 39139
rect 76 39086 92 39105
rect 126 39086 174 39120
rect 208 39086 232 39105
rect 76 39069 232 39086
rect 110 39048 198 39069
rect 76 39014 92 39035
rect 126 39014 174 39048
rect 208 39014 232 39035
rect 76 38999 232 39014
rect 110 38976 198 38999
rect 76 38942 92 38965
rect 126 38942 174 38976
rect 208 38942 232 38965
rect 76 38929 232 38942
rect 110 38904 198 38929
rect 76 38870 92 38895
rect 126 38870 174 38904
rect 208 38870 232 38895
rect 76 38859 232 38870
rect 110 38832 198 38859
rect 76 38798 92 38825
rect 126 38798 174 38832
rect 208 38798 232 38825
rect 76 38789 232 38798
rect 110 38760 198 38789
rect 76 38726 92 38755
rect 126 38726 174 38760
rect 208 38726 232 38755
rect 76 38719 232 38726
rect 110 38688 198 38719
rect 76 38654 92 38685
rect 126 38654 174 38688
rect 208 38654 232 38685
rect 76 38649 232 38654
rect 110 38616 198 38649
rect 76 38582 92 38615
rect 126 38582 174 38616
rect 208 38582 232 38615
rect 76 38579 232 38582
rect 110 38545 198 38579
rect 76 38544 232 38545
rect 76 38510 92 38544
rect 126 38510 174 38544
rect 208 38510 232 38544
rect 76 38509 232 38510
rect 110 38475 198 38509
rect 76 38472 232 38475
rect 76 38439 92 38472
rect 126 38438 174 38472
rect 208 38439 232 38472
rect 110 38405 198 38438
rect 76 38400 232 38405
rect 76 38369 92 38400
rect 126 38366 174 38400
rect 208 38369 232 38400
rect 110 38335 198 38366
rect 76 38328 232 38335
rect 76 38299 92 38328
rect 126 38294 174 38328
rect 208 38299 232 38328
rect 110 38265 198 38294
rect 76 38256 232 38265
rect 76 38229 92 38256
rect 126 38222 174 38256
rect 208 38229 232 38256
rect 110 38195 198 38222
rect 76 38184 232 38195
rect 76 38159 92 38184
rect 126 38150 174 38184
rect 208 38159 232 38184
rect 110 38125 198 38150
rect 76 38111 232 38125
rect 76 38089 92 38111
rect 126 38077 174 38111
rect 208 38089 232 38111
rect 110 38055 198 38077
rect 76 38038 232 38055
rect 76 38031 92 38038
rect 126 38004 174 38038
rect 208 38031 232 38038
rect 203 37804 331 37836
rect 203 37770 209 37804
rect 243 37770 291 37804
rect 325 37770 331 37804
rect 203 37732 331 37770
rect 203 37698 209 37732
rect 243 37698 291 37732
rect 325 37698 331 37732
rect 203 37660 331 37698
rect 203 37626 209 37660
rect 243 37626 291 37660
rect 325 37626 331 37660
rect 203 37588 331 37626
rect 203 37554 209 37588
rect 243 37554 291 37588
rect 325 37554 331 37588
rect 203 37516 331 37554
rect 24069 37674 27021 37677
rect 24069 37640 24093 37674
rect 24127 37640 24162 37674
rect 24196 37640 24231 37674
rect 24265 37640 24300 37674
rect 24334 37640 24369 37674
rect 24403 37640 24438 37674
rect 24472 37640 24507 37674
rect 24541 37640 24576 37674
rect 24610 37640 24645 37674
rect 24679 37640 24714 37674
rect 24748 37640 24783 37674
rect 24817 37640 24852 37674
rect 24886 37640 24921 37674
rect 24955 37640 24990 37674
rect 25024 37640 25059 37674
rect 25093 37640 25127 37674
rect 25161 37640 25195 37674
rect 25229 37640 25263 37674
rect 25297 37640 25331 37674
rect 25365 37640 25399 37674
rect 25433 37640 25467 37674
rect 25501 37640 25535 37674
rect 25569 37640 25603 37674
rect 25637 37640 25671 37674
rect 25705 37640 25739 37674
rect 25773 37640 25807 37674
rect 25841 37640 25875 37674
rect 25909 37640 25943 37674
rect 25977 37640 26011 37674
rect 26045 37640 26079 37674
rect 26113 37640 26147 37674
rect 26181 37640 26215 37674
rect 26249 37640 26283 37674
rect 26317 37640 26351 37674
rect 26385 37640 26419 37674
rect 26453 37640 26487 37674
rect 26521 37640 26555 37674
rect 26589 37640 26623 37674
rect 26657 37640 26691 37674
rect 26725 37640 26759 37674
rect 26793 37640 26827 37674
rect 26861 37640 26895 37674
rect 26929 37640 26963 37674
rect 26997 37640 27021 37674
rect 24069 37596 27021 37640
rect 24069 37562 24093 37596
rect 24127 37562 24162 37596
rect 24196 37562 24231 37596
rect 24265 37562 24300 37596
rect 24334 37562 24369 37596
rect 24403 37562 24438 37596
rect 24472 37562 24507 37596
rect 24541 37562 24576 37596
rect 24610 37562 24645 37596
rect 24679 37562 24714 37596
rect 24748 37562 24783 37596
rect 24817 37562 24852 37596
rect 24886 37562 24921 37596
rect 24955 37562 24990 37596
rect 25024 37562 25059 37596
rect 25093 37562 25127 37596
rect 25161 37562 25195 37596
rect 25229 37562 25263 37596
rect 25297 37562 25331 37596
rect 25365 37562 25399 37596
rect 25433 37562 25467 37596
rect 25501 37562 25535 37596
rect 25569 37562 25603 37596
rect 25637 37562 25671 37596
rect 25705 37562 25739 37596
rect 25773 37562 25807 37596
rect 25841 37562 25875 37596
rect 25909 37562 25943 37596
rect 25977 37562 26011 37596
rect 26045 37562 26079 37596
rect 26113 37562 26147 37596
rect 26181 37562 26215 37596
rect 26249 37562 26283 37596
rect 26317 37562 26351 37596
rect 26385 37562 26419 37596
rect 26453 37562 26487 37596
rect 26521 37562 26555 37596
rect 26589 37562 26623 37596
rect 26657 37562 26691 37596
rect 26725 37562 26759 37596
rect 26793 37562 26827 37596
rect 26861 37562 26895 37596
rect 26929 37562 26963 37596
rect 26997 37562 27021 37596
rect 24069 37541 27021 37562
rect 203 37482 209 37516
rect 243 37484 291 37516
rect 325 37508 331 37516
rect 22823 37540 27021 37541
rect 22823 37517 23711 37540
rect 325 37484 339 37508
rect 253 37482 291 37484
rect 203 37450 219 37482
rect 253 37450 305 37482
rect 203 37444 339 37450
rect 203 37410 209 37444
rect 243 37415 291 37444
rect 325 37415 339 37444
rect 253 37410 291 37415
rect 203 37381 219 37410
rect 253 37381 305 37410
rect 203 37372 339 37381
rect 203 37338 209 37372
rect 243 37346 291 37372
rect 325 37346 339 37372
rect 253 37338 291 37346
rect 203 37312 219 37338
rect 253 37312 305 37338
rect 203 37300 339 37312
rect 203 37266 209 37300
rect 243 37277 291 37300
rect 325 37277 339 37300
rect 253 37266 291 37277
rect 203 37243 219 37266
rect 253 37243 305 37266
rect 203 37228 339 37243
rect 203 37194 209 37228
rect 243 37208 291 37228
rect 325 37208 339 37228
rect 253 37194 291 37208
rect 203 37174 219 37194
rect 253 37174 305 37194
rect 203 37156 339 37174
rect 203 37122 209 37156
rect 243 37139 291 37156
rect 325 37139 339 37156
rect 253 37122 291 37139
rect 203 37105 219 37122
rect 253 37105 305 37122
rect 203 37084 339 37105
rect 203 37050 209 37084
rect 243 37070 291 37084
rect 325 37070 339 37084
rect 253 37050 291 37070
rect 203 37036 219 37050
rect 253 37036 305 37050
rect 203 37012 339 37036
rect 203 36978 209 37012
rect 243 37001 291 37012
rect 325 37001 339 37012
rect 253 36978 291 37001
rect 203 36967 219 36978
rect 253 36967 305 36978
rect 203 36940 339 36967
rect 203 36906 209 36940
rect 243 36932 291 36940
rect 325 36932 339 36940
rect 253 36906 291 36932
rect 203 36898 219 36906
rect 253 36898 305 36906
rect 203 36868 339 36898
rect 203 36834 209 36868
rect 243 36863 291 36868
rect 325 36863 339 36868
rect 253 36834 291 36863
rect 203 36829 219 36834
rect 253 36829 305 36834
rect 203 36796 339 36829
rect 203 36762 209 36796
rect 243 36794 291 36796
rect 325 36794 339 36796
rect 253 36762 291 36794
rect 203 36760 219 36762
rect 253 36760 305 36762
rect 203 36725 339 36760
rect 203 36724 219 36725
rect 253 36724 305 36725
rect 203 36690 209 36724
rect 253 36691 291 36724
rect 243 36690 291 36691
rect 325 36690 339 36691
rect 203 36655 339 36690
rect 203 36652 219 36655
rect 253 36652 305 36655
rect 203 36618 209 36652
rect 253 36621 291 36652
rect 243 36618 291 36621
rect 325 36618 339 36621
rect 203 36585 339 36618
rect 203 36580 219 36585
rect 253 36580 305 36585
rect 203 36546 209 36580
rect 253 36551 291 36580
rect 243 36546 291 36551
rect 325 36546 339 36551
rect 203 36515 339 36546
rect 203 36508 219 36515
rect 253 36508 305 36515
rect 203 36474 209 36508
rect 253 36481 291 36508
rect 243 36474 291 36481
rect 325 36474 339 36481
rect 203 36445 339 36474
rect 203 36436 219 36445
rect 253 36436 305 36445
rect 203 36402 209 36436
rect 253 36411 291 36436
rect 243 36402 291 36411
rect 325 36402 339 36411
rect 203 36375 339 36402
rect 203 36364 219 36375
rect 253 36364 305 36375
rect 203 36330 209 36364
rect 253 36341 291 36364
rect 243 36330 291 36341
rect 325 36330 339 36341
rect 203 36305 339 36330
rect 203 36292 219 36305
rect 253 36292 305 36305
rect 203 36258 209 36292
rect 253 36271 291 36292
rect 243 36258 291 36271
rect 325 36258 339 36271
rect 203 36235 339 36258
rect 203 36220 219 36235
rect 253 36220 305 36235
rect 203 36186 209 36220
rect 253 36201 291 36220
rect 243 36186 291 36201
rect 325 36186 339 36201
rect 203 36165 339 36186
rect 203 36148 219 36165
rect 253 36148 305 36165
rect 203 36114 209 36148
rect 253 36131 291 36148
rect 243 36114 291 36131
rect 325 36114 339 36131
rect 203 36095 339 36114
rect 203 36076 219 36095
rect 253 36076 305 36095
rect 203 36042 209 36076
rect 253 36061 291 36076
rect 243 36042 291 36061
rect 325 36042 339 36061
rect 203 36025 339 36042
rect 203 36004 219 36025
rect 253 36004 305 36025
rect 203 35970 209 36004
rect 253 35991 291 36004
rect 243 35970 291 35991
rect 325 35970 339 35991
rect 203 35932 339 35970
rect 203 35898 209 35932
rect 243 35898 291 35932
rect 325 35898 339 35932
rect 203 35891 339 35898
rect 203 35860 278 35891
rect 312 35860 339 35891
rect 203 35826 209 35860
rect 243 35857 278 35860
rect 243 35826 291 35857
rect 325 35826 339 35860
rect 203 35823 339 35826
rect 203 35789 278 35823
rect 312 35789 339 35823
rect 203 35788 339 35789
rect 203 35754 209 35788
rect 243 35755 291 35788
rect 243 35754 278 35755
rect 325 35754 339 35788
rect 203 35721 278 35754
rect 312 35721 339 35754
rect 203 35716 339 35721
rect 203 35682 209 35716
rect 243 35687 291 35716
rect 243 35682 278 35687
rect 325 35682 339 35716
rect 203 35653 278 35682
rect 312 35673 339 35682
rect 22823 37483 22827 37517
rect 22861 37483 22897 37517
rect 22931 37483 22967 37517
rect 23001 37483 23037 37517
rect 23071 37483 23107 37517
rect 23141 37483 23177 37517
rect 23211 37483 23247 37517
rect 23281 37483 23317 37517
rect 23351 37483 23387 37517
rect 23421 37483 23457 37517
rect 23491 37483 23527 37517
rect 23561 37483 23597 37517
rect 23631 37506 23711 37517
rect 23745 37506 23794 37540
rect 23828 37506 23877 37540
rect 23911 37506 23959 37540
rect 23993 37518 27021 37540
rect 23993 37506 24093 37518
rect 23631 37484 24093 37506
rect 24127 37484 24162 37518
rect 24196 37484 24231 37518
rect 24265 37484 24300 37518
rect 24334 37484 24369 37518
rect 24403 37484 24438 37518
rect 24472 37484 24507 37518
rect 24541 37484 24576 37518
rect 24610 37484 24645 37518
rect 24679 37484 24714 37518
rect 24748 37484 24783 37518
rect 24817 37484 24852 37518
rect 24886 37484 24921 37518
rect 24955 37484 24990 37518
rect 25024 37484 25059 37518
rect 25093 37484 25127 37518
rect 25161 37484 25195 37518
rect 25229 37484 25263 37518
rect 25297 37484 25331 37518
rect 25365 37484 25399 37518
rect 25433 37484 25467 37518
rect 25501 37484 25535 37518
rect 25569 37484 25603 37518
rect 25637 37484 25671 37518
rect 25705 37484 25739 37518
rect 25773 37484 25807 37518
rect 25841 37484 25875 37518
rect 25909 37484 25943 37518
rect 25977 37484 26011 37518
rect 26045 37484 26079 37518
rect 26113 37484 26147 37518
rect 26181 37484 26215 37518
rect 26249 37484 26283 37518
rect 26317 37484 26351 37518
rect 26385 37484 26419 37518
rect 26453 37484 26487 37518
rect 26521 37484 26555 37518
rect 26589 37484 26623 37518
rect 26657 37484 26691 37518
rect 26725 37484 26759 37518
rect 26793 37484 26827 37518
rect 26861 37484 26895 37518
rect 26929 37484 26963 37518
rect 26997 37484 27021 37518
rect 23631 37483 27021 37484
rect 22823 37454 27021 37483
rect 22823 37449 23711 37454
rect 22823 37415 22827 37449
rect 22861 37415 22897 37449
rect 22931 37415 22967 37449
rect 23001 37415 23037 37449
rect 23071 37415 23107 37449
rect 23141 37415 23177 37449
rect 23211 37415 23247 37449
rect 23281 37415 23317 37449
rect 23351 37415 23387 37449
rect 23421 37415 23457 37449
rect 23491 37415 23527 37449
rect 23561 37415 23597 37449
rect 23631 37420 23711 37449
rect 23745 37420 23794 37454
rect 23828 37420 23877 37454
rect 23911 37420 23959 37454
rect 23993 37440 27021 37454
rect 23993 37420 24093 37440
rect 23631 37415 24093 37420
rect 22823 37406 24093 37415
rect 24127 37406 24162 37440
rect 24196 37406 24231 37440
rect 24265 37406 24300 37440
rect 24334 37406 24369 37440
rect 24403 37406 24438 37440
rect 24472 37406 24507 37440
rect 24541 37406 24576 37440
rect 24610 37406 24645 37440
rect 24679 37406 24714 37440
rect 24748 37406 24783 37440
rect 24817 37406 24852 37440
rect 24886 37406 24921 37440
rect 24955 37406 24990 37440
rect 25024 37406 25059 37440
rect 25093 37406 25127 37440
rect 25161 37406 25195 37440
rect 25229 37406 25263 37440
rect 25297 37406 25331 37440
rect 25365 37406 25399 37440
rect 25433 37406 25467 37440
rect 25501 37406 25535 37440
rect 25569 37406 25603 37440
rect 25637 37406 25671 37440
rect 25705 37406 25739 37440
rect 25773 37406 25807 37440
rect 25841 37406 25875 37440
rect 25909 37406 25943 37440
rect 25977 37406 26011 37440
rect 26045 37406 26079 37440
rect 26113 37406 26147 37440
rect 26181 37406 26215 37440
rect 26249 37406 26283 37440
rect 26317 37406 26351 37440
rect 26385 37406 26419 37440
rect 26453 37406 26487 37440
rect 26521 37406 26555 37440
rect 26589 37406 26623 37440
rect 26657 37406 26691 37440
rect 26725 37406 26759 37440
rect 26793 37406 26827 37440
rect 26861 37406 26895 37440
rect 26929 37406 26963 37440
rect 26997 37406 27021 37440
rect 22823 37381 27021 37406
rect 22823 37347 22827 37381
rect 22861 37347 22897 37381
rect 22931 37347 22967 37381
rect 23001 37347 23037 37381
rect 23071 37347 23107 37381
rect 23141 37347 23177 37381
rect 23211 37347 23247 37381
rect 23281 37347 23317 37381
rect 23351 37347 23387 37381
rect 23421 37347 23457 37381
rect 23491 37347 23527 37381
rect 23561 37347 23597 37381
rect 23631 37368 27021 37381
rect 23631 37347 23711 37368
rect 22823 37334 23711 37347
rect 23745 37334 23794 37368
rect 23828 37334 23877 37368
rect 23911 37334 23959 37368
rect 23993 37362 27021 37368
rect 23993 37334 24093 37362
rect 22823 37328 24093 37334
rect 24127 37328 24162 37362
rect 24196 37328 24231 37362
rect 24265 37328 24300 37362
rect 24334 37328 24369 37362
rect 24403 37328 24438 37362
rect 24472 37328 24507 37362
rect 24541 37328 24576 37362
rect 24610 37328 24645 37362
rect 24679 37328 24714 37362
rect 24748 37328 24783 37362
rect 24817 37328 24852 37362
rect 24886 37328 24921 37362
rect 24955 37328 24990 37362
rect 25024 37328 25059 37362
rect 25093 37328 25127 37362
rect 25161 37328 25195 37362
rect 25229 37328 25263 37362
rect 25297 37328 25331 37362
rect 25365 37328 25399 37362
rect 25433 37328 25467 37362
rect 25501 37328 25535 37362
rect 25569 37328 25603 37362
rect 25637 37328 25671 37362
rect 25705 37328 25739 37362
rect 25773 37328 25807 37362
rect 25841 37328 25875 37362
rect 25909 37328 25943 37362
rect 25977 37328 26011 37362
rect 26045 37328 26079 37362
rect 26113 37328 26147 37362
rect 26181 37328 26215 37362
rect 26249 37328 26283 37362
rect 26317 37328 26351 37362
rect 26385 37328 26419 37362
rect 26453 37328 26487 37362
rect 26521 37328 26555 37362
rect 26589 37328 26623 37362
rect 26657 37328 26691 37362
rect 26725 37328 26759 37362
rect 26793 37328 26827 37362
rect 26861 37328 26895 37362
rect 26929 37328 26963 37362
rect 26997 37328 27021 37362
rect 22823 37313 27021 37328
rect 22823 37279 22827 37313
rect 22861 37279 22897 37313
rect 22931 37279 22967 37313
rect 23001 37279 23037 37313
rect 23071 37279 23107 37313
rect 23141 37279 23177 37313
rect 23211 37279 23247 37313
rect 23281 37279 23317 37313
rect 23351 37279 23387 37313
rect 23421 37279 23457 37313
rect 23491 37279 23527 37313
rect 23561 37279 23597 37313
rect 23631 37284 27021 37313
rect 23631 37282 24093 37284
rect 23631 37279 23711 37282
rect 22823 37248 23711 37279
rect 23745 37248 23794 37282
rect 23828 37248 23877 37282
rect 23911 37248 23959 37282
rect 23993 37250 24093 37282
rect 24127 37250 24162 37284
rect 24196 37250 24231 37284
rect 24265 37250 24300 37284
rect 24334 37250 24369 37284
rect 24403 37250 24438 37284
rect 24472 37250 24507 37284
rect 24541 37250 24576 37284
rect 24610 37250 24645 37284
rect 24679 37250 24714 37284
rect 24748 37250 24783 37284
rect 24817 37250 24852 37284
rect 24886 37250 24921 37284
rect 24955 37250 24990 37284
rect 25024 37250 25059 37284
rect 25093 37250 25127 37284
rect 25161 37250 25195 37284
rect 25229 37250 25263 37284
rect 25297 37250 25331 37284
rect 25365 37250 25399 37284
rect 25433 37250 25467 37284
rect 25501 37250 25535 37284
rect 25569 37250 25603 37284
rect 25637 37250 25671 37284
rect 25705 37250 25739 37284
rect 25773 37250 25807 37284
rect 25841 37250 25875 37284
rect 25909 37250 25943 37284
rect 25977 37250 26011 37284
rect 26045 37250 26079 37284
rect 26113 37250 26147 37284
rect 26181 37250 26215 37284
rect 26249 37250 26283 37284
rect 26317 37250 26351 37284
rect 26385 37250 26419 37284
rect 26453 37250 26487 37284
rect 26521 37250 26555 37284
rect 26589 37250 26623 37284
rect 26657 37250 26691 37284
rect 26725 37250 26759 37284
rect 26793 37250 26827 37284
rect 26861 37250 26895 37284
rect 26929 37250 26963 37284
rect 26997 37250 27021 37284
rect 23993 37248 27021 37250
rect 22823 37247 27021 37248
rect 22823 37245 23635 37247
rect 22823 37211 22827 37245
rect 22861 37211 22897 37245
rect 22931 37211 22967 37245
rect 23001 37211 23037 37245
rect 23071 37211 23107 37245
rect 23141 37211 23177 37245
rect 23211 37211 23247 37245
rect 23281 37211 23317 37245
rect 23351 37211 23387 37245
rect 23421 37211 23457 37245
rect 23491 37211 23527 37245
rect 23561 37211 23597 37245
rect 23631 37211 23635 37245
rect 22823 37177 23635 37211
rect 22823 37143 22827 37177
rect 22861 37143 22897 37177
rect 22931 37143 22967 37177
rect 23001 37143 23037 37177
rect 23071 37143 23107 37177
rect 23141 37143 23177 37177
rect 23211 37143 23247 37177
rect 23281 37143 23317 37177
rect 23351 37143 23387 37177
rect 23421 37143 23457 37177
rect 23491 37143 23527 37177
rect 23561 37143 23597 37177
rect 23631 37143 23635 37177
rect 22823 37109 23635 37143
rect 22823 37075 22827 37109
rect 22861 37075 22897 37109
rect 22931 37075 22967 37109
rect 23001 37075 23037 37109
rect 23071 37075 23107 37109
rect 23141 37075 23177 37109
rect 23211 37075 23247 37109
rect 23281 37075 23317 37109
rect 23351 37075 23387 37109
rect 23421 37075 23457 37109
rect 23491 37075 23527 37109
rect 23561 37075 23597 37109
rect 23631 37075 23635 37109
rect 22823 37041 23635 37075
rect 22823 37007 22827 37041
rect 22861 37007 22897 37041
rect 22931 37007 22967 37041
rect 23001 37007 23037 37041
rect 23071 37007 23107 37041
rect 23141 37007 23177 37041
rect 23211 37007 23247 37041
rect 23281 37007 23317 37041
rect 23351 37007 23387 37041
rect 23421 37007 23457 37041
rect 23491 37007 23527 37041
rect 23561 37007 23597 37041
rect 23631 37007 23635 37041
rect 22823 36973 23635 37007
rect 22823 36939 22827 36973
rect 22861 36939 22897 36973
rect 22931 36939 22967 36973
rect 23001 36939 23037 36973
rect 23071 36939 23107 36973
rect 23141 36939 23177 36973
rect 23211 36939 23247 36973
rect 23281 36939 23317 36973
rect 23351 36939 23387 36973
rect 23421 36939 23457 36973
rect 23491 36939 23527 36973
rect 23561 36939 23597 36973
rect 23631 36939 23635 36973
rect 22823 36905 23635 36939
rect 22823 36871 22827 36905
rect 22861 36871 22897 36905
rect 22931 36871 22967 36905
rect 23001 36871 23037 36905
rect 23071 36871 23107 36905
rect 23141 36871 23177 36905
rect 23211 36871 23247 36905
rect 23281 36871 23317 36905
rect 23351 36871 23387 36905
rect 23421 36871 23457 36905
rect 23491 36871 23527 36905
rect 23561 36871 23597 36905
rect 23631 36871 23635 36905
rect 22823 36837 23635 36871
rect 22823 36803 22827 36837
rect 22861 36803 22897 36837
rect 22931 36803 22967 36837
rect 23001 36803 23037 36837
rect 23071 36803 23107 36837
rect 23141 36803 23177 36837
rect 23211 36803 23247 36837
rect 23281 36803 23317 36837
rect 23351 36803 23387 36837
rect 23421 36803 23457 36837
rect 23491 36803 23527 36837
rect 23561 36803 23597 36837
rect 23631 36803 23635 36837
rect 22823 36769 23635 36803
rect 22823 36735 22827 36769
rect 22861 36735 22897 36769
rect 22931 36735 22967 36769
rect 23001 36735 23037 36769
rect 23071 36735 23107 36769
rect 23141 36735 23177 36769
rect 23211 36735 23247 36769
rect 23281 36735 23317 36769
rect 23351 36735 23387 36769
rect 23421 36735 23457 36769
rect 23491 36735 23527 36769
rect 23561 36735 23597 36769
rect 23631 36735 23635 36769
rect 22823 36701 23635 36735
rect 22823 36667 22827 36701
rect 22861 36667 22897 36701
rect 22931 36667 22967 36701
rect 23001 36667 23037 36701
rect 23071 36667 23107 36701
rect 23141 36667 23177 36701
rect 23211 36667 23247 36701
rect 23281 36667 23317 36701
rect 23351 36667 23387 36701
rect 23421 36667 23457 36701
rect 23491 36667 23527 36701
rect 23561 36667 23597 36701
rect 23631 36667 23635 36701
rect 22823 36633 23635 36667
rect 22823 36599 22827 36633
rect 22861 36599 22897 36633
rect 22931 36599 22967 36633
rect 23001 36599 23037 36633
rect 23071 36599 23107 36633
rect 23141 36599 23177 36633
rect 23211 36599 23247 36633
rect 23281 36599 23317 36633
rect 23351 36599 23387 36633
rect 23421 36599 23457 36633
rect 23491 36599 23527 36633
rect 23561 36599 23597 36633
rect 23631 36599 23635 36633
rect 22823 36565 23635 36599
rect 22823 36531 22827 36565
rect 22861 36531 22897 36565
rect 22931 36531 22967 36565
rect 23001 36531 23037 36565
rect 23071 36531 23107 36565
rect 23141 36531 23177 36565
rect 23211 36531 23247 36565
rect 23281 36531 23317 36565
rect 23351 36531 23387 36565
rect 23421 36531 23457 36565
rect 23491 36531 23527 36565
rect 23561 36531 23597 36565
rect 23631 36531 23635 36565
rect 22823 36497 23635 36531
rect 22823 36463 22827 36497
rect 22861 36463 22897 36497
rect 22931 36463 22967 36497
rect 23001 36463 23037 36497
rect 23071 36463 23107 36497
rect 23141 36463 23177 36497
rect 23211 36463 23247 36497
rect 23281 36463 23317 36497
rect 23351 36463 23387 36497
rect 23421 36463 23457 36497
rect 23491 36463 23527 36497
rect 23561 36463 23597 36497
rect 23631 36463 23635 36497
rect 22823 36429 23635 36463
rect 22823 36395 22827 36429
rect 22861 36395 22897 36429
rect 22931 36395 22967 36429
rect 23001 36395 23037 36429
rect 23071 36395 23107 36429
rect 23141 36395 23177 36429
rect 23211 36395 23247 36429
rect 23281 36395 23317 36429
rect 23351 36395 23387 36429
rect 23421 36395 23457 36429
rect 23491 36395 23527 36429
rect 23561 36395 23597 36429
rect 23631 36395 23635 36429
rect 22823 36384 23635 36395
rect 22823 36361 22829 36384
rect 22863 36361 22911 36384
rect 22945 36361 22993 36384
rect 23027 36361 23075 36384
rect 23109 36361 23157 36384
rect 23191 36361 23239 36384
rect 23273 36361 23635 36384
rect 22823 36327 22827 36361
rect 22863 36350 22897 36361
rect 22945 36350 22967 36361
rect 23027 36350 23037 36361
rect 22861 36327 22897 36350
rect 22931 36327 22967 36350
rect 23001 36327 23037 36350
rect 23071 36350 23075 36361
rect 23141 36350 23157 36361
rect 23211 36350 23239 36361
rect 23071 36327 23107 36350
rect 23141 36327 23177 36350
rect 23211 36327 23247 36350
rect 23281 36327 23317 36361
rect 23351 36327 23387 36361
rect 23421 36327 23457 36361
rect 23491 36327 23527 36361
rect 23561 36327 23597 36361
rect 23631 36327 23635 36361
rect 22823 36312 23635 36327
rect 22823 36293 22829 36312
rect 22863 36293 22911 36312
rect 22945 36293 22993 36312
rect 23027 36293 23075 36312
rect 23109 36293 23157 36312
rect 23191 36293 23239 36312
rect 23273 36293 23635 36312
rect 22823 36259 22827 36293
rect 22863 36278 22897 36293
rect 22945 36278 22967 36293
rect 23027 36278 23037 36293
rect 22861 36259 22897 36278
rect 22931 36259 22967 36278
rect 23001 36259 23037 36278
rect 23071 36278 23075 36293
rect 23141 36278 23157 36293
rect 23211 36278 23239 36293
rect 23071 36259 23107 36278
rect 23141 36259 23177 36278
rect 23211 36259 23247 36278
rect 23281 36259 23317 36293
rect 23351 36259 23387 36293
rect 23421 36259 23457 36293
rect 23491 36259 23527 36293
rect 23561 36259 23597 36293
rect 23631 36259 23635 36293
rect 22823 36240 23635 36259
rect 22823 36225 22829 36240
rect 22863 36225 22911 36240
rect 22945 36225 22993 36240
rect 23027 36225 23075 36240
rect 23109 36225 23157 36240
rect 23191 36225 23239 36240
rect 23273 36225 23635 36240
rect 22823 36191 22827 36225
rect 22863 36206 22897 36225
rect 22945 36206 22967 36225
rect 23027 36206 23037 36225
rect 22861 36191 22897 36206
rect 22931 36191 22967 36206
rect 23001 36191 23037 36206
rect 23071 36206 23075 36225
rect 23141 36206 23157 36225
rect 23211 36206 23239 36225
rect 23071 36191 23107 36206
rect 23141 36191 23177 36206
rect 23211 36191 23247 36206
rect 23281 36191 23317 36225
rect 23351 36191 23387 36225
rect 23421 36191 23457 36225
rect 23491 36191 23527 36225
rect 23561 36191 23597 36225
rect 23631 36191 23635 36225
rect 22823 36168 23635 36191
rect 22823 36157 22829 36168
rect 22863 36157 22911 36168
rect 22945 36157 22993 36168
rect 23027 36157 23075 36168
rect 23109 36157 23157 36168
rect 23191 36157 23239 36168
rect 23273 36157 23635 36168
rect 22823 36123 22827 36157
rect 22863 36134 22897 36157
rect 22945 36134 22967 36157
rect 23027 36134 23037 36157
rect 22861 36123 22897 36134
rect 22931 36123 22967 36134
rect 23001 36123 23037 36134
rect 23071 36134 23075 36157
rect 23141 36134 23157 36157
rect 23211 36134 23239 36157
rect 23071 36123 23107 36134
rect 23141 36123 23177 36134
rect 23211 36123 23247 36134
rect 23281 36123 23317 36157
rect 23351 36123 23387 36157
rect 23421 36123 23457 36157
rect 23491 36123 23527 36157
rect 23561 36123 23597 36157
rect 23631 36123 23635 36157
rect 22823 36096 23635 36123
rect 22823 36089 22829 36096
rect 22863 36089 22911 36096
rect 22945 36089 22993 36096
rect 23027 36089 23075 36096
rect 23109 36089 23157 36096
rect 23191 36089 23239 36096
rect 23273 36089 23635 36096
rect 22823 36055 22827 36089
rect 22863 36062 22897 36089
rect 22945 36062 22967 36089
rect 23027 36062 23037 36089
rect 22861 36055 22897 36062
rect 22931 36055 22967 36062
rect 23001 36055 23037 36062
rect 23071 36062 23075 36089
rect 23141 36062 23157 36089
rect 23211 36062 23239 36089
rect 23071 36055 23107 36062
rect 23141 36055 23177 36062
rect 23211 36055 23247 36062
rect 23281 36055 23317 36089
rect 23351 36055 23387 36089
rect 23421 36055 23457 36089
rect 23491 36055 23527 36089
rect 23561 36055 23597 36089
rect 23631 36055 23635 36089
rect 22823 36024 23635 36055
rect 22823 36021 22829 36024
rect 22863 36021 22911 36024
rect 22945 36021 22993 36024
rect 23027 36021 23075 36024
rect 23109 36021 23157 36024
rect 23191 36021 23239 36024
rect 23273 36021 23635 36024
rect 22823 35987 22827 36021
rect 22863 35990 22897 36021
rect 22945 35990 22967 36021
rect 23027 35990 23037 36021
rect 22861 35987 22897 35990
rect 22931 35987 22967 35990
rect 23001 35987 23037 35990
rect 23071 35990 23075 36021
rect 23141 35990 23157 36021
rect 23211 35990 23239 36021
rect 23071 35987 23107 35990
rect 23141 35987 23177 35990
rect 23211 35987 23247 35990
rect 23281 35987 23317 36021
rect 23351 35987 23387 36021
rect 23421 35987 23457 36021
rect 23491 35987 23527 36021
rect 23561 35987 23597 36021
rect 23631 35987 23635 36021
rect 22823 35953 23635 35987
rect 22823 35919 22827 35953
rect 22861 35952 22897 35953
rect 22931 35952 22967 35953
rect 23001 35952 23037 35953
rect 22863 35919 22897 35952
rect 22945 35919 22967 35952
rect 23027 35919 23037 35952
rect 23071 35952 23107 35953
rect 23141 35952 23177 35953
rect 23211 35952 23247 35953
rect 23071 35919 23075 35952
rect 23141 35919 23157 35952
rect 23211 35919 23239 35952
rect 23281 35919 23317 35953
rect 23351 35919 23387 35953
rect 23421 35919 23457 35953
rect 23491 35919 23527 35953
rect 23561 35919 23597 35953
rect 23631 35919 23635 35953
rect 22823 35918 22829 35919
rect 22863 35918 22911 35919
rect 22945 35918 22993 35919
rect 23027 35918 23075 35919
rect 23109 35918 23157 35919
rect 23191 35918 23239 35919
rect 23273 35918 23635 35919
rect 22823 35885 23635 35918
rect 22823 35851 22827 35885
rect 22861 35880 22897 35885
rect 22931 35880 22967 35885
rect 23001 35880 23037 35885
rect 22863 35851 22897 35880
rect 22945 35851 22967 35880
rect 23027 35851 23037 35880
rect 23071 35880 23107 35885
rect 23141 35880 23177 35885
rect 23211 35880 23247 35885
rect 23071 35851 23075 35880
rect 23141 35851 23157 35880
rect 23211 35851 23239 35880
rect 23281 35851 23317 35885
rect 23351 35851 23387 35885
rect 23421 35851 23457 35885
rect 23491 35851 23527 35885
rect 23561 35851 23597 35885
rect 23631 35851 23635 35885
rect 22823 35846 22829 35851
rect 22863 35846 22911 35851
rect 22945 35846 22993 35851
rect 23027 35846 23075 35851
rect 23109 35846 23157 35851
rect 23191 35846 23239 35851
rect 23273 35846 23635 35851
rect 22823 35817 23635 35846
rect 22823 35783 22827 35817
rect 22861 35808 22897 35817
rect 22931 35808 22967 35817
rect 23001 35808 23037 35817
rect 22863 35783 22897 35808
rect 22945 35783 22967 35808
rect 23027 35783 23037 35808
rect 23071 35808 23107 35817
rect 23141 35808 23177 35817
rect 23211 35808 23247 35817
rect 23071 35783 23075 35808
rect 23141 35783 23157 35808
rect 23211 35783 23239 35808
rect 23281 35783 23317 35817
rect 23351 35783 23387 35817
rect 23421 35783 23457 35817
rect 23491 35783 23527 35817
rect 23561 35783 23597 35817
rect 23631 35783 23635 35817
rect 22823 35774 22829 35783
rect 22863 35774 22911 35783
rect 22945 35774 22993 35783
rect 23027 35774 23075 35783
rect 23109 35774 23157 35783
rect 23191 35774 23239 35783
rect 23273 35774 23635 35783
rect 22823 35749 23635 35774
rect 22823 35715 22827 35749
rect 22861 35736 22897 35749
rect 22931 35736 22967 35749
rect 23001 35736 23037 35749
rect 22863 35715 22897 35736
rect 22945 35715 22967 35736
rect 23027 35715 23037 35736
rect 23071 35736 23107 35749
rect 23141 35736 23177 35749
rect 23211 35736 23247 35749
rect 23071 35715 23075 35736
rect 23141 35715 23157 35736
rect 23211 35715 23239 35736
rect 23281 35715 23317 35749
rect 23351 35715 23387 35749
rect 23421 35715 23457 35749
rect 23491 35715 23527 35749
rect 23561 35715 23597 35749
rect 23631 35715 23635 35749
rect 22823 35702 22829 35715
rect 22863 35702 22911 35715
rect 22945 35702 22993 35715
rect 23027 35702 23075 35715
rect 23109 35702 23157 35715
rect 23191 35702 23239 35715
rect 23273 35702 23635 35715
rect 22823 35681 23635 35702
rect 312 35653 331 35673
rect 203 35644 331 35653
rect 203 35610 209 35644
rect 243 35619 291 35644
rect 243 35610 278 35619
rect 325 35610 331 35644
rect 203 35585 278 35610
rect 312 35585 331 35610
rect 203 35572 331 35585
rect 203 35538 209 35572
rect 243 35551 291 35572
rect 243 35538 278 35551
rect 325 35538 331 35572
rect 203 35517 278 35538
rect 312 35517 331 35538
rect 203 35500 331 35517
rect 203 35466 209 35500
rect 243 35483 291 35500
rect 243 35466 278 35483
rect 325 35466 331 35500
rect 203 35449 278 35466
rect 312 35449 331 35466
rect 203 35427 331 35449
rect 203 35393 209 35427
rect 243 35415 291 35427
rect 243 35393 278 35415
rect 325 35393 331 35427
rect 203 35381 278 35393
rect 312 35381 331 35393
rect 203 35354 331 35381
rect 203 35320 209 35354
rect 243 35347 291 35354
rect 243 35320 278 35347
rect 325 35320 331 35354
rect 203 35313 278 35320
rect 312 35313 331 35320
rect 203 35281 331 35313
rect 203 35247 209 35281
rect 243 35279 291 35281
rect 243 35247 278 35279
rect 325 35247 331 35281
rect 203 35245 278 35247
rect 312 35245 331 35247
rect 203 35211 331 35245
rect 203 35208 278 35211
rect 312 35208 331 35211
rect 203 35174 209 35208
rect 243 35177 278 35208
rect 243 35174 291 35177
rect 325 35174 331 35208
rect 203 35143 331 35174
rect 203 35135 278 35143
rect 312 35135 331 35143
rect 203 35101 209 35135
rect 243 35109 278 35135
rect 243 35101 291 35109
rect 325 35101 331 35135
rect 203 35075 331 35101
rect 203 35062 278 35075
rect 312 35062 331 35075
rect 203 35028 209 35062
rect 243 35041 278 35062
rect 243 35028 291 35041
rect 325 35028 331 35062
rect 203 35006 331 35028
rect 203 34989 278 35006
rect 312 34989 331 35006
rect 203 34955 209 34989
rect 243 34972 278 34989
rect 243 34955 291 34972
rect 325 34955 331 34989
rect 203 34937 331 34955
rect 203 34916 278 34937
rect 312 34916 331 34937
rect 203 34882 209 34916
rect 243 34903 278 34916
rect 243 34882 291 34903
rect 325 34882 331 34916
rect 203 34868 331 34882
rect 203 34843 278 34868
rect 312 34843 331 34868
rect 203 34809 209 34843
rect 243 34834 278 34843
rect 243 34809 291 34834
rect 325 34809 331 34843
rect 203 34799 331 34809
rect 203 34770 278 34799
rect 312 34770 331 34799
rect 203 34736 209 34770
rect 243 34765 278 34770
rect 243 34736 291 34765
rect 325 34736 331 34770
rect 203 34730 331 34736
rect 203 34697 278 34730
rect 312 34697 331 34730
rect 203 34663 209 34697
rect 243 34696 278 34697
rect 243 34663 291 34696
rect 325 34663 331 34697
rect 203 34661 331 34663
rect 203 34627 278 34661
rect 312 34627 331 34661
rect 203 34624 331 34627
rect 203 34590 209 34624
rect 243 34592 291 34624
rect 243 34590 278 34592
rect 325 34590 331 34624
rect 203 34558 278 34590
rect 312 34558 331 34590
rect 203 34551 331 34558
rect 203 34517 209 34551
rect 243 34523 291 34551
rect 243 34517 278 34523
rect 325 34517 331 34551
rect 203 34489 278 34517
rect 312 34489 331 34517
rect 203 34478 331 34489
rect 203 34444 209 34478
rect 243 34454 291 34478
rect 243 34444 278 34454
rect 325 34444 331 34478
rect 203 34420 278 34444
rect 312 34420 331 34444
rect 203 34405 331 34420
rect 203 34371 209 34405
rect 243 34385 291 34405
rect 243 34371 278 34385
rect 325 34371 331 34405
rect 203 34351 278 34371
rect 312 34351 331 34371
rect 203 34332 331 34351
rect 203 34298 209 34332
rect 243 34316 291 34332
rect 243 34298 278 34316
rect 325 34298 331 34332
rect 203 34282 278 34298
rect 312 34282 331 34298
rect 203 34259 331 34282
rect 203 34225 209 34259
rect 243 34247 291 34259
rect 243 34225 278 34247
rect 325 34225 331 34259
rect 203 34213 278 34225
rect 312 34213 331 34225
rect 203 34186 331 34213
rect 203 34152 209 34186
rect 243 34178 291 34186
rect 243 34152 278 34178
rect 325 34152 331 34186
rect 203 34144 278 34152
rect 312 34144 331 34152
rect 203 34113 331 34144
rect 203 34079 209 34113
rect 243 34109 291 34113
rect 243 34079 278 34109
rect 325 34079 331 34113
rect 203 34075 278 34079
rect 312 34075 331 34079
rect 203 34040 331 34075
rect 203 34006 209 34040
rect 243 34006 278 34040
rect 325 34006 331 34040
rect 203 33971 331 34006
rect 203 33967 278 33971
rect 312 33967 331 33971
rect 203 33933 209 33967
rect 243 33937 278 33967
rect 243 33933 291 33937
rect 325 33933 331 33967
rect 203 33902 331 33933
rect 203 33894 278 33902
rect 312 33894 331 33902
rect 203 33860 209 33894
rect 243 33868 278 33894
rect 243 33860 291 33868
rect 325 33860 331 33894
rect 203 33833 331 33860
rect 203 33821 278 33833
rect 312 33821 331 33833
rect 203 33787 209 33821
rect 243 33799 278 33821
rect 243 33787 291 33799
rect 325 33787 331 33821
rect 203 33764 331 33787
rect 203 33748 278 33764
rect 312 33748 331 33764
rect 203 33714 209 33748
rect 243 33730 278 33748
rect 243 33714 291 33730
rect 325 33714 331 33748
rect 203 33695 331 33714
rect 203 33675 278 33695
rect 312 33675 331 33695
rect 203 33641 209 33675
rect 243 33661 278 33675
rect 243 33641 291 33661
rect 325 33641 331 33675
rect 203 33626 331 33641
rect 203 33602 278 33626
rect 312 33602 331 33626
rect 203 33568 209 33602
rect 243 33592 278 33602
rect 243 33568 291 33592
rect 325 33568 331 33602
rect 203 33557 331 33568
rect 203 33529 278 33557
rect 312 33529 331 33557
rect 203 33495 209 33529
rect 243 33523 278 33529
rect 243 33495 291 33523
rect 325 33495 331 33529
rect 203 33488 331 33495
rect 203 33456 278 33488
rect 312 33456 331 33488
rect 203 33422 209 33456
rect 243 33454 278 33456
rect 243 33422 291 33454
rect 325 33422 331 33456
rect 203 33419 331 33422
rect 203 33385 278 33419
rect 312 33385 331 33419
rect 203 33383 331 33385
rect 203 33349 209 33383
rect 243 33350 291 33383
rect 243 33349 278 33350
rect 325 33349 331 33383
rect 203 33316 278 33349
rect 312 33316 331 33349
rect 22823 35647 22827 35681
rect 22861 35664 22897 35681
rect 22931 35664 22967 35681
rect 23001 35664 23037 35681
rect 22863 35647 22897 35664
rect 22945 35647 22967 35664
rect 23027 35647 23037 35664
rect 23071 35664 23107 35681
rect 23141 35664 23177 35681
rect 23211 35664 23247 35681
rect 23071 35647 23075 35664
rect 23141 35647 23157 35664
rect 23211 35647 23239 35664
rect 23281 35647 23317 35681
rect 23351 35647 23387 35681
rect 23421 35647 23457 35681
rect 23491 35647 23527 35681
rect 23561 35647 23597 35681
rect 23631 35647 23635 35681
rect 22823 35630 22829 35647
rect 22863 35630 22911 35647
rect 22945 35630 22993 35647
rect 23027 35630 23075 35647
rect 23109 35630 23157 35647
rect 23191 35630 23239 35647
rect 23273 35630 23635 35647
rect 22823 35613 23635 35630
rect 22823 35579 22827 35613
rect 22861 35592 22897 35613
rect 22931 35592 22967 35613
rect 23001 35592 23037 35613
rect 22863 35579 22897 35592
rect 22945 35579 22967 35592
rect 23027 35579 23037 35592
rect 23071 35592 23107 35613
rect 23141 35592 23177 35613
rect 23211 35592 23247 35613
rect 23071 35579 23075 35592
rect 23141 35579 23157 35592
rect 23211 35579 23239 35592
rect 23281 35579 23317 35613
rect 23351 35579 23387 35613
rect 23421 35579 23457 35613
rect 23491 35579 23527 35613
rect 23561 35579 23597 35613
rect 23631 35579 23635 35613
rect 22823 35558 22829 35579
rect 22863 35558 22911 35579
rect 22945 35558 22993 35579
rect 23027 35558 23075 35579
rect 23109 35558 23157 35579
rect 23191 35558 23239 35579
rect 23273 35558 23635 35579
rect 22823 35545 23635 35558
rect 22823 35511 22827 35545
rect 22861 35520 22897 35545
rect 22931 35520 22967 35545
rect 23001 35520 23037 35545
rect 22863 35511 22897 35520
rect 22945 35511 22967 35520
rect 23027 35511 23037 35520
rect 23071 35520 23107 35545
rect 23141 35520 23177 35545
rect 23211 35520 23247 35545
rect 23071 35511 23075 35520
rect 23141 35511 23157 35520
rect 23211 35511 23239 35520
rect 23281 35511 23317 35545
rect 23351 35511 23387 35545
rect 23421 35511 23457 35545
rect 23491 35511 23527 35545
rect 23561 35511 23597 35545
rect 23631 35511 23635 35545
rect 22823 35486 22829 35511
rect 22863 35486 22911 35511
rect 22945 35486 22993 35511
rect 23027 35486 23075 35511
rect 23109 35486 23157 35511
rect 23191 35486 23239 35511
rect 23273 35486 23635 35511
rect 22823 35477 23635 35486
rect 22823 35443 22827 35477
rect 22861 35448 22897 35477
rect 22931 35448 22967 35477
rect 23001 35448 23037 35477
rect 22863 35443 22897 35448
rect 22945 35443 22967 35448
rect 23027 35443 23037 35448
rect 23071 35448 23107 35477
rect 23141 35448 23177 35477
rect 23211 35448 23247 35477
rect 23071 35443 23075 35448
rect 23141 35443 23157 35448
rect 23211 35443 23239 35448
rect 23281 35443 23317 35477
rect 23351 35443 23387 35477
rect 23421 35443 23457 35477
rect 23491 35443 23527 35477
rect 23561 35443 23597 35477
rect 23631 35443 23635 35477
rect 22823 35414 22829 35443
rect 22863 35414 22911 35443
rect 22945 35414 22993 35443
rect 23027 35414 23075 35443
rect 23109 35414 23157 35443
rect 23191 35414 23239 35443
rect 23273 35414 23635 35443
rect 22823 35409 23635 35414
rect 22823 35375 22827 35409
rect 22861 35376 22897 35409
rect 22931 35376 22967 35409
rect 23001 35376 23037 35409
rect 22863 35375 22897 35376
rect 22945 35375 22967 35376
rect 23027 35375 23037 35376
rect 23071 35376 23107 35409
rect 23141 35376 23177 35409
rect 23211 35376 23247 35409
rect 23071 35375 23075 35376
rect 23141 35375 23157 35376
rect 23211 35375 23239 35376
rect 23281 35375 23317 35409
rect 23351 35375 23387 35409
rect 23421 35375 23457 35409
rect 23491 35375 23527 35409
rect 23561 35375 23597 35409
rect 23631 35375 23635 35409
rect 22823 35342 22829 35375
rect 22863 35342 22911 35375
rect 22945 35342 22993 35375
rect 23027 35342 23075 35375
rect 23109 35342 23157 35375
rect 23191 35342 23239 35375
rect 23273 35342 23635 35375
rect 22823 35341 23635 35342
rect 22823 35307 22827 35341
rect 22861 35307 22897 35341
rect 22931 35307 22967 35341
rect 23001 35307 23037 35341
rect 23071 35307 23107 35341
rect 23141 35307 23177 35341
rect 23211 35307 23247 35341
rect 23281 35307 23317 35341
rect 23351 35307 23387 35341
rect 23421 35307 23457 35341
rect 23491 35307 23527 35341
rect 23561 35307 23597 35341
rect 23631 35307 23635 35341
rect 22823 35304 23635 35307
rect 22823 35273 22829 35304
rect 22863 35273 22911 35304
rect 22945 35273 22993 35304
rect 23027 35273 23075 35304
rect 23109 35273 23157 35304
rect 23191 35273 23239 35304
rect 23273 35273 23635 35304
rect 22823 35239 22827 35273
rect 22863 35270 22897 35273
rect 22945 35270 22967 35273
rect 23027 35270 23037 35273
rect 22861 35239 22897 35270
rect 22931 35239 22967 35270
rect 23001 35239 23037 35270
rect 23071 35270 23075 35273
rect 23141 35270 23157 35273
rect 23211 35270 23239 35273
rect 23071 35239 23107 35270
rect 23141 35239 23177 35270
rect 23211 35239 23247 35270
rect 23281 35239 23317 35273
rect 23351 35239 23387 35273
rect 23421 35239 23457 35273
rect 23491 35239 23527 35273
rect 23561 35239 23597 35273
rect 23631 35239 23635 35273
rect 22823 35232 23635 35239
rect 22823 35205 22829 35232
rect 22863 35205 22911 35232
rect 22945 35205 22993 35232
rect 23027 35205 23075 35232
rect 23109 35205 23157 35232
rect 23191 35205 23239 35232
rect 23273 35205 23635 35232
rect 22823 35171 22827 35205
rect 22863 35198 22897 35205
rect 22945 35198 22967 35205
rect 23027 35198 23037 35205
rect 22861 35171 22897 35198
rect 22931 35171 22967 35198
rect 23001 35171 23037 35198
rect 23071 35198 23075 35205
rect 23141 35198 23157 35205
rect 23211 35198 23239 35205
rect 23071 35171 23107 35198
rect 23141 35171 23177 35198
rect 23211 35171 23247 35198
rect 23281 35171 23317 35205
rect 23351 35171 23387 35205
rect 23421 35171 23457 35205
rect 23491 35171 23527 35205
rect 23561 35171 23597 35205
rect 23631 35171 23635 35205
rect 22823 35160 23635 35171
rect 22823 35137 22829 35160
rect 22863 35137 22911 35160
rect 22945 35137 22993 35160
rect 23027 35137 23075 35160
rect 23109 35137 23157 35160
rect 23191 35137 23239 35160
rect 23273 35137 23635 35160
rect 22823 35103 22827 35137
rect 22863 35126 22897 35137
rect 22945 35126 22967 35137
rect 23027 35126 23037 35137
rect 22861 35103 22897 35126
rect 22931 35103 22967 35126
rect 23001 35103 23037 35126
rect 23071 35126 23075 35137
rect 23141 35126 23157 35137
rect 23211 35126 23239 35137
rect 23071 35103 23107 35126
rect 23141 35103 23177 35126
rect 23211 35103 23247 35126
rect 23281 35103 23317 35137
rect 23351 35103 23387 35137
rect 23421 35103 23457 35137
rect 23491 35103 23527 35137
rect 23561 35103 23597 35137
rect 23631 35103 23635 35137
rect 22823 35088 23635 35103
rect 22823 35069 22829 35088
rect 22863 35069 22911 35088
rect 22945 35069 22993 35088
rect 23027 35069 23075 35088
rect 23109 35069 23157 35088
rect 23191 35069 23239 35088
rect 23273 35069 23635 35088
rect 22823 35035 22827 35069
rect 22863 35054 22897 35069
rect 22945 35054 22967 35069
rect 23027 35054 23037 35069
rect 22861 35035 22897 35054
rect 22931 35035 22967 35054
rect 23001 35035 23037 35054
rect 23071 35054 23075 35069
rect 23141 35054 23157 35069
rect 23211 35054 23239 35069
rect 23071 35035 23107 35054
rect 23141 35035 23177 35054
rect 23211 35035 23247 35054
rect 23281 35035 23317 35069
rect 23351 35035 23387 35069
rect 23421 35035 23457 35069
rect 23491 35035 23527 35069
rect 23561 35035 23597 35069
rect 23631 35035 23635 35069
rect 22823 35016 23635 35035
rect 22823 35001 22829 35016
rect 22863 35001 22911 35016
rect 22945 35001 22993 35016
rect 23027 35001 23075 35016
rect 23109 35001 23157 35016
rect 23191 35001 23239 35016
rect 23273 35001 23635 35016
rect 22823 34967 22827 35001
rect 22863 34982 22897 35001
rect 22945 34982 22967 35001
rect 23027 34982 23037 35001
rect 22861 34967 22897 34982
rect 22931 34967 22967 34982
rect 23001 34967 23037 34982
rect 23071 34982 23075 35001
rect 23141 34982 23157 35001
rect 23211 34982 23239 35001
rect 23071 34967 23107 34982
rect 23141 34967 23177 34982
rect 23211 34967 23247 34982
rect 23281 34967 23317 35001
rect 23351 34967 23387 35001
rect 23421 34967 23457 35001
rect 23491 34967 23527 35001
rect 23561 34967 23597 35001
rect 23631 34967 23635 35001
rect 22823 34944 23635 34967
rect 22823 34933 22829 34944
rect 22863 34933 22911 34944
rect 22945 34933 22993 34944
rect 23027 34933 23075 34944
rect 23109 34933 23157 34944
rect 23191 34933 23239 34944
rect 23273 34933 23635 34944
rect 22823 34899 22827 34933
rect 22863 34910 22897 34933
rect 22945 34910 22967 34933
rect 23027 34910 23037 34933
rect 22861 34899 22897 34910
rect 22931 34899 22967 34910
rect 23001 34899 23037 34910
rect 23071 34910 23075 34933
rect 23141 34910 23157 34933
rect 23211 34910 23239 34933
rect 23071 34899 23107 34910
rect 23141 34899 23177 34910
rect 23211 34899 23247 34910
rect 23281 34899 23317 34933
rect 23351 34899 23387 34933
rect 23421 34899 23457 34933
rect 23491 34899 23527 34933
rect 23561 34899 23597 34933
rect 23631 34899 23635 34933
rect 22823 34872 23635 34899
rect 22823 34865 22829 34872
rect 22863 34865 22911 34872
rect 22945 34865 22993 34872
rect 23027 34865 23075 34872
rect 23109 34865 23157 34872
rect 23191 34865 23239 34872
rect 23273 34865 23635 34872
rect 22823 34831 22827 34865
rect 22863 34838 22897 34865
rect 22945 34838 22967 34865
rect 23027 34838 23037 34865
rect 22861 34831 22897 34838
rect 22931 34831 22967 34838
rect 23001 34831 23037 34838
rect 23071 34838 23075 34865
rect 23141 34838 23157 34865
rect 23211 34838 23239 34865
rect 23071 34831 23107 34838
rect 23141 34831 23177 34838
rect 23211 34831 23247 34838
rect 23281 34831 23317 34865
rect 23351 34831 23387 34865
rect 23421 34831 23457 34865
rect 23491 34831 23527 34865
rect 23561 34831 23597 34865
rect 23631 34831 23635 34865
rect 22823 34800 23635 34831
rect 22823 34797 22829 34800
rect 22863 34797 22911 34800
rect 22945 34797 22993 34800
rect 23027 34797 23075 34800
rect 23109 34797 23157 34800
rect 23191 34797 23239 34800
rect 23273 34797 23635 34800
rect 22823 34763 22827 34797
rect 22863 34766 22897 34797
rect 22945 34766 22967 34797
rect 23027 34766 23037 34797
rect 22861 34763 22897 34766
rect 22931 34763 22967 34766
rect 23001 34763 23037 34766
rect 23071 34766 23075 34797
rect 23141 34766 23157 34797
rect 23211 34766 23239 34797
rect 23071 34763 23107 34766
rect 23141 34763 23177 34766
rect 23211 34763 23247 34766
rect 23281 34763 23317 34797
rect 23351 34763 23387 34797
rect 23421 34763 23457 34797
rect 23491 34763 23527 34797
rect 23561 34763 23597 34797
rect 23631 34763 23635 34797
rect 22823 34729 23635 34763
rect 22823 34695 22827 34729
rect 22861 34728 22897 34729
rect 22931 34728 22967 34729
rect 23001 34728 23037 34729
rect 22863 34695 22897 34728
rect 22945 34695 22967 34728
rect 23027 34695 23037 34728
rect 23071 34728 23107 34729
rect 23141 34728 23177 34729
rect 23211 34728 23247 34729
rect 23071 34695 23075 34728
rect 23141 34695 23157 34728
rect 23211 34695 23239 34728
rect 23281 34695 23317 34729
rect 23351 34695 23387 34729
rect 23421 34695 23457 34729
rect 23491 34695 23527 34729
rect 23561 34695 23597 34729
rect 23631 34695 23635 34729
rect 22823 34694 22829 34695
rect 22863 34694 22911 34695
rect 22945 34694 22993 34695
rect 23027 34694 23075 34695
rect 23109 34694 23157 34695
rect 23191 34694 23239 34695
rect 23273 34694 23635 34695
rect 22823 34661 23635 34694
rect 22823 34627 22827 34661
rect 22861 34656 22897 34661
rect 22931 34656 22967 34661
rect 23001 34656 23037 34661
rect 22863 34627 22897 34656
rect 22945 34627 22967 34656
rect 23027 34627 23037 34656
rect 23071 34656 23107 34661
rect 23141 34656 23177 34661
rect 23211 34656 23247 34661
rect 23071 34627 23075 34656
rect 23141 34627 23157 34656
rect 23211 34627 23239 34656
rect 23281 34627 23317 34661
rect 23351 34627 23387 34661
rect 23421 34627 23457 34661
rect 23491 34627 23527 34661
rect 23561 34627 23597 34661
rect 23631 34627 23635 34661
rect 22823 34622 22829 34627
rect 22863 34622 22911 34627
rect 22945 34622 22993 34627
rect 23027 34622 23075 34627
rect 23109 34622 23157 34627
rect 23191 34622 23239 34627
rect 23273 34622 23635 34627
rect 22823 34593 23635 34622
rect 22823 34559 22827 34593
rect 22861 34584 22897 34593
rect 22931 34584 22967 34593
rect 23001 34584 23037 34593
rect 22863 34559 22897 34584
rect 22945 34559 22967 34584
rect 23027 34559 23037 34584
rect 23071 34584 23107 34593
rect 23141 34584 23177 34593
rect 23211 34584 23247 34593
rect 23071 34559 23075 34584
rect 23141 34559 23157 34584
rect 23211 34559 23239 34584
rect 23281 34559 23317 34593
rect 23351 34559 23387 34593
rect 23421 34559 23457 34593
rect 23491 34559 23527 34593
rect 23561 34559 23597 34593
rect 23631 34559 23635 34593
rect 22823 34550 22829 34559
rect 22863 34550 22911 34559
rect 22945 34550 22993 34559
rect 23027 34550 23075 34559
rect 23109 34550 23157 34559
rect 23191 34550 23239 34559
rect 23273 34550 23635 34559
rect 22823 34525 23635 34550
rect 22823 34491 22827 34525
rect 22861 34512 22897 34525
rect 22931 34512 22967 34525
rect 23001 34512 23037 34525
rect 22863 34491 22897 34512
rect 22945 34491 22967 34512
rect 23027 34491 23037 34512
rect 23071 34512 23107 34525
rect 23141 34512 23177 34525
rect 23211 34512 23247 34525
rect 23071 34491 23075 34512
rect 23141 34491 23157 34512
rect 23211 34491 23239 34512
rect 23281 34491 23317 34525
rect 23351 34491 23387 34525
rect 23421 34491 23457 34525
rect 23491 34491 23527 34525
rect 23561 34491 23597 34525
rect 23631 34491 23635 34525
rect 22823 34478 22829 34491
rect 22863 34478 22911 34491
rect 22945 34478 22993 34491
rect 23027 34478 23075 34491
rect 23109 34478 23157 34491
rect 23191 34478 23239 34491
rect 23273 34478 23635 34491
rect 22823 34457 23635 34478
rect 22823 34423 22827 34457
rect 22861 34440 22897 34457
rect 22931 34440 22967 34457
rect 23001 34440 23037 34457
rect 22863 34423 22897 34440
rect 22945 34423 22967 34440
rect 23027 34423 23037 34440
rect 23071 34440 23107 34457
rect 23141 34440 23177 34457
rect 23211 34440 23247 34457
rect 23071 34423 23075 34440
rect 23141 34423 23157 34440
rect 23211 34423 23239 34440
rect 23281 34423 23317 34457
rect 23351 34423 23387 34457
rect 23421 34423 23457 34457
rect 23491 34423 23527 34457
rect 23561 34423 23597 34457
rect 23631 34423 23635 34457
rect 22823 34406 22829 34423
rect 22863 34406 22911 34423
rect 22945 34406 22993 34423
rect 23027 34406 23075 34423
rect 23109 34406 23157 34423
rect 23191 34406 23239 34423
rect 23273 34406 23635 34423
rect 22823 34389 23635 34406
rect 22823 34355 22827 34389
rect 22861 34368 22897 34389
rect 22931 34368 22967 34389
rect 23001 34368 23037 34389
rect 22863 34355 22897 34368
rect 22945 34355 22967 34368
rect 23027 34355 23037 34368
rect 23071 34368 23107 34389
rect 23141 34368 23177 34389
rect 23211 34368 23247 34389
rect 23071 34355 23075 34368
rect 23141 34355 23157 34368
rect 23211 34355 23239 34368
rect 23281 34355 23317 34389
rect 23351 34355 23387 34389
rect 23421 34355 23457 34389
rect 23491 34355 23527 34389
rect 23561 34355 23597 34389
rect 23631 34355 23635 34389
rect 22823 34334 22829 34355
rect 22863 34334 22911 34355
rect 22945 34334 22993 34355
rect 23027 34334 23075 34355
rect 23109 34334 23157 34355
rect 23191 34334 23239 34355
rect 23273 34334 23635 34355
rect 22823 34321 23635 34334
rect 22823 34287 22827 34321
rect 22861 34295 22897 34321
rect 22931 34295 22967 34321
rect 23001 34295 23037 34321
rect 22863 34287 22897 34295
rect 22945 34287 22967 34295
rect 23027 34287 23037 34295
rect 23071 34295 23107 34321
rect 23141 34295 23177 34321
rect 23211 34295 23247 34321
rect 23071 34287 23075 34295
rect 23141 34287 23157 34295
rect 23211 34287 23239 34295
rect 23281 34287 23317 34321
rect 23351 34287 23387 34321
rect 23421 34287 23457 34321
rect 23491 34287 23527 34321
rect 23561 34287 23597 34321
rect 23631 34287 23635 34321
rect 22823 34261 22829 34287
rect 22863 34261 22911 34287
rect 22945 34261 22993 34287
rect 23027 34261 23075 34287
rect 23109 34261 23157 34287
rect 23191 34261 23239 34287
rect 23273 34261 23635 34287
rect 22823 34253 23635 34261
rect 22823 34219 22827 34253
rect 22861 34222 22897 34253
rect 22931 34222 22967 34253
rect 23001 34222 23037 34253
rect 22863 34219 22897 34222
rect 22945 34219 22967 34222
rect 23027 34219 23037 34222
rect 23071 34222 23107 34253
rect 23141 34222 23177 34253
rect 23211 34222 23247 34253
rect 23071 34219 23075 34222
rect 23141 34219 23157 34222
rect 23211 34219 23239 34222
rect 23281 34219 23317 34253
rect 23351 34219 23387 34253
rect 23421 34219 23457 34253
rect 23491 34219 23527 34253
rect 23561 34219 23597 34253
rect 23631 34219 23635 34253
rect 22823 34188 22829 34219
rect 22863 34188 22911 34219
rect 22945 34188 22993 34219
rect 23027 34188 23075 34219
rect 23109 34188 23157 34219
rect 23191 34188 23239 34219
rect 23273 34188 23635 34219
rect 22823 34185 23635 34188
rect 22823 34151 22827 34185
rect 22861 34151 22897 34185
rect 22931 34151 22967 34185
rect 23001 34151 23037 34185
rect 23071 34151 23107 34185
rect 23141 34151 23177 34185
rect 23211 34151 23247 34185
rect 23281 34151 23317 34185
rect 23351 34151 23387 34185
rect 23421 34151 23457 34185
rect 23491 34151 23527 34185
rect 23561 34151 23597 34185
rect 23631 34151 23635 34185
rect 22823 34149 23635 34151
rect 22823 34117 22829 34149
rect 22863 34117 22911 34149
rect 22945 34117 22993 34149
rect 23027 34117 23075 34149
rect 23109 34117 23157 34149
rect 23191 34117 23239 34149
rect 23273 34117 23635 34149
rect 22823 34083 22827 34117
rect 22863 34115 22897 34117
rect 22945 34115 22967 34117
rect 23027 34115 23037 34117
rect 22861 34083 22897 34115
rect 22931 34083 22967 34115
rect 23001 34083 23037 34115
rect 23071 34115 23075 34117
rect 23141 34115 23157 34117
rect 23211 34115 23239 34117
rect 23071 34083 23107 34115
rect 23141 34083 23177 34115
rect 23211 34083 23247 34115
rect 23281 34083 23317 34117
rect 23351 34083 23387 34117
rect 23421 34083 23457 34117
rect 23491 34083 23527 34117
rect 23561 34083 23597 34117
rect 23631 34083 23635 34117
rect 22823 34076 23635 34083
rect 22823 34049 22829 34076
rect 22863 34049 22911 34076
rect 22945 34049 22993 34076
rect 23027 34049 23075 34076
rect 23109 34049 23157 34076
rect 23191 34049 23239 34076
rect 23273 34049 23635 34076
rect 22823 34015 22827 34049
rect 22863 34042 22897 34049
rect 22945 34042 22967 34049
rect 23027 34042 23037 34049
rect 22861 34015 22897 34042
rect 22931 34015 22967 34042
rect 23001 34015 23037 34042
rect 23071 34042 23075 34049
rect 23141 34042 23157 34049
rect 23211 34042 23239 34049
rect 23071 34015 23107 34042
rect 23141 34015 23177 34042
rect 23211 34015 23247 34042
rect 23281 34015 23317 34049
rect 23351 34015 23387 34049
rect 23421 34015 23457 34049
rect 23491 34015 23527 34049
rect 23561 34015 23597 34049
rect 23631 34015 23635 34049
rect 22823 34003 23635 34015
rect 22823 33981 22829 34003
rect 22863 33981 22911 34003
rect 22945 33981 22993 34003
rect 23027 33981 23075 34003
rect 23109 33981 23157 34003
rect 23191 33981 23239 34003
rect 23273 33981 23635 34003
rect 22823 33947 22827 33981
rect 22863 33969 22897 33981
rect 22945 33969 22967 33981
rect 23027 33969 23037 33981
rect 22861 33947 22897 33969
rect 22931 33947 22967 33969
rect 23001 33947 23037 33969
rect 23071 33969 23075 33981
rect 23141 33969 23157 33981
rect 23211 33969 23239 33981
rect 23071 33947 23107 33969
rect 23141 33947 23177 33969
rect 23211 33947 23247 33969
rect 23281 33947 23317 33981
rect 23351 33947 23387 33981
rect 23421 33947 23457 33981
rect 23491 33947 23527 33981
rect 23561 33947 23597 33981
rect 23631 33947 23635 33981
rect 22823 33930 23635 33947
rect 22823 33913 22829 33930
rect 22863 33913 22911 33930
rect 22945 33913 22993 33930
rect 23027 33913 23075 33930
rect 23109 33913 23157 33930
rect 23191 33913 23239 33930
rect 23273 33913 23635 33930
rect 22823 33879 22827 33913
rect 22863 33896 22897 33913
rect 22945 33896 22967 33913
rect 23027 33896 23037 33913
rect 22861 33879 22897 33896
rect 22931 33879 22967 33896
rect 23001 33879 23037 33896
rect 23071 33896 23075 33913
rect 23141 33896 23157 33913
rect 23211 33896 23239 33913
rect 23071 33879 23107 33896
rect 23141 33879 23177 33896
rect 23211 33879 23247 33896
rect 23281 33879 23317 33913
rect 23351 33879 23387 33913
rect 23421 33879 23457 33913
rect 23491 33879 23527 33913
rect 23561 33879 23597 33913
rect 23631 33879 23635 33913
rect 22823 33857 23635 33879
rect 22823 33845 22829 33857
rect 22863 33845 22911 33857
rect 22945 33845 22993 33857
rect 23027 33845 23075 33857
rect 23109 33845 23157 33857
rect 23191 33845 23239 33857
rect 23273 33845 23635 33857
rect 22823 33811 22827 33845
rect 22863 33823 22897 33845
rect 22945 33823 22967 33845
rect 23027 33823 23037 33845
rect 22861 33811 22897 33823
rect 22931 33811 22967 33823
rect 23001 33811 23037 33823
rect 23071 33823 23075 33845
rect 23141 33823 23157 33845
rect 23211 33823 23239 33845
rect 23071 33811 23107 33823
rect 23141 33811 23177 33823
rect 23211 33811 23247 33823
rect 23281 33811 23317 33845
rect 23351 33811 23387 33845
rect 23421 33811 23457 33845
rect 23491 33811 23527 33845
rect 23561 33811 23597 33845
rect 23631 33811 23635 33845
rect 22823 33784 23635 33811
rect 22823 33777 22829 33784
rect 22863 33777 22911 33784
rect 22945 33777 22993 33784
rect 23027 33777 23075 33784
rect 23109 33777 23157 33784
rect 23191 33777 23239 33784
rect 23273 33777 23635 33784
rect 22823 33743 22827 33777
rect 22863 33750 22897 33777
rect 22945 33750 22967 33777
rect 23027 33750 23037 33777
rect 22861 33743 22897 33750
rect 22931 33743 22967 33750
rect 23001 33743 23037 33750
rect 23071 33750 23075 33777
rect 23141 33750 23157 33777
rect 23211 33750 23239 33777
rect 23071 33743 23107 33750
rect 23141 33743 23177 33750
rect 23211 33743 23247 33750
rect 23281 33743 23317 33777
rect 23351 33743 23387 33777
rect 23421 33743 23457 33777
rect 23491 33743 23527 33777
rect 23561 33743 23597 33777
rect 23631 33743 23635 33777
rect 22823 33711 23635 33743
rect 22823 33709 22829 33711
rect 22863 33709 22911 33711
rect 22945 33709 22993 33711
rect 23027 33709 23075 33711
rect 23109 33709 23157 33711
rect 23191 33709 23239 33711
rect 23273 33709 23635 33711
rect 22823 33675 22827 33709
rect 22863 33677 22897 33709
rect 22945 33677 22967 33709
rect 23027 33677 23037 33709
rect 22861 33675 22897 33677
rect 22931 33675 22967 33677
rect 23001 33675 23037 33677
rect 23071 33677 23075 33709
rect 23141 33677 23157 33709
rect 23211 33677 23239 33709
rect 23071 33675 23107 33677
rect 23141 33675 23177 33677
rect 23211 33675 23247 33677
rect 23281 33675 23317 33709
rect 23351 33675 23387 33709
rect 23421 33675 23457 33709
rect 23491 33675 23527 33709
rect 23561 33675 23597 33709
rect 23631 33675 23635 33709
rect 22823 33641 23635 33675
rect 22823 33607 22827 33641
rect 22861 33638 22897 33641
rect 22931 33638 22967 33641
rect 23001 33638 23037 33641
rect 22863 33607 22897 33638
rect 22945 33607 22967 33638
rect 23027 33607 23037 33638
rect 23071 33638 23107 33641
rect 23141 33638 23177 33641
rect 23211 33638 23247 33641
rect 23071 33607 23075 33638
rect 23141 33607 23157 33638
rect 23211 33607 23239 33638
rect 23281 33607 23317 33641
rect 23351 33607 23387 33641
rect 23421 33607 23457 33641
rect 23491 33607 23527 33641
rect 23561 33607 23597 33641
rect 23631 33607 23635 33641
rect 22823 33604 22829 33607
rect 22863 33604 22911 33607
rect 22945 33604 22993 33607
rect 23027 33604 23075 33607
rect 23109 33604 23157 33607
rect 23191 33604 23239 33607
rect 23273 33604 23635 33607
rect 22823 33573 23635 33604
rect 22823 33539 22827 33573
rect 22861 33565 22897 33573
rect 22931 33565 22967 33573
rect 23001 33565 23037 33573
rect 22863 33539 22897 33565
rect 22945 33539 22967 33565
rect 23027 33539 23037 33565
rect 23071 33565 23107 33573
rect 23141 33565 23177 33573
rect 23211 33565 23247 33573
rect 23071 33539 23075 33565
rect 23141 33539 23157 33565
rect 23211 33539 23239 33565
rect 23281 33539 23317 33573
rect 23351 33539 23387 33573
rect 23421 33539 23457 33573
rect 23491 33539 23527 33573
rect 23561 33539 23597 33573
rect 23631 33539 23635 33573
rect 22823 33531 22829 33539
rect 22863 33531 22911 33539
rect 22945 33531 22993 33539
rect 23027 33531 23075 33539
rect 23109 33531 23157 33539
rect 23191 33531 23239 33539
rect 23273 33531 23635 33539
rect 22823 33505 23635 33531
rect 22823 33471 22827 33505
rect 22861 33492 22897 33505
rect 22931 33492 22967 33505
rect 23001 33492 23037 33505
rect 22863 33471 22897 33492
rect 22945 33471 22967 33492
rect 23027 33471 23037 33492
rect 23071 33492 23107 33505
rect 23141 33492 23177 33505
rect 23211 33492 23247 33505
rect 23071 33471 23075 33492
rect 23141 33471 23157 33492
rect 23211 33471 23239 33492
rect 23281 33471 23317 33505
rect 23351 33471 23387 33505
rect 23421 33471 23457 33505
rect 23491 33471 23527 33505
rect 23561 33471 23597 33505
rect 23631 33471 23635 33505
rect 22823 33458 22829 33471
rect 22863 33458 22911 33471
rect 22945 33458 22993 33471
rect 23027 33458 23075 33471
rect 23109 33458 23157 33471
rect 23191 33458 23239 33471
rect 23273 33458 23635 33471
rect 22823 33437 23635 33458
rect 22823 33403 22827 33437
rect 22861 33419 22897 33437
rect 22931 33419 22967 33437
rect 23001 33419 23037 33437
rect 22863 33403 22897 33419
rect 22945 33403 22967 33419
rect 23027 33403 23037 33419
rect 23071 33419 23107 33437
rect 23141 33419 23177 33437
rect 23211 33419 23247 33437
rect 23071 33403 23075 33419
rect 23141 33403 23157 33419
rect 23211 33403 23239 33419
rect 23281 33403 23317 33437
rect 23351 33403 23387 33437
rect 23421 33403 23457 33437
rect 23491 33403 23527 33437
rect 23561 33403 23597 33437
rect 23631 33403 23635 33437
rect 22823 33385 22829 33403
rect 22863 33385 22911 33403
rect 22945 33385 22993 33403
rect 23027 33385 23075 33403
rect 23109 33385 23157 33403
rect 23191 33385 23239 33403
rect 23273 33385 23635 33403
rect 22823 33369 23635 33385
rect 22823 33335 22827 33369
rect 22861 33346 22897 33369
rect 22931 33346 22967 33369
rect 23001 33346 23037 33369
rect 22863 33335 22897 33346
rect 22945 33335 22967 33346
rect 23027 33335 23037 33346
rect 23071 33346 23107 33369
rect 23141 33346 23177 33369
rect 23211 33346 23247 33369
rect 23071 33335 23075 33346
rect 23141 33335 23157 33346
rect 23211 33335 23239 33346
rect 23281 33335 23317 33369
rect 23351 33335 23387 33369
rect 23421 33335 23457 33369
rect 23491 33335 23527 33369
rect 23561 33335 23597 33369
rect 23631 33335 23635 33369
rect 18022 33328 18442 33331
rect 203 33310 331 33316
rect 203 33276 209 33310
rect 243 33281 291 33310
rect 243 33276 278 33281
rect 325 33276 331 33310
rect 203 33247 278 33276
rect 312 33247 331 33276
rect 203 33237 331 33247
rect 203 33203 209 33237
rect 243 33212 291 33237
rect 243 33203 278 33212
rect 325 33203 331 33237
rect 203 33178 278 33203
rect 312 33178 331 33203
rect 203 33164 331 33178
rect 203 33130 209 33164
rect 243 33143 291 33164
rect 243 33130 278 33143
rect 325 33130 331 33164
rect 203 33109 278 33130
rect 312 33109 331 33130
rect 203 33091 331 33109
rect 203 33057 209 33091
rect 243 33074 291 33091
rect 243 33057 278 33074
rect 325 33057 331 33091
rect 203 33040 278 33057
rect 312 33040 331 33057
rect 203 33018 331 33040
rect 203 32984 209 33018
rect 243 33005 291 33018
rect 243 32984 278 33005
rect 325 32984 331 33018
rect 203 32971 278 32984
rect 312 32971 331 32984
rect 203 32945 331 32971
rect 203 32911 209 32945
rect 243 32936 291 32945
rect 243 32911 278 32936
rect 325 32911 331 32945
rect 203 32902 278 32911
rect 312 32902 331 32911
rect 203 32872 331 32902
rect 203 32838 209 32872
rect 243 32867 291 32872
rect 243 32838 278 32867
rect 325 32838 331 32872
rect 203 32833 278 32838
rect 312 32833 331 32838
rect 203 32799 331 32833
rect 203 32765 209 32799
rect 243 32798 291 32799
rect 243 32765 278 32798
rect 325 32765 331 32799
rect 203 32764 278 32765
rect 312 32764 331 32765
rect 203 32729 331 32764
rect 203 32726 278 32729
rect 312 32726 331 32729
rect 203 32692 209 32726
rect 243 32695 278 32726
rect 243 32692 291 32695
rect 325 32692 331 32726
rect 203 32660 331 32692
rect 203 32653 278 32660
rect 312 32653 331 32660
rect 203 32619 209 32653
rect 243 32626 278 32653
rect 243 32619 291 32626
rect 325 32619 331 32653
rect 203 32591 331 32619
rect 203 32580 278 32591
rect 312 32580 331 32591
rect 203 32546 209 32580
rect 243 32557 278 32580
rect 243 32546 291 32557
rect 325 32546 331 32580
rect 203 32522 331 32546
rect 203 32507 278 32522
rect 312 32507 331 32522
rect 203 32473 209 32507
rect 243 32488 278 32507
rect 243 32473 291 32488
rect 325 32473 331 32507
rect 203 32453 331 32473
rect 203 32434 278 32453
rect 312 32434 331 32453
rect 203 32400 209 32434
rect 243 32419 278 32434
rect 243 32400 291 32419
rect 325 32400 331 32434
rect 203 32384 331 32400
rect 203 32361 278 32384
rect 312 32361 331 32384
rect 203 32327 209 32361
rect 243 32350 278 32361
rect 243 32327 291 32350
rect 325 32327 331 32361
rect 203 32316 331 32327
rect 18021 33294 18022 33328
rect 18056 33307 18108 33328
rect 18142 33307 18194 33328
rect 18228 33307 18280 33328
rect 18314 33307 18366 33328
rect 18021 33273 18025 33294
rect 18059 33273 18101 33307
rect 18142 33294 18177 33307
rect 18228 33294 18253 33307
rect 18314 33294 18329 33307
rect 18135 33273 18177 33294
rect 18211 33273 18253 33294
rect 18287 33273 18329 33294
rect 18363 33294 18366 33307
rect 18400 33307 18442 33328
rect 18400 33294 18405 33307
rect 18363 33273 18405 33294
rect 18439 33273 18442 33307
rect 18021 33256 18442 33273
rect 18021 33222 18022 33256
rect 18056 33239 18108 33256
rect 18142 33239 18194 33256
rect 18228 33239 18280 33256
rect 18314 33239 18366 33256
rect 18021 33205 18025 33222
rect 18059 33205 18101 33239
rect 18142 33222 18177 33239
rect 18228 33222 18253 33239
rect 18314 33222 18329 33239
rect 18135 33205 18177 33222
rect 18211 33205 18253 33222
rect 18287 33205 18329 33222
rect 18363 33222 18366 33239
rect 18400 33239 18442 33256
rect 18400 33222 18405 33239
rect 18363 33205 18405 33222
rect 18439 33205 18442 33239
rect 18021 33184 18442 33205
rect 18021 33150 18022 33184
rect 18056 33171 18108 33184
rect 18142 33171 18194 33184
rect 18228 33171 18280 33184
rect 18314 33171 18366 33184
rect 18021 33137 18025 33150
rect 18059 33137 18101 33171
rect 18142 33150 18177 33171
rect 18228 33150 18253 33171
rect 18314 33150 18329 33171
rect 18135 33137 18177 33150
rect 18211 33137 18253 33150
rect 18287 33137 18329 33150
rect 18363 33150 18366 33171
rect 18400 33171 18442 33184
rect 18400 33150 18405 33171
rect 18363 33137 18405 33150
rect 18439 33137 18442 33171
rect 18021 33112 18442 33137
rect 18021 33078 18022 33112
rect 18056 33103 18108 33112
rect 18142 33103 18194 33112
rect 18228 33103 18280 33112
rect 18314 33103 18366 33112
rect 18021 33069 18025 33078
rect 18059 33069 18101 33103
rect 18142 33078 18177 33103
rect 18228 33078 18253 33103
rect 18314 33078 18329 33103
rect 18135 33069 18177 33078
rect 18211 33069 18253 33078
rect 18287 33069 18329 33078
rect 18363 33078 18366 33103
rect 18400 33103 18442 33112
rect 18400 33078 18405 33103
rect 18363 33069 18405 33078
rect 18439 33069 18442 33103
rect 18021 33040 18442 33069
rect 18021 33006 18022 33040
rect 18056 33035 18108 33040
rect 18142 33035 18194 33040
rect 18228 33035 18280 33040
rect 18314 33035 18366 33040
rect 18021 33001 18025 33006
rect 18059 33001 18101 33035
rect 18142 33006 18177 33035
rect 18228 33006 18253 33035
rect 18314 33006 18329 33035
rect 18135 33001 18177 33006
rect 18211 33001 18253 33006
rect 18287 33001 18329 33006
rect 18363 33006 18366 33035
rect 18400 33035 18442 33040
rect 18400 33006 18405 33035
rect 18363 33001 18405 33006
rect 18439 33001 18442 33035
rect 18021 32968 18442 33001
rect 18021 32934 18022 32968
rect 18056 32967 18108 32968
rect 18142 32967 18194 32968
rect 18228 32967 18280 32968
rect 18314 32967 18366 32968
rect 18021 32933 18025 32934
rect 18059 32933 18101 32967
rect 18142 32934 18177 32967
rect 18228 32934 18253 32967
rect 18314 32934 18329 32967
rect 18135 32933 18177 32934
rect 18211 32933 18253 32934
rect 18287 32933 18329 32934
rect 18363 32934 18366 32967
rect 18400 32967 18442 32968
rect 18400 32934 18405 32967
rect 18363 32933 18405 32934
rect 18439 32933 18442 32967
rect 18021 32899 18442 32933
rect 18021 32896 18025 32899
rect 18021 32862 18022 32896
rect 18059 32865 18101 32899
rect 18135 32896 18177 32899
rect 18211 32896 18253 32899
rect 18287 32896 18329 32899
rect 18142 32865 18177 32896
rect 18228 32865 18253 32896
rect 18314 32865 18329 32896
rect 18363 32896 18405 32899
rect 18363 32865 18366 32896
rect 18056 32862 18108 32865
rect 18142 32862 18194 32865
rect 18228 32862 18280 32865
rect 18314 32862 18366 32865
rect 18400 32865 18405 32896
rect 18439 32865 18442 32899
rect 18400 32862 18442 32865
rect 18021 32831 18442 32862
rect 18021 32824 18025 32831
rect 18021 32790 18022 32824
rect 18059 32797 18101 32831
rect 18135 32824 18177 32831
rect 18211 32824 18253 32831
rect 18287 32824 18329 32831
rect 18142 32797 18177 32824
rect 18228 32797 18253 32824
rect 18314 32797 18329 32824
rect 18363 32824 18405 32831
rect 18363 32797 18366 32824
rect 18056 32790 18108 32797
rect 18142 32790 18194 32797
rect 18228 32790 18280 32797
rect 18314 32790 18366 32797
rect 18400 32797 18405 32824
rect 18439 32797 18442 32831
rect 18400 32790 18442 32797
rect 18021 32763 18442 32790
rect 18021 32752 18025 32763
rect 18021 32718 18022 32752
rect 18059 32729 18101 32763
rect 18135 32752 18177 32763
rect 18211 32752 18253 32763
rect 18287 32752 18329 32763
rect 18142 32729 18177 32752
rect 18228 32729 18253 32752
rect 18314 32729 18329 32752
rect 18363 32752 18405 32763
rect 18363 32729 18366 32752
rect 18056 32718 18108 32729
rect 18142 32718 18194 32729
rect 18228 32718 18280 32729
rect 18314 32718 18366 32729
rect 18400 32729 18405 32752
rect 18439 32729 18442 32763
rect 18400 32718 18442 32729
rect 18021 32695 18442 32718
rect 18021 32680 18025 32695
rect 18021 32646 18022 32680
rect 18059 32661 18101 32695
rect 18135 32680 18177 32695
rect 18211 32680 18253 32695
rect 18287 32680 18329 32695
rect 18142 32661 18177 32680
rect 18228 32661 18253 32680
rect 18314 32661 18329 32680
rect 18363 32680 18405 32695
rect 18363 32661 18366 32680
rect 18056 32646 18108 32661
rect 18142 32646 18194 32661
rect 18228 32646 18280 32661
rect 18314 32646 18366 32661
rect 18400 32661 18405 32680
rect 18439 32661 18442 32695
rect 18400 32646 18442 32661
rect 18021 32627 18442 32646
rect 18021 32608 18025 32627
rect 18021 32574 18022 32608
rect 18059 32593 18101 32627
rect 18135 32608 18177 32627
rect 18211 32608 18253 32627
rect 18287 32608 18329 32627
rect 18142 32593 18177 32608
rect 18228 32593 18253 32608
rect 18314 32593 18329 32608
rect 18363 32608 18405 32627
rect 18363 32593 18366 32608
rect 18056 32574 18108 32593
rect 18142 32574 18194 32593
rect 18228 32574 18280 32593
rect 18314 32574 18366 32593
rect 18400 32593 18405 32608
rect 18439 32593 18442 32627
rect 18400 32574 18442 32593
rect 18021 32559 18442 32574
rect 18021 32536 18025 32559
rect 18021 32502 18022 32536
rect 18059 32525 18101 32559
rect 18135 32536 18177 32559
rect 18211 32536 18253 32559
rect 18287 32536 18329 32559
rect 18142 32525 18177 32536
rect 18228 32525 18253 32536
rect 18314 32525 18329 32536
rect 18363 32536 18405 32559
rect 18363 32525 18366 32536
rect 18056 32502 18108 32525
rect 18142 32502 18194 32525
rect 18228 32502 18280 32525
rect 18314 32502 18366 32525
rect 18400 32525 18405 32536
rect 18439 32525 18442 32559
rect 18400 32502 18442 32525
rect 18021 32491 18442 32502
rect 18021 32464 18025 32491
rect 18021 32430 18022 32464
rect 18059 32457 18101 32491
rect 18135 32464 18177 32491
rect 18211 32464 18253 32491
rect 18287 32464 18329 32491
rect 18142 32457 18177 32464
rect 18228 32457 18253 32464
rect 18314 32457 18329 32464
rect 18363 32464 18405 32491
rect 18363 32457 18366 32464
rect 18056 32430 18108 32457
rect 18142 32430 18194 32457
rect 18228 32430 18280 32457
rect 18314 32430 18366 32457
rect 18400 32457 18405 32464
rect 18439 32457 18442 32491
rect 18400 32430 18442 32457
rect 18021 32423 18442 32430
rect 18021 32392 18025 32423
rect 18021 32358 18022 32392
rect 18059 32389 18101 32423
rect 18135 32392 18177 32423
rect 18211 32392 18253 32423
rect 18287 32392 18329 32423
rect 18142 32389 18177 32392
rect 18228 32389 18253 32392
rect 18314 32389 18329 32392
rect 18363 32392 18405 32423
rect 18363 32389 18366 32392
rect 18056 32358 18108 32389
rect 18142 32358 18194 32389
rect 18228 32358 18280 32389
rect 18314 32358 18366 32389
rect 18400 32389 18405 32392
rect 18439 32389 18442 32423
rect 18400 32358 18442 32389
rect 18021 32355 18442 32358
rect 18021 32321 18025 32355
rect 18059 32321 18101 32355
rect 18135 32321 18177 32355
rect 18211 32321 18253 32355
rect 18287 32321 18329 32355
rect 18363 32321 18405 32355
rect 18439 32321 18442 32355
rect 18021 32320 18442 32321
rect 203 32315 912 32316
rect 203 32288 278 32315
rect 312 32288 912 32315
rect 203 32254 209 32288
rect 243 32281 278 32288
rect 325 32282 912 32288
rect 243 32254 291 32281
rect 325 32254 368 32282
rect 203 32248 368 32254
rect 402 32248 440 32282
rect 474 32248 512 32282
rect 546 32248 584 32282
rect 618 32248 656 32282
rect 690 32248 728 32282
rect 762 32248 800 32282
rect 834 32248 872 32282
rect 906 32248 912 32282
rect 203 32246 912 32248
rect 203 32215 278 32246
rect 312 32215 912 32246
rect 203 32181 209 32215
rect 243 32212 278 32215
rect 243 32181 291 32212
rect 325 32206 912 32215
rect 325 32181 368 32206
rect 203 32177 368 32181
rect 203 32143 278 32177
rect 312 32172 368 32177
rect 402 32172 440 32206
rect 474 32172 512 32206
rect 546 32172 584 32206
rect 618 32172 656 32206
rect 690 32172 728 32206
rect 762 32172 800 32206
rect 834 32172 872 32206
rect 906 32172 912 32206
rect 312 32143 912 32172
rect 203 32142 912 32143
rect 203 32108 209 32142
rect 243 32108 291 32142
rect 325 32130 912 32142
rect 325 32108 368 32130
rect 203 32074 278 32108
rect 312 32096 368 32108
rect 402 32096 440 32130
rect 474 32096 512 32130
rect 546 32096 584 32130
rect 618 32096 656 32130
rect 690 32096 728 32130
rect 762 32096 800 32130
rect 834 32096 872 32130
rect 906 32096 912 32130
rect 312 32074 912 32096
rect 203 32064 912 32074
rect 203 32030 218 32064
rect 252 32054 912 32064
rect 252 32039 368 32054
rect 252 32030 278 32039
rect 203 32005 278 32030
rect 312 32020 368 32039
rect 402 32020 440 32054
rect 474 32020 512 32054
rect 546 32020 584 32054
rect 618 32020 656 32054
rect 690 32020 728 32054
rect 762 32020 800 32054
rect 834 32020 872 32054
rect 906 32020 912 32054
rect 312 32005 912 32020
rect 203 31992 912 32005
rect 203 31958 218 31992
rect 252 31978 912 31992
rect 252 31970 368 31978
rect 252 31958 278 31970
rect 203 31936 278 31958
rect 312 31944 368 31970
rect 402 31944 440 31978
rect 474 31944 512 31978
rect 546 31944 584 31978
rect 618 31944 656 31978
rect 690 31944 728 31978
rect 762 31944 800 31978
rect 834 31944 872 31978
rect 906 31944 912 31978
rect 312 31936 912 31944
rect 203 31920 912 31936
rect 203 31886 218 31920
rect 252 31902 912 31920
rect 252 31901 368 31902
rect 252 31886 278 31901
rect 203 31867 278 31886
rect 312 31868 368 31901
rect 402 31868 440 31902
rect 474 31868 512 31902
rect 546 31868 584 31902
rect 618 31868 656 31902
rect 690 31868 728 31902
rect 762 31868 800 31902
rect 834 31868 872 31902
rect 906 31868 912 31902
rect 312 31867 912 31868
rect 203 31848 912 31867
rect 203 31814 218 31848
rect 252 31832 912 31848
rect 252 31814 278 31832
rect 203 31798 278 31814
rect 312 31825 912 31832
rect 312 31798 368 31825
rect 203 31791 368 31798
rect 402 31791 440 31825
rect 474 31791 512 31825
rect 546 31791 584 31825
rect 618 31791 656 31825
rect 690 31791 728 31825
rect 762 31791 800 31825
rect 834 31791 872 31825
rect 906 31791 912 31825
rect 203 31776 912 31791
rect 203 31742 218 31776
rect 252 31763 912 31776
rect 252 31742 278 31763
rect 203 31729 278 31742
rect 312 31729 912 31763
rect 203 31705 912 31729
rect 18021 32286 18022 32320
rect 18056 32287 18108 32320
rect 18142 32287 18194 32320
rect 18228 32287 18280 32320
rect 18314 32287 18366 32320
rect 18021 32253 18025 32286
rect 18059 32253 18101 32287
rect 18142 32286 18177 32287
rect 18228 32286 18253 32287
rect 18314 32286 18329 32287
rect 18135 32253 18177 32286
rect 18211 32253 18253 32286
rect 18287 32253 18329 32286
rect 18363 32286 18366 32287
rect 18400 32287 18442 32320
rect 18400 32286 18405 32287
rect 18363 32253 18405 32286
rect 18439 32253 18442 32287
rect 18021 32248 18442 32253
rect 18021 32214 18022 32248
rect 18056 32219 18108 32248
rect 18142 32219 18194 32248
rect 18228 32219 18280 32248
rect 18314 32219 18366 32248
rect 18021 32185 18025 32214
rect 18059 32185 18101 32219
rect 18142 32214 18177 32219
rect 18228 32214 18253 32219
rect 18314 32214 18329 32219
rect 18135 32185 18177 32214
rect 18211 32185 18253 32214
rect 18287 32185 18329 32214
rect 18363 32214 18366 32219
rect 18400 32219 18442 32248
rect 18400 32214 18405 32219
rect 18363 32185 18405 32214
rect 18439 32185 18442 32219
rect 18021 32176 18442 32185
rect 18021 32142 18022 32176
rect 18056 32151 18108 32176
rect 18142 32151 18194 32176
rect 18228 32151 18280 32176
rect 18314 32151 18366 32176
rect 18021 32117 18025 32142
rect 18059 32117 18101 32151
rect 18142 32142 18177 32151
rect 18228 32142 18253 32151
rect 18314 32142 18329 32151
rect 18135 32117 18177 32142
rect 18211 32117 18253 32142
rect 18287 32117 18329 32142
rect 18363 32142 18366 32151
rect 18400 32151 18442 32176
rect 18400 32142 18405 32151
rect 18363 32117 18405 32142
rect 18439 32117 18442 32151
rect 18021 32104 18442 32117
rect 18021 32070 18022 32104
rect 18056 32083 18108 32104
rect 18142 32083 18194 32104
rect 18228 32083 18280 32104
rect 18314 32083 18366 32104
rect 18021 32049 18025 32070
rect 18059 32049 18101 32083
rect 18142 32070 18177 32083
rect 18228 32070 18253 32083
rect 18314 32070 18329 32083
rect 18135 32049 18177 32070
rect 18211 32049 18253 32070
rect 18287 32049 18329 32070
rect 18363 32070 18366 32083
rect 18400 32083 18442 32104
rect 18400 32070 18405 32083
rect 18363 32049 18405 32070
rect 18439 32049 18442 32083
rect 18021 32032 18442 32049
rect 18021 31998 18022 32032
rect 18056 32015 18108 32032
rect 18142 32015 18194 32032
rect 18228 32015 18280 32032
rect 18314 32015 18366 32032
rect 18021 31981 18025 31998
rect 18059 31981 18101 32015
rect 18142 31998 18177 32015
rect 18228 31998 18253 32015
rect 18314 31998 18329 32015
rect 18135 31981 18177 31998
rect 18211 31981 18253 31998
rect 18287 31981 18329 31998
rect 18363 31998 18366 32015
rect 18400 32015 18442 32032
rect 18400 31998 18405 32015
rect 18363 31981 18405 31998
rect 18439 31981 18442 32015
rect 18021 31960 18442 31981
rect 18021 31926 18022 31960
rect 18056 31947 18108 31960
rect 18142 31947 18194 31960
rect 18228 31947 18280 31960
rect 18314 31947 18366 31960
rect 18021 31913 18025 31926
rect 18059 31913 18101 31947
rect 18142 31926 18177 31947
rect 18228 31926 18253 31947
rect 18314 31926 18329 31947
rect 18135 31913 18177 31926
rect 18211 31913 18253 31926
rect 18287 31913 18329 31926
rect 18363 31926 18366 31947
rect 18400 31947 18442 31960
rect 18400 31926 18405 31947
rect 18363 31913 18405 31926
rect 18439 31913 18442 31947
rect 18021 31888 18442 31913
rect 18021 31854 18022 31888
rect 18056 31879 18108 31888
rect 18142 31879 18194 31888
rect 18228 31879 18280 31888
rect 18314 31879 18366 31888
rect 18021 31845 18025 31854
rect 18059 31845 18101 31879
rect 18142 31854 18177 31879
rect 18228 31854 18253 31879
rect 18314 31854 18329 31879
rect 18135 31845 18177 31854
rect 18211 31845 18253 31854
rect 18287 31845 18329 31854
rect 18363 31854 18366 31879
rect 18400 31879 18442 31888
rect 18400 31854 18405 31879
rect 18363 31845 18405 31854
rect 18439 31845 18442 31879
rect 18021 31816 18442 31845
rect 18021 31782 18022 31816
rect 18056 31811 18108 31816
rect 18142 31811 18194 31816
rect 18228 31811 18280 31816
rect 18314 31811 18366 31816
rect 18021 31777 18025 31782
rect 18059 31777 18101 31811
rect 18142 31782 18177 31811
rect 18228 31782 18253 31811
rect 18314 31782 18329 31811
rect 18135 31777 18177 31782
rect 18211 31777 18253 31782
rect 18287 31777 18329 31782
rect 18363 31782 18366 31811
rect 18400 31811 18442 31816
rect 18400 31782 18405 31811
rect 18363 31777 18405 31782
rect 18439 31777 18442 31811
rect 18021 31744 18442 31777
rect 18021 31710 18022 31744
rect 18056 31743 18108 31744
rect 18142 31743 18194 31744
rect 18228 31743 18280 31744
rect 18314 31743 18366 31744
rect 18021 31709 18025 31710
rect 18059 31709 18101 31743
rect 18142 31710 18177 31743
rect 18228 31710 18253 31743
rect 18314 31710 18329 31743
rect 18135 31709 18177 31710
rect 18211 31709 18253 31710
rect 18287 31709 18329 31710
rect 18363 31710 18366 31743
rect 18400 31743 18442 31744
rect 18400 31710 18405 31743
rect 18363 31709 18405 31710
rect 18439 31709 18442 31743
rect 203 31704 332 31705
rect 203 31670 218 31704
rect 252 31670 332 31704
rect 203 31632 332 31670
rect 203 31598 218 31632
rect 252 31598 332 31632
rect 203 31560 332 31598
rect 203 31526 218 31560
rect 252 31526 332 31560
rect 203 31488 332 31526
rect 203 31454 218 31488
rect 252 31454 332 31488
rect 203 31416 332 31454
rect 203 31382 218 31416
rect 252 31382 332 31416
rect 203 31344 332 31382
rect 203 31310 218 31344
rect 252 31310 332 31344
rect 203 31272 332 31310
rect 203 31238 218 31272
rect 252 31238 332 31272
rect 203 31200 332 31238
rect 203 31166 218 31200
rect 252 31166 332 31200
rect 203 31128 332 31166
rect 203 31094 218 31128
rect 252 31094 332 31128
rect 203 31056 332 31094
rect 203 31022 218 31056
rect 252 31022 332 31056
rect 203 30984 332 31022
rect 203 30950 218 30984
rect 252 30950 332 30984
rect 203 30912 332 30950
rect 203 30878 218 30912
rect 252 30878 332 30912
rect 203 30840 332 30878
rect 203 30806 218 30840
rect 252 30806 332 30840
rect 203 30768 332 30806
rect 203 30734 218 30768
rect 252 30734 332 30768
rect 203 30696 332 30734
rect 203 30662 218 30696
rect 252 30662 332 30696
rect 203 30624 332 30662
rect 203 30590 218 30624
rect 252 30590 332 30624
rect 203 30552 332 30590
rect 203 30518 218 30552
rect 252 30518 332 30552
rect 203 30480 332 30518
rect 203 30446 218 30480
rect 252 30446 332 30480
rect 203 30408 332 30446
rect 203 30374 218 30408
rect 252 30374 332 30408
rect 203 30336 332 30374
rect 203 30302 218 30336
rect 252 30302 332 30336
rect 203 30264 332 30302
rect 203 30230 218 30264
rect 252 30230 332 30264
rect 203 30192 332 30230
rect 203 30158 218 30192
rect 252 30158 332 30192
rect 203 30120 332 30158
rect 203 30086 218 30120
rect 252 30086 332 30120
rect 203 30048 332 30086
rect 203 30014 218 30048
rect 252 30014 332 30048
rect 203 29976 332 30014
rect 203 29942 218 29976
rect 252 29942 332 29976
rect 203 29904 332 29942
rect 203 29870 218 29904
rect 252 29870 332 29904
rect 203 29832 332 29870
rect 203 29798 218 29832
rect 252 29798 332 29832
rect 203 29760 332 29798
rect 203 29726 218 29760
rect 252 29726 332 29760
rect 203 29688 332 29726
rect 203 29654 218 29688
rect 252 29654 332 29688
rect 203 29616 332 29654
rect 203 29582 218 29616
rect 252 29582 332 29616
rect 203 29544 332 29582
rect 203 29510 218 29544
rect 252 29510 332 29544
rect 203 29472 332 29510
rect 203 29438 218 29472
rect 252 29438 332 29472
rect 203 29400 332 29438
rect 203 29366 218 29400
rect 252 29366 332 29400
rect 203 29328 332 29366
rect 203 29294 218 29328
rect 252 29294 332 29328
rect 203 29256 332 29294
rect 203 29222 218 29256
rect 252 29222 332 29256
rect 203 29184 332 29222
rect 203 29150 218 29184
rect 252 29150 332 29184
rect 203 29112 332 29150
rect 203 29078 218 29112
rect 252 29078 332 29112
rect 203 29040 332 29078
rect 203 29006 218 29040
rect 252 29006 332 29040
rect 203 28968 332 29006
rect 203 28934 218 28968
rect 252 28934 332 28968
rect 203 28896 332 28934
rect 203 28862 218 28896
rect 252 28862 332 28896
rect 203 28824 332 28862
rect 203 28790 218 28824
rect 252 28790 332 28824
rect 203 28752 332 28790
rect 203 28718 218 28752
rect 252 28718 332 28752
rect 203 28680 332 28718
rect 203 28646 218 28680
rect 252 28646 332 28680
rect 203 28608 332 28646
rect 203 28574 218 28608
rect 252 28574 332 28608
rect 203 28535 332 28574
rect 203 28501 218 28535
rect 252 28501 332 28535
rect 203 28462 332 28501
rect 203 28428 218 28462
rect 252 28428 332 28462
rect 203 28389 332 28428
rect 203 28355 218 28389
rect 252 28355 332 28389
rect 203 28316 332 28355
rect 203 28282 218 28316
rect 252 28282 332 28316
rect 203 28243 332 28282
rect 203 28209 218 28243
rect 252 28209 332 28243
rect 203 28170 332 28209
rect 203 28136 218 28170
rect 252 28136 332 28170
rect 203 28097 332 28136
rect 203 28063 218 28097
rect 252 28063 332 28097
rect 203 28024 332 28063
rect 203 27990 218 28024
rect 252 27990 332 28024
rect 203 27951 332 27990
rect 203 27917 218 27951
rect 252 27917 332 27951
rect 203 27878 332 27917
rect 203 27844 218 27878
rect 252 27844 332 27878
rect 203 27805 332 27844
rect 203 27771 218 27805
rect 252 27771 332 27805
rect 203 27732 332 27771
rect 203 27698 218 27732
rect 252 27698 332 27732
rect 203 27659 332 27698
rect 203 27625 218 27659
rect 252 27625 332 27659
rect 203 27586 332 27625
rect 203 27552 218 27586
rect 252 27552 332 27586
rect 203 27513 332 27552
rect 203 27479 218 27513
rect 252 27479 332 27513
rect 203 27440 332 27479
rect 203 27406 218 27440
rect 252 27406 332 27440
rect 203 27367 332 27406
rect 203 27333 218 27367
rect 252 27333 332 27367
rect 203 27294 332 27333
rect 203 27260 218 27294
rect 252 27260 332 27294
rect 203 27221 332 27260
rect 203 27187 218 27221
rect 252 27187 332 27221
rect 203 27148 332 27187
rect 203 27114 218 27148
rect 252 27114 332 27148
rect 203 27075 332 27114
rect 203 27041 218 27075
rect 252 27041 332 27075
rect 203 27002 332 27041
rect 203 26968 218 27002
rect 252 26968 332 27002
rect 203 26929 332 26968
rect 203 26895 218 26929
rect 252 26895 332 26929
rect 203 26856 332 26895
rect 203 26822 218 26856
rect 252 26822 332 26856
rect 203 26783 332 26822
rect 203 26749 218 26783
rect 252 26749 332 26783
rect 203 26710 332 26749
rect 203 26676 218 26710
rect 252 26676 332 26710
rect 203 26637 332 26676
rect 203 26603 218 26637
rect 252 26603 332 26637
rect 203 26564 332 26603
rect 203 26530 218 26564
rect 252 26530 332 26564
rect 203 26491 332 26530
rect 203 26457 218 26491
rect 252 26457 332 26491
rect 203 26418 332 26457
rect 203 26384 218 26418
rect 252 26384 332 26418
rect 203 26345 332 26384
rect 203 26311 218 26345
rect 252 26311 332 26345
rect 203 26272 332 26311
rect 203 26238 218 26272
rect 252 26238 332 26272
rect 203 26199 332 26238
rect 203 26165 218 26199
rect 252 26165 332 26199
rect 203 26126 332 26165
rect 203 26092 218 26126
rect 252 26092 332 26126
rect 203 26053 332 26092
rect 203 26019 218 26053
rect 252 26019 332 26053
rect 203 25980 332 26019
rect 203 25946 218 25980
rect 252 25946 332 25980
rect 203 25907 332 25946
rect 203 25873 218 25907
rect 252 25873 332 25907
rect 203 25834 332 25873
rect 203 25800 218 25834
rect 252 25800 332 25834
rect 203 25761 332 25800
rect 203 25727 218 25761
rect 252 25727 332 25761
rect 203 25688 332 25727
rect 203 25654 218 25688
rect 252 25654 332 25688
rect 203 25615 332 25654
rect 203 25581 218 25615
rect 252 25581 332 25615
rect 203 25542 332 25581
rect 203 25508 218 25542
rect 252 25508 332 25542
rect 203 25469 332 25508
rect 203 25435 218 25469
rect 252 25435 332 25469
rect 203 25396 332 25435
rect 203 25362 218 25396
rect 252 25362 332 25396
rect 203 25323 332 25362
rect 203 25289 218 25323
rect 252 25289 332 25323
rect 203 25250 332 25289
rect 203 25216 218 25250
rect 252 25216 332 25250
rect 203 25177 332 25216
rect 203 25143 218 25177
rect 252 25143 332 25177
rect 203 25104 332 25143
rect 203 25070 218 25104
rect 252 25070 332 25104
rect 203 25031 332 25070
rect 203 24997 218 25031
rect 252 24997 332 25031
rect 203 24958 332 24997
rect 203 24924 218 24958
rect 252 24924 332 24958
rect 203 24885 332 24924
rect 203 24851 218 24885
rect 252 24851 332 24885
rect 203 24812 332 24851
rect 203 24778 218 24812
rect 252 24778 332 24812
rect 203 24739 332 24778
rect 203 24705 218 24739
rect 252 24705 332 24739
rect 203 24666 332 24705
rect 203 24632 218 24666
rect 252 24632 332 24666
rect 203 24593 332 24632
rect 203 24559 218 24593
rect 252 24559 332 24593
rect 203 24520 332 24559
rect 203 24486 218 24520
rect 252 24486 332 24520
rect 203 24447 332 24486
rect 203 24413 218 24447
rect 252 24413 332 24447
rect 203 24374 332 24413
rect 203 24340 218 24374
rect 252 24340 332 24374
rect 203 24301 332 24340
rect 203 24267 218 24301
rect 252 24267 332 24301
rect 203 24228 332 24267
rect 203 24194 218 24228
rect 252 24194 332 24228
rect 203 24155 332 24194
rect 203 24121 218 24155
rect 252 24121 332 24155
rect 203 24082 332 24121
rect 203 24048 218 24082
rect 252 24048 332 24082
rect 203 24009 332 24048
rect 203 23975 218 24009
rect 252 23975 332 24009
rect 203 23936 332 23975
rect 203 23902 218 23936
rect 252 23902 332 23936
rect 203 23863 332 23902
rect 203 23829 218 23863
rect 252 23829 332 23863
rect 999 31671 1313 31705
rect 999 31637 1051 31671
rect 1085 31637 1127 31671
rect 1161 31637 1203 31671
rect 1237 31637 1279 31671
rect 999 31603 1313 31637
rect 999 31569 1051 31603
rect 1085 31569 1127 31603
rect 1161 31569 1203 31603
rect 1237 31569 1279 31603
rect 999 31535 1313 31569
rect 999 31501 1051 31535
rect 1085 31501 1127 31535
rect 1161 31501 1203 31535
rect 1237 31501 1279 31535
rect 999 31467 1313 31501
rect 999 31433 1051 31467
rect 1085 31433 1127 31467
rect 1161 31433 1203 31467
rect 1237 31433 1279 31467
rect 999 31399 1313 31433
rect 999 31365 1051 31399
rect 1085 31365 1127 31399
rect 1161 31365 1203 31399
rect 1237 31365 1279 31399
rect 999 31331 1313 31365
rect 999 31297 1051 31331
rect 1085 31297 1127 31331
rect 1161 31297 1203 31331
rect 1237 31297 1279 31331
rect 999 31263 1313 31297
rect 999 31229 1051 31263
rect 1085 31229 1127 31263
rect 1161 31229 1203 31263
rect 1237 31229 1279 31263
rect 999 31195 1313 31229
rect 999 31161 1051 31195
rect 1085 31161 1127 31195
rect 1161 31161 1203 31195
rect 1237 31161 1279 31195
rect 999 31127 1313 31161
rect 999 31093 1051 31127
rect 1085 31093 1127 31127
rect 1161 31093 1203 31127
rect 1237 31093 1279 31127
rect 999 31059 1313 31093
rect 999 31025 1051 31059
rect 1085 31025 1127 31059
rect 1161 31025 1203 31059
rect 1237 31025 1279 31059
rect 999 30991 1313 31025
rect 999 30957 1051 30991
rect 1085 30957 1127 30991
rect 1161 30957 1203 30991
rect 1237 30957 1279 30991
rect 999 30923 1313 30957
rect 999 30889 1051 30923
rect 1085 30889 1127 30923
rect 1161 30889 1203 30923
rect 1237 30889 1279 30923
rect 999 30855 1313 30889
rect 999 30821 1051 30855
rect 1085 30821 1127 30855
rect 1161 30821 1203 30855
rect 1237 30821 1279 30855
rect 999 30787 1313 30821
rect 999 30753 1051 30787
rect 1085 30753 1127 30787
rect 1161 30753 1203 30787
rect 1237 30753 1279 30787
rect 999 30719 1313 30753
rect 999 30685 1051 30719
rect 1085 30685 1127 30719
rect 1161 30685 1203 30719
rect 1237 30685 1279 30719
rect 999 30651 1313 30685
rect 999 30617 1051 30651
rect 1085 30617 1127 30651
rect 1161 30617 1203 30651
rect 1237 30617 1279 30651
rect 999 30583 1313 30617
rect 999 30549 1051 30583
rect 1085 30549 1127 30583
rect 1161 30549 1203 30583
rect 1237 30549 1279 30583
rect 999 30515 1313 30549
rect 999 30481 1051 30515
rect 1085 30481 1127 30515
rect 1161 30481 1203 30515
rect 1237 30481 1279 30515
rect 999 30447 1313 30481
rect 999 30413 1051 30447
rect 1085 30413 1127 30447
rect 1161 30413 1203 30447
rect 1237 30413 1279 30447
rect 999 30379 1313 30413
rect 999 30345 1051 30379
rect 1085 30345 1127 30379
rect 1161 30345 1203 30379
rect 1237 30345 1279 30379
rect 999 30311 1313 30345
rect 999 30277 1051 30311
rect 1085 30277 1127 30311
rect 1161 30277 1203 30311
rect 1237 30277 1279 30311
rect 999 30243 1313 30277
rect 999 30209 1051 30243
rect 1085 30209 1127 30243
rect 1161 30209 1203 30243
rect 1237 30209 1279 30243
rect 999 30175 1313 30209
rect 999 30141 1051 30175
rect 1085 30141 1127 30175
rect 1161 30141 1203 30175
rect 1237 30141 1279 30175
rect 999 30107 1313 30141
rect 999 30073 1051 30107
rect 1085 30073 1127 30107
rect 1161 30073 1203 30107
rect 1237 30073 1279 30107
rect 999 30039 1313 30073
rect 999 30005 1051 30039
rect 1085 30005 1127 30039
rect 1161 30005 1203 30039
rect 1237 30005 1279 30039
rect 999 29971 1313 30005
rect 999 29937 1051 29971
rect 1085 29937 1127 29971
rect 1161 29937 1203 29971
rect 1237 29937 1279 29971
rect 999 29903 1313 29937
rect 999 29869 1051 29903
rect 1085 29869 1127 29903
rect 1161 29869 1203 29903
rect 1237 29869 1279 29903
rect 999 29835 1313 29869
rect 999 29801 1051 29835
rect 1085 29801 1127 29835
rect 1161 29801 1203 29835
rect 1237 29801 1279 29835
rect 999 29767 1313 29801
rect 999 29733 1051 29767
rect 1085 29733 1127 29767
rect 1161 29733 1203 29767
rect 1237 29733 1279 29767
rect 999 29699 1313 29733
rect 999 29665 1051 29699
rect 1085 29665 1127 29699
rect 1161 29665 1203 29699
rect 1237 29665 1279 29699
rect 999 29631 1313 29665
rect 999 29597 1051 29631
rect 1085 29597 1127 29631
rect 1161 29597 1203 29631
rect 1237 29597 1279 29631
rect 999 29563 1313 29597
rect 999 29529 1051 29563
rect 1085 29529 1127 29563
rect 1161 29529 1203 29563
rect 1237 29529 1279 29563
rect 999 29495 1313 29529
rect 999 29461 1051 29495
rect 1085 29461 1127 29495
rect 1161 29461 1203 29495
rect 1237 29461 1279 29495
rect 999 29427 1313 29461
rect 999 29393 1051 29427
rect 1085 29393 1127 29427
rect 1161 29393 1203 29427
rect 1237 29393 1279 29427
rect 999 29359 1313 29393
rect 999 29325 1051 29359
rect 1085 29325 1127 29359
rect 1161 29325 1203 29359
rect 1237 29325 1279 29359
rect 999 29291 1313 29325
rect 999 29257 1051 29291
rect 1085 29257 1127 29291
rect 1161 29257 1203 29291
rect 1237 29257 1279 29291
rect 999 29223 1313 29257
rect 999 29189 1051 29223
rect 1085 29189 1127 29223
rect 1161 29189 1203 29223
rect 1237 29189 1279 29223
rect 999 29155 1313 29189
rect 999 29121 1051 29155
rect 1085 29121 1127 29155
rect 1161 29121 1203 29155
rect 1237 29121 1279 29155
rect 999 29086 1313 29121
rect 999 29052 1051 29086
rect 1085 29052 1127 29086
rect 1161 29052 1203 29086
rect 1237 29052 1279 29086
rect 999 29017 1313 29052
rect 999 28983 1051 29017
rect 1085 28983 1127 29017
rect 1161 28983 1203 29017
rect 1237 28983 1279 29017
rect 999 28948 1313 28983
rect 999 28914 1051 28948
rect 1085 28914 1127 28948
rect 1161 28914 1203 28948
rect 1237 28914 1279 28948
rect 999 28879 1313 28914
rect 999 28845 1051 28879
rect 1085 28845 1127 28879
rect 1161 28845 1203 28879
rect 1237 28845 1279 28879
rect 999 28810 1313 28845
rect 999 28776 1051 28810
rect 1085 28776 1127 28810
rect 1161 28776 1203 28810
rect 1237 28776 1279 28810
rect 999 28741 1313 28776
rect 999 28707 1051 28741
rect 1085 28707 1127 28741
rect 1161 28707 1203 28741
rect 1237 28707 1279 28741
rect 999 28672 1313 28707
rect 999 28638 1051 28672
rect 1085 28638 1127 28672
rect 1161 28638 1203 28672
rect 1237 28638 1279 28672
rect 999 28603 1313 28638
rect 999 28569 1051 28603
rect 1085 28569 1127 28603
rect 1161 28569 1203 28603
rect 1237 28569 1279 28603
rect 999 28534 1313 28569
rect 999 28500 1051 28534
rect 1085 28500 1127 28534
rect 1161 28500 1203 28534
rect 1237 28500 1279 28534
rect 999 28465 1313 28500
rect 999 28431 1051 28465
rect 1085 28431 1127 28465
rect 1161 28431 1203 28465
rect 1237 28431 1279 28465
rect 999 28396 1313 28431
rect 999 28362 1051 28396
rect 1085 28362 1127 28396
rect 1161 28362 1203 28396
rect 1237 28362 1279 28396
rect 999 28327 1313 28362
rect 999 28293 1051 28327
rect 1085 28293 1127 28327
rect 1161 28293 1203 28327
rect 1237 28293 1279 28327
rect 999 28258 1313 28293
rect 999 28224 1051 28258
rect 1085 28224 1127 28258
rect 1161 28224 1203 28258
rect 1237 28224 1279 28258
rect 999 28189 1313 28224
rect 999 28155 1051 28189
rect 1085 28155 1127 28189
rect 1161 28155 1203 28189
rect 1237 28155 1279 28189
rect 999 28120 1313 28155
rect 999 28086 1051 28120
rect 1085 28086 1127 28120
rect 1161 28086 1203 28120
rect 1237 28086 1279 28120
rect 999 28051 1313 28086
rect 999 28017 1051 28051
rect 1085 28017 1127 28051
rect 1161 28017 1203 28051
rect 1237 28017 1279 28051
rect 999 27982 1313 28017
rect 999 27948 1051 27982
rect 1085 27948 1127 27982
rect 1161 27948 1203 27982
rect 1237 27948 1279 27982
rect 999 27913 1313 27948
rect 999 27879 1051 27913
rect 1085 27879 1127 27913
rect 1161 27879 1203 27913
rect 1237 27879 1279 27913
rect 999 27844 1313 27879
rect 999 27810 1051 27844
rect 1085 27810 1127 27844
rect 1161 27810 1203 27844
rect 1237 27810 1279 27844
rect 999 27775 1313 27810
rect 999 27741 1051 27775
rect 1085 27741 1127 27775
rect 1161 27741 1203 27775
rect 1237 27741 1279 27775
rect 999 27706 1313 27741
rect 999 27672 1051 27706
rect 1085 27672 1127 27706
rect 1161 27672 1203 27706
rect 1237 27672 1279 27706
rect 999 27637 1313 27672
rect 999 27603 1051 27637
rect 1085 27603 1127 27637
rect 1161 27603 1203 27637
rect 1237 27603 1279 27637
rect 999 27568 1313 27603
rect 999 27534 1051 27568
rect 1085 27534 1127 27568
rect 1161 27534 1203 27568
rect 1237 27534 1279 27568
rect 999 27499 1313 27534
rect 999 27465 1051 27499
rect 1085 27465 1127 27499
rect 1161 27465 1203 27499
rect 1237 27465 1279 27499
rect 999 27430 1313 27465
rect 999 27396 1051 27430
rect 1085 27396 1127 27430
rect 1161 27396 1203 27430
rect 1237 27396 1279 27430
rect 999 27361 1313 27396
rect 999 27327 1051 27361
rect 1085 27327 1127 27361
rect 1161 27327 1203 27361
rect 1237 27327 1279 27361
rect 999 27292 1313 27327
rect 999 27258 1051 27292
rect 1085 27258 1127 27292
rect 1161 27258 1203 27292
rect 1237 27258 1279 27292
rect 999 27223 1313 27258
rect 999 27189 1051 27223
rect 1085 27189 1127 27223
rect 1161 27189 1203 27223
rect 1237 27189 1279 27223
rect 999 27103 1313 27189
rect 18021 31675 18442 31709
rect 18021 31672 18025 31675
rect 18021 31638 18022 31672
rect 18059 31641 18101 31675
rect 18135 31672 18177 31675
rect 18211 31672 18253 31675
rect 18287 31672 18329 31675
rect 18142 31641 18177 31672
rect 18228 31641 18253 31672
rect 18314 31641 18329 31672
rect 18363 31672 18405 31675
rect 18363 31641 18366 31672
rect 18056 31638 18108 31641
rect 18142 31638 18194 31641
rect 18228 31638 18280 31641
rect 18314 31638 18366 31641
rect 18400 31641 18405 31672
rect 18439 31641 18442 31675
rect 18400 31638 18442 31641
rect 18021 31607 18442 31638
rect 18021 31600 18025 31607
rect 18021 31566 18022 31600
rect 18059 31573 18101 31607
rect 18135 31600 18177 31607
rect 18211 31600 18253 31607
rect 18287 31600 18329 31607
rect 18142 31573 18177 31600
rect 18228 31573 18253 31600
rect 18314 31573 18329 31600
rect 18363 31600 18405 31607
rect 18363 31573 18366 31600
rect 18056 31566 18108 31573
rect 18142 31566 18194 31573
rect 18228 31566 18280 31573
rect 18314 31566 18366 31573
rect 18400 31573 18405 31600
rect 18439 31573 18442 31607
rect 18400 31566 18442 31573
rect 18021 31539 18442 31566
rect 18021 31528 18025 31539
rect 18021 31494 18022 31528
rect 18059 31505 18101 31539
rect 18135 31528 18177 31539
rect 18211 31528 18253 31539
rect 18287 31528 18329 31539
rect 18142 31505 18177 31528
rect 18228 31505 18253 31528
rect 18314 31505 18329 31528
rect 18363 31528 18405 31539
rect 18363 31505 18366 31528
rect 18056 31494 18108 31505
rect 18142 31494 18194 31505
rect 18228 31494 18280 31505
rect 18314 31494 18366 31505
rect 18400 31505 18405 31528
rect 18439 31505 18442 31539
rect 18400 31494 18442 31505
rect 18021 31471 18442 31494
rect 18021 31456 18025 31471
rect 18021 31422 18022 31456
rect 18059 31437 18101 31471
rect 18135 31456 18177 31471
rect 18211 31456 18253 31471
rect 18287 31456 18329 31471
rect 18142 31437 18177 31456
rect 18228 31437 18253 31456
rect 18314 31437 18329 31456
rect 18363 31456 18405 31471
rect 18363 31437 18366 31456
rect 18056 31422 18108 31437
rect 18142 31422 18194 31437
rect 18228 31422 18280 31437
rect 18314 31422 18366 31437
rect 18400 31437 18405 31456
rect 18439 31437 18442 31471
rect 18400 31422 18442 31437
rect 18021 31403 18442 31422
rect 18021 31384 18025 31403
rect 18021 31350 18022 31384
rect 18059 31369 18101 31403
rect 18135 31384 18177 31403
rect 18211 31384 18253 31403
rect 18287 31384 18329 31403
rect 18142 31369 18177 31384
rect 18228 31369 18253 31384
rect 18314 31369 18329 31384
rect 18363 31384 18405 31403
rect 18363 31369 18366 31384
rect 18056 31350 18108 31369
rect 18142 31350 18194 31369
rect 18228 31350 18280 31369
rect 18314 31350 18366 31369
rect 18400 31369 18405 31384
rect 18439 31369 18442 31403
rect 18400 31350 18442 31369
rect 18021 31335 18442 31350
rect 18021 31312 18025 31335
rect 18021 31278 18022 31312
rect 18059 31301 18101 31335
rect 18135 31312 18177 31335
rect 18211 31312 18253 31335
rect 18287 31312 18329 31335
rect 18142 31301 18177 31312
rect 18228 31301 18253 31312
rect 18314 31301 18329 31312
rect 18363 31312 18405 31335
rect 18363 31301 18366 31312
rect 18056 31278 18108 31301
rect 18142 31278 18194 31301
rect 18228 31278 18280 31301
rect 18314 31278 18366 31301
rect 18400 31301 18405 31312
rect 18439 31301 18442 31335
rect 18400 31278 18442 31301
rect 18021 31267 18442 31278
rect 18021 31240 18025 31267
rect 18021 31206 18022 31240
rect 18059 31233 18101 31267
rect 18135 31240 18177 31267
rect 18211 31240 18253 31267
rect 18287 31240 18329 31267
rect 18142 31233 18177 31240
rect 18228 31233 18253 31240
rect 18314 31233 18329 31240
rect 18363 31240 18405 31267
rect 18363 31233 18366 31240
rect 18056 31206 18108 31233
rect 18142 31206 18194 31233
rect 18228 31206 18280 31233
rect 18314 31206 18366 31233
rect 18400 31233 18405 31240
rect 18439 31233 18442 31267
rect 18400 31206 18442 31233
rect 18021 31199 18442 31206
rect 18021 31168 18025 31199
rect 18021 31134 18022 31168
rect 18059 31165 18101 31199
rect 18135 31168 18177 31199
rect 18211 31168 18253 31199
rect 18287 31168 18329 31199
rect 18142 31165 18177 31168
rect 18228 31165 18253 31168
rect 18314 31165 18329 31168
rect 18363 31168 18405 31199
rect 18363 31165 18366 31168
rect 18056 31134 18108 31165
rect 18142 31134 18194 31165
rect 18228 31134 18280 31165
rect 18314 31134 18366 31165
rect 18400 31165 18405 31168
rect 18439 31165 18442 31199
rect 18400 31134 18442 31165
rect 18021 31131 18442 31134
rect 18021 31097 18025 31131
rect 18059 31097 18101 31131
rect 18135 31097 18177 31131
rect 18211 31097 18253 31131
rect 18287 31097 18329 31131
rect 18363 31097 18405 31131
rect 18439 31097 18442 31131
rect 18021 31096 18442 31097
rect 18021 31062 18022 31096
rect 18056 31063 18108 31096
rect 18142 31063 18194 31096
rect 18228 31063 18280 31096
rect 18314 31063 18366 31096
rect 18021 31029 18025 31062
rect 18059 31029 18101 31063
rect 18142 31062 18177 31063
rect 18228 31062 18253 31063
rect 18314 31062 18329 31063
rect 18135 31029 18177 31062
rect 18211 31029 18253 31062
rect 18287 31029 18329 31062
rect 18363 31062 18366 31063
rect 18400 31063 18442 31096
rect 18400 31062 18405 31063
rect 18363 31029 18405 31062
rect 18439 31029 18442 31063
rect 18021 31024 18442 31029
rect 18021 30990 18022 31024
rect 18056 30995 18108 31024
rect 18142 30995 18194 31024
rect 18228 30995 18280 31024
rect 18314 30995 18366 31024
rect 18021 30961 18025 30990
rect 18059 30961 18101 30995
rect 18142 30990 18177 30995
rect 18228 30990 18253 30995
rect 18314 30990 18329 30995
rect 18135 30961 18177 30990
rect 18211 30961 18253 30990
rect 18287 30961 18329 30990
rect 18363 30990 18366 30995
rect 18400 30995 18442 31024
rect 18400 30990 18405 30995
rect 18363 30961 18405 30990
rect 18439 30961 18442 30995
rect 18021 30952 18442 30961
rect 18021 30918 18022 30952
rect 18056 30927 18108 30952
rect 18142 30927 18194 30952
rect 18228 30927 18280 30952
rect 18314 30927 18366 30952
rect 18021 30893 18025 30918
rect 18059 30893 18101 30927
rect 18142 30918 18177 30927
rect 18228 30918 18253 30927
rect 18314 30918 18329 30927
rect 18135 30893 18177 30918
rect 18211 30893 18253 30918
rect 18287 30893 18329 30918
rect 18363 30918 18366 30927
rect 18400 30927 18442 30952
rect 18400 30918 18405 30927
rect 18363 30893 18405 30918
rect 18439 30893 18442 30927
rect 18021 30880 18442 30893
rect 18021 30846 18022 30880
rect 18056 30859 18108 30880
rect 18142 30859 18194 30880
rect 18228 30859 18280 30880
rect 18314 30859 18366 30880
rect 18021 30825 18025 30846
rect 18059 30825 18101 30859
rect 18142 30846 18177 30859
rect 18228 30846 18253 30859
rect 18314 30846 18329 30859
rect 18135 30825 18177 30846
rect 18211 30825 18253 30846
rect 18287 30825 18329 30846
rect 18363 30846 18366 30859
rect 18400 30859 18442 30880
rect 18400 30846 18405 30859
rect 18363 30825 18405 30846
rect 18439 30825 18442 30859
rect 18021 30808 18442 30825
rect 18021 30774 18022 30808
rect 18056 30791 18108 30808
rect 18142 30791 18194 30808
rect 18228 30791 18280 30808
rect 18314 30791 18366 30808
rect 18021 30757 18025 30774
rect 18059 30757 18101 30791
rect 18142 30774 18177 30791
rect 18228 30774 18253 30791
rect 18314 30774 18329 30791
rect 18135 30757 18177 30774
rect 18211 30757 18253 30774
rect 18287 30757 18329 30774
rect 18363 30774 18366 30791
rect 18400 30791 18442 30808
rect 18400 30774 18405 30791
rect 18363 30757 18405 30774
rect 18439 30757 18442 30791
rect 18021 30736 18442 30757
rect 18021 30702 18022 30736
rect 18056 30723 18108 30736
rect 18142 30723 18194 30736
rect 18228 30723 18280 30736
rect 18314 30723 18366 30736
rect 18021 30689 18025 30702
rect 18059 30689 18101 30723
rect 18142 30702 18177 30723
rect 18228 30702 18253 30723
rect 18314 30702 18329 30723
rect 18135 30689 18177 30702
rect 18211 30689 18253 30702
rect 18287 30689 18329 30702
rect 18363 30702 18366 30723
rect 18400 30723 18442 30736
rect 18400 30702 18405 30723
rect 18363 30689 18405 30702
rect 18439 30705 18442 30723
rect 22823 33312 22829 33335
rect 22863 33312 22911 33335
rect 22945 33312 22993 33335
rect 23027 33312 23075 33335
rect 23109 33312 23157 33335
rect 23191 33312 23239 33335
rect 23273 33312 23635 33335
rect 22823 33301 23635 33312
rect 22823 33267 22827 33301
rect 22861 33273 22897 33301
rect 22931 33273 22967 33301
rect 23001 33273 23037 33301
rect 22863 33267 22897 33273
rect 22945 33267 22967 33273
rect 23027 33267 23037 33273
rect 23071 33273 23107 33301
rect 23141 33273 23177 33301
rect 23211 33273 23247 33301
rect 23071 33267 23075 33273
rect 23141 33267 23157 33273
rect 23211 33267 23239 33273
rect 23281 33267 23317 33301
rect 23351 33267 23387 33301
rect 23421 33267 23457 33301
rect 23491 33267 23527 33301
rect 23561 33267 23597 33301
rect 23631 33267 23635 33301
rect 22823 33239 22829 33267
rect 22863 33239 22911 33267
rect 22945 33239 22993 33267
rect 23027 33239 23075 33267
rect 23109 33239 23157 33267
rect 23191 33239 23239 33267
rect 23273 33239 23635 33267
rect 22823 33233 23635 33239
rect 22823 33199 22827 33233
rect 22861 33200 22897 33233
rect 22931 33200 22967 33233
rect 23001 33200 23037 33233
rect 22863 33199 22897 33200
rect 22945 33199 22967 33200
rect 23027 33199 23037 33200
rect 23071 33200 23107 33233
rect 23141 33200 23177 33233
rect 23211 33200 23247 33233
rect 23071 33199 23075 33200
rect 23141 33199 23157 33200
rect 23211 33199 23239 33200
rect 23281 33199 23317 33233
rect 23351 33199 23387 33233
rect 23421 33199 23457 33233
rect 23491 33199 23527 33233
rect 23561 33199 23597 33233
rect 23631 33199 23635 33233
rect 22823 33166 22829 33199
rect 22863 33166 22911 33199
rect 22945 33166 22993 33199
rect 23027 33166 23075 33199
rect 23109 33166 23157 33199
rect 23191 33166 23239 33199
rect 23273 33166 23635 33199
rect 22823 33165 23635 33166
rect 22823 33131 22827 33165
rect 22861 33131 22897 33165
rect 22931 33131 22967 33165
rect 23001 33131 23037 33165
rect 23071 33131 23107 33165
rect 23141 33131 23177 33165
rect 23211 33131 23247 33165
rect 23281 33131 23317 33165
rect 23351 33131 23387 33165
rect 23421 33131 23457 33165
rect 23491 33131 23527 33165
rect 23561 33131 23597 33165
rect 23631 33131 23635 33165
rect 22823 33127 23635 33131
rect 22823 33097 22829 33127
rect 22863 33097 22911 33127
rect 22945 33097 22993 33127
rect 23027 33097 23075 33127
rect 23109 33097 23157 33127
rect 23191 33097 23239 33127
rect 23273 33097 23635 33127
rect 22823 33063 22827 33097
rect 22863 33093 22897 33097
rect 22945 33093 22967 33097
rect 23027 33093 23037 33097
rect 22861 33063 22897 33093
rect 22931 33063 22967 33093
rect 23001 33063 23037 33093
rect 23071 33093 23075 33097
rect 23141 33093 23157 33097
rect 23211 33093 23239 33097
rect 23071 33063 23107 33093
rect 23141 33063 23177 33093
rect 23211 33063 23247 33093
rect 23281 33063 23317 33097
rect 23351 33063 23387 33097
rect 23421 33063 23457 33097
rect 23491 33063 23527 33097
rect 23561 33063 23597 33097
rect 23631 33063 23635 33097
rect 22823 33054 23635 33063
rect 22823 33029 22829 33054
rect 22863 33029 22911 33054
rect 22945 33029 22993 33054
rect 23027 33029 23075 33054
rect 23109 33029 23157 33054
rect 23191 33029 23239 33054
rect 23273 33029 23635 33054
rect 22823 32995 22827 33029
rect 22863 33020 22897 33029
rect 22945 33020 22967 33029
rect 23027 33020 23037 33029
rect 22861 32995 22897 33020
rect 22931 32995 22967 33020
rect 23001 32995 23037 33020
rect 23071 33020 23075 33029
rect 23141 33020 23157 33029
rect 23211 33020 23239 33029
rect 23071 32995 23107 33020
rect 23141 32995 23177 33020
rect 23211 32995 23247 33020
rect 23281 32995 23317 33029
rect 23351 32995 23387 33029
rect 23421 32995 23457 33029
rect 23491 32995 23527 33029
rect 23561 32995 23597 33029
rect 23631 32995 23635 33029
rect 22823 32981 23635 32995
rect 22823 32961 22829 32981
rect 22863 32961 22911 32981
rect 22945 32961 22993 32981
rect 23027 32961 23075 32981
rect 23109 32961 23157 32981
rect 23191 32961 23239 32981
rect 23273 32961 23635 32981
rect 22823 32927 22827 32961
rect 22863 32947 22897 32961
rect 22945 32947 22967 32961
rect 23027 32947 23037 32961
rect 22861 32927 22897 32947
rect 22931 32927 22967 32947
rect 23001 32927 23037 32947
rect 23071 32947 23075 32961
rect 23141 32947 23157 32961
rect 23211 32947 23239 32961
rect 23071 32927 23107 32947
rect 23141 32927 23177 32947
rect 23211 32927 23247 32947
rect 23281 32927 23317 32961
rect 23351 32927 23387 32961
rect 23421 32927 23457 32961
rect 23491 32927 23527 32961
rect 23561 32927 23597 32961
rect 23631 32927 23635 32961
rect 22823 32908 23635 32927
rect 22823 32893 22829 32908
rect 22863 32893 22911 32908
rect 22945 32893 22993 32908
rect 23027 32893 23075 32908
rect 23109 32893 23157 32908
rect 23191 32893 23239 32908
rect 23273 32893 23635 32908
rect 22823 32859 22827 32893
rect 22863 32874 22897 32893
rect 22945 32874 22967 32893
rect 23027 32874 23037 32893
rect 22861 32859 22897 32874
rect 22931 32859 22967 32874
rect 23001 32859 23037 32874
rect 23071 32874 23075 32893
rect 23141 32874 23157 32893
rect 23211 32874 23239 32893
rect 23071 32859 23107 32874
rect 23141 32859 23177 32874
rect 23211 32859 23247 32874
rect 23281 32859 23317 32893
rect 23351 32859 23387 32893
rect 23421 32859 23457 32893
rect 23491 32859 23527 32893
rect 23561 32859 23597 32893
rect 23631 32859 23635 32893
rect 22823 32835 23635 32859
rect 22823 32825 22829 32835
rect 22863 32825 22911 32835
rect 22945 32825 22993 32835
rect 23027 32825 23075 32835
rect 23109 32825 23157 32835
rect 23191 32825 23239 32835
rect 23273 32825 23635 32835
rect 22823 32791 22827 32825
rect 22863 32801 22897 32825
rect 22945 32801 22967 32825
rect 23027 32801 23037 32825
rect 22861 32791 22897 32801
rect 22931 32791 22967 32801
rect 23001 32791 23037 32801
rect 23071 32801 23075 32825
rect 23141 32801 23157 32825
rect 23211 32801 23239 32825
rect 23071 32791 23107 32801
rect 23141 32791 23177 32801
rect 23211 32791 23247 32801
rect 23281 32791 23317 32825
rect 23351 32791 23387 32825
rect 23421 32791 23457 32825
rect 23491 32791 23527 32825
rect 23561 32791 23597 32825
rect 23631 32791 23635 32825
rect 22823 32762 23635 32791
rect 22823 32757 22829 32762
rect 22863 32757 22911 32762
rect 22945 32757 22993 32762
rect 23027 32757 23075 32762
rect 23109 32757 23157 32762
rect 23191 32757 23239 32762
rect 23273 32757 23635 32762
rect 22823 32723 22827 32757
rect 22863 32728 22897 32757
rect 22945 32728 22967 32757
rect 23027 32728 23037 32757
rect 22861 32723 22897 32728
rect 22931 32723 22967 32728
rect 23001 32723 23037 32728
rect 23071 32728 23075 32757
rect 23141 32728 23157 32757
rect 23211 32728 23239 32757
rect 23071 32723 23107 32728
rect 23141 32723 23177 32728
rect 23211 32723 23247 32728
rect 23281 32723 23317 32757
rect 23351 32723 23387 32757
rect 23421 32723 23457 32757
rect 23491 32723 23527 32757
rect 23561 32723 23597 32757
rect 23631 32723 23635 32757
rect 22823 32689 23635 32723
rect 22823 32655 22827 32689
rect 22863 32655 22897 32689
rect 22945 32655 22967 32689
rect 23027 32655 23037 32689
rect 23071 32655 23075 32689
rect 23141 32655 23157 32689
rect 23211 32655 23239 32689
rect 23281 32655 23317 32689
rect 23351 32655 23387 32689
rect 23421 32655 23457 32689
rect 23491 32655 23527 32689
rect 23561 32655 23597 32689
rect 23631 32655 23635 32689
rect 22823 32621 23635 32655
rect 22823 32587 22827 32621
rect 22861 32616 22897 32621
rect 22931 32616 22967 32621
rect 23001 32616 23037 32621
rect 22863 32587 22897 32616
rect 22945 32587 22967 32616
rect 23027 32587 23037 32616
rect 23071 32616 23107 32621
rect 23141 32616 23177 32621
rect 23211 32616 23247 32621
rect 23071 32587 23075 32616
rect 23141 32587 23157 32616
rect 23211 32587 23239 32616
rect 23281 32587 23317 32621
rect 23351 32587 23387 32621
rect 23421 32587 23457 32621
rect 23491 32587 23527 32621
rect 23561 32587 23597 32621
rect 23631 32587 23635 32621
rect 22823 32582 22829 32587
rect 22863 32582 22911 32587
rect 22945 32582 22993 32587
rect 23027 32582 23075 32587
rect 23109 32582 23157 32587
rect 23191 32582 23239 32587
rect 23273 32582 23635 32587
rect 22823 32553 23635 32582
rect 22823 32519 22827 32553
rect 22861 32543 22897 32553
rect 22931 32543 22967 32553
rect 23001 32543 23037 32553
rect 22863 32519 22897 32543
rect 22945 32519 22967 32543
rect 23027 32519 23037 32543
rect 23071 32543 23107 32553
rect 23141 32543 23177 32553
rect 23211 32543 23247 32553
rect 23071 32519 23075 32543
rect 23141 32519 23157 32543
rect 23211 32519 23239 32543
rect 23281 32519 23317 32553
rect 23351 32519 23387 32553
rect 23421 32519 23457 32553
rect 23491 32519 23527 32553
rect 23561 32519 23597 32553
rect 23631 32519 23635 32553
rect 22823 32509 22829 32519
rect 22863 32509 22911 32519
rect 22945 32509 22993 32519
rect 23027 32509 23075 32519
rect 23109 32509 23157 32519
rect 23191 32509 23239 32519
rect 23273 32509 23635 32519
rect 22823 32485 23635 32509
rect 22823 32451 22827 32485
rect 22861 32470 22897 32485
rect 22931 32470 22967 32485
rect 23001 32470 23037 32485
rect 22863 32451 22897 32470
rect 22945 32451 22967 32470
rect 23027 32451 23037 32470
rect 23071 32470 23107 32485
rect 23141 32470 23177 32485
rect 23211 32470 23247 32485
rect 23071 32451 23075 32470
rect 23141 32451 23157 32470
rect 23211 32451 23239 32470
rect 23281 32451 23317 32485
rect 23351 32451 23387 32485
rect 23421 32451 23457 32485
rect 23491 32451 23527 32485
rect 23561 32451 23597 32485
rect 23631 32451 23635 32485
rect 22823 32436 22829 32451
rect 22863 32436 22911 32451
rect 22945 32436 22993 32451
rect 23027 32436 23075 32451
rect 23109 32436 23157 32451
rect 23191 32436 23239 32451
rect 23273 32436 23635 32451
rect 22823 32417 23635 32436
rect 22823 32383 22827 32417
rect 22861 32397 22897 32417
rect 22931 32397 22967 32417
rect 23001 32397 23037 32417
rect 22863 32383 22897 32397
rect 22945 32383 22967 32397
rect 23027 32383 23037 32397
rect 23071 32397 23107 32417
rect 23141 32397 23177 32417
rect 23211 32397 23247 32417
rect 23071 32383 23075 32397
rect 23141 32383 23157 32397
rect 23211 32383 23239 32397
rect 23281 32383 23317 32417
rect 23351 32383 23387 32417
rect 23421 32383 23457 32417
rect 23491 32383 23527 32417
rect 23561 32383 23597 32417
rect 23631 32383 23635 32417
rect 22823 32363 22829 32383
rect 22863 32363 22911 32383
rect 22945 32363 22993 32383
rect 23027 32363 23075 32383
rect 23109 32363 23157 32383
rect 23191 32363 23239 32383
rect 23273 32363 23635 32383
rect 22823 32349 23635 32363
rect 22823 32315 22827 32349
rect 22861 32324 22897 32349
rect 22931 32324 22967 32349
rect 23001 32324 23037 32349
rect 22863 32315 22897 32324
rect 22945 32315 22967 32324
rect 23027 32315 23037 32324
rect 23071 32324 23107 32349
rect 23141 32324 23177 32349
rect 23211 32324 23247 32349
rect 23071 32315 23075 32324
rect 23141 32315 23157 32324
rect 23211 32315 23239 32324
rect 23281 32315 23317 32349
rect 23351 32315 23387 32349
rect 23421 32315 23457 32349
rect 23491 32315 23527 32349
rect 23561 32315 23597 32349
rect 23631 32315 23635 32349
rect 22823 32290 22829 32315
rect 22863 32290 22911 32315
rect 22945 32290 22993 32315
rect 23027 32290 23075 32315
rect 23109 32290 23157 32315
rect 23191 32290 23239 32315
rect 23273 32290 23635 32315
rect 22823 32281 23635 32290
rect 22823 32247 22827 32281
rect 22861 32251 22897 32281
rect 22931 32251 22967 32281
rect 23001 32251 23037 32281
rect 22863 32247 22897 32251
rect 22945 32247 22967 32251
rect 23027 32247 23037 32251
rect 23071 32251 23107 32281
rect 23141 32251 23177 32281
rect 23211 32251 23247 32281
rect 23071 32247 23075 32251
rect 23141 32247 23157 32251
rect 23211 32247 23239 32251
rect 23281 32247 23317 32281
rect 23351 32247 23387 32281
rect 23421 32247 23457 32281
rect 23491 32247 23527 32281
rect 23561 32247 23597 32281
rect 23631 32247 23635 32281
rect 22823 32217 22829 32247
rect 22863 32217 22911 32247
rect 22945 32217 22993 32247
rect 23027 32217 23075 32247
rect 23109 32217 23157 32247
rect 23191 32217 23239 32247
rect 23273 32217 23635 32247
rect 22823 32213 23635 32217
rect 22823 32179 22827 32213
rect 22861 32179 22897 32213
rect 22931 32179 22967 32213
rect 23001 32179 23037 32213
rect 23071 32179 23107 32213
rect 23141 32179 23177 32213
rect 23211 32179 23247 32213
rect 23281 32179 23317 32213
rect 23351 32179 23387 32213
rect 23421 32179 23457 32213
rect 23491 32179 23527 32213
rect 23561 32179 23597 32213
rect 23631 32179 23635 32213
rect 22823 32178 23635 32179
rect 22823 32145 22829 32178
rect 22863 32145 22911 32178
rect 22945 32145 22993 32178
rect 23027 32145 23075 32178
rect 23109 32145 23157 32178
rect 23191 32145 23239 32178
rect 23273 32145 23635 32178
rect 22823 32111 22827 32145
rect 22863 32144 22897 32145
rect 22945 32144 22967 32145
rect 23027 32144 23037 32145
rect 22861 32111 22897 32144
rect 22931 32111 22967 32144
rect 23001 32111 23037 32144
rect 23071 32144 23075 32145
rect 23141 32144 23157 32145
rect 23211 32144 23239 32145
rect 23071 32111 23107 32144
rect 23141 32111 23177 32144
rect 23211 32111 23247 32144
rect 23281 32111 23317 32145
rect 23351 32111 23387 32145
rect 23421 32111 23457 32145
rect 23491 32111 23527 32145
rect 23561 32111 23597 32145
rect 23631 32111 23635 32145
rect 22823 32105 23635 32111
rect 22823 32077 22829 32105
rect 22863 32077 22911 32105
rect 22945 32077 22993 32105
rect 23027 32077 23075 32105
rect 23109 32077 23157 32105
rect 23191 32077 23239 32105
rect 23273 32077 23635 32105
rect 22823 32043 22827 32077
rect 22863 32071 22897 32077
rect 22945 32071 22967 32077
rect 23027 32071 23037 32077
rect 22861 32043 22897 32071
rect 22931 32043 22967 32071
rect 23001 32043 23037 32071
rect 23071 32071 23075 32077
rect 23141 32071 23157 32077
rect 23211 32071 23239 32077
rect 23071 32043 23107 32071
rect 23141 32043 23177 32071
rect 23211 32043 23247 32071
rect 23281 32043 23317 32077
rect 23351 32043 23387 32077
rect 23421 32043 23457 32077
rect 23491 32043 23527 32077
rect 23561 32043 23597 32077
rect 23631 32043 23635 32077
rect 22823 32032 23635 32043
rect 22823 32009 22829 32032
rect 22863 32009 22911 32032
rect 22945 32009 22993 32032
rect 23027 32009 23075 32032
rect 23109 32009 23157 32032
rect 23191 32009 23239 32032
rect 23273 32009 23635 32032
rect 22823 31975 22827 32009
rect 22863 31998 22897 32009
rect 22945 31998 22967 32009
rect 23027 31998 23037 32009
rect 22861 31975 22897 31998
rect 22931 31975 22967 31998
rect 23001 31975 23037 31998
rect 23071 31998 23075 32009
rect 23141 31998 23157 32009
rect 23211 31998 23239 32009
rect 23071 31975 23107 31998
rect 23141 31975 23177 31998
rect 23211 31975 23247 31998
rect 23281 31975 23317 32009
rect 23351 31975 23387 32009
rect 23421 31975 23457 32009
rect 23491 31975 23527 32009
rect 23561 31975 23597 32009
rect 23631 31975 23635 32009
rect 22823 31959 23635 31975
rect 22823 31941 22829 31959
rect 22863 31941 22911 31959
rect 22945 31941 22993 31959
rect 23027 31941 23075 31959
rect 23109 31941 23157 31959
rect 23191 31941 23239 31959
rect 23273 31941 23635 31959
rect 22823 31907 22827 31941
rect 22863 31925 22897 31941
rect 22945 31925 22967 31941
rect 23027 31925 23037 31941
rect 22861 31907 22897 31925
rect 22931 31907 22967 31925
rect 23001 31907 23037 31925
rect 23071 31925 23075 31941
rect 23141 31925 23157 31941
rect 23211 31925 23239 31941
rect 23071 31907 23107 31925
rect 23141 31907 23177 31925
rect 23211 31907 23247 31925
rect 23281 31907 23317 31941
rect 23351 31907 23387 31941
rect 23421 31907 23457 31941
rect 23491 31907 23527 31941
rect 23561 31907 23597 31941
rect 23631 31907 23635 31941
rect 22823 31886 23635 31907
rect 22823 31873 22829 31886
rect 22863 31873 22911 31886
rect 22945 31873 22993 31886
rect 23027 31873 23075 31886
rect 23109 31873 23157 31886
rect 23191 31873 23239 31886
rect 23273 31873 23635 31886
rect 22823 31839 22827 31873
rect 22863 31852 22897 31873
rect 22945 31852 22967 31873
rect 23027 31852 23037 31873
rect 22861 31839 22897 31852
rect 22931 31839 22967 31852
rect 23001 31839 23037 31852
rect 23071 31852 23075 31873
rect 23141 31852 23157 31873
rect 23211 31852 23239 31873
rect 23071 31839 23107 31852
rect 23141 31839 23177 31852
rect 23211 31839 23247 31852
rect 23281 31839 23317 31873
rect 23351 31839 23387 31873
rect 23421 31839 23457 31873
rect 23491 31839 23527 31873
rect 23561 31839 23597 31873
rect 23631 31839 23635 31873
rect 22823 31813 23635 31839
rect 22823 31805 22829 31813
rect 22863 31805 22911 31813
rect 22945 31805 22993 31813
rect 23027 31805 23075 31813
rect 23109 31805 23157 31813
rect 23191 31805 23239 31813
rect 23273 31805 23635 31813
rect 22823 31771 22827 31805
rect 22863 31779 22897 31805
rect 22945 31779 22967 31805
rect 23027 31779 23037 31805
rect 22861 31771 22897 31779
rect 22931 31771 22967 31779
rect 23001 31771 23037 31779
rect 23071 31779 23075 31805
rect 23141 31779 23157 31805
rect 23211 31779 23239 31805
rect 23071 31771 23107 31779
rect 23141 31771 23177 31779
rect 23211 31771 23247 31779
rect 23281 31771 23317 31805
rect 23351 31771 23387 31805
rect 23421 31771 23457 31805
rect 23491 31771 23527 31805
rect 23561 31771 23597 31805
rect 23631 31771 23635 31805
rect 22823 31740 23635 31771
rect 22823 31737 22829 31740
rect 22863 31737 22911 31740
rect 22945 31737 22993 31740
rect 23027 31737 23075 31740
rect 23109 31737 23157 31740
rect 23191 31737 23239 31740
rect 23273 31737 23635 31740
rect 22823 31703 22827 31737
rect 22863 31706 22897 31737
rect 22945 31706 22967 31737
rect 23027 31706 23037 31737
rect 22861 31703 22897 31706
rect 22931 31703 22967 31706
rect 23001 31703 23037 31706
rect 23071 31706 23075 31737
rect 23141 31706 23157 31737
rect 23211 31706 23239 31737
rect 23071 31703 23107 31706
rect 23141 31703 23177 31706
rect 23211 31703 23247 31706
rect 23281 31703 23317 31737
rect 23351 31703 23387 31737
rect 23421 31703 23457 31737
rect 23491 31703 23527 31737
rect 23561 31703 23597 31737
rect 23631 31703 23635 31737
rect 22823 31669 23635 31703
rect 22823 31635 22827 31669
rect 22861 31642 22897 31669
rect 22864 31635 22897 31642
rect 22931 31642 22967 31669
rect 22931 31635 22932 31642
rect 22823 31608 22830 31635
rect 22864 31608 22932 31635
rect 22966 31635 22967 31642
rect 23001 31642 23037 31669
rect 23001 31635 23034 31642
rect 23071 31635 23107 31669
rect 23141 31635 23177 31669
rect 23211 31635 23247 31669
rect 23281 31635 23317 31669
rect 23351 31635 23387 31669
rect 23421 31635 23457 31669
rect 23491 31635 23527 31669
rect 23561 31635 23597 31669
rect 23631 31635 23635 31669
rect 22966 31608 23034 31635
rect 23068 31608 23635 31635
rect 22823 31601 23635 31608
rect 22823 31567 22827 31601
rect 22861 31568 22897 31601
rect 22864 31567 22897 31568
rect 22931 31568 22967 31601
rect 22931 31567 22932 31568
rect 22823 31534 22830 31567
rect 22864 31534 22932 31567
rect 22966 31567 22967 31568
rect 23001 31568 23037 31601
rect 23001 31567 23034 31568
rect 23071 31567 23107 31601
rect 23141 31567 23177 31601
rect 23211 31567 23247 31601
rect 23281 31567 23317 31601
rect 23351 31567 23387 31601
rect 23421 31567 23457 31601
rect 23491 31567 23527 31601
rect 23561 31567 23597 31601
rect 23631 31567 23635 31601
rect 22966 31534 23034 31567
rect 23068 31534 23635 31567
rect 22823 31533 23635 31534
rect 22823 31499 22827 31533
rect 22861 31499 22897 31533
rect 22931 31499 22967 31533
rect 23001 31499 23037 31533
rect 23071 31499 23107 31533
rect 23141 31499 23177 31533
rect 23211 31499 23247 31533
rect 23281 31499 23317 31533
rect 23351 31499 23387 31533
rect 23421 31499 23457 31533
rect 23491 31499 23527 31533
rect 23561 31499 23597 31533
rect 23631 31499 23635 31533
rect 22823 31494 23635 31499
rect 22823 31465 22830 31494
rect 22864 31465 22932 31494
rect 22823 31431 22827 31465
rect 22864 31460 22897 31465
rect 22861 31431 22897 31460
rect 22931 31460 22932 31465
rect 22966 31465 23034 31494
rect 23068 31465 23635 31494
rect 22966 31460 22967 31465
rect 22931 31431 22967 31460
rect 23001 31460 23034 31465
rect 23001 31431 23037 31460
rect 23071 31431 23107 31465
rect 23141 31431 23177 31465
rect 23211 31431 23247 31465
rect 23281 31431 23317 31465
rect 23351 31431 23387 31465
rect 23421 31431 23457 31465
rect 23491 31431 23527 31465
rect 23561 31431 23597 31465
rect 23631 31431 23635 31465
rect 22823 31420 23635 31431
rect 22823 31397 22830 31420
rect 22864 31397 22932 31420
rect 22823 31363 22827 31397
rect 22864 31386 22897 31397
rect 22861 31363 22897 31386
rect 22931 31386 22932 31397
rect 22966 31397 23034 31420
rect 23068 31397 23635 31420
rect 22966 31386 22967 31397
rect 22931 31363 22967 31386
rect 23001 31386 23034 31397
rect 23001 31363 23037 31386
rect 23071 31363 23107 31397
rect 23141 31363 23177 31397
rect 23211 31363 23247 31397
rect 23281 31363 23317 31397
rect 23351 31363 23387 31397
rect 23421 31363 23457 31397
rect 23491 31363 23527 31397
rect 23561 31363 23597 31397
rect 23631 31363 23635 31397
rect 22823 31346 23635 31363
rect 22823 31329 22830 31346
rect 22864 31329 22932 31346
rect 22823 31295 22827 31329
rect 22864 31312 22897 31329
rect 22861 31295 22897 31312
rect 22931 31312 22932 31329
rect 22966 31329 23034 31346
rect 23068 31329 23635 31346
rect 22966 31312 22967 31329
rect 22931 31295 22967 31312
rect 23001 31312 23034 31329
rect 23001 31295 23037 31312
rect 23071 31295 23107 31329
rect 23141 31295 23177 31329
rect 23211 31295 23247 31329
rect 23281 31295 23317 31329
rect 23351 31295 23387 31329
rect 23421 31295 23457 31329
rect 23491 31295 23527 31329
rect 23561 31295 23597 31329
rect 23631 31295 23635 31329
rect 22823 31271 23635 31295
rect 22823 31261 22830 31271
rect 22864 31261 22932 31271
rect 22823 31227 22827 31261
rect 22864 31237 22897 31261
rect 22861 31227 22897 31237
rect 22931 31237 22932 31261
rect 22966 31261 23034 31271
rect 23068 31261 23635 31271
rect 22966 31237 22967 31261
rect 22931 31227 22967 31237
rect 23001 31237 23034 31261
rect 23001 31227 23037 31237
rect 23071 31227 23107 31261
rect 23141 31227 23177 31261
rect 23211 31227 23247 31261
rect 23281 31227 23317 31261
rect 23351 31227 23387 31261
rect 23421 31227 23457 31261
rect 23491 31227 23527 31261
rect 23561 31227 23597 31261
rect 23631 31227 23635 31261
rect 22823 31196 23635 31227
rect 22823 31193 22830 31196
rect 22864 31193 22932 31196
rect 22823 31159 22827 31193
rect 22864 31162 22897 31193
rect 22861 31159 22897 31162
rect 22931 31162 22932 31193
rect 22966 31193 23034 31196
rect 23068 31193 23635 31196
rect 22966 31162 22967 31193
rect 22931 31159 22967 31162
rect 23001 31162 23034 31193
rect 23001 31159 23037 31162
rect 23071 31159 23107 31193
rect 23141 31159 23177 31193
rect 23211 31159 23247 31193
rect 23281 31159 23317 31193
rect 23351 31159 23387 31193
rect 23421 31159 23457 31193
rect 23491 31159 23527 31193
rect 23561 31159 23597 31193
rect 23631 31159 23635 31193
rect 22823 31125 23635 31159
rect 22823 31091 22827 31125
rect 22861 31121 22897 31125
rect 22864 31091 22897 31121
rect 22931 31121 22967 31125
rect 22931 31091 22932 31121
rect 22823 31087 22830 31091
rect 22864 31087 22932 31091
rect 22966 31091 22967 31121
rect 23001 31121 23037 31125
rect 23001 31091 23034 31121
rect 23071 31091 23107 31125
rect 23141 31091 23177 31125
rect 23211 31091 23247 31125
rect 23281 31091 23317 31125
rect 23351 31091 23387 31125
rect 23421 31091 23457 31125
rect 23491 31091 23527 31125
rect 23561 31091 23597 31125
rect 23631 31091 23635 31125
rect 22966 31087 23034 31091
rect 23068 31087 23635 31091
rect 22823 31057 23635 31087
rect 22823 31023 22827 31057
rect 22861 31046 22897 31057
rect 22864 31023 22897 31046
rect 22931 31046 22967 31057
rect 22931 31023 22932 31046
rect 22823 31012 22830 31023
rect 22864 31012 22932 31023
rect 22966 31023 22967 31046
rect 23001 31046 23037 31057
rect 23001 31023 23034 31046
rect 23071 31023 23107 31057
rect 23141 31023 23177 31057
rect 23211 31023 23247 31057
rect 23281 31023 23317 31057
rect 23351 31023 23387 31057
rect 23421 31023 23457 31057
rect 23491 31023 23527 31057
rect 23561 31023 23597 31057
rect 23631 31023 23635 31057
rect 22966 31012 23034 31023
rect 23068 31012 23635 31023
rect 22823 30989 23635 31012
rect 22823 30955 22827 30989
rect 22861 30971 22897 30989
rect 22864 30955 22897 30971
rect 22931 30971 22967 30989
rect 22931 30955 22932 30971
rect 22823 30937 22830 30955
rect 22864 30937 22932 30955
rect 22966 30955 22967 30971
rect 23001 30971 23037 30989
rect 23001 30955 23034 30971
rect 23071 30955 23107 30989
rect 23141 30955 23177 30989
rect 23211 30955 23247 30989
rect 23281 30955 23317 30989
rect 23351 30955 23387 30989
rect 23421 30955 23457 30989
rect 23491 30955 23527 30989
rect 23561 30955 23597 30989
rect 23631 30955 23635 30989
rect 22966 30937 23034 30955
rect 23068 30937 23635 30955
rect 22823 30921 23635 30937
rect 22823 30887 22827 30921
rect 22861 30896 22897 30921
rect 22864 30887 22897 30896
rect 22931 30896 22967 30921
rect 22931 30887 22932 30896
rect 22823 30862 22830 30887
rect 22864 30862 22932 30887
rect 22966 30887 22967 30896
rect 23001 30896 23037 30921
rect 23001 30887 23034 30896
rect 23071 30887 23107 30921
rect 23141 30887 23177 30921
rect 23211 30887 23247 30921
rect 23281 30887 23317 30921
rect 23351 30887 23387 30921
rect 23421 30887 23457 30921
rect 23491 30887 23527 30921
rect 23561 30887 23597 30921
rect 23631 30887 23635 30921
rect 22966 30862 23034 30887
rect 23068 30862 23635 30887
rect 22823 30853 23635 30862
rect 22823 30819 22827 30853
rect 22861 30821 22897 30853
rect 22864 30819 22897 30821
rect 22931 30821 22967 30853
rect 22931 30819 22932 30821
rect 22823 30787 22830 30819
rect 22864 30787 22932 30819
rect 22966 30819 22967 30821
rect 23001 30821 23037 30853
rect 23001 30819 23034 30821
rect 23071 30819 23107 30853
rect 23141 30819 23177 30853
rect 23211 30819 23247 30853
rect 23281 30819 23317 30853
rect 23351 30819 23387 30853
rect 23421 30819 23457 30853
rect 23491 30819 23527 30853
rect 23561 30819 23597 30853
rect 23631 30819 23635 30853
rect 22966 30787 23034 30819
rect 23068 30787 23635 30819
rect 22823 30785 23635 30787
rect 22823 30751 22827 30785
rect 22861 30751 22897 30785
rect 22931 30751 22967 30785
rect 23001 30751 23037 30785
rect 23071 30751 23107 30785
rect 23141 30751 23177 30785
rect 23211 30751 23247 30785
rect 23281 30751 23317 30785
rect 23351 30751 23387 30785
rect 23421 30751 23457 30785
rect 23491 30751 23527 30785
rect 23561 30751 23597 30785
rect 23631 30751 23635 30785
rect 22823 30746 23635 30751
rect 22823 30717 22830 30746
rect 22864 30717 22932 30746
rect 18439 30689 19012 30705
rect 18021 30671 19012 30689
rect 18021 30664 18486 30671
rect 18021 30630 18022 30664
rect 18056 30655 18108 30664
rect 18142 30655 18194 30664
rect 18228 30655 18280 30664
rect 18314 30655 18366 30664
rect 18021 30621 18025 30630
rect 18059 30621 18101 30655
rect 18142 30630 18177 30655
rect 18228 30630 18253 30655
rect 18314 30630 18329 30655
rect 18135 30621 18177 30630
rect 18211 30621 18253 30630
rect 18287 30621 18329 30630
rect 18363 30630 18366 30655
rect 18400 30655 18486 30664
rect 18400 30630 18405 30655
rect 18363 30621 18405 30630
rect 18439 30637 18486 30655
rect 18520 30637 18556 30671
rect 18590 30637 18626 30671
rect 18660 30637 18696 30671
rect 18730 30637 18766 30671
rect 18800 30637 18836 30671
rect 18870 30637 18906 30671
rect 18940 30637 18976 30671
rect 19010 30637 19012 30671
rect 18439 30621 19012 30637
rect 18021 30603 19012 30621
rect 18021 30592 18486 30603
rect 18021 30558 18022 30592
rect 18056 30587 18108 30592
rect 18142 30587 18194 30592
rect 18228 30587 18280 30592
rect 18314 30587 18366 30592
rect 18021 30553 18025 30558
rect 18059 30553 18101 30587
rect 18142 30558 18177 30587
rect 18228 30558 18253 30587
rect 18314 30558 18329 30587
rect 18135 30553 18177 30558
rect 18211 30553 18253 30558
rect 18287 30553 18329 30558
rect 18363 30558 18366 30587
rect 18400 30587 18486 30592
rect 18400 30558 18405 30587
rect 18363 30553 18405 30558
rect 18439 30569 18486 30587
rect 18520 30569 18556 30603
rect 18590 30569 18626 30603
rect 18660 30569 18696 30603
rect 18730 30569 18766 30603
rect 18800 30569 18836 30603
rect 18870 30569 18906 30603
rect 18940 30569 18976 30603
rect 19010 30569 19012 30603
rect 18439 30553 19012 30569
rect 18021 30535 19012 30553
rect 18021 30520 18486 30535
rect 18021 30486 18022 30520
rect 18056 30519 18108 30520
rect 18142 30519 18194 30520
rect 18228 30519 18280 30520
rect 18314 30519 18366 30520
rect 18021 30485 18025 30486
rect 18059 30485 18101 30519
rect 18142 30486 18177 30519
rect 18228 30486 18253 30519
rect 18314 30486 18329 30519
rect 18135 30485 18177 30486
rect 18211 30485 18253 30486
rect 18287 30485 18329 30486
rect 18363 30486 18366 30519
rect 18400 30519 18486 30520
rect 18400 30486 18405 30519
rect 18363 30485 18405 30486
rect 18439 30501 18486 30519
rect 18520 30501 18556 30535
rect 18590 30501 18626 30535
rect 18660 30501 18696 30535
rect 18730 30501 18766 30535
rect 18800 30501 18836 30535
rect 18870 30501 18906 30535
rect 18940 30501 18976 30535
rect 19010 30501 19012 30535
rect 18439 30485 19012 30501
rect 18021 30467 19012 30485
rect 18021 30451 18486 30467
rect 18021 30448 18025 30451
rect 18021 30414 18022 30448
rect 18059 30417 18101 30451
rect 18135 30448 18177 30451
rect 18211 30448 18253 30451
rect 18287 30448 18329 30451
rect 18142 30417 18177 30448
rect 18228 30417 18253 30448
rect 18314 30417 18329 30448
rect 18363 30448 18405 30451
rect 18363 30417 18366 30448
rect 18056 30414 18108 30417
rect 18142 30414 18194 30417
rect 18228 30414 18280 30417
rect 18314 30414 18366 30417
rect 18400 30417 18405 30448
rect 18439 30433 18486 30451
rect 18520 30433 18556 30467
rect 18590 30433 18626 30467
rect 18660 30433 18696 30467
rect 18730 30433 18766 30467
rect 18800 30433 18836 30467
rect 18870 30433 18906 30467
rect 18940 30433 18976 30467
rect 19010 30433 19012 30467
rect 18439 30417 19012 30433
rect 18400 30414 19012 30417
rect 18021 30399 19012 30414
rect 18021 30383 18486 30399
rect 18021 30376 18025 30383
rect 18021 30342 18022 30376
rect 18059 30349 18101 30383
rect 18135 30376 18177 30383
rect 18211 30376 18253 30383
rect 18287 30376 18329 30383
rect 18142 30349 18177 30376
rect 18228 30349 18253 30376
rect 18314 30349 18329 30376
rect 18363 30376 18405 30383
rect 18363 30349 18366 30376
rect 18056 30342 18108 30349
rect 18142 30342 18194 30349
rect 18228 30342 18280 30349
rect 18314 30342 18366 30349
rect 18400 30349 18405 30376
rect 18439 30365 18486 30383
rect 18520 30365 18556 30399
rect 18590 30365 18626 30399
rect 18660 30365 18696 30399
rect 18730 30365 18766 30399
rect 18800 30365 18836 30399
rect 18870 30365 18906 30399
rect 18940 30365 18976 30399
rect 19010 30365 19012 30399
rect 18439 30349 19012 30365
rect 18400 30342 19012 30349
rect 18021 30331 19012 30342
rect 18021 30315 18486 30331
rect 18021 30304 18025 30315
rect 18021 30270 18022 30304
rect 18059 30281 18101 30315
rect 18135 30304 18177 30315
rect 18211 30304 18253 30315
rect 18287 30304 18329 30315
rect 18142 30281 18177 30304
rect 18228 30281 18253 30304
rect 18314 30281 18329 30304
rect 18363 30304 18405 30315
rect 18363 30281 18366 30304
rect 18056 30270 18108 30281
rect 18142 30270 18194 30281
rect 18228 30270 18280 30281
rect 18314 30270 18366 30281
rect 18400 30281 18405 30304
rect 18439 30297 18486 30315
rect 18520 30297 18556 30331
rect 18590 30297 18626 30331
rect 18660 30297 18696 30331
rect 18730 30297 18766 30331
rect 18800 30297 18836 30331
rect 18870 30297 18906 30331
rect 18940 30297 18976 30331
rect 19010 30297 19012 30331
rect 18439 30281 19012 30297
rect 18400 30270 19012 30281
rect 18021 30263 19012 30270
rect 18021 30247 18486 30263
rect 18021 30232 18025 30247
rect 18021 30198 18022 30232
rect 18059 30213 18101 30247
rect 18135 30232 18177 30247
rect 18211 30232 18253 30247
rect 18287 30232 18329 30247
rect 18142 30213 18177 30232
rect 18228 30213 18253 30232
rect 18314 30213 18329 30232
rect 18363 30232 18405 30247
rect 18363 30213 18366 30232
rect 18056 30198 18108 30213
rect 18142 30198 18194 30213
rect 18228 30198 18280 30213
rect 18314 30198 18366 30213
rect 18400 30213 18405 30232
rect 18439 30229 18486 30247
rect 18520 30229 18556 30263
rect 18590 30229 18626 30263
rect 18660 30229 18696 30263
rect 18730 30229 18766 30263
rect 18800 30229 18836 30263
rect 18870 30229 18906 30263
rect 18940 30229 18976 30263
rect 19010 30229 19012 30263
rect 18439 30213 19012 30229
rect 18400 30198 19012 30213
rect 18021 30195 19012 30198
rect 18021 30179 18486 30195
rect 18021 30160 18025 30179
rect 18021 30126 18022 30160
rect 18059 30145 18101 30179
rect 18135 30160 18177 30179
rect 18211 30160 18253 30179
rect 18287 30160 18329 30179
rect 18142 30145 18177 30160
rect 18228 30145 18253 30160
rect 18314 30145 18329 30160
rect 18363 30160 18405 30179
rect 18363 30145 18366 30160
rect 18056 30126 18108 30145
rect 18142 30126 18194 30145
rect 18228 30126 18280 30145
rect 18314 30126 18366 30145
rect 18400 30145 18405 30160
rect 18439 30161 18486 30179
rect 18520 30161 18556 30195
rect 18590 30161 18626 30195
rect 18660 30161 18696 30195
rect 18730 30161 18766 30195
rect 18800 30161 18836 30195
rect 18870 30161 18906 30195
rect 18940 30161 18976 30195
rect 19010 30161 19012 30195
rect 18439 30145 19012 30161
rect 18400 30127 19012 30145
rect 18400 30126 18486 30127
rect 18021 30111 18486 30126
rect 18021 30088 18025 30111
rect 18021 30054 18022 30088
rect 18059 30077 18101 30111
rect 18135 30088 18177 30111
rect 18211 30088 18253 30111
rect 18287 30088 18329 30111
rect 18142 30077 18177 30088
rect 18228 30077 18253 30088
rect 18314 30077 18329 30088
rect 18363 30088 18405 30111
rect 18363 30077 18366 30088
rect 18056 30054 18108 30077
rect 18142 30054 18194 30077
rect 18228 30054 18280 30077
rect 18314 30054 18366 30077
rect 18400 30077 18405 30088
rect 18439 30093 18486 30111
rect 18520 30093 18556 30127
rect 18590 30093 18626 30127
rect 18660 30093 18696 30127
rect 18730 30093 18766 30127
rect 18800 30093 18836 30127
rect 18870 30093 18906 30127
rect 18940 30093 18976 30127
rect 19010 30093 19012 30127
rect 18439 30077 19012 30093
rect 18400 30059 19012 30077
rect 18400 30054 18486 30059
rect 18021 30043 18486 30054
rect 18021 30016 18025 30043
rect 18021 29982 18022 30016
rect 18059 30009 18101 30043
rect 18135 30016 18177 30043
rect 18211 30016 18253 30043
rect 18287 30016 18329 30043
rect 18142 30009 18177 30016
rect 18228 30009 18253 30016
rect 18314 30009 18329 30016
rect 18363 30016 18405 30043
rect 18363 30009 18366 30016
rect 18056 29982 18108 30009
rect 18142 29982 18194 30009
rect 18228 29982 18280 30009
rect 18314 29982 18366 30009
rect 18400 30009 18405 30016
rect 18439 30025 18486 30043
rect 18520 30025 18556 30059
rect 18590 30025 18626 30059
rect 18660 30025 18696 30059
rect 18730 30025 18766 30059
rect 18800 30025 18836 30059
rect 18870 30025 18906 30059
rect 18940 30025 18976 30059
rect 19010 30025 19012 30059
rect 18439 30009 19012 30025
rect 18400 29991 19012 30009
rect 18400 29982 18486 29991
rect 18021 29975 18486 29982
rect 18021 29944 18025 29975
rect 18021 29910 18022 29944
rect 18059 29941 18101 29975
rect 18135 29944 18177 29975
rect 18211 29944 18253 29975
rect 18287 29944 18329 29975
rect 18142 29941 18177 29944
rect 18228 29941 18253 29944
rect 18314 29941 18329 29944
rect 18363 29944 18405 29975
rect 18363 29941 18366 29944
rect 18056 29910 18108 29941
rect 18142 29910 18194 29941
rect 18228 29910 18280 29941
rect 18314 29910 18366 29941
rect 18400 29941 18405 29944
rect 18439 29957 18486 29975
rect 18520 29957 18556 29991
rect 18590 29957 18626 29991
rect 18660 29957 18696 29991
rect 18730 29957 18766 29991
rect 18800 29957 18836 29991
rect 18870 29957 18906 29991
rect 18940 29957 18976 29991
rect 19010 29957 19012 29991
rect 18439 29941 19012 29957
rect 18400 29923 19012 29941
rect 18400 29910 18486 29923
rect 18021 29907 18486 29910
rect 18021 29873 18025 29907
rect 18059 29873 18101 29907
rect 18135 29873 18177 29907
rect 18211 29873 18253 29907
rect 18287 29873 18329 29907
rect 18363 29873 18405 29907
rect 18439 29889 18486 29907
rect 18520 29889 18556 29923
rect 18590 29889 18626 29923
rect 18660 29889 18696 29923
rect 18730 29889 18766 29923
rect 18800 29889 18836 29923
rect 18870 29889 18906 29923
rect 18940 29889 18976 29923
rect 19010 29889 19012 29923
rect 18439 29873 19012 29889
rect 18021 29872 19012 29873
rect 18021 29838 18022 29872
rect 18056 29839 18108 29872
rect 18142 29839 18194 29872
rect 18228 29839 18280 29872
rect 18314 29839 18366 29872
rect 18021 29805 18025 29838
rect 18059 29805 18101 29839
rect 18142 29838 18177 29839
rect 18228 29838 18253 29839
rect 18314 29838 18329 29839
rect 18135 29805 18177 29838
rect 18211 29805 18253 29838
rect 18287 29805 18329 29838
rect 18363 29838 18366 29839
rect 18400 29855 19012 29872
rect 18400 29839 18486 29855
rect 18400 29838 18405 29839
rect 18363 29805 18405 29838
rect 18439 29821 18486 29839
rect 18520 29821 18556 29855
rect 18590 29821 18626 29855
rect 18660 29821 18696 29855
rect 18730 29821 18766 29855
rect 18800 29821 18836 29855
rect 18870 29821 18906 29855
rect 18940 29821 18976 29855
rect 19010 29821 19012 29855
rect 18439 29805 19012 29821
rect 18021 29800 19012 29805
rect 18021 29766 18022 29800
rect 18056 29771 18108 29800
rect 18142 29771 18194 29800
rect 18228 29771 18280 29800
rect 18314 29771 18366 29800
rect 18021 29737 18025 29766
rect 18059 29737 18101 29771
rect 18142 29766 18177 29771
rect 18228 29766 18253 29771
rect 18314 29766 18329 29771
rect 18135 29737 18177 29766
rect 18211 29737 18253 29766
rect 18287 29737 18329 29766
rect 18363 29766 18366 29771
rect 18400 29787 19012 29800
rect 18400 29771 18486 29787
rect 18400 29766 18405 29771
rect 18363 29737 18405 29766
rect 18439 29753 18486 29771
rect 18520 29753 18556 29787
rect 18590 29753 18626 29787
rect 18660 29753 18696 29787
rect 18730 29753 18766 29787
rect 18800 29753 18836 29787
rect 18870 29753 18906 29787
rect 18940 29753 18976 29787
rect 19010 29753 19012 29787
rect 18439 29737 19012 29753
rect 18021 29728 19012 29737
rect 18021 29694 18022 29728
rect 18056 29703 18108 29728
rect 18142 29703 18194 29728
rect 18228 29703 18280 29728
rect 18314 29703 18366 29728
rect 18021 29669 18025 29694
rect 18059 29669 18101 29703
rect 18142 29694 18177 29703
rect 18228 29694 18253 29703
rect 18314 29694 18329 29703
rect 18135 29669 18177 29694
rect 18211 29669 18253 29694
rect 18287 29669 18329 29694
rect 18363 29694 18366 29703
rect 18400 29719 19012 29728
rect 18400 29703 18486 29719
rect 18400 29694 18405 29703
rect 18363 29669 18405 29694
rect 18439 29685 18486 29703
rect 18520 29685 18556 29719
rect 18590 29685 18626 29719
rect 18660 29685 18696 29719
rect 18730 29685 18766 29719
rect 18800 29685 18836 29719
rect 18870 29685 18906 29719
rect 18940 29685 18976 29719
rect 19010 29685 19012 29719
rect 18439 29669 19012 29685
rect 18021 29656 19012 29669
rect 18021 29622 18022 29656
rect 18056 29635 18108 29656
rect 18142 29635 18194 29656
rect 18228 29635 18280 29656
rect 18314 29635 18366 29656
rect 18021 29601 18025 29622
rect 18059 29601 18101 29635
rect 18142 29622 18177 29635
rect 18228 29622 18253 29635
rect 18314 29622 18329 29635
rect 18135 29601 18177 29622
rect 18211 29601 18253 29622
rect 18287 29601 18329 29622
rect 18363 29622 18366 29635
rect 18400 29651 19012 29656
rect 18400 29635 18486 29651
rect 18400 29622 18405 29635
rect 18363 29601 18405 29622
rect 18439 29617 18486 29635
rect 18520 29617 18556 29651
rect 18590 29617 18626 29651
rect 18660 29617 18696 29651
rect 18730 29617 18766 29651
rect 18800 29617 18836 29651
rect 18870 29617 18906 29651
rect 18940 29617 18976 29651
rect 19010 29617 19012 29651
rect 18439 29601 19012 29617
rect 18021 29584 19012 29601
rect 18021 29550 18022 29584
rect 18056 29567 18108 29584
rect 18142 29567 18194 29584
rect 18228 29567 18280 29584
rect 18314 29567 18366 29584
rect 18021 29533 18025 29550
rect 18059 29533 18101 29567
rect 18142 29550 18177 29567
rect 18228 29550 18253 29567
rect 18314 29550 18329 29567
rect 18135 29533 18177 29550
rect 18211 29533 18253 29550
rect 18287 29533 18329 29550
rect 18363 29550 18366 29567
rect 18400 29583 19012 29584
rect 18400 29567 18486 29583
rect 18400 29550 18405 29567
rect 18363 29533 18405 29550
rect 18439 29549 18486 29567
rect 18520 29549 18556 29583
rect 18590 29549 18626 29583
rect 18660 29549 18696 29583
rect 18730 29549 18766 29583
rect 18800 29549 18836 29583
rect 18870 29549 18906 29583
rect 18940 29549 18976 29583
rect 19010 29549 19012 29583
rect 18439 29533 19012 29549
rect 18021 29515 19012 29533
rect 18021 29512 18486 29515
rect 18021 29478 18022 29512
rect 18056 29499 18108 29512
rect 18142 29499 18194 29512
rect 18228 29499 18280 29512
rect 18314 29499 18366 29512
rect 18021 29465 18025 29478
rect 18059 29465 18101 29499
rect 18142 29478 18177 29499
rect 18228 29478 18253 29499
rect 18314 29478 18329 29499
rect 18135 29465 18177 29478
rect 18211 29465 18253 29478
rect 18287 29465 18329 29478
rect 18363 29478 18366 29499
rect 18400 29499 18486 29512
rect 18400 29478 18405 29499
rect 18363 29465 18405 29478
rect 18439 29481 18486 29499
rect 18520 29481 18556 29515
rect 18590 29481 18626 29515
rect 18660 29481 18696 29515
rect 18730 29481 18766 29515
rect 18800 29481 18836 29515
rect 18870 29481 18906 29515
rect 18940 29481 18976 29515
rect 19010 29481 19012 29515
rect 18439 29465 19012 29481
rect 18021 29447 19012 29465
rect 18021 29440 18486 29447
rect 18021 29406 18022 29440
rect 18056 29431 18108 29440
rect 18142 29431 18194 29440
rect 18228 29431 18280 29440
rect 18314 29431 18366 29440
rect 18021 29397 18025 29406
rect 18059 29397 18101 29431
rect 18142 29406 18177 29431
rect 18228 29406 18253 29431
rect 18314 29406 18329 29431
rect 18135 29397 18177 29406
rect 18211 29397 18253 29406
rect 18287 29397 18329 29406
rect 18363 29406 18366 29431
rect 18400 29431 18486 29440
rect 18400 29406 18405 29431
rect 18363 29397 18405 29406
rect 18439 29413 18486 29431
rect 18520 29413 18556 29447
rect 18590 29413 18626 29447
rect 18660 29413 18696 29447
rect 18730 29413 18766 29447
rect 18800 29413 18836 29447
rect 18870 29413 18906 29447
rect 18940 29413 18976 29447
rect 19010 29413 19012 29447
rect 18439 29397 19012 29413
rect 18021 29379 19012 29397
rect 18021 29368 18486 29379
rect 18021 29334 18022 29368
rect 18056 29363 18108 29368
rect 18142 29363 18194 29368
rect 18228 29363 18280 29368
rect 18314 29363 18366 29368
rect 18021 29329 18025 29334
rect 18059 29329 18101 29363
rect 18142 29334 18177 29363
rect 18228 29334 18253 29363
rect 18314 29334 18329 29363
rect 18135 29329 18177 29334
rect 18211 29329 18253 29334
rect 18287 29329 18329 29334
rect 18363 29334 18366 29363
rect 18400 29363 18486 29368
rect 18400 29334 18405 29363
rect 18363 29329 18405 29334
rect 18439 29345 18486 29363
rect 18520 29345 18556 29379
rect 18590 29345 18626 29379
rect 18660 29345 18696 29379
rect 18730 29345 18766 29379
rect 18800 29345 18836 29379
rect 18870 29345 18906 29379
rect 18940 29345 18976 29379
rect 19010 29345 19012 29379
rect 18439 29329 19012 29345
rect 18021 29311 19012 29329
rect 18021 29296 18486 29311
rect 18021 29262 18022 29296
rect 18056 29295 18108 29296
rect 18142 29295 18194 29296
rect 18228 29295 18280 29296
rect 18314 29295 18366 29296
rect 18021 29261 18025 29262
rect 18059 29261 18101 29295
rect 18142 29262 18177 29295
rect 18228 29262 18253 29295
rect 18314 29262 18329 29295
rect 18135 29261 18177 29262
rect 18211 29261 18253 29262
rect 18287 29261 18329 29262
rect 18363 29262 18366 29295
rect 18400 29295 18486 29296
rect 18400 29262 18405 29295
rect 18363 29261 18405 29262
rect 18439 29277 18486 29295
rect 18520 29277 18556 29311
rect 18590 29277 18626 29311
rect 18660 29277 18696 29311
rect 18730 29277 18766 29311
rect 18800 29277 18836 29311
rect 18870 29277 18906 29311
rect 18940 29277 18976 29311
rect 19010 29277 19012 29311
rect 18439 29261 19012 29277
rect 18021 29243 19012 29261
rect 18021 29227 18486 29243
rect 18021 29224 18025 29227
rect 18021 29190 18022 29224
rect 18059 29193 18101 29227
rect 18135 29224 18177 29227
rect 18211 29224 18253 29227
rect 18287 29224 18329 29227
rect 18142 29193 18177 29224
rect 18228 29193 18253 29224
rect 18314 29193 18329 29224
rect 18363 29224 18405 29227
rect 18363 29193 18366 29224
rect 18056 29190 18108 29193
rect 18142 29190 18194 29193
rect 18228 29190 18280 29193
rect 18314 29190 18366 29193
rect 18400 29193 18405 29224
rect 18439 29209 18486 29227
rect 18520 29209 18556 29243
rect 18590 29209 18626 29243
rect 18660 29209 18696 29243
rect 18730 29209 18766 29243
rect 18800 29209 18836 29243
rect 18870 29209 18906 29243
rect 18940 29209 18976 29243
rect 19010 29209 19012 29243
rect 18439 29193 19012 29209
rect 18400 29190 19012 29193
rect 18021 29175 19012 29190
rect 18021 29159 18486 29175
rect 18021 29152 18025 29159
rect 18021 29118 18022 29152
rect 18059 29125 18101 29159
rect 18135 29152 18177 29159
rect 18211 29152 18253 29159
rect 18287 29152 18329 29159
rect 18142 29125 18177 29152
rect 18228 29125 18253 29152
rect 18314 29125 18329 29152
rect 18363 29152 18405 29159
rect 18363 29125 18366 29152
rect 18056 29118 18108 29125
rect 18142 29118 18194 29125
rect 18228 29118 18280 29125
rect 18314 29118 18366 29125
rect 18400 29125 18405 29152
rect 18439 29141 18486 29159
rect 18520 29141 18556 29175
rect 18590 29141 18626 29175
rect 18660 29141 18696 29175
rect 18730 29141 18766 29175
rect 18800 29141 18836 29175
rect 18870 29141 18906 29175
rect 18940 29141 18976 29175
rect 19010 29141 19012 29175
rect 18439 29125 19012 29141
rect 18400 29118 19012 29125
rect 18021 29107 19012 29118
rect 18021 29091 18486 29107
rect 18021 29080 18025 29091
rect 18021 29046 18022 29080
rect 18059 29057 18101 29091
rect 18135 29080 18177 29091
rect 18211 29080 18253 29091
rect 18287 29080 18329 29091
rect 18142 29057 18177 29080
rect 18228 29057 18253 29080
rect 18314 29057 18329 29080
rect 18363 29080 18405 29091
rect 18363 29057 18366 29080
rect 18056 29046 18108 29057
rect 18142 29046 18194 29057
rect 18228 29046 18280 29057
rect 18314 29046 18366 29057
rect 18400 29057 18405 29080
rect 18439 29073 18486 29091
rect 18520 29073 18556 29107
rect 18590 29073 18626 29107
rect 18660 29073 18696 29107
rect 18730 29073 18766 29107
rect 18800 29073 18836 29107
rect 18870 29073 18906 29107
rect 18940 29073 18976 29107
rect 19010 29073 19012 29107
rect 18439 29057 19012 29073
rect 18400 29046 19012 29057
rect 18021 29039 19012 29046
rect 18021 29023 18486 29039
rect 18021 29008 18025 29023
rect 18021 28974 18022 29008
rect 18059 28989 18101 29023
rect 18135 29008 18177 29023
rect 18211 29008 18253 29023
rect 18287 29008 18329 29023
rect 18142 28989 18177 29008
rect 18228 28989 18253 29008
rect 18314 28989 18329 29008
rect 18363 29008 18405 29023
rect 18363 28989 18366 29008
rect 18056 28974 18108 28989
rect 18142 28974 18194 28989
rect 18228 28974 18280 28989
rect 18314 28974 18366 28989
rect 18400 28989 18405 29008
rect 18439 29005 18486 29023
rect 18520 29005 18556 29039
rect 18590 29005 18626 29039
rect 18660 29005 18696 29039
rect 18730 29005 18766 29039
rect 18800 29005 18836 29039
rect 18870 29005 18906 29039
rect 18940 29005 18976 29039
rect 19010 29005 19012 29039
rect 18439 28989 19012 29005
rect 18400 28974 19012 28989
rect 18021 28971 19012 28974
rect 18021 28955 18486 28971
rect 18021 28936 18025 28955
rect 18021 28902 18022 28936
rect 18059 28921 18101 28955
rect 18135 28936 18177 28955
rect 18211 28936 18253 28955
rect 18287 28936 18329 28955
rect 18142 28921 18177 28936
rect 18228 28921 18253 28936
rect 18314 28921 18329 28936
rect 18363 28936 18405 28955
rect 18363 28921 18366 28936
rect 18056 28902 18108 28921
rect 18142 28902 18194 28921
rect 18228 28902 18280 28921
rect 18314 28902 18366 28921
rect 18400 28921 18405 28936
rect 18439 28937 18486 28955
rect 18520 28937 18556 28971
rect 18590 28937 18626 28971
rect 18660 28937 18696 28971
rect 18730 28937 18766 28971
rect 18800 28937 18836 28971
rect 18870 28937 18906 28971
rect 18940 28937 18976 28971
rect 19010 28937 19012 28971
rect 18439 28921 19012 28937
rect 18400 28903 19012 28921
rect 18400 28902 18486 28903
rect 18021 28887 18486 28902
rect 18021 28864 18025 28887
rect 18021 28830 18022 28864
rect 18059 28853 18101 28887
rect 18135 28864 18177 28887
rect 18211 28864 18253 28887
rect 18287 28864 18329 28887
rect 18142 28853 18177 28864
rect 18228 28853 18253 28864
rect 18314 28853 18329 28864
rect 18363 28864 18405 28887
rect 18363 28853 18366 28864
rect 18056 28830 18108 28853
rect 18142 28830 18194 28853
rect 18228 28830 18280 28853
rect 18314 28830 18366 28853
rect 18400 28853 18405 28864
rect 18439 28869 18486 28887
rect 18520 28869 18556 28903
rect 18590 28869 18626 28903
rect 18660 28869 18696 28903
rect 18730 28869 18766 28903
rect 18800 28869 18836 28903
rect 18870 28869 18906 28903
rect 18940 28869 18976 28903
rect 19010 28869 19012 28903
rect 18439 28853 19012 28869
rect 18400 28835 19012 28853
rect 18400 28830 18486 28835
rect 18021 28819 18486 28830
rect 18021 28792 18025 28819
rect 18021 28758 18022 28792
rect 18059 28785 18101 28819
rect 18135 28792 18177 28819
rect 18211 28792 18253 28819
rect 18287 28792 18329 28819
rect 18142 28785 18177 28792
rect 18228 28785 18253 28792
rect 18314 28785 18329 28792
rect 18363 28792 18405 28819
rect 18363 28785 18366 28792
rect 18056 28758 18108 28785
rect 18142 28758 18194 28785
rect 18228 28758 18280 28785
rect 18314 28758 18366 28785
rect 18400 28785 18405 28792
rect 18439 28801 18486 28819
rect 18520 28801 18556 28835
rect 18590 28801 18626 28835
rect 18660 28801 18696 28835
rect 18730 28801 18766 28835
rect 18800 28801 18836 28835
rect 18870 28801 18906 28835
rect 18940 28801 18976 28835
rect 19010 28801 19012 28835
rect 18439 28785 19012 28801
rect 18400 28767 19012 28785
rect 18400 28758 18486 28767
rect 18021 28751 18486 28758
rect 18021 28720 18025 28751
rect 18021 28686 18022 28720
rect 18059 28717 18101 28751
rect 18135 28720 18177 28751
rect 18211 28720 18253 28751
rect 18287 28720 18329 28751
rect 18142 28717 18177 28720
rect 18228 28717 18253 28720
rect 18314 28717 18329 28720
rect 18363 28720 18405 28751
rect 18363 28717 18366 28720
rect 18056 28686 18108 28717
rect 18142 28686 18194 28717
rect 18228 28686 18280 28717
rect 18314 28686 18366 28717
rect 18400 28717 18405 28720
rect 18439 28733 18486 28751
rect 18520 28733 18556 28767
rect 18590 28733 18626 28767
rect 18660 28733 18696 28767
rect 18730 28733 18766 28767
rect 18800 28733 18836 28767
rect 18870 28733 18906 28767
rect 18940 28733 18976 28767
rect 19010 28733 19012 28767
rect 18439 28717 19012 28733
rect 18400 28699 19012 28717
rect 18400 28686 18486 28699
rect 18021 28683 18486 28686
rect 18021 28649 18025 28683
rect 18059 28649 18101 28683
rect 18135 28649 18177 28683
rect 18211 28649 18253 28683
rect 18287 28649 18329 28683
rect 18363 28649 18405 28683
rect 18439 28665 18486 28683
rect 18520 28665 18556 28699
rect 18590 28665 18626 28699
rect 18660 28665 18696 28699
rect 18730 28665 18766 28699
rect 18800 28665 18836 28699
rect 18870 28665 18906 28699
rect 18940 28665 18976 28699
rect 19010 28665 19012 28699
rect 18439 28649 19012 28665
rect 18021 28648 19012 28649
rect 18021 28614 18022 28648
rect 18056 28615 18108 28648
rect 18142 28615 18194 28648
rect 18228 28615 18280 28648
rect 18314 28615 18366 28648
rect 18021 28581 18025 28614
rect 18059 28581 18101 28615
rect 18142 28614 18177 28615
rect 18228 28614 18253 28615
rect 18314 28614 18329 28615
rect 18135 28581 18177 28614
rect 18211 28581 18253 28614
rect 18287 28581 18329 28614
rect 18363 28614 18366 28615
rect 18400 28631 19012 28648
rect 18400 28615 18486 28631
rect 18400 28614 18405 28615
rect 18363 28581 18405 28614
rect 18439 28597 18486 28615
rect 18520 28597 18556 28631
rect 18590 28597 18626 28631
rect 18660 28597 18696 28631
rect 18730 28597 18766 28631
rect 18800 28597 18836 28631
rect 18870 28597 18906 28631
rect 18940 28597 18976 28631
rect 19010 28597 19012 28631
rect 18439 28581 19012 28597
rect 18021 28576 19012 28581
rect 18021 28542 18022 28576
rect 18056 28547 18108 28576
rect 18142 28547 18194 28576
rect 18228 28547 18280 28576
rect 18314 28547 18366 28576
rect 18021 28513 18025 28542
rect 18059 28513 18101 28547
rect 18142 28542 18177 28547
rect 18228 28542 18253 28547
rect 18314 28542 18329 28547
rect 18135 28513 18177 28542
rect 18211 28513 18253 28542
rect 18287 28513 18329 28542
rect 18363 28542 18366 28547
rect 18400 28563 19012 28576
rect 18400 28547 18486 28563
rect 18400 28542 18405 28547
rect 18363 28513 18405 28542
rect 18439 28529 18486 28547
rect 18520 28529 18556 28563
rect 18590 28529 18626 28563
rect 18660 28529 18696 28563
rect 18730 28529 18766 28563
rect 18800 28529 18836 28563
rect 18870 28529 18906 28563
rect 18940 28529 18976 28563
rect 19010 28529 19012 28563
rect 18439 28513 19012 28529
rect 18021 28504 19012 28513
rect 18021 28470 18022 28504
rect 18056 28479 18108 28504
rect 18142 28479 18194 28504
rect 18228 28479 18280 28504
rect 18314 28479 18366 28504
rect 18021 28445 18025 28470
rect 18059 28445 18101 28479
rect 18142 28470 18177 28479
rect 18228 28470 18253 28479
rect 18314 28470 18329 28479
rect 18135 28445 18177 28470
rect 18211 28445 18253 28470
rect 18287 28445 18329 28470
rect 18363 28470 18366 28479
rect 18400 28495 19012 28504
rect 18400 28479 18486 28495
rect 18400 28470 18405 28479
rect 18363 28445 18405 28470
rect 18439 28461 18486 28479
rect 18520 28461 18556 28495
rect 18590 28461 18626 28495
rect 18660 28461 18696 28495
rect 18730 28461 18766 28495
rect 18800 28461 18836 28495
rect 18870 28461 18906 28495
rect 18940 28461 18976 28495
rect 19010 28461 19012 28495
rect 18439 28445 19012 28461
rect 18021 28432 19012 28445
rect 18021 28398 18022 28432
rect 18056 28411 18108 28432
rect 18142 28411 18194 28432
rect 18228 28411 18280 28432
rect 18314 28411 18366 28432
rect 18021 28377 18025 28398
rect 18059 28377 18101 28411
rect 18142 28398 18177 28411
rect 18228 28398 18253 28411
rect 18314 28398 18329 28411
rect 18135 28377 18177 28398
rect 18211 28377 18253 28398
rect 18287 28377 18329 28398
rect 18363 28398 18366 28411
rect 18400 28427 19012 28432
rect 18400 28411 18486 28427
rect 18400 28398 18405 28411
rect 18363 28377 18405 28398
rect 18439 28393 18486 28411
rect 18520 28393 18556 28427
rect 18590 28393 18626 28427
rect 18660 28393 18696 28427
rect 18730 28393 18766 28427
rect 18800 28393 18836 28427
rect 18870 28393 18906 28427
rect 18940 28393 18976 28427
rect 19010 28393 19012 28427
rect 18439 28377 19012 28393
rect 18021 28360 19012 28377
rect 18021 28326 18022 28360
rect 18056 28343 18108 28360
rect 18142 28343 18194 28360
rect 18228 28343 18280 28360
rect 18314 28343 18366 28360
rect 18021 28309 18025 28326
rect 18059 28309 18101 28343
rect 18142 28326 18177 28343
rect 18228 28326 18253 28343
rect 18314 28326 18329 28343
rect 18135 28309 18177 28326
rect 18211 28309 18253 28326
rect 18287 28309 18329 28326
rect 18363 28326 18366 28343
rect 18400 28359 19012 28360
rect 18400 28343 18486 28359
rect 18400 28326 18405 28343
rect 18363 28309 18405 28326
rect 18439 28325 18486 28343
rect 18520 28325 18556 28359
rect 18590 28325 18626 28359
rect 18660 28325 18696 28359
rect 18730 28325 18766 28359
rect 18800 28325 18836 28359
rect 18870 28325 18906 28359
rect 18940 28325 18976 28359
rect 19010 28325 19012 28359
rect 18439 28309 19012 28325
rect 18021 28291 19012 28309
rect 18021 28288 18486 28291
rect 18021 28254 18022 28288
rect 18056 28275 18108 28288
rect 18142 28275 18194 28288
rect 18228 28275 18280 28288
rect 18314 28275 18366 28288
rect 18021 28241 18025 28254
rect 18059 28241 18101 28275
rect 18142 28254 18177 28275
rect 18228 28254 18253 28275
rect 18314 28254 18329 28275
rect 18135 28241 18177 28254
rect 18211 28241 18253 28254
rect 18287 28241 18329 28254
rect 18363 28254 18366 28275
rect 18400 28275 18486 28288
rect 18400 28254 18405 28275
rect 18363 28241 18405 28254
rect 18439 28257 18486 28275
rect 18520 28257 18556 28291
rect 18590 28257 18626 28291
rect 18660 28257 18696 28291
rect 18730 28257 18766 28291
rect 18800 28257 18836 28291
rect 18870 28257 18906 28291
rect 18940 28257 18976 28291
rect 19010 28257 19012 28291
rect 18439 28241 19012 28257
rect 18021 28223 19012 28241
rect 18021 28216 18486 28223
rect 18021 28182 18022 28216
rect 18056 28207 18108 28216
rect 18142 28207 18194 28216
rect 18228 28207 18280 28216
rect 18314 28207 18366 28216
rect 18021 28173 18025 28182
rect 18059 28173 18101 28207
rect 18142 28182 18177 28207
rect 18228 28182 18253 28207
rect 18314 28182 18329 28207
rect 18135 28173 18177 28182
rect 18211 28173 18253 28182
rect 18287 28173 18329 28182
rect 18363 28182 18366 28207
rect 18400 28207 18486 28216
rect 18400 28182 18405 28207
rect 18363 28173 18405 28182
rect 18439 28189 18486 28207
rect 18520 28189 18556 28223
rect 18590 28189 18626 28223
rect 18660 28189 18696 28223
rect 18730 28189 18766 28223
rect 18800 28189 18836 28223
rect 18870 28189 18906 28223
rect 18940 28189 18976 28223
rect 19010 28189 19012 28223
rect 18439 28173 19012 28189
rect 18021 28155 19012 28173
rect 18021 28144 18486 28155
rect 18021 28110 18022 28144
rect 18056 28139 18108 28144
rect 18142 28139 18194 28144
rect 18228 28139 18280 28144
rect 18314 28139 18366 28144
rect 18021 28105 18025 28110
rect 18059 28105 18101 28139
rect 18142 28110 18177 28139
rect 18228 28110 18253 28139
rect 18314 28110 18329 28139
rect 18135 28105 18177 28110
rect 18211 28105 18253 28110
rect 18287 28105 18329 28110
rect 18363 28110 18366 28139
rect 18400 28139 18486 28144
rect 18400 28110 18405 28139
rect 18363 28105 18405 28110
rect 18439 28121 18486 28139
rect 18520 28121 18556 28155
rect 18590 28121 18626 28155
rect 18660 28121 18696 28155
rect 18730 28121 18766 28155
rect 18800 28121 18836 28155
rect 18870 28121 18906 28155
rect 18940 28121 18976 28155
rect 19010 28121 19012 28155
rect 18439 28105 19012 28121
rect 18021 28087 19012 28105
rect 18021 28072 18486 28087
rect 18021 28038 18022 28072
rect 18056 28071 18108 28072
rect 18142 28071 18194 28072
rect 18228 28071 18280 28072
rect 18314 28071 18366 28072
rect 18021 28037 18025 28038
rect 18059 28037 18101 28071
rect 18142 28038 18177 28071
rect 18228 28038 18253 28071
rect 18314 28038 18329 28071
rect 18135 28037 18177 28038
rect 18211 28037 18253 28038
rect 18287 28037 18329 28038
rect 18363 28038 18366 28071
rect 18400 28071 18486 28072
rect 18400 28038 18405 28071
rect 18363 28037 18405 28038
rect 18439 28053 18486 28071
rect 18520 28053 18556 28087
rect 18590 28053 18626 28087
rect 18660 28053 18696 28087
rect 18730 28053 18766 28087
rect 18800 28053 18836 28087
rect 18870 28053 18906 28087
rect 18940 28053 18976 28087
rect 19010 28053 19012 28087
rect 18439 28037 19012 28053
rect 18021 28019 19012 28037
rect 18021 28003 18486 28019
rect 18021 28000 18025 28003
rect 18021 27966 18022 28000
rect 18059 27969 18101 28003
rect 18135 28000 18177 28003
rect 18211 28000 18253 28003
rect 18287 28000 18329 28003
rect 18142 27969 18177 28000
rect 18228 27969 18253 28000
rect 18314 27969 18329 28000
rect 18363 28000 18405 28003
rect 18363 27969 18366 28000
rect 18056 27966 18108 27969
rect 18142 27966 18194 27969
rect 18228 27966 18280 27969
rect 18314 27966 18366 27969
rect 18400 27969 18405 28000
rect 18439 27985 18486 28003
rect 18520 27985 18556 28019
rect 18590 27985 18626 28019
rect 18660 27985 18696 28019
rect 18730 27985 18766 28019
rect 18800 27985 18836 28019
rect 18870 27985 18906 28019
rect 18940 27985 18976 28019
rect 19010 27985 19012 28019
rect 18439 27969 19012 27985
rect 18400 27966 19012 27969
rect 18021 27951 19012 27966
rect 18021 27935 18486 27951
rect 18021 27928 18025 27935
rect 18021 27894 18022 27928
rect 18059 27901 18101 27935
rect 18135 27928 18177 27935
rect 18211 27928 18253 27935
rect 18287 27928 18329 27935
rect 18142 27901 18177 27928
rect 18228 27901 18253 27928
rect 18314 27901 18329 27928
rect 18363 27928 18405 27935
rect 18363 27901 18366 27928
rect 18056 27894 18108 27901
rect 18142 27894 18194 27901
rect 18228 27894 18280 27901
rect 18314 27894 18366 27901
rect 18400 27901 18405 27928
rect 18439 27917 18486 27935
rect 18520 27917 18556 27951
rect 18590 27917 18626 27951
rect 18660 27917 18696 27951
rect 18730 27917 18766 27951
rect 18800 27917 18836 27951
rect 18870 27917 18906 27951
rect 18940 27917 18976 27951
rect 19010 27917 19012 27951
rect 18439 27901 19012 27917
rect 18400 27894 19012 27901
rect 18021 27883 19012 27894
rect 18021 27867 18486 27883
rect 18021 27856 18025 27867
rect 18021 27822 18022 27856
rect 18059 27833 18101 27867
rect 18135 27856 18177 27867
rect 18211 27856 18253 27867
rect 18287 27856 18329 27867
rect 18142 27833 18177 27856
rect 18228 27833 18253 27856
rect 18314 27833 18329 27856
rect 18363 27856 18405 27867
rect 18363 27833 18366 27856
rect 18056 27822 18108 27833
rect 18142 27822 18194 27833
rect 18228 27822 18280 27833
rect 18314 27822 18366 27833
rect 18400 27833 18405 27856
rect 18439 27849 18486 27867
rect 18520 27849 18556 27883
rect 18590 27849 18626 27883
rect 18660 27849 18696 27883
rect 18730 27849 18766 27883
rect 18800 27849 18836 27883
rect 18870 27849 18906 27883
rect 18940 27849 18976 27883
rect 19010 27849 19012 27883
rect 18439 27833 19012 27849
rect 18400 27822 19012 27833
rect 18021 27815 19012 27822
rect 18021 27799 18486 27815
rect 18021 27784 18025 27799
rect 18021 27750 18022 27784
rect 18059 27765 18101 27799
rect 18135 27784 18177 27799
rect 18211 27784 18253 27799
rect 18287 27784 18329 27799
rect 18142 27765 18177 27784
rect 18228 27765 18253 27784
rect 18314 27765 18329 27784
rect 18363 27784 18405 27799
rect 18363 27765 18366 27784
rect 18056 27750 18108 27765
rect 18142 27750 18194 27765
rect 18228 27750 18280 27765
rect 18314 27750 18366 27765
rect 18400 27765 18405 27784
rect 18439 27781 18486 27799
rect 18520 27781 18556 27815
rect 18590 27781 18626 27815
rect 18660 27781 18696 27815
rect 18730 27781 18766 27815
rect 18800 27781 18836 27815
rect 18870 27781 18906 27815
rect 18940 27781 18976 27815
rect 19010 27781 19012 27815
rect 18439 27765 19012 27781
rect 18400 27750 19012 27765
rect 18021 27747 19012 27750
rect 18021 27731 18486 27747
rect 18021 27712 18025 27731
rect 18021 27678 18022 27712
rect 18059 27697 18101 27731
rect 18135 27712 18177 27731
rect 18211 27712 18253 27731
rect 18287 27712 18329 27731
rect 18142 27697 18177 27712
rect 18228 27697 18253 27712
rect 18314 27697 18329 27712
rect 18363 27712 18405 27731
rect 18363 27697 18366 27712
rect 18056 27678 18108 27697
rect 18142 27678 18194 27697
rect 18228 27678 18280 27697
rect 18314 27678 18366 27697
rect 18400 27697 18405 27712
rect 18439 27713 18486 27731
rect 18520 27713 18556 27747
rect 18590 27713 18626 27747
rect 18660 27713 18696 27747
rect 18730 27713 18766 27747
rect 18800 27713 18836 27747
rect 18870 27713 18906 27747
rect 18940 27713 18976 27747
rect 19010 27713 19012 27747
rect 18439 27697 19012 27713
rect 18400 27679 19012 27697
rect 18400 27678 18486 27679
rect 18021 27663 18486 27678
rect 18021 27640 18025 27663
rect 18021 27606 18022 27640
rect 18059 27629 18101 27663
rect 18135 27640 18177 27663
rect 18211 27640 18253 27663
rect 18287 27640 18329 27663
rect 18142 27629 18177 27640
rect 18228 27629 18253 27640
rect 18314 27629 18329 27640
rect 18363 27640 18405 27663
rect 18363 27629 18366 27640
rect 18056 27606 18108 27629
rect 18142 27606 18194 27629
rect 18228 27606 18280 27629
rect 18314 27606 18366 27629
rect 18400 27629 18405 27640
rect 18439 27645 18486 27663
rect 18520 27645 18556 27679
rect 18590 27645 18626 27679
rect 18660 27645 18696 27679
rect 18730 27645 18766 27679
rect 18800 27645 18836 27679
rect 18870 27645 18906 27679
rect 18940 27645 18976 27679
rect 19010 27645 19012 27679
rect 18439 27629 19012 27645
rect 18400 27611 19012 27629
rect 18400 27606 18486 27611
rect 18021 27595 18486 27606
rect 18021 27568 18025 27595
rect 18021 27534 18022 27568
rect 18059 27561 18101 27595
rect 18135 27568 18177 27595
rect 18211 27568 18253 27595
rect 18287 27568 18329 27595
rect 18142 27561 18177 27568
rect 18228 27561 18253 27568
rect 18314 27561 18329 27568
rect 18363 27568 18405 27595
rect 18363 27561 18366 27568
rect 18056 27534 18108 27561
rect 18142 27534 18194 27561
rect 18228 27534 18280 27561
rect 18314 27534 18366 27561
rect 18400 27561 18405 27568
rect 18439 27577 18486 27595
rect 18520 27577 18556 27611
rect 18590 27577 18626 27611
rect 18660 27577 18696 27611
rect 18730 27577 18766 27611
rect 18800 27577 18836 27611
rect 18870 27577 18906 27611
rect 18940 27577 18976 27611
rect 19010 27577 19012 27611
rect 18439 27561 19012 27577
rect 18400 27543 19012 27561
rect 18400 27534 18486 27543
rect 18021 27527 18486 27534
rect 18021 27496 18025 27527
rect 18021 27462 18022 27496
rect 18059 27493 18101 27527
rect 18135 27496 18177 27527
rect 18211 27496 18253 27527
rect 18287 27496 18329 27527
rect 18142 27493 18177 27496
rect 18228 27493 18253 27496
rect 18314 27493 18329 27496
rect 18363 27496 18405 27527
rect 18363 27493 18366 27496
rect 18056 27462 18108 27493
rect 18142 27462 18194 27493
rect 18228 27462 18280 27493
rect 18314 27462 18366 27493
rect 18400 27493 18405 27496
rect 18439 27509 18486 27527
rect 18520 27509 18556 27543
rect 18590 27509 18626 27543
rect 18660 27509 18696 27543
rect 18730 27509 18766 27543
rect 18800 27509 18836 27543
rect 18870 27509 18906 27543
rect 18940 27509 18976 27543
rect 19010 27509 19012 27543
rect 18439 27493 19012 27509
rect 18400 27475 19012 27493
rect 18400 27462 18486 27475
rect 18021 27459 18486 27462
rect 18021 27425 18025 27459
rect 18059 27425 18101 27459
rect 18135 27425 18177 27459
rect 18211 27425 18253 27459
rect 18287 27425 18329 27459
rect 18363 27425 18405 27459
rect 18439 27441 18486 27459
rect 18520 27441 18556 27475
rect 18590 27441 18626 27475
rect 18660 27441 18696 27475
rect 18730 27441 18766 27475
rect 18800 27441 18836 27475
rect 18870 27441 18906 27475
rect 18940 27441 18976 27475
rect 19010 27441 19012 27475
rect 18439 27425 19012 27441
rect 18021 27424 19012 27425
rect 18021 27390 18022 27424
rect 18056 27391 18108 27424
rect 18142 27391 18194 27424
rect 18228 27391 18280 27424
rect 18314 27391 18366 27424
rect 18021 27357 18025 27390
rect 18059 27357 18101 27391
rect 18142 27390 18177 27391
rect 18228 27390 18253 27391
rect 18314 27390 18329 27391
rect 18135 27357 18177 27390
rect 18211 27357 18253 27390
rect 18287 27357 18329 27390
rect 18363 27390 18366 27391
rect 18400 27407 19012 27424
rect 18400 27391 18486 27407
rect 18400 27390 18405 27391
rect 18363 27357 18405 27390
rect 18439 27373 18486 27391
rect 18520 27373 18556 27407
rect 18590 27373 18626 27407
rect 18660 27373 18696 27407
rect 18730 27373 18766 27407
rect 18800 27373 18836 27407
rect 18870 27373 18906 27407
rect 18940 27373 18976 27407
rect 19010 27373 19012 27407
rect 18439 27357 19012 27373
rect 18021 27352 19012 27357
rect 18021 27318 18022 27352
rect 18056 27323 18108 27352
rect 18142 27323 18194 27352
rect 18228 27323 18280 27352
rect 18314 27323 18366 27352
rect 18021 27289 18025 27318
rect 18059 27289 18101 27323
rect 18142 27318 18177 27323
rect 18228 27318 18253 27323
rect 18314 27318 18329 27323
rect 18135 27289 18177 27318
rect 18211 27289 18253 27318
rect 18287 27289 18329 27318
rect 18363 27318 18366 27323
rect 18400 27339 19012 27352
rect 18400 27323 18486 27339
rect 18400 27318 18405 27323
rect 18363 27289 18405 27318
rect 18439 27305 18486 27323
rect 18520 27305 18556 27339
rect 18590 27305 18626 27339
rect 18660 27305 18696 27339
rect 18730 27305 18766 27339
rect 18800 27305 18836 27339
rect 18870 27305 18906 27339
rect 18940 27305 18976 27339
rect 19010 27305 19012 27339
rect 18439 27289 19012 27305
rect 18021 27280 19012 27289
rect 18021 27246 18022 27280
rect 18056 27255 18108 27280
rect 18142 27255 18194 27280
rect 18228 27255 18280 27280
rect 18314 27255 18366 27280
rect 18021 27221 18025 27246
rect 18059 27221 18101 27255
rect 18142 27246 18177 27255
rect 18228 27246 18253 27255
rect 18314 27246 18329 27255
rect 18135 27221 18177 27246
rect 18211 27221 18253 27246
rect 18287 27221 18329 27246
rect 18363 27246 18366 27255
rect 18400 27271 19012 27280
rect 18400 27255 18486 27271
rect 18400 27246 18405 27255
rect 18363 27221 18405 27246
rect 18439 27237 18486 27255
rect 18520 27237 18556 27271
rect 18590 27237 18626 27271
rect 18660 27237 18696 27271
rect 18730 27237 18766 27271
rect 18800 27237 18836 27271
rect 18870 27237 18906 27271
rect 18940 27237 18976 27271
rect 19010 27237 19012 27271
rect 18439 27221 19012 27237
rect 18021 27208 19012 27221
rect 18021 27174 18022 27208
rect 18056 27187 18108 27208
rect 18142 27187 18194 27208
rect 18228 27187 18280 27208
rect 18314 27187 18366 27208
rect 18021 27153 18025 27174
rect 18059 27153 18101 27187
rect 18142 27174 18177 27187
rect 18228 27174 18253 27187
rect 18314 27174 18329 27187
rect 18135 27153 18177 27174
rect 18211 27153 18253 27174
rect 18287 27153 18329 27174
rect 18363 27174 18366 27187
rect 18400 27203 19012 27208
rect 18400 27187 18486 27203
rect 18400 27174 18405 27187
rect 18363 27153 18405 27174
rect 18439 27169 18486 27187
rect 18520 27169 18556 27203
rect 18590 27169 18626 27203
rect 18660 27169 18696 27203
rect 18730 27169 18766 27203
rect 18800 27169 18836 27203
rect 18870 27169 18906 27203
rect 18940 27169 18976 27203
rect 19010 27169 19012 27203
rect 18439 27153 19012 27169
rect 18021 27136 19012 27153
rect 999 27079 1758 27103
rect 999 27045 1057 27079
rect 1091 27045 1125 27079
rect 1159 27045 1193 27079
rect 1227 27045 1261 27079
rect 1295 27045 1329 27079
rect 1363 27045 1397 27079
rect 1431 27045 1465 27079
rect 1499 27045 1533 27079
rect 1567 27045 1601 27079
rect 1635 27045 1669 27079
rect 1703 27045 1758 27079
rect 999 27015 1758 27045
rect 999 27010 1470 27015
rect 1504 27010 1544 27015
rect 1578 27010 1618 27015
rect 1652 27010 1692 27015
rect 999 26976 1057 27010
rect 1091 26976 1125 27010
rect 1159 26976 1193 27010
rect 1227 26976 1261 27010
rect 1295 26976 1329 27010
rect 1363 27006 1397 27010
rect 1363 26976 1395 27006
rect 1431 26976 1465 27010
rect 1504 26981 1533 27010
rect 1578 26981 1601 27010
rect 1652 26981 1669 27010
rect 1726 26981 1758 27015
rect 1499 26976 1533 26981
rect 1567 26976 1601 26981
rect 1635 26976 1669 26981
rect 1703 26976 1758 26981
rect 999 26972 1395 26976
rect 1429 26972 1758 26976
rect 999 26943 1758 26972
rect 999 26941 1470 26943
rect 1504 26941 1544 26943
rect 1578 26941 1618 26943
rect 1652 26941 1692 26943
rect 999 26907 1057 26941
rect 1091 26907 1125 26941
rect 1159 26907 1193 26941
rect 1227 26907 1261 26941
rect 1295 26907 1329 26941
rect 1363 26932 1397 26941
rect 1363 26907 1395 26932
rect 1431 26907 1465 26941
rect 1504 26909 1533 26941
rect 1578 26909 1601 26941
rect 1652 26909 1669 26941
rect 1726 26909 1758 26943
rect 1499 26907 1533 26909
rect 1567 26907 1601 26909
rect 1635 26907 1669 26909
rect 1703 26907 1758 26909
rect 999 26898 1395 26907
rect 1429 26898 1758 26907
rect 999 26872 1758 26898
rect 999 26838 1057 26872
rect 1091 26838 1125 26872
rect 1159 26838 1193 26872
rect 1227 26838 1261 26872
rect 1295 26838 1329 26872
rect 1363 26858 1397 26872
rect 1363 26838 1395 26858
rect 1431 26838 1465 26872
rect 1499 26871 1533 26872
rect 1567 26871 1601 26872
rect 1635 26871 1669 26872
rect 1703 26871 1758 26872
rect 1504 26838 1533 26871
rect 1578 26838 1601 26871
rect 1652 26838 1669 26871
rect 999 26824 1395 26838
rect 1429 26837 1470 26838
rect 1504 26837 1544 26838
rect 1578 26837 1618 26838
rect 1652 26837 1692 26838
rect 1726 26837 1758 26871
rect 1429 26824 1758 26837
rect 999 26803 1758 26824
rect 999 26769 1057 26803
rect 1091 26769 1125 26803
rect 1159 26769 1193 26803
rect 1227 26769 1261 26803
rect 1295 26769 1329 26803
rect 1363 26784 1397 26803
rect 1363 26769 1395 26784
rect 1431 26769 1465 26803
rect 1499 26799 1533 26803
rect 1567 26799 1601 26803
rect 1635 26799 1669 26803
rect 1703 26799 1758 26803
rect 1504 26769 1533 26799
rect 1578 26769 1601 26799
rect 1652 26769 1669 26799
rect 999 26750 1395 26769
rect 1429 26765 1470 26769
rect 1504 26765 1544 26769
rect 1578 26765 1618 26769
rect 1652 26765 1692 26769
rect 1726 26765 1758 26799
rect 1429 26750 1758 26765
rect 999 26734 1758 26750
rect 999 26700 1057 26734
rect 1091 26700 1125 26734
rect 1159 26700 1193 26734
rect 1227 26700 1261 26734
rect 1295 26700 1329 26734
rect 1363 26710 1397 26734
rect 1363 26700 1395 26710
rect 1431 26700 1465 26734
rect 1499 26727 1533 26734
rect 1567 26727 1601 26734
rect 1635 26727 1669 26734
rect 1703 26727 1758 26734
rect 1504 26700 1533 26727
rect 1578 26700 1601 26727
rect 1652 26700 1669 26727
rect 999 26676 1395 26700
rect 1429 26693 1470 26700
rect 1504 26693 1544 26700
rect 1578 26693 1618 26700
rect 1652 26693 1692 26700
rect 1726 26693 1758 26727
rect 1429 26676 1758 26693
rect 999 26665 1758 26676
rect 999 26631 1057 26665
rect 1091 26631 1125 26665
rect 1159 26631 1193 26665
rect 1227 26631 1261 26665
rect 1295 26631 1329 26665
rect 1363 26636 1397 26665
rect 1363 26631 1395 26636
rect 1431 26631 1465 26665
rect 1499 26655 1533 26665
rect 1567 26655 1601 26665
rect 1635 26655 1669 26665
rect 1703 26655 1758 26665
rect 1504 26631 1533 26655
rect 1578 26631 1601 26655
rect 1652 26631 1669 26655
rect 999 26602 1395 26631
rect 1429 26621 1470 26631
rect 1504 26621 1544 26631
rect 1578 26621 1618 26631
rect 1652 26621 1692 26631
rect 1726 26621 1758 26655
rect 1429 26602 1758 26621
rect 999 26596 1758 26602
rect 999 26562 1057 26596
rect 1091 26562 1125 26596
rect 1159 26562 1193 26596
rect 1227 26562 1261 26596
rect 1295 26562 1329 26596
rect 1363 26562 1397 26596
rect 1431 26562 1465 26596
rect 1499 26583 1533 26596
rect 1567 26583 1601 26596
rect 1635 26583 1669 26596
rect 1703 26583 1758 26596
rect 1504 26562 1533 26583
rect 1578 26562 1601 26583
rect 1652 26562 1669 26583
rect 999 26528 1395 26562
rect 1429 26549 1470 26562
rect 1504 26549 1544 26562
rect 1578 26549 1618 26562
rect 1652 26549 1692 26562
rect 1726 26549 1758 26583
rect 1429 26528 1758 26549
rect 999 26527 1758 26528
rect 999 26493 1057 26527
rect 1091 26493 1125 26527
rect 1159 26493 1193 26527
rect 1227 26493 1261 26527
rect 1295 26493 1329 26527
rect 1363 26493 1397 26527
rect 1431 26493 1465 26527
rect 1499 26511 1533 26527
rect 1567 26511 1601 26527
rect 1635 26511 1669 26527
rect 1703 26511 1758 26527
rect 1504 26493 1533 26511
rect 1578 26493 1601 26511
rect 1652 26493 1669 26511
rect 999 26488 1470 26493
rect 999 26458 1395 26488
rect 1429 26477 1470 26488
rect 1504 26477 1544 26493
rect 1578 26477 1618 26493
rect 1652 26477 1692 26493
rect 1726 26477 1758 26511
rect 1429 26458 1758 26477
rect 999 26424 1057 26458
rect 1091 26424 1125 26458
rect 1159 26424 1193 26458
rect 1227 26424 1261 26458
rect 1295 26424 1329 26458
rect 1363 26454 1395 26458
rect 1363 26424 1397 26454
rect 1431 26424 1465 26458
rect 1499 26439 1533 26458
rect 1567 26439 1601 26458
rect 1635 26439 1669 26458
rect 1703 26439 1758 26458
rect 1504 26424 1533 26439
rect 1578 26424 1601 26439
rect 1652 26424 1669 26439
rect 999 26414 1470 26424
rect 999 26389 1395 26414
rect 1429 26405 1470 26414
rect 1504 26405 1544 26424
rect 1578 26405 1618 26424
rect 1652 26405 1692 26424
rect 1726 26405 1758 26439
rect 1429 26389 1758 26405
rect 999 26355 1057 26389
rect 1091 26355 1125 26389
rect 1159 26355 1193 26389
rect 1227 26355 1261 26389
rect 1295 26355 1329 26389
rect 1363 26380 1395 26389
rect 1363 26355 1397 26380
rect 1431 26355 1465 26389
rect 1499 26367 1533 26389
rect 1567 26367 1601 26389
rect 1635 26367 1669 26389
rect 1703 26367 1758 26389
rect 1504 26355 1533 26367
rect 1578 26355 1601 26367
rect 1652 26355 1669 26367
rect 999 26340 1470 26355
rect 999 26320 1395 26340
rect 1429 26333 1470 26340
rect 1504 26333 1544 26355
rect 1578 26333 1618 26355
rect 1652 26333 1692 26355
rect 1726 26333 1758 26367
rect 1429 26320 1758 26333
rect 999 26286 1057 26320
rect 1091 26286 1125 26320
rect 1159 26286 1193 26320
rect 1227 26286 1261 26320
rect 1295 26286 1329 26320
rect 1363 26306 1395 26320
rect 1363 26286 1397 26306
rect 1431 26286 1465 26320
rect 1499 26295 1533 26320
rect 1567 26295 1601 26320
rect 1635 26295 1669 26320
rect 1703 26295 1758 26320
rect 1504 26286 1533 26295
rect 1578 26286 1601 26295
rect 1652 26286 1669 26295
rect 999 26266 1470 26286
rect 999 26251 1395 26266
rect 1429 26261 1470 26266
rect 1504 26261 1544 26286
rect 1578 26261 1618 26286
rect 1652 26261 1692 26286
rect 1726 26261 1758 26295
rect 1429 26251 1758 26261
rect 999 26217 1057 26251
rect 1091 26217 1125 26251
rect 1159 26217 1193 26251
rect 1227 26217 1261 26251
rect 1295 26217 1329 26251
rect 1363 26232 1395 26251
rect 1363 26217 1397 26232
rect 1431 26217 1465 26251
rect 1499 26223 1533 26251
rect 1567 26223 1601 26251
rect 1635 26223 1669 26251
rect 1703 26223 1758 26251
rect 1504 26217 1533 26223
rect 1578 26217 1601 26223
rect 1652 26217 1669 26223
rect 999 26193 1470 26217
rect 999 26182 1395 26193
rect 1429 26189 1470 26193
rect 1504 26189 1544 26217
rect 1578 26189 1618 26217
rect 1652 26189 1692 26217
rect 1726 26189 1758 26223
rect 1429 26182 1758 26189
rect 999 26148 1057 26182
rect 1091 26148 1125 26182
rect 1159 26148 1193 26182
rect 1227 26148 1261 26182
rect 1295 26148 1329 26182
rect 1363 26159 1395 26182
rect 1363 26148 1397 26159
rect 1431 26148 1465 26182
rect 1499 26151 1533 26182
rect 1567 26151 1601 26182
rect 1635 26151 1669 26182
rect 1703 26151 1758 26182
rect 1504 26148 1533 26151
rect 1578 26148 1601 26151
rect 1652 26148 1669 26151
rect 999 26120 1470 26148
rect 999 26113 1395 26120
rect 1429 26117 1470 26120
rect 1504 26117 1544 26148
rect 1578 26117 1618 26148
rect 1652 26117 1692 26148
rect 1726 26117 1758 26151
rect 1429 26113 1758 26117
rect 999 26079 1057 26113
rect 1091 26079 1125 26113
rect 1159 26079 1193 26113
rect 1227 26079 1261 26113
rect 1295 26079 1329 26113
rect 1363 26086 1395 26113
rect 1363 26079 1397 26086
rect 1431 26079 1465 26113
rect 1499 26079 1533 26113
rect 1567 26079 1601 26113
rect 1635 26079 1669 26113
rect 1703 26079 1758 26113
rect 999 26047 1470 26079
rect 999 26044 1395 26047
rect 1429 26045 1470 26047
rect 1504 26045 1544 26079
rect 1578 26045 1618 26079
rect 1652 26045 1692 26079
rect 1726 26045 1758 26079
rect 1429 26044 1758 26045
rect 999 26010 1057 26044
rect 1091 26010 1125 26044
rect 1159 26010 1193 26044
rect 1227 26010 1261 26044
rect 1295 26010 1329 26044
rect 1363 26013 1395 26044
rect 1363 26010 1397 26013
rect 1431 26010 1465 26044
rect 1499 26010 1533 26044
rect 1567 26010 1601 26044
rect 1635 26010 1669 26044
rect 1703 26010 1758 26044
rect 999 26007 1758 26010
rect 999 25975 1470 26007
rect 1504 25975 1544 26007
rect 1578 25975 1618 26007
rect 1652 25975 1692 26007
rect 999 25941 1057 25975
rect 1091 25941 1125 25975
rect 1159 25941 1193 25975
rect 1227 25941 1261 25975
rect 1295 25941 1329 25975
rect 1363 25974 1397 25975
rect 1363 25941 1395 25974
rect 1431 25941 1465 25975
rect 1504 25973 1533 25975
rect 1578 25973 1601 25975
rect 1652 25973 1669 25975
rect 1726 25973 1758 26007
rect 1499 25941 1533 25973
rect 1567 25941 1601 25973
rect 1635 25941 1669 25973
rect 1703 25941 1758 25973
rect 999 25940 1395 25941
rect 1429 25940 1758 25941
rect 999 25935 1758 25940
rect 999 25906 1470 25935
rect 1504 25906 1544 25935
rect 1578 25906 1618 25935
rect 1652 25906 1692 25935
rect 999 25872 1057 25906
rect 1091 25872 1125 25906
rect 1159 25872 1193 25906
rect 1227 25872 1261 25906
rect 1295 25872 1329 25906
rect 1363 25901 1397 25906
rect 1363 25872 1395 25901
rect 1431 25872 1465 25906
rect 1504 25901 1533 25906
rect 1578 25901 1601 25906
rect 1652 25901 1669 25906
rect 1726 25901 1758 25935
rect 1499 25872 1533 25901
rect 1567 25872 1601 25901
rect 1635 25872 1669 25901
rect 1703 25872 1758 25901
rect 999 25867 1395 25872
rect 1429 25867 1758 25872
rect 999 25863 1758 25867
rect 999 25837 1470 25863
rect 1504 25837 1544 25863
rect 1578 25837 1618 25863
rect 1652 25837 1692 25863
rect 999 25803 1057 25837
rect 1091 25803 1125 25837
rect 1159 25803 1193 25837
rect 1227 25803 1261 25837
rect 1295 25803 1329 25837
rect 1363 25828 1397 25837
rect 1363 25803 1395 25828
rect 1431 25803 1465 25837
rect 1504 25829 1533 25837
rect 1578 25829 1601 25837
rect 1652 25829 1669 25837
rect 1726 25829 1758 25863
rect 1499 25803 1533 25829
rect 1567 25803 1601 25829
rect 1635 25803 1669 25829
rect 1703 25803 1758 25829
rect 999 25794 1395 25803
rect 1429 25794 1758 25803
rect 999 25791 1758 25794
rect 999 25768 1470 25791
rect 1504 25768 1544 25791
rect 1578 25768 1618 25791
rect 1652 25768 1692 25791
rect 999 25734 1057 25768
rect 1091 25734 1125 25768
rect 1159 25734 1193 25768
rect 1227 25734 1261 25768
rect 1295 25734 1329 25768
rect 1363 25755 1397 25768
rect 1363 25734 1395 25755
rect 1431 25734 1465 25768
rect 1504 25757 1533 25768
rect 1578 25757 1601 25768
rect 1652 25757 1669 25768
rect 1726 25757 1758 25791
rect 1499 25734 1533 25757
rect 1567 25734 1601 25757
rect 1635 25734 1669 25757
rect 1703 25734 1758 25757
rect 999 25721 1395 25734
rect 1429 25721 1758 25734
rect 999 25719 1758 25721
rect 999 25699 1470 25719
rect 1504 25699 1544 25719
rect 1578 25699 1618 25719
rect 1652 25699 1692 25719
rect 999 25665 1057 25699
rect 1091 25665 1125 25699
rect 1159 25665 1193 25699
rect 1227 25665 1261 25699
rect 1295 25665 1329 25699
rect 1363 25682 1397 25699
rect 1363 25665 1395 25682
rect 1431 25665 1465 25699
rect 1504 25685 1533 25699
rect 1578 25685 1601 25699
rect 1652 25685 1669 25699
rect 1726 25685 1758 25719
rect 1499 25665 1533 25685
rect 1567 25665 1601 25685
rect 1635 25665 1669 25685
rect 1703 25665 1758 25685
rect 999 25648 1395 25665
rect 1429 25648 1758 25665
rect 999 25647 1758 25648
rect 999 25630 1470 25647
rect 1504 25630 1544 25647
rect 1578 25630 1618 25647
rect 1652 25630 1692 25647
rect 999 25596 1057 25630
rect 1091 25596 1125 25630
rect 1159 25596 1193 25630
rect 1227 25596 1261 25630
rect 1295 25596 1329 25630
rect 1363 25609 1397 25630
rect 1363 25596 1395 25609
rect 1431 25596 1465 25630
rect 1504 25613 1533 25630
rect 1578 25613 1601 25630
rect 1652 25613 1669 25630
rect 1726 25613 1758 25647
rect 1499 25596 1533 25613
rect 1567 25596 1601 25613
rect 1635 25596 1669 25613
rect 1703 25596 1758 25613
rect 999 25575 1395 25596
rect 1429 25575 1758 25596
rect 999 25561 1470 25575
rect 1504 25561 1544 25575
rect 1578 25561 1618 25575
rect 1652 25561 1692 25575
rect 999 25527 1057 25561
rect 1091 25527 1125 25561
rect 1159 25527 1193 25561
rect 1227 25527 1261 25561
rect 1295 25527 1329 25561
rect 1363 25527 1397 25561
rect 1431 25527 1465 25561
rect 1504 25541 1533 25561
rect 1578 25541 1601 25561
rect 1652 25541 1669 25561
rect 1726 25541 1758 25575
rect 1499 25527 1533 25541
rect 1567 25527 1601 25541
rect 1635 25527 1669 25541
rect 1703 25527 1758 25541
rect 999 25502 1758 25527
rect 999 25492 1470 25502
rect 1504 25492 1544 25502
rect 1578 25492 1618 25502
rect 1652 25492 1692 25502
rect 999 25458 1057 25492
rect 1091 25458 1125 25492
rect 1159 25458 1193 25492
rect 1227 25458 1261 25492
rect 1295 25458 1329 25492
rect 1363 25458 1397 25492
rect 1431 25458 1465 25492
rect 1504 25468 1533 25492
rect 1578 25468 1601 25492
rect 1652 25468 1669 25492
rect 1726 25468 1758 25502
rect 1499 25458 1533 25468
rect 1567 25458 1601 25468
rect 1635 25458 1669 25468
rect 1703 25458 1758 25468
rect 999 25429 1758 25458
rect 999 25423 1470 25429
rect 1504 25423 1544 25429
rect 1578 25423 1618 25429
rect 1652 25423 1692 25429
rect 999 25389 1057 25423
rect 1091 25389 1125 25423
rect 1159 25389 1193 25423
rect 1227 25389 1261 25423
rect 1295 25389 1329 25423
rect 1363 25389 1397 25423
rect 1431 25389 1465 25423
rect 1504 25395 1533 25423
rect 1578 25395 1601 25423
rect 1652 25395 1669 25423
rect 1726 25395 1758 25429
rect 1499 25389 1533 25395
rect 1567 25389 1601 25395
rect 1635 25389 1669 25395
rect 1703 25389 1758 25395
rect 999 25356 1758 25389
rect 999 25354 1470 25356
rect 1504 25354 1544 25356
rect 1578 25354 1618 25356
rect 1652 25354 1692 25356
rect 999 25320 1057 25354
rect 1091 25320 1125 25354
rect 1159 25320 1193 25354
rect 1227 25320 1261 25354
rect 1295 25320 1329 25354
rect 1363 25320 1397 25354
rect 1431 25320 1465 25354
rect 1504 25322 1533 25354
rect 1578 25322 1601 25354
rect 1652 25322 1669 25354
rect 1726 25322 1758 25356
rect 1499 25320 1533 25322
rect 1567 25320 1601 25322
rect 1635 25320 1669 25322
rect 1703 25320 1758 25322
rect 999 25285 1758 25320
rect 999 25251 1057 25285
rect 1091 25251 1125 25285
rect 1159 25251 1193 25285
rect 1227 25251 1261 25285
rect 1295 25251 1329 25285
rect 1363 25251 1397 25285
rect 1431 25251 1465 25285
rect 1499 25251 1533 25285
rect 1567 25251 1601 25285
rect 1635 25251 1669 25285
rect 1703 25251 1758 25285
rect 999 25216 1758 25251
rect 999 25182 1057 25216
rect 1091 25209 1125 25216
rect 1159 25209 1193 25216
rect 1227 25209 1261 25216
rect 1295 25209 1329 25216
rect 1363 25209 1397 25216
rect 1431 25209 1465 25216
rect 1093 25182 1125 25209
rect 1167 25182 1193 25209
rect 1241 25182 1261 25209
rect 1315 25182 1329 25209
rect 1389 25182 1397 25209
rect 1463 25182 1465 25209
rect 1499 25209 1533 25216
rect 1567 25209 1601 25216
rect 1635 25209 1669 25216
rect 1499 25182 1503 25209
rect 1567 25182 1577 25209
rect 1635 25182 1651 25209
rect 1703 25182 1758 25216
rect 999 25175 1059 25182
rect 1093 25175 1133 25182
rect 1167 25175 1207 25182
rect 1241 25175 1281 25182
rect 1315 25175 1355 25182
rect 1389 25175 1429 25182
rect 1463 25175 1503 25182
rect 1537 25175 1577 25182
rect 1611 25175 1651 25182
rect 1685 25175 1758 25182
rect 999 25147 1758 25175
rect 999 25113 1057 25147
rect 1091 25134 1125 25147
rect 1159 25134 1193 25147
rect 1227 25134 1261 25147
rect 1295 25134 1329 25147
rect 1363 25134 1397 25147
rect 1431 25134 1465 25147
rect 1093 25113 1125 25134
rect 1167 25113 1193 25134
rect 1241 25113 1261 25134
rect 1315 25113 1329 25134
rect 1389 25113 1397 25134
rect 1463 25113 1465 25134
rect 1499 25134 1533 25147
rect 1567 25134 1601 25147
rect 1635 25134 1669 25147
rect 1499 25113 1503 25134
rect 1567 25113 1577 25134
rect 1635 25113 1651 25134
rect 1703 25113 1758 25147
rect 999 25100 1059 25113
rect 1093 25100 1133 25113
rect 1167 25100 1207 25113
rect 1241 25100 1281 25113
rect 1315 25100 1355 25113
rect 1389 25100 1429 25113
rect 1463 25100 1503 25113
rect 1537 25100 1577 25113
rect 1611 25100 1651 25113
rect 1685 25100 1758 25113
rect 999 25077 1758 25100
rect 999 25043 1057 25077
rect 1091 25059 1125 25077
rect 1159 25059 1193 25077
rect 1227 25059 1261 25077
rect 1295 25059 1329 25077
rect 1363 25059 1397 25077
rect 1431 25059 1465 25077
rect 1093 25043 1125 25059
rect 1167 25043 1193 25059
rect 1241 25043 1261 25059
rect 1315 25043 1329 25059
rect 1389 25043 1397 25059
rect 1463 25043 1465 25059
rect 1499 25059 1533 25077
rect 1567 25059 1601 25077
rect 1635 25059 1669 25077
rect 1499 25043 1503 25059
rect 1567 25043 1577 25059
rect 1635 25043 1651 25059
rect 1703 25043 1758 25077
rect 999 25025 1059 25043
rect 1093 25025 1133 25043
rect 1167 25025 1207 25043
rect 1241 25025 1281 25043
rect 1315 25025 1355 25043
rect 1389 25025 1429 25043
rect 1463 25025 1503 25043
rect 1537 25025 1577 25043
rect 1611 25025 1651 25043
rect 1685 25025 1758 25043
rect 999 25007 1758 25025
rect 999 24973 1057 25007
rect 1091 24984 1125 25007
rect 1159 24984 1193 25007
rect 1227 24984 1261 25007
rect 1295 24984 1329 25007
rect 1363 24984 1397 25007
rect 1431 24984 1465 25007
rect 1093 24973 1125 24984
rect 1167 24973 1193 24984
rect 1241 24973 1261 24984
rect 1315 24973 1329 24984
rect 1389 24973 1397 24984
rect 1463 24973 1465 24984
rect 1499 24984 1533 25007
rect 1567 24984 1601 25007
rect 1635 24984 1669 25007
rect 1499 24973 1503 24984
rect 1567 24973 1577 24984
rect 1635 24973 1651 24984
rect 1703 24973 1758 25007
rect 999 24950 1059 24973
rect 1093 24950 1133 24973
rect 1167 24950 1207 24973
rect 1241 24950 1281 24973
rect 1315 24950 1355 24973
rect 1389 24950 1429 24973
rect 1463 24950 1503 24973
rect 1537 24950 1577 24973
rect 1611 24950 1651 24973
rect 1685 24950 1758 24973
rect 999 24937 1758 24950
rect 999 24903 1057 24937
rect 1091 24909 1125 24937
rect 1159 24909 1193 24937
rect 1227 24909 1261 24937
rect 1295 24909 1329 24937
rect 1363 24909 1397 24937
rect 1431 24909 1465 24937
rect 1093 24903 1125 24909
rect 1167 24903 1193 24909
rect 1241 24903 1261 24909
rect 1315 24903 1329 24909
rect 1389 24903 1397 24909
rect 1463 24903 1465 24909
rect 1499 24909 1533 24937
rect 1567 24909 1601 24937
rect 1635 24909 1669 24937
rect 1499 24903 1503 24909
rect 1567 24903 1577 24909
rect 1635 24903 1651 24909
rect 1703 24903 1758 24937
rect 999 24875 1059 24903
rect 1093 24875 1133 24903
rect 1167 24875 1207 24903
rect 1241 24875 1281 24903
rect 1315 24875 1355 24903
rect 1389 24875 1429 24903
rect 1463 24875 1503 24903
rect 1537 24875 1577 24903
rect 1611 24875 1651 24903
rect 1685 24875 1758 24903
rect 999 24867 1758 24875
rect 999 24833 1057 24867
rect 1091 24834 1125 24867
rect 1159 24834 1193 24867
rect 1227 24834 1261 24867
rect 1295 24834 1329 24867
rect 1363 24834 1397 24867
rect 1431 24834 1465 24867
rect 1093 24833 1125 24834
rect 1167 24833 1193 24834
rect 1241 24833 1261 24834
rect 1315 24833 1329 24834
rect 1389 24833 1397 24834
rect 1463 24833 1465 24834
rect 1499 24834 1533 24867
rect 1567 24834 1601 24867
rect 1635 24834 1669 24867
rect 1499 24833 1503 24834
rect 1567 24833 1577 24834
rect 1635 24833 1651 24834
rect 1703 24833 1758 24867
rect 999 24800 1059 24833
rect 1093 24800 1133 24833
rect 1167 24800 1207 24833
rect 1241 24800 1281 24833
rect 1315 24800 1355 24833
rect 1389 24800 1429 24833
rect 1463 24800 1503 24833
rect 1537 24800 1577 24833
rect 1611 24800 1651 24833
rect 1685 24800 1758 24833
rect 999 24797 1758 24800
rect 999 24763 1057 24797
rect 1091 24763 1125 24797
rect 1159 24763 1193 24797
rect 1227 24763 1261 24797
rect 1295 24763 1329 24797
rect 1363 24763 1397 24797
rect 1431 24763 1465 24797
rect 1499 24763 1533 24797
rect 1567 24763 1601 24797
rect 1635 24763 1669 24797
rect 1703 24763 1758 24797
rect 999 24759 1758 24763
rect 999 24727 1059 24759
rect 1093 24727 1133 24759
rect 1167 24727 1207 24759
rect 1241 24727 1281 24759
rect 1315 24727 1355 24759
rect 1389 24727 1429 24759
rect 1463 24727 1503 24759
rect 1537 24727 1577 24759
rect 1611 24727 1651 24759
rect 1685 24727 1758 24759
rect 999 24693 1057 24727
rect 1093 24725 1125 24727
rect 1167 24725 1193 24727
rect 1241 24725 1261 24727
rect 1315 24725 1329 24727
rect 1389 24725 1397 24727
rect 1463 24725 1465 24727
rect 1091 24693 1125 24725
rect 1159 24693 1193 24725
rect 1227 24693 1261 24725
rect 1295 24693 1329 24725
rect 1363 24693 1397 24725
rect 1431 24693 1465 24725
rect 1499 24725 1503 24727
rect 1567 24725 1577 24727
rect 1635 24725 1651 24727
rect 1499 24693 1533 24725
rect 1567 24693 1601 24725
rect 1635 24693 1669 24725
rect 1703 24693 1758 24727
rect 999 24684 1758 24693
rect 999 24657 1059 24684
rect 1093 24657 1133 24684
rect 1167 24657 1207 24684
rect 1241 24657 1281 24684
rect 1315 24657 1355 24684
rect 1389 24657 1429 24684
rect 1463 24657 1503 24684
rect 1537 24657 1577 24684
rect 1611 24657 1651 24684
rect 1685 24657 1758 24684
rect 999 24623 1057 24657
rect 1093 24650 1125 24657
rect 1167 24650 1193 24657
rect 1241 24650 1261 24657
rect 1315 24650 1329 24657
rect 1389 24650 1397 24657
rect 1463 24650 1465 24657
rect 1091 24623 1125 24650
rect 1159 24623 1193 24650
rect 1227 24623 1261 24650
rect 1295 24623 1329 24650
rect 1363 24623 1397 24650
rect 1431 24623 1465 24650
rect 1499 24650 1503 24657
rect 1567 24650 1577 24657
rect 1635 24650 1651 24657
rect 1499 24623 1533 24650
rect 1567 24623 1601 24650
rect 1635 24623 1669 24650
rect 1703 24623 1758 24657
rect 999 24609 1758 24623
rect 999 24587 1059 24609
rect 1093 24587 1133 24609
rect 1167 24587 1207 24609
rect 1241 24587 1281 24609
rect 1315 24587 1355 24609
rect 1389 24587 1429 24609
rect 1463 24587 1503 24609
rect 1537 24587 1577 24609
rect 1611 24587 1651 24609
rect 1685 24587 1758 24609
rect 999 24553 1057 24587
rect 1093 24575 1125 24587
rect 1167 24575 1193 24587
rect 1241 24575 1261 24587
rect 1315 24575 1329 24587
rect 1389 24575 1397 24587
rect 1463 24575 1465 24587
rect 1091 24553 1125 24575
rect 1159 24553 1193 24575
rect 1227 24553 1261 24575
rect 1295 24553 1329 24575
rect 1363 24553 1397 24575
rect 1431 24553 1465 24575
rect 1499 24575 1503 24587
rect 1567 24575 1577 24587
rect 1635 24575 1651 24587
rect 1499 24553 1533 24575
rect 1567 24553 1601 24575
rect 1635 24553 1669 24575
rect 1703 24553 1758 24587
rect 999 24533 1758 24553
rect 999 24517 1059 24533
rect 1093 24517 1133 24533
rect 1167 24517 1207 24533
rect 1241 24517 1281 24533
rect 1315 24517 1355 24533
rect 1389 24517 1429 24533
rect 1463 24517 1503 24533
rect 1537 24517 1577 24533
rect 1611 24517 1651 24533
rect 1685 24517 1758 24533
rect 999 24483 1057 24517
rect 1093 24499 1125 24517
rect 1167 24499 1193 24517
rect 1241 24499 1261 24517
rect 1315 24499 1329 24517
rect 1389 24499 1397 24517
rect 1463 24499 1465 24517
rect 1091 24483 1125 24499
rect 1159 24483 1193 24499
rect 1227 24483 1261 24499
rect 1295 24483 1329 24499
rect 1363 24483 1397 24499
rect 1431 24483 1465 24499
rect 1499 24499 1503 24517
rect 1567 24499 1577 24517
rect 1635 24499 1651 24517
rect 1499 24483 1533 24499
rect 1567 24483 1601 24499
rect 1635 24483 1669 24499
rect 1703 24483 1758 24517
rect 999 24457 1758 24483
rect 999 24447 1059 24457
rect 1093 24447 1133 24457
rect 1167 24447 1207 24457
rect 1241 24447 1281 24457
rect 1315 24447 1355 24457
rect 1389 24447 1429 24457
rect 1463 24447 1503 24457
rect 1537 24447 1577 24457
rect 1611 24447 1651 24457
rect 1685 24447 1758 24457
rect 999 24413 1057 24447
rect 1093 24423 1125 24447
rect 1167 24423 1193 24447
rect 1241 24423 1261 24447
rect 1315 24423 1329 24447
rect 1389 24423 1397 24447
rect 1463 24423 1465 24447
rect 1091 24413 1125 24423
rect 1159 24413 1193 24423
rect 1227 24413 1261 24423
rect 1295 24413 1329 24423
rect 1363 24413 1397 24423
rect 1431 24413 1465 24423
rect 1499 24423 1503 24447
rect 1567 24423 1577 24447
rect 1635 24423 1651 24447
rect 1499 24413 1533 24423
rect 1567 24413 1601 24423
rect 1635 24413 1669 24423
rect 1703 24413 1758 24447
rect 999 24381 1758 24413
rect 999 24377 1059 24381
rect 1093 24377 1133 24381
rect 1167 24377 1207 24381
rect 1241 24377 1281 24381
rect 1315 24377 1355 24381
rect 1389 24377 1429 24381
rect 1463 24377 1503 24381
rect 1537 24377 1577 24381
rect 1611 24377 1651 24381
rect 1685 24377 1758 24381
rect 999 24343 1057 24377
rect 1093 24347 1125 24377
rect 1167 24347 1193 24377
rect 1241 24347 1261 24377
rect 1315 24347 1329 24377
rect 1389 24347 1397 24377
rect 1463 24347 1465 24377
rect 1091 24343 1125 24347
rect 1159 24343 1193 24347
rect 1227 24343 1261 24347
rect 1295 24343 1329 24347
rect 1363 24343 1397 24347
rect 1431 24343 1465 24347
rect 1499 24347 1503 24377
rect 1567 24347 1577 24377
rect 1635 24347 1651 24377
rect 1499 24343 1533 24347
rect 1567 24343 1601 24347
rect 1635 24343 1669 24347
rect 1703 24343 1758 24377
rect 999 24307 1758 24343
rect 999 24273 1057 24307
rect 1091 24305 1125 24307
rect 1159 24305 1193 24307
rect 1227 24305 1261 24307
rect 1295 24305 1329 24307
rect 1363 24305 1397 24307
rect 1431 24305 1465 24307
rect 1093 24273 1125 24305
rect 1167 24273 1193 24305
rect 1241 24273 1261 24305
rect 1315 24273 1329 24305
rect 1389 24273 1397 24305
rect 1463 24273 1465 24305
rect 1499 24305 1533 24307
rect 1567 24305 1601 24307
rect 1635 24305 1669 24307
rect 1499 24273 1503 24305
rect 1567 24273 1577 24305
rect 1635 24273 1651 24305
rect 1703 24273 1758 24307
rect 999 24271 1059 24273
rect 1093 24271 1133 24273
rect 1167 24271 1207 24273
rect 1241 24271 1281 24273
rect 1315 24271 1355 24273
rect 1389 24271 1429 24273
rect 1463 24271 1503 24273
rect 1537 24271 1577 24273
rect 1611 24271 1651 24273
rect 1685 24271 1758 24273
rect 999 24237 1758 24271
rect 999 24203 1057 24237
rect 1091 24229 1125 24237
rect 1159 24229 1193 24237
rect 1227 24229 1261 24237
rect 1295 24229 1329 24237
rect 1363 24229 1397 24237
rect 1431 24229 1465 24237
rect 1093 24203 1125 24229
rect 1167 24203 1193 24229
rect 1241 24203 1261 24229
rect 1315 24203 1329 24229
rect 1389 24203 1397 24229
rect 1463 24203 1465 24229
rect 1499 24229 1533 24237
rect 1567 24229 1601 24237
rect 1635 24229 1669 24237
rect 1499 24203 1503 24229
rect 1567 24203 1577 24229
rect 1635 24203 1651 24229
rect 1703 24203 1758 24237
rect 999 24195 1059 24203
rect 1093 24195 1133 24203
rect 1167 24195 1207 24203
rect 1241 24195 1281 24203
rect 1315 24195 1355 24203
rect 1389 24195 1429 24203
rect 1463 24195 1503 24203
rect 1537 24195 1577 24203
rect 1611 24195 1651 24203
rect 1685 24195 1758 24203
rect 999 24167 1758 24195
rect 999 24133 1057 24167
rect 1091 24153 1125 24167
rect 1159 24153 1193 24167
rect 1227 24153 1261 24167
rect 1295 24153 1329 24167
rect 1363 24153 1397 24167
rect 1431 24153 1465 24167
rect 1093 24133 1125 24153
rect 1167 24133 1193 24153
rect 1241 24133 1261 24153
rect 1315 24133 1329 24153
rect 1389 24133 1397 24153
rect 1463 24133 1465 24153
rect 1499 24153 1533 24167
rect 1567 24153 1601 24167
rect 1635 24153 1669 24167
rect 1499 24133 1503 24153
rect 1567 24133 1577 24153
rect 1635 24133 1651 24153
rect 1703 24133 1758 24167
rect 999 24119 1059 24133
rect 1093 24119 1133 24133
rect 1167 24119 1207 24133
rect 1241 24119 1281 24133
rect 1315 24119 1355 24133
rect 1389 24119 1429 24133
rect 1463 24119 1503 24133
rect 1537 24119 1577 24133
rect 1611 24119 1651 24133
rect 1685 24119 1758 24133
rect 999 24097 1758 24119
rect 999 24063 1057 24097
rect 1091 24077 1125 24097
rect 1159 24077 1193 24097
rect 1227 24077 1261 24097
rect 1295 24077 1329 24097
rect 1363 24077 1397 24097
rect 1431 24077 1465 24097
rect 1093 24063 1125 24077
rect 1167 24063 1193 24077
rect 1241 24063 1261 24077
rect 1315 24063 1329 24077
rect 1389 24063 1397 24077
rect 1463 24063 1465 24077
rect 1499 24077 1533 24097
rect 1567 24077 1601 24097
rect 1635 24077 1669 24097
rect 1499 24063 1503 24077
rect 1567 24063 1577 24077
rect 1635 24063 1651 24077
rect 1703 24063 1758 24097
rect 999 24043 1059 24063
rect 1093 24043 1133 24063
rect 1167 24043 1207 24063
rect 1241 24043 1281 24063
rect 1315 24043 1355 24063
rect 1389 24043 1429 24063
rect 1463 24043 1503 24063
rect 1537 24043 1577 24063
rect 1611 24043 1651 24063
rect 1685 24043 1758 24063
rect 999 24027 1758 24043
rect 999 23993 1057 24027
rect 1091 24001 1125 24027
rect 1159 24001 1193 24027
rect 1227 24001 1261 24027
rect 1295 24001 1329 24027
rect 1363 24001 1397 24027
rect 1431 24001 1465 24027
rect 1093 23993 1125 24001
rect 1167 23993 1193 24001
rect 1241 23993 1261 24001
rect 1315 23993 1329 24001
rect 1389 23993 1397 24001
rect 1463 23993 1465 24001
rect 1499 24001 1533 24027
rect 1567 24001 1601 24027
rect 1635 24001 1669 24027
rect 1499 23993 1503 24001
rect 1567 23993 1577 24001
rect 1635 23993 1651 24001
rect 1703 23993 1758 24027
rect 999 23967 1059 23993
rect 1093 23967 1133 23993
rect 1167 23967 1207 23993
rect 1241 23967 1281 23993
rect 1315 23967 1355 23993
rect 1389 23967 1429 23993
rect 1463 23967 1503 23993
rect 1537 23967 1577 23993
rect 1611 23967 1651 23993
rect 1685 23967 1758 23993
rect 999 23957 1758 23967
rect 999 23923 1057 23957
rect 1091 23925 1125 23957
rect 1159 23925 1193 23957
rect 1227 23925 1261 23957
rect 1295 23925 1329 23957
rect 1363 23925 1397 23957
rect 1431 23925 1465 23957
rect 1093 23923 1125 23925
rect 1167 23923 1193 23925
rect 1241 23923 1261 23925
rect 1315 23923 1329 23925
rect 1389 23923 1397 23925
rect 1463 23923 1465 23925
rect 1499 23925 1533 23957
rect 1567 23925 1601 23957
rect 1635 23925 1669 23957
rect 1499 23923 1503 23925
rect 1567 23923 1577 23925
rect 1635 23923 1651 23925
rect 1703 23923 1758 23957
rect 999 23891 1059 23923
rect 1093 23891 1133 23923
rect 1167 23891 1207 23923
rect 1241 23891 1281 23923
rect 1315 23891 1355 23923
rect 1389 23891 1429 23923
rect 1463 23891 1503 23923
rect 1537 23891 1577 23923
rect 1611 23891 1651 23923
rect 1685 23891 1758 23923
rect 999 23887 1758 23891
rect 999 23853 1057 23887
rect 1091 23853 1125 23887
rect 1159 23853 1193 23887
rect 1227 23853 1261 23887
rect 1295 23853 1329 23887
rect 1363 23853 1397 23887
rect 1431 23853 1465 23887
rect 1499 23853 1533 23887
rect 1567 23853 1601 23887
rect 1635 23853 1669 23887
rect 1703 23853 1758 23887
rect 999 23849 1758 23853
rect 999 23829 1059 23849
rect 211 23815 1059 23829
rect 1093 23815 1133 23849
rect 1167 23815 1207 23849
rect 1241 23815 1281 23849
rect 1315 23815 1355 23849
rect 1389 23815 1429 23849
rect 1463 23815 1503 23849
rect 1537 23815 1577 23849
rect 1611 23815 1651 23849
rect 1685 23815 1758 23849
rect 211 23753 1758 23815
rect 211 23724 314 23753
rect 348 23724 384 23753
rect 418 23724 454 23753
rect 211 23690 212 23724
rect 246 23690 288 23724
rect 348 23719 364 23724
rect 418 23719 440 23724
rect 488 23719 524 23753
rect 558 23719 594 23753
rect 628 23719 664 23753
rect 698 23719 734 23753
rect 768 23719 804 23753
rect 838 23719 874 23753
rect 908 23719 944 23753
rect 978 23719 1014 23753
rect 1048 23719 1084 23753
rect 1118 23719 1154 23753
rect 1188 23719 1224 23753
rect 1258 23719 1294 23753
rect 1328 23719 1364 23753
rect 1398 23719 1434 23753
rect 1468 23719 1545 23753
rect 1579 23719 1613 23753
rect 1647 23719 1681 23753
rect 1715 23719 1758 23753
rect 322 23690 364 23719
rect 398 23690 440 23719
rect 474 23703 1758 23719
rect 474 23690 513 23703
rect 211 23683 513 23690
rect 547 23683 590 23703
rect 624 23683 667 23703
rect 701 23683 744 23703
rect 778 23683 821 23703
rect 855 23683 898 23703
rect 932 23683 975 23703
rect 1009 23683 1052 23703
rect 1086 23683 1129 23703
rect 1163 23683 1206 23703
rect 1240 23683 1283 23703
rect 1317 23683 1360 23703
rect 1394 23683 1437 23703
rect 211 23652 314 23683
rect 348 23652 384 23683
rect 418 23652 454 23683
rect 488 23669 513 23683
rect 558 23669 590 23683
rect 211 23618 212 23652
rect 246 23618 288 23652
rect 348 23649 364 23652
rect 418 23649 440 23652
rect 488 23649 524 23669
rect 558 23649 594 23669
rect 628 23649 664 23683
rect 701 23669 734 23683
rect 778 23669 804 23683
rect 855 23669 874 23683
rect 932 23669 944 23683
rect 1009 23669 1014 23683
rect 698 23649 734 23669
rect 768 23649 804 23669
rect 838 23649 874 23669
rect 908 23649 944 23669
rect 978 23649 1014 23669
rect 1048 23669 1052 23683
rect 1118 23669 1129 23683
rect 1188 23669 1206 23683
rect 1258 23669 1283 23683
rect 1328 23669 1360 23683
rect 1048 23649 1084 23669
rect 1118 23649 1154 23669
rect 1188 23649 1224 23669
rect 1258 23649 1294 23669
rect 1328 23649 1364 23669
rect 1398 23649 1434 23683
rect 1471 23669 1758 23703
rect 1468 23650 1758 23669
rect 1468 23649 1545 23650
rect 322 23618 364 23649
rect 398 23618 440 23649
rect 474 23623 1545 23649
rect 474 23618 513 23623
rect 211 23613 513 23618
rect 547 23613 590 23623
rect 624 23613 667 23623
rect 701 23613 744 23623
rect 778 23613 821 23623
rect 855 23613 898 23623
rect 932 23613 975 23623
rect 1009 23613 1052 23623
rect 1086 23613 1129 23623
rect 1163 23613 1206 23623
rect 1240 23613 1283 23623
rect 1317 23613 1360 23623
rect 1394 23613 1437 23623
rect 1471 23616 1545 23623
rect 1579 23616 1613 23650
rect 1647 23616 1681 23650
rect 1715 23616 1758 23650
rect 211 23580 314 23613
rect 348 23580 384 23613
rect 418 23580 454 23613
rect 488 23589 513 23613
rect 558 23589 590 23613
rect 211 23546 212 23580
rect 246 23546 288 23580
rect 348 23579 364 23580
rect 418 23579 440 23580
rect 488 23579 524 23589
rect 558 23579 594 23589
rect 628 23579 664 23613
rect 701 23589 734 23613
rect 778 23589 804 23613
rect 855 23589 874 23613
rect 932 23589 944 23613
rect 1009 23589 1014 23613
rect 698 23579 734 23589
rect 768 23579 804 23589
rect 838 23579 874 23589
rect 908 23579 944 23589
rect 978 23579 1014 23589
rect 1048 23589 1052 23613
rect 1118 23589 1129 23613
rect 1188 23589 1206 23613
rect 1258 23589 1283 23613
rect 1328 23589 1360 23613
rect 1048 23579 1084 23589
rect 1118 23579 1154 23589
rect 1188 23579 1224 23589
rect 1258 23579 1294 23589
rect 1328 23579 1364 23589
rect 1398 23579 1434 23613
rect 1471 23592 1758 23616
rect 18021 27102 18022 27136
rect 18056 27119 18108 27136
rect 18142 27119 18194 27136
rect 18228 27119 18280 27136
rect 18314 27119 18366 27136
rect 18021 27085 18025 27102
rect 18059 27085 18101 27119
rect 18142 27102 18177 27119
rect 18228 27102 18253 27119
rect 18314 27102 18329 27119
rect 18135 27085 18177 27102
rect 18211 27085 18253 27102
rect 18287 27085 18329 27102
rect 18363 27102 18366 27119
rect 18400 27135 19012 27136
rect 18400 27119 18486 27135
rect 18400 27102 18405 27119
rect 18363 27085 18405 27102
rect 18439 27101 18486 27119
rect 18520 27101 18556 27135
rect 18590 27101 18626 27135
rect 18660 27101 18696 27135
rect 18730 27101 18766 27135
rect 18800 27101 18836 27135
rect 18870 27101 18906 27135
rect 18940 27101 18976 27135
rect 19010 27101 19012 27135
rect 18439 27085 19012 27101
rect 18021 27067 19012 27085
rect 18021 27064 18486 27067
rect 18021 27030 18022 27064
rect 18056 27051 18108 27064
rect 18142 27051 18194 27064
rect 18228 27051 18280 27064
rect 18314 27051 18366 27064
rect 18021 27017 18025 27030
rect 18059 27017 18101 27051
rect 18142 27030 18177 27051
rect 18228 27030 18253 27051
rect 18314 27030 18329 27051
rect 18135 27017 18177 27030
rect 18211 27017 18253 27030
rect 18287 27017 18329 27030
rect 18363 27030 18366 27051
rect 18400 27051 18486 27064
rect 18400 27030 18405 27051
rect 18363 27017 18405 27030
rect 18439 27033 18486 27051
rect 18520 27033 18556 27067
rect 18590 27033 18626 27067
rect 18660 27033 18696 27067
rect 18730 27033 18766 27067
rect 18800 27033 18836 27067
rect 18870 27033 18906 27067
rect 18940 27033 18976 27067
rect 19010 27033 19012 27067
rect 18439 27017 19012 27033
rect 18021 26999 19012 27017
rect 18021 26992 18486 26999
rect 18021 26958 18022 26992
rect 18056 26983 18108 26992
rect 18142 26983 18194 26992
rect 18228 26983 18280 26992
rect 18314 26983 18366 26992
rect 18021 26949 18025 26958
rect 18059 26949 18101 26983
rect 18142 26958 18177 26983
rect 18228 26958 18253 26983
rect 18314 26958 18329 26983
rect 18135 26949 18177 26958
rect 18211 26949 18253 26958
rect 18287 26949 18329 26958
rect 18363 26958 18366 26983
rect 18400 26983 18486 26992
rect 18400 26958 18405 26983
rect 18363 26949 18405 26958
rect 18439 26965 18486 26983
rect 18520 26965 18556 26999
rect 18590 26965 18626 26999
rect 18660 26965 18696 26999
rect 18730 26965 18766 26999
rect 18800 26965 18836 26999
rect 18870 26965 18906 26999
rect 18940 26965 18976 26999
rect 19010 26965 19012 26999
rect 18439 26949 19012 26965
rect 18021 26931 19012 26949
rect 18021 26920 18486 26931
rect 18021 26886 18022 26920
rect 18056 26915 18108 26920
rect 18142 26915 18194 26920
rect 18228 26915 18280 26920
rect 18314 26915 18366 26920
rect 18021 26881 18025 26886
rect 18059 26881 18101 26915
rect 18142 26886 18177 26915
rect 18228 26886 18253 26915
rect 18314 26886 18329 26915
rect 18135 26881 18177 26886
rect 18211 26881 18253 26886
rect 18287 26881 18329 26886
rect 18363 26886 18366 26915
rect 18400 26915 18486 26920
rect 18400 26886 18405 26915
rect 18363 26881 18405 26886
rect 18439 26897 18486 26915
rect 18520 26897 18556 26931
rect 18590 26897 18626 26931
rect 18660 26897 18696 26931
rect 18730 26897 18766 26931
rect 18800 26897 18836 26931
rect 18870 26897 18906 26931
rect 18940 26897 18976 26931
rect 19010 26897 19012 26931
rect 18439 26881 19012 26897
rect 18021 26863 19012 26881
rect 18021 26848 18486 26863
rect 18021 26814 18022 26848
rect 18056 26847 18108 26848
rect 18142 26847 18194 26848
rect 18228 26847 18280 26848
rect 18314 26847 18366 26848
rect 18021 26813 18025 26814
rect 18059 26813 18101 26847
rect 18142 26814 18177 26847
rect 18228 26814 18253 26847
rect 18314 26814 18329 26847
rect 18135 26813 18177 26814
rect 18211 26813 18253 26814
rect 18287 26813 18329 26814
rect 18363 26814 18366 26847
rect 18400 26847 18486 26848
rect 18400 26814 18405 26847
rect 18363 26813 18405 26814
rect 18439 26829 18486 26847
rect 18520 26829 18556 26863
rect 18590 26829 18626 26863
rect 18660 26829 18696 26863
rect 18730 26829 18766 26863
rect 18800 26829 18836 26863
rect 18870 26829 18906 26863
rect 18940 26829 18976 26863
rect 19010 26829 19012 26863
rect 18439 26813 19012 26829
rect 18021 26795 19012 26813
rect 18021 26779 18486 26795
rect 18021 26776 18025 26779
rect 18021 26742 18022 26776
rect 18059 26745 18101 26779
rect 18135 26776 18177 26779
rect 18211 26776 18253 26779
rect 18287 26776 18329 26779
rect 18142 26745 18177 26776
rect 18228 26745 18253 26776
rect 18314 26745 18329 26776
rect 18363 26776 18405 26779
rect 18363 26745 18366 26776
rect 18056 26742 18108 26745
rect 18142 26742 18194 26745
rect 18228 26742 18280 26745
rect 18314 26742 18366 26745
rect 18400 26745 18405 26776
rect 18439 26761 18486 26779
rect 18520 26761 18556 26795
rect 18590 26761 18626 26795
rect 18660 26761 18696 26795
rect 18730 26761 18766 26795
rect 18800 26761 18836 26795
rect 18870 26761 18906 26795
rect 18940 26761 18976 26795
rect 19010 26761 19012 26795
rect 18439 26745 19012 26761
rect 18400 26742 19012 26745
rect 18021 26727 19012 26742
rect 18021 26711 18486 26727
rect 18021 26704 18025 26711
rect 18021 26670 18022 26704
rect 18059 26677 18101 26711
rect 18135 26704 18177 26711
rect 18211 26704 18253 26711
rect 18287 26704 18329 26711
rect 18142 26677 18177 26704
rect 18228 26677 18253 26704
rect 18314 26677 18329 26704
rect 18363 26704 18405 26711
rect 18363 26677 18366 26704
rect 18056 26670 18108 26677
rect 18142 26670 18194 26677
rect 18228 26670 18280 26677
rect 18314 26670 18366 26677
rect 18400 26677 18405 26704
rect 18439 26693 18486 26711
rect 18520 26693 18556 26727
rect 18590 26693 18626 26727
rect 18660 26693 18696 26727
rect 18730 26693 18766 26727
rect 18800 26693 18836 26727
rect 18870 26693 18906 26727
rect 18940 26693 18976 26727
rect 19010 26693 19012 26727
rect 18439 26677 19012 26693
rect 18400 26670 19012 26677
rect 18021 26659 19012 26670
rect 18021 26643 18486 26659
rect 18021 26632 18025 26643
rect 18021 26598 18022 26632
rect 18059 26609 18101 26643
rect 18135 26632 18177 26643
rect 18211 26632 18253 26643
rect 18287 26632 18329 26643
rect 18142 26609 18177 26632
rect 18228 26609 18253 26632
rect 18314 26609 18329 26632
rect 18363 26632 18405 26643
rect 18363 26609 18366 26632
rect 18056 26598 18108 26609
rect 18142 26598 18194 26609
rect 18228 26598 18280 26609
rect 18314 26598 18366 26609
rect 18400 26609 18405 26632
rect 18439 26625 18486 26643
rect 18520 26625 18556 26659
rect 18590 26625 18626 26659
rect 18660 26625 18696 26659
rect 18730 26625 18766 26659
rect 18800 26625 18836 26659
rect 18870 26625 18906 26659
rect 18940 26625 18976 26659
rect 19010 26625 19012 26659
rect 18439 26609 19012 26625
rect 18400 26598 19012 26609
rect 18021 26591 19012 26598
rect 18021 26575 18486 26591
rect 18021 26560 18025 26575
rect 18021 26526 18022 26560
rect 18059 26541 18101 26575
rect 18135 26560 18177 26575
rect 18211 26560 18253 26575
rect 18287 26560 18329 26575
rect 18142 26541 18177 26560
rect 18228 26541 18253 26560
rect 18314 26541 18329 26560
rect 18363 26560 18405 26575
rect 18363 26541 18366 26560
rect 18056 26526 18108 26541
rect 18142 26526 18194 26541
rect 18228 26526 18280 26541
rect 18314 26526 18366 26541
rect 18400 26541 18405 26560
rect 18439 26557 18486 26575
rect 18520 26557 18556 26591
rect 18590 26557 18626 26591
rect 18660 26557 18696 26591
rect 18730 26557 18766 26591
rect 18800 26557 18836 26591
rect 18870 26557 18906 26591
rect 18940 26557 18976 26591
rect 19010 26557 19012 26591
rect 18439 26541 19012 26557
rect 18400 26526 19012 26541
rect 18021 26523 19012 26526
rect 18021 26507 18486 26523
rect 18021 26488 18025 26507
rect 18021 26454 18022 26488
rect 18059 26473 18101 26507
rect 18135 26488 18177 26507
rect 18211 26488 18253 26507
rect 18287 26488 18329 26507
rect 18142 26473 18177 26488
rect 18228 26473 18253 26488
rect 18314 26473 18329 26488
rect 18363 26488 18405 26507
rect 18363 26473 18366 26488
rect 18056 26454 18108 26473
rect 18142 26454 18194 26473
rect 18228 26454 18280 26473
rect 18314 26454 18366 26473
rect 18400 26473 18405 26488
rect 18439 26489 18486 26507
rect 18520 26489 18556 26523
rect 18590 26489 18626 26523
rect 18660 26489 18696 26523
rect 18730 26489 18766 26523
rect 18800 26489 18836 26523
rect 18870 26489 18906 26523
rect 18940 26489 18976 26523
rect 19010 26489 19012 26523
rect 18439 26473 19012 26489
rect 18400 26455 19012 26473
rect 18400 26454 18486 26455
rect 18021 26439 18486 26454
rect 18021 26416 18025 26439
rect 18021 26382 18022 26416
rect 18059 26405 18101 26439
rect 18135 26416 18177 26439
rect 18211 26416 18253 26439
rect 18287 26416 18329 26439
rect 18142 26405 18177 26416
rect 18228 26405 18253 26416
rect 18314 26405 18329 26416
rect 18363 26416 18405 26439
rect 18363 26405 18366 26416
rect 18056 26382 18108 26405
rect 18142 26382 18194 26405
rect 18228 26382 18280 26405
rect 18314 26382 18366 26405
rect 18400 26405 18405 26416
rect 18439 26421 18486 26439
rect 18520 26421 18556 26455
rect 18590 26421 18626 26455
rect 18660 26421 18696 26455
rect 18730 26421 18766 26455
rect 18800 26421 18836 26455
rect 18870 26421 18906 26455
rect 18940 26421 18976 26455
rect 19010 26421 19012 26455
rect 18439 26405 19012 26421
rect 18400 26387 19012 26405
rect 18400 26382 18486 26387
rect 18021 26371 18486 26382
rect 18021 26344 18025 26371
rect 18021 26310 18022 26344
rect 18059 26337 18101 26371
rect 18135 26344 18177 26371
rect 18211 26344 18253 26371
rect 18287 26344 18329 26371
rect 18142 26337 18177 26344
rect 18228 26337 18253 26344
rect 18314 26337 18329 26344
rect 18363 26344 18405 26371
rect 18363 26337 18366 26344
rect 18056 26310 18108 26337
rect 18142 26310 18194 26337
rect 18228 26310 18280 26337
rect 18314 26310 18366 26337
rect 18400 26337 18405 26344
rect 18439 26353 18486 26371
rect 18520 26353 18556 26387
rect 18590 26353 18626 26387
rect 18660 26353 18696 26387
rect 18730 26353 18766 26387
rect 18800 26353 18836 26387
rect 18870 26353 18906 26387
rect 18940 26353 18976 26387
rect 19010 26353 19012 26387
rect 18439 26337 19012 26353
rect 18400 26319 19012 26337
rect 18400 26310 18486 26319
rect 18021 26303 18486 26310
rect 18021 26272 18025 26303
rect 18021 26238 18022 26272
rect 18059 26269 18101 26303
rect 18135 26272 18177 26303
rect 18211 26272 18253 26303
rect 18287 26272 18329 26303
rect 18142 26269 18177 26272
rect 18228 26269 18253 26272
rect 18314 26269 18329 26272
rect 18363 26272 18405 26303
rect 18363 26269 18366 26272
rect 18056 26238 18108 26269
rect 18142 26238 18194 26269
rect 18228 26238 18280 26269
rect 18314 26238 18366 26269
rect 18400 26269 18405 26272
rect 18439 26285 18486 26303
rect 18520 26285 18556 26319
rect 18590 26285 18626 26319
rect 18660 26285 18696 26319
rect 18730 26285 18766 26319
rect 18800 26285 18836 26319
rect 18870 26285 18906 26319
rect 18940 26285 18976 26319
rect 19010 26285 19012 26319
rect 18439 26269 19012 26285
rect 18400 26251 19012 26269
rect 18400 26238 18486 26251
rect 18021 26235 18486 26238
rect 18021 26201 18025 26235
rect 18059 26201 18101 26235
rect 18135 26201 18177 26235
rect 18211 26201 18253 26235
rect 18287 26201 18329 26235
rect 18363 26201 18405 26235
rect 18439 26217 18486 26235
rect 18520 26217 18556 26251
rect 18590 26217 18626 26251
rect 18660 26217 18696 26251
rect 18730 26217 18766 26251
rect 18800 26217 18836 26251
rect 18870 26217 18906 26251
rect 18940 26217 18976 26251
rect 19010 26217 19012 26251
rect 18439 26201 19012 26217
rect 18021 26200 19012 26201
rect 18021 26166 18022 26200
rect 18056 26167 18108 26200
rect 18142 26167 18194 26200
rect 18228 26167 18280 26200
rect 18314 26167 18366 26200
rect 18021 26133 18025 26166
rect 18059 26133 18101 26167
rect 18142 26166 18177 26167
rect 18228 26166 18253 26167
rect 18314 26166 18329 26167
rect 18135 26133 18177 26166
rect 18211 26133 18253 26166
rect 18287 26133 18329 26166
rect 18363 26166 18366 26167
rect 18400 26183 19012 26200
rect 18400 26167 18486 26183
rect 18400 26166 18405 26167
rect 18363 26133 18405 26166
rect 18439 26149 18486 26167
rect 18520 26149 18556 26183
rect 18590 26149 18626 26183
rect 18660 26149 18696 26183
rect 18730 26149 18766 26183
rect 18800 26149 18836 26183
rect 18870 26149 18906 26183
rect 18940 26149 18976 26183
rect 19010 26149 19012 26183
rect 18439 26133 19012 26149
rect 18021 26128 19012 26133
rect 18021 26094 18022 26128
rect 18056 26099 18108 26128
rect 18142 26099 18194 26128
rect 18228 26099 18280 26128
rect 18314 26099 18366 26128
rect 18021 26065 18025 26094
rect 18059 26065 18101 26099
rect 18142 26094 18177 26099
rect 18228 26094 18253 26099
rect 18314 26094 18329 26099
rect 18135 26065 18177 26094
rect 18211 26065 18253 26094
rect 18287 26065 18329 26094
rect 18363 26094 18366 26099
rect 18400 26115 19012 26128
rect 18400 26099 18486 26115
rect 18400 26094 18405 26099
rect 18363 26065 18405 26094
rect 18439 26081 18486 26099
rect 18520 26081 18556 26115
rect 18590 26081 18626 26115
rect 18660 26081 18696 26115
rect 18730 26081 18766 26115
rect 18800 26081 18836 26115
rect 18870 26081 18906 26115
rect 18940 26081 18976 26115
rect 19010 26081 19012 26115
rect 18439 26065 19012 26081
rect 18021 26056 19012 26065
rect 18021 26022 18022 26056
rect 18056 26031 18108 26056
rect 18142 26031 18194 26056
rect 18228 26031 18280 26056
rect 18314 26031 18366 26056
rect 18021 25997 18025 26022
rect 18059 25997 18101 26031
rect 18142 26022 18177 26031
rect 18228 26022 18253 26031
rect 18314 26022 18329 26031
rect 18135 25997 18177 26022
rect 18211 25997 18253 26022
rect 18287 25997 18329 26022
rect 18363 26022 18366 26031
rect 18400 26047 19012 26056
rect 18400 26031 18486 26047
rect 18400 26022 18405 26031
rect 18363 25997 18405 26022
rect 18439 26013 18486 26031
rect 18520 26013 18556 26047
rect 18590 26013 18626 26047
rect 18660 26013 18696 26047
rect 18730 26013 18766 26047
rect 18800 26013 18836 26047
rect 18870 26013 18906 26047
rect 18940 26013 18976 26047
rect 19010 26013 19012 26047
rect 18439 25997 19012 26013
rect 18021 25984 19012 25997
rect 18021 25950 18022 25984
rect 18056 25963 18108 25984
rect 18142 25963 18194 25984
rect 18228 25963 18280 25984
rect 18314 25963 18366 25984
rect 18021 25929 18025 25950
rect 18059 25929 18101 25963
rect 18142 25950 18177 25963
rect 18228 25950 18253 25963
rect 18314 25950 18329 25963
rect 18135 25929 18177 25950
rect 18211 25929 18253 25950
rect 18287 25929 18329 25950
rect 18363 25950 18366 25963
rect 18400 25979 19012 25984
rect 18400 25963 18486 25979
rect 18400 25950 18405 25963
rect 18363 25929 18405 25950
rect 18439 25945 18486 25963
rect 18520 25945 18556 25979
rect 18590 25945 18626 25979
rect 18660 25945 18696 25979
rect 18730 25945 18766 25979
rect 18800 25945 18836 25979
rect 18870 25945 18906 25979
rect 18940 25945 18976 25979
rect 19010 25945 19012 25979
rect 18439 25929 19012 25945
rect 18021 25912 19012 25929
rect 18021 25878 18022 25912
rect 18056 25895 18108 25912
rect 18142 25895 18194 25912
rect 18228 25895 18280 25912
rect 18314 25895 18366 25912
rect 18021 25861 18025 25878
rect 18059 25861 18101 25895
rect 18142 25878 18177 25895
rect 18228 25878 18253 25895
rect 18314 25878 18329 25895
rect 18135 25861 18177 25878
rect 18211 25861 18253 25878
rect 18287 25861 18329 25878
rect 18363 25878 18366 25895
rect 18400 25911 19012 25912
rect 18400 25895 18486 25911
rect 18400 25878 18405 25895
rect 18363 25861 18405 25878
rect 18439 25877 18486 25895
rect 18520 25877 18556 25911
rect 18590 25877 18626 25911
rect 18660 25877 18696 25911
rect 18730 25877 18766 25911
rect 18800 25877 18836 25911
rect 18870 25877 18906 25911
rect 18940 25877 18976 25911
rect 19010 25877 19012 25911
rect 18439 25861 19012 25877
rect 18021 25843 19012 25861
rect 18021 25840 18486 25843
rect 18021 25806 18022 25840
rect 18056 25827 18108 25840
rect 18142 25827 18194 25840
rect 18228 25827 18280 25840
rect 18314 25827 18366 25840
rect 18021 25793 18025 25806
rect 18059 25793 18101 25827
rect 18142 25806 18177 25827
rect 18228 25806 18253 25827
rect 18314 25806 18329 25827
rect 18135 25793 18177 25806
rect 18211 25793 18253 25806
rect 18287 25793 18329 25806
rect 18363 25806 18366 25827
rect 18400 25827 18486 25840
rect 18400 25806 18405 25827
rect 18363 25793 18405 25806
rect 18439 25809 18486 25827
rect 18520 25809 18556 25843
rect 18590 25809 18626 25843
rect 18660 25809 18696 25843
rect 18730 25809 18766 25843
rect 18800 25809 18836 25843
rect 18870 25809 18906 25843
rect 18940 25809 18976 25843
rect 19010 25809 19012 25843
rect 18439 25793 19012 25809
rect 18021 25775 19012 25793
rect 18021 25768 18486 25775
rect 18021 25734 18022 25768
rect 18056 25759 18108 25768
rect 18142 25759 18194 25768
rect 18228 25759 18280 25768
rect 18314 25759 18366 25768
rect 18021 25725 18025 25734
rect 18059 25725 18101 25759
rect 18142 25734 18177 25759
rect 18228 25734 18253 25759
rect 18314 25734 18329 25759
rect 18135 25725 18177 25734
rect 18211 25725 18253 25734
rect 18287 25725 18329 25734
rect 18363 25734 18366 25759
rect 18400 25759 18486 25768
rect 18400 25734 18405 25759
rect 18363 25725 18405 25734
rect 18439 25741 18486 25759
rect 18520 25741 18556 25775
rect 18590 25741 18626 25775
rect 18660 25741 18696 25775
rect 18730 25741 18766 25775
rect 18800 25741 18836 25775
rect 18870 25741 18906 25775
rect 18940 25741 18976 25775
rect 19010 25741 19012 25775
rect 18439 25725 19012 25741
rect 18021 25707 19012 25725
rect 18021 25696 18486 25707
rect 18021 25662 18022 25696
rect 18056 25691 18108 25696
rect 18142 25691 18194 25696
rect 18228 25691 18280 25696
rect 18314 25691 18366 25696
rect 18021 25657 18025 25662
rect 18059 25657 18101 25691
rect 18142 25662 18177 25691
rect 18228 25662 18253 25691
rect 18314 25662 18329 25691
rect 18135 25657 18177 25662
rect 18211 25657 18253 25662
rect 18287 25657 18329 25662
rect 18363 25662 18366 25691
rect 18400 25691 18486 25696
rect 18400 25662 18405 25691
rect 18363 25657 18405 25662
rect 18439 25673 18486 25691
rect 18520 25673 18556 25707
rect 18590 25673 18626 25707
rect 18660 25673 18696 25707
rect 18730 25673 18766 25707
rect 18800 25673 18836 25707
rect 18870 25673 18906 25707
rect 18940 25673 18976 25707
rect 19010 25673 19012 25707
rect 18439 25657 19012 25673
rect 18021 25638 19012 25657
rect 18021 25624 18486 25638
rect 18021 25590 18022 25624
rect 18056 25623 18108 25624
rect 18142 25623 18194 25624
rect 18228 25623 18280 25624
rect 18314 25623 18366 25624
rect 18021 25589 18025 25590
rect 18059 25589 18101 25623
rect 18142 25590 18177 25623
rect 18228 25590 18253 25623
rect 18314 25590 18329 25623
rect 18135 25589 18177 25590
rect 18211 25589 18253 25590
rect 18287 25589 18329 25590
rect 18363 25590 18366 25623
rect 18400 25623 18486 25624
rect 18400 25590 18405 25623
rect 18363 25589 18405 25590
rect 18439 25604 18486 25623
rect 18520 25604 18556 25638
rect 18590 25604 18626 25638
rect 18660 25604 18696 25638
rect 18730 25604 18766 25638
rect 18800 25604 18836 25638
rect 18870 25604 18906 25638
rect 18940 25604 18976 25638
rect 19010 25604 19012 25638
rect 18439 25589 19012 25604
rect 18021 25569 19012 25589
rect 18021 25555 18486 25569
rect 18021 25552 18025 25555
rect 18021 25518 18022 25552
rect 18059 25521 18101 25555
rect 18135 25552 18177 25555
rect 18211 25552 18253 25555
rect 18287 25552 18329 25555
rect 18142 25521 18177 25552
rect 18228 25521 18253 25552
rect 18314 25521 18329 25552
rect 18363 25552 18405 25555
rect 18363 25521 18366 25552
rect 18056 25518 18108 25521
rect 18142 25518 18194 25521
rect 18228 25518 18280 25521
rect 18314 25518 18366 25521
rect 18400 25521 18405 25552
rect 18439 25535 18486 25555
rect 18520 25535 18556 25569
rect 18590 25535 18626 25569
rect 18660 25535 18696 25569
rect 18730 25535 18766 25569
rect 18800 25535 18836 25569
rect 18870 25535 18906 25569
rect 18940 25535 18976 25569
rect 19010 25535 19012 25569
rect 18439 25521 19012 25535
rect 18400 25518 19012 25521
rect 18021 25500 19012 25518
rect 18021 25487 18486 25500
rect 18021 25480 18025 25487
rect 18021 25446 18022 25480
rect 18059 25453 18101 25487
rect 18135 25480 18177 25487
rect 18211 25480 18253 25487
rect 18287 25480 18329 25487
rect 18142 25453 18177 25480
rect 18228 25453 18253 25480
rect 18314 25453 18329 25480
rect 18363 25480 18405 25487
rect 18363 25453 18366 25480
rect 18056 25446 18108 25453
rect 18142 25446 18194 25453
rect 18228 25446 18280 25453
rect 18314 25446 18366 25453
rect 18400 25453 18405 25480
rect 18439 25466 18486 25487
rect 18520 25466 18556 25500
rect 18590 25466 18626 25500
rect 18660 25466 18696 25500
rect 18730 25466 18766 25500
rect 18800 25466 18836 25500
rect 18870 25466 18906 25500
rect 18940 25466 18976 25500
rect 19010 25466 19012 25500
rect 18439 25453 19012 25466
rect 18400 25446 19012 25453
rect 18021 25431 19012 25446
rect 18021 25419 18486 25431
rect 18021 25408 18025 25419
rect 18021 25374 18022 25408
rect 18059 25385 18101 25419
rect 18135 25408 18177 25419
rect 18211 25408 18253 25419
rect 18287 25408 18329 25419
rect 18142 25385 18177 25408
rect 18228 25385 18253 25408
rect 18314 25385 18329 25408
rect 18363 25408 18405 25419
rect 18363 25385 18366 25408
rect 18056 25374 18108 25385
rect 18142 25374 18194 25385
rect 18228 25374 18280 25385
rect 18314 25374 18366 25385
rect 18400 25385 18405 25408
rect 18439 25397 18486 25419
rect 18520 25397 18556 25431
rect 18590 25397 18626 25431
rect 18660 25397 18696 25431
rect 18730 25397 18766 25431
rect 18800 25397 18836 25431
rect 18870 25397 18906 25431
rect 18940 25397 18976 25431
rect 19010 25397 19012 25431
rect 18439 25385 19012 25397
rect 18400 25374 19012 25385
rect 18021 25362 19012 25374
rect 18021 25351 18486 25362
rect 18021 25336 18025 25351
rect 18021 25302 18022 25336
rect 18059 25317 18101 25351
rect 18135 25336 18177 25351
rect 18211 25336 18253 25351
rect 18287 25336 18329 25351
rect 18142 25317 18177 25336
rect 18228 25317 18253 25336
rect 18314 25317 18329 25336
rect 18363 25336 18405 25351
rect 18363 25317 18366 25336
rect 18056 25302 18108 25317
rect 18142 25302 18194 25317
rect 18228 25302 18280 25317
rect 18314 25302 18366 25317
rect 18400 25317 18405 25336
rect 18439 25328 18486 25351
rect 18520 25328 18556 25362
rect 18590 25328 18626 25362
rect 18660 25328 18696 25362
rect 18730 25328 18766 25362
rect 18800 25328 18836 25362
rect 18870 25328 18906 25362
rect 18940 25328 18976 25362
rect 19010 25328 19012 25362
rect 18439 25317 19012 25328
rect 18400 25302 19012 25317
rect 18021 25293 19012 25302
rect 18021 25283 18486 25293
rect 18021 25264 18025 25283
rect 18021 25230 18022 25264
rect 18059 25249 18101 25283
rect 18135 25264 18177 25283
rect 18211 25264 18253 25283
rect 18287 25264 18329 25283
rect 18142 25249 18177 25264
rect 18228 25249 18253 25264
rect 18314 25249 18329 25264
rect 18363 25264 18405 25283
rect 18363 25249 18366 25264
rect 18056 25230 18108 25249
rect 18142 25230 18194 25249
rect 18228 25230 18280 25249
rect 18314 25230 18366 25249
rect 18400 25249 18405 25264
rect 18439 25259 18486 25283
rect 18520 25259 18556 25293
rect 18590 25259 18626 25293
rect 18660 25259 18696 25293
rect 18730 25259 18766 25293
rect 18800 25259 18836 25293
rect 18870 25259 18906 25293
rect 18940 25259 18976 25293
rect 19010 25259 19012 25293
rect 18439 25249 19012 25259
rect 18400 25230 19012 25249
rect 18021 25224 19012 25230
rect 18021 25214 18486 25224
rect 18021 25192 18025 25214
rect 18021 25158 18022 25192
rect 18059 25180 18101 25214
rect 18135 25192 18177 25214
rect 18211 25192 18253 25214
rect 18287 25192 18329 25214
rect 18142 25180 18177 25192
rect 18228 25180 18253 25192
rect 18314 25180 18329 25192
rect 18363 25192 18405 25214
rect 18363 25180 18366 25192
rect 18056 25158 18108 25180
rect 18142 25158 18194 25180
rect 18228 25158 18280 25180
rect 18314 25158 18366 25180
rect 18400 25180 18405 25192
rect 18439 25190 18486 25214
rect 18520 25190 18556 25224
rect 18590 25190 18626 25224
rect 18660 25190 18696 25224
rect 18730 25190 18766 25224
rect 18800 25190 18836 25224
rect 18870 25190 18906 25224
rect 18940 25190 18976 25224
rect 19010 25190 19012 25224
rect 18439 25180 19012 25190
rect 18400 25158 19012 25180
rect 18021 25155 19012 25158
rect 18021 25145 18486 25155
rect 18021 25120 18025 25145
rect 18021 25086 18022 25120
rect 18059 25111 18101 25145
rect 18135 25120 18177 25145
rect 18211 25120 18253 25145
rect 18287 25120 18329 25145
rect 18142 25111 18177 25120
rect 18228 25111 18253 25120
rect 18314 25111 18329 25120
rect 18363 25120 18405 25145
rect 18363 25111 18366 25120
rect 18056 25086 18108 25111
rect 18142 25086 18194 25111
rect 18228 25086 18280 25111
rect 18314 25086 18366 25111
rect 18400 25111 18405 25120
rect 18439 25121 18486 25145
rect 18520 25121 18556 25155
rect 18590 25121 18626 25155
rect 18660 25121 18696 25155
rect 18730 25121 18766 25155
rect 18800 25121 18836 25155
rect 18870 25121 18906 25155
rect 18940 25121 18976 25155
rect 19010 25121 19012 25155
rect 18439 25111 19012 25121
rect 18400 25086 19012 25111
rect 18021 25076 18486 25086
rect 18021 25048 18025 25076
rect 18021 25014 18022 25048
rect 18059 25042 18101 25076
rect 18135 25048 18177 25076
rect 18211 25048 18253 25076
rect 18287 25048 18329 25076
rect 18142 25042 18177 25048
rect 18228 25042 18253 25048
rect 18314 25042 18329 25048
rect 18363 25048 18405 25076
rect 18363 25042 18366 25048
rect 18056 25014 18108 25042
rect 18142 25014 18194 25042
rect 18228 25014 18280 25042
rect 18314 25014 18366 25042
rect 18400 25042 18405 25048
rect 18439 25052 18486 25076
rect 18520 25052 18556 25086
rect 18590 25052 18626 25086
rect 18660 25052 18696 25086
rect 18730 25052 18766 25086
rect 18800 25052 18836 25086
rect 18870 25052 18906 25086
rect 18940 25052 18976 25086
rect 19010 25052 19012 25086
rect 18439 25042 19012 25052
rect 18400 25017 19012 25042
rect 18400 25014 18486 25017
rect 18021 25007 18486 25014
rect 18021 24976 18025 25007
rect 18021 24942 18022 24976
rect 18059 24973 18101 25007
rect 18135 24976 18177 25007
rect 18211 24976 18253 25007
rect 18287 24976 18329 25007
rect 18142 24973 18177 24976
rect 18228 24973 18253 24976
rect 18314 24973 18329 24976
rect 18363 24976 18405 25007
rect 18363 24973 18366 24976
rect 18056 24942 18108 24973
rect 18142 24942 18194 24973
rect 18228 24942 18280 24973
rect 18314 24942 18366 24973
rect 18400 24973 18405 24976
rect 18439 24983 18486 25007
rect 18520 24983 18556 25017
rect 18590 24983 18626 25017
rect 18660 24983 18696 25017
rect 18730 24983 18766 25017
rect 18800 24983 18836 25017
rect 18870 24983 18906 25017
rect 18940 24983 18976 25017
rect 19010 24983 19012 25017
rect 18439 24973 19012 24983
rect 18400 24948 19012 24973
rect 18400 24942 18486 24948
rect 18021 24938 18486 24942
rect 18021 24904 18025 24938
rect 18059 24904 18101 24938
rect 18135 24904 18177 24938
rect 18211 24904 18253 24938
rect 18287 24904 18329 24938
rect 18363 24904 18405 24938
rect 18439 24914 18486 24938
rect 18520 24914 18556 24948
rect 18590 24914 18626 24948
rect 18660 24914 18696 24948
rect 18730 24914 18766 24948
rect 18800 24914 18836 24948
rect 18870 24914 18906 24948
rect 18940 24914 18976 24948
rect 19010 24914 19012 24948
rect 18439 24904 19012 24914
rect 18021 24870 18022 24904
rect 18056 24870 18108 24904
rect 18142 24870 18194 24904
rect 18228 24870 18280 24904
rect 18314 24870 18366 24904
rect 18400 24879 19012 24904
rect 18400 24870 18486 24879
rect 18021 24869 18486 24870
rect 18021 24835 18025 24869
rect 18059 24835 18101 24869
rect 18135 24835 18177 24869
rect 18211 24835 18253 24869
rect 18287 24835 18329 24869
rect 18363 24835 18405 24869
rect 18439 24845 18486 24869
rect 18520 24845 18556 24879
rect 18590 24845 18626 24879
rect 18660 24845 18696 24879
rect 18730 24845 18766 24879
rect 18800 24845 18836 24879
rect 18870 24845 18906 24879
rect 18940 24845 18976 24879
rect 19010 24845 19012 24879
rect 18439 24835 19012 24845
rect 18021 24832 19012 24835
rect 18021 24798 18022 24832
rect 18056 24800 18108 24832
rect 18142 24800 18194 24832
rect 18228 24800 18280 24832
rect 18314 24800 18366 24832
rect 18021 24766 18025 24798
rect 18059 24766 18101 24800
rect 18142 24798 18177 24800
rect 18228 24798 18253 24800
rect 18314 24798 18329 24800
rect 18135 24766 18177 24798
rect 18211 24766 18253 24798
rect 18287 24766 18329 24798
rect 18363 24798 18366 24800
rect 18400 24810 19012 24832
rect 18400 24800 18486 24810
rect 18400 24798 18405 24800
rect 18363 24766 18405 24798
rect 18439 24776 18486 24800
rect 18520 24776 18556 24810
rect 18590 24776 18626 24810
rect 18660 24776 18696 24810
rect 18730 24776 18766 24810
rect 18800 24776 18836 24810
rect 18870 24776 18906 24810
rect 18940 24776 18976 24810
rect 19010 24776 19012 24810
rect 18439 24766 19012 24776
rect 18021 24760 19012 24766
rect 18021 24726 18022 24760
rect 18056 24731 18108 24760
rect 18142 24731 18194 24760
rect 18228 24731 18280 24760
rect 18314 24731 18366 24760
rect 18021 24697 18025 24726
rect 18059 24697 18101 24731
rect 18142 24726 18177 24731
rect 18228 24726 18253 24731
rect 18314 24726 18329 24731
rect 18135 24697 18177 24726
rect 18211 24697 18253 24726
rect 18287 24697 18329 24726
rect 18363 24726 18366 24731
rect 18400 24741 19012 24760
rect 18400 24731 18486 24741
rect 18400 24726 18405 24731
rect 18363 24697 18405 24726
rect 18439 24707 18486 24731
rect 18520 24707 18556 24741
rect 18590 24707 18626 24741
rect 18660 24707 18696 24741
rect 18730 24707 18766 24741
rect 18800 24707 18836 24741
rect 18870 24707 18906 24741
rect 18940 24707 18976 24741
rect 19010 24707 19012 24741
rect 18439 24697 19012 24707
rect 18021 24688 19012 24697
rect 18021 24654 18022 24688
rect 18056 24662 18108 24688
rect 18142 24662 18194 24688
rect 18228 24662 18280 24688
rect 18314 24662 18366 24688
rect 18021 24628 18025 24654
rect 18059 24628 18101 24662
rect 18142 24654 18177 24662
rect 18228 24654 18253 24662
rect 18314 24654 18329 24662
rect 18135 24628 18177 24654
rect 18211 24628 18253 24654
rect 18287 24628 18329 24654
rect 18363 24654 18366 24662
rect 18400 24672 19012 24688
rect 18400 24662 18486 24672
rect 18400 24654 18405 24662
rect 18363 24628 18405 24654
rect 18439 24638 18486 24662
rect 18520 24638 18556 24672
rect 18590 24638 18626 24672
rect 18660 24638 18696 24672
rect 18730 24638 18766 24672
rect 18800 24638 18836 24672
rect 18870 24638 18906 24672
rect 18940 24638 18976 24672
rect 19010 24638 19012 24672
rect 18439 24628 19012 24638
rect 18021 24616 19012 24628
rect 18021 24582 18022 24616
rect 18056 24593 18108 24616
rect 18142 24593 18194 24616
rect 18228 24593 18280 24616
rect 18314 24593 18366 24616
rect 18021 24559 18025 24582
rect 18059 24559 18101 24593
rect 18142 24582 18177 24593
rect 18228 24582 18253 24593
rect 18314 24582 18329 24593
rect 18135 24559 18177 24582
rect 18211 24559 18253 24582
rect 18287 24559 18329 24582
rect 18363 24582 18366 24593
rect 18400 24603 19012 24616
rect 18400 24593 18486 24603
rect 18400 24582 18405 24593
rect 18363 24559 18405 24582
rect 18439 24569 18486 24593
rect 18520 24569 18556 24603
rect 18590 24569 18626 24603
rect 18660 24569 18696 24603
rect 18730 24569 18766 24603
rect 18800 24569 18836 24603
rect 18870 24569 18906 24603
rect 18940 24569 18976 24603
rect 19010 24569 19012 24603
rect 18439 24559 19012 24569
rect 18021 24544 19012 24559
rect 18021 24510 18022 24544
rect 18056 24524 18108 24544
rect 18142 24524 18194 24544
rect 18228 24524 18280 24544
rect 18314 24524 18366 24544
rect 18021 24490 18025 24510
rect 18059 24490 18101 24524
rect 18142 24510 18177 24524
rect 18228 24510 18253 24524
rect 18314 24510 18329 24524
rect 18135 24490 18177 24510
rect 18211 24490 18253 24510
rect 18287 24490 18329 24510
rect 18363 24510 18366 24524
rect 18400 24534 19012 24544
rect 18400 24524 18486 24534
rect 18400 24510 18405 24524
rect 18363 24490 18405 24510
rect 18439 24500 18486 24524
rect 18520 24500 18556 24534
rect 18590 24500 18626 24534
rect 18660 24500 18696 24534
rect 18730 24500 18766 24534
rect 18800 24500 18836 24534
rect 18870 24500 18906 24534
rect 18940 24500 18976 24534
rect 19010 24500 19012 24534
rect 18439 24490 19012 24500
rect 18021 24472 19012 24490
rect 18021 24438 18022 24472
rect 18056 24455 18108 24472
rect 18142 24455 18194 24472
rect 18228 24455 18280 24472
rect 18314 24455 18366 24472
rect 18021 24421 18025 24438
rect 18059 24421 18101 24455
rect 18142 24438 18177 24455
rect 18228 24438 18253 24455
rect 18314 24438 18329 24455
rect 18135 24421 18177 24438
rect 18211 24421 18253 24438
rect 18287 24421 18329 24438
rect 18363 24438 18366 24455
rect 18400 24465 19012 24472
rect 18400 24455 18486 24465
rect 18400 24438 18405 24455
rect 18363 24421 18405 24438
rect 18439 24431 18486 24455
rect 18520 24431 18556 24465
rect 18590 24431 18626 24465
rect 18660 24431 18696 24465
rect 18730 24431 18766 24465
rect 18800 24431 18836 24465
rect 18870 24431 18906 24465
rect 18940 24431 18976 24465
rect 19010 24431 19012 24465
rect 18439 24421 19012 24431
rect 18021 24400 19012 24421
rect 18021 24366 18022 24400
rect 18056 24386 18108 24400
rect 18142 24386 18194 24400
rect 18228 24386 18280 24400
rect 18314 24386 18366 24400
rect 18021 24352 18025 24366
rect 18059 24352 18101 24386
rect 18142 24366 18177 24386
rect 18228 24366 18253 24386
rect 18314 24366 18329 24386
rect 18135 24352 18177 24366
rect 18211 24352 18253 24366
rect 18287 24352 18329 24366
rect 18363 24366 18366 24386
rect 18400 24396 19012 24400
rect 18400 24386 18486 24396
rect 18400 24366 18405 24386
rect 18363 24352 18405 24366
rect 18439 24362 18486 24386
rect 18520 24362 18556 24396
rect 18590 24362 18626 24396
rect 18660 24362 18696 24396
rect 18730 24362 18766 24396
rect 18800 24362 18836 24396
rect 18870 24362 18906 24396
rect 18940 24362 18976 24396
rect 19010 24362 19012 24396
rect 18439 24352 19012 24362
rect 18021 24328 19012 24352
rect 18021 24294 18022 24328
rect 18056 24317 18108 24328
rect 18142 24317 18194 24328
rect 18228 24317 18280 24328
rect 18314 24317 18366 24328
rect 18021 24283 18025 24294
rect 18059 24283 18101 24317
rect 18142 24294 18177 24317
rect 18228 24294 18253 24317
rect 18314 24294 18329 24317
rect 18135 24283 18177 24294
rect 18211 24283 18253 24294
rect 18287 24283 18329 24294
rect 18363 24294 18366 24317
rect 18400 24327 19012 24328
rect 18400 24317 18486 24327
rect 18400 24294 18405 24317
rect 18363 24283 18405 24294
rect 18439 24293 18486 24317
rect 18520 24293 18556 24327
rect 18590 24293 18626 24327
rect 18660 24293 18696 24327
rect 18730 24293 18766 24327
rect 18800 24293 18836 24327
rect 18870 24293 18906 24327
rect 18940 24293 18976 24327
rect 19010 24293 19012 24327
rect 18439 24283 19012 24293
rect 18021 24258 19012 24283
rect 18021 24256 18486 24258
rect 18021 24222 18022 24256
rect 18056 24248 18108 24256
rect 18142 24248 18194 24256
rect 18228 24248 18280 24256
rect 18314 24248 18366 24256
rect 18021 24214 18025 24222
rect 18059 24214 18101 24248
rect 18142 24222 18177 24248
rect 18228 24222 18253 24248
rect 18314 24222 18329 24248
rect 18135 24214 18177 24222
rect 18211 24214 18253 24222
rect 18287 24214 18329 24222
rect 18363 24222 18366 24248
rect 18400 24248 18486 24256
rect 18400 24222 18405 24248
rect 18363 24214 18405 24222
rect 18439 24224 18486 24248
rect 18520 24224 18556 24258
rect 18590 24224 18626 24258
rect 18660 24224 18696 24258
rect 18730 24224 18766 24258
rect 18800 24224 18836 24258
rect 18870 24224 18906 24258
rect 18940 24224 18976 24258
rect 19010 24224 19012 24258
rect 18439 24214 19012 24224
rect 18021 24189 19012 24214
rect 18021 24184 18486 24189
rect 18021 24150 18022 24184
rect 18056 24179 18108 24184
rect 18142 24179 18194 24184
rect 18228 24179 18280 24184
rect 18314 24179 18366 24184
rect 18021 24145 18025 24150
rect 18059 24145 18101 24179
rect 18142 24150 18177 24179
rect 18228 24150 18253 24179
rect 18314 24150 18329 24179
rect 18135 24145 18177 24150
rect 18211 24145 18253 24150
rect 18287 24145 18329 24150
rect 18363 24150 18366 24179
rect 18400 24179 18486 24184
rect 18400 24150 18405 24179
rect 18363 24145 18405 24150
rect 18439 24155 18486 24179
rect 18520 24155 18556 24189
rect 18590 24155 18626 24189
rect 18660 24155 18696 24189
rect 18730 24155 18766 24189
rect 18800 24155 18836 24189
rect 18870 24155 18906 24189
rect 18940 24155 18976 24189
rect 19010 24155 19012 24189
rect 18439 24145 19012 24155
rect 18021 24120 19012 24145
rect 18021 24112 18486 24120
rect 18021 24078 18022 24112
rect 18056 24110 18108 24112
rect 18142 24110 18194 24112
rect 18228 24110 18280 24112
rect 18314 24110 18366 24112
rect 18021 24076 18025 24078
rect 18059 24076 18101 24110
rect 18142 24078 18177 24110
rect 18228 24078 18253 24110
rect 18314 24078 18329 24110
rect 18135 24076 18177 24078
rect 18211 24076 18253 24078
rect 18287 24076 18329 24078
rect 18363 24078 18366 24110
rect 18400 24110 18486 24112
rect 18400 24078 18405 24110
rect 18363 24076 18405 24078
rect 18439 24086 18486 24110
rect 18520 24086 18556 24120
rect 18590 24086 18626 24120
rect 18660 24086 18696 24120
rect 18730 24086 18766 24120
rect 18800 24086 18836 24120
rect 18870 24086 18906 24120
rect 18940 24086 18976 24120
rect 19010 24086 19012 24120
rect 18439 24076 19012 24086
rect 18021 24051 19012 24076
rect 18021 24041 18486 24051
rect 18021 24040 18025 24041
rect 18021 24006 18022 24040
rect 18059 24007 18101 24041
rect 18135 24040 18177 24041
rect 18211 24040 18253 24041
rect 18287 24040 18329 24041
rect 18142 24007 18177 24040
rect 18228 24007 18253 24040
rect 18314 24007 18329 24040
rect 18363 24040 18405 24041
rect 18363 24007 18366 24040
rect 18056 24006 18108 24007
rect 18142 24006 18194 24007
rect 18228 24006 18280 24007
rect 18314 24006 18366 24007
rect 18400 24007 18405 24040
rect 18439 24017 18486 24041
rect 18520 24017 18556 24051
rect 18590 24017 18626 24051
rect 18660 24017 18696 24051
rect 18730 24017 18766 24051
rect 18800 24017 18836 24051
rect 18870 24017 18906 24051
rect 18940 24017 18976 24051
rect 19010 24017 19012 24051
rect 18439 24007 19012 24017
rect 18400 24006 19012 24007
rect 18021 23982 19012 24006
rect 18021 23972 18486 23982
rect 18021 23968 18025 23972
rect 18021 23934 18022 23968
rect 18059 23938 18101 23972
rect 18135 23968 18177 23972
rect 18211 23968 18253 23972
rect 18287 23968 18329 23972
rect 18142 23938 18177 23968
rect 18228 23938 18253 23968
rect 18314 23938 18329 23968
rect 18363 23968 18405 23972
rect 18363 23938 18366 23968
rect 18056 23934 18108 23938
rect 18142 23934 18194 23938
rect 18228 23934 18280 23938
rect 18314 23934 18366 23938
rect 18400 23938 18405 23968
rect 18439 23948 18486 23972
rect 18520 23948 18556 23982
rect 18590 23948 18626 23982
rect 18660 23948 18696 23982
rect 18730 23948 18766 23982
rect 18800 23948 18836 23982
rect 18870 23948 18906 23982
rect 18940 23948 18976 23982
rect 19010 23948 19012 23982
rect 18439 23938 19012 23948
rect 18400 23934 19012 23938
rect 18021 23913 19012 23934
rect 18021 23903 18486 23913
rect 18021 23896 18025 23903
rect 18021 23862 18022 23896
rect 18059 23869 18101 23903
rect 18135 23896 18177 23903
rect 18211 23896 18253 23903
rect 18287 23896 18329 23903
rect 18142 23869 18177 23896
rect 18228 23869 18253 23896
rect 18314 23869 18329 23896
rect 18363 23896 18405 23903
rect 18363 23869 18366 23896
rect 18056 23862 18108 23869
rect 18142 23862 18194 23869
rect 18228 23862 18280 23869
rect 18314 23862 18366 23869
rect 18400 23869 18405 23896
rect 18439 23879 18486 23903
rect 18520 23879 18556 23913
rect 18590 23879 18626 23913
rect 18660 23879 18696 23913
rect 18730 23879 18766 23913
rect 18800 23879 18836 23913
rect 18870 23879 18906 23913
rect 18940 23879 18976 23913
rect 19010 23879 19012 23913
rect 18439 23869 19012 23879
rect 18400 23862 19012 23869
rect 18021 23844 19012 23862
rect 18021 23834 18486 23844
rect 18021 23824 18025 23834
rect 18021 23790 18022 23824
rect 18059 23800 18101 23834
rect 18135 23824 18177 23834
rect 18211 23824 18253 23834
rect 18287 23824 18329 23834
rect 18142 23800 18177 23824
rect 18228 23800 18253 23824
rect 18314 23800 18329 23824
rect 18363 23824 18405 23834
rect 18363 23800 18366 23824
rect 18056 23790 18108 23800
rect 18142 23790 18194 23800
rect 18228 23790 18280 23800
rect 18314 23790 18366 23800
rect 18400 23800 18405 23824
rect 18439 23810 18486 23834
rect 18520 23810 18556 23844
rect 18590 23810 18626 23844
rect 18660 23810 18696 23844
rect 18730 23810 18766 23844
rect 18800 23810 18836 23844
rect 18870 23810 18906 23844
rect 18940 23810 18976 23844
rect 19010 23810 19012 23844
rect 18439 23800 19012 23810
rect 18400 23790 19012 23800
rect 18021 23775 19012 23790
rect 18021 23765 18486 23775
rect 18021 23752 18025 23765
rect 18021 23718 18022 23752
rect 18059 23731 18101 23765
rect 18135 23752 18177 23765
rect 18211 23752 18253 23765
rect 18287 23752 18329 23765
rect 18142 23731 18177 23752
rect 18228 23731 18253 23752
rect 18314 23731 18329 23752
rect 18363 23752 18405 23765
rect 18363 23731 18366 23752
rect 18056 23718 18108 23731
rect 18142 23718 18194 23731
rect 18228 23718 18280 23731
rect 18314 23718 18366 23731
rect 18400 23731 18405 23752
rect 18439 23741 18486 23765
rect 18520 23741 18556 23775
rect 18590 23741 18626 23775
rect 18660 23741 18696 23775
rect 18730 23741 18766 23775
rect 18800 23741 18836 23775
rect 18870 23741 18906 23775
rect 18940 23741 18976 23775
rect 19010 23741 19012 23775
rect 18439 23731 19012 23741
rect 18400 23718 19012 23731
rect 18021 23706 19012 23718
rect 18021 23696 18486 23706
rect 18021 23680 18025 23696
rect 18021 23646 18022 23680
rect 18059 23662 18101 23696
rect 18135 23680 18177 23696
rect 18211 23680 18253 23696
rect 18287 23680 18329 23696
rect 18142 23662 18177 23680
rect 18228 23662 18253 23680
rect 18314 23662 18329 23680
rect 18363 23680 18405 23696
rect 18363 23662 18366 23680
rect 18056 23646 18108 23662
rect 18142 23646 18194 23662
rect 18228 23646 18280 23662
rect 18314 23646 18366 23662
rect 18400 23662 18405 23680
rect 18439 23672 18486 23696
rect 18520 23672 18556 23706
rect 18590 23672 18626 23706
rect 18660 23672 18696 23706
rect 18730 23672 18766 23706
rect 18800 23672 18836 23706
rect 18870 23672 18906 23706
rect 18940 23672 18976 23706
rect 19010 23672 19012 23706
rect 18439 23662 19012 23672
rect 18400 23646 19012 23662
rect 18021 23637 19012 23646
rect 18021 23627 18486 23637
rect 18021 23607 18025 23627
rect 1471 23589 1503 23592
rect 1468 23579 1503 23589
rect 322 23546 364 23579
rect 398 23546 440 23579
rect 474 23546 1503 23579
rect 211 23543 1503 23546
rect 211 23509 314 23543
rect 348 23509 384 23543
rect 418 23509 454 23543
rect 488 23509 513 23543
rect 558 23509 590 23543
rect 628 23509 664 23543
rect 701 23509 734 23543
rect 778 23509 804 23543
rect 855 23509 874 23543
rect 932 23509 944 23543
rect 1009 23509 1014 23543
rect 1048 23509 1052 23543
rect 1118 23509 1129 23543
rect 1188 23509 1206 23543
rect 1258 23509 1283 23543
rect 1328 23509 1360 23543
rect 1398 23509 1434 23543
rect 1471 23509 1503 23543
rect 211 23508 1503 23509
rect 211 23474 212 23508
rect 246 23474 288 23508
rect 322 23474 364 23508
rect 398 23474 440 23508
rect 474 23474 1503 23508
rect 18021 23573 18022 23607
rect 18059 23593 18101 23627
rect 18135 23607 18177 23627
rect 18211 23607 18253 23627
rect 18287 23607 18329 23627
rect 18142 23593 18177 23607
rect 18228 23593 18253 23607
rect 18314 23593 18329 23607
rect 18363 23607 18405 23627
rect 18363 23593 18366 23607
rect 18056 23573 18108 23593
rect 18142 23573 18194 23593
rect 18228 23573 18280 23593
rect 18314 23573 18366 23593
rect 18400 23593 18405 23607
rect 18439 23603 18486 23627
rect 18520 23603 18556 23637
rect 18590 23603 18626 23637
rect 18660 23603 18696 23637
rect 18730 23603 18766 23637
rect 18800 23603 18836 23637
rect 18870 23603 18906 23637
rect 18940 23603 18976 23637
rect 19010 23603 19012 23637
rect 18439 23593 19012 23603
rect 18400 23573 19012 23593
rect 18021 23568 19012 23573
rect 18021 23558 18486 23568
rect 18021 23534 18025 23558
rect 18021 23500 18022 23534
rect 18059 23524 18101 23558
rect 18135 23534 18177 23558
rect 18211 23534 18253 23558
rect 18287 23534 18329 23558
rect 18142 23524 18177 23534
rect 18228 23524 18253 23534
rect 18314 23524 18329 23534
rect 18363 23534 18405 23558
rect 18363 23524 18366 23534
rect 18056 23500 18108 23524
rect 18142 23500 18194 23524
rect 18228 23500 18280 23524
rect 18314 23500 18366 23524
rect 18400 23524 18405 23534
rect 18439 23534 18486 23558
rect 18520 23534 18556 23568
rect 18590 23534 18626 23568
rect 18660 23534 18696 23568
rect 18730 23534 18766 23568
rect 18800 23534 18836 23568
rect 18870 23534 18906 23568
rect 18940 23534 18976 23568
rect 19010 23534 19012 23568
rect 18439 23524 19012 23534
rect 18400 23500 19012 23524
rect 22823 30683 22827 30717
rect 22864 30712 22897 30717
rect 22861 30683 22897 30712
rect 22931 30712 22932 30717
rect 22966 30717 23034 30746
rect 23068 30717 23635 30746
rect 22966 30712 22967 30717
rect 22931 30683 22967 30712
rect 23001 30712 23034 30717
rect 23001 30683 23037 30712
rect 23071 30683 23107 30717
rect 23141 30683 23177 30717
rect 23211 30683 23247 30717
rect 23281 30683 23317 30717
rect 23351 30683 23387 30717
rect 23421 30683 23457 30717
rect 23491 30683 23527 30717
rect 23561 30683 23597 30717
rect 23631 30683 23635 30717
rect 22823 30671 23635 30683
rect 22823 30649 22830 30671
rect 22864 30649 22932 30671
rect 22823 30615 22827 30649
rect 22864 30637 22897 30649
rect 22861 30615 22897 30637
rect 22931 30637 22932 30649
rect 22966 30649 23034 30671
rect 23068 30649 23635 30671
rect 22966 30637 22967 30649
rect 22931 30615 22967 30637
rect 23001 30637 23034 30649
rect 23001 30615 23037 30637
rect 23071 30615 23107 30649
rect 23141 30615 23177 30649
rect 23211 30615 23247 30649
rect 23281 30615 23317 30649
rect 23351 30615 23387 30649
rect 23421 30615 23457 30649
rect 23491 30615 23527 30649
rect 23561 30615 23597 30649
rect 23631 30615 23635 30649
rect 22823 30596 23635 30615
rect 22823 30581 22830 30596
rect 22864 30581 22932 30596
rect 22823 30547 22827 30581
rect 22864 30562 22897 30581
rect 22861 30547 22897 30562
rect 22931 30562 22932 30581
rect 22966 30581 23034 30596
rect 23068 30581 23635 30596
rect 22966 30562 22967 30581
rect 22931 30547 22967 30562
rect 23001 30562 23034 30581
rect 23001 30547 23037 30562
rect 23071 30547 23107 30581
rect 23141 30547 23177 30581
rect 23211 30547 23247 30581
rect 23281 30547 23317 30581
rect 23351 30547 23387 30581
rect 23421 30547 23457 30581
rect 23491 30547 23527 30581
rect 23561 30547 23597 30581
rect 23631 30547 23635 30581
rect 22823 30521 23635 30547
rect 22823 30513 22830 30521
rect 22864 30513 22932 30521
rect 22823 30479 22827 30513
rect 22864 30487 22897 30513
rect 22861 30479 22897 30487
rect 22931 30487 22932 30513
rect 22966 30513 23034 30521
rect 23068 30513 23635 30521
rect 22966 30487 22967 30513
rect 22931 30479 22967 30487
rect 23001 30487 23034 30513
rect 23001 30479 23037 30487
rect 23071 30479 23107 30513
rect 23141 30479 23177 30513
rect 23211 30479 23247 30513
rect 23281 30479 23317 30513
rect 23351 30479 23387 30513
rect 23421 30479 23457 30513
rect 23491 30479 23527 30513
rect 23561 30479 23597 30513
rect 23631 30479 23635 30513
rect 22823 30446 23635 30479
rect 22823 30445 22830 30446
rect 22864 30445 22932 30446
rect 22823 30411 22827 30445
rect 22864 30412 22897 30445
rect 22861 30411 22897 30412
rect 22931 30412 22932 30445
rect 22966 30445 23034 30446
rect 23068 30445 23635 30446
rect 22966 30412 22967 30445
rect 22931 30411 22967 30412
rect 23001 30412 23034 30445
rect 23001 30411 23037 30412
rect 23071 30411 23107 30445
rect 23141 30411 23177 30445
rect 23211 30411 23247 30445
rect 23281 30411 23317 30445
rect 23351 30411 23387 30445
rect 23421 30411 23457 30445
rect 23491 30411 23527 30445
rect 23561 30411 23597 30445
rect 23631 30411 23635 30445
rect 22823 30377 23635 30411
rect 22823 30343 22827 30377
rect 22861 30371 22897 30377
rect 22864 30343 22897 30371
rect 22931 30371 22967 30377
rect 22931 30343 22932 30371
rect 22823 30337 22830 30343
rect 22864 30337 22932 30343
rect 22966 30343 22967 30371
rect 23001 30371 23037 30377
rect 23001 30343 23034 30371
rect 23071 30343 23107 30377
rect 23141 30343 23177 30377
rect 23211 30343 23247 30377
rect 23281 30343 23317 30377
rect 23351 30343 23387 30377
rect 23421 30343 23457 30377
rect 23491 30343 23527 30377
rect 23561 30343 23597 30377
rect 23631 30343 23635 30377
rect 22966 30337 23034 30343
rect 23068 30337 23635 30343
rect 22823 30309 23635 30337
rect 22823 30275 22827 30309
rect 22861 30296 22897 30309
rect 22864 30275 22897 30296
rect 22931 30296 22967 30309
rect 22931 30275 22932 30296
rect 22823 30262 22830 30275
rect 22864 30262 22932 30275
rect 22966 30275 22967 30296
rect 23001 30296 23037 30309
rect 23001 30275 23034 30296
rect 23071 30275 23107 30309
rect 23141 30275 23177 30309
rect 23211 30275 23247 30309
rect 23281 30275 23317 30309
rect 23351 30275 23387 30309
rect 23421 30275 23457 30309
rect 23491 30275 23527 30309
rect 23561 30275 23597 30309
rect 23631 30275 23635 30309
rect 22966 30262 23034 30275
rect 23068 30262 23635 30275
rect 22823 30241 23635 30262
rect 22823 30207 22827 30241
rect 22861 30221 22897 30241
rect 22864 30207 22897 30221
rect 22931 30221 22967 30241
rect 22931 30207 22932 30221
rect 22823 30187 22830 30207
rect 22864 30187 22932 30207
rect 22966 30207 22967 30221
rect 23001 30221 23037 30241
rect 23001 30207 23034 30221
rect 23071 30207 23107 30241
rect 23141 30207 23177 30241
rect 23211 30207 23247 30241
rect 23281 30207 23317 30241
rect 23351 30207 23387 30241
rect 23421 30207 23457 30241
rect 23491 30207 23527 30241
rect 23561 30207 23597 30241
rect 23631 30207 23635 30241
rect 22966 30187 23034 30207
rect 23068 30187 23635 30207
rect 22823 30173 23635 30187
rect 22823 30139 22827 30173
rect 22861 30146 22897 30173
rect 22864 30139 22897 30146
rect 22931 30146 22967 30173
rect 22931 30139 22932 30146
rect 22823 30112 22830 30139
rect 22864 30112 22932 30139
rect 22966 30139 22967 30146
rect 23001 30146 23037 30173
rect 23001 30139 23034 30146
rect 23071 30139 23107 30173
rect 23141 30139 23177 30173
rect 23211 30139 23247 30173
rect 23281 30139 23317 30173
rect 23351 30139 23387 30173
rect 23421 30139 23457 30173
rect 23491 30139 23527 30173
rect 23561 30139 23597 30173
rect 23631 30139 23635 30173
rect 22966 30112 23034 30139
rect 23068 30112 23635 30139
rect 22823 30105 23635 30112
rect 22823 30071 22827 30105
rect 22861 30071 22897 30105
rect 22931 30071 22967 30105
rect 23001 30071 23037 30105
rect 23071 30071 23107 30105
rect 23141 30071 23177 30105
rect 23211 30071 23247 30105
rect 23281 30071 23317 30105
rect 23351 30071 23387 30105
rect 23421 30071 23457 30105
rect 23491 30071 23527 30105
rect 23561 30071 23597 30105
rect 23631 30071 23635 30105
rect 22823 30037 22830 30071
rect 22864 30037 22932 30071
rect 22966 30037 23034 30071
rect 23068 30037 23635 30071
rect 22823 30003 22827 30037
rect 22861 30003 22897 30037
rect 22931 30003 22967 30037
rect 23001 30003 23037 30037
rect 23071 30003 23107 30037
rect 23141 30003 23177 30037
rect 23211 30003 23247 30037
rect 23281 30003 23317 30037
rect 23351 30003 23387 30037
rect 23421 30003 23457 30037
rect 23491 30003 23527 30037
rect 23561 30003 23597 30037
rect 23631 30003 23635 30037
rect 22823 29996 23635 30003
rect 22823 29969 22830 29996
rect 22864 29969 22932 29996
rect 22823 29935 22827 29969
rect 22864 29962 22897 29969
rect 22861 29935 22897 29962
rect 22931 29962 22932 29969
rect 22966 29969 23034 29996
rect 23068 29969 23635 29996
rect 22966 29962 22967 29969
rect 22931 29935 22967 29962
rect 23001 29962 23034 29969
rect 23001 29935 23037 29962
rect 23071 29935 23107 29969
rect 23141 29935 23177 29969
rect 23211 29935 23247 29969
rect 23281 29935 23317 29969
rect 23351 29935 23387 29969
rect 23421 29935 23457 29969
rect 23491 29935 23527 29969
rect 23561 29935 23597 29969
rect 23631 29935 23635 29969
rect 22823 29921 23635 29935
rect 22823 29901 22830 29921
rect 22864 29901 22932 29921
rect 22823 29867 22827 29901
rect 22864 29887 22897 29901
rect 22861 29867 22897 29887
rect 22931 29887 22932 29901
rect 22966 29901 23034 29921
rect 23068 29901 23635 29921
rect 22966 29887 22967 29901
rect 22931 29867 22967 29887
rect 23001 29887 23034 29901
rect 23001 29867 23037 29887
rect 23071 29867 23107 29901
rect 23141 29867 23177 29901
rect 23211 29867 23247 29901
rect 23281 29867 23317 29901
rect 23351 29867 23387 29901
rect 23421 29867 23457 29901
rect 23491 29867 23527 29901
rect 23561 29867 23597 29901
rect 23631 29867 23635 29901
rect 22823 29846 23635 29867
rect 22823 29833 22830 29846
rect 22864 29833 22932 29846
rect 22823 29799 22827 29833
rect 22864 29812 22897 29833
rect 22861 29799 22897 29812
rect 22931 29812 22932 29833
rect 22966 29833 23034 29846
rect 23068 29833 23635 29846
rect 22966 29812 22967 29833
rect 22931 29799 22967 29812
rect 23001 29812 23034 29833
rect 23001 29799 23037 29812
rect 23071 29799 23107 29833
rect 23141 29799 23177 29833
rect 23211 29799 23247 29833
rect 23281 29799 23317 29833
rect 23351 29799 23387 29833
rect 23421 29799 23457 29833
rect 23491 29799 23527 29833
rect 23561 29799 23597 29833
rect 23631 29799 23635 29833
rect 22823 29771 23635 29799
rect 22823 29765 22830 29771
rect 22864 29765 22932 29771
rect 22823 29731 22827 29765
rect 22864 29737 22897 29765
rect 22861 29731 22897 29737
rect 22931 29737 22932 29765
rect 22966 29765 23034 29771
rect 23068 29765 23635 29771
rect 22966 29737 22967 29765
rect 22931 29731 22967 29737
rect 23001 29737 23034 29765
rect 23001 29731 23037 29737
rect 23071 29731 23107 29765
rect 23141 29731 23177 29765
rect 23211 29731 23247 29765
rect 23281 29731 23317 29765
rect 23351 29731 23387 29765
rect 23421 29731 23457 29765
rect 23491 29731 23527 29765
rect 23561 29731 23597 29765
rect 23631 29731 23635 29765
rect 22823 29697 23635 29731
rect 22823 29663 22827 29697
rect 22861 29693 22897 29697
rect 22876 29663 22897 29693
rect 22931 29663 22967 29697
rect 23001 29663 23037 29697
rect 23071 29663 23107 29697
rect 23141 29663 23177 29697
rect 23211 29663 23247 29697
rect 23281 29663 23317 29697
rect 23351 29663 23387 29697
rect 23421 29663 23457 29697
rect 23491 29663 23527 29697
rect 23561 29663 23597 29697
rect 23631 29663 23635 29697
rect 22823 29659 22842 29663
rect 22876 29659 23635 29663
rect 22823 29629 23635 29659
rect 22823 29595 22827 29629
rect 22861 29621 22897 29629
rect 22876 29595 22897 29621
rect 22931 29595 22967 29629
rect 23001 29595 23037 29629
rect 23071 29595 23107 29629
rect 23141 29595 23177 29629
rect 23211 29595 23247 29629
rect 23281 29595 23317 29629
rect 23351 29595 23387 29629
rect 23421 29595 23457 29629
rect 23491 29595 23527 29629
rect 23561 29595 23597 29629
rect 23631 29595 23635 29629
rect 22823 29587 22842 29595
rect 22876 29587 23635 29595
rect 22823 29561 23635 29587
rect 22823 29527 22827 29561
rect 22861 29549 22897 29561
rect 22876 29527 22897 29549
rect 22931 29527 22967 29561
rect 23001 29527 23037 29561
rect 23071 29527 23107 29561
rect 23141 29527 23177 29561
rect 23211 29527 23247 29561
rect 23281 29527 23317 29561
rect 23351 29527 23387 29561
rect 23421 29527 23457 29561
rect 23491 29527 23527 29561
rect 23561 29527 23597 29561
rect 23631 29527 23635 29561
rect 22823 29515 22842 29527
rect 22876 29515 23635 29527
rect 22823 29493 23635 29515
rect 22823 29459 22827 29493
rect 22861 29477 22897 29493
rect 22876 29459 22897 29477
rect 22931 29459 22967 29493
rect 23001 29459 23037 29493
rect 23071 29459 23107 29493
rect 23141 29459 23177 29493
rect 23211 29459 23247 29493
rect 23281 29459 23317 29493
rect 23351 29459 23387 29493
rect 23421 29459 23457 29493
rect 23491 29459 23527 29493
rect 23561 29459 23597 29493
rect 23631 29459 23635 29493
rect 22823 29443 22842 29459
rect 22876 29443 23635 29459
rect 22823 29425 23635 29443
rect 22823 29391 22827 29425
rect 22861 29405 22897 29425
rect 22876 29391 22897 29405
rect 22931 29391 22967 29425
rect 23001 29391 23037 29425
rect 23071 29391 23107 29425
rect 23141 29391 23177 29425
rect 23211 29391 23247 29425
rect 23281 29391 23317 29425
rect 23351 29391 23387 29425
rect 23421 29391 23457 29425
rect 23491 29391 23527 29425
rect 23561 29391 23597 29425
rect 23631 29391 23635 29425
rect 22823 29371 22842 29391
rect 22876 29371 23635 29391
rect 22823 29357 23635 29371
rect 22823 29323 22827 29357
rect 22861 29333 22897 29357
rect 22876 29323 22897 29333
rect 22931 29323 22967 29357
rect 23001 29323 23037 29357
rect 23071 29323 23107 29357
rect 23141 29323 23177 29357
rect 23211 29323 23247 29357
rect 23281 29323 23317 29357
rect 23351 29323 23387 29357
rect 23421 29323 23457 29357
rect 23491 29323 23527 29357
rect 23561 29323 23597 29357
rect 23631 29323 23635 29357
rect 22823 29299 22842 29323
rect 22876 29299 23635 29323
rect 22823 29289 23635 29299
rect 22823 29255 22827 29289
rect 22861 29261 22897 29289
rect 22876 29255 22897 29261
rect 22931 29255 22967 29289
rect 23001 29255 23037 29289
rect 23071 29255 23107 29289
rect 23141 29255 23177 29289
rect 23211 29255 23247 29289
rect 23281 29255 23317 29289
rect 23351 29255 23387 29289
rect 23421 29255 23457 29289
rect 23491 29255 23527 29289
rect 23561 29255 23597 29289
rect 23631 29255 23635 29289
rect 22823 29227 22842 29255
rect 22876 29227 23635 29255
rect 22823 29221 23635 29227
rect 22823 29187 22827 29221
rect 22861 29189 22897 29221
rect 22876 29187 22897 29189
rect 22931 29187 22967 29221
rect 23001 29187 23037 29221
rect 23071 29187 23107 29221
rect 23141 29187 23177 29221
rect 23211 29187 23247 29221
rect 23281 29187 23317 29221
rect 23351 29187 23387 29221
rect 23421 29187 23457 29221
rect 23491 29187 23527 29221
rect 23561 29187 23597 29221
rect 23631 29187 23635 29221
rect 22823 29155 22842 29187
rect 22876 29155 23635 29187
rect 22823 29153 23635 29155
rect 22823 29119 22827 29153
rect 22861 29119 22897 29153
rect 22931 29119 22967 29153
rect 23001 29119 23037 29153
rect 23071 29119 23107 29153
rect 23141 29119 23177 29153
rect 23211 29119 23247 29153
rect 23281 29119 23317 29153
rect 23351 29119 23387 29153
rect 23421 29119 23457 29153
rect 23491 29119 23527 29153
rect 23561 29119 23597 29153
rect 23631 29119 23635 29153
rect 22823 29117 23635 29119
rect 22823 29085 22842 29117
rect 22876 29085 23635 29117
rect 22823 29051 22827 29085
rect 22876 29083 22897 29085
rect 22861 29051 22897 29083
rect 22931 29051 22967 29085
rect 23001 29051 23037 29085
rect 23071 29051 23107 29085
rect 23141 29051 23177 29085
rect 23211 29051 23247 29085
rect 23281 29051 23317 29085
rect 23351 29051 23387 29085
rect 23421 29051 23457 29085
rect 23491 29051 23527 29085
rect 23561 29051 23597 29085
rect 23631 29051 23635 29085
rect 22823 29045 23635 29051
rect 22823 29017 22842 29045
rect 22876 29017 23635 29045
rect 22823 28983 22827 29017
rect 22876 29011 22897 29017
rect 22861 28983 22897 29011
rect 22931 28983 22967 29017
rect 23001 28983 23037 29017
rect 23071 28983 23107 29017
rect 23141 28983 23177 29017
rect 23211 28983 23247 29017
rect 23281 28983 23317 29017
rect 23351 28983 23387 29017
rect 23421 28983 23457 29017
rect 23491 28983 23527 29017
rect 23561 28983 23597 29017
rect 23631 28983 23635 29017
rect 22823 28973 23635 28983
rect 22823 28949 22842 28973
rect 22876 28949 23635 28973
rect 22823 28915 22827 28949
rect 22876 28939 22897 28949
rect 22861 28915 22897 28939
rect 22931 28915 22967 28949
rect 23001 28915 23037 28949
rect 23071 28915 23107 28949
rect 23141 28915 23177 28949
rect 23211 28915 23247 28949
rect 23281 28915 23317 28949
rect 23351 28915 23387 28949
rect 23421 28915 23457 28949
rect 23491 28915 23527 28949
rect 23561 28915 23597 28949
rect 23631 28915 23635 28949
rect 22823 28901 23635 28915
rect 22823 28881 22842 28901
rect 22876 28881 23635 28901
rect 22823 28847 22827 28881
rect 22876 28867 22897 28881
rect 22861 28847 22897 28867
rect 22931 28847 22967 28881
rect 23001 28847 23037 28881
rect 23071 28847 23107 28881
rect 23141 28847 23177 28881
rect 23211 28847 23247 28881
rect 23281 28847 23317 28881
rect 23351 28847 23387 28881
rect 23421 28847 23457 28881
rect 23491 28847 23527 28881
rect 23561 28847 23597 28881
rect 23631 28847 23635 28881
rect 22823 28829 23635 28847
rect 22823 28813 22842 28829
rect 22876 28813 23635 28829
rect 22823 28779 22827 28813
rect 22876 28795 22897 28813
rect 22861 28779 22897 28795
rect 22931 28779 22967 28813
rect 23001 28779 23037 28813
rect 23071 28779 23107 28813
rect 23141 28779 23177 28813
rect 23211 28779 23247 28813
rect 23281 28779 23317 28813
rect 23351 28779 23387 28813
rect 23421 28779 23457 28813
rect 23491 28779 23527 28813
rect 23561 28779 23597 28813
rect 23631 28779 23635 28813
rect 22823 28757 23635 28779
rect 22823 28745 22842 28757
rect 22876 28745 23635 28757
rect 22823 28711 22827 28745
rect 22876 28723 22897 28745
rect 22861 28711 22897 28723
rect 22931 28711 22967 28745
rect 23001 28711 23037 28745
rect 23071 28711 23107 28745
rect 23141 28711 23177 28745
rect 23211 28711 23247 28745
rect 23281 28711 23317 28745
rect 23351 28711 23387 28745
rect 23421 28711 23457 28745
rect 23491 28711 23527 28745
rect 23561 28711 23597 28745
rect 23631 28711 23635 28745
rect 22823 28685 23635 28711
rect 22823 28677 22842 28685
rect 22876 28677 23635 28685
rect 22823 28643 22827 28677
rect 22876 28651 22897 28677
rect 22861 28643 22897 28651
rect 22931 28643 22967 28677
rect 23001 28643 23037 28677
rect 23071 28643 23107 28677
rect 23141 28643 23177 28677
rect 23211 28643 23247 28677
rect 23281 28643 23317 28677
rect 23351 28643 23387 28677
rect 23421 28643 23457 28677
rect 23491 28643 23527 28677
rect 23561 28643 23597 28677
rect 23631 28643 23635 28677
rect 22823 28613 23635 28643
rect 22823 28609 22842 28613
rect 22876 28609 23635 28613
rect 22823 28575 22827 28609
rect 22876 28579 22897 28609
rect 22861 28575 22897 28579
rect 22931 28575 22967 28609
rect 23001 28575 23037 28609
rect 23071 28575 23107 28609
rect 23141 28575 23177 28609
rect 23211 28575 23247 28609
rect 23281 28575 23317 28609
rect 23351 28575 23387 28609
rect 23421 28575 23457 28609
rect 23491 28575 23527 28609
rect 23561 28575 23597 28609
rect 23631 28575 23635 28609
rect 22823 28541 23635 28575
rect 22823 28507 22827 28541
rect 22876 28507 22897 28541
rect 22931 28507 22967 28541
rect 23001 28507 23037 28541
rect 23071 28507 23107 28541
rect 23141 28507 23177 28541
rect 23211 28507 23247 28541
rect 23281 28507 23317 28541
rect 23351 28507 23387 28541
rect 23421 28507 23457 28541
rect 23491 28507 23527 28541
rect 23561 28507 23597 28541
rect 23631 28507 23635 28541
rect 22823 28473 23635 28507
rect 22823 28439 22827 28473
rect 22861 28469 22897 28473
rect 22876 28439 22897 28469
rect 22931 28439 22967 28473
rect 23001 28439 23037 28473
rect 23071 28439 23107 28473
rect 23141 28439 23177 28473
rect 23211 28439 23247 28473
rect 23281 28439 23317 28473
rect 23351 28439 23387 28473
rect 23421 28439 23457 28473
rect 23491 28439 23527 28473
rect 23561 28439 23597 28473
rect 23631 28439 23635 28473
rect 22823 28435 22842 28439
rect 22876 28435 23635 28439
rect 22823 28405 23635 28435
rect 22823 28371 22827 28405
rect 22861 28397 22897 28405
rect 22876 28371 22897 28397
rect 22931 28371 22967 28405
rect 23001 28371 23037 28405
rect 23071 28371 23107 28405
rect 23141 28371 23177 28405
rect 23211 28371 23247 28405
rect 23281 28371 23317 28405
rect 23351 28371 23387 28405
rect 23421 28371 23457 28405
rect 23491 28371 23527 28405
rect 23561 28371 23597 28405
rect 23631 28371 23635 28405
rect 22823 28363 22842 28371
rect 22876 28363 23635 28371
rect 22823 28337 23635 28363
rect 22823 28303 22827 28337
rect 22861 28325 22897 28337
rect 22876 28303 22897 28325
rect 22931 28303 22967 28337
rect 23001 28303 23037 28337
rect 23071 28303 23107 28337
rect 23141 28303 23177 28337
rect 23211 28303 23247 28337
rect 23281 28303 23317 28337
rect 23351 28303 23387 28337
rect 23421 28303 23457 28337
rect 23491 28303 23527 28337
rect 23561 28303 23597 28337
rect 23631 28303 23635 28337
rect 22823 28291 22842 28303
rect 22876 28291 23635 28303
rect 22823 28269 23635 28291
rect 22823 28235 22827 28269
rect 22861 28253 22897 28269
rect 22876 28235 22897 28253
rect 22931 28235 22967 28269
rect 23001 28235 23037 28269
rect 23071 28235 23107 28269
rect 23141 28235 23177 28269
rect 23211 28235 23247 28269
rect 23281 28235 23317 28269
rect 23351 28235 23387 28269
rect 23421 28235 23457 28269
rect 23491 28235 23527 28269
rect 23561 28235 23597 28269
rect 23631 28235 23635 28269
rect 22823 28219 22842 28235
rect 22876 28219 23635 28235
rect 22823 28201 23635 28219
rect 22823 28167 22827 28201
rect 22861 28181 22897 28201
rect 22876 28167 22897 28181
rect 22931 28167 22967 28201
rect 23001 28167 23037 28201
rect 23071 28167 23107 28201
rect 23141 28167 23177 28201
rect 23211 28167 23247 28201
rect 23281 28167 23317 28201
rect 23351 28167 23387 28201
rect 23421 28167 23457 28201
rect 23491 28167 23527 28201
rect 23561 28167 23597 28201
rect 23631 28167 23635 28201
rect 22823 28147 22842 28167
rect 22876 28147 23635 28167
rect 22823 28133 23635 28147
rect 22823 28099 22827 28133
rect 22861 28109 22897 28133
rect 22876 28099 22897 28109
rect 22931 28099 22967 28133
rect 23001 28099 23037 28133
rect 23071 28099 23107 28133
rect 23141 28099 23177 28133
rect 23211 28099 23247 28133
rect 23281 28099 23317 28133
rect 23351 28099 23387 28133
rect 23421 28099 23457 28133
rect 23491 28099 23527 28133
rect 23561 28099 23597 28133
rect 23631 28099 23635 28133
rect 22823 28075 22842 28099
rect 22876 28075 23635 28099
rect 22823 28065 23635 28075
rect 22823 28031 22827 28065
rect 22861 28037 22897 28065
rect 22876 28031 22897 28037
rect 22931 28031 22967 28065
rect 23001 28031 23037 28065
rect 23071 28031 23107 28065
rect 23141 28031 23177 28065
rect 23211 28031 23247 28065
rect 23281 28031 23317 28065
rect 23351 28031 23387 28065
rect 23421 28031 23457 28065
rect 23491 28031 23527 28065
rect 23561 28031 23597 28065
rect 23631 28031 23635 28065
rect 22823 28003 22842 28031
rect 22876 28003 23635 28031
rect 22823 27997 23635 28003
rect 22823 27963 22827 27997
rect 22861 27965 22897 27997
rect 22876 27963 22897 27965
rect 22931 27963 22967 27997
rect 23001 27963 23037 27997
rect 23071 27963 23107 27997
rect 23141 27963 23177 27997
rect 23211 27963 23247 27997
rect 23281 27963 23317 27997
rect 23351 27963 23387 27997
rect 23421 27963 23457 27997
rect 23491 27963 23527 27997
rect 23561 27963 23597 27997
rect 23631 27963 23635 27997
rect 22823 27931 22842 27963
rect 22876 27931 23635 27963
rect 22823 27929 23635 27931
rect 22823 27895 22827 27929
rect 22861 27895 22897 27929
rect 22931 27895 22967 27929
rect 23001 27895 23037 27929
rect 23071 27895 23107 27929
rect 23141 27895 23177 27929
rect 23211 27895 23247 27929
rect 23281 27895 23317 27929
rect 23351 27895 23387 27929
rect 23421 27895 23457 27929
rect 23491 27895 23527 27929
rect 23561 27895 23597 27929
rect 23631 27895 23635 27929
rect 22823 27893 23635 27895
rect 22823 27861 22842 27893
rect 22876 27861 23635 27893
rect 22823 27827 22827 27861
rect 22876 27859 22897 27861
rect 22861 27827 22897 27859
rect 22931 27827 22967 27861
rect 23001 27827 23037 27861
rect 23071 27827 23107 27861
rect 23141 27827 23177 27861
rect 23211 27827 23247 27861
rect 23281 27827 23317 27861
rect 23351 27827 23387 27861
rect 23421 27827 23457 27861
rect 23491 27827 23527 27861
rect 23561 27827 23597 27861
rect 23631 27827 23635 27861
rect 22823 27821 23635 27827
rect 22823 27793 22842 27821
rect 22876 27793 23635 27821
rect 22823 27759 22827 27793
rect 22876 27787 22897 27793
rect 22861 27759 22897 27787
rect 22931 27759 22967 27793
rect 23001 27759 23037 27793
rect 23071 27759 23107 27793
rect 23141 27759 23177 27793
rect 23211 27759 23247 27793
rect 23281 27759 23317 27793
rect 23351 27759 23387 27793
rect 23421 27759 23457 27793
rect 23491 27759 23527 27793
rect 23561 27759 23597 27793
rect 23631 27759 23635 27793
rect 22823 27749 23635 27759
rect 22823 27725 22842 27749
rect 22876 27725 23635 27749
rect 22823 27691 22827 27725
rect 22876 27715 22897 27725
rect 22861 27691 22897 27715
rect 22931 27691 22967 27725
rect 23001 27691 23037 27725
rect 23071 27691 23107 27725
rect 23141 27691 23177 27725
rect 23211 27691 23247 27725
rect 23281 27691 23317 27725
rect 23351 27691 23387 27725
rect 23421 27691 23457 27725
rect 23491 27691 23527 27725
rect 23561 27691 23597 27725
rect 23631 27691 23635 27725
rect 22823 27677 23635 27691
rect 22823 27657 22842 27677
rect 22876 27657 23635 27677
rect 22823 27623 22827 27657
rect 22876 27643 22897 27657
rect 22861 27623 22897 27643
rect 22931 27623 22967 27657
rect 23001 27623 23037 27657
rect 23071 27623 23107 27657
rect 23141 27623 23177 27657
rect 23211 27623 23247 27657
rect 23281 27623 23317 27657
rect 23351 27623 23387 27657
rect 23421 27623 23457 27657
rect 23491 27623 23527 27657
rect 23561 27623 23597 27657
rect 23631 27623 23635 27657
rect 22823 27605 23635 27623
rect 22823 27589 22842 27605
rect 22876 27589 23635 27605
rect 22823 27555 22827 27589
rect 22876 27571 22897 27589
rect 22861 27555 22897 27571
rect 22931 27555 22967 27589
rect 23001 27555 23037 27589
rect 23071 27555 23107 27589
rect 23141 27555 23177 27589
rect 23211 27555 23247 27589
rect 23281 27555 23317 27589
rect 23351 27555 23387 27589
rect 23421 27555 23457 27589
rect 23491 27555 23527 27589
rect 23561 27555 23597 27589
rect 23631 27555 23635 27589
rect 22823 27533 23635 27555
rect 22823 27521 22842 27533
rect 22876 27521 23635 27533
rect 22823 27487 22827 27521
rect 22876 27499 22897 27521
rect 22861 27487 22897 27499
rect 22931 27487 22967 27521
rect 23001 27487 23037 27521
rect 23071 27487 23107 27521
rect 23141 27487 23177 27521
rect 23211 27487 23247 27521
rect 23281 27487 23317 27521
rect 23351 27487 23387 27521
rect 23421 27487 23457 27521
rect 23491 27487 23527 27521
rect 23561 27487 23597 27521
rect 23631 27487 23635 27521
rect 22823 27461 23635 27487
rect 22823 27453 22842 27461
rect 22876 27453 23635 27461
rect 22823 27419 22827 27453
rect 22876 27427 22897 27453
rect 22861 27419 22897 27427
rect 22931 27419 22967 27453
rect 23001 27419 23037 27453
rect 23071 27419 23107 27453
rect 23141 27419 23177 27453
rect 23211 27419 23247 27453
rect 23281 27419 23317 27453
rect 23351 27419 23387 27453
rect 23421 27419 23457 27453
rect 23491 27419 23527 27453
rect 23561 27419 23597 27453
rect 23631 27419 23635 27453
rect 22823 27389 23635 27419
rect 22823 27385 22842 27389
rect 22876 27385 23635 27389
rect 22823 27351 22827 27385
rect 22876 27355 22897 27385
rect 22861 27351 22897 27355
rect 22931 27351 22967 27385
rect 23001 27351 23037 27385
rect 23071 27351 23107 27385
rect 23141 27351 23177 27385
rect 23211 27351 23247 27385
rect 23281 27351 23317 27385
rect 23351 27351 23387 27385
rect 23421 27351 23457 27385
rect 23491 27351 23527 27385
rect 23561 27351 23597 27385
rect 23631 27351 23635 27385
rect 22823 27317 23635 27351
rect 22823 27283 22827 27317
rect 22876 27283 22897 27317
rect 22931 27283 22967 27317
rect 23001 27283 23037 27317
rect 23071 27283 23107 27317
rect 23141 27283 23177 27317
rect 23211 27283 23247 27317
rect 23281 27283 23317 27317
rect 23351 27283 23387 27317
rect 23421 27283 23457 27317
rect 23491 27283 23527 27317
rect 23561 27283 23597 27317
rect 23631 27283 23635 27317
rect 22823 27249 23635 27283
rect 22823 27215 22827 27249
rect 22861 27245 22897 27249
rect 22876 27215 22897 27245
rect 22931 27215 22967 27249
rect 23001 27215 23037 27249
rect 23071 27215 23107 27249
rect 23141 27215 23177 27249
rect 23211 27215 23247 27249
rect 23281 27215 23317 27249
rect 23351 27215 23387 27249
rect 23421 27215 23457 27249
rect 23491 27215 23527 27249
rect 23561 27215 23597 27249
rect 23631 27215 23635 27249
rect 22823 27211 22842 27215
rect 22876 27211 23635 27215
rect 22823 27181 23635 27211
rect 22823 27147 22827 27181
rect 22861 27173 22897 27181
rect 22876 27147 22897 27173
rect 22931 27147 22967 27181
rect 23001 27147 23037 27181
rect 23071 27147 23107 27181
rect 23141 27147 23177 27181
rect 23211 27147 23247 27181
rect 23281 27147 23317 27181
rect 23351 27147 23387 27181
rect 23421 27147 23457 27181
rect 23491 27147 23527 27181
rect 23561 27147 23597 27181
rect 23631 27147 23635 27181
rect 22823 27139 22842 27147
rect 22876 27139 23635 27147
rect 22823 27113 23635 27139
rect 22823 27079 22827 27113
rect 22861 27101 22897 27113
rect 22876 27079 22897 27101
rect 22931 27079 22967 27113
rect 23001 27079 23037 27113
rect 23071 27079 23107 27113
rect 23141 27079 23177 27113
rect 23211 27079 23247 27113
rect 23281 27079 23317 27113
rect 23351 27079 23387 27113
rect 23421 27079 23457 27113
rect 23491 27079 23527 27113
rect 23561 27079 23597 27113
rect 23631 27079 23635 27113
rect 22823 27067 22842 27079
rect 22876 27067 23635 27079
rect 22823 27045 23635 27067
rect 22823 27011 22827 27045
rect 22861 27029 22897 27045
rect 22876 27011 22897 27029
rect 22931 27011 22967 27045
rect 23001 27011 23037 27045
rect 23071 27011 23107 27045
rect 23141 27011 23177 27045
rect 23211 27011 23247 27045
rect 23281 27011 23317 27045
rect 23351 27011 23387 27045
rect 23421 27011 23457 27045
rect 23491 27011 23527 27045
rect 23561 27011 23597 27045
rect 23631 27011 23635 27045
rect 22823 26995 22842 27011
rect 22876 26995 23635 27011
rect 22823 26977 23635 26995
rect 22823 26943 22827 26977
rect 22861 26957 22897 26977
rect 22876 26943 22897 26957
rect 22931 26943 22967 26977
rect 23001 26943 23037 26977
rect 23071 26943 23107 26977
rect 23141 26943 23177 26977
rect 23211 26943 23247 26977
rect 23281 26943 23317 26977
rect 23351 26943 23387 26977
rect 23421 26943 23457 26977
rect 23491 26943 23527 26977
rect 23561 26943 23597 26977
rect 23631 26943 23635 26977
rect 22823 26923 22842 26943
rect 22876 26923 23635 26943
rect 22823 26909 23635 26923
rect 22823 26875 22827 26909
rect 22861 26885 22897 26909
rect 22876 26875 22897 26885
rect 22931 26875 22967 26909
rect 23001 26875 23037 26909
rect 23071 26875 23107 26909
rect 23141 26875 23177 26909
rect 23211 26875 23247 26909
rect 23281 26875 23317 26909
rect 23351 26875 23387 26909
rect 23421 26875 23457 26909
rect 23491 26875 23527 26909
rect 23561 26875 23597 26909
rect 23631 26875 23635 26909
rect 22823 26851 22842 26875
rect 22876 26851 23635 26875
rect 22823 26841 23635 26851
rect 22823 26807 22827 26841
rect 22861 26813 22897 26841
rect 22876 26807 22897 26813
rect 22931 26807 22967 26841
rect 23001 26807 23037 26841
rect 23071 26807 23107 26841
rect 23141 26807 23177 26841
rect 23211 26807 23247 26841
rect 23281 26807 23317 26841
rect 23351 26807 23387 26841
rect 23421 26807 23457 26841
rect 23491 26807 23527 26841
rect 23561 26807 23597 26841
rect 23631 26807 23635 26841
rect 22823 26779 22842 26807
rect 22876 26779 23635 26807
rect 22823 26773 23635 26779
rect 22823 26739 22827 26773
rect 22861 26741 22897 26773
rect 22876 26739 22897 26741
rect 22931 26739 22967 26773
rect 23001 26739 23037 26773
rect 23071 26739 23107 26773
rect 23141 26739 23177 26773
rect 23211 26739 23247 26773
rect 23281 26739 23317 26773
rect 23351 26739 23387 26773
rect 23421 26739 23457 26773
rect 23491 26739 23527 26773
rect 23561 26739 23597 26773
rect 23631 26739 23635 26773
rect 22823 26707 22842 26739
rect 22876 26707 23635 26739
rect 22823 26705 23635 26707
rect 22823 26671 22827 26705
rect 22861 26671 22897 26705
rect 22931 26671 22967 26705
rect 23001 26671 23037 26705
rect 23071 26671 23107 26705
rect 23141 26671 23177 26705
rect 23211 26671 23247 26705
rect 23281 26671 23317 26705
rect 23351 26671 23387 26705
rect 23421 26671 23457 26705
rect 23491 26671 23527 26705
rect 23561 26671 23597 26705
rect 23631 26671 23635 26705
rect 22823 26669 23635 26671
rect 22823 26637 22842 26669
rect 22876 26637 23635 26669
rect 22823 26603 22827 26637
rect 22876 26635 22897 26637
rect 22861 26603 22897 26635
rect 22931 26603 22967 26637
rect 23001 26603 23037 26637
rect 23071 26603 23107 26637
rect 23141 26603 23177 26637
rect 23211 26603 23247 26637
rect 23281 26603 23317 26637
rect 23351 26603 23387 26637
rect 23421 26603 23457 26637
rect 23491 26603 23527 26637
rect 23561 26603 23597 26637
rect 23631 26603 23635 26637
rect 22823 26597 23635 26603
rect 22823 26569 22842 26597
rect 22876 26569 23635 26597
rect 22823 26535 22827 26569
rect 22876 26563 22897 26569
rect 22861 26535 22897 26563
rect 22931 26535 22967 26569
rect 23001 26535 23037 26569
rect 23071 26535 23107 26569
rect 23141 26535 23177 26569
rect 23211 26535 23247 26569
rect 23281 26535 23317 26569
rect 23351 26535 23387 26569
rect 23421 26535 23457 26569
rect 23491 26535 23527 26569
rect 23561 26535 23597 26569
rect 23631 26535 23635 26569
rect 22823 26525 23635 26535
rect 22823 26501 22842 26525
rect 22876 26501 23635 26525
rect 22823 26467 22827 26501
rect 22876 26491 22897 26501
rect 22861 26467 22897 26491
rect 22931 26467 22967 26501
rect 23001 26467 23037 26501
rect 23071 26467 23107 26501
rect 23141 26467 23177 26501
rect 23211 26467 23247 26501
rect 23281 26467 23317 26501
rect 23351 26467 23387 26501
rect 23421 26467 23457 26501
rect 23491 26467 23527 26501
rect 23561 26467 23597 26501
rect 23631 26467 23635 26501
rect 22823 26453 23635 26467
rect 22823 26433 22842 26453
rect 22876 26433 23635 26453
rect 22823 26399 22827 26433
rect 22876 26419 22897 26433
rect 22861 26399 22897 26419
rect 22931 26399 22967 26433
rect 23001 26399 23037 26433
rect 23071 26399 23107 26433
rect 23141 26399 23177 26433
rect 23211 26399 23247 26433
rect 23281 26399 23317 26433
rect 23351 26399 23387 26433
rect 23421 26399 23457 26433
rect 23491 26399 23527 26433
rect 23561 26399 23597 26433
rect 23631 26399 23635 26433
rect 22823 26381 23635 26399
rect 22823 26365 22842 26381
rect 22876 26365 23635 26381
rect 22823 26331 22827 26365
rect 22876 26347 22897 26365
rect 22861 26331 22897 26347
rect 22931 26331 22967 26365
rect 23001 26331 23037 26365
rect 23071 26331 23107 26365
rect 23141 26331 23177 26365
rect 23211 26331 23247 26365
rect 23281 26331 23317 26365
rect 23351 26331 23387 26365
rect 23421 26331 23457 26365
rect 23491 26331 23527 26365
rect 23561 26331 23597 26365
rect 23631 26331 23635 26365
rect 22823 26309 23635 26331
rect 22823 26297 22842 26309
rect 22876 26297 23635 26309
rect 22823 26263 22827 26297
rect 22876 26275 22897 26297
rect 22861 26263 22897 26275
rect 22931 26263 22967 26297
rect 23001 26263 23037 26297
rect 23071 26263 23107 26297
rect 23141 26263 23177 26297
rect 23211 26263 23247 26297
rect 23281 26263 23317 26297
rect 23351 26263 23387 26297
rect 23421 26263 23457 26297
rect 23491 26263 23527 26297
rect 23561 26263 23597 26297
rect 23631 26263 23635 26297
rect 22823 26237 23635 26263
rect 22823 26229 22842 26237
rect 22876 26229 23635 26237
rect 22823 26195 22827 26229
rect 22876 26203 22897 26229
rect 22861 26195 22897 26203
rect 22931 26195 22967 26229
rect 23001 26195 23037 26229
rect 23071 26195 23107 26229
rect 23141 26195 23177 26229
rect 23211 26195 23247 26229
rect 23281 26195 23317 26229
rect 23351 26195 23387 26229
rect 23421 26195 23457 26229
rect 23491 26195 23527 26229
rect 23561 26195 23597 26229
rect 23631 26195 23635 26229
rect 22823 26165 23635 26195
rect 22823 26161 22842 26165
rect 22876 26161 23635 26165
rect 22823 26127 22827 26161
rect 22876 26131 22897 26161
rect 22861 26127 22897 26131
rect 22931 26127 22967 26161
rect 23001 26127 23037 26161
rect 23071 26127 23107 26161
rect 23141 26127 23177 26161
rect 23211 26127 23247 26161
rect 23281 26127 23317 26161
rect 23351 26127 23387 26161
rect 23421 26127 23457 26161
rect 23491 26127 23527 26161
rect 23561 26127 23597 26161
rect 23631 26127 23635 26161
rect 22823 26093 23635 26127
rect 22823 26059 22827 26093
rect 22876 26059 22897 26093
rect 22931 26059 22967 26093
rect 23001 26059 23037 26093
rect 23071 26059 23107 26093
rect 23141 26059 23177 26093
rect 23211 26059 23247 26093
rect 23281 26059 23317 26093
rect 23351 26059 23387 26093
rect 23421 26059 23457 26093
rect 23491 26059 23527 26093
rect 23561 26059 23597 26093
rect 23631 26059 23635 26093
rect 22823 26025 23635 26059
rect 22823 25991 22827 26025
rect 22861 26021 22897 26025
rect 22876 25991 22897 26021
rect 22931 25991 22967 26025
rect 23001 25991 23037 26025
rect 23071 25991 23107 26025
rect 23141 25991 23177 26025
rect 23211 25991 23247 26025
rect 23281 25991 23317 26025
rect 23351 25991 23387 26025
rect 23421 25991 23457 26025
rect 23491 25991 23527 26025
rect 23561 25991 23597 26025
rect 23631 25991 23635 26025
rect 22823 25987 22842 25991
rect 22876 25987 23635 25991
rect 22823 25957 23635 25987
rect 22823 25923 22827 25957
rect 22861 25949 22897 25957
rect 22876 25923 22897 25949
rect 22931 25923 22967 25957
rect 23001 25923 23037 25957
rect 23071 25923 23107 25957
rect 23141 25923 23177 25957
rect 23211 25923 23247 25957
rect 23281 25923 23317 25957
rect 23351 25923 23387 25957
rect 23421 25923 23457 25957
rect 23491 25923 23527 25957
rect 23561 25923 23597 25957
rect 23631 25923 23635 25957
rect 22823 25915 22842 25923
rect 22876 25915 23635 25923
rect 22823 25889 23635 25915
rect 22823 25855 22827 25889
rect 22861 25877 22897 25889
rect 22876 25855 22897 25877
rect 22931 25855 22967 25889
rect 23001 25855 23037 25889
rect 23071 25855 23107 25889
rect 23141 25855 23177 25889
rect 23211 25855 23247 25889
rect 23281 25855 23317 25889
rect 23351 25855 23387 25889
rect 23421 25855 23457 25889
rect 23491 25855 23527 25889
rect 23561 25855 23597 25889
rect 23631 25855 23635 25889
rect 22823 25843 22842 25855
rect 22876 25843 23635 25855
rect 22823 25821 23635 25843
rect 22823 25787 22827 25821
rect 22861 25805 22897 25821
rect 22876 25787 22897 25805
rect 22931 25787 22967 25821
rect 23001 25787 23037 25821
rect 23071 25787 23107 25821
rect 23141 25787 23177 25821
rect 23211 25787 23247 25821
rect 23281 25787 23317 25821
rect 23351 25787 23387 25821
rect 23421 25787 23457 25821
rect 23491 25787 23527 25821
rect 23561 25787 23597 25821
rect 23631 25787 23635 25821
rect 22823 25771 22842 25787
rect 22876 25771 23635 25787
rect 22823 25753 23635 25771
rect 22823 25719 22827 25753
rect 22861 25733 22897 25753
rect 22876 25719 22897 25733
rect 22931 25719 22967 25753
rect 23001 25719 23037 25753
rect 23071 25719 23107 25753
rect 23141 25719 23177 25753
rect 23211 25719 23247 25753
rect 23281 25719 23317 25753
rect 23351 25719 23387 25753
rect 23421 25719 23457 25753
rect 23491 25719 23527 25753
rect 23561 25719 23597 25753
rect 23631 25719 23635 25753
rect 22823 25699 22842 25719
rect 22876 25699 23635 25719
rect 22823 25685 23635 25699
rect 22823 25651 22827 25685
rect 22861 25661 22897 25685
rect 22876 25651 22897 25661
rect 22931 25651 22967 25685
rect 23001 25651 23037 25685
rect 23071 25651 23107 25685
rect 23141 25651 23177 25685
rect 23211 25651 23247 25685
rect 23281 25651 23317 25685
rect 23351 25651 23387 25685
rect 23421 25651 23457 25685
rect 23491 25651 23527 25685
rect 23561 25651 23597 25685
rect 23631 25651 23635 25685
rect 22823 25627 22842 25651
rect 22876 25627 23635 25651
rect 22823 25617 23635 25627
rect 22823 25583 22827 25617
rect 22861 25589 22897 25617
rect 22876 25583 22897 25589
rect 22931 25583 22967 25617
rect 23001 25583 23037 25617
rect 23071 25583 23107 25617
rect 23141 25583 23177 25617
rect 23211 25583 23247 25617
rect 23281 25583 23317 25617
rect 23351 25583 23387 25617
rect 23421 25583 23457 25617
rect 23491 25583 23527 25617
rect 23561 25583 23597 25617
rect 23631 25583 23635 25617
rect 22823 25555 22842 25583
rect 22876 25555 23635 25583
rect 22823 25549 23635 25555
rect 22823 25515 22827 25549
rect 22861 25517 22897 25549
rect 22876 25515 22897 25517
rect 22931 25515 22967 25549
rect 23001 25515 23037 25549
rect 23071 25515 23107 25549
rect 23141 25515 23177 25549
rect 23211 25515 23247 25549
rect 23281 25515 23317 25549
rect 23351 25515 23387 25549
rect 23421 25515 23457 25549
rect 23491 25515 23527 25549
rect 23561 25515 23597 25549
rect 23631 25515 23635 25549
rect 22823 25483 22842 25515
rect 22876 25483 23635 25515
rect 22823 25481 23635 25483
rect 22823 25447 22827 25481
rect 22861 25447 22897 25481
rect 22931 25447 22967 25481
rect 23001 25447 23037 25481
rect 23071 25447 23107 25481
rect 23141 25447 23177 25481
rect 23211 25447 23247 25481
rect 23281 25447 23317 25481
rect 23351 25447 23387 25481
rect 23421 25447 23457 25481
rect 23491 25447 23527 25481
rect 23561 25447 23597 25481
rect 23631 25447 23635 25481
rect 22823 25445 23635 25447
rect 22823 25413 22842 25445
rect 22876 25413 23635 25445
rect 22823 25379 22827 25413
rect 22876 25411 22897 25413
rect 22861 25379 22897 25411
rect 22931 25379 22967 25413
rect 23001 25379 23037 25413
rect 23071 25379 23107 25413
rect 23141 25379 23177 25413
rect 23211 25379 23247 25413
rect 23281 25379 23317 25413
rect 23351 25379 23387 25413
rect 23421 25379 23457 25413
rect 23491 25379 23527 25413
rect 23561 25379 23597 25413
rect 23631 25379 23635 25413
rect 22823 25373 23635 25379
rect 22823 25345 22842 25373
rect 22876 25345 23635 25373
rect 22823 25311 22827 25345
rect 22876 25339 22897 25345
rect 22861 25311 22897 25339
rect 22931 25311 22967 25345
rect 23001 25311 23037 25345
rect 23071 25311 23107 25345
rect 23141 25311 23177 25345
rect 23211 25311 23247 25345
rect 23281 25311 23317 25345
rect 23351 25311 23387 25345
rect 23421 25311 23457 25345
rect 23491 25311 23527 25345
rect 23561 25311 23597 25345
rect 23631 25311 23635 25345
rect 22823 25300 23635 25311
rect 22823 25277 22842 25300
rect 22876 25277 23635 25300
rect 22823 25243 22827 25277
rect 22876 25266 22897 25277
rect 22861 25243 22897 25266
rect 22931 25243 22967 25277
rect 23001 25243 23037 25277
rect 23071 25243 23107 25277
rect 23141 25243 23177 25277
rect 23211 25243 23247 25277
rect 23281 25243 23317 25277
rect 23351 25243 23387 25277
rect 23421 25243 23457 25277
rect 23491 25243 23527 25277
rect 23561 25243 23597 25277
rect 23631 25243 23635 25277
rect 22823 25227 23635 25243
rect 22823 25209 22842 25227
rect 22876 25209 23635 25227
rect 22823 25175 22827 25209
rect 22876 25193 22897 25209
rect 22861 25175 22897 25193
rect 22931 25175 22967 25209
rect 23001 25175 23037 25209
rect 23071 25175 23107 25209
rect 23141 25175 23177 25209
rect 23211 25175 23247 25209
rect 23281 25175 23317 25209
rect 23351 25175 23387 25209
rect 23421 25175 23457 25209
rect 23491 25175 23527 25209
rect 23561 25175 23597 25209
rect 23631 25175 23635 25209
rect 22823 25154 23635 25175
rect 22823 25140 22842 25154
rect 22876 25140 23635 25154
rect 22823 25106 22827 25140
rect 22876 25120 22897 25140
rect 22861 25106 22897 25120
rect 22931 25106 22967 25140
rect 23001 25106 23037 25140
rect 23071 25106 23107 25140
rect 23141 25106 23177 25140
rect 23211 25106 23247 25140
rect 23281 25106 23317 25140
rect 23351 25106 23387 25140
rect 23421 25106 23457 25140
rect 23491 25106 23527 25140
rect 23561 25106 23597 25140
rect 23631 25106 23635 25140
rect 22823 25081 23635 25106
rect 22823 25071 22842 25081
rect 22876 25071 23635 25081
rect 22823 25037 22827 25071
rect 22876 25047 22897 25071
rect 22861 25037 22897 25047
rect 22931 25037 22967 25071
rect 23001 25037 23037 25071
rect 23071 25037 23107 25071
rect 23141 25037 23177 25071
rect 23211 25037 23247 25071
rect 23281 25037 23317 25071
rect 23351 25037 23387 25071
rect 23421 25037 23457 25071
rect 23491 25037 23527 25071
rect 23561 25037 23597 25071
rect 23631 25037 23635 25071
rect 22823 25008 23635 25037
rect 22823 25002 22842 25008
rect 22876 25002 23635 25008
rect 22823 24968 22827 25002
rect 22876 24974 22897 25002
rect 22861 24968 22897 24974
rect 22931 24968 22967 25002
rect 23001 24968 23037 25002
rect 23071 24968 23107 25002
rect 23141 24968 23177 25002
rect 23211 24968 23247 25002
rect 23281 24968 23317 25002
rect 23351 24968 23387 25002
rect 23421 24968 23457 25002
rect 23491 24968 23527 25002
rect 23561 24968 23597 25002
rect 23631 24968 23635 25002
rect 22823 24935 23635 24968
rect 22823 24933 22842 24935
rect 22876 24933 23635 24935
rect 22823 24899 22827 24933
rect 22876 24901 22897 24933
rect 22861 24899 22897 24901
rect 22931 24899 22967 24933
rect 23001 24899 23037 24933
rect 23071 24899 23107 24933
rect 23141 24899 23177 24933
rect 23211 24899 23247 24933
rect 23281 24899 23317 24933
rect 23351 24899 23387 24933
rect 23421 24899 23457 24933
rect 23491 24899 23527 24933
rect 23561 24899 23597 24933
rect 23631 24899 23635 24933
rect 22823 24864 23635 24899
rect 22823 24830 22827 24864
rect 22861 24862 22897 24864
rect 22876 24830 22897 24862
rect 22931 24830 22967 24864
rect 23001 24830 23037 24864
rect 23071 24830 23107 24864
rect 23141 24830 23177 24864
rect 23211 24830 23247 24864
rect 23281 24830 23317 24864
rect 23351 24830 23387 24864
rect 23421 24830 23457 24864
rect 23491 24830 23527 24864
rect 23561 24830 23597 24864
rect 23631 24830 23635 24864
rect 22823 24828 22842 24830
rect 22876 24828 23635 24830
rect 22823 24795 23635 24828
rect 22823 24761 22827 24795
rect 22861 24789 22897 24795
rect 22876 24761 22897 24789
rect 22931 24761 22967 24795
rect 23001 24761 23037 24795
rect 23071 24761 23107 24795
rect 23141 24761 23177 24795
rect 23211 24761 23247 24795
rect 23281 24761 23317 24795
rect 23351 24761 23387 24795
rect 23421 24761 23457 24795
rect 23491 24761 23527 24795
rect 23561 24761 23597 24795
rect 23631 24761 23635 24795
rect 22823 24755 22842 24761
rect 22876 24755 23635 24761
rect 22823 24726 23635 24755
rect 22823 24692 22827 24726
rect 22861 24716 22897 24726
rect 22876 24692 22897 24716
rect 22931 24692 22967 24726
rect 23001 24692 23037 24726
rect 23071 24692 23107 24726
rect 23141 24692 23177 24726
rect 23211 24692 23247 24726
rect 23281 24692 23317 24726
rect 23351 24692 23387 24726
rect 23421 24692 23457 24726
rect 23491 24692 23527 24726
rect 23561 24692 23597 24726
rect 23631 24692 23635 24726
rect 22823 24682 22842 24692
rect 22876 24682 23635 24692
rect 22823 24657 23635 24682
rect 22823 24623 22827 24657
rect 22861 24643 22897 24657
rect 22876 24623 22897 24643
rect 22931 24623 22967 24657
rect 23001 24623 23037 24657
rect 23071 24623 23107 24657
rect 23141 24623 23177 24657
rect 23211 24623 23247 24657
rect 23281 24623 23317 24657
rect 23351 24623 23387 24657
rect 23421 24623 23457 24657
rect 23491 24623 23527 24657
rect 23561 24623 23597 24657
rect 23631 24623 23635 24657
rect 22823 24609 22842 24623
rect 22876 24609 23635 24623
rect 22823 24588 23635 24609
rect 22823 24554 22827 24588
rect 22861 24570 22897 24588
rect 22876 24554 22897 24570
rect 22931 24554 22967 24588
rect 23001 24554 23037 24588
rect 23071 24554 23107 24588
rect 23141 24554 23177 24588
rect 23211 24554 23247 24588
rect 23281 24554 23317 24588
rect 23351 24554 23387 24588
rect 23421 24554 23457 24588
rect 23491 24554 23527 24588
rect 23561 24554 23597 24588
rect 23631 24554 23635 24588
rect 22823 24536 22842 24554
rect 22876 24536 23635 24554
rect 22823 24519 23635 24536
rect 22823 24485 22827 24519
rect 22861 24497 22897 24519
rect 22876 24485 22897 24497
rect 22931 24485 22967 24519
rect 23001 24485 23037 24519
rect 23071 24485 23107 24519
rect 23141 24485 23177 24519
rect 23211 24485 23247 24519
rect 23281 24485 23317 24519
rect 23351 24485 23387 24519
rect 23421 24485 23457 24519
rect 23491 24485 23527 24519
rect 23561 24485 23597 24519
rect 23631 24485 23635 24519
rect 22823 24463 22842 24485
rect 22876 24463 23635 24485
rect 22823 24450 23635 24463
rect 22823 24416 22827 24450
rect 22861 24424 22897 24450
rect 22876 24416 22897 24424
rect 22931 24416 22967 24450
rect 23001 24416 23037 24450
rect 23071 24416 23107 24450
rect 23141 24416 23177 24450
rect 23211 24416 23247 24450
rect 23281 24416 23317 24450
rect 23351 24416 23387 24450
rect 23421 24416 23457 24450
rect 23491 24416 23527 24450
rect 23561 24416 23597 24450
rect 23631 24416 23635 24450
rect 22823 24390 22842 24416
rect 22876 24390 23635 24416
rect 22823 24381 23635 24390
rect 22823 24347 22827 24381
rect 22861 24351 22897 24381
rect 22876 24347 22897 24351
rect 22931 24347 22967 24381
rect 23001 24347 23037 24381
rect 23071 24347 23107 24381
rect 23141 24347 23177 24381
rect 23211 24347 23247 24381
rect 23281 24347 23317 24381
rect 23351 24347 23387 24381
rect 23421 24347 23457 24381
rect 23491 24347 23527 24381
rect 23561 24347 23597 24381
rect 23631 24347 23635 24381
rect 22823 24317 22842 24347
rect 22876 24317 23635 24347
rect 22823 24312 23635 24317
rect 22823 24278 22827 24312
rect 22861 24278 22897 24312
rect 22931 24278 22967 24312
rect 23001 24278 23037 24312
rect 23071 24278 23107 24312
rect 23141 24278 23177 24312
rect 23211 24278 23247 24312
rect 23281 24278 23317 24312
rect 23351 24278 23387 24312
rect 23421 24278 23457 24312
rect 23491 24278 23527 24312
rect 23561 24278 23597 24312
rect 23631 24278 23635 24312
rect 22823 24244 22842 24278
rect 22876 24244 23635 24278
rect 22823 24243 23635 24244
rect 22823 24209 22827 24243
rect 22861 24209 22897 24243
rect 22931 24209 22967 24243
rect 23001 24209 23037 24243
rect 23071 24209 23107 24243
rect 23141 24209 23177 24243
rect 23211 24209 23247 24243
rect 23281 24209 23317 24243
rect 23351 24209 23387 24243
rect 23421 24209 23457 24243
rect 23491 24209 23527 24243
rect 23561 24209 23597 24243
rect 23631 24209 23635 24243
rect 22823 24205 23635 24209
rect 22823 24174 22842 24205
rect 22876 24174 23635 24205
rect 22823 24140 22827 24174
rect 22876 24171 22897 24174
rect 22861 24140 22897 24171
rect 22931 24140 22967 24174
rect 23001 24140 23037 24174
rect 23071 24140 23107 24174
rect 23141 24140 23177 24174
rect 23211 24140 23247 24174
rect 23281 24140 23317 24174
rect 23351 24140 23387 24174
rect 23421 24140 23457 24174
rect 23491 24140 23527 24174
rect 23561 24140 23597 24174
rect 23631 24140 23635 24174
rect 22823 24132 23635 24140
rect 22823 24105 22842 24132
rect 22876 24105 23635 24132
rect 22823 24071 22827 24105
rect 22876 24098 22897 24105
rect 22861 24071 22897 24098
rect 22931 24071 22967 24105
rect 23001 24071 23037 24105
rect 23071 24071 23107 24105
rect 23141 24071 23177 24105
rect 23211 24071 23247 24105
rect 23281 24071 23317 24105
rect 23351 24071 23387 24105
rect 23421 24071 23457 24105
rect 23491 24071 23527 24105
rect 23561 24071 23597 24105
rect 23631 24071 23635 24105
rect 22823 24059 23635 24071
rect 22823 24036 22842 24059
rect 22876 24036 23635 24059
rect 22823 24002 22827 24036
rect 22876 24025 22897 24036
rect 22861 24002 22897 24025
rect 22931 24002 22967 24036
rect 23001 24002 23037 24036
rect 23071 24002 23107 24036
rect 23141 24002 23177 24036
rect 23211 24002 23247 24036
rect 23281 24002 23317 24036
rect 23351 24002 23387 24036
rect 23421 24002 23457 24036
rect 23491 24002 23527 24036
rect 23561 24002 23597 24036
rect 23631 24002 23635 24036
rect 22823 23986 23635 24002
rect 22823 23967 22842 23986
rect 22876 23967 23635 23986
rect 22823 23933 22827 23967
rect 22876 23952 22897 23967
rect 22861 23933 22897 23952
rect 22931 23933 22967 23967
rect 23001 23933 23037 23967
rect 23071 23933 23107 23967
rect 23141 23933 23177 23967
rect 23211 23933 23247 23967
rect 23281 23933 23317 23967
rect 23351 23933 23387 23967
rect 23421 23933 23457 23967
rect 23491 23933 23527 23967
rect 23561 23933 23597 23967
rect 23631 23933 23635 23967
rect 22823 23913 23635 23933
rect 22823 23898 22842 23913
rect 22876 23898 23635 23913
rect 22823 23864 22827 23898
rect 22876 23879 22897 23898
rect 22861 23864 22897 23879
rect 22931 23864 22967 23898
rect 23001 23864 23037 23898
rect 23071 23864 23107 23898
rect 23141 23864 23177 23898
rect 23211 23864 23247 23898
rect 23281 23864 23317 23898
rect 23351 23864 23387 23898
rect 23421 23864 23457 23898
rect 23491 23864 23527 23898
rect 23561 23864 23597 23898
rect 23631 23864 23635 23898
rect 22823 23840 23635 23864
rect 22823 23829 22842 23840
rect 22876 23829 23635 23840
rect 22823 23795 22827 23829
rect 22876 23806 22897 23829
rect 22861 23795 22897 23806
rect 22931 23795 22967 23829
rect 23001 23795 23037 23829
rect 23071 23795 23107 23829
rect 23141 23795 23177 23829
rect 23211 23795 23247 23829
rect 23281 23795 23317 23829
rect 23351 23795 23387 23829
rect 23421 23795 23457 23829
rect 23491 23795 23527 23829
rect 23561 23795 23597 23829
rect 23631 23795 23635 23829
rect 22823 23767 23635 23795
rect 22823 23760 22842 23767
rect 22876 23760 23635 23767
rect 22823 23726 22827 23760
rect 22876 23733 22897 23760
rect 22861 23726 22897 23733
rect 22931 23726 22967 23760
rect 23001 23726 23037 23760
rect 23071 23726 23107 23760
rect 23141 23726 23177 23760
rect 23211 23726 23247 23760
rect 23281 23726 23317 23760
rect 23351 23726 23387 23760
rect 23421 23726 23457 23760
rect 23491 23726 23527 23760
rect 23561 23726 23597 23760
rect 23631 23726 23635 23760
rect 22823 23694 23635 23726
rect 22823 23691 22842 23694
rect 22876 23691 23635 23694
rect 22823 23657 22827 23691
rect 22876 23660 22897 23691
rect 22861 23657 22897 23660
rect 22931 23657 22967 23691
rect 23001 23657 23037 23691
rect 23071 23657 23107 23691
rect 23141 23657 23177 23691
rect 23211 23657 23247 23691
rect 23281 23657 23317 23691
rect 23351 23657 23387 23691
rect 23421 23657 23457 23691
rect 23491 23657 23527 23691
rect 23561 23657 23597 23691
rect 23631 23657 23635 23691
rect 22823 23622 23635 23657
rect 22823 23588 22827 23622
rect 22861 23621 22897 23622
rect 22876 23588 22897 23621
rect 22931 23588 22967 23622
rect 23001 23588 23037 23622
rect 23071 23588 23107 23622
rect 23141 23588 23177 23622
rect 23211 23588 23247 23622
rect 23281 23588 23317 23622
rect 23351 23588 23387 23622
rect 23421 23588 23457 23622
rect 23491 23588 23527 23622
rect 23561 23588 23597 23622
rect 23631 23588 23635 23622
rect 22823 23587 22842 23588
rect 22876 23587 23635 23588
rect 22823 23553 23635 23587
rect 22823 23519 22827 23553
rect 22861 23548 22897 23553
rect 22876 23519 22897 23548
rect 22931 23519 22967 23553
rect 23001 23519 23037 23553
rect 23071 23519 23107 23553
rect 23141 23519 23177 23553
rect 23211 23519 23247 23553
rect 23281 23519 23317 23553
rect 23351 23519 23387 23553
rect 23421 23519 23457 23553
rect 23491 23519 23527 23553
rect 23561 23519 23597 23553
rect 23631 23519 23635 23553
rect 22823 23514 22842 23519
rect 22876 23514 23635 23519
rect 211 23473 1503 23474
rect 211 23439 314 23473
rect 348 23439 384 23473
rect 418 23439 454 23473
rect 488 23463 524 23473
rect 558 23463 594 23473
rect 488 23439 513 23463
rect 558 23439 590 23463
rect 628 23439 664 23473
rect 698 23463 734 23473
rect 768 23463 804 23473
rect 838 23463 874 23473
rect 908 23463 944 23473
rect 978 23463 1014 23473
rect 701 23439 734 23463
rect 778 23439 804 23463
rect 855 23439 874 23463
rect 932 23439 944 23463
rect 1009 23439 1014 23463
rect 1048 23463 1084 23473
rect 1118 23463 1154 23473
rect 1188 23463 1224 23473
rect 1258 23463 1294 23473
rect 1328 23463 1364 23473
rect 1048 23439 1052 23463
rect 1118 23439 1129 23463
rect 1188 23439 1206 23463
rect 1258 23439 1283 23463
rect 1328 23439 1360 23463
rect 1398 23439 1434 23473
rect 1468 23463 1503 23473
rect 211 23436 513 23439
rect 211 23402 212 23436
rect 246 23402 288 23436
rect 322 23403 364 23436
rect 398 23403 440 23436
rect 474 23429 513 23436
rect 547 23429 590 23439
rect 624 23429 667 23439
rect 701 23429 744 23439
rect 778 23429 821 23439
rect 855 23429 898 23439
rect 932 23429 975 23439
rect 1009 23429 1052 23439
rect 1086 23429 1129 23439
rect 1163 23429 1206 23439
rect 1240 23429 1283 23439
rect 1317 23429 1360 23439
rect 1394 23429 1437 23439
rect 1471 23429 1503 23463
rect 474 23403 1503 23429
rect 348 23402 364 23403
rect 418 23402 440 23403
rect 211 23369 314 23402
rect 348 23369 384 23402
rect 418 23369 454 23402
rect 488 23383 524 23403
rect 558 23383 594 23403
rect 488 23369 513 23383
rect 558 23369 590 23383
rect 628 23369 664 23403
rect 698 23383 734 23403
rect 768 23383 804 23403
rect 838 23383 874 23403
rect 908 23383 944 23403
rect 978 23383 1014 23403
rect 701 23369 734 23383
rect 778 23369 804 23383
rect 855 23369 874 23383
rect 932 23369 944 23383
rect 1009 23369 1014 23383
rect 1048 23383 1084 23403
rect 1118 23383 1154 23403
rect 1188 23383 1224 23403
rect 1258 23383 1294 23403
rect 1328 23383 1364 23403
rect 1048 23369 1052 23383
rect 1118 23369 1129 23383
rect 1188 23369 1206 23383
rect 1258 23369 1283 23383
rect 1328 23369 1360 23383
rect 1398 23369 1434 23403
rect 1468 23383 1503 23403
rect 211 23364 513 23369
rect 211 23330 212 23364
rect 246 23330 288 23364
rect 322 23333 364 23364
rect 398 23333 440 23364
rect 474 23349 513 23364
rect 547 23349 590 23369
rect 624 23349 667 23369
rect 701 23349 744 23369
rect 778 23349 821 23369
rect 855 23349 898 23369
rect 932 23349 975 23369
rect 1009 23349 1052 23369
rect 1086 23349 1129 23369
rect 1163 23349 1206 23369
rect 1240 23349 1283 23369
rect 1317 23349 1360 23369
rect 1394 23349 1437 23369
rect 1471 23349 1503 23383
rect 474 23333 1503 23349
rect 348 23330 364 23333
rect 418 23330 440 23333
rect 211 23299 314 23330
rect 348 23299 384 23330
rect 418 23299 454 23330
rect 488 23303 524 23333
rect 558 23303 594 23333
rect 488 23299 513 23303
rect 558 23299 590 23303
rect 628 23299 664 23333
rect 698 23303 734 23333
rect 768 23303 804 23333
rect 838 23303 874 23333
rect 908 23303 944 23333
rect 978 23303 1014 23333
rect 701 23299 734 23303
rect 778 23299 804 23303
rect 855 23299 874 23303
rect 932 23299 944 23303
rect 1009 23299 1014 23303
rect 1048 23303 1084 23333
rect 1118 23303 1154 23333
rect 1188 23303 1224 23333
rect 1258 23303 1294 23333
rect 1328 23303 1364 23333
rect 1048 23299 1052 23303
rect 1118 23299 1129 23303
rect 1188 23299 1206 23303
rect 1258 23299 1283 23303
rect 1328 23299 1360 23303
rect 1398 23299 1434 23333
rect 1468 23303 1503 23333
rect 211 23292 513 23299
rect 211 23258 212 23292
rect 246 23258 288 23292
rect 322 23263 364 23292
rect 398 23263 440 23292
rect 474 23269 513 23292
rect 547 23269 590 23299
rect 624 23269 667 23299
rect 701 23269 744 23299
rect 778 23269 821 23299
rect 855 23269 898 23299
rect 932 23269 975 23299
rect 1009 23269 1052 23299
rect 1086 23269 1129 23299
rect 1163 23269 1206 23299
rect 1240 23269 1283 23299
rect 1317 23269 1360 23299
rect 1394 23269 1437 23299
rect 1471 23269 1503 23303
rect 474 23263 1503 23269
rect 348 23258 364 23263
rect 418 23258 440 23263
rect 211 23229 314 23258
rect 348 23229 384 23258
rect 418 23229 454 23258
rect 488 23229 524 23263
rect 558 23229 594 23263
rect 628 23229 664 23263
rect 698 23229 734 23263
rect 768 23229 804 23263
rect 838 23229 874 23263
rect 908 23229 944 23263
rect 978 23229 1014 23263
rect 1048 23229 1084 23263
rect 1118 23229 1154 23263
rect 1188 23229 1224 23263
rect 1258 23229 1294 23263
rect 1328 23229 1364 23263
rect 1398 23229 1434 23263
rect 1468 23229 1503 23263
rect 211 23223 1503 23229
rect 211 23220 513 23223
rect 211 23186 212 23220
rect 246 23186 288 23220
rect 322 23193 364 23220
rect 398 23193 440 23220
rect 474 23193 513 23220
rect 547 23193 590 23223
rect 624 23193 667 23223
rect 701 23193 744 23223
rect 778 23193 821 23223
rect 855 23193 898 23223
rect 932 23193 975 23223
rect 1009 23193 1052 23223
rect 1086 23193 1129 23223
rect 1163 23193 1206 23223
rect 1240 23193 1283 23223
rect 1317 23193 1360 23223
rect 1394 23193 1437 23223
rect 348 23186 364 23193
rect 418 23186 440 23193
rect 488 23189 513 23193
rect 558 23189 590 23193
rect 211 23159 314 23186
rect 348 23159 384 23186
rect 418 23159 454 23186
rect 488 23159 524 23189
rect 558 23159 594 23189
rect 628 23159 664 23193
rect 701 23189 734 23193
rect 778 23189 804 23193
rect 855 23189 874 23193
rect 932 23189 944 23193
rect 1009 23189 1014 23193
rect 698 23159 734 23189
rect 768 23159 804 23189
rect 838 23159 874 23189
rect 908 23159 944 23189
rect 978 23159 1014 23189
rect 1048 23189 1052 23193
rect 1118 23189 1129 23193
rect 1188 23189 1206 23193
rect 1258 23189 1283 23193
rect 1328 23189 1360 23193
rect 1048 23159 1084 23189
rect 1118 23159 1154 23189
rect 1188 23159 1224 23189
rect 1258 23159 1294 23189
rect 1328 23159 1364 23189
rect 1398 23159 1434 23193
rect 1471 23189 1503 23223
rect 1468 23180 1503 23189
rect 22823 23484 23635 23514
rect 22823 23450 22827 23484
rect 22861 23475 22897 23484
rect 22876 23450 22897 23475
rect 22931 23450 22967 23484
rect 23001 23450 23037 23484
rect 23071 23450 23107 23484
rect 23141 23450 23177 23484
rect 23211 23450 23247 23484
rect 23281 23450 23317 23484
rect 23351 23450 23387 23484
rect 23421 23450 23457 23484
rect 23491 23450 23527 23484
rect 23561 23450 23597 23484
rect 23631 23450 23635 23484
rect 22823 23441 22842 23450
rect 22876 23441 23635 23450
rect 22823 23415 23635 23441
rect 22823 23381 22827 23415
rect 22861 23402 22897 23415
rect 22876 23381 22897 23402
rect 22931 23381 22967 23415
rect 23001 23381 23037 23415
rect 23071 23381 23107 23415
rect 23141 23381 23177 23415
rect 23211 23381 23247 23415
rect 23281 23381 23317 23415
rect 23351 23381 23387 23415
rect 23421 23381 23457 23415
rect 23491 23381 23527 23415
rect 23561 23381 23597 23415
rect 23631 23381 23635 23415
rect 22823 23368 22842 23381
rect 22876 23368 23635 23381
rect 22823 23346 23635 23368
rect 22823 23312 22827 23346
rect 22861 23329 22897 23346
rect 22876 23312 22897 23329
rect 22931 23312 22967 23346
rect 23001 23312 23037 23346
rect 23071 23312 23107 23346
rect 23141 23312 23177 23346
rect 23211 23312 23247 23346
rect 23281 23312 23317 23346
rect 23351 23312 23387 23346
rect 23421 23312 23457 23346
rect 23491 23312 23527 23346
rect 23561 23312 23597 23346
rect 23631 23312 23635 23346
rect 22823 23295 22842 23312
rect 22876 23295 23635 23312
rect 22823 23277 23635 23295
rect 22823 23243 22827 23277
rect 22861 23256 22897 23277
rect 22876 23243 22897 23256
rect 22931 23243 22967 23277
rect 23001 23243 23037 23277
rect 23071 23243 23107 23277
rect 23141 23243 23177 23277
rect 23211 23243 23247 23277
rect 23281 23243 23317 23277
rect 23351 23243 23387 23277
rect 23421 23243 23457 23277
rect 23491 23243 23527 23277
rect 23561 23243 23597 23277
rect 23631 23243 23635 23277
rect 22823 23222 22842 23243
rect 22876 23222 23635 23243
rect 22823 23208 23635 23222
rect 1468 23159 1502 23180
rect 211 23148 1502 23159
rect 211 23114 212 23148
rect 246 23114 288 23148
rect 322 23123 364 23148
rect 398 23123 440 23148
rect 474 23123 1502 23148
rect 348 23114 364 23123
rect 418 23114 440 23123
rect 211 23089 314 23114
rect 348 23089 384 23114
rect 418 23089 454 23114
rect 488 23089 524 23123
rect 558 23089 594 23123
rect 628 23089 664 23123
rect 698 23089 734 23123
rect 768 23089 804 23123
rect 838 23089 874 23123
rect 908 23089 944 23123
rect 978 23089 1014 23123
rect 1048 23089 1084 23123
rect 1118 23089 1154 23123
rect 1188 23089 1224 23123
rect 1258 23089 1294 23123
rect 1328 23089 1364 23123
rect 1398 23089 1434 23123
rect 1468 23089 1502 23123
rect 211 23076 1502 23089
rect 211 23042 212 23076
rect 246 23042 288 23076
rect 322 23053 364 23076
rect 398 23053 440 23076
rect 474 23053 1502 23076
rect 348 23042 364 23053
rect 418 23042 440 23053
rect 211 23019 314 23042
rect 348 23019 384 23042
rect 418 23019 454 23042
rect 488 23019 524 23053
rect 558 23019 594 23053
rect 628 23019 664 23053
rect 698 23019 734 23053
rect 768 23019 804 23053
rect 838 23019 874 23053
rect 908 23019 944 23053
rect 978 23019 1014 23053
rect 1048 23019 1084 23053
rect 1118 23019 1154 23053
rect 1188 23019 1224 23053
rect 1258 23019 1294 23053
rect 1328 23019 1364 23053
rect 1398 23019 1434 23053
rect 1468 23019 1502 23053
rect 211 23004 1502 23019
rect 211 22970 212 23004
rect 246 22970 288 23004
rect 322 22983 364 23004
rect 398 22983 440 23004
rect 474 22983 1502 23004
rect 348 22970 364 22983
rect 418 22970 440 22983
rect 211 22949 314 22970
rect 348 22949 384 22970
rect 418 22949 454 22970
rect 488 22949 524 22983
rect 558 22949 594 22983
rect 628 22949 664 22983
rect 698 22949 734 22983
rect 768 22949 804 22983
rect 838 22949 874 22983
rect 908 22949 944 22983
rect 978 22949 1014 22983
rect 1048 22949 1084 22983
rect 1118 22949 1154 22983
rect 1188 22949 1224 22983
rect 1258 22949 1294 22983
rect 1328 22949 1364 22983
rect 1398 22949 1434 22983
rect 1468 22949 1502 22983
rect 211 22932 1502 22949
rect 211 22898 212 22932
rect 246 22898 288 22932
rect 322 22913 364 22932
rect 398 22913 440 22932
rect 474 22913 1502 22932
rect 348 22898 364 22913
rect 418 22898 440 22913
rect 211 22879 314 22898
rect 348 22879 384 22898
rect 418 22879 454 22898
rect 488 22879 524 22913
rect 558 22879 594 22913
rect 628 22879 664 22913
rect 698 22879 734 22913
rect 768 22879 804 22913
rect 838 22879 874 22913
rect 908 22879 944 22913
rect 978 22879 1014 22913
rect 1048 22879 1084 22913
rect 1118 22879 1154 22913
rect 1188 22879 1224 22913
rect 1258 22879 1294 22913
rect 1328 22879 1364 22913
rect 1398 22879 1434 22913
rect 1468 22879 1502 22913
rect 211 22860 1502 22879
rect 211 22826 212 22860
rect 246 22826 288 22860
rect 322 22843 364 22860
rect 398 22843 440 22860
rect 474 22843 1502 22860
rect 348 22826 364 22843
rect 418 22826 440 22843
rect 211 22809 314 22826
rect 348 22809 384 22826
rect 418 22809 454 22826
rect 488 22809 524 22843
rect 558 22809 594 22843
rect 628 22809 664 22843
rect 698 22809 734 22843
rect 768 22809 804 22843
rect 838 22809 874 22843
rect 908 22809 944 22843
rect 978 22809 1014 22843
rect 1048 22809 1084 22843
rect 1118 22809 1154 22843
rect 1188 22809 1224 22843
rect 1258 22809 1294 22843
rect 1328 22809 1364 22843
rect 1398 22809 1434 22843
rect 1468 22809 1502 22843
rect 211 22788 1502 22809
rect 211 22754 212 22788
rect 246 22754 288 22788
rect 322 22773 364 22788
rect 398 22773 440 22788
rect 474 22773 1502 22788
rect 348 22754 364 22773
rect 418 22754 440 22773
rect 211 22739 314 22754
rect 348 22739 384 22754
rect 418 22739 454 22754
rect 488 22739 524 22773
rect 558 22739 594 22773
rect 628 22739 664 22773
rect 698 22739 734 22773
rect 768 22739 804 22773
rect 838 22739 874 22773
rect 908 22739 944 22773
rect 978 22739 1014 22773
rect 1048 22739 1084 22773
rect 1118 22739 1154 22773
rect 1188 22739 1224 22773
rect 1258 22739 1294 22773
rect 1328 22739 1364 22773
rect 1398 22739 1434 22773
rect 1468 22739 1502 22773
rect 211 22715 1502 22739
rect 211 22681 212 22715
rect 246 22681 288 22715
rect 322 22702 364 22715
rect 398 22702 440 22715
rect 474 22702 1502 22715
rect 348 22681 364 22702
rect 418 22681 440 22702
rect 211 22668 314 22681
rect 348 22668 384 22681
rect 418 22668 454 22681
rect 488 22668 524 22702
rect 558 22668 594 22702
rect 628 22668 664 22702
rect 698 22668 734 22702
rect 768 22668 804 22702
rect 838 22668 874 22702
rect 908 22668 944 22702
rect 978 22668 1014 22702
rect 1048 22668 1084 22702
rect 1118 22668 1154 22702
rect 1188 22668 1224 22702
rect 1258 22668 1294 22702
rect 1328 22668 1364 22702
rect 1398 22668 1434 22702
rect 1468 22668 1502 22702
rect 211 22642 1502 22668
rect 211 22608 212 22642
rect 246 22608 288 22642
rect 322 22631 364 22642
rect 398 22631 440 22642
rect 474 22631 1502 22642
rect 348 22608 364 22631
rect 418 22608 440 22631
rect 211 22597 314 22608
rect 348 22597 384 22608
rect 418 22597 454 22608
rect 488 22597 524 22631
rect 558 22597 594 22631
rect 628 22597 664 22631
rect 698 22597 734 22631
rect 768 22597 804 22631
rect 838 22597 874 22631
rect 908 22597 944 22631
rect 978 22597 1014 22631
rect 1048 22597 1084 22631
rect 1118 22597 1154 22631
rect 1188 22597 1224 22631
rect 1258 22597 1294 22631
rect 1328 22597 1364 22631
rect 1398 22597 1434 22631
rect 1468 22597 1502 22631
rect 211 22569 1502 22597
rect 211 22535 212 22569
rect 246 22535 288 22569
rect 322 22560 364 22569
rect 398 22560 440 22569
rect 474 22560 1502 22569
rect 348 22535 364 22560
rect 418 22535 440 22560
rect 280 22526 314 22535
rect 348 22526 384 22535
rect 418 22526 454 22535
rect 488 22526 524 22560
rect 558 22526 594 22560
rect 628 22526 664 22560
rect 698 22526 734 22560
rect 768 22526 804 22560
rect 838 22526 874 22560
rect 908 22526 944 22560
rect 978 22526 1014 22560
rect 1048 22526 1084 22560
rect 1118 22526 1154 22560
rect 1188 22526 1224 22560
rect 1258 22526 1294 22560
rect 1328 22526 1364 22560
rect 1398 22526 1434 22560
rect 1468 22526 1502 22560
rect 280 22489 1502 22526
rect 280 22455 314 22489
rect 348 22455 384 22489
rect 418 22455 454 22489
rect 488 22455 524 22489
rect 558 22455 594 22489
rect 628 22482 664 22489
rect 698 22482 734 22489
rect 628 22455 649 22482
rect 698 22455 729 22482
rect 768 22455 804 22489
rect 838 22482 874 22489
rect 908 22482 944 22489
rect 978 22482 1014 22489
rect 843 22455 874 22482
rect 923 22455 944 22482
rect 1003 22455 1014 22482
rect 1048 22482 1084 22489
rect 1048 22455 1049 22482
rect 280 22448 649 22455
rect 683 22448 729 22455
rect 763 22448 809 22455
rect 843 22448 889 22455
rect 923 22448 969 22455
rect 1003 22448 1049 22455
rect 1083 22455 1084 22482
rect 1118 22455 1154 22489
rect 1188 22455 1224 22489
rect 1258 22455 1294 22489
rect 1328 22455 1364 22489
rect 1398 22455 1434 22489
rect 1468 22455 1502 22489
rect 1083 22448 1502 22455
rect 280 22418 1502 22448
rect 280 22384 314 22418
rect 348 22384 384 22418
rect 418 22384 454 22418
rect 488 22384 524 22418
rect 558 22384 594 22418
rect 628 22410 664 22418
rect 698 22410 734 22418
rect 628 22384 649 22410
rect 698 22384 729 22410
rect 768 22384 804 22418
rect 838 22410 874 22418
rect 908 22410 944 22418
rect 978 22410 1014 22418
rect 843 22384 874 22410
rect 923 22384 944 22410
rect 1003 22384 1014 22410
rect 1048 22410 1084 22418
rect 1048 22384 1049 22410
rect 280 22376 649 22384
rect 683 22376 729 22384
rect 763 22376 809 22384
rect 843 22376 889 22384
rect 923 22376 969 22384
rect 1003 22376 1049 22384
rect 1083 22384 1084 22410
rect 1118 22384 1154 22418
rect 1188 22384 1224 22418
rect 1258 22384 1294 22418
rect 1328 22384 1364 22418
rect 1398 22384 1434 22418
rect 1468 22384 1502 22418
rect 1083 22376 1502 22384
rect 280 22347 1502 22376
rect 280 22313 314 22347
rect 348 22313 384 22347
rect 418 22313 454 22347
rect 488 22313 524 22347
rect 558 22313 594 22347
rect 628 22338 664 22347
rect 698 22338 734 22347
rect 628 22313 649 22338
rect 698 22313 729 22338
rect 768 22313 804 22347
rect 838 22338 874 22347
rect 908 22338 944 22347
rect 978 22338 1014 22347
rect 843 22313 874 22338
rect 923 22313 944 22338
rect 1003 22313 1014 22338
rect 1048 22338 1084 22347
rect 1048 22313 1049 22338
rect 280 22304 649 22313
rect 683 22304 729 22313
rect 763 22304 809 22313
rect 843 22304 889 22313
rect 923 22304 969 22313
rect 1003 22304 1049 22313
rect 1083 22313 1084 22338
rect 1118 22313 1154 22347
rect 1188 22313 1224 22347
rect 1258 22313 1294 22347
rect 1328 22313 1364 22347
rect 1398 22313 1434 22347
rect 1468 22313 1502 22347
rect 1083 22304 1502 22313
rect 280 22289 1502 22304
rect 22823 23174 22827 23208
rect 22861 23183 22897 23208
rect 22876 23174 22897 23183
rect 22931 23174 22967 23208
rect 23001 23174 23037 23208
rect 23071 23174 23107 23208
rect 23141 23174 23177 23208
rect 23211 23174 23247 23208
rect 23281 23174 23317 23208
rect 23351 23174 23387 23208
rect 23421 23174 23457 23208
rect 23491 23174 23527 23208
rect 23561 23174 23597 23208
rect 23631 23174 23635 23208
rect 22823 23149 22842 23174
rect 22876 23149 23635 23174
rect 22823 23139 23635 23149
rect 22823 23105 22827 23139
rect 22861 23110 22897 23139
rect 22876 23105 22897 23110
rect 22931 23105 22967 23139
rect 23001 23105 23037 23139
rect 23071 23105 23107 23139
rect 23141 23105 23177 23139
rect 23211 23105 23247 23139
rect 23281 23105 23317 23139
rect 23351 23105 23387 23139
rect 23421 23105 23457 23139
rect 23491 23105 23527 23139
rect 23561 23105 23597 23139
rect 23631 23105 23635 23139
rect 22823 23076 22842 23105
rect 22876 23076 23635 23105
rect 22823 23070 23635 23076
rect 22823 23036 22827 23070
rect 22861 23037 22897 23070
rect 22876 23036 22897 23037
rect 22931 23036 22967 23070
rect 23001 23036 23037 23070
rect 23071 23036 23107 23070
rect 23141 23036 23177 23070
rect 23211 23036 23247 23070
rect 23281 23036 23317 23070
rect 23351 23036 23387 23070
rect 23421 23036 23457 23070
rect 23491 23036 23527 23070
rect 23561 23036 23597 23070
rect 23631 23036 23635 23070
rect 22823 23003 22842 23036
rect 22876 23003 23635 23036
rect 22823 23001 23635 23003
rect 22823 22967 22827 23001
rect 22861 22967 22897 23001
rect 22931 22967 22967 23001
rect 23001 22967 23037 23001
rect 23071 22967 23107 23001
rect 23141 22967 23177 23001
rect 23211 22967 23247 23001
rect 23281 22967 23317 23001
rect 23351 22967 23387 23001
rect 23421 22967 23457 23001
rect 23491 22967 23527 23001
rect 23561 22967 23597 23001
rect 23631 22967 23635 23001
rect 22823 22964 23635 22967
rect 22823 22932 22842 22964
rect 22876 22932 23635 22964
rect 22823 22898 22827 22932
rect 22876 22930 22897 22932
rect 22861 22898 22897 22930
rect 22931 22898 22967 22932
rect 23001 22898 23037 22932
rect 23071 22898 23107 22932
rect 23141 22898 23177 22932
rect 23211 22898 23247 22932
rect 23281 22898 23317 22932
rect 23351 22898 23387 22932
rect 23421 22898 23457 22932
rect 23491 22898 23527 22932
rect 23561 22898 23597 22932
rect 23631 22898 23635 22932
rect 22823 22891 23635 22898
rect 22823 22863 22842 22891
rect 22876 22863 23635 22891
rect 22823 22829 22827 22863
rect 22876 22857 22897 22863
rect 22861 22829 22897 22857
rect 22931 22829 22967 22863
rect 23001 22829 23037 22863
rect 23071 22829 23107 22863
rect 23141 22829 23177 22863
rect 23211 22829 23247 22863
rect 23281 22829 23317 22863
rect 23351 22829 23387 22863
rect 23421 22829 23457 22863
rect 23491 22829 23527 22863
rect 23561 22829 23597 22863
rect 23631 22829 23635 22863
rect 22823 22818 23635 22829
rect 22823 22794 22842 22818
rect 22876 22794 23635 22818
rect 22823 22760 22827 22794
rect 22876 22784 22897 22794
rect 22861 22760 22897 22784
rect 22931 22760 22967 22794
rect 23001 22760 23037 22794
rect 23071 22760 23107 22794
rect 23141 22760 23177 22794
rect 23211 22760 23247 22794
rect 23281 22760 23317 22794
rect 23351 22760 23387 22794
rect 23421 22760 23457 22794
rect 23491 22760 23527 22794
rect 23561 22760 23597 22794
rect 23631 22760 23635 22794
rect 22823 22745 23635 22760
rect 22823 22725 22842 22745
rect 22876 22725 23635 22745
rect 22823 22691 22827 22725
rect 22876 22711 22897 22725
rect 22861 22691 22897 22711
rect 22931 22691 22967 22725
rect 23001 22691 23037 22725
rect 23071 22691 23107 22725
rect 23141 22691 23177 22725
rect 23211 22691 23247 22725
rect 23281 22691 23317 22725
rect 23351 22691 23387 22725
rect 23421 22691 23457 22725
rect 23491 22691 23527 22725
rect 23561 22691 23597 22725
rect 23631 22691 23635 22725
rect 22823 22672 23635 22691
rect 22823 22656 22842 22672
rect 22876 22656 23635 22672
rect 22823 22622 22827 22656
rect 22876 22638 22897 22656
rect 22861 22622 22897 22638
rect 22931 22622 22967 22656
rect 23001 22622 23037 22656
rect 23071 22622 23107 22656
rect 23141 22622 23177 22656
rect 23211 22622 23247 22656
rect 23281 22622 23317 22656
rect 23351 22622 23387 22656
rect 23421 22622 23457 22656
rect 23491 22622 23527 22656
rect 23561 22622 23597 22656
rect 23631 22622 23635 22656
rect 22823 22599 23635 22622
rect 22823 22587 22842 22599
rect 22876 22587 23635 22599
rect 22823 22553 22827 22587
rect 22876 22565 22897 22587
rect 22861 22553 22897 22565
rect 22931 22553 22967 22587
rect 23001 22553 23037 22587
rect 23071 22553 23107 22587
rect 23141 22553 23177 22587
rect 23211 22553 23247 22587
rect 23281 22553 23317 22587
rect 23351 22553 23387 22587
rect 23421 22553 23457 22587
rect 23491 22553 23527 22587
rect 23561 22553 23597 22587
rect 23631 22553 23635 22587
rect 22823 22526 23635 22553
rect 22823 22518 22842 22526
rect 22876 22518 23635 22526
rect 22823 22484 22827 22518
rect 22876 22492 22897 22518
rect 22861 22484 22897 22492
rect 22931 22484 22967 22518
rect 23001 22484 23037 22518
rect 23071 22484 23107 22518
rect 23141 22484 23177 22518
rect 23211 22484 23247 22518
rect 23281 22484 23317 22518
rect 23351 22484 23387 22518
rect 23421 22484 23457 22518
rect 23491 22484 23527 22518
rect 23561 22484 23597 22518
rect 23631 22484 23635 22518
rect 22823 22453 23635 22484
rect 22823 22449 22842 22453
rect 22876 22449 23635 22453
rect 22823 22415 22827 22449
rect 22876 22419 22897 22449
rect 22861 22415 22897 22419
rect 22931 22415 22967 22449
rect 23001 22415 23037 22449
rect 23071 22415 23107 22449
rect 23141 22415 23177 22449
rect 23211 22415 23247 22449
rect 23281 22415 23317 22449
rect 23351 22415 23387 22449
rect 23421 22415 23457 22449
rect 23491 22415 23527 22449
rect 23561 22415 23597 22449
rect 23631 22415 23635 22449
rect 22823 22380 23635 22415
rect 22823 22346 22827 22380
rect 22876 22346 22897 22380
rect 22931 22346 22967 22380
rect 23001 22346 23037 22380
rect 23071 22346 23107 22380
rect 23141 22346 23177 22380
rect 23211 22346 23247 22380
rect 23281 22346 23317 22380
rect 23351 22346 23387 22380
rect 23421 22346 23457 22380
rect 23491 22346 23527 22380
rect 23561 22346 23597 22380
rect 23631 22346 23635 22380
rect 22823 22311 23635 22346
rect 649 22266 1083 22289
rect 683 22232 729 22266
rect 763 22232 809 22266
rect 843 22232 889 22266
rect 923 22232 969 22266
rect 1003 22232 1049 22266
rect 649 22213 1083 22232
rect 649 22194 714 22213
rect 1020 22194 1083 22213
rect 683 22160 714 22194
rect 1020 22160 1049 22194
rect 649 22122 714 22160
rect 1020 22122 1083 22160
rect 683 22088 714 22122
rect 1020 22088 1049 22122
rect 22823 22277 22827 22311
rect 22861 22307 22897 22311
rect 22876 22277 22897 22307
rect 22931 22277 22967 22311
rect 23001 22277 23037 22311
rect 23071 22277 23107 22311
rect 23141 22277 23177 22311
rect 23211 22277 23247 22311
rect 23281 22277 23317 22311
rect 23351 22277 23387 22311
rect 23421 22277 23457 22311
rect 23491 22277 23527 22311
rect 23561 22277 23597 22311
rect 23631 22277 23635 22311
rect 22823 22273 22842 22277
rect 22876 22273 23635 22277
rect 22823 22242 23635 22273
rect 22823 22208 22827 22242
rect 22861 22234 22897 22242
rect 22876 22208 22897 22234
rect 22931 22208 22967 22242
rect 23001 22208 23037 22242
rect 23071 22208 23107 22242
rect 23141 22208 23177 22242
rect 23211 22208 23247 22242
rect 23281 22208 23317 22242
rect 23351 22208 23387 22242
rect 23421 22208 23457 22242
rect 23491 22208 23527 22242
rect 23561 22208 23597 22242
rect 23631 22208 23635 22242
rect 22823 22200 22842 22208
rect 22876 22200 23635 22208
rect 22823 22173 23635 22200
rect 22823 22139 22827 22173
rect 22861 22161 22897 22173
rect 22876 22139 22897 22161
rect 22931 22139 22967 22173
rect 23001 22139 23037 22173
rect 23071 22139 23107 22173
rect 23141 22139 23177 22173
rect 23211 22139 23247 22173
rect 23281 22139 23317 22173
rect 23351 22139 23387 22173
rect 23421 22139 23457 22173
rect 23491 22139 23527 22173
rect 23561 22139 23597 22173
rect 23631 22139 23635 22173
rect 22823 22127 22842 22139
rect 22876 22127 23635 22139
rect 22823 22115 23635 22127
rect 649 22050 714 22088
rect 1020 22050 1083 22088
rect 683 22016 714 22050
rect 1020 22016 1049 22050
rect 649 21978 714 22016
rect 1020 21978 1083 22016
rect 683 21944 714 21978
rect 1020 21944 1049 21978
rect 649 21906 714 21944
rect 1020 21906 1083 21944
rect 683 21872 714 21906
rect 1020 21872 1049 21906
rect 649 21834 714 21872
rect 1020 21834 1083 21872
rect 683 21800 714 21834
rect 1020 21800 1049 21834
rect 649 21762 714 21800
rect 1020 21762 1083 21800
rect 683 21728 714 21762
rect 1020 21728 1049 21762
rect 649 21690 714 21728
rect 1020 21690 1083 21728
rect 683 21656 714 21690
rect 1020 21656 1049 21690
rect 649 21618 714 21656
rect 1020 21618 1083 21656
rect 683 21584 714 21618
rect 1020 21584 1049 21618
rect 649 21546 714 21584
rect 1020 21546 1083 21584
rect 683 21512 714 21546
rect 1020 21512 1049 21546
rect 649 21474 714 21512
rect 1020 21474 1083 21512
rect 683 21440 714 21474
rect 1020 21440 1049 21474
rect 649 21402 714 21440
rect 1020 21402 1083 21440
rect 683 21368 714 21402
rect 1020 21368 1049 21402
rect 649 21330 714 21368
rect 1020 21330 1083 21368
rect 683 21296 714 21330
rect 1020 21296 1049 21330
rect 649 21258 714 21296
rect 1020 21258 1083 21296
rect 683 21224 714 21258
rect 1020 21224 1049 21258
rect 649 21186 714 21224
rect 1020 21186 1083 21224
rect 683 21152 714 21186
rect 1020 21152 1049 21186
rect 649 21114 714 21152
rect 1020 21114 1083 21152
rect 683 21080 714 21114
rect 1020 21080 1049 21114
rect 649 21042 714 21080
rect 1020 21042 1083 21080
rect 683 21008 714 21042
rect 1020 21008 1049 21042
rect 649 20970 714 21008
rect 1020 20970 1083 21008
rect 683 20936 714 20970
rect 1020 20936 1049 20970
rect 649 20898 714 20936
rect 1020 20898 1083 20936
rect 683 20864 714 20898
rect 1020 20864 1049 20898
rect 649 20826 714 20864
rect 1020 20826 1083 20864
rect 683 20792 714 20826
rect 1020 20792 1049 20826
rect 649 20754 714 20792
rect 1020 20754 1083 20792
rect 683 20720 714 20754
rect 1020 20720 1049 20754
rect 649 20682 714 20720
rect 1020 20682 1083 20720
rect 683 20648 714 20682
rect 1020 20648 1049 20682
rect 649 20610 714 20648
rect 1020 20610 1083 20648
rect 683 20576 714 20610
rect 1020 20576 1049 20610
rect 649 20538 714 20576
rect 1020 20538 1083 20576
rect 683 20504 714 20538
rect 1020 20504 1049 20538
rect 649 20466 714 20504
rect 1020 20466 1083 20504
rect 683 20432 714 20466
rect 1020 20432 1049 20466
rect 649 20394 714 20432
rect 1020 20394 1083 20432
rect 2335 20750 3196 20804
rect 2335 20716 2401 20750
rect 2435 20716 2474 20750
rect 2508 20716 2547 20750
rect 2581 20716 2620 20750
rect 2654 20716 2693 20750
rect 2727 20716 2766 20750
rect 2800 20716 2839 20750
rect 2873 20716 2912 20750
rect 2946 20716 2984 20750
rect 3018 20716 3056 20750
rect 3090 20716 3128 20750
rect 3162 20716 3196 20750
rect 2335 20672 3196 20716
rect 2335 20638 2401 20672
rect 2435 20638 2474 20672
rect 2508 20638 2547 20672
rect 2581 20638 2620 20672
rect 2654 20638 2693 20672
rect 2727 20638 2766 20672
rect 2800 20638 2839 20672
rect 2873 20638 2912 20672
rect 2946 20638 2984 20672
rect 3018 20638 3056 20672
rect 3090 20638 3128 20672
rect 3162 20638 3196 20672
rect 2335 20594 3196 20638
rect 2335 20560 2401 20594
rect 2435 20560 2474 20594
rect 2508 20560 2547 20594
rect 2581 20560 2620 20594
rect 2654 20560 2693 20594
rect 2727 20560 2766 20594
rect 2800 20560 2839 20594
rect 2873 20560 2912 20594
rect 2946 20560 2984 20594
rect 3018 20560 3056 20594
rect 3090 20560 3128 20594
rect 3162 20560 3196 20594
rect 2335 20538 3196 20560
rect 2335 20504 2377 20538
rect 2411 20516 2453 20538
rect 2487 20516 2529 20538
rect 2563 20516 2605 20538
rect 2639 20516 2680 20538
rect 2714 20516 2755 20538
rect 2789 20516 2830 20538
rect 2864 20516 2905 20538
rect 2939 20516 2980 20538
rect 3014 20516 3055 20538
rect 3089 20516 3130 20538
rect 2435 20504 2453 20516
rect 2508 20504 2529 20516
rect 2581 20504 2605 20516
rect 2654 20504 2680 20516
rect 2727 20504 2755 20516
rect 2800 20504 2830 20516
rect 2873 20504 2905 20516
rect 2946 20504 2980 20516
rect 3018 20504 3055 20516
rect 2335 20482 2401 20504
rect 2435 20482 2474 20504
rect 2508 20482 2547 20504
rect 2581 20482 2620 20504
rect 2654 20482 2693 20504
rect 2727 20482 2766 20504
rect 2800 20482 2839 20504
rect 2873 20482 2912 20504
rect 2946 20482 2984 20504
rect 3018 20482 3056 20504
rect 3090 20482 3128 20516
rect 3164 20504 3196 20538
rect 3162 20482 3196 20504
rect 2335 20452 3196 20482
rect 2335 20418 2377 20452
rect 2411 20438 2453 20452
rect 2487 20438 2529 20452
rect 2563 20438 2605 20452
rect 2639 20438 2680 20452
rect 2714 20438 2755 20452
rect 2789 20438 2830 20452
rect 2864 20438 2905 20452
rect 2939 20438 2980 20452
rect 3014 20438 3055 20452
rect 3089 20438 3130 20452
rect 2435 20418 2453 20438
rect 2508 20418 2529 20438
rect 2581 20418 2605 20438
rect 2654 20418 2680 20438
rect 2727 20418 2755 20438
rect 2800 20418 2830 20438
rect 2873 20418 2905 20438
rect 2946 20418 2980 20438
rect 3018 20418 3055 20438
rect 2335 20404 2401 20418
rect 2435 20404 2474 20418
rect 2508 20404 2547 20418
rect 2581 20404 2620 20418
rect 2654 20404 2693 20418
rect 2727 20404 2766 20418
rect 2800 20404 2839 20418
rect 2873 20404 2912 20418
rect 2946 20404 2984 20418
rect 3018 20404 3056 20418
rect 3090 20404 3128 20438
rect 3164 20418 3196 20452
rect 3162 20404 3196 20418
rect 26366 20718 26986 20793
rect 26366 20684 26371 20718
rect 26405 20684 26441 20718
rect 26475 20684 26511 20718
rect 26545 20684 26581 20718
rect 26615 20684 26651 20718
rect 26685 20684 26721 20718
rect 26755 20684 26791 20718
rect 26825 20684 26861 20718
rect 26895 20684 26986 20718
rect 26366 20647 26986 20684
rect 26366 20613 26371 20647
rect 26405 20613 26441 20647
rect 26475 20613 26511 20647
rect 26545 20613 26581 20647
rect 26615 20613 26651 20647
rect 26685 20613 26721 20647
rect 26755 20613 26791 20647
rect 26825 20613 26861 20647
rect 26895 20613 26986 20647
rect 26366 20576 26986 20613
rect 26366 20542 26371 20576
rect 26405 20542 26441 20576
rect 26475 20542 26511 20576
rect 26545 20542 26581 20576
rect 26615 20542 26651 20576
rect 26685 20542 26721 20576
rect 26755 20542 26791 20576
rect 26825 20542 26861 20576
rect 26895 20542 26986 20576
rect 26366 20505 26986 20542
rect 26366 20471 26371 20505
rect 26405 20471 26441 20505
rect 26475 20471 26511 20505
rect 26545 20471 26581 20505
rect 26615 20471 26651 20505
rect 26685 20471 26721 20505
rect 26755 20471 26791 20505
rect 26825 20471 26861 20505
rect 26895 20471 26986 20505
rect 26366 20439 27043 20471
rect 26366 20434 26921 20439
rect 683 20360 714 20394
rect 1020 20360 1049 20394
rect 649 20322 714 20360
rect 1020 20322 1083 20360
rect 683 20288 714 20322
rect 1020 20288 1049 20322
rect 649 20250 714 20288
rect 1020 20250 1083 20288
rect 683 20216 714 20250
rect 1020 20216 1049 20250
rect 649 20178 714 20216
rect 1020 20178 1083 20216
rect 683 20144 714 20178
rect 1020 20144 1049 20178
rect 649 20106 714 20144
rect 1020 20106 1083 20144
rect 683 20072 714 20106
rect 1020 20072 1049 20106
rect 649 20034 714 20072
rect 1020 20034 1083 20072
rect 683 20000 714 20034
rect 1020 20000 1049 20034
rect 26366 20400 26371 20434
rect 26405 20400 26441 20434
rect 26475 20400 26511 20434
rect 26545 20400 26581 20434
rect 26615 20400 26651 20434
rect 26685 20400 26721 20434
rect 26755 20400 26791 20434
rect 26825 20400 26861 20434
rect 26895 20405 26921 20434
rect 26955 20405 27003 20439
rect 27037 20405 27043 20439
rect 26895 20400 27043 20405
rect 26366 20363 27043 20400
rect 26366 20329 26371 20363
rect 26405 20329 26441 20363
rect 26475 20329 26511 20363
rect 26545 20329 26581 20363
rect 26615 20329 26651 20363
rect 26685 20329 26721 20363
rect 26755 20329 26791 20363
rect 26825 20329 26861 20363
rect 26895 20362 27043 20363
rect 26895 20329 26921 20362
rect 26366 20328 26921 20329
rect 26955 20328 27003 20362
rect 27037 20328 27043 20362
rect 26366 20296 27043 20328
rect 26366 20292 26986 20296
rect 26366 20258 26371 20292
rect 26405 20260 26441 20292
rect 26366 20226 26405 20258
rect 26439 20258 26441 20260
rect 26475 20260 26511 20292
rect 26545 20260 26581 20292
rect 26615 20260 26651 20292
rect 26685 20260 26721 20292
rect 26755 20260 26791 20292
rect 26475 20258 26481 20260
rect 26545 20258 26557 20260
rect 26615 20258 26633 20260
rect 26685 20258 26709 20260
rect 26755 20258 26785 20260
rect 26825 20258 26861 20292
rect 26895 20267 26986 20292
rect 26895 20260 27078 20267
rect 26439 20226 26481 20258
rect 26515 20226 26557 20258
rect 26591 20226 26633 20258
rect 26667 20226 26709 20258
rect 26743 20226 26785 20258
rect 26819 20226 26861 20258
rect 26895 20226 26937 20260
rect 26971 20226 27012 20260
rect 27046 20226 27078 20260
rect 26366 20221 27078 20226
rect 26366 20187 26371 20221
rect 26405 20187 26441 20221
rect 26475 20187 26511 20221
rect 26545 20187 26581 20221
rect 26615 20187 26651 20221
rect 26685 20187 26721 20221
rect 26755 20187 26791 20221
rect 26825 20187 26861 20221
rect 26895 20187 27078 20221
rect 26366 20176 27078 20187
rect 26366 20150 26405 20176
rect 26366 20116 26371 20150
rect 26439 20150 26481 20176
rect 26515 20150 26557 20176
rect 26591 20150 26633 20176
rect 26667 20150 26709 20176
rect 26743 20150 26785 20176
rect 26819 20150 26861 20176
rect 26439 20142 26441 20150
rect 26405 20116 26441 20142
rect 26475 20142 26481 20150
rect 26545 20142 26557 20150
rect 26615 20142 26633 20150
rect 26685 20142 26709 20150
rect 26755 20142 26785 20150
rect 26475 20116 26511 20142
rect 26545 20116 26581 20142
rect 26615 20116 26651 20142
rect 26685 20116 26721 20142
rect 26755 20116 26791 20142
rect 26825 20116 26861 20150
rect 26895 20142 26937 20176
rect 26971 20142 27012 20176
rect 27046 20142 27078 20176
rect 26895 20116 27078 20142
rect 26366 20092 27078 20116
rect 26366 20078 26405 20092
rect 26366 20044 26371 20078
rect 26439 20078 26481 20092
rect 26515 20078 26557 20092
rect 26591 20078 26633 20092
rect 26667 20078 26709 20092
rect 26743 20078 26785 20092
rect 26819 20078 26861 20092
rect 26439 20058 26441 20078
rect 26405 20044 26441 20058
rect 26475 20058 26481 20078
rect 26545 20058 26557 20078
rect 26615 20058 26633 20078
rect 26685 20058 26709 20078
rect 26755 20058 26785 20078
rect 26475 20044 26511 20058
rect 26545 20044 26581 20058
rect 26615 20044 26651 20058
rect 26685 20044 26721 20058
rect 26755 20044 26791 20058
rect 26825 20044 26861 20078
rect 26895 20058 26937 20092
rect 26971 20058 27012 20092
rect 27046 20058 27078 20092
rect 26895 20051 27078 20058
rect 26895 20044 26986 20051
rect 26366 20010 26986 20044
rect 649 19962 714 20000
rect 1020 19962 1083 20000
rect 683 19928 714 19962
rect 1020 19928 1049 19962
rect 649 19890 714 19928
rect 1020 19890 1083 19928
rect 683 19856 714 19890
rect 1020 19856 1049 19890
rect 649 19818 714 19856
rect 1020 19818 1083 19856
rect 683 19784 714 19818
rect 1020 19784 1049 19818
rect 649 19746 714 19784
rect 1020 19746 1083 19784
rect 683 19712 714 19746
rect 1020 19712 1049 19746
rect 649 19674 714 19712
rect 1020 19674 1083 19712
rect 683 19640 714 19674
rect 1020 19640 1049 19674
rect 649 19602 714 19640
rect 1020 19602 1083 19640
rect 683 19568 714 19602
rect 1020 19568 1049 19602
rect 649 19530 714 19568
rect 1020 19530 1083 19568
rect 683 19496 714 19530
rect 1020 19496 1049 19530
rect 649 19458 714 19496
rect 1020 19458 1083 19496
rect 683 19424 714 19458
rect 1020 19424 1049 19458
rect 649 19386 714 19424
rect 1020 19386 1083 19424
rect 683 19352 714 19386
rect 1020 19352 1049 19386
rect 649 19314 714 19352
rect 1020 19314 1083 19352
rect 683 19280 714 19314
rect 1020 19280 1049 19314
rect 649 19242 714 19280
rect 1020 19242 1083 19280
rect 683 19208 714 19242
rect 1020 19208 1049 19242
rect 649 19170 714 19208
rect 1020 19170 1083 19208
rect 683 19136 714 19170
rect 1020 19136 1049 19170
rect 649 19098 714 19136
rect 1020 19098 1083 19136
rect 683 19064 714 19098
rect 1020 19064 1049 19098
rect 649 19026 714 19064
rect 1020 19026 1083 19064
rect 683 18992 714 19026
rect 1020 18992 1049 19026
rect 649 18954 714 18992
rect 1020 18954 1083 18992
rect 683 18920 714 18954
rect 1020 18920 1049 18954
rect 649 18882 714 18920
rect 1020 18882 1083 18920
rect 683 18848 714 18882
rect 1020 18848 1049 18882
rect 649 18810 714 18848
rect 1020 18810 1083 18848
rect 683 18776 714 18810
rect 1020 18776 1049 18810
rect 649 18738 714 18776
rect 1020 18738 1083 18776
rect 683 18704 714 18738
rect 1020 18704 1049 18738
rect 649 18666 714 18704
rect 1020 18666 1083 18704
rect 683 18632 714 18666
rect 1020 18632 1049 18666
rect 649 18594 714 18632
rect 1020 18594 1083 18632
rect 683 18560 714 18594
rect 1020 18560 1049 18594
rect 649 18522 714 18560
rect 1020 18522 1083 18560
rect 683 18488 714 18522
rect 1020 18488 1049 18522
rect 649 18450 714 18488
rect 1020 18450 1083 18488
rect 683 18416 714 18450
rect 1020 18416 1049 18450
rect 649 18378 714 18416
rect 1020 18378 1083 18416
rect 683 18344 714 18378
rect 1020 18344 1049 18378
rect 649 18306 714 18344
rect 1020 18306 1083 18344
rect 683 18272 714 18306
rect 1020 18272 1049 18306
rect 649 18234 714 18272
rect 1020 18234 1083 18272
rect 683 18200 714 18234
rect 1020 18200 1049 18234
rect 649 18162 714 18200
rect 1020 18162 1083 18200
rect 683 18128 714 18162
rect 1020 18128 1049 18162
rect 649 18090 714 18128
rect 1020 18090 1083 18128
rect 683 18056 714 18090
rect 1020 18056 1049 18090
rect 649 18018 714 18056
rect 1020 18018 1083 18056
rect 683 17984 714 18018
rect 1020 17984 1049 18018
rect 649 17946 714 17984
rect 1020 17946 1083 17984
rect 683 17912 714 17946
rect 1020 17912 1049 17946
rect 649 17874 714 17912
rect 1020 17874 1083 17912
rect 683 17840 714 17874
rect 1020 17840 1049 17874
rect 649 17802 714 17840
rect 1020 17802 1083 17840
rect 683 17768 714 17802
rect 1020 17768 1049 17802
rect 649 17730 714 17768
rect 1020 17730 1083 17768
rect 683 17696 714 17730
rect 1020 17696 1049 17730
rect 649 17658 714 17696
rect 1020 17658 1083 17696
rect 683 17624 714 17658
rect 1020 17624 1049 17658
rect 649 17586 714 17624
rect 1020 17586 1083 17624
rect 683 17552 714 17586
rect 1020 17552 1049 17586
rect 649 17514 714 17552
rect 1020 17514 1083 17552
rect 683 17480 714 17514
rect 1020 17480 1049 17514
rect 649 17442 714 17480
rect 1020 17442 1083 17480
rect 683 17419 714 17442
rect 1020 17419 1049 17442
rect 683 17408 729 17419
rect 763 17408 809 17419
rect 843 17408 889 17419
rect 923 17408 969 17419
rect 1003 17408 1049 17419
rect 649 17384 1083 17408
rect 649 17370 714 17384
rect 748 17370 782 17384
rect 816 17370 850 17384
rect 683 17350 714 17370
rect 763 17350 782 17370
rect 843 17350 850 17370
rect 884 17370 918 17384
rect 952 17370 986 17384
rect 1020 17370 1083 17384
rect 884 17350 889 17370
rect 952 17350 969 17370
rect 1020 17350 1049 17370
rect 683 17336 729 17350
rect 763 17336 809 17350
rect 843 17336 889 17350
rect 923 17336 969 17350
rect 1003 17336 1049 17350
rect 649 17315 1083 17336
rect 649 17298 714 17315
rect 748 17298 782 17315
rect 816 17298 850 17315
rect 683 17281 714 17298
rect 763 17281 782 17298
rect 843 17281 850 17298
rect 884 17298 918 17315
rect 952 17298 986 17315
rect 1020 17298 1083 17315
rect 884 17281 889 17298
rect 952 17281 969 17298
rect 1020 17281 1049 17298
rect 683 17264 729 17281
rect 763 17264 809 17281
rect 843 17264 889 17281
rect 923 17264 969 17281
rect 1003 17264 1049 17281
rect 649 17246 1083 17264
rect 649 17226 714 17246
rect 748 17226 782 17246
rect 816 17226 850 17246
rect 683 17212 714 17226
rect 763 17212 782 17226
rect 843 17212 850 17226
rect 884 17226 918 17246
rect 952 17226 986 17246
rect 1020 17226 1083 17246
rect 884 17212 889 17226
rect 952 17212 969 17226
rect 1020 17212 1049 17226
rect 683 17192 729 17212
rect 763 17192 809 17212
rect 843 17192 889 17212
rect 923 17192 969 17212
rect 1003 17192 1049 17212
rect 649 17177 1083 17192
rect 649 17154 714 17177
rect 748 17154 782 17177
rect 816 17154 850 17177
rect 683 17143 714 17154
rect 763 17143 782 17154
rect 843 17143 850 17154
rect 884 17154 918 17177
rect 952 17154 986 17177
rect 1020 17154 1083 17177
rect 884 17143 889 17154
rect 952 17143 969 17154
rect 1020 17143 1049 17154
rect 683 17120 729 17143
rect 763 17120 809 17143
rect 843 17120 889 17143
rect 923 17120 969 17143
rect 1003 17120 1049 17143
rect 649 17108 1083 17120
rect 649 17082 714 17108
rect 748 17082 782 17108
rect 816 17082 850 17108
rect 683 17074 714 17082
rect 763 17074 782 17082
rect 843 17074 850 17082
rect 884 17082 918 17108
rect 952 17082 986 17108
rect 1020 17082 1083 17108
rect 884 17074 889 17082
rect 952 17074 969 17082
rect 1020 17074 1049 17082
rect 683 17048 729 17074
rect 763 17048 809 17074
rect 843 17048 889 17074
rect 923 17048 969 17074
rect 1003 17048 1049 17074
rect 649 17039 1083 17048
rect 649 17010 714 17039
rect 748 17010 782 17039
rect 816 17010 850 17039
rect 683 17005 714 17010
rect 763 17005 782 17010
rect 843 17005 850 17010
rect 884 17010 918 17039
rect 952 17010 986 17039
rect 1020 17010 1083 17039
rect 884 17005 889 17010
rect 952 17005 969 17010
rect 1020 17005 1049 17010
rect 683 16976 729 17005
rect 763 16976 809 17005
rect 843 16976 889 17005
rect 923 16976 969 17005
rect 1003 16976 1049 17005
rect 649 16970 1083 16976
rect 649 16937 714 16970
rect 748 16937 782 16970
rect 816 16937 850 16970
rect 683 16936 714 16937
rect 763 16936 782 16937
rect 843 16936 850 16937
rect 884 16937 918 16970
rect 952 16937 986 16970
rect 1020 16937 1083 16970
rect 884 16936 889 16937
rect 952 16936 969 16937
rect 1020 16936 1049 16937
rect 683 16903 729 16936
rect 763 16903 809 16936
rect 843 16903 889 16936
rect 923 16903 969 16936
rect 1003 16903 1049 16936
rect 649 16901 1083 16903
rect 649 16867 714 16901
rect 748 16867 782 16901
rect 816 16867 850 16901
rect 884 16867 918 16901
rect 952 16867 986 16901
rect 1020 16867 1083 16901
rect 649 16864 1083 16867
rect 683 16832 729 16864
rect 763 16832 809 16864
rect 843 16832 889 16864
rect 923 16832 969 16864
rect 1003 16832 1049 16864
rect 683 16830 714 16832
rect 763 16830 782 16832
rect 843 16830 850 16832
rect 649 16798 714 16830
rect 748 16798 782 16830
rect 816 16798 850 16830
rect 884 16830 889 16832
rect 952 16830 969 16832
rect 1020 16830 1049 16832
rect 884 16798 918 16830
rect 952 16798 986 16830
rect 1020 16798 1083 16830
rect 649 16791 1083 16798
rect 683 16763 729 16791
rect 763 16763 809 16791
rect 843 16763 889 16791
rect 923 16763 969 16791
rect 1003 16763 1049 16791
rect 683 16757 714 16763
rect 763 16757 782 16763
rect 843 16757 850 16763
rect 649 16729 714 16757
rect 748 16729 782 16757
rect 816 16729 850 16757
rect 884 16757 889 16763
rect 952 16757 969 16763
rect 1020 16757 1049 16763
rect 884 16729 918 16757
rect 952 16729 986 16757
rect 1020 16729 1083 16757
rect 649 16718 1083 16729
rect 683 16694 729 16718
rect 763 16694 809 16718
rect 843 16694 889 16718
rect 923 16694 969 16718
rect 1003 16694 1049 16718
rect 683 16684 714 16694
rect 763 16684 782 16694
rect 843 16684 850 16694
rect 649 16660 714 16684
rect 748 16660 782 16684
rect 816 16660 850 16684
rect 884 16684 889 16694
rect 952 16684 969 16694
rect 1020 16684 1049 16694
rect 884 16660 918 16684
rect 952 16660 986 16684
rect 1020 16660 1083 16684
rect 649 16645 1083 16660
rect 683 16625 729 16645
rect 763 16625 809 16645
rect 843 16625 889 16645
rect 923 16625 969 16645
rect 1003 16625 1049 16645
rect 683 16611 714 16625
rect 763 16611 782 16625
rect 843 16611 850 16625
rect 649 16591 714 16611
rect 748 16591 782 16611
rect 816 16591 850 16611
rect 884 16611 889 16625
rect 952 16611 969 16625
rect 1020 16611 1049 16625
rect 884 16591 918 16611
rect 952 16591 986 16611
rect 1020 16591 1083 16611
rect 649 16572 1083 16591
rect 683 16556 729 16572
rect 763 16556 809 16572
rect 843 16556 889 16572
rect 923 16556 969 16572
rect 1003 16556 1049 16572
rect 683 16538 714 16556
rect 763 16538 782 16556
rect 843 16538 850 16556
rect 649 16522 714 16538
rect 748 16522 782 16538
rect 816 16522 850 16538
rect 884 16538 889 16556
rect 952 16538 969 16556
rect 1020 16538 1049 16556
rect 3484 19551 4095 19585
rect 3484 19517 3485 19551
rect 3519 19517 3561 19551
rect 3595 19517 3637 19551
rect 3671 19517 3713 19551
rect 3747 19517 3789 19551
rect 3823 19517 3865 19551
rect 3899 19517 3941 19551
rect 3975 19517 4017 19551
rect 4051 19517 4095 19551
rect 3484 19483 4095 19517
rect 3484 19449 3485 19483
rect 3519 19449 3561 19483
rect 3595 19449 3637 19483
rect 3671 19449 3713 19483
rect 3747 19449 3789 19483
rect 3823 19449 3865 19483
rect 3899 19449 3941 19483
rect 3975 19449 4017 19483
rect 4051 19449 4095 19483
rect 3484 19415 4095 19449
rect 3484 19381 3485 19415
rect 3519 19381 3561 19415
rect 3595 19381 3637 19415
rect 3671 19381 3713 19415
rect 3747 19381 3789 19415
rect 3823 19381 3865 19415
rect 3899 19381 3941 19415
rect 3975 19381 4017 19415
rect 4051 19381 4095 19415
rect 3484 19347 4095 19381
rect 3484 19313 3485 19347
rect 3519 19313 3561 19347
rect 3595 19313 3637 19347
rect 3671 19313 3713 19347
rect 3747 19313 3789 19347
rect 3823 19313 3865 19347
rect 3899 19313 3941 19347
rect 3975 19313 4017 19347
rect 4051 19313 4095 19347
rect 3484 19279 4095 19313
rect 3484 19245 3485 19279
rect 3519 19245 3561 19279
rect 3595 19245 3637 19279
rect 3671 19245 3713 19279
rect 3747 19245 3789 19279
rect 3823 19245 3865 19279
rect 3899 19245 3941 19279
rect 3975 19245 4017 19279
rect 4051 19245 4095 19279
rect 3484 19210 4095 19245
rect 3484 19176 3485 19210
rect 3519 19176 3561 19210
rect 3595 19176 3637 19210
rect 3671 19176 3713 19210
rect 3747 19176 3789 19210
rect 3823 19176 3865 19210
rect 3899 19176 3941 19210
rect 3975 19176 4017 19210
rect 4051 19176 4095 19210
rect 3484 19141 4095 19176
rect 3484 19107 3485 19141
rect 3519 19107 3561 19141
rect 3595 19107 3637 19141
rect 3671 19107 3713 19141
rect 3747 19107 3789 19141
rect 3823 19107 3865 19141
rect 3899 19107 3941 19141
rect 3975 19107 4017 19141
rect 4051 19107 4095 19141
rect 3484 19072 4095 19107
rect 3484 19038 3485 19072
rect 3519 19038 3561 19072
rect 3595 19038 3637 19072
rect 3671 19038 3713 19072
rect 3747 19038 3789 19072
rect 3823 19038 3865 19072
rect 3899 19038 3941 19072
rect 3975 19038 4017 19072
rect 4051 19038 4095 19072
rect 3484 19003 4095 19038
rect 3484 18969 3485 19003
rect 3519 18969 3561 19003
rect 3595 18969 3637 19003
rect 3671 18969 3713 19003
rect 3747 18969 3789 19003
rect 3823 18969 3865 19003
rect 3899 18969 3941 19003
rect 3975 18969 4017 19003
rect 4051 18969 4095 19003
rect 3484 18934 4095 18969
rect 3484 18900 3485 18934
rect 3519 18900 3561 18934
rect 3595 18900 3637 18934
rect 3671 18900 3713 18934
rect 3747 18900 3789 18934
rect 3823 18900 3865 18934
rect 3899 18900 3941 18934
rect 3975 18900 4017 18934
rect 4051 18900 4095 18934
rect 3484 18865 4095 18900
rect 3484 18831 3485 18865
rect 3519 18831 3561 18865
rect 3595 18831 3637 18865
rect 3671 18831 3713 18865
rect 3747 18831 3789 18865
rect 3823 18831 3865 18865
rect 3899 18831 3941 18865
rect 3975 18831 4017 18865
rect 4051 18831 4095 18865
rect 3484 18796 4095 18831
rect 3484 18762 3485 18796
rect 3519 18762 3561 18796
rect 3595 18762 3637 18796
rect 3671 18762 3713 18796
rect 3747 18762 3789 18796
rect 3823 18762 3865 18796
rect 3899 18762 3941 18796
rect 3975 18762 4017 18796
rect 4051 18762 4095 18796
rect 3484 18727 4095 18762
rect 3484 18693 3485 18727
rect 3519 18693 3561 18727
rect 3595 18693 3637 18727
rect 3671 18693 3713 18727
rect 3747 18693 3789 18727
rect 3823 18693 3865 18727
rect 3899 18693 3941 18727
rect 3975 18693 4017 18727
rect 4051 18693 4095 18727
rect 3484 18658 4095 18693
rect 3484 18624 3485 18658
rect 3519 18624 3561 18658
rect 3595 18624 3637 18658
rect 3671 18624 3713 18658
rect 3747 18624 3789 18658
rect 3823 18624 3865 18658
rect 3899 18624 3941 18658
rect 3975 18624 4017 18658
rect 4051 18624 4095 18658
rect 3484 18589 4095 18624
rect 3484 18555 3485 18589
rect 3519 18555 3561 18589
rect 3595 18555 3637 18589
rect 3671 18555 3713 18589
rect 3747 18555 3789 18589
rect 3823 18555 3865 18589
rect 3899 18555 3941 18589
rect 3975 18555 4017 18589
rect 4051 18555 4095 18589
rect 3484 18520 4095 18555
rect 3484 18486 3485 18520
rect 3519 18486 3561 18520
rect 3595 18486 3637 18520
rect 3671 18486 3713 18520
rect 3747 18486 3789 18520
rect 3823 18486 3865 18520
rect 3899 18486 3941 18520
rect 3975 18486 4017 18520
rect 4051 18486 4095 18520
rect 3484 18451 4095 18486
rect 3484 18417 3485 18451
rect 3519 18417 3561 18451
rect 3595 18417 3637 18451
rect 3671 18417 3713 18451
rect 3747 18417 3789 18451
rect 3823 18417 3865 18451
rect 3899 18417 3941 18451
rect 3975 18417 4017 18451
rect 4051 18417 4095 18451
rect 3484 18382 4095 18417
rect 3484 18348 3485 18382
rect 3519 18348 3561 18382
rect 3595 18348 3637 18382
rect 3671 18348 3713 18382
rect 3747 18348 3789 18382
rect 3823 18348 3865 18382
rect 3899 18348 3941 18382
rect 3975 18348 4017 18382
rect 4051 18348 4095 18382
rect 3484 18313 4095 18348
rect 3484 18279 3485 18313
rect 3519 18279 3561 18313
rect 3595 18279 3637 18313
rect 3671 18279 3713 18313
rect 3747 18279 3789 18313
rect 3823 18279 3865 18313
rect 3899 18279 3941 18313
rect 3975 18279 4017 18313
rect 4051 18279 4095 18313
rect 3484 18244 4095 18279
rect 3484 18210 3485 18244
rect 3519 18210 3561 18244
rect 3595 18210 3637 18244
rect 3671 18210 3713 18244
rect 3747 18210 3789 18244
rect 3823 18210 3865 18244
rect 3899 18210 3941 18244
rect 3975 18210 4017 18244
rect 4051 18210 4095 18244
rect 3484 18175 4095 18210
rect 3484 18141 3485 18175
rect 3519 18141 3561 18175
rect 3595 18141 3637 18175
rect 3671 18141 3713 18175
rect 3747 18141 3789 18175
rect 3823 18141 3865 18175
rect 3899 18141 3941 18175
rect 3975 18141 4017 18175
rect 4051 18141 4095 18175
rect 3484 18106 4095 18141
rect 3484 18072 3485 18106
rect 3519 18072 3561 18106
rect 3595 18072 3637 18106
rect 3671 18072 3713 18106
rect 3747 18072 3789 18106
rect 3823 18072 3865 18106
rect 3899 18072 3941 18106
rect 3975 18072 4017 18106
rect 4051 18072 4095 18106
rect 3484 18037 4095 18072
rect 3484 18003 3485 18037
rect 3519 18003 3561 18037
rect 3595 18003 3637 18037
rect 3671 18003 3713 18037
rect 3747 18003 3789 18037
rect 3823 18003 3865 18037
rect 3899 18003 3941 18037
rect 3975 18003 4017 18037
rect 4051 18003 4095 18037
rect 3484 17968 4095 18003
rect 3484 17934 3485 17968
rect 3519 17934 3561 17968
rect 3595 17934 3637 17968
rect 3671 17934 3713 17968
rect 3747 17934 3789 17968
rect 3823 17934 3865 17968
rect 3899 17934 3941 17968
rect 3975 17934 4017 17968
rect 4051 17934 4095 17968
rect 3484 17899 4095 17934
rect 3484 17865 3485 17899
rect 3519 17865 3561 17899
rect 3595 17865 3637 17899
rect 3671 17865 3713 17899
rect 3747 17865 3789 17899
rect 3823 17865 3865 17899
rect 3899 17865 3941 17899
rect 3975 17865 4017 17899
rect 4051 17865 4095 17899
rect 3484 17830 4095 17865
rect 3484 17796 3485 17830
rect 3519 17796 3561 17830
rect 3595 17796 3637 17830
rect 3671 17796 3713 17830
rect 3747 17796 3789 17830
rect 3823 17796 3865 17830
rect 3899 17796 3941 17830
rect 3975 17796 4017 17830
rect 4051 17796 4095 17830
rect 3484 17761 4095 17796
rect 3484 17727 3485 17761
rect 3519 17727 3561 17761
rect 3595 17727 3637 17761
rect 3671 17727 3713 17761
rect 3747 17727 3789 17761
rect 3823 17727 3865 17761
rect 3899 17727 3941 17761
rect 3975 17727 4017 17761
rect 4051 17727 4095 17761
rect 3484 17692 4095 17727
rect 3484 17658 3485 17692
rect 3519 17658 3561 17692
rect 3595 17658 3637 17692
rect 3671 17658 3713 17692
rect 3747 17658 3789 17692
rect 3823 17658 3865 17692
rect 3899 17658 3941 17692
rect 3975 17658 4017 17692
rect 4051 17658 4095 17692
rect 3484 17623 4095 17658
rect 3484 17589 3485 17623
rect 3519 17589 3561 17623
rect 3595 17589 3637 17623
rect 3671 17589 3713 17623
rect 3747 17589 3789 17623
rect 3823 17589 3865 17623
rect 3899 17589 3941 17623
rect 3975 17589 4017 17623
rect 4051 17589 4095 17623
rect 3484 17554 4095 17589
rect 3484 17520 3485 17554
rect 3519 17520 3561 17554
rect 3595 17520 3637 17554
rect 3671 17520 3713 17554
rect 3747 17520 3789 17554
rect 3823 17520 3865 17554
rect 3899 17520 3941 17554
rect 3975 17520 4017 17554
rect 4051 17520 4095 17554
rect 3484 17485 4095 17520
rect 3484 17451 3485 17485
rect 3519 17451 3561 17485
rect 3595 17451 3637 17485
rect 3671 17451 3713 17485
rect 3747 17451 3789 17485
rect 3823 17451 3865 17485
rect 3899 17451 3941 17485
rect 3975 17451 4017 17485
rect 4051 17451 4095 17485
rect 3484 17416 4095 17451
rect 3484 17382 3485 17416
rect 3519 17382 3561 17416
rect 3595 17382 3637 17416
rect 3671 17382 3713 17416
rect 3747 17382 3789 17416
rect 3823 17382 3865 17416
rect 3899 17382 3941 17416
rect 3975 17382 4017 17416
rect 4051 17382 4095 17416
rect 3484 17347 4095 17382
rect 3484 17313 3485 17347
rect 3519 17313 3561 17347
rect 3595 17313 3637 17347
rect 3671 17313 3713 17347
rect 3747 17313 3789 17347
rect 3823 17313 3865 17347
rect 3899 17313 3941 17347
rect 3975 17313 4017 17347
rect 4051 17313 4095 17347
rect 3484 17278 4095 17313
rect 3484 17244 3485 17278
rect 3519 17244 3561 17278
rect 3595 17244 3637 17278
rect 3671 17244 3713 17278
rect 3747 17244 3789 17278
rect 3823 17244 3865 17278
rect 3899 17244 3941 17278
rect 3975 17244 4017 17278
rect 4051 17244 4095 17278
rect 3484 17209 4095 17244
rect 3484 17175 3485 17209
rect 3519 17175 3561 17209
rect 3595 17175 3637 17209
rect 3671 17175 3713 17209
rect 3747 17175 3789 17209
rect 3823 17175 3865 17209
rect 3899 17175 3941 17209
rect 3975 17175 4017 17209
rect 4051 17175 4095 17209
rect 3484 17140 4095 17175
rect 3484 17106 3485 17140
rect 3519 17106 3561 17140
rect 3595 17106 3637 17140
rect 3671 17106 3713 17140
rect 3747 17106 3789 17140
rect 3823 17106 3865 17140
rect 3899 17106 3941 17140
rect 3975 17106 4017 17140
rect 4051 17106 4095 17140
rect 3484 17047 4095 17106
rect 3484 17013 3767 17047
rect 3801 17013 3835 17047
rect 3869 17013 3903 17047
rect 3937 17013 3971 17047
rect 4005 17013 4039 17047
rect 4073 17013 4095 17047
rect 3484 16973 4095 17013
rect 3484 16939 3767 16973
rect 3801 16939 3835 16973
rect 3869 16939 3903 16973
rect 3937 16939 3971 16973
rect 4005 16939 4039 16973
rect 4073 16939 4095 16973
rect 3484 16899 4095 16939
rect 3484 16865 3767 16899
rect 3801 16865 3835 16899
rect 3869 16865 3903 16899
rect 3937 16865 3971 16899
rect 4005 16865 4039 16899
rect 4073 16865 4095 16899
rect 3484 16825 4095 16865
rect 3484 16791 3767 16825
rect 3801 16791 3835 16825
rect 3869 16791 3903 16825
rect 3937 16791 3971 16825
rect 4005 16791 4039 16825
rect 4073 16791 4095 16825
rect 3484 16751 4095 16791
rect 3484 16717 3767 16751
rect 3801 16717 3835 16751
rect 3869 16717 3903 16751
rect 3937 16717 3971 16751
rect 4005 16717 4039 16751
rect 4073 16717 4095 16751
rect 3484 16677 4095 16717
rect 3484 16643 3767 16677
rect 3801 16643 3835 16677
rect 3869 16643 3903 16677
rect 3937 16643 3971 16677
rect 4005 16643 4039 16677
rect 4073 16643 4095 16677
rect 3484 16603 4095 16643
rect 3484 16569 3767 16603
rect 3801 16569 3835 16603
rect 3869 16569 3903 16603
rect 3937 16569 3971 16603
rect 4005 16569 4039 16603
rect 4073 16569 4095 16603
rect 3484 16561 4095 16569
rect 884 16522 918 16538
rect 952 16522 986 16538
rect 1020 16522 1083 16538
rect 649 16499 1083 16522
rect 683 16487 729 16499
rect 763 16487 809 16499
rect 843 16487 889 16499
rect 923 16487 969 16499
rect 1003 16487 1049 16499
rect 683 16465 714 16487
rect 763 16465 782 16487
rect 843 16465 850 16487
rect 649 16453 714 16465
rect 748 16453 782 16465
rect 816 16453 850 16465
rect 884 16465 889 16487
rect 952 16465 969 16487
rect 1020 16465 1049 16487
rect 884 16453 918 16465
rect 952 16453 986 16465
rect 1020 16453 1083 16465
rect 649 16426 1083 16453
rect 3451 16527 3493 16561
rect 3527 16527 3569 16561
rect 3603 16529 4095 16561
rect 3603 16527 3767 16529
rect 3417 16495 3767 16527
rect 3801 16495 3835 16529
rect 3869 16495 3903 16529
rect 3937 16495 3971 16529
rect 4005 16495 4039 16529
rect 4073 16495 4095 16529
rect 3417 16483 4095 16495
rect 3451 16449 3493 16483
rect 3527 16449 3569 16483
rect 3603 16455 4095 16483
rect 3603 16449 3767 16455
rect 683 16418 729 16426
rect 763 16418 809 16426
rect 843 16418 889 16426
rect 923 16418 969 16426
rect 1003 16418 1049 16426
rect 683 16392 714 16418
rect 763 16392 782 16418
rect 843 16392 850 16418
rect 748 16384 782 16392
rect 816 16384 850 16392
rect 884 16392 889 16418
rect 952 16392 969 16418
rect 1020 16392 1049 16418
rect 3484 16421 3767 16449
rect 3801 16421 3835 16455
rect 3869 16421 3903 16455
rect 3937 16421 3971 16455
rect 4005 16421 4039 16455
rect 4073 16421 4095 16455
rect 884 16384 918 16392
rect 952 16384 986 16392
rect 714 16349 1020 16384
rect 748 16315 782 16349
rect 816 16315 850 16349
rect 884 16315 918 16349
rect 952 16315 986 16349
rect 714 16280 1020 16315
rect 3484 16380 4095 16421
rect 3484 16346 3767 16380
rect 3801 16346 3835 16380
rect 3869 16346 3903 16380
rect 3937 16346 3971 16380
rect 4005 16346 4039 16380
rect 4073 16346 4095 16380
rect 3484 16312 4095 16346
rect 3484 16294 3732 16312
rect 748 16246 782 16280
rect 816 16246 850 16280
rect 884 16246 918 16280
rect 952 16246 986 16280
rect 714 16222 1020 16246
rect 2950 16260 3732 16294
rect 2984 16226 3018 16260
rect 3052 16226 3086 16260
rect 3120 16226 3154 16260
rect 3188 16226 3222 16260
rect 3256 16226 3290 16260
rect 3324 16226 3358 16260
rect 3392 16226 3426 16260
rect 3460 16226 3494 16260
rect 3528 16226 3562 16260
rect 3596 16226 3630 16260
rect 3664 16226 3698 16260
rect 2950 16188 3732 16226
rect 2984 16154 3018 16188
rect 3052 16154 3086 16188
rect 3120 16154 3154 16188
rect 3188 16154 3222 16188
rect 3256 16154 3290 16188
rect 3324 16154 3358 16188
rect 3392 16154 3426 16188
rect 3460 16154 3494 16188
rect 3528 16154 3562 16188
rect 3596 16154 3630 16188
rect 3664 16154 3698 16188
rect 2950 16116 3732 16154
rect 2984 16082 3018 16116
rect 3052 16082 3086 16116
rect 3120 16082 3154 16116
rect 3188 16082 3222 16116
rect 3256 16082 3290 16116
rect 3324 16082 3358 16116
rect 3392 16082 3426 16116
rect 3460 16082 3494 16116
rect 3528 16082 3562 16116
rect 3596 16082 3630 16116
rect 3664 16082 3698 16116
rect 2950 16044 3732 16082
rect 2984 16010 3018 16044
rect 3052 16010 3086 16044
rect 3120 16010 3154 16044
rect 3188 16010 3222 16044
rect 3256 16010 3290 16044
rect 3324 16010 3358 16044
rect 3392 16010 3426 16044
rect 3460 16010 3494 16044
rect 3528 16010 3562 16044
rect 3596 16010 3630 16044
rect 3664 16010 3698 16044
rect 2950 15972 3732 16010
rect 2984 15938 3018 15972
rect 3052 15938 3086 15972
rect 3120 15938 3154 15972
rect 3188 15938 3222 15972
rect 3256 15938 3290 15972
rect 3324 15938 3358 15972
rect 3392 15938 3426 15972
rect 3460 15938 3494 15972
rect 3528 15938 3562 15972
rect 3596 15938 3630 15972
rect 3664 15938 3698 15972
rect 2950 15900 3732 15938
rect 2984 15866 3018 15900
rect 3052 15866 3086 15900
rect 3120 15866 3154 15900
rect 3188 15866 3222 15900
rect 3256 15866 3290 15900
rect 3324 15866 3358 15900
rect 3392 15866 3426 15900
rect 3460 15866 3494 15900
rect 3528 15866 3562 15900
rect 3596 15866 3630 15900
rect 3664 15866 3698 15900
rect 2950 15828 3732 15866
rect 2984 15794 3018 15828
rect 3052 15794 3086 15828
rect 3120 15794 3154 15828
rect 3188 15794 3222 15828
rect 3256 15794 3290 15828
rect 3324 15794 3358 15828
rect 3392 15794 3426 15828
rect 3460 15794 3494 15828
rect 3528 15794 3562 15828
rect 3596 15794 3630 15828
rect 3664 15794 3698 15828
rect 2950 15756 3732 15794
rect 2984 15722 3018 15756
rect 3052 15722 3086 15756
rect 3120 15722 3154 15756
rect 3188 15722 3222 15756
rect 3256 15722 3290 15756
rect 3324 15722 3358 15756
rect 3392 15722 3426 15756
rect 3460 15722 3494 15756
rect 3528 15722 3562 15756
rect 3596 15722 3630 15756
rect 3664 15722 3698 15756
rect 2950 15684 3732 15722
rect 2984 15650 3018 15684
rect 3052 15650 3086 15684
rect 3120 15650 3154 15684
rect 3188 15650 3222 15684
rect 3256 15650 3290 15684
rect 3324 15650 3358 15684
rect 3392 15650 3426 15684
rect 3460 15650 3494 15684
rect 3528 15650 3562 15684
rect 3596 15650 3630 15684
rect 3664 15650 3698 15684
rect 2950 15612 3732 15650
rect 2984 15578 3018 15612
rect 3052 15578 3086 15612
rect 3120 15578 3154 15612
rect 3188 15578 3222 15612
rect 3256 15578 3290 15612
rect 3324 15578 3358 15612
rect 3392 15578 3426 15612
rect 3460 15578 3494 15612
rect 3528 15578 3562 15612
rect 3596 15578 3630 15612
rect 3664 15578 3698 15612
rect 2950 15540 3732 15578
rect 2984 15506 3018 15540
rect 3052 15506 3086 15540
rect 3120 15506 3154 15540
rect 3188 15506 3222 15540
rect 3256 15506 3290 15540
rect 3324 15506 3358 15540
rect 3392 15506 3426 15540
rect 3460 15506 3494 15540
rect 3528 15506 3562 15540
rect 3596 15506 3630 15540
rect 3664 15506 3698 15540
rect 2950 15468 3732 15506
rect 2984 15434 3018 15468
rect 3052 15434 3086 15468
rect 3120 15434 3154 15468
rect 3188 15434 3222 15468
rect 3256 15434 3290 15468
rect 3324 15434 3358 15468
rect 3392 15434 3426 15468
rect 3460 15434 3494 15468
rect 3528 15434 3562 15468
rect 3596 15434 3630 15468
rect 3664 15434 3698 15468
rect 2950 15400 3732 15434
rect 7855 16278 8275 16312
rect 7855 16244 7858 16278
rect 7892 16244 7934 16278
rect 7968 16244 8010 16278
rect 8044 16272 8086 16278
rect 8072 16244 8086 16272
rect 8120 16272 8162 16278
rect 8120 16244 8138 16272
rect 8196 16244 8238 16278
rect 7855 16238 8038 16244
rect 8072 16238 8138 16244
rect 8172 16238 8238 16244
rect 8272 16238 8275 16278
rect 7855 16209 8275 16238
rect 7855 16175 7858 16209
rect 7892 16175 7934 16209
rect 7968 16175 8010 16209
rect 8044 16189 8086 16209
rect 8072 16175 8086 16189
rect 8120 16189 8162 16209
rect 8120 16175 8138 16189
rect 8196 16175 8238 16209
rect 7855 16155 8038 16175
rect 8072 16155 8138 16175
rect 8172 16155 8238 16175
rect 8272 16155 8275 16209
rect 7855 16140 8275 16155
rect 7855 16106 7858 16140
rect 7892 16106 7934 16140
rect 7968 16106 8010 16140
rect 8044 16106 8086 16140
rect 8120 16106 8162 16140
rect 8196 16106 8238 16140
rect 7855 16072 8038 16106
rect 8072 16072 8138 16106
rect 8172 16072 8238 16106
rect 8272 16072 8275 16140
rect 7855 16071 8275 16072
rect 7855 16037 7858 16071
rect 7892 16037 7934 16071
rect 7968 16037 8010 16071
rect 8044 16037 8086 16071
rect 8120 16037 8162 16071
rect 8196 16037 8238 16071
rect 8272 16037 8275 16071
rect 7855 16023 8275 16037
rect 7855 16002 8038 16023
rect 8072 16002 8138 16023
rect 8172 16002 8238 16023
rect 7855 15968 7858 16002
rect 7892 15968 7934 16002
rect 7968 15968 8010 16002
rect 8072 15989 8086 16002
rect 8044 15968 8086 15989
rect 8120 15989 8138 16002
rect 8120 15968 8162 15989
rect 8196 15968 8238 16002
rect 8272 15968 8275 16023
rect 7855 15939 8275 15968
rect 7855 15933 8038 15939
rect 8072 15933 8138 15939
rect 8172 15933 8238 15939
rect 7855 15899 7858 15933
rect 7892 15899 7934 15933
rect 7968 15899 8010 15933
rect 8072 15905 8086 15933
rect 8044 15899 8086 15905
rect 8120 15905 8138 15933
rect 8120 15899 8162 15905
rect 8196 15899 8238 15933
rect 8272 15899 8275 15939
rect 7855 15864 8275 15899
rect 7855 15830 7858 15864
rect 7892 15830 7934 15864
rect 7968 15830 8010 15864
rect 8044 15855 8086 15864
rect 8072 15830 8086 15855
rect 8120 15855 8162 15864
rect 8120 15830 8138 15855
rect 8196 15830 8238 15864
rect 7855 15821 8038 15830
rect 8072 15821 8138 15830
rect 8172 15821 8238 15830
rect 8272 15821 8275 15864
rect 7855 15795 8275 15821
rect 7855 15761 7858 15795
rect 7892 15761 7934 15795
rect 7968 15761 8010 15795
rect 8044 15761 8086 15795
rect 8120 15761 8162 15795
rect 8196 15761 8238 15795
rect 8272 15761 8275 15795
rect 7855 15726 8275 15761
rect 7855 15692 7858 15726
rect 7892 15692 7934 15726
rect 7968 15692 8010 15726
rect 8044 15692 8086 15726
rect 8120 15692 8162 15726
rect 8196 15692 8238 15726
rect 8272 15692 8275 15726
rect 7855 15657 8275 15692
rect 7855 15623 7858 15657
rect 7892 15623 7934 15657
rect 7968 15623 8010 15657
rect 8044 15623 8086 15657
rect 8120 15623 8162 15657
rect 8196 15623 8238 15657
rect 8272 15623 8275 15657
rect 7855 15588 8275 15623
rect 7855 15554 7858 15588
rect 7892 15554 7934 15588
rect 7968 15554 8010 15588
rect 8044 15554 8086 15588
rect 8120 15554 8162 15588
rect 8196 15554 8238 15588
rect 8272 15554 8275 15588
rect 7855 15519 8275 15554
rect 7855 15485 7858 15519
rect 7892 15485 7934 15519
rect 7968 15485 8010 15519
rect 8044 15485 8086 15519
rect 8120 15485 8162 15519
rect 8196 15485 8238 15519
rect 8272 15485 8275 15519
rect 7855 15449 8275 15485
rect 7855 15415 7858 15449
rect 7892 15415 7934 15449
rect 7968 15415 8010 15449
rect 8044 15415 8086 15449
rect 8120 15415 8162 15449
rect 8196 15415 8238 15449
rect 8272 15415 8275 15449
rect 7855 15381 8275 15415
rect 226 12948 1226 12972
rect 226 12914 233 12948
rect 267 12940 301 12948
rect 335 12940 369 12948
rect 403 12940 437 12948
rect 471 12940 505 12948
rect 269 12914 301 12940
rect 347 12914 369 12940
rect 425 12914 437 12940
rect 503 12914 505 12940
rect 539 12940 573 12948
rect 607 12940 641 12948
rect 539 12914 547 12940
rect 607 12914 625 12940
rect 675 12914 709 12948
rect 743 12914 777 12948
rect 811 12914 845 12948
rect 879 12914 913 12948
rect 947 12914 981 12948
rect 1015 12914 1049 12948
rect 1083 12914 1117 12948
rect 1151 12914 1185 12948
rect 1219 12914 1226 12948
rect 226 12906 235 12914
rect 269 12906 313 12914
rect 347 12906 391 12914
rect 425 12906 469 12914
rect 503 12906 547 12914
rect 581 12906 625 12914
rect 659 12906 1226 12914
rect 226 12877 1226 12906
rect 226 12843 233 12877
rect 267 12868 301 12877
rect 335 12868 369 12877
rect 403 12868 437 12877
rect 471 12868 505 12877
rect 269 12843 301 12868
rect 347 12843 369 12868
rect 425 12843 437 12868
rect 503 12843 505 12868
rect 539 12868 573 12877
rect 607 12868 641 12877
rect 539 12843 547 12868
rect 607 12843 625 12868
rect 675 12843 709 12877
rect 743 12843 777 12877
rect 811 12843 845 12877
rect 879 12843 913 12877
rect 947 12843 981 12877
rect 1015 12843 1049 12877
rect 1083 12843 1117 12877
rect 1151 12843 1185 12877
rect 1219 12843 1226 12877
rect 226 12834 235 12843
rect 269 12834 313 12843
rect 347 12834 391 12843
rect 425 12834 469 12843
rect 503 12834 547 12843
rect 581 12834 625 12843
rect 659 12834 1226 12843
rect 226 12806 1226 12834
rect 226 12772 233 12806
rect 267 12796 301 12806
rect 335 12796 369 12806
rect 403 12796 437 12806
rect 471 12796 505 12806
rect 269 12772 301 12796
rect 347 12772 369 12796
rect 425 12772 437 12796
rect 503 12772 505 12796
rect 539 12796 573 12806
rect 607 12796 641 12806
rect 539 12772 547 12796
rect 607 12772 625 12796
rect 675 12772 709 12806
rect 743 12772 777 12806
rect 811 12772 845 12806
rect 879 12772 913 12806
rect 947 12772 981 12806
rect 1015 12772 1049 12806
rect 1083 12772 1117 12806
rect 1151 12772 1185 12806
rect 1219 12772 1226 12806
rect 226 12762 235 12772
rect 269 12762 313 12772
rect 347 12762 391 12772
rect 425 12762 469 12772
rect 503 12762 547 12772
rect 581 12762 625 12772
rect 659 12762 1226 12772
rect 226 12735 1226 12762
rect 226 12701 233 12735
rect 267 12724 301 12735
rect 335 12724 369 12735
rect 403 12724 437 12735
rect 471 12724 505 12735
rect 269 12701 301 12724
rect 347 12701 369 12724
rect 425 12701 437 12724
rect 503 12701 505 12724
rect 539 12724 573 12735
rect 607 12724 641 12735
rect 539 12701 547 12724
rect 607 12701 625 12724
rect 675 12701 709 12735
rect 743 12701 777 12735
rect 811 12701 845 12735
rect 879 12701 913 12735
rect 947 12701 981 12735
rect 1015 12701 1049 12735
rect 1083 12701 1117 12735
rect 1151 12701 1185 12735
rect 1219 12701 1226 12735
rect 226 12690 235 12701
rect 269 12690 313 12701
rect 347 12690 391 12701
rect 425 12690 469 12701
rect 503 12690 547 12701
rect 581 12690 625 12701
rect 659 12690 1226 12701
rect 226 12664 1226 12690
rect 226 12630 233 12664
rect 267 12652 301 12664
rect 335 12652 369 12664
rect 403 12652 437 12664
rect 471 12652 505 12664
rect 269 12630 301 12652
rect 347 12630 369 12652
rect 425 12630 437 12652
rect 503 12630 505 12652
rect 539 12652 573 12664
rect 607 12652 641 12664
rect 539 12630 547 12652
rect 607 12630 625 12652
rect 675 12630 709 12664
rect 743 12630 777 12664
rect 811 12630 845 12664
rect 879 12630 913 12664
rect 947 12630 981 12664
rect 1015 12630 1049 12664
rect 1083 12630 1117 12664
rect 1151 12630 1185 12664
rect 1219 12630 1226 12664
rect 226 12618 235 12630
rect 269 12618 313 12630
rect 347 12618 391 12630
rect 425 12618 469 12630
rect 503 12618 547 12630
rect 581 12618 625 12630
rect 659 12618 1226 12630
rect 226 12593 1226 12618
rect 226 12559 233 12593
rect 267 12579 301 12593
rect 335 12579 369 12593
rect 403 12579 437 12593
rect 471 12579 505 12593
rect 269 12559 301 12579
rect 347 12559 369 12579
rect 425 12559 437 12579
rect 503 12559 505 12579
rect 539 12579 573 12593
rect 607 12579 641 12593
rect 539 12559 547 12579
rect 607 12559 625 12579
rect 675 12559 709 12593
rect 743 12559 777 12593
rect 811 12559 845 12593
rect 879 12559 913 12593
rect 947 12559 981 12593
rect 1015 12559 1049 12593
rect 1083 12559 1117 12593
rect 1151 12559 1185 12593
rect 1219 12559 1226 12593
rect 226 12545 235 12559
rect 269 12545 313 12559
rect 347 12545 391 12559
rect 425 12545 469 12559
rect 503 12545 547 12559
rect 581 12545 625 12559
rect 659 12545 1226 12559
rect 226 12522 1226 12545
rect 226 12488 233 12522
rect 267 12506 301 12522
rect 335 12506 369 12522
rect 403 12506 437 12522
rect 471 12506 505 12522
rect 269 12488 301 12506
rect 347 12488 369 12506
rect 425 12488 437 12506
rect 503 12488 505 12506
rect 539 12506 573 12522
rect 607 12506 641 12522
rect 539 12488 547 12506
rect 607 12488 625 12506
rect 675 12488 709 12522
rect 743 12488 777 12522
rect 811 12488 845 12522
rect 879 12488 913 12522
rect 947 12488 981 12522
rect 1015 12488 1049 12522
rect 1083 12488 1117 12522
rect 1151 12488 1185 12522
rect 1219 12488 1226 12522
rect 226 12472 235 12488
rect 269 12472 313 12488
rect 347 12472 391 12488
rect 425 12472 469 12488
rect 503 12472 547 12488
rect 581 12472 625 12488
rect 659 12472 1226 12488
rect 226 12451 1226 12472
rect 226 12417 233 12451
rect 267 12417 301 12451
rect 335 12417 369 12451
rect 403 12417 437 12451
rect 471 12417 505 12451
rect 539 12417 573 12451
rect 607 12417 641 12451
rect 675 12417 709 12451
rect 743 12417 777 12451
rect 811 12417 845 12451
rect 879 12417 913 12451
rect 947 12417 981 12451
rect 1015 12417 1049 12451
rect 1083 12417 1117 12451
rect 1151 12417 1185 12451
rect 1219 12417 1226 12451
rect 226 12413 1226 12417
rect 226 12380 236 12413
rect 270 12380 309 12413
rect 343 12380 382 12413
rect 416 12380 455 12413
rect 489 12380 527 12413
rect 561 12380 599 12413
rect 633 12380 671 12413
rect 705 12380 743 12413
rect 226 12346 233 12380
rect 270 12379 301 12380
rect 343 12379 369 12380
rect 416 12379 437 12380
rect 489 12379 505 12380
rect 561 12379 573 12380
rect 633 12379 641 12380
rect 705 12379 709 12380
rect 267 12346 301 12379
rect 335 12346 369 12379
rect 403 12346 437 12379
rect 471 12346 505 12379
rect 539 12346 573 12379
rect 607 12346 641 12379
rect 675 12346 709 12379
rect 777 12380 815 12413
rect 849 12380 887 12413
rect 921 12380 959 12413
rect 993 12380 1031 12413
rect 1065 12380 1103 12413
rect 1137 12380 1175 12413
rect 1209 12380 1226 12413
rect 743 12346 777 12379
rect 811 12379 815 12380
rect 879 12379 887 12380
rect 947 12379 959 12380
rect 1015 12379 1031 12380
rect 1083 12379 1103 12380
rect 1151 12379 1175 12380
rect 811 12346 845 12379
rect 879 12346 913 12379
rect 947 12346 981 12379
rect 1015 12346 1049 12379
rect 1083 12346 1117 12379
rect 1151 12346 1185 12379
rect 1219 12346 1226 12380
rect 226 12339 1226 12346
rect 226 12309 236 12339
rect 270 12309 309 12339
rect 343 12309 382 12339
rect 416 12309 455 12339
rect 489 12309 527 12339
rect 561 12309 599 12339
rect 633 12309 671 12339
rect 705 12309 743 12339
rect 226 12275 233 12309
rect 270 12305 301 12309
rect 343 12305 369 12309
rect 416 12305 437 12309
rect 489 12305 505 12309
rect 561 12305 573 12309
rect 633 12305 641 12309
rect 705 12305 709 12309
rect 267 12275 301 12305
rect 335 12275 369 12305
rect 403 12275 437 12305
rect 471 12275 505 12305
rect 539 12275 573 12305
rect 607 12275 641 12305
rect 675 12275 709 12305
rect 777 12309 815 12339
rect 849 12309 887 12339
rect 921 12309 959 12339
rect 993 12309 1031 12339
rect 1065 12309 1103 12339
rect 1137 12309 1175 12339
rect 1209 12309 1226 12339
rect 743 12275 777 12305
rect 811 12305 815 12309
rect 879 12305 887 12309
rect 947 12305 959 12309
rect 1015 12305 1031 12309
rect 1083 12305 1103 12309
rect 1151 12305 1175 12309
rect 811 12275 845 12305
rect 879 12275 913 12305
rect 947 12275 981 12305
rect 1015 12275 1049 12305
rect 1083 12275 1117 12305
rect 1151 12275 1185 12305
rect 1219 12275 1226 12309
rect 226 12265 1226 12275
rect 226 12238 236 12265
rect 270 12238 309 12265
rect 343 12238 382 12265
rect 416 12238 455 12265
rect 489 12238 527 12265
rect 561 12238 599 12265
rect 633 12238 671 12265
rect 705 12238 743 12265
rect 226 12204 233 12238
rect 270 12231 301 12238
rect 343 12231 369 12238
rect 416 12231 437 12238
rect 489 12231 505 12238
rect 561 12231 573 12238
rect 633 12231 641 12238
rect 705 12231 709 12238
rect 267 12204 301 12231
rect 335 12204 369 12231
rect 403 12204 437 12231
rect 471 12204 505 12231
rect 539 12204 573 12231
rect 607 12204 641 12231
rect 675 12204 709 12231
rect 777 12238 815 12265
rect 849 12238 887 12265
rect 921 12238 959 12265
rect 993 12238 1031 12265
rect 1065 12238 1103 12265
rect 1137 12238 1175 12265
rect 1209 12238 1226 12265
rect 743 12204 777 12231
rect 811 12231 815 12238
rect 879 12231 887 12238
rect 947 12231 959 12238
rect 1015 12231 1031 12238
rect 1083 12231 1103 12238
rect 1151 12231 1175 12238
rect 811 12204 845 12231
rect 879 12204 913 12231
rect 947 12204 981 12231
rect 1015 12204 1049 12231
rect 1083 12204 1117 12231
rect 1151 12204 1185 12231
rect 1219 12204 1226 12238
rect 226 12191 1226 12204
rect 226 12167 236 12191
rect 270 12167 309 12191
rect 343 12167 382 12191
rect 416 12167 455 12191
rect 489 12167 527 12191
rect 561 12167 599 12191
rect 633 12167 671 12191
rect 705 12167 743 12191
rect 226 12133 233 12167
rect 270 12157 301 12167
rect 343 12157 369 12167
rect 416 12157 437 12167
rect 489 12157 505 12167
rect 561 12157 573 12167
rect 633 12157 641 12167
rect 705 12157 709 12167
rect 267 12133 301 12157
rect 335 12133 369 12157
rect 403 12133 437 12157
rect 471 12133 505 12157
rect 539 12133 573 12157
rect 607 12133 641 12157
rect 675 12133 709 12157
rect 777 12167 815 12191
rect 849 12167 887 12191
rect 921 12167 959 12191
rect 993 12167 1031 12191
rect 1065 12167 1103 12191
rect 1137 12167 1175 12191
rect 1209 12167 1226 12191
rect 743 12133 777 12157
rect 811 12157 815 12167
rect 879 12157 887 12167
rect 947 12157 959 12167
rect 1015 12157 1031 12167
rect 1083 12157 1103 12167
rect 1151 12157 1175 12167
rect 811 12133 845 12157
rect 879 12133 913 12157
rect 947 12133 981 12157
rect 1015 12133 1049 12157
rect 1083 12133 1117 12157
rect 1151 12133 1185 12157
rect 1219 12133 1226 12167
rect 226 12117 1226 12133
rect 226 12096 236 12117
rect 270 12096 309 12117
rect 343 12096 382 12117
rect 416 12096 455 12117
rect 489 12096 527 12117
rect 561 12096 599 12117
rect 633 12096 671 12117
rect 705 12096 743 12117
rect 226 12062 233 12096
rect 270 12083 301 12096
rect 343 12083 369 12096
rect 416 12083 437 12096
rect 489 12083 505 12096
rect 561 12083 573 12096
rect 633 12083 641 12096
rect 705 12083 709 12096
rect 267 12062 301 12083
rect 335 12062 369 12083
rect 403 12062 437 12083
rect 471 12062 505 12083
rect 539 12062 573 12083
rect 607 12062 641 12083
rect 675 12062 709 12083
rect 777 12096 815 12117
rect 849 12096 887 12117
rect 921 12096 959 12117
rect 993 12096 1031 12117
rect 1065 12096 1103 12117
rect 1137 12096 1175 12117
rect 1209 12096 1226 12117
rect 743 12062 777 12083
rect 811 12083 815 12096
rect 879 12083 887 12096
rect 947 12083 959 12096
rect 1015 12083 1031 12096
rect 1083 12083 1103 12096
rect 1151 12083 1175 12096
rect 811 12062 845 12083
rect 879 12062 913 12083
rect 947 12062 981 12083
rect 1015 12062 1049 12083
rect 1083 12062 1117 12083
rect 1151 12062 1185 12083
rect 1219 12062 1226 12096
rect 226 12043 1226 12062
rect 226 12025 236 12043
rect 270 12025 309 12043
rect 343 12025 382 12043
rect 416 12025 455 12043
rect 489 12025 527 12043
rect 561 12025 599 12043
rect 633 12025 671 12043
rect 705 12025 743 12043
rect 226 11991 233 12025
rect 270 12009 301 12025
rect 343 12009 369 12025
rect 416 12009 437 12025
rect 489 12009 505 12025
rect 561 12009 573 12025
rect 633 12009 641 12025
rect 705 12009 709 12025
rect 267 11991 301 12009
rect 335 11991 369 12009
rect 403 11991 437 12009
rect 471 11991 505 12009
rect 539 11991 573 12009
rect 607 11991 641 12009
rect 675 11991 709 12009
rect 777 12025 815 12043
rect 849 12025 887 12043
rect 921 12025 959 12043
rect 993 12025 1031 12043
rect 1065 12025 1103 12043
rect 1137 12025 1175 12043
rect 1209 12025 1226 12043
rect 743 11991 777 12009
rect 811 12009 815 12025
rect 879 12009 887 12025
rect 947 12009 959 12025
rect 1015 12009 1031 12025
rect 1083 12009 1103 12025
rect 1151 12009 1175 12025
rect 811 11991 845 12009
rect 879 11991 913 12009
rect 947 11991 981 12009
rect 1015 11991 1049 12009
rect 1083 11991 1117 12009
rect 1151 11991 1185 12009
rect 1219 11991 1226 12025
rect 226 11969 1226 11991
rect 226 11954 236 11969
rect 270 11954 309 11969
rect 343 11954 382 11969
rect 416 11954 455 11969
rect 489 11954 527 11969
rect 561 11954 599 11969
rect 633 11954 671 11969
rect 705 11954 743 11969
rect 226 11920 233 11954
rect 270 11935 301 11954
rect 343 11935 369 11954
rect 416 11935 437 11954
rect 489 11935 505 11954
rect 561 11935 573 11954
rect 633 11935 641 11954
rect 705 11935 709 11954
rect 267 11920 301 11935
rect 335 11920 369 11935
rect 403 11920 437 11935
rect 471 11920 505 11935
rect 539 11920 573 11935
rect 607 11920 641 11935
rect 675 11920 709 11935
rect 777 11954 815 11969
rect 849 11954 887 11969
rect 921 11954 959 11969
rect 993 11954 1031 11969
rect 1065 11954 1103 11969
rect 1137 11954 1175 11969
rect 1209 11954 1226 11969
rect 743 11920 777 11935
rect 811 11935 815 11954
rect 879 11935 887 11954
rect 947 11935 959 11954
rect 1015 11935 1031 11954
rect 1083 11935 1103 11954
rect 1151 11935 1175 11954
rect 811 11920 845 11935
rect 879 11920 913 11935
rect 947 11920 981 11935
rect 1015 11920 1049 11935
rect 1083 11920 1117 11935
rect 1151 11920 1185 11935
rect 1219 11920 1226 11954
rect 226 11895 1226 11920
rect 226 11883 236 11895
rect 270 11883 309 11895
rect 343 11883 382 11895
rect 416 11883 455 11895
rect 489 11883 527 11895
rect 561 11883 599 11895
rect 633 11883 671 11895
rect 705 11883 743 11895
rect 226 11849 233 11883
rect 270 11861 301 11883
rect 343 11861 369 11883
rect 416 11861 437 11883
rect 489 11861 505 11883
rect 561 11861 573 11883
rect 633 11861 641 11883
rect 705 11861 709 11883
rect 267 11849 301 11861
rect 335 11849 369 11861
rect 403 11849 437 11861
rect 471 11849 505 11861
rect 539 11849 573 11861
rect 607 11849 641 11861
rect 675 11849 709 11861
rect 777 11883 815 11895
rect 849 11883 887 11895
rect 921 11883 959 11895
rect 993 11883 1031 11895
rect 1065 11883 1103 11895
rect 1137 11883 1175 11895
rect 1209 11883 1226 11895
rect 743 11849 777 11861
rect 811 11861 815 11883
rect 879 11861 887 11883
rect 947 11861 959 11883
rect 1015 11861 1031 11883
rect 1083 11861 1103 11883
rect 1151 11861 1175 11883
rect 811 11849 845 11861
rect 879 11849 913 11861
rect 947 11849 981 11861
rect 1015 11849 1049 11861
rect 1083 11849 1117 11861
rect 1151 11849 1185 11861
rect 1219 11849 1226 11883
rect 226 11821 1226 11849
rect 226 11812 236 11821
rect 270 11812 309 11821
rect 343 11812 382 11821
rect 416 11812 455 11821
rect 489 11812 527 11821
rect 561 11812 599 11821
rect 633 11812 671 11821
rect 705 11812 743 11821
rect 226 11778 233 11812
rect 270 11787 301 11812
rect 343 11787 369 11812
rect 416 11787 437 11812
rect 489 11787 505 11812
rect 561 11787 573 11812
rect 633 11787 641 11812
rect 705 11787 709 11812
rect 267 11778 301 11787
rect 335 11778 369 11787
rect 403 11778 437 11787
rect 471 11778 505 11787
rect 539 11778 573 11787
rect 607 11778 641 11787
rect 675 11778 709 11787
rect 777 11812 815 11821
rect 849 11812 887 11821
rect 921 11812 959 11821
rect 993 11812 1031 11821
rect 1065 11812 1103 11821
rect 1137 11812 1175 11821
rect 1209 11812 1226 11821
rect 743 11778 777 11787
rect 811 11787 815 11812
rect 879 11787 887 11812
rect 947 11787 959 11812
rect 1015 11787 1031 11812
rect 1083 11787 1103 11812
rect 1151 11787 1175 11812
rect 811 11778 845 11787
rect 879 11778 913 11787
rect 947 11778 981 11787
rect 1015 11778 1049 11787
rect 1083 11778 1117 11787
rect 1151 11778 1185 11787
rect 1219 11778 1226 11812
rect 226 11747 1226 11778
rect 226 11741 236 11747
rect 270 11741 309 11747
rect 343 11741 382 11747
rect 416 11741 455 11747
rect 489 11741 527 11747
rect 561 11741 599 11747
rect 633 11741 671 11747
rect 705 11741 743 11747
rect 226 11707 233 11741
rect 270 11713 301 11741
rect 343 11713 369 11741
rect 416 11713 437 11741
rect 489 11713 505 11741
rect 561 11713 573 11741
rect 633 11713 641 11741
rect 705 11713 709 11741
rect 267 11707 301 11713
rect 335 11707 369 11713
rect 403 11707 437 11713
rect 471 11707 505 11713
rect 539 11707 573 11713
rect 607 11707 641 11713
rect 675 11707 709 11713
rect 777 11741 815 11747
rect 849 11741 887 11747
rect 921 11741 959 11747
rect 993 11741 1031 11747
rect 1065 11741 1103 11747
rect 1137 11741 1175 11747
rect 1209 11741 1226 11747
rect 743 11707 777 11713
rect 811 11713 815 11741
rect 879 11713 887 11741
rect 947 11713 959 11741
rect 1015 11713 1031 11741
rect 1083 11713 1103 11741
rect 1151 11713 1175 11741
rect 811 11707 845 11713
rect 879 11707 913 11713
rect 947 11707 981 11713
rect 1015 11707 1049 11713
rect 1083 11707 1117 11713
rect 1151 11707 1185 11713
rect 1219 11707 1226 11741
rect 226 11673 1226 11707
rect 226 11670 236 11673
rect 270 11670 309 11673
rect 343 11670 382 11673
rect 416 11670 455 11673
rect 489 11670 527 11673
rect 561 11670 599 11673
rect 633 11670 671 11673
rect 705 11670 743 11673
rect 226 11636 233 11670
rect 270 11639 301 11670
rect 343 11639 369 11670
rect 416 11639 437 11670
rect 489 11639 505 11670
rect 561 11639 573 11670
rect 633 11639 641 11670
rect 705 11639 709 11670
rect 267 11636 301 11639
rect 335 11636 369 11639
rect 403 11636 437 11639
rect 471 11636 505 11639
rect 539 11636 573 11639
rect 607 11636 641 11639
rect 675 11636 709 11639
rect 777 11670 815 11673
rect 849 11670 887 11673
rect 921 11670 959 11673
rect 993 11670 1031 11673
rect 1065 11670 1103 11673
rect 1137 11670 1175 11673
rect 1209 11670 1226 11673
rect 743 11636 777 11639
rect 811 11639 815 11670
rect 879 11639 887 11670
rect 947 11639 959 11670
rect 1015 11639 1031 11670
rect 1083 11639 1103 11670
rect 1151 11639 1175 11670
rect 811 11636 845 11639
rect 879 11636 913 11639
rect 947 11636 981 11639
rect 1015 11636 1049 11639
rect 1083 11636 1117 11639
rect 1151 11636 1185 11639
rect 1219 11636 1226 11670
rect 226 11599 1226 11636
rect 6819 11694 6859 11728
rect 6893 11694 6932 11728
rect 6966 11694 7005 11728
rect 7039 11694 7078 11728
rect 7112 11694 7151 11728
rect 7185 11694 7224 11728
rect 7258 11694 7297 11728
rect 7331 11694 7370 11728
rect 7404 11694 7443 11728
rect 7477 11694 7516 11728
rect 7550 11694 7589 11728
rect 7623 11694 7662 11728
rect 6785 11656 7696 11694
rect 6819 11622 6859 11656
rect 6893 11622 6932 11656
rect 6966 11622 7005 11656
rect 7039 11622 7078 11656
rect 7112 11622 7151 11656
rect 7185 11622 7224 11656
rect 7258 11622 7297 11656
rect 7331 11622 7370 11656
rect 7404 11622 7443 11656
rect 7477 11622 7516 11656
rect 7550 11622 7589 11656
rect 7623 11622 7662 11656
rect 226 11598 236 11599
rect 270 11598 309 11599
rect 343 11598 382 11599
rect 416 11598 455 11599
rect 489 11598 527 11599
rect 561 11598 599 11599
rect 633 11598 671 11599
rect 705 11598 743 11599
rect 226 11564 233 11598
rect 270 11565 301 11598
rect 343 11565 369 11598
rect 416 11565 437 11598
rect 489 11565 505 11598
rect 561 11565 573 11598
rect 633 11565 641 11598
rect 705 11565 709 11598
rect 267 11564 301 11565
rect 335 11564 369 11565
rect 403 11564 437 11565
rect 471 11564 505 11565
rect 539 11564 573 11565
rect 607 11564 641 11565
rect 675 11564 709 11565
rect 777 11598 815 11599
rect 849 11598 887 11599
rect 921 11598 959 11599
rect 993 11598 1031 11599
rect 1065 11598 1103 11599
rect 1137 11598 1175 11599
rect 1209 11598 1226 11599
rect 743 11564 777 11565
rect 811 11565 815 11598
rect 879 11565 887 11598
rect 947 11565 959 11598
rect 1015 11565 1031 11598
rect 1083 11565 1103 11598
rect 1151 11565 1175 11598
rect 811 11564 845 11565
rect 879 11564 913 11565
rect 947 11564 981 11565
rect 1015 11564 1049 11565
rect 1083 11564 1117 11565
rect 1151 11564 1185 11565
rect 1219 11564 1226 11598
rect 226 11526 1226 11564
rect 226 11492 233 11526
rect 267 11525 301 11526
rect 335 11525 369 11526
rect 403 11525 437 11526
rect 471 11525 505 11526
rect 539 11525 573 11526
rect 607 11525 641 11526
rect 675 11525 709 11526
rect 270 11492 301 11525
rect 343 11492 369 11525
rect 416 11492 437 11525
rect 489 11492 505 11525
rect 561 11492 573 11525
rect 633 11492 641 11525
rect 705 11492 709 11525
rect 743 11525 777 11526
rect 226 11491 236 11492
rect 270 11491 309 11492
rect 343 11491 382 11492
rect 416 11491 455 11492
rect 489 11491 527 11492
rect 561 11491 599 11492
rect 633 11491 671 11492
rect 705 11491 743 11492
rect 811 11525 845 11526
rect 879 11525 913 11526
rect 947 11525 981 11526
rect 1015 11525 1049 11526
rect 1083 11525 1117 11526
rect 1151 11525 1185 11526
rect 811 11492 815 11525
rect 879 11492 887 11525
rect 947 11492 959 11525
rect 1015 11492 1031 11525
rect 1083 11492 1103 11525
rect 1151 11492 1175 11525
rect 1219 11492 1226 11526
rect 777 11491 815 11492
rect 849 11491 887 11492
rect 921 11491 959 11492
rect 993 11491 1031 11492
rect 1065 11491 1103 11492
rect 1137 11491 1175 11492
rect 1209 11491 1226 11492
rect 226 11468 1226 11491
rect 6746 11618 16309 11622
rect 6746 11584 6770 11618
rect 6804 11584 6839 11618
rect 6873 11584 6908 11618
rect 6942 11584 6977 11618
rect 7011 11584 7046 11618
rect 7080 11584 7115 11618
rect 7149 11584 7184 11618
rect 7218 11584 7253 11618
rect 7287 11584 7322 11618
rect 7356 11584 7391 11618
rect 7425 11584 7460 11618
rect 7494 11584 7529 11618
rect 7563 11584 7598 11618
rect 7632 11584 7667 11618
rect 7701 11584 7736 11618
rect 7770 11584 7805 11618
rect 7839 11584 7874 11618
rect 7908 11584 7943 11618
rect 7977 11584 8012 11618
rect 8046 11584 8081 11618
rect 8115 11584 8150 11618
rect 8184 11584 8219 11618
rect 8253 11584 8288 11618
rect 8322 11584 8357 11618
rect 8391 11584 8426 11618
rect 8460 11584 8495 11618
rect 8529 11584 8564 11618
rect 8598 11584 8633 11618
rect 8667 11584 8702 11618
rect 8736 11584 8771 11618
rect 8805 11584 8840 11618
rect 8874 11584 8909 11618
rect 8943 11584 8978 11618
rect 9012 11584 9046 11618
rect 9080 11584 9114 11618
rect 9148 11584 9182 11618
rect 9216 11584 9250 11618
rect 9284 11584 9318 11618
rect 9352 11584 9386 11618
rect 9420 11584 9454 11618
rect 9488 11584 9522 11618
rect 9556 11584 9590 11618
rect 9624 11584 9658 11618
rect 9692 11584 9726 11618
rect 9760 11584 9794 11618
rect 9828 11584 9862 11618
rect 9896 11584 9930 11618
rect 9964 11584 9998 11618
rect 10032 11584 10066 11618
rect 10100 11584 10134 11618
rect 10168 11584 10202 11618
rect 10236 11584 10270 11618
rect 10304 11588 16309 11618
rect 16343 11588 16379 11622
rect 16413 11588 16449 11622
rect 16483 11588 16519 11622
rect 16553 11588 16589 11622
rect 16623 11588 16658 11622
rect 16692 11588 16727 11622
rect 16761 11588 16796 11622
rect 16830 11588 16865 11622
rect 16899 11588 16934 11622
rect 16968 11588 17003 11622
rect 17037 11588 17072 11622
rect 17106 11588 17141 11622
rect 17175 11588 17210 11622
rect 17244 11588 17279 11622
rect 17313 11588 17348 11622
rect 17382 11588 17417 11622
rect 17451 11617 17486 11622
rect 17479 11588 17486 11617
rect 17520 11617 17555 11622
rect 17589 11617 17624 11622
rect 17658 11617 17693 11622
rect 17520 11588 17525 11617
rect 17589 11588 17605 11617
rect 17658 11588 17684 11617
rect 17727 11588 17762 11622
rect 17796 11617 17831 11622
rect 17865 11617 17900 11622
rect 17934 11617 17969 11622
rect 18003 11617 18038 11622
rect 17797 11588 17831 11617
rect 17876 11588 17900 11617
rect 17955 11588 17969 11617
rect 18034 11588 18038 11617
rect 18072 11617 18107 11622
rect 18141 11617 18176 11622
rect 18072 11588 18079 11617
rect 18141 11588 18158 11617
rect 18210 11588 18245 11622
rect 18279 11588 18314 11622
rect 18348 11588 18383 11622
rect 18417 11588 18452 11622
rect 18486 11615 18521 11622
rect 18555 11615 18590 11622
rect 18486 11588 18500 11615
rect 18555 11588 18585 11615
rect 18624 11588 18659 11622
rect 18693 11615 18728 11622
rect 18762 11615 18797 11622
rect 18703 11588 18728 11615
rect 18787 11588 18797 11615
rect 18831 11615 18866 11622
rect 18900 11615 18935 11622
rect 18831 11588 18837 11615
rect 18900 11588 18921 11615
rect 18969 11588 19004 11622
rect 19038 11588 19073 11622
rect 19107 11588 19142 11622
rect 19176 11588 19211 11622
rect 19245 11588 19280 11622
rect 19314 11588 19349 11622
rect 19383 11588 19418 11622
rect 19452 11588 19487 11622
rect 19521 11588 19556 11622
rect 19590 11588 19625 11622
rect 19659 11621 19683 11622
rect 19773 11621 19797 11629
rect 19659 11595 19797 11621
rect 19831 11595 19866 11629
rect 19900 11595 19935 11629
rect 19969 11595 20004 11629
rect 20038 11595 20073 11629
rect 20107 11595 20142 11629
rect 20176 11595 20211 11629
rect 20245 11595 20280 11629
rect 20314 11595 20349 11629
rect 20383 11595 20418 11629
rect 20452 11595 20487 11629
rect 20521 11595 20556 11629
rect 20590 11595 20625 11629
rect 20659 11595 20694 11629
rect 20728 11595 20763 11629
rect 20797 11595 20832 11629
rect 20866 11595 20901 11629
rect 20935 11595 20970 11629
rect 21004 11595 21039 11629
rect 21073 11595 21108 11629
rect 21142 11595 21177 11629
rect 21211 11595 21246 11629
rect 21280 11595 21315 11629
rect 21349 11595 21384 11629
rect 21418 11595 21453 11629
rect 21487 11595 21522 11629
rect 21556 11595 21591 11629
rect 21625 11595 21660 11629
rect 21694 11595 21729 11629
rect 21763 11595 21798 11629
rect 21832 11595 21866 11629
rect 21900 11595 21934 11629
rect 21968 11595 22002 11629
rect 22036 11595 22070 11629
rect 22104 11595 22138 11629
rect 22172 11595 22206 11629
rect 22240 11595 22274 11629
rect 22308 11595 22342 11629
rect 22376 11595 22410 11629
rect 22444 11595 22478 11629
rect 22512 11595 22546 11629
rect 22580 11595 22614 11629
rect 22648 11595 22682 11629
rect 22716 11595 22750 11629
rect 22784 11595 22818 11629
rect 22852 11595 22886 11629
rect 22920 11595 22954 11629
rect 22988 11595 23022 11629
rect 23056 11595 23090 11629
rect 23124 11595 23158 11629
rect 23192 11595 23226 11629
rect 23260 11595 23294 11629
rect 23328 11595 23362 11629
rect 23396 11595 23430 11629
rect 23464 11595 23498 11629
rect 23532 11595 23566 11629
rect 23600 11595 23634 11629
rect 23668 11595 23702 11629
rect 23736 11595 23770 11629
rect 23804 11595 23838 11629
rect 23872 11595 23906 11629
rect 23940 11595 23974 11629
rect 24008 11595 24042 11629
rect 24076 11595 24110 11629
rect 24144 11595 24178 11629
rect 24212 11595 24246 11629
rect 24280 11595 24314 11629
rect 24348 11595 24382 11629
rect 24416 11595 24450 11629
rect 24484 11595 24518 11629
rect 24552 11595 24586 11629
rect 24620 11595 24654 11629
rect 24688 11595 24722 11629
rect 24756 11595 24790 11629
rect 24824 11595 24858 11629
rect 24892 11595 24926 11629
rect 24960 11595 24994 11629
rect 25028 11595 25062 11629
rect 25096 11595 25130 11629
rect 25164 11595 25198 11629
rect 25232 11595 25266 11629
rect 25300 11595 25334 11629
rect 25368 11595 25402 11629
rect 25436 11595 25470 11629
rect 25504 11595 25528 11629
rect 19659 11588 20283 11595
rect 10304 11584 17445 11588
rect 6746 11583 17445 11584
rect 17479 11583 17525 11588
rect 17559 11583 17605 11588
rect 17639 11583 17684 11588
rect 17718 11583 17763 11588
rect 17797 11583 17842 11588
rect 17876 11583 17921 11588
rect 17955 11583 18000 11588
rect 18034 11583 18079 11588
rect 18113 11583 18158 11588
rect 18192 11583 18500 11588
rect 6746 11581 18500 11583
rect 18534 11581 18585 11588
rect 18619 11581 18669 11588
rect 18703 11581 18753 11588
rect 18787 11581 18837 11588
rect 18871 11581 18921 11588
rect 18955 11581 25528 11588
rect 6746 11579 25528 11581
rect 6746 11546 6779 11579
rect 6813 11546 6867 11579
rect 6901 11546 6955 11579
rect 6989 11546 7043 11579
rect 7077 11546 7131 11579
rect 7165 11577 25528 11579
rect 7165 11546 7577 11577
rect 7611 11546 7651 11577
rect 7685 11546 7725 11577
rect 7759 11546 7799 11577
rect 7833 11546 7873 11577
rect 7907 11546 7947 11577
rect 7981 11546 8021 11577
rect 8055 11546 8095 11577
rect 8129 11546 8169 11577
rect 8203 11546 8243 11577
rect 8277 11546 8317 11577
rect 8351 11546 8391 11577
rect 6746 11512 6770 11546
rect 6813 11545 6839 11546
rect 6901 11545 6908 11546
rect 6804 11512 6839 11545
rect 6873 11512 6908 11545
rect 6942 11545 6955 11546
rect 7011 11545 7043 11546
rect 6942 11512 6977 11545
rect 7011 11512 7046 11545
rect 7080 11512 7115 11546
rect 7165 11545 7184 11546
rect 7149 11512 7184 11545
rect 7218 11512 7253 11546
rect 7287 11512 7322 11546
rect 7356 11512 7391 11546
rect 7425 11512 7460 11546
rect 7494 11512 7529 11546
rect 7563 11543 7577 11546
rect 7632 11543 7651 11546
rect 7701 11543 7725 11546
rect 7770 11543 7799 11546
rect 7839 11543 7873 11546
rect 7563 11512 7598 11543
rect 7632 11512 7667 11543
rect 7701 11512 7736 11543
rect 7770 11512 7805 11543
rect 7839 11512 7874 11543
rect 7908 11512 7943 11546
rect 7981 11543 8012 11546
rect 8055 11543 8081 11546
rect 8129 11543 8150 11546
rect 8203 11543 8219 11546
rect 8277 11543 8288 11546
rect 8351 11543 8357 11546
rect 7977 11512 8012 11543
rect 8046 11512 8081 11543
rect 8115 11512 8150 11543
rect 8184 11512 8219 11543
rect 8253 11512 8288 11543
rect 8322 11512 8357 11543
rect 8425 11546 8465 11577
rect 8499 11546 8539 11577
rect 8573 11546 8613 11577
rect 8647 11546 8687 11577
rect 8721 11546 8761 11577
rect 8795 11546 8835 11577
rect 8869 11546 8909 11577
rect 8943 11546 8983 11577
rect 9017 11546 9058 11577
rect 9092 11546 9133 11577
rect 9167 11546 9208 11577
rect 9242 11546 9283 11577
rect 9317 11546 9358 11577
rect 9392 11546 9433 11577
rect 9467 11546 9508 11577
rect 9542 11546 10404 11577
rect 8425 11543 8426 11546
rect 8391 11512 8426 11543
rect 8460 11543 8465 11546
rect 8529 11543 8539 11546
rect 8598 11543 8613 11546
rect 8667 11543 8687 11546
rect 8736 11543 8761 11546
rect 8805 11543 8835 11546
rect 8460 11512 8495 11543
rect 8529 11512 8564 11543
rect 8598 11512 8633 11543
rect 8667 11512 8702 11543
rect 8736 11512 8771 11543
rect 8805 11512 8840 11543
rect 8874 11512 8909 11546
rect 8943 11512 8978 11546
rect 9017 11543 9046 11546
rect 9092 11543 9114 11546
rect 9167 11543 9182 11546
rect 9242 11543 9250 11546
rect 9317 11543 9318 11546
rect 9012 11512 9046 11543
rect 9080 11512 9114 11543
rect 9148 11512 9182 11543
rect 9216 11512 9250 11543
rect 9284 11512 9318 11543
rect 9352 11543 9358 11546
rect 9420 11543 9433 11546
rect 9488 11543 9508 11546
rect 9352 11512 9386 11543
rect 9420 11512 9454 11543
rect 9488 11512 9522 11543
rect 9556 11512 9590 11546
rect 9624 11512 9658 11546
rect 9692 11512 9726 11546
rect 9760 11512 9794 11546
rect 9828 11512 9862 11546
rect 9896 11512 9930 11546
rect 9964 11512 9998 11546
rect 10032 11512 10066 11546
rect 10100 11512 10134 11546
rect 10168 11512 10202 11546
rect 10236 11512 10270 11546
rect 10304 11543 10404 11546
rect 10438 11543 10473 11577
rect 10507 11543 10542 11577
rect 10576 11543 10611 11577
rect 10645 11543 10680 11577
rect 10714 11543 10749 11577
rect 10783 11543 10818 11577
rect 10852 11543 10887 11577
rect 10921 11543 10956 11577
rect 10990 11543 11025 11577
rect 11059 11543 11094 11577
rect 11128 11543 11163 11577
rect 11197 11543 11232 11577
rect 11266 11543 11301 11577
rect 11335 11543 11370 11577
rect 11404 11543 11439 11577
rect 11473 11543 11508 11577
rect 11542 11543 11577 11577
rect 11611 11543 11646 11577
rect 11680 11543 11715 11577
rect 11749 11543 11784 11577
rect 11818 11543 11853 11577
rect 11887 11543 11922 11577
rect 11956 11543 11991 11577
rect 12025 11543 12060 11577
rect 12094 11543 12129 11577
rect 12163 11543 12198 11577
rect 12232 11543 12267 11577
rect 12301 11543 12336 11577
rect 12370 11543 12405 11577
rect 12439 11543 12474 11577
rect 12508 11543 12543 11577
rect 12577 11543 12612 11577
rect 12646 11543 12681 11577
rect 12715 11543 12750 11577
rect 12784 11543 12819 11577
rect 12853 11543 12888 11577
rect 12922 11543 12957 11577
rect 12991 11543 13026 11577
rect 13060 11543 13095 11577
rect 13129 11543 13164 11577
rect 13198 11543 13233 11577
rect 13267 11543 13302 11577
rect 13336 11543 13371 11577
rect 10304 11512 13371 11543
rect 6746 11509 13371 11512
rect 6746 11507 10404 11509
rect 6746 11474 6779 11507
rect 6813 11474 6867 11507
rect 6901 11474 6955 11507
rect 6989 11474 7043 11507
rect 7077 11474 7131 11507
rect 7165 11489 10404 11507
rect 7165 11474 7577 11489
rect 7611 11474 7651 11489
rect 7685 11474 7725 11489
rect 7759 11474 7799 11489
rect 7833 11474 7873 11489
rect 7907 11474 7947 11489
rect 7981 11474 8021 11489
rect 8055 11474 8095 11489
rect 8129 11474 8169 11489
rect 8203 11474 8243 11489
rect 8277 11474 8317 11489
rect 8351 11474 8391 11489
rect 6746 11440 6770 11474
rect 6813 11473 6839 11474
rect 6901 11473 6908 11474
rect 6804 11440 6839 11473
rect 6873 11440 6908 11473
rect 6942 11473 6955 11474
rect 7011 11473 7043 11474
rect 6942 11440 6977 11473
rect 7011 11440 7046 11473
rect 7080 11440 7115 11474
rect 7165 11473 7184 11474
rect 7149 11440 7184 11473
rect 7218 11440 7253 11474
rect 7287 11440 7322 11474
rect 7356 11440 7391 11474
rect 7425 11440 7460 11474
rect 7494 11440 7529 11474
rect 7563 11455 7577 11474
rect 7632 11455 7651 11474
rect 7701 11455 7725 11474
rect 7770 11455 7799 11474
rect 7839 11455 7873 11474
rect 7563 11440 7598 11455
rect 7632 11440 7667 11455
rect 7701 11440 7736 11455
rect 7770 11440 7805 11455
rect 7839 11440 7874 11455
rect 7908 11440 7943 11474
rect 7981 11455 8012 11474
rect 8055 11455 8081 11474
rect 8129 11455 8150 11474
rect 8203 11455 8219 11474
rect 8277 11455 8288 11474
rect 8351 11455 8357 11474
rect 7977 11440 8012 11455
rect 8046 11440 8081 11455
rect 8115 11440 8150 11455
rect 8184 11440 8219 11455
rect 8253 11440 8288 11455
rect 8322 11440 8357 11455
rect 8425 11474 8465 11489
rect 8499 11474 8539 11489
rect 8573 11474 8613 11489
rect 8647 11474 8687 11489
rect 8721 11474 8761 11489
rect 8795 11474 8835 11489
rect 8869 11474 8909 11489
rect 8943 11474 8983 11489
rect 9017 11474 9058 11489
rect 9092 11474 9133 11489
rect 9167 11474 9208 11489
rect 9242 11474 9283 11489
rect 9317 11474 9358 11489
rect 9392 11474 9433 11489
rect 9467 11474 9508 11489
rect 9542 11475 10404 11489
rect 10438 11475 10473 11509
rect 10507 11475 10542 11509
rect 10576 11475 10611 11509
rect 10645 11475 10680 11509
rect 10714 11475 10749 11509
rect 10783 11475 10818 11509
rect 10852 11475 10887 11509
rect 10921 11475 10956 11509
rect 10990 11475 11025 11509
rect 11059 11475 11094 11509
rect 11128 11475 11163 11509
rect 11197 11475 11232 11509
rect 11266 11475 11301 11509
rect 11335 11475 11370 11509
rect 11404 11475 11439 11509
rect 11473 11475 11508 11509
rect 11542 11475 11577 11509
rect 11611 11475 11646 11509
rect 11680 11475 11715 11509
rect 11749 11475 11784 11509
rect 11818 11475 11853 11509
rect 11887 11475 11922 11509
rect 11956 11475 11991 11509
rect 12025 11475 12060 11509
rect 12094 11475 12129 11509
rect 12163 11475 12198 11509
rect 12232 11475 12267 11509
rect 12301 11475 12336 11509
rect 12370 11475 12405 11509
rect 12439 11475 12474 11509
rect 12508 11475 12543 11509
rect 12577 11475 12612 11509
rect 12646 11475 12681 11509
rect 12715 11475 12750 11509
rect 12784 11475 12819 11509
rect 12853 11475 12888 11509
rect 12922 11475 12957 11509
rect 12991 11475 13026 11509
rect 13060 11475 13095 11509
rect 13129 11475 13164 11509
rect 13198 11475 13233 11509
rect 13267 11475 13302 11509
rect 13336 11475 13371 11509
rect 9542 11474 13371 11475
rect 8425 11455 8426 11474
rect 8391 11440 8426 11455
rect 8460 11455 8465 11474
rect 8529 11455 8539 11474
rect 8598 11455 8613 11474
rect 8667 11455 8687 11474
rect 8736 11455 8761 11474
rect 8805 11455 8835 11474
rect 8460 11440 8495 11455
rect 8529 11440 8564 11455
rect 8598 11440 8633 11455
rect 8667 11440 8702 11455
rect 8736 11440 8771 11455
rect 8805 11440 8840 11455
rect 8874 11440 8909 11474
rect 8943 11440 8978 11474
rect 9017 11455 9046 11474
rect 9092 11455 9114 11474
rect 9167 11455 9182 11474
rect 9242 11455 9250 11474
rect 9317 11455 9318 11474
rect 9012 11440 9046 11455
rect 9080 11440 9114 11455
rect 9148 11440 9182 11455
rect 9216 11440 9250 11455
rect 9284 11440 9318 11455
rect 9352 11455 9358 11474
rect 9420 11455 9433 11474
rect 9488 11455 9508 11474
rect 9352 11440 9386 11455
rect 9420 11440 9454 11455
rect 9488 11440 9522 11455
rect 9556 11440 9590 11474
rect 9624 11440 9658 11474
rect 9692 11440 9726 11474
rect 9760 11440 9794 11474
rect 9828 11440 9862 11474
rect 9896 11440 9930 11474
rect 9964 11440 9998 11474
rect 10032 11440 10066 11474
rect 10100 11440 10134 11474
rect 10168 11440 10202 11474
rect 10236 11440 10270 11474
rect 10304 11452 13371 11474
rect 16261 11554 25528 11577
rect 16261 11520 16309 11554
rect 16343 11520 16379 11554
rect 16413 11520 16449 11554
rect 16483 11520 16519 11554
rect 16553 11520 16589 11554
rect 16623 11520 16658 11554
rect 16692 11520 16727 11554
rect 16761 11520 16796 11554
rect 16830 11520 16865 11554
rect 16899 11520 16934 11554
rect 16968 11520 17003 11554
rect 17037 11520 17072 11554
rect 17106 11520 17141 11554
rect 17175 11520 17210 11554
rect 17244 11520 17279 11554
rect 17313 11520 17348 11554
rect 17382 11520 17417 11554
rect 17451 11545 17486 11554
rect 17479 11520 17486 11545
rect 17520 11545 17555 11554
rect 17589 11545 17624 11554
rect 17658 11545 17693 11554
rect 17520 11520 17525 11545
rect 17589 11520 17605 11545
rect 17658 11520 17684 11545
rect 17727 11520 17762 11554
rect 17796 11545 17831 11554
rect 17865 11545 17900 11554
rect 17934 11545 17969 11554
rect 18003 11545 18038 11554
rect 17797 11520 17831 11545
rect 17876 11520 17900 11545
rect 17955 11520 17969 11545
rect 18034 11520 18038 11545
rect 18072 11545 18107 11554
rect 18141 11545 18176 11554
rect 18072 11520 18079 11545
rect 18141 11520 18158 11545
rect 18210 11520 18245 11554
rect 18279 11520 18314 11554
rect 18348 11520 18383 11554
rect 18417 11520 18452 11554
rect 18486 11543 18521 11554
rect 18555 11543 18590 11554
rect 18486 11520 18500 11543
rect 18555 11520 18585 11543
rect 18624 11520 18659 11554
rect 18693 11543 18728 11554
rect 18762 11543 18797 11554
rect 18703 11520 18728 11543
rect 18787 11520 18797 11543
rect 18831 11543 18866 11554
rect 18900 11543 18935 11554
rect 18831 11520 18837 11543
rect 18900 11520 18921 11543
rect 18969 11520 19004 11554
rect 19038 11520 19073 11554
rect 19107 11520 19142 11554
rect 19176 11520 19211 11554
rect 19245 11520 19280 11554
rect 19314 11520 19349 11554
rect 19383 11520 19418 11554
rect 19452 11520 19487 11554
rect 19521 11520 19556 11554
rect 19590 11520 19625 11554
rect 19659 11536 25528 11554
rect 19659 11527 20283 11536
rect 19659 11520 19683 11527
rect 16261 11511 17445 11520
rect 17479 11511 17525 11520
rect 17559 11511 17605 11520
rect 17639 11511 17684 11520
rect 17718 11511 17763 11520
rect 17797 11511 17842 11520
rect 17876 11511 17921 11520
rect 17955 11511 18000 11520
rect 18034 11511 18079 11520
rect 18113 11511 18158 11520
rect 18192 11511 18500 11520
rect 16261 11509 18500 11511
rect 18534 11509 18585 11520
rect 18619 11509 18669 11520
rect 18703 11509 18753 11520
rect 18787 11509 18837 11520
rect 18871 11509 18921 11520
rect 18955 11509 19683 11520
rect 16261 11486 19683 11509
rect 16261 11452 16309 11486
rect 16343 11452 16379 11486
rect 16413 11452 16449 11486
rect 16483 11452 16519 11486
rect 16553 11452 16589 11486
rect 16623 11452 16658 11486
rect 16692 11452 16727 11486
rect 16761 11452 16796 11486
rect 16830 11452 16865 11486
rect 16899 11452 16934 11486
rect 16968 11452 17003 11486
rect 17037 11452 17072 11486
rect 17106 11452 17141 11486
rect 17175 11452 17210 11486
rect 17244 11452 17279 11486
rect 17313 11452 17348 11486
rect 17382 11452 17417 11486
rect 17451 11473 17486 11486
rect 17479 11452 17486 11473
rect 17520 11473 17555 11486
rect 17589 11473 17624 11486
rect 17658 11473 17693 11486
rect 17520 11452 17525 11473
rect 17589 11452 17605 11473
rect 17658 11452 17684 11473
rect 17727 11452 17762 11486
rect 17796 11473 17831 11486
rect 17865 11473 17900 11486
rect 17934 11473 17969 11486
rect 18003 11473 18038 11486
rect 17797 11452 17831 11473
rect 17876 11452 17900 11473
rect 17955 11452 17969 11473
rect 18034 11452 18038 11473
rect 18072 11473 18107 11486
rect 18141 11473 18176 11486
rect 18072 11452 18079 11473
rect 18141 11452 18158 11473
rect 18210 11452 18245 11486
rect 18279 11452 18314 11486
rect 18348 11452 18383 11486
rect 18417 11452 18452 11486
rect 18486 11471 18521 11486
rect 18555 11471 18590 11486
rect 18486 11452 18500 11471
rect 18555 11452 18585 11471
rect 18624 11452 18659 11486
rect 18693 11471 18728 11486
rect 18762 11471 18797 11486
rect 18703 11452 18728 11471
rect 18787 11452 18797 11471
rect 18831 11471 18866 11486
rect 18900 11471 18935 11486
rect 18831 11452 18837 11471
rect 18900 11452 18921 11471
rect 18969 11452 19004 11486
rect 19038 11452 19073 11486
rect 19107 11452 19142 11486
rect 19176 11452 19211 11486
rect 19245 11452 19280 11486
rect 19314 11452 19349 11486
rect 19383 11452 19418 11486
rect 19452 11452 19487 11486
rect 19521 11452 19556 11486
rect 19590 11452 19625 11486
rect 19659 11452 19683 11486
rect 10304 11441 10456 11452
rect 10490 11441 10529 11452
rect 10563 11441 10602 11452
rect 10636 11441 10675 11452
rect 10709 11441 10748 11452
rect 10782 11441 10821 11452
rect 10855 11441 10893 11452
rect 10927 11441 10965 11452
rect 10999 11441 11037 11452
rect 11071 11441 11109 11452
rect 11143 11441 11181 11452
rect 11215 11441 11253 11452
rect 11287 11441 11325 11452
rect 11359 11441 11397 11452
rect 11431 11441 11469 11452
rect 11503 11441 11541 11452
rect 11575 11441 11613 11452
rect 11647 11441 11685 11452
rect 11719 11441 11757 11452
rect 11791 11441 11829 11452
rect 11863 11441 11901 11452
rect 11935 11441 11973 11452
rect 12007 11441 12045 11452
rect 12079 11441 12117 11452
rect 12151 11441 12189 11452
rect 12223 11441 12261 11452
rect 12295 11441 12333 11452
rect 12367 11441 13371 11452
rect 10304 11440 10404 11441
rect 6746 11435 10404 11440
rect 6746 11402 6779 11435
rect 6813 11402 6867 11435
rect 6901 11402 6955 11435
rect 6989 11402 7043 11435
rect 7077 11402 7131 11435
rect 7165 11407 10404 11435
rect 10438 11418 10456 11441
rect 10507 11418 10529 11441
rect 10576 11418 10602 11441
rect 10645 11418 10675 11441
rect 10714 11418 10748 11441
rect 10438 11407 10473 11418
rect 10507 11407 10542 11418
rect 10576 11407 10611 11418
rect 10645 11407 10680 11418
rect 10714 11407 10749 11418
rect 10783 11407 10818 11441
rect 10855 11418 10887 11441
rect 10927 11418 10956 11441
rect 10999 11418 11025 11441
rect 11071 11418 11094 11441
rect 11143 11418 11163 11441
rect 11215 11418 11232 11441
rect 11287 11418 11301 11441
rect 11359 11418 11370 11441
rect 11431 11418 11439 11441
rect 11503 11418 11508 11441
rect 11575 11418 11577 11441
rect 10852 11407 10887 11418
rect 10921 11407 10956 11418
rect 10990 11407 11025 11418
rect 11059 11407 11094 11418
rect 11128 11407 11163 11418
rect 11197 11407 11232 11418
rect 11266 11407 11301 11418
rect 11335 11407 11370 11418
rect 11404 11407 11439 11418
rect 11473 11407 11508 11418
rect 11542 11407 11577 11418
rect 11611 11418 11613 11441
rect 11680 11418 11685 11441
rect 11749 11418 11757 11441
rect 11818 11418 11829 11441
rect 11887 11418 11901 11441
rect 11956 11418 11973 11441
rect 12025 11418 12045 11441
rect 12094 11418 12117 11441
rect 12163 11418 12189 11441
rect 12232 11418 12261 11441
rect 12301 11418 12333 11441
rect 11611 11407 11646 11418
rect 11680 11407 11715 11418
rect 11749 11407 11784 11418
rect 11818 11407 11853 11418
rect 11887 11407 11922 11418
rect 11956 11407 11991 11418
rect 12025 11407 12060 11418
rect 12094 11407 12129 11418
rect 12163 11407 12198 11418
rect 12232 11407 12267 11418
rect 12301 11407 12336 11418
rect 12370 11407 12405 11441
rect 12439 11407 12474 11441
rect 12508 11407 12543 11441
rect 12577 11407 12612 11441
rect 12646 11407 12681 11441
rect 12715 11407 12750 11441
rect 12784 11407 12819 11441
rect 12853 11407 12888 11441
rect 12922 11407 12957 11441
rect 12991 11407 13026 11441
rect 13060 11407 13095 11441
rect 13129 11407 13164 11441
rect 13198 11407 13233 11441
rect 13267 11407 13302 11441
rect 13336 11407 13371 11441
rect 16261 11439 17445 11452
rect 17479 11439 17525 11452
rect 17559 11439 17605 11452
rect 17639 11439 17684 11452
rect 17718 11439 17763 11452
rect 17797 11439 17842 11452
rect 17876 11439 17921 11452
rect 17955 11439 18000 11452
rect 18034 11439 18079 11452
rect 18113 11439 18158 11452
rect 18192 11439 18500 11452
rect 16261 11437 18500 11439
rect 18534 11437 18585 11452
rect 18619 11437 18669 11452
rect 18703 11437 18753 11452
rect 18787 11437 18837 11452
rect 18871 11437 18921 11452
rect 18955 11437 19683 11452
rect 16261 11418 19683 11437
rect 16261 11407 16309 11418
rect 7165 11402 16309 11407
rect 6746 11368 6770 11402
rect 6813 11401 6839 11402
rect 6901 11401 6908 11402
rect 6804 11368 6839 11401
rect 6873 11368 6908 11401
rect 6942 11401 6955 11402
rect 7011 11401 7043 11402
rect 6942 11368 6977 11401
rect 7011 11368 7046 11401
rect 7080 11368 7115 11402
rect 7165 11401 7184 11402
rect 7149 11368 7184 11401
rect 7218 11368 7253 11402
rect 7287 11368 7322 11402
rect 7356 11368 7391 11402
rect 7425 11368 7460 11402
rect 7494 11368 7529 11402
rect 7563 11401 7598 11402
rect 7632 11401 7667 11402
rect 7701 11401 7736 11402
rect 7770 11401 7805 11402
rect 7839 11401 7874 11402
rect 7563 11368 7577 11401
rect 7632 11368 7651 11401
rect 7701 11368 7725 11401
rect 7770 11368 7799 11401
rect 7839 11368 7873 11401
rect 7908 11368 7943 11402
rect 7977 11401 8012 11402
rect 8046 11401 8081 11402
rect 8115 11401 8150 11402
rect 8184 11401 8219 11402
rect 8253 11401 8288 11402
rect 8322 11401 8357 11402
rect 7981 11368 8012 11401
rect 8055 11368 8081 11401
rect 8129 11368 8150 11401
rect 8203 11368 8219 11401
rect 8277 11368 8288 11401
rect 8351 11368 8357 11401
rect 8391 11401 8426 11402
rect 6746 11367 7577 11368
rect 7611 11367 7651 11368
rect 7685 11367 7725 11368
rect 7759 11367 7799 11368
rect 7833 11367 7873 11368
rect 7907 11367 7947 11368
rect 7981 11367 8021 11368
rect 8055 11367 8095 11368
rect 8129 11367 8169 11368
rect 8203 11367 8243 11368
rect 8277 11367 8317 11368
rect 8351 11367 8391 11368
rect 8425 11368 8426 11401
rect 8460 11401 8495 11402
rect 8529 11401 8564 11402
rect 8598 11401 8633 11402
rect 8667 11401 8702 11402
rect 8736 11401 8771 11402
rect 8805 11401 8840 11402
rect 8460 11368 8465 11401
rect 8529 11368 8539 11401
rect 8598 11368 8613 11401
rect 8667 11368 8687 11401
rect 8736 11368 8761 11401
rect 8805 11368 8835 11401
rect 8874 11368 8909 11402
rect 8943 11368 8978 11402
rect 9012 11401 9046 11402
rect 9080 11401 9114 11402
rect 9148 11401 9182 11402
rect 9216 11401 9250 11402
rect 9284 11401 9318 11402
rect 9017 11368 9046 11401
rect 9092 11368 9114 11401
rect 9167 11368 9182 11401
rect 9242 11368 9250 11401
rect 9317 11368 9318 11401
rect 9352 11401 9386 11402
rect 9420 11401 9454 11402
rect 9488 11401 9522 11402
rect 9352 11368 9358 11401
rect 9420 11368 9433 11401
rect 9488 11368 9508 11401
rect 9556 11368 9590 11402
rect 9624 11368 9658 11402
rect 9692 11368 9726 11402
rect 9760 11368 9794 11402
rect 9828 11368 9862 11402
rect 9896 11368 9930 11402
rect 9964 11368 9998 11402
rect 10032 11368 10066 11402
rect 10100 11368 10134 11402
rect 10168 11368 10202 11402
rect 10236 11368 10270 11402
rect 10304 11384 16309 11402
rect 16343 11384 16379 11418
rect 16413 11384 16449 11418
rect 16483 11384 16519 11418
rect 16553 11384 16589 11418
rect 16623 11384 16658 11418
rect 16692 11384 16727 11418
rect 16761 11384 16796 11418
rect 16830 11384 16865 11418
rect 16899 11384 16934 11418
rect 16968 11384 17003 11418
rect 17037 11384 17072 11418
rect 17106 11384 17141 11418
rect 17175 11384 17210 11418
rect 17244 11384 17279 11418
rect 17313 11384 17348 11418
rect 17382 11384 17417 11418
rect 17451 11401 17486 11418
rect 17479 11384 17486 11401
rect 17520 11401 17555 11418
rect 17589 11401 17624 11418
rect 17658 11401 17693 11418
rect 17520 11384 17525 11401
rect 17589 11384 17605 11401
rect 17658 11384 17684 11401
rect 17727 11384 17762 11418
rect 17796 11401 17831 11418
rect 17865 11401 17900 11418
rect 17934 11401 17969 11418
rect 18003 11401 18038 11418
rect 17797 11384 17831 11401
rect 17876 11384 17900 11401
rect 17955 11384 17969 11401
rect 18034 11384 18038 11401
rect 18072 11401 18107 11418
rect 18141 11401 18176 11418
rect 18072 11384 18079 11401
rect 18141 11384 18158 11401
rect 18210 11384 18245 11418
rect 18279 11384 18314 11418
rect 18348 11384 18383 11418
rect 18417 11384 18452 11418
rect 18486 11399 18521 11418
rect 18555 11399 18590 11418
rect 18486 11384 18500 11399
rect 18555 11384 18585 11399
rect 18624 11384 18659 11418
rect 18693 11399 18728 11418
rect 18762 11399 18797 11418
rect 18703 11384 18728 11399
rect 18787 11384 18797 11399
rect 18831 11399 18866 11418
rect 18900 11399 18935 11418
rect 18831 11384 18837 11399
rect 18900 11384 18921 11399
rect 18969 11384 19004 11418
rect 19038 11384 19073 11418
rect 19107 11384 19142 11418
rect 19176 11384 19211 11418
rect 19245 11384 19280 11418
rect 19314 11384 19349 11418
rect 19383 11384 19418 11418
rect 19452 11384 19487 11418
rect 19521 11384 19556 11418
rect 19590 11384 19625 11418
rect 19659 11384 19683 11418
rect 10304 11368 17445 11384
rect 8425 11367 8465 11368
rect 8499 11367 8539 11368
rect 8573 11367 8613 11368
rect 8647 11367 8687 11368
rect 8721 11367 8761 11368
rect 8795 11367 8835 11368
rect 8869 11367 8909 11368
rect 8943 11367 8983 11368
rect 9017 11367 9058 11368
rect 9092 11367 9133 11368
rect 9167 11367 9208 11368
rect 9242 11367 9283 11368
rect 9317 11367 9358 11368
rect 9392 11367 9433 11368
rect 9467 11367 9508 11368
rect 9542 11367 17445 11368
rect 17479 11367 17525 11384
rect 17559 11367 17605 11384
rect 17639 11367 17684 11384
rect 17718 11367 17763 11384
rect 17797 11367 17842 11384
rect 17876 11367 17921 11384
rect 17955 11367 18000 11384
rect 18034 11367 18079 11384
rect 18113 11367 18158 11384
rect 18192 11367 18500 11384
rect 6746 11365 18500 11367
rect 18534 11365 18585 11384
rect 18619 11365 18669 11384
rect 18703 11365 18753 11384
rect 18787 11365 18837 11384
rect 18871 11365 18921 11384
rect 18955 11365 19382 11384
rect 6746 11363 19382 11365
rect 6746 11330 6779 11363
rect 6813 11330 6867 11363
rect 6901 11330 6955 11363
rect 6989 11330 7043 11363
rect 7077 11330 7131 11363
rect 7165 11350 19382 11363
rect 7165 11338 16319 11350
rect 7165 11330 10456 11338
rect 6746 11296 6770 11330
rect 6813 11329 6839 11330
rect 6901 11329 6908 11330
rect 6804 11296 6839 11329
rect 6873 11296 6908 11329
rect 6942 11329 6955 11330
rect 7011 11329 7043 11330
rect 6942 11296 6977 11329
rect 7011 11296 7046 11329
rect 7080 11296 7115 11330
rect 7165 11329 7184 11330
rect 7149 11296 7184 11329
rect 7218 11296 7253 11330
rect 7287 11296 7322 11330
rect 7356 11296 7391 11330
rect 7425 11296 7460 11330
rect 7494 11296 7529 11330
rect 7563 11313 7598 11330
rect 7632 11313 7667 11330
rect 7701 11313 7736 11330
rect 7770 11313 7805 11330
rect 7839 11313 7874 11330
rect 7563 11296 7577 11313
rect 7632 11296 7651 11313
rect 7701 11296 7725 11313
rect 7770 11296 7799 11313
rect 7839 11296 7873 11313
rect 7908 11296 7943 11330
rect 7977 11313 8012 11330
rect 8046 11313 8081 11330
rect 8115 11313 8150 11330
rect 8184 11313 8219 11330
rect 8253 11313 8288 11330
rect 8322 11313 8357 11330
rect 7981 11296 8012 11313
rect 8055 11296 8081 11313
rect 8129 11296 8150 11313
rect 8203 11296 8219 11313
rect 8277 11296 8288 11313
rect 8351 11296 8357 11313
rect 8391 11313 8426 11330
rect 6746 11291 7577 11296
rect 6746 11258 6779 11291
rect 6813 11258 6867 11291
rect 6901 11258 6955 11291
rect 6989 11258 7043 11291
rect 7077 11258 7131 11291
rect 7165 11279 7577 11291
rect 7611 11279 7651 11296
rect 7685 11279 7725 11296
rect 7759 11279 7799 11296
rect 7833 11279 7873 11296
rect 7907 11279 7947 11296
rect 7981 11279 8021 11296
rect 8055 11279 8095 11296
rect 8129 11279 8169 11296
rect 8203 11279 8243 11296
rect 8277 11279 8317 11296
rect 8351 11279 8391 11296
rect 8425 11296 8426 11313
rect 8460 11313 8495 11330
rect 8529 11313 8564 11330
rect 8598 11313 8633 11330
rect 8667 11313 8702 11330
rect 8736 11313 8771 11330
rect 8805 11313 8840 11330
rect 8460 11296 8465 11313
rect 8529 11296 8539 11313
rect 8598 11296 8613 11313
rect 8667 11296 8687 11313
rect 8736 11296 8761 11313
rect 8805 11296 8835 11313
rect 8874 11296 8909 11330
rect 8943 11296 8978 11330
rect 9012 11313 9046 11330
rect 9080 11313 9114 11330
rect 9148 11313 9182 11330
rect 9216 11313 9250 11330
rect 9284 11313 9318 11330
rect 9017 11296 9046 11313
rect 9092 11296 9114 11313
rect 9167 11296 9182 11313
rect 9242 11296 9250 11313
rect 9317 11296 9318 11313
rect 9352 11313 9386 11330
rect 9420 11313 9454 11330
rect 9488 11313 9522 11330
rect 9352 11296 9358 11313
rect 9420 11296 9433 11313
rect 9488 11296 9508 11313
rect 9556 11296 9590 11330
rect 9624 11296 9658 11330
rect 9692 11296 9726 11330
rect 9760 11296 9794 11330
rect 9828 11296 9862 11330
rect 9896 11296 9930 11330
rect 9964 11296 9998 11330
rect 10032 11296 10066 11330
rect 10100 11296 10134 11330
rect 10168 11296 10202 11330
rect 10236 11296 10270 11330
rect 10304 11304 10456 11330
rect 10490 11304 10529 11338
rect 10563 11304 10602 11338
rect 10636 11304 10675 11338
rect 10709 11304 10748 11338
rect 10782 11304 10821 11338
rect 10855 11304 10893 11338
rect 10927 11304 10965 11338
rect 10999 11304 11037 11338
rect 11071 11304 11109 11338
rect 11143 11304 11181 11338
rect 11215 11304 11253 11338
rect 11287 11304 11325 11338
rect 11359 11304 11397 11338
rect 11431 11304 11469 11338
rect 11503 11304 11541 11338
rect 11575 11304 11613 11338
rect 11647 11304 11685 11338
rect 11719 11304 11757 11338
rect 11791 11304 11829 11338
rect 11863 11304 11901 11338
rect 11935 11304 11973 11338
rect 12007 11304 12045 11338
rect 12079 11304 12117 11338
rect 12151 11304 12189 11338
rect 12223 11304 12261 11338
rect 12295 11304 12333 11338
rect 12367 11304 13411 11338
rect 13445 11304 13485 11338
rect 13519 11304 13559 11338
rect 13593 11304 13633 11338
rect 13667 11304 13707 11338
rect 13741 11304 13781 11338
rect 13815 11304 13855 11338
rect 13889 11304 13929 11338
rect 13963 11304 14003 11338
rect 14037 11304 14077 11338
rect 14111 11304 14151 11338
rect 14185 11304 14225 11338
rect 14259 11304 14299 11338
rect 14333 11304 14372 11338
rect 14406 11304 14445 11338
rect 14479 11304 14518 11338
rect 14552 11304 14591 11338
rect 14625 11304 14664 11338
rect 14698 11304 14737 11338
rect 14771 11304 14810 11338
rect 14844 11304 14883 11338
rect 14917 11304 14956 11338
rect 14990 11304 15029 11338
rect 15063 11304 15102 11338
rect 15136 11304 15175 11338
rect 15209 11304 15248 11338
rect 15282 11304 15321 11338
rect 15355 11304 15394 11338
rect 15428 11304 15467 11338
rect 15501 11304 15540 11338
rect 15574 11304 15613 11338
rect 15647 11316 16319 11338
rect 16353 11316 16388 11350
rect 16422 11316 16457 11350
rect 16491 11316 16526 11350
rect 16560 11316 16594 11350
rect 16628 11316 16662 11350
rect 16696 11316 16730 11350
rect 16764 11316 16798 11350
rect 16832 11316 16866 11350
rect 16900 11316 16934 11350
rect 16968 11316 17002 11350
rect 17036 11316 17070 11350
rect 17104 11316 17138 11350
rect 17172 11316 17206 11350
rect 17240 11316 17274 11350
rect 17308 11316 17342 11350
rect 17376 11316 17410 11350
rect 17444 11329 17478 11350
rect 17512 11329 17546 11350
rect 17580 11329 17614 11350
rect 17444 11316 17445 11329
rect 17512 11316 17525 11329
rect 17580 11316 17605 11329
rect 17648 11316 17682 11350
rect 17716 11329 17750 11350
rect 17784 11329 17818 11350
rect 17852 11329 17886 11350
rect 17718 11316 17750 11329
rect 17797 11316 17818 11329
rect 17876 11316 17886 11329
rect 17920 11329 17954 11350
rect 17988 11329 18022 11350
rect 18056 11329 18090 11350
rect 17920 11316 17921 11329
rect 17988 11316 18000 11329
rect 18056 11316 18079 11329
rect 18124 11316 18158 11350
rect 18192 11316 18226 11350
rect 18260 11316 18294 11350
rect 18328 11316 18362 11350
rect 18396 11316 18430 11350
rect 18464 11316 18498 11350
rect 18532 11327 18566 11350
rect 18600 11327 18634 11350
rect 18534 11316 18566 11327
rect 18619 11316 18634 11327
rect 18668 11327 18702 11350
rect 18736 11327 18770 11350
rect 18804 11327 18838 11350
rect 18668 11316 18669 11327
rect 18736 11316 18753 11327
rect 18804 11316 18837 11327
rect 18872 11316 18906 11350
rect 18940 11327 18974 11350
rect 18955 11316 18974 11327
rect 19008 11316 19042 11350
rect 19076 11316 19110 11350
rect 19144 11316 19178 11350
rect 19212 11316 19246 11350
rect 19280 11316 19314 11350
rect 19348 11316 19382 11350
rect 10304 11296 14092 11304
rect 8425 11279 8465 11296
rect 8499 11279 8539 11296
rect 8573 11279 8613 11296
rect 8647 11279 8687 11296
rect 8721 11279 8761 11296
rect 8795 11279 8835 11296
rect 8869 11279 8909 11296
rect 8943 11279 8983 11296
rect 9017 11279 9058 11296
rect 9092 11279 9133 11296
rect 9167 11279 9208 11296
rect 9242 11279 9283 11296
rect 9317 11279 9358 11296
rect 9392 11279 9433 11296
rect 9467 11279 9508 11296
rect 9542 11279 14092 11296
rect 7165 11258 14092 11279
rect 6746 11224 6770 11258
rect 6813 11257 6839 11258
rect 6901 11257 6908 11258
rect 6804 11224 6839 11257
rect 6873 11224 6908 11257
rect 6942 11257 6955 11258
rect 7011 11257 7043 11258
rect 6942 11224 6977 11257
rect 7011 11224 7046 11257
rect 7080 11224 7115 11258
rect 7165 11257 7184 11258
rect 7149 11224 7184 11257
rect 7218 11224 7253 11258
rect 7287 11224 7322 11258
rect 7356 11224 7391 11258
rect 7425 11224 7460 11258
rect 7494 11224 7529 11258
rect 7563 11225 7598 11258
rect 7632 11225 7667 11258
rect 7701 11225 7736 11258
rect 7770 11225 7805 11258
rect 7839 11225 7874 11258
rect 7563 11224 7577 11225
rect 7632 11224 7651 11225
rect 7701 11224 7725 11225
rect 7770 11224 7799 11225
rect 7839 11224 7873 11225
rect 7908 11224 7943 11258
rect 7977 11225 8012 11258
rect 8046 11225 8081 11258
rect 8115 11225 8150 11258
rect 8184 11225 8219 11258
rect 8253 11225 8288 11258
rect 8322 11225 8357 11258
rect 7981 11224 8012 11225
rect 8055 11224 8081 11225
rect 8129 11224 8150 11225
rect 8203 11224 8219 11225
rect 8277 11224 8288 11225
rect 8351 11224 8357 11225
rect 8391 11225 8426 11258
rect 6746 11219 7577 11224
rect 6746 11186 6779 11219
rect 6813 11186 6867 11219
rect 6901 11186 6955 11219
rect 6989 11186 7043 11219
rect 7077 11186 7131 11219
rect 7165 11191 7577 11219
rect 7611 11191 7651 11224
rect 7685 11191 7725 11224
rect 7759 11191 7799 11224
rect 7833 11191 7873 11224
rect 7907 11191 7947 11224
rect 7981 11191 8021 11224
rect 8055 11191 8095 11224
rect 8129 11191 8169 11224
rect 8203 11191 8243 11224
rect 8277 11191 8317 11224
rect 8351 11191 8391 11224
rect 8425 11224 8426 11225
rect 8460 11225 8495 11258
rect 8529 11225 8564 11258
rect 8598 11225 8633 11258
rect 8667 11225 8702 11258
rect 8736 11225 8771 11258
rect 8805 11225 8840 11258
rect 8460 11224 8465 11225
rect 8529 11224 8539 11225
rect 8598 11224 8613 11225
rect 8667 11224 8687 11225
rect 8736 11224 8761 11225
rect 8805 11224 8835 11225
rect 8874 11224 8909 11258
rect 8943 11224 8978 11258
rect 9012 11225 9046 11258
rect 9080 11225 9114 11258
rect 9148 11225 9182 11258
rect 9216 11225 9250 11258
rect 9284 11225 9318 11258
rect 9017 11224 9046 11225
rect 9092 11224 9114 11225
rect 9167 11224 9182 11225
rect 9242 11224 9250 11225
rect 9317 11224 9318 11225
rect 9352 11225 9386 11258
rect 9420 11225 9454 11258
rect 9488 11225 9522 11258
rect 9352 11224 9358 11225
rect 9420 11224 9433 11225
rect 9488 11224 9508 11225
rect 9556 11224 9590 11258
rect 9624 11224 9658 11258
rect 9692 11224 9726 11258
rect 9760 11224 9794 11258
rect 9828 11224 9862 11258
rect 9896 11224 9930 11258
rect 9964 11224 9998 11258
rect 10032 11224 10066 11258
rect 10100 11224 10134 11258
rect 10168 11224 10202 11258
rect 10236 11224 10270 11258
rect 10304 11231 14092 11258
rect 16285 11295 17445 11316
rect 17479 11295 17525 11316
rect 17559 11295 17605 11316
rect 17639 11295 17684 11316
rect 17718 11295 17763 11316
rect 17797 11295 17842 11316
rect 17876 11295 17921 11316
rect 17955 11295 18000 11316
rect 18034 11295 18079 11316
rect 18113 11295 18158 11316
rect 18192 11295 18500 11316
rect 16285 11293 18500 11295
rect 18534 11293 18585 11316
rect 18619 11293 18669 11316
rect 18703 11293 18753 11316
rect 18787 11293 18837 11316
rect 18871 11293 18921 11316
rect 18955 11293 19382 11316
rect 16285 11278 19382 11293
rect 16285 11244 16319 11278
rect 16353 11244 16388 11278
rect 16422 11244 16457 11278
rect 16491 11244 16526 11278
rect 16560 11244 16594 11278
rect 16628 11244 16662 11278
rect 16696 11244 16730 11278
rect 16764 11244 16798 11278
rect 16832 11244 16866 11278
rect 16900 11244 16934 11278
rect 16968 11244 17002 11278
rect 17036 11244 17070 11278
rect 17104 11244 17138 11278
rect 17172 11244 17206 11278
rect 17240 11244 17274 11278
rect 17308 11244 17342 11278
rect 17376 11244 17410 11278
rect 17444 11257 17478 11278
rect 17512 11257 17546 11278
rect 17580 11257 17614 11278
rect 17444 11244 17445 11257
rect 17512 11244 17525 11257
rect 17580 11244 17605 11257
rect 17648 11244 17682 11278
rect 17716 11257 17750 11278
rect 17784 11257 17818 11278
rect 17852 11257 17886 11278
rect 17718 11244 17750 11257
rect 17797 11244 17818 11257
rect 17876 11244 17886 11257
rect 17920 11257 17954 11278
rect 17988 11257 18022 11278
rect 18056 11257 18090 11278
rect 17920 11244 17921 11257
rect 17988 11244 18000 11257
rect 18056 11244 18079 11257
rect 18124 11244 18158 11278
rect 18192 11244 18226 11278
rect 18260 11244 18294 11278
rect 18328 11244 18362 11278
rect 18396 11244 18430 11278
rect 18464 11244 18498 11278
rect 18532 11255 18566 11278
rect 18600 11255 18634 11278
rect 18534 11244 18566 11255
rect 18619 11244 18634 11255
rect 18668 11255 18702 11278
rect 18736 11255 18770 11278
rect 18804 11255 18838 11278
rect 18668 11244 18669 11255
rect 18736 11244 18753 11255
rect 18804 11244 18837 11255
rect 18872 11244 18906 11278
rect 18940 11255 18974 11278
rect 18955 11244 18974 11255
rect 19008 11244 19042 11278
rect 19076 11244 19110 11278
rect 19144 11244 19178 11278
rect 19212 11244 19246 11278
rect 19280 11244 19314 11278
rect 19348 11244 19382 11278
rect 10304 11224 10328 11231
rect 8425 11191 8465 11224
rect 8499 11191 8539 11224
rect 8573 11191 8613 11224
rect 8647 11191 8687 11224
rect 8721 11191 8761 11224
rect 8795 11191 8835 11224
rect 8869 11191 8909 11224
rect 8943 11191 8983 11224
rect 9017 11191 9058 11224
rect 9092 11191 9133 11224
rect 9167 11191 9208 11224
rect 9242 11191 9283 11224
rect 9317 11191 9358 11224
rect 9392 11191 9433 11224
rect 9467 11191 9508 11224
rect 9542 11191 10328 11224
rect 7165 11186 10328 11191
rect 6746 11152 6770 11186
rect 6813 11185 6839 11186
rect 6901 11185 6908 11186
rect 6804 11152 6839 11185
rect 6873 11152 6908 11185
rect 6942 11185 6955 11186
rect 7011 11185 7043 11186
rect 6942 11152 6977 11185
rect 7011 11152 7046 11185
rect 7080 11152 7115 11186
rect 7165 11185 7184 11186
rect 7149 11152 7184 11185
rect 7218 11152 7253 11186
rect 7287 11152 7322 11186
rect 7356 11152 7391 11186
rect 7425 11152 7460 11186
rect 7494 11152 7529 11186
rect 7563 11152 7598 11186
rect 7632 11152 7667 11186
rect 7701 11152 7736 11186
rect 7770 11152 7805 11186
rect 7839 11152 7874 11186
rect 7908 11152 7943 11186
rect 7977 11152 8012 11186
rect 8046 11152 8081 11186
rect 8115 11152 8150 11186
rect 8184 11152 8219 11186
rect 8253 11152 8288 11186
rect 8322 11152 8357 11186
rect 8391 11152 8426 11186
rect 8460 11152 8495 11186
rect 8529 11152 8564 11186
rect 8598 11152 8633 11186
rect 8667 11152 8702 11186
rect 8736 11152 8771 11186
rect 8805 11152 8840 11186
rect 8874 11152 8909 11186
rect 8943 11152 8978 11186
rect 9012 11152 9046 11186
rect 9080 11152 9114 11186
rect 9148 11152 9182 11186
rect 9216 11152 9250 11186
rect 9284 11152 9318 11186
rect 9352 11152 9386 11186
rect 9420 11152 9454 11186
rect 9488 11152 9522 11186
rect 9556 11152 9590 11186
rect 9624 11152 9658 11186
rect 9692 11152 9726 11186
rect 9760 11152 9794 11186
rect 9828 11152 9862 11186
rect 9896 11152 9930 11186
rect 9964 11152 9998 11186
rect 10032 11152 10066 11186
rect 10100 11152 10134 11186
rect 10168 11152 10202 11186
rect 10236 11152 10270 11186
rect 10304 11152 10328 11186
rect 6746 11148 10328 11152
rect 16285 11223 17445 11244
rect 17479 11223 17525 11244
rect 17559 11223 17605 11244
rect 17639 11223 17684 11244
rect 17718 11223 17763 11244
rect 17797 11223 17842 11244
rect 17876 11223 17921 11244
rect 17955 11223 18000 11244
rect 18034 11223 18079 11244
rect 18113 11223 18158 11244
rect 18192 11223 18500 11244
rect 16285 11221 18500 11223
rect 18534 11221 18585 11244
rect 18619 11221 18669 11244
rect 18703 11221 18753 11244
rect 18787 11221 18837 11244
rect 18871 11221 18921 11244
rect 18955 11221 19382 11244
rect 16285 11206 19382 11221
rect 16285 11172 16319 11206
rect 16353 11172 16388 11206
rect 16422 11172 16457 11206
rect 16491 11172 16526 11206
rect 16560 11172 16594 11206
rect 16628 11172 16662 11206
rect 16696 11172 16730 11206
rect 16764 11172 16798 11206
rect 16832 11172 16866 11206
rect 16900 11172 16934 11206
rect 16968 11172 17002 11206
rect 17036 11172 17070 11206
rect 17104 11172 17138 11206
rect 17172 11172 17206 11206
rect 17240 11172 17274 11206
rect 17308 11172 17342 11206
rect 17376 11172 17410 11206
rect 17444 11185 17478 11206
rect 17512 11185 17546 11206
rect 17580 11185 17614 11206
rect 17444 11172 17445 11185
rect 17512 11172 17525 11185
rect 17580 11172 17605 11185
rect 17648 11172 17682 11206
rect 17716 11185 17750 11206
rect 17784 11185 17818 11206
rect 17852 11185 17886 11206
rect 17718 11172 17750 11185
rect 17797 11172 17818 11185
rect 17876 11172 17886 11185
rect 17920 11185 17954 11206
rect 17988 11185 18022 11206
rect 18056 11185 18090 11206
rect 17920 11172 17921 11185
rect 17988 11172 18000 11185
rect 18056 11172 18079 11185
rect 18124 11172 18158 11206
rect 18192 11172 18226 11206
rect 18260 11172 18294 11206
rect 18328 11172 18362 11206
rect 18396 11172 18430 11206
rect 18464 11172 18498 11206
rect 18532 11183 18566 11206
rect 18600 11183 18634 11206
rect 18534 11172 18566 11183
rect 18619 11172 18634 11183
rect 18668 11183 18702 11206
rect 18736 11183 18770 11206
rect 18804 11183 18838 11206
rect 18668 11172 18669 11183
rect 18736 11172 18753 11183
rect 18804 11172 18837 11183
rect 18872 11172 18906 11206
rect 18940 11183 18974 11206
rect 18955 11172 18974 11183
rect 19008 11172 19042 11206
rect 19076 11172 19110 11206
rect 19144 11172 19178 11206
rect 19212 11172 19246 11206
rect 19280 11172 19314 11206
rect 19348 11172 19382 11206
rect 16285 11151 17445 11172
rect 17479 11151 17525 11172
rect 17559 11151 17605 11172
rect 17639 11151 17684 11172
rect 17718 11151 17763 11172
rect 17797 11151 17842 11172
rect 17876 11151 17921 11172
rect 17955 11151 18000 11172
rect 18034 11151 18079 11172
rect 18113 11151 18158 11172
rect 18192 11151 18500 11172
rect 16285 11149 18500 11151
rect 18534 11149 18585 11172
rect 18619 11149 18669 11172
rect 18703 11149 18753 11172
rect 18787 11149 18837 11172
rect 18871 11149 18921 11172
rect 18955 11149 19382 11172
rect 6746 11147 7246 11148
rect 6746 11113 6779 11147
rect 6813 11113 6867 11147
rect 6901 11113 6955 11147
rect 6989 11113 7043 11147
rect 7077 11113 7131 11147
rect 7165 11113 7246 11147
rect 6746 11075 7246 11113
rect 6746 11072 6779 11075
rect 6813 11072 6867 11075
rect 6746 11038 6751 11072
rect 6813 11041 6827 11072
rect 6785 11038 6827 11041
rect 6861 11041 6867 11072
rect 6901 11072 6955 11075
rect 6989 11072 7043 11075
rect 7077 11072 7131 11075
rect 7165 11072 7246 11075
rect 6901 11041 6903 11072
rect 6861 11038 6903 11041
rect 6937 11041 6955 11072
rect 7013 11041 7043 11072
rect 6937 11038 6979 11041
rect 7013 11038 7055 11041
rect 7089 11038 7131 11072
rect 7165 11038 7207 11072
rect 7241 11038 7246 11072
rect 6746 11004 7246 11038
rect 6746 10970 6751 11004
rect 6785 11002 6827 11004
rect 6813 10970 6827 11002
rect 6861 11002 6903 11004
rect 6861 10970 6867 11002
rect 6746 10968 6779 10970
rect 6813 10968 6867 10970
rect 6901 10970 6903 11002
rect 6937 11002 6979 11004
rect 7013 11002 7055 11004
rect 6937 10970 6955 11002
rect 7013 10970 7043 11002
rect 7089 10970 7131 11004
rect 7165 10970 7207 11004
rect 7241 10970 7246 11004
rect 6901 10968 6955 10970
rect 6989 10968 7043 10970
rect 7077 10968 7131 10970
rect 7165 10968 7246 10970
rect 6746 10936 7246 10968
rect 6746 10902 6751 10936
rect 6785 10929 6827 10936
rect 6813 10902 6827 10929
rect 6861 10929 6903 10936
rect 6861 10902 6867 10929
rect 6746 10895 6779 10902
rect 6813 10895 6867 10902
rect 6901 10902 6903 10929
rect 6937 10929 6979 10936
rect 7013 10929 7055 10936
rect 6937 10902 6955 10929
rect 7013 10902 7043 10929
rect 7089 10902 7131 10936
rect 7165 10902 7207 10936
rect 7241 10902 7246 10936
rect 6901 10895 6955 10902
rect 6989 10895 7043 10902
rect 7077 10895 7131 10902
rect 7165 10895 7246 10902
rect 6746 10868 7246 10895
rect 6746 10834 6751 10868
rect 6785 10856 6827 10868
rect 6813 10834 6827 10856
rect 6861 10856 6903 10868
rect 6861 10834 6867 10856
rect 6746 10822 6779 10834
rect 6813 10822 6867 10834
rect 6901 10834 6903 10856
rect 6937 10856 6979 10868
rect 7013 10856 7055 10868
rect 6937 10834 6955 10856
rect 7013 10834 7043 10856
rect 7089 10834 7131 10868
rect 7165 10834 7207 10868
rect 7241 10834 7246 10868
rect 6901 10822 6955 10834
rect 6989 10822 7043 10834
rect 7077 10822 7131 10834
rect 7165 10822 7246 10834
rect 6746 10800 7246 10822
rect 6746 10766 6751 10800
rect 6785 10783 6827 10800
rect 6813 10766 6827 10783
rect 6861 10783 6903 10800
rect 6861 10766 6867 10783
rect 6746 10749 6779 10766
rect 6813 10749 6867 10766
rect 6901 10766 6903 10783
rect 6937 10783 6979 10800
rect 7013 10783 7055 10800
rect 6937 10766 6955 10783
rect 7013 10766 7043 10783
rect 7089 10766 7131 10800
rect 7165 10766 7207 10800
rect 7241 10766 7246 10800
rect 6901 10749 6955 10766
rect 6989 10749 7043 10766
rect 7077 10749 7131 10766
rect 7165 10749 7246 10766
rect 6746 10732 7246 10749
rect 6746 10698 6751 10732
rect 6785 10698 6827 10732
rect 6861 10698 6903 10732
rect 6937 10698 6979 10732
rect 7013 10698 7055 10732
rect 7089 10698 7131 10732
rect 7165 10698 7207 10732
rect 7241 10698 7246 10732
rect 6746 10696 7246 10698
rect 6746 10664 7155 10696
rect 7189 10664 7246 10696
rect 6746 10630 6751 10664
rect 6785 10630 6827 10664
rect 6861 10630 6903 10664
rect 6937 10630 6979 10664
rect 7013 10630 7055 10664
rect 7089 10630 7131 10664
rect 7189 10662 7207 10664
rect 7165 10630 7207 10662
rect 7241 10630 7246 10664
rect 6746 10620 7246 10630
rect 6746 10596 7155 10620
rect 7189 10596 7246 10620
rect 6746 10562 6751 10596
rect 6785 10562 6827 10596
rect 6861 10562 6903 10596
rect 6937 10562 6979 10596
rect 7013 10562 7055 10596
rect 7089 10562 7131 10596
rect 7189 10586 7207 10596
rect 7165 10562 7207 10586
rect 7241 10562 7246 10596
rect 6746 10544 7246 10562
rect 6746 10528 7155 10544
rect 7189 10528 7246 10544
rect 6746 10494 6751 10528
rect 6785 10494 6827 10528
rect 6861 10494 6903 10528
rect 6937 10494 6979 10528
rect 7013 10494 7055 10528
rect 7089 10494 7131 10528
rect 7189 10510 7207 10528
rect 7165 10494 7207 10510
rect 7241 10494 7246 10528
rect 6746 10468 7246 10494
rect 6746 10460 7155 10468
rect 7189 10460 7246 10468
rect 6746 10426 6751 10460
rect 6785 10426 6827 10460
rect 6861 10426 6903 10460
rect 6937 10426 6979 10460
rect 7013 10426 7055 10460
rect 7089 10426 7131 10460
rect 7189 10434 7207 10460
rect 7165 10426 7207 10434
rect 7241 10426 7246 10460
rect 6746 10392 7246 10426
rect 6746 10358 6751 10392
rect 6785 10358 6827 10392
rect 6861 10358 6903 10392
rect 6937 10358 6979 10392
rect 7013 10358 7055 10392
rect 7089 10358 7131 10392
rect 7189 10358 7207 10392
rect 7241 10358 7246 10392
rect 6746 10324 7246 10358
rect 6746 10290 6751 10324
rect 6785 10290 6827 10324
rect 6861 10290 6903 10324
rect 6937 10290 6979 10324
rect 7013 10290 7055 10324
rect 7089 10290 7131 10324
rect 7165 10316 7207 10324
rect 7189 10290 7207 10316
rect 7241 10290 7246 10324
rect 6746 10282 7155 10290
rect 7189 10282 7246 10290
rect 6746 10261 7246 10282
rect 10049 11096 10313 11148
rect 16285 11134 19382 11149
rect 16285 11100 16319 11134
rect 16353 11100 16388 11134
rect 16422 11100 16457 11134
rect 16491 11100 16526 11134
rect 16560 11100 16594 11134
rect 16628 11100 16662 11134
rect 16696 11100 16730 11134
rect 16764 11100 16798 11134
rect 16832 11100 16866 11134
rect 16900 11100 16934 11134
rect 16968 11100 17002 11134
rect 17036 11100 17070 11134
rect 17104 11100 17138 11134
rect 17172 11100 17206 11134
rect 17240 11100 17274 11134
rect 17308 11100 17342 11134
rect 17376 11100 17410 11134
rect 17444 11100 17478 11134
rect 17512 11100 17546 11134
rect 17580 11100 17614 11134
rect 17648 11100 17682 11134
rect 17716 11100 17750 11134
rect 17784 11100 17818 11134
rect 17852 11100 17886 11134
rect 17920 11100 17954 11134
rect 17988 11100 18022 11134
rect 18056 11100 18090 11134
rect 18124 11100 18158 11134
rect 18192 11100 18226 11134
rect 18260 11100 18294 11134
rect 18328 11100 18362 11134
rect 18396 11100 18430 11134
rect 18464 11100 18498 11134
rect 18532 11100 18566 11134
rect 18600 11100 18634 11134
rect 18668 11100 18702 11134
rect 18736 11100 18770 11134
rect 18804 11100 18838 11134
rect 18872 11100 18906 11134
rect 18940 11100 18974 11134
rect 19008 11100 19042 11134
rect 19076 11100 19110 11134
rect 19144 11100 19178 11134
rect 19212 11100 19246 11134
rect 19280 11100 19314 11134
rect 19348 11100 19382 11134
rect 10049 11072 10219 11096
rect 16285 11062 19382 11100
rect 16285 11028 16319 11062
rect 16353 11028 16388 11062
rect 16422 11028 16457 11062
rect 16491 11028 16526 11062
rect 16560 11028 16594 11062
rect 16628 11028 16662 11062
rect 16696 11028 16730 11062
rect 16764 11028 16798 11062
rect 16832 11028 16866 11062
rect 16900 11028 16934 11062
rect 16968 11028 17002 11062
rect 17036 11028 17070 11062
rect 17104 11028 17138 11062
rect 17172 11028 17206 11062
rect 17240 11028 17274 11062
rect 17308 11028 17342 11062
rect 17376 11028 17410 11062
rect 17444 11028 17478 11062
rect 17512 11028 17546 11062
rect 17580 11028 17614 11062
rect 17648 11028 17682 11062
rect 17716 11028 17750 11062
rect 17784 11028 17818 11062
rect 17852 11028 17886 11062
rect 17920 11028 17954 11062
rect 17988 11028 18022 11062
rect 18056 11028 18090 11062
rect 18124 11028 18158 11062
rect 18192 11028 18226 11062
rect 18260 11028 18294 11062
rect 18328 11028 18362 11062
rect 18396 11028 18430 11062
rect 18464 11028 18498 11062
rect 18532 11028 18566 11062
rect 18600 11028 18634 11062
rect 18668 11028 18702 11062
rect 18736 11028 18770 11062
rect 18804 11028 18838 11062
rect 18872 11028 18906 11062
rect 18940 11028 18974 11062
rect 19008 11028 19042 11062
rect 19076 11028 19110 11062
rect 19144 11028 19178 11062
rect 19212 11028 19246 11062
rect 19280 11028 19314 11062
rect 19348 11028 19382 11062
rect 16285 11025 19382 11028
rect 19548 11317 19650 11384
rect 19548 11283 19581 11317
rect 19615 11283 19650 11317
rect 19548 11242 19650 11283
rect 25100 11355 25528 11422
rect 25100 11321 25124 11355
rect 25158 11321 25196 11355
rect 25230 11321 25268 11355
rect 25302 11321 25340 11355
rect 25374 11321 25412 11355
rect 25446 11321 25484 11355
rect 25518 11321 25556 11355
rect 25590 11321 25627 11355
rect 25661 11321 25698 11355
rect 25732 11321 25769 11355
rect 25803 11321 25840 11355
rect 25874 11321 25911 11355
rect 25945 11321 25982 11355
rect 26016 11321 26053 11355
rect 26087 11321 26124 11355
rect 26158 11321 26195 11355
rect 26229 11321 26253 11355
rect 25100 11287 26253 11321
rect 25100 11253 25124 11287
rect 25158 11253 25196 11287
rect 25230 11253 25268 11287
rect 25302 11253 25340 11287
rect 25374 11253 25412 11287
rect 25446 11253 25484 11287
rect 25518 11253 25556 11287
rect 25590 11253 25627 11287
rect 25661 11253 25698 11287
rect 25732 11253 25769 11287
rect 25803 11253 25840 11287
rect 25874 11253 25911 11287
rect 25945 11253 25982 11287
rect 26016 11253 26053 11287
rect 26087 11253 26124 11287
rect 26158 11253 26195 11287
rect 26229 11253 26253 11287
rect 19548 11208 19581 11242
rect 19615 11208 19650 11242
rect 19548 11167 19650 11208
rect 19548 11133 19581 11167
rect 19615 11133 19650 11167
rect 19548 11091 19650 11133
rect 19548 11057 19581 11091
rect 19615 11057 19650 11091
rect 19548 11036 19650 11057
rect 6746 10256 7266 10261
rect 6746 10222 6751 10256
rect 6785 10222 6827 10256
rect 6861 10222 6903 10256
rect 6937 10222 6979 10256
rect 7013 10222 7055 10256
rect 7089 10222 7131 10256
rect 7165 10240 7207 10256
rect 7189 10222 7207 10240
rect 7241 10227 7266 10256
rect 7300 10227 7323 10261
rect 7241 10222 7323 10227
rect 6746 10206 7155 10222
rect 7189 10206 7323 10222
rect 6746 10189 7323 10206
rect 6746 10188 7266 10189
rect 6746 10154 6751 10188
rect 6785 10154 6827 10188
rect 6861 10154 6903 10188
rect 6937 10154 6979 10188
rect 7013 10154 7055 10188
rect 7089 10154 7131 10188
rect 7165 10164 7207 10188
rect 7189 10154 7207 10164
rect 7241 10155 7266 10188
rect 7300 10155 7323 10189
rect 7241 10154 7323 10155
rect 6746 10130 7155 10154
rect 7189 10130 7323 10154
rect 6746 10120 7323 10130
rect 6746 10086 6751 10120
rect 6785 10086 6827 10120
rect 6861 10086 6903 10120
rect 6937 10086 6979 10120
rect 7013 10086 7055 10120
rect 7089 10086 7131 10120
rect 7165 10088 7207 10120
rect 7189 10086 7207 10088
rect 7241 10117 7323 10120
rect 7241 10086 7266 10117
rect 6746 10054 7155 10086
rect 7189 10083 7266 10086
rect 7300 10083 7323 10117
rect 7189 10054 7323 10083
rect 6746 10052 7323 10054
rect 6746 10018 6751 10052
rect 6785 10018 6827 10052
rect 6861 10018 6903 10052
rect 6937 10018 6979 10052
rect 7013 10018 7055 10052
rect 7089 10018 7131 10052
rect 7165 10018 7207 10052
rect 7241 10045 7323 10052
rect 7241 10018 7266 10045
rect 6746 10012 7266 10018
rect 6746 9984 7155 10012
rect 7189 10011 7266 10012
rect 7300 10011 7323 10045
rect 7189 9984 7323 10011
rect 6746 9950 6751 9984
rect 6785 9950 6827 9984
rect 6861 9950 6903 9984
rect 6937 9950 6979 9984
rect 7013 9950 7055 9984
rect 7089 9950 7131 9984
rect 7189 9978 7207 9984
rect 7165 9950 7207 9978
rect 7241 9973 7323 9984
rect 7241 9950 7266 9973
rect 6746 9939 7266 9950
rect 7300 9939 7323 9973
rect 6746 9935 7323 9939
rect 6746 9916 7155 9935
rect 7189 9916 7323 9935
rect 6746 9882 6751 9916
rect 6785 9882 6827 9916
rect 6861 9882 6903 9916
rect 6937 9882 6979 9916
rect 7013 9882 7055 9916
rect 7089 9882 7131 9916
rect 7189 9901 7207 9916
rect 7165 9882 7207 9901
rect 7241 9901 7323 9916
rect 7241 9882 7266 9901
rect 6746 9867 7266 9882
rect 7300 9867 7323 9901
rect 6746 9858 7323 9867
rect 6746 9848 7155 9858
rect 7189 9848 7323 9858
rect 6746 9814 6751 9848
rect 6785 9814 6827 9848
rect 6861 9814 6903 9848
rect 6937 9814 6979 9848
rect 7013 9814 7055 9848
rect 7089 9814 7131 9848
rect 7189 9824 7207 9848
rect 7165 9814 7207 9824
rect 7241 9829 7323 9848
rect 7241 9814 7266 9829
rect 6746 9795 7266 9814
rect 7300 9795 7323 9829
rect 6746 9781 7323 9795
rect 6746 9780 7155 9781
rect 7189 9780 7323 9781
rect 6746 9746 6751 9780
rect 6785 9746 6827 9780
rect 6861 9746 6903 9780
rect 6937 9746 6979 9780
rect 7013 9746 7055 9780
rect 7089 9746 7131 9780
rect 7189 9747 7207 9780
rect 7165 9746 7207 9747
rect 7241 9757 7323 9780
rect 7241 9746 7266 9757
rect 6746 9723 7266 9746
rect 7300 9723 7323 9757
rect 6746 9712 7323 9723
rect 6746 9678 6751 9712
rect 6785 9678 6827 9712
rect 6861 9678 6903 9712
rect 6937 9678 6979 9712
rect 7013 9678 7055 9712
rect 7089 9678 7131 9712
rect 7165 9704 7207 9712
rect 7189 9678 7207 9704
rect 7241 9699 7323 9712
rect 10049 10255 10219 10290
rect 19582 11015 19616 11036
rect 19615 11002 19616 11015
rect 19548 10981 19581 11002
rect 19615 10981 19650 11002
rect 19548 10939 19650 10981
rect 19548 10933 19581 10939
rect 19615 10933 19650 10939
rect 19615 10905 19616 10933
rect 19582 10899 19616 10905
rect 19548 10863 19650 10899
rect 19548 10830 19581 10863
rect 19615 10830 19650 10863
rect 19615 10829 19616 10830
rect 19582 10796 19616 10829
rect 19548 10787 19650 10796
rect 19548 10753 19581 10787
rect 19615 10753 19650 10787
rect 19548 10727 19650 10753
rect 19582 10711 19616 10727
rect 19615 10693 19616 10711
rect 19548 10677 19581 10693
rect 19615 10677 19650 10693
rect 19548 10635 19650 10677
rect 19548 10623 19581 10635
rect 19615 10623 19650 10635
rect 19615 10601 19616 10623
rect 19582 10589 19616 10601
rect 19548 10559 19650 10589
rect 19548 10525 19581 10559
rect 19615 10525 19650 10559
rect 19548 10519 19650 10525
rect 19582 10485 19616 10519
rect 19548 10483 19650 10485
rect 19548 10449 19581 10483
rect 19615 10449 19650 10483
rect 19548 10415 19650 10449
rect 19582 10407 19616 10415
rect 19615 10381 19616 10407
rect 19548 10373 19581 10381
rect 19615 10373 19650 10381
rect 19548 10331 19650 10373
rect 19548 10311 19581 10331
rect 19615 10311 19650 10331
rect 19615 10297 19616 10311
rect 10106 10221 10117 10255
rect 10151 10221 10178 10255
rect 10049 10186 10219 10221
rect 10083 10183 10117 10186
rect 10106 10152 10117 10183
rect 10151 10183 10185 10186
rect 10151 10152 10178 10183
rect 10049 10149 10072 10152
rect 10106 10149 10178 10152
rect 10212 10149 10219 10152
rect 10049 10117 10219 10149
rect 10083 10111 10117 10117
rect 10106 10083 10117 10111
rect 10151 10111 10185 10117
rect 10151 10083 10178 10111
rect 10049 10077 10072 10083
rect 10106 10077 10178 10083
rect 10212 10077 10219 10083
rect 10049 10048 10219 10077
rect 10083 10039 10117 10048
rect 10106 10014 10117 10039
rect 10151 10039 10185 10048
rect 10151 10014 10178 10039
rect 10049 10005 10072 10014
rect 10106 10005 10178 10014
rect 10212 10005 10219 10014
rect 10049 9979 10219 10005
rect 10083 9967 10117 9979
rect 10106 9945 10117 9967
rect 10151 9967 10185 9979
rect 10151 9945 10178 9967
rect 10049 9933 10072 9945
rect 10106 9933 10178 9945
rect 10212 9933 10219 9945
rect 10049 9910 10219 9933
rect 10083 9895 10117 9910
rect 10106 9876 10117 9895
rect 10151 9895 10185 9910
rect 10151 9876 10178 9895
rect 10049 9861 10072 9876
rect 10106 9861 10178 9876
rect 10212 9861 10219 9876
rect 10049 9841 10219 9861
rect 10083 9823 10117 9841
rect 10106 9807 10117 9823
rect 10151 9823 10185 9841
rect 10151 9807 10178 9823
rect 10049 9789 10072 9807
rect 10106 9789 10178 9807
rect 10212 9789 10219 9807
rect 10049 9772 10219 9789
rect 10083 9751 10117 9772
rect 10106 9738 10117 9751
rect 10151 9751 10185 9772
rect 10151 9738 10178 9751
rect 10049 9717 10072 9738
rect 10106 9717 10178 9738
rect 10212 9717 10219 9738
rect 10049 9703 10219 9717
rect 7241 9685 7360 9699
rect 7241 9678 7266 9685
rect 6746 9670 7155 9678
rect 7189 9670 7266 9678
rect 6746 9651 7266 9670
rect 7300 9665 7360 9685
rect 7394 9665 7435 9699
rect 7469 9665 7510 9699
rect 7544 9665 7585 9699
rect 7619 9665 7660 9699
rect 7694 9665 7735 9699
rect 7769 9665 7810 9699
rect 7844 9665 7885 9699
rect 7919 9665 7960 9699
rect 7994 9665 8035 9699
rect 8069 9665 8110 9699
rect 8144 9665 8185 9699
rect 8219 9665 8260 9699
rect 8294 9665 8335 9699
rect 8369 9665 8410 9699
rect 8444 9665 8485 9699
rect 8519 9665 8559 9699
rect 8593 9665 8633 9699
rect 8667 9665 8707 9699
rect 8741 9665 8781 9699
rect 8815 9665 8855 9699
rect 8889 9665 8929 9699
rect 8963 9665 9003 9699
rect 9037 9665 9077 9699
rect 9111 9665 9151 9699
rect 10083 9678 10117 9703
rect 10106 9669 10117 9678
rect 10151 9678 10185 9703
rect 10151 9669 10178 9678
rect 7300 9651 7323 9665
rect 6746 9644 7323 9651
rect 6746 9610 6751 9644
rect 6785 9610 6827 9644
rect 6861 9610 6903 9644
rect 6937 9610 6979 9644
rect 7013 9610 7055 9644
rect 7089 9610 7131 9644
rect 7165 9627 7207 9644
rect 7189 9610 7207 9627
rect 7241 9613 7323 9644
rect 7241 9610 7266 9613
rect 6746 9593 7155 9610
rect 7189 9593 7266 9610
rect 6746 9579 7266 9593
rect 7300 9589 7323 9613
rect 10049 9644 10072 9669
rect 10106 9644 10178 9669
rect 10212 9644 10219 9669
rect 10049 9634 10219 9644
rect 10083 9605 10117 9634
rect 10106 9600 10117 9605
rect 10151 9605 10185 9634
rect 10151 9600 10178 9605
rect 7300 9588 8333 9589
rect 8367 9588 8406 9592
rect 8440 9588 8479 9592
rect 8513 9588 8553 9592
rect 8587 9588 8627 9592
rect 10049 9589 10072 9600
rect 8661 9588 10072 9589
rect 7300 9579 7332 9588
rect 6746 9576 7332 9579
rect 6746 9542 6751 9576
rect 6785 9542 6827 9576
rect 6861 9542 6903 9576
rect 6937 9542 6979 9576
rect 7013 9542 7055 9576
rect 7089 9542 7131 9576
rect 7165 9542 7207 9576
rect 7241 9554 7332 9576
rect 7366 9554 7401 9588
rect 7435 9554 7470 9588
rect 7504 9554 7539 9588
rect 7573 9554 7608 9588
rect 7642 9554 7677 9588
rect 7711 9554 7746 9588
rect 7780 9554 7815 9588
rect 7849 9582 7884 9588
rect 7849 9554 7883 9582
rect 7918 9554 7953 9588
rect 7987 9582 8022 9588
rect 7987 9554 8011 9582
rect 8056 9554 8091 9588
rect 8125 9554 8160 9588
rect 8194 9554 8229 9588
rect 8263 9554 8297 9588
rect 8331 9558 8333 9588
rect 8399 9558 8406 9588
rect 8467 9558 8479 9588
rect 8535 9558 8553 9588
rect 8603 9558 8627 9588
rect 8331 9554 8365 9558
rect 8399 9554 8433 9558
rect 8467 9554 8501 9558
rect 8535 9554 8569 9558
rect 8603 9554 8637 9558
rect 8671 9554 8705 9588
rect 8739 9554 8773 9588
rect 8807 9554 8841 9588
rect 8875 9554 8909 9588
rect 8943 9554 8977 9588
rect 9011 9554 9045 9588
rect 9079 9582 9113 9588
rect 9091 9554 9113 9582
rect 9147 9554 9181 9588
rect 9215 9582 9249 9588
rect 9219 9554 9249 9582
rect 9283 9554 9317 9588
rect 9351 9554 9385 9588
rect 9419 9554 9453 9588
rect 9487 9554 9521 9588
rect 9555 9554 9589 9588
rect 9623 9554 9657 9588
rect 9691 9554 9725 9588
rect 9759 9554 9793 9588
rect 9827 9554 9861 9588
rect 9895 9554 9929 9588
rect 9963 9571 10072 9588
rect 10106 9571 10178 9600
rect 10212 9571 10219 9600
rect 9963 9565 10219 9571
rect 9963 9554 10049 9565
rect 7241 9548 7883 9554
rect 7917 9548 8011 9554
rect 8045 9548 9057 9554
rect 9091 9548 9185 9554
rect 9219 9548 10049 9554
rect 7241 9542 10049 9548
rect 6746 9541 10049 9542
rect 6746 9508 7266 9541
rect 6746 9474 6751 9508
rect 6785 9474 6827 9508
rect 6861 9474 6903 9508
rect 6937 9474 6979 9508
rect 7013 9474 7055 9508
rect 7089 9474 7131 9508
rect 7165 9474 7207 9508
rect 7241 9507 7266 9508
rect 7300 9531 10049 9541
rect 10083 9532 10117 9565
rect 10106 9531 10117 9532
rect 10151 9532 10185 9565
rect 16563 10255 16887 10279
rect 16597 10221 16631 10255
rect 16665 10221 16699 10255
rect 16733 10221 16767 10255
rect 16801 10221 16887 10255
rect 16563 10182 16887 10221
rect 16597 10148 16631 10182
rect 16665 10148 16699 10182
rect 16733 10154 16767 10182
rect 16801 10154 16887 10182
rect 19582 10277 19616 10297
rect 19548 10255 19650 10277
rect 19548 10221 19581 10255
rect 19615 10221 19650 10255
rect 19548 10207 19650 10221
rect 19582 10179 19616 10207
rect 19615 10173 19616 10179
rect 16742 10148 16767 10154
rect 16563 10120 16708 10148
rect 16742 10120 16781 10148
rect 16815 10120 16854 10154
rect 16563 10109 16888 10120
rect 16597 10075 16631 10109
rect 16665 10075 16699 10109
rect 16733 10082 16767 10109
rect 16801 10082 16888 10109
rect 16742 10075 16767 10082
rect 16563 10048 16708 10075
rect 16742 10048 16781 10075
rect 16815 10048 16854 10082
rect 19548 10145 19581 10173
rect 19615 10145 19650 10173
rect 19548 10103 19650 10145
rect 19615 10069 19616 10103
rect 16563 10036 16887 10048
rect 16597 10002 16631 10036
rect 16665 10002 16699 10036
rect 16733 10002 16767 10036
rect 16801 10002 16887 10036
rect 16563 9962 16887 10002
rect 16597 9928 16631 9962
rect 16665 9928 16699 9962
rect 16733 9928 16767 9962
rect 16801 9928 16887 9962
rect 16563 9888 16887 9928
rect 16597 9854 16631 9888
rect 16665 9854 16699 9888
rect 16733 9854 16767 9888
rect 16801 9854 16887 9888
rect 16563 9814 16887 9854
rect 19548 10027 19650 10069
rect 19548 9999 19581 10027
rect 19615 9999 19650 10027
rect 19615 9993 19616 9999
rect 19582 9965 19616 9993
rect 19548 9951 19650 9965
rect 19548 9917 19581 9951
rect 19615 9917 19650 9951
rect 19548 9895 19650 9917
rect 19582 9861 19616 9895
rect 19548 9837 19650 9861
rect 26253 10336 26277 10370
rect 26311 10336 26348 10370
rect 26382 10336 26419 10370
rect 26453 10336 26490 10370
rect 26524 10336 26561 10370
rect 26595 10336 26632 10370
rect 26666 10336 26703 10370
rect 26737 10336 26774 10370
rect 26808 10336 26845 10370
rect 26879 10336 26916 10370
rect 26950 10336 26986 10370
rect 27020 10336 27056 10370
rect 27090 10336 27126 10370
rect 27160 10336 27196 10370
rect 27230 10336 27266 10370
rect 27300 10336 27336 10370
rect 27370 10336 27406 10370
rect 27440 10346 27974 10370
rect 27440 10341 27547 10346
rect 27581 10341 27615 10346
rect 27649 10341 27683 10346
rect 27440 10336 27501 10341
rect 26253 10332 27501 10336
rect 26253 10298 26272 10332
rect 26306 10302 26348 10332
rect 26382 10302 26424 10332
rect 26458 10302 26500 10332
rect 26534 10302 26576 10332
rect 26610 10302 26652 10332
rect 26686 10302 26727 10332
rect 26761 10302 26802 10332
rect 26836 10302 26877 10332
rect 26911 10302 26952 10332
rect 26253 10268 26277 10298
rect 26311 10268 26348 10302
rect 26382 10268 26419 10302
rect 26458 10298 26490 10302
rect 26534 10298 26561 10302
rect 26610 10298 26632 10302
rect 26686 10298 26703 10302
rect 26761 10298 26774 10302
rect 26836 10298 26845 10302
rect 26911 10298 26916 10302
rect 26453 10268 26490 10298
rect 26524 10268 26561 10298
rect 26595 10268 26632 10298
rect 26666 10268 26703 10298
rect 26737 10268 26774 10298
rect 26808 10268 26845 10298
rect 26879 10268 26916 10298
rect 26950 10298 26952 10302
rect 26986 10302 27027 10332
rect 27061 10302 27102 10332
rect 27136 10302 27177 10332
rect 27211 10302 27252 10332
rect 27286 10302 27327 10332
rect 27361 10302 27402 10332
rect 27436 10307 27501 10332
rect 27535 10312 27547 10341
rect 27607 10312 27615 10341
rect 27679 10312 27683 10341
rect 27717 10341 27751 10346
rect 27535 10307 27573 10312
rect 27607 10307 27645 10312
rect 27679 10307 27717 10312
rect 27785 10341 27819 10346
rect 27853 10341 27974 10346
rect 27785 10312 27789 10341
rect 27853 10312 27861 10341
rect 27751 10307 27789 10312
rect 27823 10307 27861 10312
rect 27895 10307 27974 10341
rect 27436 10302 27974 10307
rect 26950 10268 26986 10298
rect 27020 10298 27027 10302
rect 27090 10298 27102 10302
rect 27160 10298 27177 10302
rect 27230 10298 27252 10302
rect 27300 10298 27327 10302
rect 27370 10298 27402 10302
rect 27020 10268 27056 10298
rect 27090 10268 27126 10298
rect 27160 10268 27196 10298
rect 27230 10268 27266 10298
rect 27300 10268 27336 10298
rect 27370 10268 27406 10298
rect 27440 10277 27974 10302
rect 27440 10268 27547 10277
rect 27581 10268 27615 10277
rect 27649 10268 27683 10277
rect 26253 10260 27501 10268
rect 26253 10226 26272 10260
rect 26306 10234 26348 10260
rect 26382 10234 26424 10260
rect 26458 10234 26500 10260
rect 26534 10234 26576 10260
rect 26610 10234 26652 10260
rect 26686 10234 26727 10260
rect 26761 10234 26802 10260
rect 26836 10234 26877 10260
rect 26911 10234 26952 10260
rect 26253 10200 26277 10226
rect 26311 10200 26348 10234
rect 26382 10200 26419 10234
rect 26458 10226 26490 10234
rect 26534 10226 26561 10234
rect 26610 10226 26632 10234
rect 26686 10226 26703 10234
rect 26761 10226 26774 10234
rect 26836 10226 26845 10234
rect 26911 10226 26916 10234
rect 26453 10200 26490 10226
rect 26524 10200 26561 10226
rect 26595 10200 26632 10226
rect 26666 10200 26703 10226
rect 26737 10200 26774 10226
rect 26808 10200 26845 10226
rect 26879 10200 26916 10226
rect 26950 10226 26952 10234
rect 26986 10234 27027 10260
rect 27061 10234 27102 10260
rect 27136 10234 27177 10260
rect 27211 10234 27252 10260
rect 27286 10234 27327 10260
rect 27361 10234 27402 10260
rect 27436 10234 27501 10260
rect 27535 10243 27547 10268
rect 27607 10243 27615 10268
rect 27679 10243 27683 10268
rect 27717 10268 27751 10277
rect 27535 10234 27573 10243
rect 27607 10234 27645 10243
rect 27679 10234 27717 10243
rect 27785 10268 27819 10277
rect 27853 10268 27974 10277
rect 27785 10243 27789 10268
rect 27853 10243 27861 10268
rect 27751 10234 27789 10243
rect 27823 10234 27861 10243
rect 27895 10234 27974 10268
rect 26950 10200 26986 10226
rect 27020 10226 27027 10234
rect 27090 10226 27102 10234
rect 27160 10226 27177 10234
rect 27230 10226 27252 10234
rect 27300 10226 27327 10234
rect 27370 10226 27402 10234
rect 27020 10200 27056 10226
rect 27090 10200 27126 10226
rect 27160 10200 27196 10226
rect 27230 10200 27266 10226
rect 27300 10200 27336 10226
rect 27370 10200 27406 10226
rect 27440 10208 27974 10234
rect 27440 10200 27547 10208
rect 26253 10195 27547 10200
rect 27581 10195 27615 10208
rect 27649 10195 27683 10208
rect 26253 10188 27501 10195
rect 26253 10154 26272 10188
rect 26306 10166 26348 10188
rect 26382 10166 26424 10188
rect 26458 10166 26500 10188
rect 26534 10166 26576 10188
rect 26610 10166 26652 10188
rect 26686 10166 26727 10188
rect 26761 10166 26802 10188
rect 26836 10166 26877 10188
rect 26911 10166 26952 10188
rect 26253 10132 26277 10154
rect 26311 10132 26348 10166
rect 26382 10132 26419 10166
rect 26458 10154 26490 10166
rect 26534 10154 26561 10166
rect 26610 10154 26632 10166
rect 26686 10154 26703 10166
rect 26761 10154 26774 10166
rect 26836 10154 26845 10166
rect 26911 10154 26916 10166
rect 26453 10132 26490 10154
rect 26524 10132 26561 10154
rect 26595 10132 26632 10154
rect 26666 10132 26703 10154
rect 26737 10132 26774 10154
rect 26808 10132 26845 10154
rect 26879 10132 26916 10154
rect 26950 10154 26952 10166
rect 26986 10166 27027 10188
rect 27061 10166 27102 10188
rect 27136 10166 27177 10188
rect 27211 10166 27252 10188
rect 27286 10166 27327 10188
rect 27361 10166 27402 10188
rect 27436 10166 27501 10188
rect 26950 10132 26986 10154
rect 27020 10154 27027 10166
rect 27090 10154 27102 10166
rect 27160 10154 27177 10166
rect 27230 10154 27252 10166
rect 27300 10154 27327 10166
rect 27370 10154 27402 10166
rect 27440 10161 27501 10166
rect 27535 10174 27547 10195
rect 27607 10174 27615 10195
rect 27679 10174 27683 10195
rect 27717 10195 27751 10208
rect 27535 10161 27573 10174
rect 27607 10161 27645 10174
rect 27679 10161 27717 10174
rect 27785 10195 27819 10208
rect 27853 10195 27974 10208
rect 27785 10174 27789 10195
rect 27853 10174 27861 10195
rect 27751 10161 27789 10174
rect 27823 10161 27861 10174
rect 27895 10161 27974 10195
rect 27020 10132 27056 10154
rect 27090 10132 27126 10154
rect 27160 10132 27196 10154
rect 27230 10132 27266 10154
rect 27300 10132 27336 10154
rect 27370 10132 27406 10154
rect 27440 10139 27974 10161
rect 27440 10132 27547 10139
rect 26253 10122 27547 10132
rect 27581 10122 27615 10139
rect 27649 10122 27683 10139
rect 26253 10116 27501 10122
rect 26253 10082 26272 10116
rect 26306 10098 26348 10116
rect 26382 10098 26424 10116
rect 26458 10098 26500 10116
rect 26534 10098 26576 10116
rect 26610 10098 26652 10116
rect 26686 10098 26727 10116
rect 26761 10098 26802 10116
rect 26836 10098 26877 10116
rect 26911 10098 26952 10116
rect 26253 10064 26277 10082
rect 26311 10064 26348 10098
rect 26382 10064 26419 10098
rect 26458 10082 26490 10098
rect 26534 10082 26561 10098
rect 26610 10082 26632 10098
rect 26686 10082 26703 10098
rect 26761 10082 26774 10098
rect 26836 10082 26845 10098
rect 26911 10082 26916 10098
rect 26453 10064 26490 10082
rect 26524 10064 26561 10082
rect 26595 10064 26632 10082
rect 26666 10064 26703 10082
rect 26737 10064 26774 10082
rect 26808 10064 26845 10082
rect 26879 10064 26916 10082
rect 26950 10082 26952 10098
rect 26986 10098 27027 10116
rect 27061 10098 27102 10116
rect 27136 10098 27177 10116
rect 27211 10098 27252 10116
rect 27286 10098 27327 10116
rect 27361 10098 27402 10116
rect 27436 10098 27501 10116
rect 26950 10064 26986 10082
rect 27020 10082 27027 10098
rect 27090 10082 27102 10098
rect 27160 10082 27177 10098
rect 27230 10082 27252 10098
rect 27300 10082 27327 10098
rect 27370 10082 27402 10098
rect 27440 10088 27501 10098
rect 27535 10105 27547 10122
rect 27607 10105 27615 10122
rect 27679 10105 27683 10122
rect 27717 10122 27751 10139
rect 27535 10088 27573 10105
rect 27607 10088 27645 10105
rect 27679 10088 27717 10105
rect 27785 10122 27819 10139
rect 27853 10122 27974 10139
rect 27785 10105 27789 10122
rect 27853 10105 27861 10122
rect 27751 10088 27789 10105
rect 27823 10088 27861 10105
rect 27895 10088 27974 10122
rect 27020 10064 27056 10082
rect 27090 10064 27126 10082
rect 27160 10064 27196 10082
rect 27230 10064 27266 10082
rect 27300 10064 27336 10082
rect 27370 10064 27406 10082
rect 27440 10070 27974 10088
rect 27440 10064 27547 10070
rect 26253 10049 27547 10064
rect 27581 10049 27615 10070
rect 27649 10049 27683 10070
rect 26253 10044 27501 10049
rect 26253 10010 26272 10044
rect 26306 10030 26348 10044
rect 26382 10030 26424 10044
rect 26458 10030 26500 10044
rect 26534 10030 26576 10044
rect 26610 10030 26652 10044
rect 26686 10030 26727 10044
rect 26761 10030 26802 10044
rect 26836 10030 26877 10044
rect 26911 10030 26952 10044
rect 26253 9996 26277 10010
rect 26311 9996 26348 10030
rect 26382 9996 26419 10030
rect 26458 10010 26490 10030
rect 26534 10010 26561 10030
rect 26610 10010 26632 10030
rect 26686 10010 26703 10030
rect 26761 10010 26774 10030
rect 26836 10010 26845 10030
rect 26911 10010 26916 10030
rect 26453 9996 26490 10010
rect 26524 9996 26561 10010
rect 26595 9996 26632 10010
rect 26666 9996 26703 10010
rect 26737 9996 26774 10010
rect 26808 9996 26845 10010
rect 26879 9996 26916 10010
rect 26950 10010 26952 10030
rect 26986 10030 27027 10044
rect 27061 10030 27102 10044
rect 27136 10030 27177 10044
rect 27211 10030 27252 10044
rect 27286 10030 27327 10044
rect 27361 10030 27402 10044
rect 27436 10030 27501 10044
rect 26950 9996 26986 10010
rect 27020 10010 27027 10030
rect 27090 10010 27102 10030
rect 27160 10010 27177 10030
rect 27230 10010 27252 10030
rect 27300 10010 27327 10030
rect 27370 10010 27402 10030
rect 27440 10015 27501 10030
rect 27535 10036 27547 10049
rect 27607 10036 27615 10049
rect 27679 10036 27683 10049
rect 27717 10049 27751 10070
rect 27535 10015 27573 10036
rect 27607 10015 27645 10036
rect 27679 10015 27717 10036
rect 27785 10049 27819 10070
rect 27853 10049 27974 10070
rect 27785 10036 27789 10049
rect 27853 10036 27861 10049
rect 27751 10015 27789 10036
rect 27823 10015 27861 10036
rect 27895 10015 27974 10049
rect 27020 9996 27056 10010
rect 27090 9996 27126 10010
rect 27160 9996 27196 10010
rect 27230 9996 27266 10010
rect 27300 9996 27336 10010
rect 27370 9996 27406 10010
rect 27440 10001 27974 10015
rect 27440 9996 27547 10001
rect 26253 9976 27547 9996
rect 27581 9976 27615 10001
rect 27649 9976 27683 10001
rect 26253 9972 27501 9976
rect 26253 9938 26272 9972
rect 26306 9962 26348 9972
rect 26382 9962 26424 9972
rect 26458 9962 26500 9972
rect 26534 9962 26576 9972
rect 26610 9962 26652 9972
rect 26686 9962 26727 9972
rect 26761 9962 26802 9972
rect 26836 9962 26877 9972
rect 26911 9962 26952 9972
rect 26253 9928 26277 9938
rect 26311 9928 26348 9962
rect 26382 9928 26419 9962
rect 26458 9938 26490 9962
rect 26534 9938 26561 9962
rect 26610 9938 26632 9962
rect 26686 9938 26703 9962
rect 26761 9938 26774 9962
rect 26836 9938 26845 9962
rect 26911 9938 26916 9962
rect 26453 9928 26490 9938
rect 26524 9928 26561 9938
rect 26595 9928 26632 9938
rect 26666 9928 26703 9938
rect 26737 9928 26774 9938
rect 26808 9928 26845 9938
rect 26879 9928 26916 9938
rect 26950 9938 26952 9962
rect 26986 9962 27027 9972
rect 27061 9962 27102 9972
rect 27136 9962 27177 9972
rect 27211 9962 27252 9972
rect 27286 9962 27327 9972
rect 27361 9962 27402 9972
rect 27436 9962 27501 9972
rect 26950 9928 26986 9938
rect 27020 9938 27027 9962
rect 27090 9938 27102 9962
rect 27160 9938 27177 9962
rect 27230 9938 27252 9962
rect 27300 9938 27327 9962
rect 27370 9938 27402 9962
rect 27440 9942 27501 9962
rect 27535 9967 27547 9976
rect 27607 9967 27615 9976
rect 27679 9967 27683 9976
rect 27717 9976 27751 10001
rect 27535 9942 27573 9967
rect 27607 9942 27645 9967
rect 27679 9942 27717 9967
rect 27785 9976 27819 10001
rect 27853 9976 27974 10001
rect 27785 9967 27789 9976
rect 27853 9967 27861 9976
rect 27751 9942 27789 9967
rect 27823 9942 27861 9967
rect 27895 9942 27974 9976
rect 27020 9928 27056 9938
rect 27090 9928 27126 9938
rect 27160 9928 27196 9938
rect 27230 9928 27266 9938
rect 27300 9928 27336 9938
rect 27370 9928 27406 9938
rect 27440 9932 27974 9942
rect 27440 9928 27547 9932
rect 26253 9902 27547 9928
rect 27581 9902 27615 9932
rect 27649 9902 27683 9932
rect 26253 9900 27501 9902
rect 26253 9866 26272 9900
rect 26306 9894 26348 9900
rect 26382 9894 26424 9900
rect 26458 9894 26500 9900
rect 26534 9894 26576 9900
rect 26610 9894 26652 9900
rect 26686 9894 26727 9900
rect 26761 9894 26802 9900
rect 26836 9894 26877 9900
rect 26911 9894 26952 9900
rect 26253 9860 26277 9866
rect 26311 9860 26348 9894
rect 26382 9860 26419 9894
rect 26458 9866 26490 9894
rect 26534 9866 26561 9894
rect 26610 9866 26632 9894
rect 26686 9866 26703 9894
rect 26761 9866 26774 9894
rect 26836 9866 26845 9894
rect 26911 9866 26916 9894
rect 26453 9860 26490 9866
rect 26524 9860 26561 9866
rect 26595 9860 26632 9866
rect 26666 9860 26703 9866
rect 26737 9860 26774 9866
rect 26808 9860 26845 9866
rect 26879 9860 26916 9866
rect 26950 9866 26952 9894
rect 26986 9894 27027 9900
rect 27061 9894 27102 9900
rect 27136 9894 27177 9900
rect 27211 9894 27252 9900
rect 27286 9894 27327 9900
rect 27361 9894 27402 9900
rect 27436 9894 27501 9900
rect 26950 9860 26986 9866
rect 27020 9866 27027 9894
rect 27090 9866 27102 9894
rect 27160 9866 27177 9894
rect 27230 9866 27252 9894
rect 27300 9866 27327 9894
rect 27370 9866 27402 9894
rect 27440 9868 27501 9894
rect 27535 9898 27547 9902
rect 27607 9898 27615 9902
rect 27679 9898 27683 9902
rect 27717 9902 27751 9932
rect 27535 9868 27573 9898
rect 27607 9868 27645 9898
rect 27679 9868 27717 9898
rect 27785 9902 27819 9932
rect 27853 9902 27974 9932
rect 27785 9898 27789 9902
rect 27853 9898 27861 9902
rect 27751 9868 27789 9898
rect 27823 9868 27861 9898
rect 27895 9868 27974 9902
rect 27020 9860 27056 9866
rect 27090 9860 27126 9866
rect 27160 9860 27196 9866
rect 27230 9860 27266 9866
rect 27300 9860 27336 9866
rect 27370 9860 27406 9866
rect 27440 9863 27974 9868
rect 27440 9860 27547 9863
rect 16597 9780 16631 9814
rect 16665 9780 16699 9814
rect 16733 9780 16767 9814
rect 16801 9780 16887 9814
rect 16563 9740 16887 9780
rect 16597 9706 16631 9740
rect 16665 9706 16699 9740
rect 16733 9706 16767 9740
rect 16801 9706 16887 9740
rect 16563 9666 16887 9706
rect 16597 9632 16631 9666
rect 16665 9632 16699 9666
rect 16733 9632 16767 9666
rect 16801 9632 16887 9666
rect 16563 9592 16887 9632
rect 16597 9558 16631 9592
rect 16665 9558 16699 9592
rect 16733 9558 16767 9592
rect 16801 9558 16887 9592
rect 16563 9534 16887 9558
rect 27501 9829 27547 9860
rect 27581 9829 27615 9863
rect 27649 9829 27683 9863
rect 27717 9829 27751 9863
rect 27785 9829 27819 9863
rect 27853 9829 27974 9863
rect 27501 9828 27974 9829
rect 27535 9794 27573 9828
rect 27607 9794 27645 9828
rect 27679 9794 27717 9828
rect 27751 9794 27789 9828
rect 27823 9794 27861 9828
rect 27895 9794 27974 9828
rect 27501 9760 27547 9794
rect 27581 9760 27615 9794
rect 27649 9760 27683 9794
rect 27717 9760 27751 9794
rect 27785 9760 27819 9794
rect 27853 9760 27974 9794
rect 27501 9754 27974 9760
rect 27535 9724 27573 9754
rect 27607 9724 27645 9754
rect 27679 9724 27717 9754
rect 27535 9720 27547 9724
rect 27607 9720 27615 9724
rect 27679 9720 27683 9724
rect 27501 9690 27547 9720
rect 27581 9690 27615 9720
rect 27649 9690 27683 9720
rect 27751 9724 27789 9754
rect 27823 9724 27861 9754
rect 27717 9690 27751 9720
rect 27785 9720 27789 9724
rect 27853 9720 27861 9724
rect 27895 9720 27974 9754
rect 27785 9690 27819 9720
rect 27853 9690 27974 9720
rect 27501 9680 27974 9690
rect 27535 9654 27573 9680
rect 27607 9654 27645 9680
rect 27679 9654 27717 9680
rect 27535 9646 27547 9654
rect 27607 9646 27615 9654
rect 27679 9646 27683 9654
rect 27501 9620 27547 9646
rect 27581 9620 27615 9646
rect 27649 9620 27683 9646
rect 27751 9654 27789 9680
rect 27823 9654 27861 9680
rect 27717 9620 27751 9646
rect 27785 9646 27789 9654
rect 27853 9646 27861 9654
rect 27895 9646 27974 9680
rect 27785 9620 27819 9646
rect 27853 9620 27974 9646
rect 27501 9606 27974 9620
rect 27535 9584 27573 9606
rect 27607 9584 27645 9606
rect 27679 9584 27717 9606
rect 27535 9572 27547 9584
rect 27607 9572 27615 9584
rect 27679 9572 27683 9584
rect 27501 9550 27547 9572
rect 27581 9550 27615 9572
rect 27649 9550 27683 9572
rect 27751 9584 27789 9606
rect 27823 9584 27861 9606
rect 27717 9550 27751 9572
rect 27785 9572 27789 9584
rect 27853 9572 27861 9584
rect 27895 9572 27974 9606
rect 27785 9550 27819 9572
rect 27853 9550 27974 9572
rect 10151 9531 10178 9532
rect 7300 9520 10072 9531
rect 7300 9510 8333 9520
rect 7300 9507 7883 9510
rect 7241 9496 7883 9507
rect 7917 9496 8011 9510
rect 8045 9496 8333 9510
rect 8367 9496 8406 9520
rect 8440 9496 8479 9520
rect 8513 9496 8553 9520
rect 8587 9496 8627 9520
rect 8661 9508 10072 9520
rect 8661 9496 9057 9508
rect 9091 9496 9185 9508
rect 9219 9498 10072 9508
rect 10106 9498 10178 9531
rect 10212 9527 10219 9531
rect 27501 9532 27974 9550
rect 10212 9498 10305 9527
rect 9219 9496 10305 9498
rect 7241 9474 7332 9496
rect 6746 9469 7332 9474
rect 6746 9440 7266 9469
rect 6746 9406 6751 9440
rect 6785 9406 6827 9440
rect 6861 9406 6903 9440
rect 6937 9406 6979 9440
rect 7013 9406 7055 9440
rect 7089 9406 7131 9440
rect 7165 9406 7207 9440
rect 7241 9435 7266 9440
rect 7300 9462 7332 9469
rect 7366 9462 7401 9496
rect 7435 9462 7470 9496
rect 7504 9462 7539 9496
rect 7573 9462 7608 9496
rect 7642 9462 7677 9496
rect 7711 9462 7746 9496
rect 7780 9462 7815 9496
rect 7849 9476 7883 9496
rect 7849 9462 7884 9476
rect 7918 9462 7953 9496
rect 7987 9476 8011 9496
rect 7987 9462 8022 9476
rect 8056 9462 8091 9496
rect 8125 9462 8160 9496
rect 8194 9462 8229 9496
rect 8263 9462 8297 9496
rect 8331 9486 8333 9496
rect 8399 9486 8406 9496
rect 8467 9486 8479 9496
rect 8535 9486 8553 9496
rect 8603 9486 8627 9496
rect 8331 9462 8365 9486
rect 8399 9462 8433 9486
rect 8467 9462 8501 9486
rect 8535 9462 8569 9486
rect 8603 9462 8637 9486
rect 8671 9462 8705 9496
rect 8739 9462 8773 9496
rect 8807 9462 8841 9496
rect 8875 9462 8909 9496
rect 8943 9462 8977 9496
rect 9011 9462 9045 9496
rect 9091 9474 9113 9496
rect 9079 9462 9113 9474
rect 9147 9462 9181 9496
rect 9219 9474 9249 9496
rect 9215 9462 9249 9474
rect 9283 9462 9317 9496
rect 9351 9462 9385 9496
rect 9419 9462 9453 9496
rect 9487 9462 9521 9496
rect 9555 9462 9589 9496
rect 9623 9462 9657 9496
rect 9691 9462 9725 9496
rect 9759 9462 9793 9496
rect 9827 9462 9861 9496
rect 9895 9462 9929 9496
rect 9963 9462 10049 9496
rect 10083 9462 10117 9496
rect 10151 9462 10185 9496
rect 10219 9493 10305 9496
rect 10339 9493 10405 9527
rect 10439 9493 10505 9527
rect 10539 9493 10607 9527
rect 10219 9462 10607 9493
rect 7300 9459 10607 9462
rect 7300 9438 10072 9459
rect 7300 9435 7883 9438
rect 7241 9406 7883 9435
rect 6746 9404 7883 9406
rect 7917 9404 8011 9438
rect 8045 9434 10072 9438
rect 8045 9404 9057 9434
rect 9091 9404 9185 9434
rect 9219 9427 10072 9434
rect 10106 9427 10178 9459
rect 10212 9455 10607 9459
rect 10212 9427 10573 9455
rect 9219 9404 10049 9427
rect 10106 9425 10117 9427
rect 6746 9397 7332 9404
rect 6746 9372 7266 9397
rect 6746 9338 6751 9372
rect 6785 9338 6827 9372
rect 6861 9338 6903 9372
rect 6937 9338 6979 9372
rect 7013 9338 7055 9372
rect 7089 9338 7131 9372
rect 7165 9338 7207 9372
rect 7241 9363 7266 9372
rect 7300 9370 7332 9397
rect 7366 9370 7401 9404
rect 7435 9370 7470 9404
rect 7504 9370 7539 9404
rect 7573 9370 7608 9404
rect 7642 9370 7677 9404
rect 7711 9370 7746 9404
rect 7780 9370 7815 9404
rect 7849 9370 7884 9404
rect 7918 9370 7953 9404
rect 7987 9370 8022 9404
rect 8056 9370 8091 9404
rect 8125 9370 8160 9404
rect 8194 9370 8229 9404
rect 8263 9370 8297 9404
rect 8331 9370 8365 9404
rect 8399 9370 8433 9404
rect 8467 9370 8501 9404
rect 8535 9370 8569 9404
rect 8603 9370 8637 9404
rect 8671 9370 8705 9404
rect 8739 9370 8773 9404
rect 8807 9370 8841 9404
rect 8875 9370 8909 9404
rect 8943 9370 8977 9404
rect 9011 9370 9045 9404
rect 9091 9400 9113 9404
rect 9079 9370 9113 9400
rect 9147 9370 9181 9404
rect 9219 9400 9249 9404
rect 9215 9370 9249 9400
rect 9283 9370 9317 9404
rect 9351 9370 9385 9404
rect 9419 9370 9453 9404
rect 9487 9370 9521 9404
rect 9555 9370 9589 9404
rect 9623 9370 9657 9404
rect 9691 9370 9725 9404
rect 9759 9370 9793 9404
rect 9827 9370 9861 9404
rect 9895 9370 9929 9404
rect 9963 9393 10049 9404
rect 10083 9393 10117 9425
rect 10151 9425 10178 9427
rect 10151 9393 10185 9425
rect 10219 9421 10573 9427
rect 27535 9514 27573 9532
rect 27607 9514 27645 9532
rect 27679 9514 27717 9532
rect 27535 9498 27547 9514
rect 27607 9498 27615 9514
rect 27679 9498 27683 9514
rect 27501 9480 27547 9498
rect 27581 9480 27615 9498
rect 27649 9480 27683 9498
rect 27751 9514 27789 9532
rect 27823 9514 27861 9532
rect 27717 9480 27751 9498
rect 27785 9498 27789 9514
rect 27853 9498 27861 9514
rect 27895 9498 27974 9532
rect 27785 9480 27819 9498
rect 27853 9480 27974 9498
rect 27501 9458 27974 9480
rect 10219 9403 10607 9421
rect 10219 9393 10305 9403
rect 9963 9370 10305 9393
rect 7300 9369 10305 9370
rect 10339 9369 10377 9403
rect 10411 9369 10449 9403
rect 10483 9383 10607 9403
rect 10483 9369 10573 9383
rect 7300 9363 7323 9369
rect 7241 9338 7323 9363
rect 6746 9324 7323 9338
rect 6746 9304 7266 9324
rect 6746 9270 6751 9304
rect 6785 9270 6827 9304
rect 6861 9270 6903 9304
rect 6937 9270 6979 9304
rect 7013 9270 7055 9304
rect 7089 9270 7131 9304
rect 7165 9270 7207 9304
rect 7241 9290 7266 9304
rect 7300 9290 7323 9324
rect 7241 9270 7323 9290
rect 6746 9251 7323 9270
rect 6746 9250 7266 9251
rect 6746 9236 7028 9250
rect 7062 9236 7266 9250
rect 6746 9202 6751 9236
rect 6785 9202 6827 9236
rect 6861 9202 6903 9236
rect 6937 9202 6979 9236
rect 7013 9216 7028 9236
rect 7013 9202 7055 9216
rect 7089 9202 7131 9236
rect 7165 9202 7207 9236
rect 7241 9217 7266 9236
rect 7300 9217 7323 9251
rect 7241 9202 7323 9217
rect 6746 9178 7323 9202
rect 6746 9177 7266 9178
rect 6746 9168 7028 9177
rect 7062 9168 7266 9177
rect 6746 9134 6751 9168
rect 6785 9134 6827 9168
rect 6861 9134 6903 9168
rect 6937 9134 6979 9168
rect 7013 9143 7028 9168
rect 7013 9134 7055 9143
rect 7089 9134 7131 9168
rect 7165 9134 7207 9168
rect 7241 9144 7266 9168
rect 7300 9144 7323 9178
rect 7241 9134 7323 9144
rect 6746 9105 7323 9134
rect 6746 9103 7266 9105
rect 6746 9100 7028 9103
rect 7062 9100 7266 9103
rect 6746 9066 6751 9100
rect 6785 9066 6827 9100
rect 6861 9066 6903 9100
rect 6937 9066 6979 9100
rect 7013 9069 7028 9100
rect 7013 9066 7055 9069
rect 7089 9066 7131 9100
rect 7165 9066 7207 9100
rect 7241 9071 7266 9100
rect 7300 9071 7323 9105
rect 7241 9066 7323 9071
rect 6746 9032 7323 9066
rect 6746 8998 6751 9032
rect 6785 8998 6827 9032
rect 6861 8998 6903 9032
rect 6937 8998 6979 9032
rect 7013 9029 7055 9032
rect 7013 8998 7028 9029
rect 7089 8998 7131 9032
rect 7165 8998 7207 9032
rect 7241 8998 7266 9032
rect 7300 8998 7323 9032
rect 6746 8995 7028 8998
rect 7062 8995 7323 8998
rect 6746 8964 7323 8995
rect 6746 8930 6751 8964
rect 6785 8930 6827 8964
rect 6861 8930 6903 8964
rect 6937 8930 6979 8964
rect 7013 8955 7055 8964
rect 7013 8930 7028 8955
rect 7089 8930 7131 8964
rect 7165 8930 7207 8964
rect 7241 8959 7323 8964
rect 7241 8930 7266 8959
rect 6746 8921 7028 8930
rect 7062 8925 7266 8930
rect 7300 8925 7323 8959
rect 7062 8921 7323 8925
rect 6746 8896 7323 8921
rect 6746 8862 6751 8896
rect 6785 8862 6827 8896
rect 6861 8862 6903 8896
rect 6937 8876 6979 8896
rect 6965 8862 6979 8876
rect 7013 8876 7055 8896
rect 7013 8862 7051 8876
rect 7089 8862 7131 8896
rect 7165 8862 7207 8896
rect 7241 8886 7323 8896
rect 7241 8862 7266 8886
rect 168 8856 1846 8861
rect 168 8822 192 8856
rect 226 8822 262 8856
rect 296 8822 332 8856
rect 366 8822 402 8856
rect 436 8822 472 8856
rect 506 8822 542 8856
rect 576 8822 612 8856
rect 646 8822 682 8856
rect 716 8822 752 8856
rect 786 8822 822 8856
rect 856 8822 891 8856
rect 925 8822 960 8856
rect 994 8822 1029 8856
rect 1063 8822 1098 8856
rect 1132 8822 1167 8856
rect 1201 8822 1236 8856
rect 1270 8822 1305 8856
rect 1339 8822 1374 8856
rect 1408 8822 1443 8856
rect 1477 8822 1512 8856
rect 1546 8822 1581 8856
rect 1615 8822 1650 8856
rect 1684 8822 1719 8856
rect 1753 8822 1788 8856
rect 1822 8822 1846 8856
rect 168 8782 1846 8822
rect 168 8748 192 8782
rect 226 8748 262 8782
rect 296 8748 332 8782
rect 366 8748 402 8782
rect 436 8748 472 8782
rect 506 8748 542 8782
rect 576 8748 612 8782
rect 646 8748 682 8782
rect 716 8748 752 8782
rect 786 8748 822 8782
rect 856 8748 891 8782
rect 925 8748 960 8782
rect 994 8748 1029 8782
rect 1063 8748 1098 8782
rect 1132 8748 1167 8782
rect 1201 8748 1236 8782
rect 1270 8748 1305 8782
rect 1339 8748 1374 8782
rect 1408 8748 1443 8782
rect 1477 8748 1512 8782
rect 1546 8748 1581 8782
rect 1615 8748 1650 8782
rect 1684 8748 1719 8782
rect 1753 8748 1788 8782
rect 1822 8748 1846 8782
rect 168 8708 1846 8748
rect 168 8674 192 8708
rect 226 8674 262 8708
rect 296 8674 332 8708
rect 366 8674 402 8708
rect 436 8674 472 8708
rect 506 8674 542 8708
rect 576 8674 612 8708
rect 646 8674 682 8708
rect 716 8674 752 8708
rect 786 8674 822 8708
rect 856 8674 891 8708
rect 925 8674 960 8708
rect 994 8674 1029 8708
rect 1063 8674 1098 8708
rect 1132 8674 1167 8708
rect 1201 8674 1236 8708
rect 1270 8674 1305 8708
rect 1339 8674 1374 8708
rect 1408 8674 1443 8708
rect 1477 8674 1512 8708
rect 1546 8674 1581 8708
rect 1615 8674 1650 8708
rect 1684 8674 1719 8708
rect 1753 8674 1788 8708
rect 1822 8674 1846 8708
rect 168 8634 1846 8674
rect 168 8600 192 8634
rect 226 8600 262 8634
rect 296 8600 332 8634
rect 366 8600 402 8634
rect 436 8600 472 8634
rect 506 8600 542 8634
rect 576 8600 612 8634
rect 646 8600 682 8634
rect 716 8600 752 8634
rect 786 8600 822 8634
rect 856 8600 891 8634
rect 925 8600 960 8634
rect 994 8600 1029 8634
rect 1063 8600 1098 8634
rect 1132 8600 1167 8634
rect 1201 8600 1236 8634
rect 1270 8600 1305 8634
rect 1339 8600 1374 8634
rect 1408 8600 1443 8634
rect 1477 8600 1512 8634
rect 1546 8600 1581 8634
rect 1615 8600 1650 8634
rect 1684 8600 1719 8634
rect 1753 8600 1788 8634
rect 1822 8600 1846 8634
rect 168 8560 1846 8600
rect 168 8526 192 8560
rect 226 8526 262 8560
rect 296 8526 332 8560
rect 366 8526 402 8560
rect 436 8526 472 8560
rect 506 8526 542 8560
rect 576 8526 612 8560
rect 646 8526 682 8560
rect 716 8526 752 8560
rect 786 8526 822 8560
rect 856 8526 891 8560
rect 925 8526 960 8560
rect 994 8526 1029 8560
rect 1063 8526 1098 8560
rect 1132 8526 1167 8560
rect 1201 8526 1236 8560
rect 1270 8526 1305 8560
rect 1339 8526 1374 8560
rect 1408 8526 1443 8560
rect 1477 8526 1512 8560
rect 1546 8526 1581 8560
rect 1615 8526 1650 8560
rect 1684 8526 1719 8560
rect 1753 8526 1788 8560
rect 1822 8526 1846 8560
rect 168 8486 1846 8526
rect 168 8452 192 8486
rect 226 8452 262 8486
rect 296 8452 332 8486
rect 366 8452 402 8486
rect 436 8452 472 8486
rect 506 8452 542 8486
rect 576 8452 612 8486
rect 646 8452 682 8486
rect 716 8452 752 8486
rect 786 8452 822 8486
rect 856 8452 891 8486
rect 925 8452 960 8486
rect 994 8452 1029 8486
rect 1063 8452 1098 8486
rect 1132 8452 1167 8486
rect 1201 8452 1236 8486
rect 1270 8452 1305 8486
rect 1339 8452 1374 8486
rect 1408 8452 1443 8486
rect 1477 8452 1512 8486
rect 1546 8452 1581 8486
rect 1615 8452 1650 8486
rect 1684 8452 1719 8486
rect 1753 8452 1788 8486
rect 1822 8452 1846 8486
rect 168 8412 1846 8452
rect 168 8378 192 8412
rect 226 8378 262 8412
rect 296 8378 332 8412
rect 366 8378 402 8412
rect 436 8378 472 8412
rect 506 8378 542 8412
rect 576 8378 612 8412
rect 646 8378 682 8412
rect 716 8378 752 8412
rect 786 8378 822 8412
rect 856 8378 891 8412
rect 925 8378 960 8412
rect 994 8378 1029 8412
rect 1063 8378 1098 8412
rect 1132 8378 1167 8412
rect 1201 8378 1236 8412
rect 1270 8378 1305 8412
rect 1339 8378 1374 8412
rect 1408 8378 1443 8412
rect 1477 8378 1512 8412
rect 1546 8378 1581 8412
rect 1615 8378 1650 8412
rect 1684 8378 1719 8412
rect 1753 8378 1788 8412
rect 1822 8378 1846 8412
rect 168 8338 1846 8378
rect 168 8304 192 8338
rect 226 8304 262 8338
rect 296 8304 332 8338
rect 366 8304 402 8338
rect 436 8304 472 8338
rect 506 8304 542 8338
rect 576 8304 612 8338
rect 646 8304 682 8338
rect 716 8304 752 8338
rect 786 8304 822 8338
rect 856 8304 891 8338
rect 925 8304 960 8338
rect 994 8304 1029 8338
rect 1063 8304 1098 8338
rect 1132 8304 1167 8338
rect 1201 8304 1236 8338
rect 1270 8304 1305 8338
rect 1339 8304 1374 8338
rect 1408 8304 1443 8338
rect 1477 8304 1512 8338
rect 1546 8304 1581 8338
rect 1615 8304 1650 8338
rect 1684 8304 1719 8338
rect 1753 8304 1788 8338
rect 1822 8304 1846 8338
rect 168 8256 1846 8304
rect 6746 8842 6931 8862
rect 6965 8842 7051 8862
rect 7085 8852 7266 8862
rect 7300 8852 7323 8886
rect 7085 8842 7323 8852
rect 6746 8828 7323 8842
rect 6746 8794 6751 8828
rect 6785 8794 6827 8828
rect 6861 8794 6903 8828
rect 6937 8794 6979 8828
rect 7013 8794 7055 8828
rect 7089 8794 7131 8828
rect 7165 8794 7207 8828
rect 7241 8813 7323 8828
rect 7241 8794 7266 8813
rect 6746 8792 7266 8794
rect 6746 8760 6931 8792
rect 6965 8760 7051 8792
rect 7085 8779 7266 8792
rect 7300 8779 7323 8813
rect 7085 8760 7323 8779
rect 6746 8726 6751 8760
rect 6785 8726 6827 8760
rect 6861 8726 6903 8760
rect 6965 8758 6979 8760
rect 6937 8726 6979 8758
rect 7013 8758 7051 8760
rect 7013 8726 7055 8758
rect 7089 8726 7131 8760
rect 7165 8726 7207 8760
rect 7241 8740 7323 8760
rect 7241 8726 7266 8740
rect 6746 8708 7266 8726
rect 6746 8692 6931 8708
rect 6965 8692 7051 8708
rect 7085 8706 7266 8708
rect 7300 8706 7323 8740
rect 7085 8692 7323 8706
rect 6746 8658 6751 8692
rect 6785 8658 6827 8692
rect 6861 8658 6903 8692
rect 6965 8674 6979 8692
rect 6937 8658 6979 8674
rect 7013 8674 7051 8692
rect 7013 8658 7055 8674
rect 7089 8658 7131 8692
rect 7165 8658 7207 8692
rect 7241 8667 7323 8692
rect 7241 8658 7266 8667
rect 6746 8633 7266 8658
rect 7300 8633 7323 8667
rect 6746 8624 7323 8633
rect 6746 8590 6751 8624
rect 6785 8590 6827 8624
rect 6861 8590 6903 8624
rect 6965 8590 6979 8624
rect 7013 8590 7051 8624
rect 7089 8590 7131 8624
rect 7165 8590 7207 8624
rect 7241 8594 7323 8624
rect 7241 8590 7266 8594
rect 6746 8584 7266 8590
rect 6746 8550 6749 8584
rect 6783 8555 6851 8584
rect 6885 8560 7266 8584
rect 7300 8560 7323 8594
rect 6885 8555 7323 8560
rect 6746 8521 6751 8550
rect 6785 8521 6827 8555
rect 6885 8550 6903 8555
rect 6861 8521 6903 8550
rect 6937 8540 6979 8555
rect 6965 8521 6979 8540
rect 7013 8540 7055 8555
rect 7013 8521 7051 8540
rect 7089 8521 7131 8555
rect 7165 8521 7207 8555
rect 7241 8521 7323 8555
rect 6746 8506 6931 8521
rect 6965 8506 7051 8521
rect 7085 8506 7266 8521
rect 6746 8505 7266 8506
rect 6746 8471 6749 8505
rect 6783 8471 6851 8505
rect 6885 8497 7266 8505
rect 6885 8471 6968 8497
rect 6746 8426 6968 8471
rect 6746 8392 6749 8426
rect 6783 8392 6851 8426
rect 6885 8392 6968 8426
rect 6746 8347 6968 8392
rect 6746 8313 6749 8347
rect 6783 8313 6851 8347
rect 6885 8313 6968 8347
rect 6746 8269 6968 8313
rect 7088 8487 7266 8497
rect 7300 8487 7323 8521
rect 10449 9349 10573 9369
rect 10449 9335 10607 9349
rect 10483 9311 10607 9335
rect 10483 9301 10573 9311
rect 10449 9277 10573 9301
rect 10449 9267 10607 9277
rect 10483 9239 10607 9267
rect 10483 9233 10573 9239
rect 10449 9205 10573 9233
rect 10449 9199 10607 9205
rect 10483 9167 10607 9199
rect 10483 9165 10573 9167
rect 10449 9133 10573 9165
rect 10449 9131 10607 9133
rect 10483 9097 10607 9131
rect 10449 9095 10607 9097
rect 10449 9063 10573 9095
rect 10483 9061 10573 9063
rect 10483 9029 10607 9061
rect 10449 9023 10607 9029
rect 10449 8995 10573 9023
rect 10483 8989 10573 8995
rect 23855 9431 24068 9434
rect 23855 9397 23879 9431
rect 23913 9397 24010 9431
rect 24044 9397 24068 9431
rect 23855 9351 24068 9397
rect 23855 9317 23879 9351
rect 23913 9317 24010 9351
rect 24044 9317 24068 9351
rect 23855 9271 24068 9317
rect 23855 9237 23879 9271
rect 23913 9237 24010 9271
rect 24044 9237 24068 9271
rect 23855 9191 24068 9237
rect 23855 9157 23879 9191
rect 23913 9157 24010 9191
rect 24044 9157 24068 9191
rect 23855 9111 24068 9157
rect 23855 9077 23879 9111
rect 23913 9077 24010 9111
rect 24044 9077 24068 9111
rect 23855 9031 24068 9077
rect 23855 9006 23879 9031
rect 10483 8961 10607 8989
rect 23566 8972 23590 9006
rect 23624 8972 23659 9006
rect 23693 8972 23728 9006
rect 23762 8972 23797 9006
rect 23831 8997 23879 9006
rect 23913 8997 24010 9031
rect 24044 8997 24068 9031
rect 23831 8994 24068 8997
rect 27535 9444 27573 9458
rect 27607 9444 27645 9458
rect 27679 9444 27717 9458
rect 27535 9424 27547 9444
rect 27607 9424 27615 9444
rect 27679 9424 27683 9444
rect 27501 9410 27547 9424
rect 27581 9410 27615 9424
rect 27649 9410 27683 9424
rect 27751 9444 27789 9458
rect 27823 9444 27861 9458
rect 27717 9410 27751 9424
rect 27785 9424 27789 9444
rect 27853 9424 27861 9444
rect 27895 9424 27974 9458
rect 27785 9410 27819 9424
rect 27853 9410 27974 9424
rect 27501 9384 27974 9410
rect 27535 9374 27573 9384
rect 27607 9374 27645 9384
rect 27679 9374 27717 9384
rect 27535 9350 27547 9374
rect 27607 9350 27615 9374
rect 27679 9350 27683 9374
rect 27501 9340 27547 9350
rect 27581 9340 27615 9350
rect 27649 9340 27683 9350
rect 27751 9374 27789 9384
rect 27823 9374 27861 9384
rect 27717 9340 27751 9350
rect 27785 9350 27789 9374
rect 27853 9350 27861 9374
rect 27895 9350 27974 9384
rect 27785 9340 27819 9350
rect 27853 9340 27974 9350
rect 27501 9310 27974 9340
rect 27535 9304 27573 9310
rect 27607 9304 27645 9310
rect 27679 9304 27717 9310
rect 27535 9276 27547 9304
rect 27607 9276 27615 9304
rect 27679 9276 27683 9304
rect 27501 9270 27547 9276
rect 27581 9270 27615 9276
rect 27649 9270 27683 9276
rect 27751 9304 27789 9310
rect 27823 9304 27861 9310
rect 27717 9270 27751 9276
rect 27785 9276 27789 9304
rect 27853 9276 27861 9304
rect 27895 9276 27974 9310
rect 27785 9270 27819 9276
rect 27853 9270 27974 9276
rect 27501 9236 27974 9270
rect 27535 9234 27573 9236
rect 27607 9234 27645 9236
rect 27679 9234 27717 9236
rect 27535 9202 27547 9234
rect 27607 9202 27615 9234
rect 27679 9202 27683 9234
rect 27501 9200 27547 9202
rect 27581 9200 27615 9202
rect 27649 9200 27683 9202
rect 27751 9234 27789 9236
rect 27823 9234 27861 9236
rect 27717 9200 27751 9202
rect 27785 9202 27789 9234
rect 27853 9202 27861 9234
rect 27895 9202 27974 9236
rect 27785 9200 27819 9202
rect 27853 9200 27974 9202
rect 27501 9164 27974 9200
rect 27501 9162 27547 9164
rect 27581 9162 27615 9164
rect 27649 9162 27683 9164
rect 27535 9130 27547 9162
rect 27607 9130 27615 9162
rect 27679 9130 27683 9162
rect 27717 9162 27751 9164
rect 27535 9128 27573 9130
rect 27607 9128 27645 9130
rect 27679 9128 27717 9130
rect 27785 9162 27819 9164
rect 27853 9162 27974 9164
rect 27785 9130 27789 9162
rect 27853 9130 27861 9162
rect 27751 9128 27789 9130
rect 27823 9128 27861 9130
rect 27895 9128 27974 9162
rect 27501 9094 27974 9128
rect 27501 9088 27547 9094
rect 27581 9088 27615 9094
rect 27649 9088 27683 9094
rect 27535 9060 27547 9088
rect 27607 9060 27615 9088
rect 27679 9060 27683 9088
rect 27717 9088 27751 9094
rect 27535 9054 27573 9060
rect 27607 9054 27645 9060
rect 27679 9054 27717 9060
rect 27785 9088 27819 9094
rect 27853 9088 27974 9094
rect 27785 9060 27789 9088
rect 27853 9060 27861 9088
rect 27751 9054 27789 9060
rect 27823 9054 27861 9060
rect 27895 9054 27974 9088
rect 27501 9024 27974 9054
rect 27501 9014 27547 9024
rect 27581 9014 27615 9024
rect 27649 9014 27683 9024
rect 23831 8972 24067 8994
rect 10449 8950 10607 8961
rect 10449 8927 10573 8950
rect 10483 8916 10573 8927
rect 23832 8942 24067 8972
rect 27535 8990 27547 9014
rect 27607 8990 27615 9014
rect 27679 8990 27683 9014
rect 27717 9014 27751 9024
rect 27535 8980 27573 8990
rect 27607 8980 27645 8990
rect 27679 8980 27717 8990
rect 27785 9014 27819 9024
rect 27853 9014 27974 9024
rect 27785 8990 27789 9014
rect 27853 8990 27861 9014
rect 27751 8980 27789 8990
rect 27823 8980 27861 8990
rect 27895 8980 27974 9014
rect 27501 8954 27974 8980
rect 10483 8893 10607 8916
rect 10449 8877 10607 8893
rect 10449 8859 10573 8877
rect 10483 8843 10573 8859
rect 10483 8825 10607 8843
rect 10449 8804 10607 8825
rect 10449 8791 10573 8804
rect 10483 8770 10573 8791
rect 10483 8757 10607 8770
rect 10449 8731 10607 8757
rect 10449 8723 10573 8731
rect 10483 8697 10573 8723
rect 10483 8689 10607 8697
rect 10449 8658 10607 8689
rect 10449 8654 10573 8658
rect 10483 8624 10573 8654
rect 10483 8620 10607 8624
rect 10449 8585 10607 8620
rect 10483 8551 10573 8585
rect 20784 8939 22923 8942
rect 23832 8941 23870 8942
rect 20784 8905 20808 8939
rect 20842 8905 20883 8939
rect 20917 8905 20958 8939
rect 20992 8905 21033 8939
rect 21067 8905 21108 8939
rect 21142 8905 21183 8939
rect 21217 8905 21258 8939
rect 21292 8905 21332 8939
rect 21366 8905 21406 8939
rect 21440 8905 21480 8939
rect 21514 8908 22923 8939
rect 23846 8908 23870 8941
rect 23904 8908 23940 8942
rect 23974 8908 24010 8942
rect 24044 8908 24068 8942
rect 27501 8940 27547 8954
rect 27581 8940 27615 8954
rect 27649 8940 27683 8954
rect 21514 8905 21572 8908
rect 20784 8874 21572 8905
rect 21606 8874 21648 8908
rect 21682 8874 21724 8908
rect 21758 8874 21800 8908
rect 21834 8874 21876 8908
rect 21910 8874 21952 8908
rect 21986 8874 22027 8908
rect 22061 8874 22102 8908
rect 22136 8890 22923 8908
rect 22136 8874 22194 8890
rect 20784 8871 22194 8874
rect 20784 8837 20808 8871
rect 20842 8837 20883 8871
rect 20917 8837 20958 8871
rect 20992 8837 21033 8871
rect 21067 8837 21108 8871
rect 21142 8837 21183 8871
rect 21217 8837 21258 8871
rect 21292 8837 21332 8871
rect 21366 8837 21406 8871
rect 21440 8837 21480 8871
rect 21514 8856 22194 8871
rect 22228 8856 22269 8890
rect 22303 8856 22344 8890
rect 22378 8856 22419 8890
rect 22453 8856 22494 8890
rect 22528 8856 22569 8890
rect 22603 8856 22643 8890
rect 22677 8856 22717 8890
rect 22751 8856 22791 8890
rect 22825 8856 22865 8890
rect 22899 8856 22923 8890
rect 21514 8840 22923 8856
rect 21514 8837 21572 8840
rect 20784 8806 21572 8837
rect 21606 8806 21648 8840
rect 21682 8806 21724 8840
rect 21758 8806 21800 8840
rect 21834 8806 21876 8840
rect 21910 8806 21952 8840
rect 21986 8806 22027 8840
rect 22061 8806 22102 8840
rect 22136 8822 22923 8840
rect 22136 8806 22194 8822
rect 20784 8803 21538 8806
rect 20784 8769 20808 8803
rect 20842 8769 20883 8803
rect 20917 8769 20958 8803
rect 20992 8769 21033 8803
rect 21067 8769 21108 8803
rect 21142 8769 21183 8803
rect 21217 8769 21258 8803
rect 21292 8769 21332 8803
rect 21366 8769 21406 8803
rect 21440 8769 21480 8803
rect 21514 8769 21538 8803
rect 20784 8735 21538 8769
rect 20784 8701 20808 8735
rect 20842 8701 20883 8735
rect 20917 8701 20958 8735
rect 20992 8701 21033 8735
rect 21067 8701 21108 8735
rect 21142 8701 21183 8735
rect 21217 8701 21258 8735
rect 21292 8701 21332 8735
rect 21366 8701 21406 8735
rect 21440 8701 21480 8735
rect 21514 8701 21538 8735
rect 20784 8667 21538 8701
rect 20784 8633 20808 8667
rect 20842 8633 20883 8667
rect 20917 8633 20958 8667
rect 20992 8633 21033 8667
rect 21067 8633 21108 8667
rect 21142 8633 21183 8667
rect 21217 8633 21258 8667
rect 21292 8633 21332 8667
rect 21366 8633 21406 8667
rect 21440 8633 21480 8667
rect 21514 8633 21538 8667
rect 20784 8599 21538 8633
rect 20784 8565 20808 8599
rect 20842 8565 20883 8599
rect 20917 8565 20958 8599
rect 20992 8565 21033 8599
rect 21067 8565 21108 8599
rect 21142 8565 21183 8599
rect 21217 8565 21258 8599
rect 21292 8565 21332 8599
rect 21366 8565 21406 8599
rect 21440 8565 21480 8599
rect 21514 8565 21538 8599
rect 22170 8788 22194 8806
rect 22228 8788 22269 8822
rect 22303 8788 22344 8822
rect 22378 8788 22419 8822
rect 22453 8788 22494 8822
rect 22528 8788 22569 8822
rect 22603 8788 22643 8822
rect 22677 8788 22717 8822
rect 22751 8788 22791 8822
rect 22825 8788 22865 8822
rect 22899 8788 22923 8822
rect 22170 8754 22923 8788
rect 22170 8720 22194 8754
rect 22228 8720 22269 8754
rect 22303 8720 22344 8754
rect 22378 8720 22419 8754
rect 22453 8720 22494 8754
rect 22528 8720 22569 8754
rect 22603 8720 22643 8754
rect 22677 8720 22717 8754
rect 22751 8720 22791 8754
rect 22825 8720 22865 8754
rect 22899 8720 22923 8754
rect 22170 8686 22923 8720
rect 22170 8652 22194 8686
rect 22228 8652 22269 8686
rect 22303 8652 22344 8686
rect 22378 8652 22419 8686
rect 22453 8652 22494 8686
rect 22528 8652 22569 8686
rect 22603 8652 22643 8686
rect 22677 8652 22717 8686
rect 22751 8652 22791 8686
rect 22825 8652 22865 8686
rect 22899 8652 22923 8686
rect 22170 8618 22923 8652
rect 22170 8584 22194 8618
rect 22228 8584 22269 8618
rect 22303 8584 22344 8618
rect 22378 8584 22419 8618
rect 22453 8584 22494 8618
rect 22528 8584 22569 8618
rect 22603 8584 22643 8618
rect 22677 8584 22717 8618
rect 22751 8584 22791 8618
rect 22825 8584 22865 8618
rect 22899 8584 22923 8618
rect 27535 8920 27547 8940
rect 27607 8920 27615 8940
rect 27679 8920 27683 8940
rect 27717 8940 27751 8954
rect 27535 8906 27573 8920
rect 27607 8906 27645 8920
rect 27679 8906 27717 8920
rect 27785 8940 27819 8954
rect 27853 8940 27974 8954
rect 27785 8920 27789 8940
rect 27853 8920 27861 8940
rect 27751 8906 27789 8920
rect 27823 8906 27861 8920
rect 27895 8906 27974 8940
rect 27501 8884 27974 8906
rect 27501 8866 27547 8884
rect 27581 8866 27615 8884
rect 27649 8866 27683 8884
rect 27535 8850 27547 8866
rect 27607 8850 27615 8866
rect 27679 8850 27683 8866
rect 27717 8866 27751 8884
rect 27535 8832 27573 8850
rect 27607 8832 27645 8850
rect 27679 8832 27717 8850
rect 27785 8866 27819 8884
rect 27853 8866 27974 8884
rect 27785 8850 27789 8866
rect 27853 8850 27861 8866
rect 27751 8832 27789 8850
rect 27823 8832 27861 8850
rect 27895 8832 27974 8866
rect 27501 8814 27974 8832
rect 27501 8792 27547 8814
rect 27581 8792 27615 8814
rect 27649 8792 27683 8814
rect 27535 8780 27547 8792
rect 27607 8780 27615 8792
rect 27679 8780 27683 8792
rect 27717 8792 27751 8814
rect 27535 8758 27573 8780
rect 27607 8758 27645 8780
rect 27679 8758 27717 8780
rect 27785 8792 27819 8814
rect 27853 8792 27974 8814
rect 27785 8780 27789 8792
rect 27853 8780 27861 8792
rect 27751 8758 27789 8780
rect 27823 8758 27861 8780
rect 27895 8758 27974 8792
rect 27501 8744 27974 8758
rect 27501 8718 27547 8744
rect 27581 8718 27615 8744
rect 27649 8718 27683 8744
rect 27535 8710 27547 8718
rect 27607 8710 27615 8718
rect 27679 8710 27683 8718
rect 27717 8718 27751 8744
rect 27535 8684 27573 8710
rect 27607 8684 27645 8710
rect 27679 8684 27717 8710
rect 27785 8718 27819 8744
rect 27853 8718 27974 8744
rect 27785 8710 27789 8718
rect 27853 8710 27861 8718
rect 27751 8684 27789 8710
rect 27823 8684 27861 8710
rect 27895 8684 27974 8718
rect 27501 8674 27974 8684
rect 27501 8644 27547 8674
rect 27581 8644 27615 8674
rect 27649 8644 27683 8674
rect 27535 8640 27547 8644
rect 27607 8640 27615 8644
rect 27679 8640 27683 8644
rect 27717 8644 27751 8674
rect 27535 8610 27573 8640
rect 27607 8610 27645 8640
rect 27679 8610 27717 8640
rect 27785 8644 27819 8674
rect 27853 8644 27974 8674
rect 27785 8640 27789 8644
rect 27853 8640 27861 8644
rect 27751 8610 27789 8640
rect 27823 8610 27861 8640
rect 27895 8610 27974 8644
rect 27501 8604 27974 8610
rect 20784 8562 21538 8565
rect 27501 8570 27547 8604
rect 27581 8570 27615 8604
rect 27649 8570 27683 8604
rect 27717 8570 27751 8604
rect 27785 8570 27819 8604
rect 27853 8570 27974 8604
rect 10449 8517 10607 8551
rect 27501 8534 27974 8570
rect 7088 8463 7323 8487
rect 7122 8429 7212 8463
rect 7246 8448 7323 8463
rect 7246 8429 7266 8448
rect 7088 8414 7266 8429
rect 7300 8414 7323 8448
rect 7088 8394 7323 8414
rect 27501 8500 27547 8534
rect 27581 8500 27615 8534
rect 27649 8500 27683 8534
rect 27717 8500 27751 8534
rect 27785 8500 27819 8534
rect 27853 8500 27974 8534
rect 27501 8464 27974 8500
rect 27501 8430 27547 8464
rect 27581 8430 27615 8464
rect 27649 8430 27683 8464
rect 27717 8430 27751 8464
rect 27785 8430 27819 8464
rect 27853 8430 27974 8464
rect 27501 8406 27974 8430
rect 7122 8360 7212 8394
rect 7246 8375 7323 8394
rect 7246 8360 7266 8375
rect 7088 8341 7266 8360
rect 7300 8341 7323 8375
rect 7088 8325 7323 8341
rect 27270 8395 27974 8406
rect 27270 8361 27272 8395
rect 27306 8361 27344 8395
rect 27378 8361 27416 8395
rect 27450 8361 27488 8395
rect 27522 8361 27560 8395
rect 27594 8361 27632 8395
rect 27666 8361 27704 8395
rect 27738 8361 27776 8395
rect 27810 8361 27848 8395
rect 27882 8361 27920 8395
rect 27954 8361 27974 8395
rect 27270 8354 27974 8361
rect 7122 8291 7212 8325
rect 7246 8302 7323 8325
rect 15743 8302 15782 8336
rect 15816 8302 15855 8336
rect 15889 8302 15928 8336
rect 15962 8302 16000 8336
rect 16034 8302 16072 8336
rect 16106 8302 16144 8336
rect 16178 8302 16216 8336
rect 16250 8302 16288 8336
rect 16322 8302 16360 8336
rect 16394 8302 16432 8336
rect 16466 8302 16504 8336
rect 16538 8302 16576 8336
rect 27304 8320 27338 8354
rect 27372 8320 27406 8354
rect 27440 8320 27474 8354
rect 27508 8320 27542 8354
rect 27576 8320 27610 8354
rect 27644 8320 27678 8354
rect 27712 8320 27746 8354
rect 27780 8320 27814 8354
rect 27848 8320 27974 8354
rect 27270 8315 27974 8320
rect 7246 8291 7266 8302
rect 168 8222 175 8256
rect 209 8222 245 8256
rect 279 8222 315 8256
rect 349 8222 385 8256
rect 419 8222 455 8256
rect 489 8222 525 8256
rect 559 8222 595 8256
rect 629 8222 665 8256
rect 699 8222 735 8256
rect 769 8222 805 8256
rect 839 8235 1846 8256
rect 7088 8268 7266 8291
rect 7300 8268 7323 8302
rect 27270 8283 27272 8315
rect 27306 8283 27344 8315
rect 27378 8283 27416 8315
rect 27450 8283 27488 8315
rect 27522 8283 27560 8315
rect 27594 8283 27632 8315
rect 27666 8283 27704 8315
rect 27738 8283 27776 8315
rect 27810 8283 27848 8315
rect 27306 8281 27338 8283
rect 27378 8281 27406 8283
rect 27450 8281 27474 8283
rect 27522 8281 27542 8283
rect 27594 8281 27610 8283
rect 27666 8281 27678 8283
rect 27738 8281 27746 8283
rect 27810 8281 27814 8283
rect 7088 8256 7246 8268
rect 839 8222 846 8235
rect 168 8188 846 8222
rect 168 8154 175 8188
rect 209 8154 245 8188
rect 279 8154 315 8188
rect 349 8154 385 8188
rect 419 8154 455 8188
rect 489 8154 525 8188
rect 559 8154 595 8188
rect 629 8154 665 8188
rect 699 8154 735 8188
rect 769 8154 805 8188
rect 839 8154 846 8188
rect 168 8120 846 8154
rect 168 8086 175 8120
rect 209 8086 245 8120
rect 279 8086 315 8120
rect 349 8086 385 8120
rect 419 8086 455 8120
rect 489 8086 525 8120
rect 559 8086 595 8120
rect 629 8086 665 8120
rect 699 8086 735 8120
rect 769 8086 805 8120
rect 839 8086 846 8120
rect 168 8068 846 8086
rect 168 8052 179 8068
rect 213 8052 257 8068
rect 291 8052 335 8068
rect 369 8052 413 8068
rect 447 8052 491 8068
rect 168 8018 175 8052
rect 213 8034 245 8052
rect 291 8034 315 8052
rect 369 8034 385 8052
rect 447 8034 455 8052
rect 209 8018 245 8034
rect 279 8018 315 8034
rect 349 8018 385 8034
rect 419 8018 455 8034
rect 489 8034 491 8052
rect 525 8052 569 8068
rect 603 8052 647 8068
rect 681 8052 725 8068
rect 759 8052 803 8068
rect 837 8052 846 8068
rect 489 8018 525 8034
rect 559 8034 569 8052
rect 629 8034 647 8052
rect 699 8034 725 8052
rect 769 8034 803 8052
rect 559 8018 595 8034
rect 629 8018 665 8034
rect 699 8018 735 8034
rect 769 8018 805 8034
rect 839 8018 846 8052
rect 168 7996 846 8018
rect 168 7984 179 7996
rect 213 7984 257 7996
rect 291 7984 335 7996
rect 369 7984 413 7996
rect 447 7984 491 7996
rect 168 7950 175 7984
rect 213 7962 245 7984
rect 291 7962 315 7984
rect 369 7962 385 7984
rect 447 7962 455 7984
rect 209 7950 245 7962
rect 279 7950 315 7962
rect 349 7950 385 7962
rect 419 7950 455 7962
rect 489 7962 491 7984
rect 525 7984 569 7996
rect 603 7984 647 7996
rect 681 7984 725 7996
rect 759 7984 803 7996
rect 837 7984 846 7996
rect 489 7950 525 7962
rect 559 7962 569 7984
rect 629 7962 647 7984
rect 699 7962 725 7984
rect 769 7962 803 7984
rect 559 7950 595 7962
rect 629 7950 665 7962
rect 699 7950 735 7962
rect 769 7950 805 7962
rect 839 7950 846 7984
rect 168 7924 846 7950
rect 168 7915 179 7924
rect 213 7915 257 7924
rect 291 7915 335 7924
rect 369 7915 413 7924
rect 447 7915 491 7924
rect 168 7881 175 7915
rect 213 7890 245 7915
rect 291 7890 315 7915
rect 369 7890 385 7915
rect 447 7890 455 7915
rect 209 7881 245 7890
rect 279 7881 315 7890
rect 349 7881 385 7890
rect 419 7881 455 7890
rect 489 7890 491 7915
rect 525 7915 569 7924
rect 603 7915 647 7924
rect 681 7915 725 7924
rect 759 7915 803 7924
rect 837 7915 846 7924
rect 489 7881 525 7890
rect 559 7890 569 7915
rect 629 7890 647 7915
rect 699 7890 725 7915
rect 769 7890 803 7915
rect 559 7881 595 7890
rect 629 7881 665 7890
rect 699 7881 735 7890
rect 769 7881 805 7890
rect 839 7881 846 7915
rect 168 7852 846 7881
rect 168 7846 179 7852
rect 213 7846 257 7852
rect 291 7846 335 7852
rect 369 7846 413 7852
rect 447 7846 491 7852
rect 168 7812 175 7846
rect 213 7818 245 7846
rect 291 7818 315 7846
rect 369 7818 385 7846
rect 447 7818 455 7846
rect 209 7812 245 7818
rect 279 7812 315 7818
rect 349 7812 385 7818
rect 419 7812 455 7818
rect 489 7818 491 7846
rect 525 7846 569 7852
rect 603 7846 647 7852
rect 681 7846 725 7852
rect 759 7846 803 7852
rect 837 7846 846 7852
rect 489 7812 525 7818
rect 559 7818 569 7846
rect 629 7818 647 7846
rect 699 7818 725 7846
rect 769 7818 803 7846
rect 559 7812 595 7818
rect 629 7812 665 7818
rect 699 7812 735 7818
rect 769 7812 805 7818
rect 839 7812 846 7846
rect 168 7780 846 7812
rect 168 7777 179 7780
rect 213 7777 257 7780
rect 291 7777 335 7780
rect 369 7777 413 7780
rect 447 7777 491 7780
rect 168 7743 175 7777
rect 213 7746 245 7777
rect 291 7746 315 7777
rect 369 7746 385 7777
rect 447 7746 455 7777
rect 209 7743 245 7746
rect 279 7743 315 7746
rect 349 7743 385 7746
rect 419 7743 455 7746
rect 489 7746 491 7777
rect 525 7777 569 7780
rect 603 7777 647 7780
rect 681 7777 725 7780
rect 759 7777 803 7780
rect 837 7777 846 7780
rect 489 7743 525 7746
rect 559 7746 569 7777
rect 629 7746 647 7777
rect 699 7746 725 7777
rect 769 7746 803 7777
rect 559 7743 595 7746
rect 629 7743 665 7746
rect 699 7743 735 7746
rect 769 7743 805 7746
rect 839 7743 846 7777
rect 168 7708 846 7743
rect 168 7674 175 7708
rect 209 7707 245 7708
rect 279 7707 315 7708
rect 349 7707 385 7708
rect 419 7707 455 7708
rect 213 7674 245 7707
rect 291 7674 315 7707
rect 369 7674 385 7707
rect 447 7674 455 7707
rect 489 7707 525 7708
rect 489 7674 491 7707
rect 168 7673 179 7674
rect 213 7673 257 7674
rect 291 7673 335 7674
rect 369 7673 413 7674
rect 447 7673 491 7674
rect 559 7707 595 7708
rect 629 7707 665 7708
rect 699 7707 735 7708
rect 769 7707 805 7708
rect 559 7674 569 7707
rect 629 7674 647 7707
rect 699 7674 725 7707
rect 769 7674 803 7707
rect 839 7674 846 7708
rect 525 7673 569 7674
rect 603 7673 647 7674
rect 681 7673 725 7674
rect 759 7673 803 7674
rect 837 7673 846 7674
rect 168 7639 846 7673
rect 168 7605 175 7639
rect 209 7634 245 7639
rect 279 7634 315 7639
rect 349 7634 385 7639
rect 419 7634 455 7639
rect 213 7605 245 7634
rect 291 7605 315 7634
rect 369 7605 385 7634
rect 447 7605 455 7634
rect 489 7634 525 7639
rect 489 7605 491 7634
rect 168 7600 179 7605
rect 213 7600 257 7605
rect 291 7600 335 7605
rect 369 7600 413 7605
rect 447 7600 491 7605
rect 559 7634 595 7639
rect 629 7634 665 7639
rect 699 7634 735 7639
rect 769 7634 805 7639
rect 559 7605 569 7634
rect 629 7605 647 7634
rect 699 7605 725 7634
rect 769 7605 803 7634
rect 839 7605 846 7639
rect 525 7600 569 7605
rect 603 7600 647 7605
rect 681 7600 725 7605
rect 759 7600 803 7605
rect 837 7600 846 7605
rect 168 7570 846 7600
rect 168 7536 175 7570
rect 209 7561 245 7570
rect 279 7561 315 7570
rect 349 7561 385 7570
rect 419 7561 455 7570
rect 213 7536 245 7561
rect 291 7536 315 7561
rect 369 7536 385 7561
rect 447 7536 455 7561
rect 489 7561 525 7570
rect 489 7536 491 7561
rect 168 7527 179 7536
rect 213 7527 257 7536
rect 291 7527 335 7536
rect 369 7527 413 7536
rect 447 7527 491 7536
rect 559 7561 595 7570
rect 629 7561 665 7570
rect 699 7561 735 7570
rect 769 7561 805 7570
rect 559 7536 569 7561
rect 629 7536 647 7561
rect 699 7536 725 7561
rect 769 7536 803 7561
rect 839 7536 846 7570
rect 525 7527 569 7536
rect 603 7527 647 7536
rect 681 7527 725 7536
rect 759 7527 803 7536
rect 837 7527 846 7536
rect 168 7501 846 7527
rect 168 7467 175 7501
rect 209 7488 245 7501
rect 279 7488 315 7501
rect 349 7488 385 7501
rect 419 7488 455 7501
rect 213 7467 245 7488
rect 291 7467 315 7488
rect 369 7467 385 7488
rect 447 7467 455 7488
rect 489 7488 525 7501
rect 489 7467 491 7488
rect 168 7454 179 7467
rect 213 7454 257 7467
rect 291 7454 335 7467
rect 369 7454 413 7467
rect 447 7454 491 7467
rect 559 7488 595 7501
rect 629 7488 665 7501
rect 699 7488 735 7501
rect 769 7488 805 7501
rect 559 7467 569 7488
rect 629 7467 647 7488
rect 699 7467 725 7488
rect 769 7467 803 7488
rect 839 7467 846 7501
rect 525 7454 569 7467
rect 603 7454 647 7467
rect 681 7454 725 7467
rect 759 7454 803 7467
rect 837 7454 846 7467
rect 168 7432 846 7454
rect 168 7398 175 7432
rect 209 7415 245 7432
rect 279 7415 315 7432
rect 349 7415 385 7432
rect 419 7415 455 7432
rect 213 7398 245 7415
rect 291 7398 315 7415
rect 369 7398 385 7415
rect 447 7398 455 7415
rect 489 7415 525 7432
rect 489 7398 491 7415
rect 168 7381 179 7398
rect 213 7381 257 7398
rect 291 7381 335 7398
rect 369 7381 413 7398
rect 447 7381 491 7398
rect 559 7415 595 7432
rect 629 7415 665 7432
rect 699 7415 735 7432
rect 769 7415 805 7432
rect 559 7398 569 7415
rect 629 7398 647 7415
rect 699 7398 725 7415
rect 769 7398 803 7415
rect 839 7398 846 7432
rect 525 7381 569 7398
rect 603 7381 647 7398
rect 681 7381 725 7398
rect 759 7381 803 7398
rect 837 7381 846 7398
rect 168 7363 846 7381
rect 168 7329 175 7363
rect 209 7342 245 7363
rect 279 7342 315 7363
rect 349 7342 385 7363
rect 419 7342 455 7363
rect 213 7329 245 7342
rect 291 7329 315 7342
rect 369 7329 385 7342
rect 447 7329 455 7342
rect 489 7342 525 7363
rect 489 7329 491 7342
rect 168 7308 179 7329
rect 213 7308 257 7329
rect 291 7308 335 7329
rect 369 7308 413 7329
rect 447 7308 491 7329
rect 559 7342 595 7363
rect 629 7342 665 7363
rect 699 7342 735 7363
rect 769 7342 805 7363
rect 559 7329 569 7342
rect 629 7329 647 7342
rect 699 7329 725 7342
rect 769 7329 803 7342
rect 839 7329 846 7363
rect 525 7308 569 7329
rect 603 7308 647 7329
rect 681 7308 725 7329
rect 759 7308 803 7329
rect 837 7308 846 7329
rect 168 7294 846 7308
rect 168 7260 175 7294
rect 209 7269 245 7294
rect 279 7269 315 7294
rect 349 7269 385 7294
rect 419 7269 455 7294
rect 213 7260 245 7269
rect 291 7260 315 7269
rect 369 7260 385 7269
rect 447 7260 455 7269
rect 489 7269 525 7294
rect 489 7260 491 7269
rect 168 7235 179 7260
rect 213 7235 257 7260
rect 291 7235 335 7260
rect 369 7235 413 7260
rect 447 7235 491 7260
rect 559 7269 595 7294
rect 629 7269 665 7294
rect 699 7269 735 7294
rect 769 7269 805 7294
rect 559 7260 569 7269
rect 629 7260 647 7269
rect 699 7260 725 7269
rect 769 7260 803 7269
rect 839 7260 846 7294
rect 7122 8222 7212 8256
rect 7088 8212 7246 8222
rect 7088 8187 7091 8212
rect 7125 8178 7205 8212
rect 7239 8187 7246 8212
rect 7122 8153 7212 8178
rect 7088 8118 7246 8153
rect 7122 8084 7212 8118
rect 7088 8080 7246 8084
rect 7088 8048 7091 8080
rect 7125 8046 7205 8080
rect 7239 8048 7246 8080
rect 7122 8014 7212 8046
rect 7088 7978 7246 8014
rect 7122 7944 7212 7978
rect 7088 7908 7246 7944
rect 7122 7874 7212 7908
rect 7088 7838 7246 7874
rect 7122 7804 7212 7838
rect 7088 7768 7246 7804
rect 7122 7734 7212 7768
rect 7088 7698 7246 7734
rect 7122 7664 7212 7698
rect 7088 7628 7246 7664
rect 27304 8249 27338 8281
rect 27372 8249 27406 8281
rect 27440 8249 27474 8281
rect 27508 8249 27542 8281
rect 27576 8249 27610 8281
rect 27644 8249 27678 8281
rect 27712 8249 27746 8281
rect 27780 8249 27814 8281
rect 27882 8281 27920 8315
rect 27954 8281 27974 8315
rect 27848 8249 27974 8281
rect 27270 8235 27974 8249
rect 27270 8212 27272 8235
rect 27306 8212 27344 8235
rect 27378 8212 27416 8235
rect 27450 8212 27488 8235
rect 27522 8212 27560 8235
rect 27594 8212 27632 8235
rect 27666 8212 27704 8235
rect 27738 8212 27776 8235
rect 27810 8212 27848 8235
rect 27306 8201 27338 8212
rect 27378 8201 27406 8212
rect 27450 8201 27474 8212
rect 27522 8201 27542 8212
rect 27594 8201 27610 8212
rect 27666 8201 27678 8212
rect 27738 8201 27746 8212
rect 27810 8201 27814 8212
rect 27304 8178 27338 8201
rect 27372 8178 27406 8201
rect 27440 8178 27474 8201
rect 27508 8178 27542 8201
rect 27576 8178 27610 8201
rect 27644 8178 27678 8201
rect 27712 8178 27746 8201
rect 27780 8178 27814 8201
rect 27882 8201 27920 8235
rect 27954 8201 27974 8235
rect 27848 8178 27974 8201
rect 27270 8155 27974 8178
rect 27270 8141 27272 8155
rect 27306 8141 27344 8155
rect 27378 8141 27416 8155
rect 27450 8141 27488 8155
rect 27522 8141 27560 8155
rect 27594 8141 27632 8155
rect 27666 8141 27704 8155
rect 27738 8141 27776 8155
rect 27810 8141 27848 8155
rect 27306 8121 27338 8141
rect 27378 8121 27406 8141
rect 27450 8121 27474 8141
rect 27522 8121 27542 8141
rect 27594 8121 27610 8141
rect 27666 8121 27678 8141
rect 27738 8121 27746 8141
rect 27810 8121 27814 8141
rect 27304 8107 27338 8121
rect 27372 8107 27406 8121
rect 27440 8107 27474 8121
rect 27508 8107 27542 8121
rect 27576 8107 27610 8121
rect 27644 8107 27678 8121
rect 27712 8107 27746 8121
rect 27780 8107 27814 8121
rect 27882 8121 27920 8155
rect 27954 8121 27974 8155
rect 27848 8107 27974 8121
rect 27270 8074 27974 8107
rect 27270 8070 27272 8074
rect 27306 8070 27344 8074
rect 27378 8070 27416 8074
rect 27450 8070 27488 8074
rect 27522 8070 27560 8074
rect 27594 8070 27632 8074
rect 27666 8070 27704 8074
rect 27738 8070 27776 8074
rect 27810 8070 27848 8074
rect 27306 8040 27338 8070
rect 27378 8040 27406 8070
rect 27450 8040 27474 8070
rect 27522 8040 27542 8070
rect 27594 8040 27610 8070
rect 27666 8040 27678 8070
rect 27738 8040 27746 8070
rect 27810 8040 27814 8070
rect 27304 8036 27338 8040
rect 27372 8036 27406 8040
rect 27440 8036 27474 8040
rect 27508 8036 27542 8040
rect 27576 8036 27610 8040
rect 27644 8036 27678 8040
rect 27712 8036 27746 8040
rect 27780 8036 27814 8040
rect 27882 8040 27920 8074
rect 27954 8040 27974 8074
rect 27848 8036 27974 8040
rect 27270 7999 27974 8036
rect 27304 7993 27338 7999
rect 27372 7993 27406 7999
rect 27440 7993 27474 7999
rect 27508 7993 27542 7999
rect 27576 7993 27610 7999
rect 27644 7993 27678 7999
rect 27712 7993 27746 7999
rect 27780 7993 27814 7999
rect 27306 7965 27338 7993
rect 27378 7965 27406 7993
rect 27450 7965 27474 7993
rect 27522 7965 27542 7993
rect 27594 7965 27610 7993
rect 27666 7965 27678 7993
rect 27738 7965 27746 7993
rect 27810 7965 27814 7993
rect 27848 7993 27974 7999
rect 27270 7959 27272 7965
rect 27306 7959 27344 7965
rect 27378 7959 27416 7965
rect 27450 7959 27488 7965
rect 27522 7959 27560 7965
rect 27594 7959 27632 7965
rect 27666 7959 27704 7965
rect 27738 7959 27776 7965
rect 27810 7959 27848 7965
rect 27882 7959 27920 7993
rect 27954 7959 27974 7993
rect 27270 7928 27974 7959
rect 27304 7912 27338 7928
rect 27372 7912 27406 7928
rect 27440 7912 27474 7928
rect 27508 7912 27542 7928
rect 27576 7912 27610 7928
rect 27644 7912 27678 7928
rect 27712 7912 27746 7928
rect 27780 7912 27814 7928
rect 27306 7894 27338 7912
rect 27378 7894 27406 7912
rect 27450 7894 27474 7912
rect 27522 7894 27542 7912
rect 27594 7894 27610 7912
rect 27666 7894 27678 7912
rect 27738 7894 27746 7912
rect 27810 7894 27814 7912
rect 27848 7912 27974 7928
rect 27270 7878 27272 7894
rect 27306 7878 27344 7894
rect 27378 7878 27416 7894
rect 27450 7878 27488 7894
rect 27522 7878 27560 7894
rect 27594 7878 27632 7894
rect 27666 7878 27704 7894
rect 27738 7878 27776 7894
rect 27810 7878 27848 7894
rect 27882 7878 27920 7912
rect 27954 7878 27974 7912
rect 27270 7857 27974 7878
rect 27304 7831 27338 7857
rect 27372 7831 27406 7857
rect 27440 7831 27474 7857
rect 27508 7831 27542 7857
rect 27576 7831 27610 7857
rect 27644 7831 27678 7857
rect 27712 7831 27746 7857
rect 27780 7831 27814 7857
rect 27306 7823 27338 7831
rect 27378 7823 27406 7831
rect 27450 7823 27474 7831
rect 27522 7823 27542 7831
rect 27594 7823 27610 7831
rect 27666 7823 27678 7831
rect 27738 7823 27746 7831
rect 27810 7823 27814 7831
rect 27848 7831 27974 7857
rect 27270 7797 27272 7823
rect 27306 7797 27344 7823
rect 27378 7797 27416 7823
rect 27450 7797 27488 7823
rect 27522 7797 27560 7823
rect 27594 7797 27632 7823
rect 27666 7797 27704 7823
rect 27738 7797 27776 7823
rect 27810 7797 27848 7823
rect 27882 7797 27920 7831
rect 27954 7797 27974 7831
rect 27270 7786 27974 7797
rect 27304 7752 27338 7786
rect 27372 7752 27406 7786
rect 27440 7752 27474 7786
rect 27508 7752 27542 7786
rect 27576 7752 27610 7786
rect 27644 7752 27678 7786
rect 27712 7752 27746 7786
rect 27780 7752 27814 7786
rect 27848 7752 27974 7786
rect 27270 7750 27974 7752
rect 27270 7716 27272 7750
rect 27306 7716 27344 7750
rect 27378 7716 27416 7750
rect 27450 7716 27488 7750
rect 27522 7716 27560 7750
rect 27594 7716 27632 7750
rect 27666 7716 27704 7750
rect 27738 7716 27776 7750
rect 27810 7716 27848 7750
rect 27882 7716 27920 7750
rect 27954 7716 27974 7750
rect 27270 7714 27974 7716
rect 27304 7680 27338 7714
rect 27372 7680 27406 7714
rect 27440 7680 27474 7714
rect 27508 7680 27542 7714
rect 27576 7680 27610 7714
rect 27644 7680 27678 7714
rect 27712 7680 27746 7714
rect 27780 7680 27814 7714
rect 27848 7680 27974 7714
rect 27270 7656 27974 7680
rect 7122 7594 7212 7628
rect 7088 7558 7246 7594
rect 7122 7524 7212 7558
rect 7088 7488 7246 7524
rect 7122 7454 7212 7488
rect 7088 7418 7246 7454
rect 7122 7384 7212 7418
rect 7088 7348 7246 7384
rect 7122 7314 7212 7348
rect 7088 7280 7246 7314
rect 525 7235 569 7260
rect 603 7235 647 7260
rect 681 7235 725 7260
rect 759 7235 803 7260
rect 837 7235 846 7260
rect 168 7225 846 7235
rect 168 7191 175 7225
rect 209 7196 245 7225
rect 279 7196 315 7225
rect 349 7196 385 7225
rect 419 7196 455 7225
rect 213 7191 245 7196
rect 291 7191 315 7196
rect 369 7191 385 7196
rect 447 7191 455 7196
rect 489 7196 525 7225
rect 489 7191 491 7196
rect 168 7162 179 7191
rect 213 7162 257 7191
rect 291 7162 335 7191
rect 369 7162 413 7191
rect 447 7162 491 7191
rect 559 7196 595 7225
rect 629 7196 665 7225
rect 699 7196 735 7225
rect 769 7196 805 7225
rect 559 7191 569 7196
rect 629 7191 647 7196
rect 699 7191 725 7196
rect 769 7191 803 7196
rect 839 7191 846 7225
rect 525 7162 569 7191
rect 603 7162 647 7191
rect 681 7162 725 7191
rect 759 7162 803 7191
rect 837 7162 846 7191
rect 168 7156 846 7162
rect 168 7122 175 7156
rect 209 7123 245 7156
rect 279 7123 315 7156
rect 349 7123 385 7156
rect 419 7123 455 7156
rect 213 7122 245 7123
rect 291 7122 315 7123
rect 369 7122 385 7123
rect 447 7122 455 7123
rect 489 7123 525 7156
rect 489 7122 491 7123
rect 168 7089 179 7122
rect 213 7089 257 7122
rect 291 7089 335 7122
rect 369 7089 413 7122
rect 447 7089 491 7122
rect 559 7123 595 7156
rect 629 7123 665 7156
rect 699 7123 735 7156
rect 769 7123 805 7156
rect 559 7122 569 7123
rect 629 7122 647 7123
rect 699 7122 725 7123
rect 769 7122 803 7123
rect 839 7122 846 7156
rect 525 7089 569 7122
rect 603 7089 647 7122
rect 681 7089 725 7122
rect 759 7089 803 7122
rect 837 7089 846 7122
rect 168 7087 846 7089
rect 168 7053 175 7087
rect 209 7053 245 7087
rect 279 7053 315 7087
rect 349 7053 385 7087
rect 419 7053 455 7087
rect 489 7053 525 7087
rect 559 7053 595 7087
rect 629 7053 665 7087
rect 699 7053 735 7087
rect 769 7053 805 7087
rect 839 7053 846 7087
rect 168 7050 846 7053
rect 168 7018 179 7050
rect 213 7018 257 7050
rect 291 7018 335 7050
rect 369 7018 413 7050
rect 447 7018 491 7050
rect 168 6984 175 7018
rect 213 7016 245 7018
rect 291 7016 315 7018
rect 369 7016 385 7018
rect 447 7016 455 7018
rect 209 6984 245 7016
rect 279 6984 315 7016
rect 349 6984 385 7016
rect 419 6984 455 7016
rect 489 7016 491 7018
rect 525 7018 569 7050
rect 603 7018 647 7050
rect 681 7018 725 7050
rect 759 7018 803 7050
rect 837 7018 846 7050
rect 489 6984 525 7016
rect 559 7016 569 7018
rect 629 7016 647 7018
rect 699 7016 725 7018
rect 769 7016 803 7018
rect 559 6984 595 7016
rect 629 6984 665 7016
rect 699 6984 735 7016
rect 769 6984 805 7016
rect 839 6984 846 7018
rect 168 6977 846 6984
rect 168 6949 179 6977
rect 213 6949 257 6977
rect 291 6949 335 6977
rect 369 6949 413 6977
rect 447 6949 491 6977
rect 168 6915 175 6949
rect 213 6943 245 6949
rect 291 6943 315 6949
rect 369 6943 385 6949
rect 447 6943 455 6949
rect 209 6915 245 6943
rect 279 6915 315 6943
rect 349 6915 385 6943
rect 419 6915 455 6943
rect 489 6943 491 6949
rect 525 6949 569 6977
rect 603 6949 647 6977
rect 681 6949 725 6977
rect 759 6949 803 6977
rect 837 6949 846 6977
rect 489 6915 525 6943
rect 559 6943 569 6949
rect 629 6943 647 6949
rect 699 6943 725 6949
rect 769 6943 803 6949
rect 559 6915 595 6943
rect 629 6915 665 6943
rect 699 6915 735 6943
rect 769 6915 805 6943
rect 839 6915 846 6949
rect 14257 7013 14263 7037
rect 14441 7013 14763 7037
rect 15085 7013 15093 7037
rect 14257 6979 14262 7013
rect 14441 6979 14478 7013
rect 14512 6979 14550 7013
rect 14584 6979 14622 7013
rect 14656 6979 14694 7013
rect 14728 6979 14763 7013
rect 15088 6979 15093 7013
rect 14257 6940 14263 6979
rect 14441 6940 14763 6979
rect 15085 6940 15093 6979
rect 14257 6930 14262 6940
rect 168 6904 846 6915
rect 168 6880 179 6904
rect 213 6880 257 6904
rect 291 6880 335 6904
rect 369 6880 413 6904
rect 447 6880 491 6904
rect 168 6846 175 6880
rect 213 6870 245 6880
rect 291 6870 315 6880
rect 369 6870 385 6880
rect 447 6870 455 6880
rect 209 6846 245 6870
rect 279 6846 315 6870
rect 349 6846 385 6870
rect 419 6846 455 6870
rect 489 6870 491 6880
rect 525 6880 569 6904
rect 603 6880 647 6904
rect 681 6880 725 6904
rect 759 6880 803 6904
rect 837 6880 846 6904
rect 489 6846 525 6870
rect 559 6870 569 6880
rect 629 6870 647 6880
rect 699 6870 725 6880
rect 769 6870 803 6880
rect 559 6846 595 6870
rect 629 6846 665 6870
rect 699 6846 735 6870
rect 769 6846 805 6870
rect 839 6846 846 6880
rect 168 6831 846 6846
rect 168 6811 179 6831
rect 213 6811 257 6831
rect 291 6811 335 6831
rect 369 6811 413 6831
rect 447 6811 491 6831
rect 168 6777 175 6811
rect 213 6797 245 6811
rect 291 6797 315 6811
rect 369 6797 385 6811
rect 447 6797 455 6811
rect 209 6777 245 6797
rect 279 6777 315 6797
rect 349 6777 385 6797
rect 419 6777 455 6797
rect 489 6797 491 6811
rect 525 6811 569 6831
rect 603 6811 647 6831
rect 681 6811 725 6831
rect 759 6811 803 6831
rect 837 6811 846 6831
rect 489 6777 525 6797
rect 559 6797 569 6811
rect 629 6797 647 6811
rect 699 6797 725 6811
rect 769 6797 803 6811
rect 559 6777 595 6797
rect 629 6777 665 6797
rect 699 6777 735 6797
rect 769 6777 805 6797
rect 839 6777 846 6811
rect 168 6758 846 6777
rect 168 6742 179 6758
rect 213 6742 257 6758
rect 291 6742 335 6758
rect 369 6742 413 6758
rect 447 6742 491 6758
rect 168 6708 175 6742
rect 213 6724 245 6742
rect 291 6724 315 6742
rect 369 6724 385 6742
rect 447 6724 455 6742
rect 209 6708 245 6724
rect 279 6708 315 6724
rect 349 6708 385 6724
rect 419 6708 455 6724
rect 489 6724 491 6742
rect 525 6742 569 6758
rect 603 6742 647 6758
rect 681 6742 725 6758
rect 759 6742 803 6758
rect 837 6742 846 6758
rect 489 6708 525 6724
rect 559 6724 569 6742
rect 629 6724 647 6742
rect 699 6724 725 6742
rect 769 6724 803 6742
rect 559 6708 595 6724
rect 629 6708 665 6724
rect 699 6708 735 6724
rect 769 6708 805 6724
rect 839 6708 846 6742
rect 168 6685 846 6708
rect 168 6673 179 6685
rect 213 6673 257 6685
rect 291 6673 335 6685
rect 369 6673 413 6685
rect 447 6673 491 6685
rect 168 6639 175 6673
rect 213 6651 245 6673
rect 291 6651 315 6673
rect 369 6651 385 6673
rect 447 6651 455 6673
rect 209 6639 245 6651
rect 279 6639 315 6651
rect 349 6639 385 6651
rect 419 6639 455 6651
rect 489 6651 491 6673
rect 525 6673 569 6685
rect 603 6673 647 6685
rect 681 6673 725 6685
rect 759 6673 803 6685
rect 837 6673 846 6685
rect 489 6639 525 6651
rect 559 6651 569 6673
rect 629 6651 647 6673
rect 699 6651 725 6673
rect 769 6651 803 6673
rect 559 6639 595 6651
rect 629 6639 665 6651
rect 699 6639 735 6651
rect 769 6639 805 6651
rect 839 6639 846 6673
rect 168 6612 846 6639
rect 168 6604 179 6612
rect 213 6604 257 6612
rect 291 6604 335 6612
rect 369 6604 413 6612
rect 447 6604 491 6612
rect 168 6570 175 6604
rect 213 6578 245 6604
rect 291 6578 315 6604
rect 369 6578 385 6604
rect 447 6578 455 6604
rect 209 6570 245 6578
rect 279 6570 315 6578
rect 349 6570 385 6578
rect 419 6570 455 6578
rect 489 6578 491 6604
rect 525 6604 569 6612
rect 603 6604 647 6612
rect 681 6604 725 6612
rect 759 6604 803 6612
rect 837 6604 846 6612
rect 489 6570 525 6578
rect 559 6578 569 6604
rect 629 6578 647 6604
rect 699 6578 725 6604
rect 769 6578 803 6604
rect 559 6570 595 6578
rect 629 6570 665 6578
rect 699 6570 735 6578
rect 769 6570 805 6578
rect 839 6570 846 6604
rect 168 6539 846 6570
rect 168 6535 179 6539
rect 213 6535 257 6539
rect 291 6535 335 6539
rect 369 6535 413 6539
rect 447 6535 491 6539
rect 168 6501 175 6535
rect 213 6505 245 6535
rect 291 6505 315 6535
rect 369 6505 385 6535
rect 447 6505 455 6535
rect 209 6501 245 6505
rect 279 6501 315 6505
rect 349 6501 385 6505
rect 419 6501 455 6505
rect 489 6505 491 6535
rect 525 6535 569 6539
rect 603 6535 647 6539
rect 681 6535 725 6539
rect 759 6535 803 6539
rect 837 6535 846 6539
rect 489 6501 525 6505
rect 559 6505 569 6535
rect 629 6505 647 6535
rect 699 6505 725 6535
rect 769 6505 803 6535
rect 559 6501 595 6505
rect 629 6501 665 6505
rect 699 6501 735 6505
rect 769 6501 805 6505
rect 839 6501 846 6535
rect 168 6466 846 6501
rect 168 6432 175 6466
rect 213 6432 245 6466
rect 291 6432 315 6466
rect 369 6432 385 6466
rect 447 6432 455 6466
rect 489 6432 491 6466
rect 559 6432 569 6466
rect 629 6432 647 6466
rect 699 6432 725 6466
rect 769 6432 803 6466
rect 839 6432 846 6466
rect 168 6397 846 6432
rect 168 6363 175 6397
rect 209 6393 245 6397
rect 279 6393 315 6397
rect 349 6393 385 6397
rect 419 6393 455 6397
rect 213 6363 245 6393
rect 291 6363 315 6393
rect 369 6363 385 6393
rect 447 6363 455 6393
rect 489 6393 525 6397
rect 489 6363 491 6393
rect 168 6359 179 6363
rect 213 6359 257 6363
rect 291 6359 335 6363
rect 369 6359 413 6363
rect 447 6359 491 6363
rect 559 6393 595 6397
rect 629 6393 665 6397
rect 699 6393 735 6397
rect 769 6393 805 6397
rect 559 6363 569 6393
rect 629 6363 647 6393
rect 699 6363 725 6393
rect 769 6363 803 6393
rect 839 6363 846 6397
rect 525 6359 569 6363
rect 603 6359 647 6363
rect 681 6359 725 6363
rect 759 6359 803 6363
rect 837 6359 846 6363
rect 168 6328 846 6359
rect 168 6294 175 6328
rect 209 6320 245 6328
rect 279 6320 315 6328
rect 349 6320 385 6328
rect 419 6320 455 6328
rect 213 6294 245 6320
rect 291 6294 315 6320
rect 369 6294 385 6320
rect 447 6294 455 6320
rect 489 6320 525 6328
rect 489 6294 491 6320
rect 168 6286 179 6294
rect 213 6286 257 6294
rect 291 6286 335 6294
rect 369 6286 413 6294
rect 447 6286 491 6294
rect 559 6320 595 6328
rect 629 6320 665 6328
rect 699 6320 735 6328
rect 769 6320 805 6328
rect 559 6294 569 6320
rect 629 6294 647 6320
rect 699 6294 725 6320
rect 769 6294 803 6320
rect 839 6294 846 6328
rect 525 6286 569 6294
rect 603 6286 647 6294
rect 681 6286 725 6294
rect 759 6286 803 6294
rect 837 6286 846 6294
rect 13030 6923 14262 6930
rect 13030 6889 13054 6923
rect 13088 6889 13123 6923
rect 13157 6889 13192 6923
rect 13226 6889 13261 6923
rect 13295 6889 13330 6923
rect 13364 6889 13399 6923
rect 13433 6889 13467 6923
rect 13501 6889 13535 6923
rect 13569 6889 13603 6923
rect 13637 6889 13671 6923
rect 13705 6889 13739 6923
rect 13773 6889 13807 6923
rect 13841 6889 13875 6923
rect 13909 6889 13943 6923
rect 13977 6889 14011 6923
rect 14045 6889 14079 6923
rect 14113 6889 14147 6923
rect 14181 6906 14262 6923
rect 14441 6906 14478 6940
rect 14512 6906 14550 6940
rect 14584 6906 14622 6940
rect 14656 6906 14694 6940
rect 14728 6906 14763 6940
rect 15088 6906 15093 6940
rect 14181 6889 14263 6906
rect 13030 6866 14263 6889
rect 14441 6866 14763 6906
rect 15085 6866 15093 6906
rect 13030 6849 14262 6866
rect 13030 6815 13054 6849
rect 13088 6815 13123 6849
rect 13157 6828 13192 6849
rect 13226 6828 13261 6849
rect 13157 6815 13187 6828
rect 13226 6815 13260 6828
rect 13295 6815 13330 6849
rect 13364 6828 13399 6849
rect 13433 6828 13467 6849
rect 13501 6828 13535 6849
rect 13569 6828 13603 6849
rect 13637 6828 13671 6849
rect 13705 6828 13739 6849
rect 13773 6828 13807 6849
rect 13841 6828 13875 6849
rect 13367 6815 13399 6828
rect 13440 6815 13467 6828
rect 13513 6815 13535 6828
rect 13586 6815 13603 6828
rect 13658 6815 13671 6828
rect 13730 6815 13739 6828
rect 13802 6815 13807 6828
rect 13874 6815 13875 6828
rect 13909 6828 13943 6849
rect 13909 6815 13912 6828
rect 13977 6815 14011 6849
rect 14045 6815 14079 6849
rect 14113 6815 14147 6849
rect 14181 6832 14262 6849
rect 14441 6832 14478 6866
rect 14512 6832 14550 6866
rect 14584 6832 14622 6866
rect 14656 6832 14694 6866
rect 14728 6832 14763 6866
rect 15088 6832 15093 6866
rect 14181 6815 14263 6832
rect 13030 6794 13187 6815
rect 13221 6794 13260 6815
rect 13294 6794 13333 6815
rect 13367 6794 13406 6815
rect 13440 6794 13479 6815
rect 13513 6794 13552 6815
rect 13586 6794 13624 6815
rect 13658 6794 13696 6815
rect 13730 6794 13768 6815
rect 13802 6794 13840 6815
rect 13874 6794 13912 6815
rect 13946 6794 14263 6815
rect 13030 6792 14263 6794
rect 14441 6792 14763 6832
rect 15085 6792 15093 6832
rect 13030 6775 14262 6792
rect 13030 6741 13054 6775
rect 13088 6741 13123 6775
rect 13157 6750 13192 6775
rect 13226 6750 13261 6775
rect 13157 6741 13187 6750
rect 13226 6741 13260 6750
rect 13295 6741 13330 6775
rect 13364 6750 13399 6775
rect 13433 6750 13467 6775
rect 13501 6750 13535 6775
rect 13569 6750 13603 6775
rect 13637 6750 13671 6775
rect 13705 6750 13739 6775
rect 13773 6750 13807 6775
rect 13841 6750 13875 6775
rect 13367 6741 13399 6750
rect 13440 6741 13467 6750
rect 13513 6741 13535 6750
rect 13586 6741 13603 6750
rect 13658 6741 13671 6750
rect 13730 6741 13739 6750
rect 13802 6741 13807 6750
rect 13874 6741 13875 6750
rect 13909 6750 13943 6775
rect 13909 6741 13912 6750
rect 13977 6741 14011 6775
rect 14045 6741 14079 6775
rect 14113 6741 14147 6775
rect 14181 6758 14262 6775
rect 14441 6758 14478 6792
rect 14512 6758 14550 6792
rect 14584 6758 14622 6792
rect 14656 6758 14694 6792
rect 14728 6758 14763 6792
rect 15088 6758 15093 6792
rect 14181 6741 14263 6758
rect 13030 6716 13187 6741
rect 13221 6716 13260 6741
rect 13294 6716 13333 6741
rect 13367 6716 13406 6741
rect 13440 6716 13479 6741
rect 13513 6716 13552 6741
rect 13586 6716 13624 6741
rect 13658 6716 13696 6741
rect 13730 6716 13768 6741
rect 13802 6716 13840 6741
rect 13874 6716 13912 6741
rect 13946 6718 14263 6741
rect 14441 6718 14763 6758
rect 15085 6718 15093 6758
rect 13946 6716 14262 6718
rect 13030 6701 14262 6716
rect 13030 6667 13054 6701
rect 13088 6667 13123 6701
rect 13157 6672 13192 6701
rect 13226 6672 13261 6701
rect 13157 6667 13187 6672
rect 13226 6667 13260 6672
rect 13295 6667 13330 6701
rect 13364 6672 13399 6701
rect 13433 6672 13467 6701
rect 13501 6672 13535 6701
rect 13569 6672 13603 6701
rect 13637 6672 13671 6701
rect 13705 6672 13739 6701
rect 13773 6672 13807 6701
rect 13841 6672 13875 6701
rect 13367 6667 13399 6672
rect 13440 6667 13467 6672
rect 13513 6667 13535 6672
rect 13586 6667 13603 6672
rect 13658 6667 13671 6672
rect 13730 6667 13739 6672
rect 13802 6667 13807 6672
rect 13874 6667 13875 6672
rect 13909 6672 13943 6701
rect 13909 6667 13912 6672
rect 13977 6667 14011 6701
rect 14045 6667 14079 6701
rect 14113 6667 14147 6701
rect 14181 6684 14262 6701
rect 14441 6684 14478 6718
rect 14512 6684 14550 6718
rect 14584 6684 14622 6718
rect 14656 6684 14694 6718
rect 14728 6684 14763 6718
rect 15088 6684 15093 6718
rect 14181 6667 14263 6684
rect 13030 6638 13187 6667
rect 13221 6638 13260 6667
rect 13294 6638 13333 6667
rect 13367 6638 13406 6667
rect 13440 6638 13479 6667
rect 13513 6638 13552 6667
rect 13586 6638 13624 6667
rect 13658 6638 13696 6667
rect 13730 6638 13768 6667
rect 13802 6638 13840 6667
rect 13874 6638 13912 6667
rect 13946 6644 14263 6667
rect 14441 6644 14763 6684
rect 15085 6644 15093 6684
rect 13946 6638 14262 6644
rect 13030 6627 14262 6638
rect 13030 6593 13054 6627
rect 13088 6593 13123 6627
rect 13157 6594 13192 6627
rect 13226 6594 13261 6627
rect 13157 6593 13187 6594
rect 13226 6593 13260 6594
rect 13295 6593 13330 6627
rect 13364 6594 13399 6627
rect 13433 6594 13467 6627
rect 13501 6594 13535 6627
rect 13569 6594 13603 6627
rect 13637 6594 13671 6627
rect 13705 6594 13739 6627
rect 13773 6594 13807 6627
rect 13841 6594 13875 6627
rect 13367 6593 13399 6594
rect 13440 6593 13467 6594
rect 13513 6593 13535 6594
rect 13586 6593 13603 6594
rect 13658 6593 13671 6594
rect 13730 6593 13739 6594
rect 13802 6593 13807 6594
rect 13874 6593 13875 6594
rect 13909 6594 13943 6627
rect 13909 6593 13912 6594
rect 13977 6593 14011 6627
rect 14045 6593 14079 6627
rect 14113 6593 14147 6627
rect 14181 6610 14262 6627
rect 14441 6610 14478 6644
rect 14512 6610 14550 6644
rect 14584 6610 14622 6644
rect 14656 6610 14694 6644
rect 14728 6610 14763 6644
rect 15088 6610 15093 6644
rect 14181 6593 14263 6610
rect 13030 6560 13187 6593
rect 13221 6560 13260 6593
rect 13294 6560 13333 6593
rect 13367 6560 13406 6593
rect 13440 6560 13479 6593
rect 13513 6560 13552 6593
rect 13586 6560 13624 6593
rect 13658 6560 13696 6593
rect 13730 6560 13768 6593
rect 13802 6560 13840 6593
rect 13874 6560 13912 6593
rect 13946 6570 14263 6593
rect 14441 6570 14763 6610
rect 15085 6570 15093 6610
rect 13946 6560 14262 6570
rect 13030 6553 14262 6560
rect 13030 6519 13054 6553
rect 13088 6519 13123 6553
rect 13157 6519 13192 6553
rect 13226 6519 13261 6553
rect 13295 6519 13330 6553
rect 13364 6519 13399 6553
rect 13433 6519 13467 6553
rect 13501 6519 13535 6553
rect 13569 6519 13603 6553
rect 13637 6519 13671 6553
rect 13705 6519 13739 6553
rect 13773 6519 13807 6553
rect 13841 6519 13875 6553
rect 13909 6519 13943 6553
rect 13977 6519 14011 6553
rect 14045 6519 14079 6553
rect 14113 6519 14147 6553
rect 14181 6536 14262 6553
rect 14441 6536 14478 6570
rect 14512 6536 14550 6570
rect 14584 6536 14622 6570
rect 14656 6536 14694 6570
rect 14728 6536 14763 6570
rect 15088 6536 15093 6570
rect 14181 6519 14263 6536
rect 13030 6516 14263 6519
rect 13030 6482 13187 6516
rect 13221 6482 13260 6516
rect 13294 6482 13333 6516
rect 13367 6482 13406 6516
rect 13440 6482 13479 6516
rect 13513 6482 13552 6516
rect 13586 6482 13624 6516
rect 13658 6482 13696 6516
rect 13730 6482 13768 6516
rect 13802 6482 13840 6516
rect 13874 6482 13912 6516
rect 13946 6496 14263 6516
rect 14441 6496 14763 6536
rect 15085 6496 15093 6536
rect 13946 6482 14262 6496
rect 13030 6479 14262 6482
rect 13030 6445 13054 6479
rect 13088 6445 13123 6479
rect 13157 6445 13192 6479
rect 13226 6445 13261 6479
rect 13295 6445 13330 6479
rect 13364 6445 13399 6479
rect 13433 6445 13467 6479
rect 13501 6445 13535 6479
rect 13569 6445 13603 6479
rect 13637 6445 13671 6479
rect 13705 6445 13739 6479
rect 13773 6445 13807 6479
rect 13841 6445 13875 6479
rect 13909 6445 13943 6479
rect 13977 6445 14011 6479
rect 14045 6445 14079 6479
rect 14113 6445 14147 6479
rect 14181 6462 14262 6479
rect 14441 6462 14478 6496
rect 14512 6462 14550 6496
rect 14584 6462 14622 6496
rect 14656 6462 14694 6496
rect 14728 6462 14763 6496
rect 15088 6462 15093 6496
rect 14181 6448 14263 6462
rect 14441 6448 14763 6462
rect 15085 6448 15093 6462
rect 14181 6445 15093 6448
rect 13030 6438 15093 6445
rect 13030 6405 13187 6438
rect 13221 6405 13260 6438
rect 13294 6405 13333 6438
rect 13367 6405 13406 6438
rect 13440 6405 13479 6438
rect 13513 6405 13552 6438
rect 13586 6405 13624 6438
rect 13658 6405 13696 6438
rect 13730 6405 13768 6438
rect 13802 6405 13840 6438
rect 13874 6405 13912 6438
rect 13946 6422 15093 6438
rect 13946 6405 14262 6422
rect 14296 6409 14334 6422
rect 14368 6409 14406 6422
rect 14440 6409 14478 6422
rect 13030 6371 13054 6405
rect 13088 6371 13123 6405
rect 13157 6404 13187 6405
rect 13226 6404 13260 6405
rect 13157 6371 13192 6404
rect 13226 6371 13261 6404
rect 13295 6371 13330 6405
rect 13367 6404 13399 6405
rect 13440 6404 13467 6405
rect 13513 6404 13535 6405
rect 13586 6404 13603 6405
rect 13658 6404 13671 6405
rect 13730 6404 13739 6405
rect 13802 6404 13807 6405
rect 13874 6404 13875 6405
rect 13364 6371 13399 6404
rect 13433 6371 13467 6404
rect 13501 6371 13535 6404
rect 13569 6371 13603 6404
rect 13637 6371 13671 6404
rect 13705 6371 13739 6404
rect 13773 6371 13807 6404
rect 13841 6371 13875 6404
rect 13909 6404 13912 6405
rect 13909 6371 13943 6404
rect 13977 6371 14011 6405
rect 14045 6371 14079 6405
rect 14113 6371 14147 6405
rect 14181 6388 14262 6405
rect 14297 6388 14334 6409
rect 14369 6388 14406 6409
rect 14441 6388 14478 6409
rect 14512 6388 14550 6422
rect 14584 6388 14622 6422
rect 14656 6388 14694 6422
rect 14728 6409 14766 6422
rect 14800 6409 14838 6422
rect 14872 6409 14910 6422
rect 14944 6409 14982 6422
rect 15016 6409 15054 6422
rect 14728 6388 14763 6409
rect 14800 6388 14835 6409
rect 14872 6388 14907 6409
rect 14944 6388 14979 6409
rect 15016 6388 15051 6409
rect 15088 6388 15093 6422
rect 14181 6375 14263 6388
rect 14297 6375 14335 6388
rect 14369 6375 14407 6388
rect 14441 6375 14763 6388
rect 14797 6375 14835 6388
rect 14869 6375 14907 6388
rect 14941 6375 14979 6388
rect 15013 6375 15051 6388
rect 15085 6375 15093 6388
rect 14181 6371 15093 6375
rect 13030 6360 15093 6371
rect 13030 6331 13187 6360
rect 13221 6331 13260 6360
rect 13294 6331 13333 6360
rect 13367 6331 13406 6360
rect 13440 6331 13479 6360
rect 13513 6331 13552 6360
rect 13586 6331 13624 6360
rect 13658 6331 13696 6360
rect 13730 6331 13768 6360
rect 13802 6331 13840 6360
rect 13874 6331 13912 6360
rect 13946 6348 15093 6360
rect 13946 6331 14262 6348
rect 14296 6336 14334 6348
rect 14368 6336 14406 6348
rect 14440 6336 14478 6348
rect 13030 6297 13054 6331
rect 13088 6297 13123 6331
rect 13157 6326 13187 6331
rect 13226 6326 13260 6331
rect 13157 6297 13192 6326
rect 13226 6297 13261 6326
rect 13295 6297 13330 6331
rect 13367 6326 13399 6331
rect 13440 6326 13467 6331
rect 13513 6326 13535 6331
rect 13586 6326 13603 6331
rect 13658 6326 13671 6331
rect 13730 6326 13739 6331
rect 13802 6326 13807 6331
rect 13874 6326 13875 6331
rect 13364 6297 13399 6326
rect 13433 6297 13467 6326
rect 13501 6297 13535 6326
rect 13569 6297 13603 6326
rect 13637 6297 13671 6326
rect 13705 6297 13739 6326
rect 13773 6297 13807 6326
rect 13841 6297 13875 6326
rect 13909 6326 13912 6331
rect 13909 6297 13943 6326
rect 13977 6297 14011 6331
rect 14045 6297 14079 6331
rect 14113 6297 14147 6331
rect 14181 6314 14262 6331
rect 14297 6314 14334 6336
rect 14369 6314 14406 6336
rect 14441 6314 14478 6336
rect 14512 6314 14550 6348
rect 14584 6314 14622 6348
rect 14656 6314 14694 6348
rect 14728 6336 14766 6348
rect 14800 6336 14838 6348
rect 14872 6336 14910 6348
rect 14944 6336 14982 6348
rect 15016 6336 15054 6348
rect 14728 6314 14763 6336
rect 14800 6314 14835 6336
rect 14872 6314 14907 6336
rect 14944 6314 14979 6336
rect 15016 6314 15051 6336
rect 15088 6314 15093 6348
rect 14181 6302 14263 6314
rect 14297 6302 14335 6314
rect 14369 6302 14407 6314
rect 14441 6302 14763 6314
rect 14797 6302 14835 6314
rect 14869 6302 14907 6314
rect 14941 6302 14979 6314
rect 15013 6302 15051 6314
rect 15085 6302 15093 6314
rect 14181 6297 15093 6302
rect 13030 6290 15093 6297
rect 168 6259 846 6286
rect 168 6225 175 6259
rect 209 6247 245 6259
rect 279 6247 315 6259
rect 349 6247 385 6259
rect 419 6247 455 6259
rect 213 6225 245 6247
rect 291 6225 315 6247
rect 369 6225 385 6247
rect 447 6225 455 6247
rect 489 6247 525 6259
rect 489 6225 491 6247
rect 168 6213 179 6225
rect 213 6213 257 6225
rect 291 6213 335 6225
rect 369 6213 413 6225
rect 447 6213 491 6225
rect 559 6247 595 6259
rect 629 6247 665 6259
rect 699 6247 735 6259
rect 769 6247 805 6259
rect 559 6225 569 6247
rect 629 6225 647 6247
rect 699 6225 725 6247
rect 769 6225 803 6247
rect 839 6225 846 6259
rect 525 6213 569 6225
rect 603 6213 647 6225
rect 681 6213 725 6225
rect 759 6213 803 6225
rect 837 6213 846 6225
rect 168 6201 846 6213
rect 168 6166 356 6201
rect 168 6125 173 6166
rect 351 6125 356 6166
rect 168 6091 169 6125
rect 355 6091 356 6125
rect 168 6056 173 6091
rect 351 6056 356 6091
rect 168 6022 169 6056
rect 355 6022 356 6056
rect 168 5987 173 6022
rect 351 5987 356 6022
rect 168 5953 169 5987
rect 355 5953 356 5987
rect 168 5918 173 5953
rect 351 5918 356 5953
rect 168 5884 169 5918
rect 355 5884 356 5918
rect 168 5849 173 5884
rect 351 5849 356 5884
rect 168 5815 169 5849
rect 355 5815 356 5849
rect 168 5780 173 5815
rect 351 5780 356 5815
rect 168 5746 169 5780
rect 355 5746 356 5780
rect 168 5711 173 5746
rect 351 5711 356 5746
rect 168 5677 169 5711
rect 355 5677 356 5711
rect 168 5642 173 5677
rect 351 5642 356 5677
rect 168 5608 169 5642
rect 355 5608 356 5642
rect 168 5573 173 5608
rect 351 5573 356 5608
rect 168 5539 169 5573
rect 355 5539 356 5573
rect 168 5504 173 5539
rect 351 5504 356 5539
rect 168 5470 169 5504
rect 355 5470 356 5504
rect 168 5435 173 5470
rect 351 5435 356 5470
rect 168 5401 169 5435
rect 355 5401 356 5435
rect 168 5366 173 5401
rect 351 5366 356 5401
rect 168 5332 169 5366
rect 355 5332 356 5366
rect 168 5297 173 5332
rect 351 5297 356 5332
rect 168 5263 169 5297
rect 355 5263 356 5297
rect 168 5228 173 5263
rect 351 5228 356 5263
rect 168 5194 169 5228
rect 355 5194 356 5228
rect 168 5159 173 5194
rect 351 5159 356 5194
rect 168 5125 169 5159
rect 355 5125 356 5159
rect 168 5124 173 5125
rect 351 5124 356 5125
rect 168 5090 356 5124
rect 168 5056 169 5090
rect 203 5085 245 5090
rect 279 5085 321 5090
rect 168 5051 173 5056
rect 207 5051 245 5085
rect 279 5051 317 5085
rect 355 5056 356 5090
rect 351 5051 356 5056
rect 168 5021 356 5051
rect 168 4987 169 5021
rect 203 5012 245 5021
rect 279 5012 321 5021
rect 168 4978 173 4987
rect 207 4978 245 5012
rect 279 4978 317 5012
rect 355 4987 356 5021
rect 351 4978 356 4987
rect 168 4952 356 4978
rect 168 4918 169 4952
rect 203 4918 245 4952
rect 279 4918 321 4952
rect 355 4918 408 4952
rect 168 4883 408 4918
rect 168 4849 169 4883
rect 203 4849 245 4883
rect 279 4849 321 4883
rect 355 4849 408 4883
rect 168 4814 408 4849
rect 168 4780 169 4814
rect 203 4780 245 4814
rect 279 4780 321 4814
rect 355 4780 408 4814
rect 168 4745 408 4780
rect 168 4711 169 4745
rect 203 4711 245 4745
rect 279 4711 321 4745
rect 355 4711 408 4745
rect 168 4676 408 4711
rect 168 4642 169 4676
rect 203 4642 245 4676
rect 279 4642 321 4676
rect 355 4642 408 4676
rect 168 4607 408 4642
rect 168 4573 169 4607
rect 203 4573 245 4607
rect 279 4573 321 4607
rect 355 4573 408 4607
rect 168 4538 408 4573
rect 168 4504 169 4538
rect 203 4504 245 4538
rect 279 4504 321 4538
rect 355 4504 408 4538
rect 168 4469 408 4504
rect 168 4435 169 4469
rect 203 4435 245 4469
rect 279 4435 321 4469
rect 355 4435 408 4469
rect 168 4400 408 4435
rect 168 4366 169 4400
rect 203 4366 245 4400
rect 279 4366 321 4400
rect 355 4366 408 4400
rect 168 4331 408 4366
rect 168 4297 169 4331
rect 203 4297 245 4331
rect 279 4297 321 4331
rect 355 4297 408 4331
rect 168 4262 408 4297
rect 168 4228 169 4262
rect 203 4228 245 4262
rect 279 4228 321 4262
rect 355 4228 408 4262
rect 168 4193 408 4228
rect 168 4159 169 4193
rect 203 4159 245 4193
rect 279 4159 321 4193
rect 355 4159 408 4193
rect 168 4146 1048 4159
rect 168 4124 176 4146
rect 210 4124 254 4146
rect 288 4125 1048 4146
rect 288 4124 2120 4125
rect 168 4090 169 4124
rect 210 4112 245 4124
rect 288 4112 321 4124
rect 203 4090 245 4112
rect 279 4090 321 4112
rect 355 4090 2120 4124
rect 168 4081 2120 4090
rect 168 4074 442 4081
rect 168 4055 176 4074
rect 210 4055 254 4074
rect 288 4055 442 4074
rect 168 4021 169 4055
rect 210 4040 245 4055
rect 288 4040 321 4055
rect 203 4021 245 4040
rect 279 4021 321 4040
rect 355 4047 442 4055
rect 476 4047 512 4081
rect 546 4047 582 4081
rect 616 4047 652 4081
rect 686 4047 722 4081
rect 756 4047 792 4081
rect 826 4047 862 4081
rect 896 4047 932 4081
rect 966 4047 1002 4081
rect 1036 4047 1072 4081
rect 1106 4047 1142 4081
rect 1176 4047 1212 4081
rect 1246 4047 1282 4081
rect 1316 4047 1352 4081
rect 1386 4047 1422 4081
rect 1456 4047 1492 4081
rect 1526 4047 1562 4081
rect 1596 4047 1632 4081
rect 1666 4047 1702 4081
rect 1736 4047 1772 4081
rect 1806 4047 1842 4081
rect 1876 4047 1912 4081
rect 1946 4047 1982 4081
rect 2016 4047 2052 4081
rect 2086 4047 2120 4081
rect 355 4021 2120 4047
rect 168 4002 2120 4021
rect 168 3986 176 4002
rect 210 3986 254 4002
rect 288 3986 2120 4002
rect 168 3952 169 3986
rect 210 3968 245 3986
rect 288 3968 321 3986
rect 203 3952 245 3968
rect 279 3952 321 3968
rect 355 3955 2120 3986
rect 355 3952 442 3955
rect 168 3930 442 3952
rect 168 3917 176 3930
rect 210 3917 254 3930
rect 288 3921 442 3930
rect 476 3921 512 3955
rect 546 3921 582 3955
rect 616 3921 652 3955
rect 686 3921 722 3955
rect 756 3921 792 3955
rect 826 3921 862 3955
rect 896 3921 932 3955
rect 966 3921 1002 3955
rect 1036 3921 1072 3955
rect 1106 3921 1142 3955
rect 1176 3921 1212 3955
rect 1246 3921 1282 3955
rect 1316 3921 1352 3955
rect 1386 3921 1422 3955
rect 1456 3921 1492 3955
rect 1526 3921 1562 3955
rect 1596 3921 1632 3955
rect 1666 3921 1702 3955
rect 1736 3921 1772 3955
rect 1806 3921 1842 3955
rect 1876 3921 1912 3955
rect 1946 3921 1982 3955
rect 2016 3921 2052 3955
rect 2086 3921 2120 3955
rect 288 3917 668 3921
rect 168 3883 169 3917
rect 210 3896 245 3917
rect 288 3896 321 3917
rect 203 3883 245 3896
rect 279 3883 321 3896
rect 355 3883 668 3917
rect 168 3858 668 3883
rect 168 3848 176 3858
rect 210 3848 254 3858
rect 288 3848 668 3858
rect 168 3814 169 3848
rect 210 3824 245 3848
rect 288 3824 321 3848
rect 203 3814 245 3824
rect 279 3814 321 3824
rect 355 3845 668 3848
rect 355 3814 410 3845
rect 168 3811 410 3814
rect 444 3811 484 3845
rect 518 3811 558 3845
rect 592 3811 632 3845
rect 666 3811 668 3845
rect 168 3786 668 3811
rect 168 3779 176 3786
rect 210 3779 254 3786
rect 288 3779 668 3786
rect 168 3745 169 3779
rect 210 3752 245 3779
rect 288 3752 321 3779
rect 203 3745 245 3752
rect 279 3745 321 3752
rect 355 3774 668 3779
rect 355 3745 410 3774
rect 168 3740 410 3745
rect 444 3740 484 3774
rect 518 3740 558 3774
rect 592 3740 632 3774
rect 666 3740 668 3774
rect 168 3714 668 3740
rect 168 3710 176 3714
rect 210 3710 254 3714
rect 288 3710 668 3714
rect 168 3676 169 3710
rect 210 3680 245 3710
rect 288 3680 321 3710
rect 203 3676 245 3680
rect 279 3676 321 3680
rect 355 3702 668 3710
rect 355 3676 410 3702
rect 168 3668 410 3676
rect 444 3668 484 3702
rect 518 3668 558 3702
rect 592 3668 632 3702
rect 666 3668 668 3702
rect 168 3642 668 3668
rect 168 3641 176 3642
rect 210 3641 254 3642
rect 288 3641 668 3642
rect 168 3607 169 3641
rect 210 3608 245 3641
rect 288 3608 321 3641
rect 203 3607 245 3608
rect 279 3607 321 3608
rect 355 3630 668 3641
rect 355 3607 410 3630
rect 168 3596 410 3607
rect 444 3596 484 3630
rect 518 3596 558 3630
rect 592 3596 632 3630
rect 666 3596 668 3630
rect 168 3571 668 3596
rect 168 3537 169 3571
rect 203 3570 245 3571
rect 279 3570 321 3571
rect 210 3537 245 3570
rect 288 3537 321 3570
rect 355 3558 668 3571
rect 355 3537 410 3558
rect 168 3536 176 3537
rect 210 3536 254 3537
rect 288 3536 410 3537
rect 168 3524 410 3536
rect 444 3524 484 3558
rect 518 3524 558 3558
rect 592 3524 632 3558
rect 666 3524 668 3558
rect 168 3501 668 3524
rect 168 3467 169 3501
rect 203 3497 245 3501
rect 279 3497 321 3501
rect 210 3467 245 3497
rect 288 3467 321 3497
rect 355 3486 668 3501
rect 355 3467 410 3486
rect 168 3463 176 3467
rect 210 3463 254 3467
rect 288 3463 410 3467
rect 168 3452 410 3463
rect 444 3452 484 3486
rect 518 3452 558 3486
rect 592 3452 632 3486
rect 666 3452 668 3486
rect 168 3431 668 3452
rect 168 3397 169 3431
rect 203 3424 245 3431
rect 279 3424 321 3431
rect 210 3397 245 3424
rect 288 3397 321 3424
rect 355 3414 668 3431
rect 355 3397 410 3414
rect 168 3390 176 3397
rect 210 3390 254 3397
rect 288 3390 410 3397
rect 168 3380 410 3390
rect 444 3380 484 3414
rect 518 3380 558 3414
rect 592 3380 632 3414
rect 666 3380 668 3414
rect 168 3361 668 3380
rect 168 3327 169 3361
rect 203 3351 245 3361
rect 279 3351 321 3361
rect 210 3327 245 3351
rect 288 3327 321 3351
rect 355 3342 668 3361
rect 355 3327 410 3342
rect 168 3317 176 3327
rect 210 3317 254 3327
rect 288 3317 410 3327
rect 168 3308 410 3317
rect 444 3308 484 3342
rect 518 3308 558 3342
rect 592 3308 632 3342
rect 666 3308 668 3342
rect 168 3291 668 3308
rect 168 3257 169 3291
rect 203 3278 245 3291
rect 279 3278 321 3291
rect 210 3257 245 3278
rect 288 3257 321 3278
rect 355 3270 668 3291
rect 355 3257 410 3270
rect 168 3244 176 3257
rect 210 3244 254 3257
rect 288 3244 410 3257
rect 168 3236 410 3244
rect 444 3236 484 3270
rect 518 3236 558 3270
rect 592 3236 632 3270
rect 666 3236 668 3270
rect 168 3221 668 3236
rect 168 3187 169 3221
rect 203 3205 245 3221
rect 279 3205 321 3221
rect 210 3187 245 3205
rect 288 3187 321 3205
rect 355 3198 668 3221
rect 355 3187 410 3198
rect 168 3171 176 3187
rect 210 3171 254 3187
rect 288 3171 410 3187
rect 168 3164 410 3171
rect 444 3164 484 3198
rect 518 3164 558 3198
rect 592 3164 632 3198
rect 666 3164 668 3198
rect 168 3151 668 3164
rect 168 3117 169 3151
rect 203 3132 245 3151
rect 279 3132 321 3151
rect 210 3117 245 3132
rect 288 3117 321 3132
rect 355 3117 668 3151
rect 168 3098 176 3117
rect 210 3098 254 3117
rect 288 3098 668 3117
rect 168 3089 668 3098
rect 1339 3841 2120 3921
rect 1339 3807 1373 3841
rect 1407 3807 1449 3841
rect 1483 3807 1525 3841
rect 1559 3807 1601 3841
rect 1635 3807 1677 3841
rect 1711 3807 1752 3841
rect 1786 3807 1827 3841
rect 1861 3807 1902 3841
rect 1936 3807 1977 3841
rect 2011 3807 2052 3841
rect 2086 3807 2120 3841
rect 1339 3761 2120 3807
rect 1339 3727 1373 3761
rect 1407 3727 1449 3761
rect 1483 3727 1525 3761
rect 1559 3727 1601 3761
rect 1635 3727 1677 3761
rect 1711 3727 1752 3761
rect 1786 3727 1827 3761
rect 1861 3727 1902 3761
rect 1936 3727 1977 3761
rect 2011 3727 2052 3761
rect 2086 3727 2120 3761
rect 1339 3681 2120 3727
rect 1339 3647 1373 3681
rect 1407 3647 1449 3681
rect 1483 3647 1525 3681
rect 1559 3647 1601 3681
rect 1635 3647 1677 3681
rect 1711 3647 1752 3681
rect 1786 3647 1827 3681
rect 1861 3647 1902 3681
rect 1936 3647 1977 3681
rect 2011 3647 2052 3681
rect 2086 3647 2120 3681
rect 1339 3637 2120 3647
rect 1339 3603 1356 3637
rect 1390 3603 1436 3637
rect 1470 3603 1516 3637
rect 1550 3603 1596 3637
rect 1630 3603 1676 3637
rect 1710 3603 1755 3637
rect 1789 3603 1834 3637
rect 1868 3603 1913 3637
rect 1947 3603 1992 3637
rect 2026 3603 2071 3637
rect 2105 3603 2120 3637
rect 1339 3601 2120 3603
rect 1339 3567 1373 3601
rect 1407 3567 1449 3601
rect 1483 3567 1525 3601
rect 1559 3567 1601 3601
rect 1635 3567 1677 3601
rect 1711 3567 1752 3601
rect 1786 3567 1827 3601
rect 1861 3567 1902 3601
rect 1936 3567 1977 3601
rect 2011 3567 2052 3601
rect 2086 3567 2120 3601
rect 1339 3561 2120 3567
rect 1339 3527 1356 3561
rect 1390 3527 1436 3561
rect 1470 3527 1516 3561
rect 1550 3527 1596 3561
rect 1630 3527 1676 3561
rect 1710 3527 1755 3561
rect 1789 3527 1834 3561
rect 1868 3527 1913 3561
rect 1947 3527 1992 3561
rect 2026 3527 2071 3561
rect 2105 3527 2120 3561
rect 1339 3521 2120 3527
rect 1339 3487 1373 3521
rect 1407 3487 1449 3521
rect 1483 3487 1525 3521
rect 1559 3487 1601 3521
rect 1635 3487 1677 3521
rect 1711 3487 1752 3521
rect 1786 3487 1827 3521
rect 1861 3487 1902 3521
rect 1936 3487 1977 3521
rect 2011 3487 2052 3521
rect 2086 3487 2120 3521
rect 1339 3485 2120 3487
rect 1339 3451 1356 3485
rect 1390 3451 1436 3485
rect 1470 3451 1516 3485
rect 1550 3451 1596 3485
rect 1630 3451 1676 3485
rect 1710 3451 1755 3485
rect 1789 3451 1834 3485
rect 1868 3451 1913 3485
rect 1947 3451 1992 3485
rect 2026 3451 2071 3485
rect 2105 3451 2120 3485
rect 1339 3441 2120 3451
rect 1339 3407 1373 3441
rect 1407 3407 1449 3441
rect 1483 3407 1525 3441
rect 1559 3407 1601 3441
rect 1635 3407 1677 3441
rect 1711 3407 1752 3441
rect 1786 3407 1827 3441
rect 1861 3407 1902 3441
rect 1936 3407 1977 3441
rect 2011 3407 2052 3441
rect 2086 3407 2120 3441
rect 1339 3371 2120 3407
rect 1339 3337 1389 3371
rect 1423 3337 1464 3371
rect 1498 3337 1539 3371
rect 1573 3337 1614 3371
rect 1648 3337 1689 3371
rect 1723 3337 1764 3371
rect 1798 3337 1839 3371
rect 1873 3337 1914 3371
rect 1948 3337 1988 3371
rect 2022 3337 2062 3371
rect 2096 3337 2120 3371
rect 1339 3303 2120 3337
rect 1339 3269 1389 3303
rect 1423 3269 1464 3303
rect 1498 3269 1539 3303
rect 1573 3269 1614 3303
rect 1648 3269 1689 3303
rect 1723 3269 1764 3303
rect 1798 3269 1839 3303
rect 1873 3269 1914 3303
rect 1948 3269 1988 3303
rect 2022 3269 2062 3303
rect 2096 3269 2120 3303
rect 1339 3233 2120 3269
rect 1339 3199 1363 3233
rect 1397 3199 1432 3233
rect 1466 3199 1501 3233
rect 1535 3199 1570 3233
rect 1604 3199 1639 3233
rect 1673 3199 1708 3233
rect 1742 3199 1777 3233
rect 1811 3199 1846 3233
rect 1880 3199 1915 3233
rect 1949 3199 1984 3233
rect 2018 3199 2053 3233
rect 2087 3199 2122 3233
rect 2156 3199 2191 3233
rect 2225 3199 2259 3233
rect 2293 3199 2327 3233
rect 2361 3199 2395 3233
rect 2429 3199 2463 3233
rect 2497 3199 2531 3233
rect 2565 3199 2599 3233
rect 2633 3199 2667 3233
rect 2701 3199 2735 3233
rect 2769 3199 2803 3233
rect 2837 3199 2871 3233
rect 2905 3199 2939 3233
rect 2973 3199 3007 3233
rect 3041 3199 3075 3233
rect 3109 3199 3133 3233
rect 1339 3159 3133 3199
rect 1339 3125 1363 3159
rect 1397 3125 1432 3159
rect 1466 3125 1501 3159
rect 1535 3125 1570 3159
rect 1604 3125 1639 3159
rect 1673 3125 1708 3159
rect 1742 3125 1777 3159
rect 1811 3125 1846 3159
rect 1880 3125 1915 3159
rect 1949 3125 1984 3159
rect 2018 3125 2053 3159
rect 2087 3125 2122 3159
rect 2156 3125 2191 3159
rect 2225 3125 2259 3159
rect 2293 3125 2327 3159
rect 2361 3125 2395 3159
rect 2429 3125 2463 3159
rect 2497 3125 2531 3159
rect 2565 3125 2599 3159
rect 2633 3125 2667 3159
rect 2701 3125 2735 3159
rect 2769 3125 2803 3159
rect 2837 3125 2871 3159
rect 2905 3125 2939 3159
rect 2973 3125 3007 3159
rect 3041 3125 3075 3159
rect 3109 3125 3133 3159
rect 1339 3089 3133 3125
rect 168 3087 3133 3089
rect 168 3081 410 3087
rect 168 3047 169 3081
rect 203 3059 245 3081
rect 279 3059 321 3081
rect 210 3047 245 3059
rect 288 3047 321 3059
rect 355 3053 410 3081
rect 444 3053 481 3087
rect 515 3053 552 3087
rect 586 3053 623 3087
rect 657 3053 694 3087
rect 728 3053 765 3087
rect 799 3053 835 3087
rect 869 3053 905 3087
rect 939 3053 975 3087
rect 1009 3053 1045 3087
rect 1079 3053 1115 3087
rect 1149 3053 1185 3087
rect 1219 3053 1255 3087
rect 1289 3085 3133 3087
rect 1289 3053 1363 3085
rect 355 3051 1363 3053
rect 1397 3051 1432 3085
rect 1466 3051 1501 3085
rect 1535 3051 1570 3085
rect 1604 3051 1639 3085
rect 1673 3051 1708 3085
rect 1742 3051 1777 3085
rect 1811 3051 1846 3085
rect 1880 3051 1915 3085
rect 1949 3051 1984 3085
rect 2018 3051 2053 3085
rect 2087 3051 2122 3085
rect 2156 3051 2191 3085
rect 2225 3051 2259 3085
rect 2293 3051 2327 3085
rect 2361 3051 2395 3085
rect 2429 3051 2463 3085
rect 2497 3051 2531 3085
rect 2565 3051 2599 3085
rect 2633 3051 2667 3085
rect 2701 3051 2735 3085
rect 2769 3051 2803 3085
rect 2837 3051 2871 3085
rect 2905 3051 2939 3085
rect 2973 3051 3007 3085
rect 3041 3051 3075 3085
rect 3109 3051 3133 3085
rect 355 3047 3133 3051
rect 168 3025 176 3047
rect 210 3025 254 3047
rect 288 3025 3133 3047
rect 168 3013 3133 3025
rect 168 3011 410 3013
rect 168 2977 169 3011
rect 203 2986 245 3011
rect 279 2986 321 3011
rect 355 3000 410 3011
rect 444 3000 481 3013
rect 515 3000 552 3013
rect 586 3000 623 3013
rect 657 3000 694 3013
rect 728 3000 765 3013
rect 799 3000 835 3013
rect 869 3000 905 3013
rect 939 3000 975 3013
rect 1009 3000 1045 3013
rect 210 2977 245 2986
rect 288 2977 321 2986
rect 375 2979 410 3000
rect 449 2979 481 3000
rect 523 2979 552 3000
rect 597 2979 623 3000
rect 671 2979 694 3000
rect 745 2979 765 3000
rect 819 2979 835 3000
rect 893 2979 905 3000
rect 967 2979 975 3000
rect 1040 2979 1045 3000
rect 1079 2979 1115 3013
rect 1149 2979 1185 3013
rect 1219 2979 1255 3013
rect 1289 3011 3133 3013
rect 1289 2979 1363 3011
rect 168 2952 176 2977
rect 210 2952 254 2977
rect 288 2966 341 2977
rect 375 2966 415 2979
rect 449 2966 489 2979
rect 523 2966 563 2979
rect 597 2966 637 2979
rect 671 2966 711 2979
rect 745 2966 785 2979
rect 819 2966 859 2979
rect 893 2966 933 2979
rect 967 2966 1006 2979
rect 1040 2977 1363 2979
rect 1397 2977 1432 3011
rect 1466 2977 1501 3011
rect 1535 2977 1570 3011
rect 1604 2977 1639 3011
rect 1673 2977 1708 3011
rect 1742 2977 1777 3011
rect 1811 2977 1846 3011
rect 1880 2977 1915 3011
rect 1949 2977 1984 3011
rect 2018 2977 2053 3011
rect 2087 2977 2122 3011
rect 2156 2977 2191 3011
rect 2225 2977 2259 3011
rect 2293 2977 2327 3011
rect 2361 2977 2395 3011
rect 2429 2977 2463 3011
rect 2497 2977 2531 3011
rect 2565 2977 2599 3011
rect 2633 2977 2667 3011
rect 2734 2977 2735 3011
rect 2769 2977 2778 3011
rect 2837 2977 2856 3011
rect 2905 2977 2934 3011
rect 2973 2977 3007 3011
rect 3046 2977 3075 3011
rect 3124 2977 3133 3011
rect 1040 2966 3133 2977
rect 288 2952 3133 2966
rect 168 2941 3133 2952
rect 168 2907 169 2941
rect 203 2907 245 2941
rect 279 2907 321 2941
rect 355 2939 3133 2941
rect 355 2907 410 2939
rect 168 2905 410 2907
rect 444 2905 481 2939
rect 515 2905 552 2939
rect 586 2905 623 2939
rect 657 2905 694 2939
rect 728 2905 765 2939
rect 799 2905 835 2939
rect 869 2905 905 2939
rect 939 2905 975 2939
rect 1009 2905 1045 2939
rect 1079 2905 1115 2939
rect 1149 2905 1185 2939
rect 1219 2905 1255 2939
rect 1289 2937 3133 2939
rect 1289 2905 1363 2937
rect 168 2903 1363 2905
rect 1397 2903 1432 2937
rect 1466 2903 1501 2937
rect 1535 2903 1570 2937
rect 1604 2903 1639 2937
rect 1673 2903 1708 2937
rect 1742 2903 1777 2937
rect 1811 2903 1846 2937
rect 1880 2903 1915 2937
rect 1949 2903 1984 2937
rect 2018 2903 2053 2937
rect 2087 2903 2122 2937
rect 2156 2903 2191 2937
rect 2225 2903 2259 2937
rect 2293 2903 2327 2937
rect 2361 2903 2395 2937
rect 2429 2903 2463 2937
rect 2497 2903 2531 2937
rect 2565 2903 2599 2937
rect 2633 2903 2667 2937
rect 2701 2935 2735 2937
rect 2734 2903 2735 2935
rect 2769 2935 2803 2937
rect 2837 2935 2871 2937
rect 2905 2935 2939 2937
rect 2769 2903 2778 2935
rect 2837 2903 2856 2935
rect 2905 2903 2934 2935
rect 2973 2903 3007 2937
rect 3041 2935 3075 2937
rect 3109 2935 3133 2937
rect 3046 2903 3075 2935
rect 168 2901 2700 2903
rect 2734 2901 2778 2903
rect 2812 2901 2856 2903
rect 2890 2901 2934 2903
rect 2968 2901 3012 2903
rect 3046 2901 3090 2903
rect 3124 2901 3133 2935
rect 168 2871 3133 2901
rect 168 2837 169 2871
rect 203 2837 245 2871
rect 279 2837 321 2871
rect 355 2866 3133 2871
rect 375 2865 415 2866
rect 449 2865 489 2866
rect 523 2865 563 2866
rect 597 2865 637 2866
rect 671 2865 711 2866
rect 745 2865 785 2866
rect 819 2865 859 2866
rect 893 2865 933 2866
rect 967 2865 1006 2866
rect 1040 2865 3133 2866
rect 168 2832 341 2837
rect 375 2832 410 2865
rect 449 2832 481 2865
rect 523 2832 552 2865
rect 597 2832 623 2865
rect 671 2832 694 2865
rect 745 2832 765 2865
rect 819 2832 835 2865
rect 893 2832 905 2865
rect 967 2832 975 2865
rect 1040 2832 1045 2865
rect 168 2831 410 2832
rect 444 2831 481 2832
rect 515 2831 552 2832
rect 586 2831 623 2832
rect 657 2831 694 2832
rect 728 2831 765 2832
rect 799 2831 835 2832
rect 869 2831 905 2832
rect 939 2831 975 2832
rect 1009 2831 1045 2832
rect 1079 2831 1115 2865
rect 1149 2831 1185 2865
rect 1219 2831 1255 2865
rect 1289 2863 3133 2865
rect 1289 2831 1363 2863
rect 168 2829 1363 2831
rect 1397 2829 1432 2863
rect 1466 2829 1501 2863
rect 1535 2829 1570 2863
rect 1604 2829 1639 2863
rect 1673 2829 1708 2863
rect 1742 2829 1777 2863
rect 1811 2829 1846 2863
rect 1880 2829 1915 2863
rect 1949 2829 1984 2863
rect 2018 2829 2053 2863
rect 2087 2829 2122 2863
rect 2156 2829 2191 2863
rect 2225 2829 2259 2863
rect 2293 2829 2327 2863
rect 2361 2829 2395 2863
rect 2429 2829 2463 2863
rect 2497 2829 2531 2863
rect 2565 2829 2599 2863
rect 2633 2829 2667 2863
rect 2701 2859 2735 2863
rect 2734 2829 2735 2859
rect 2769 2859 2803 2863
rect 2837 2859 2871 2863
rect 2905 2859 2939 2863
rect 2769 2829 2778 2859
rect 2837 2829 2856 2859
rect 2905 2829 2934 2859
rect 2973 2829 3007 2863
rect 3041 2859 3075 2863
rect 3109 2859 3133 2863
rect 3046 2829 3075 2859
rect 168 2825 2700 2829
rect 2734 2825 2778 2829
rect 2812 2825 2856 2829
rect 2890 2825 2934 2829
rect 2968 2825 3012 2829
rect 3046 2825 3090 2829
rect 3124 2825 3133 2859
rect 168 2801 3133 2825
rect 168 2767 169 2801
rect 203 2767 245 2801
rect 279 2767 321 2801
rect 355 2791 3133 2801
rect 355 2767 410 2791
rect 168 2757 410 2767
rect 444 2757 481 2791
rect 515 2757 552 2791
rect 586 2757 623 2791
rect 657 2757 694 2791
rect 728 2757 765 2791
rect 799 2757 835 2791
rect 869 2757 905 2791
rect 939 2757 975 2791
rect 1009 2757 1045 2791
rect 1079 2757 1115 2791
rect 1149 2757 1185 2791
rect 1219 2757 1255 2791
rect 1289 2789 3133 2791
rect 1289 2757 1363 2789
rect 168 2755 1363 2757
rect 1397 2755 1432 2789
rect 1466 2755 1501 2789
rect 1535 2755 1570 2789
rect 1604 2755 1639 2789
rect 1673 2755 1708 2789
rect 1742 2755 1777 2789
rect 1811 2755 1846 2789
rect 1880 2755 1915 2789
rect 1949 2755 1984 2789
rect 2018 2755 2053 2789
rect 2087 2755 2122 2789
rect 2156 2755 2191 2789
rect 2225 2755 2259 2789
rect 2293 2755 2327 2789
rect 2361 2755 2395 2789
rect 2429 2755 2463 2789
rect 2497 2755 2531 2789
rect 2565 2755 2599 2789
rect 2633 2755 2667 2789
rect 2701 2783 2735 2789
rect 2734 2755 2735 2783
rect 2769 2783 2803 2789
rect 2837 2783 2871 2789
rect 2905 2783 2939 2789
rect 2769 2755 2778 2783
rect 2837 2755 2856 2783
rect 2905 2755 2934 2783
rect 2973 2755 3007 2789
rect 3041 2783 3075 2789
rect 3109 2783 3133 2789
rect 3046 2755 3075 2783
rect 168 2749 2700 2755
rect 2734 2749 2778 2755
rect 2812 2749 2856 2755
rect 2890 2749 2934 2755
rect 2968 2749 3012 2755
rect 3046 2749 3090 2755
rect 3124 2749 3133 2783
rect 168 2731 3133 2749
rect 168 2697 169 2731
rect 203 2697 245 2731
rect 279 2697 321 2731
rect 355 2717 3133 2731
rect 355 2697 410 2717
rect 168 2683 410 2697
rect 444 2683 481 2717
rect 515 2683 552 2717
rect 586 2683 623 2717
rect 657 2683 694 2717
rect 728 2683 765 2717
rect 799 2683 835 2717
rect 869 2683 905 2717
rect 939 2683 975 2717
rect 1009 2683 1045 2717
rect 1079 2683 1115 2717
rect 1149 2683 1185 2717
rect 1219 2683 1255 2717
rect 1289 2715 3133 2717
rect 1289 2683 1363 2715
rect 168 2681 1363 2683
rect 1397 2681 1432 2715
rect 1466 2681 1501 2715
rect 1535 2681 1570 2715
rect 1604 2681 1639 2715
rect 1673 2681 1708 2715
rect 1742 2681 1777 2715
rect 1811 2681 1846 2715
rect 1880 2681 1915 2715
rect 1949 2686 1984 2715
rect 2018 2686 2053 2715
rect 2087 2686 2122 2715
rect 2156 2686 2191 2715
rect 1949 2681 1958 2686
rect 2018 2681 2034 2686
rect 2087 2681 2110 2686
rect 2156 2681 2186 2686
rect 2225 2681 2259 2715
rect 2293 2686 2327 2715
rect 2361 2686 2395 2715
rect 2429 2686 2463 2715
rect 2497 2686 2531 2715
rect 2296 2681 2327 2686
rect 2372 2681 2395 2686
rect 2448 2681 2463 2686
rect 2524 2681 2531 2686
rect 2565 2686 2599 2715
rect 168 2661 1958 2681
rect 168 2627 169 2661
rect 203 2627 245 2661
rect 279 2627 321 2661
rect 355 2652 1958 2661
rect 1992 2652 2034 2681
rect 2068 2652 2110 2681
rect 2144 2652 2186 2681
rect 2220 2652 2262 2681
rect 2296 2652 2338 2681
rect 2372 2652 2414 2681
rect 2448 2652 2490 2681
rect 2524 2652 2565 2681
rect 2633 2686 2667 2715
rect 2701 2686 2735 2715
rect 2769 2686 2803 2715
rect 2837 2686 2871 2715
rect 2633 2681 2640 2686
rect 2701 2681 2715 2686
rect 2769 2681 2790 2686
rect 2837 2681 2865 2686
rect 2905 2681 2939 2715
rect 2973 2686 3007 2715
rect 3041 2686 3075 2715
rect 3109 2686 3133 2715
rect 2974 2681 3007 2686
rect 3049 2681 3075 2686
rect 2599 2652 2640 2681
rect 2674 2652 2715 2681
rect 2749 2652 2790 2681
rect 2824 2652 2865 2681
rect 2899 2652 2940 2681
rect 2974 2652 3015 2681
rect 3049 2652 3090 2681
rect 3124 2652 3133 2686
rect 355 2643 3133 2652
rect 355 2627 410 2643
rect 168 2609 410 2627
rect 444 2609 481 2643
rect 515 2609 552 2643
rect 586 2609 623 2643
rect 657 2609 694 2643
rect 728 2609 765 2643
rect 799 2609 835 2643
rect 869 2609 905 2643
rect 939 2609 975 2643
rect 1009 2609 1045 2643
rect 1079 2609 1115 2643
rect 1149 2609 1185 2643
rect 1219 2609 1255 2643
rect 1289 2641 3133 2643
rect 1289 2609 1363 2641
rect 168 2607 1363 2609
rect 1397 2607 1432 2641
rect 1466 2607 1501 2641
rect 1535 2607 1570 2641
rect 1604 2607 1639 2641
rect 1673 2607 1708 2641
rect 1742 2607 1777 2641
rect 1811 2607 1846 2641
rect 1880 2607 1915 2641
rect 1949 2607 1984 2641
rect 2018 2607 2053 2641
rect 2087 2607 2122 2641
rect 2156 2607 2191 2641
rect 2225 2607 2259 2641
rect 2293 2607 2327 2641
rect 2361 2607 2395 2641
rect 2429 2607 2463 2641
rect 2497 2607 2531 2641
rect 2565 2607 2599 2641
rect 2633 2607 2667 2641
rect 2701 2607 2735 2641
rect 2769 2607 2803 2641
rect 2837 2607 2871 2641
rect 2905 2607 2939 2641
rect 2973 2607 3007 2641
rect 3041 2607 3075 2641
rect 3109 2607 3133 2641
rect 168 2591 3133 2607
rect 168 2557 169 2591
rect 203 2557 245 2591
rect 279 2557 321 2591
rect 355 2576 3133 2591
rect 355 2569 1958 2576
rect 355 2557 410 2569
rect 168 2535 410 2557
rect 444 2535 481 2569
rect 515 2535 552 2569
rect 586 2535 623 2569
rect 657 2535 694 2569
rect 728 2535 765 2569
rect 799 2535 835 2569
rect 869 2535 905 2569
rect 939 2535 975 2569
rect 1009 2535 1045 2569
rect 1079 2535 1115 2569
rect 1149 2535 1185 2569
rect 1219 2535 1255 2569
rect 1289 2567 1958 2569
rect 1992 2567 2034 2576
rect 2068 2567 2110 2576
rect 2144 2567 2186 2576
rect 2220 2567 2262 2576
rect 2296 2567 2338 2576
rect 2372 2567 2414 2576
rect 2448 2567 2490 2576
rect 2524 2567 2565 2576
rect 1289 2535 1363 2567
rect 168 2533 1363 2535
rect 1397 2533 1432 2567
rect 1466 2533 1501 2567
rect 1535 2533 1570 2567
rect 1604 2533 1639 2567
rect 1673 2533 1708 2567
rect 1742 2533 1777 2567
rect 1811 2533 1846 2567
rect 1880 2533 1915 2567
rect 1949 2542 1958 2567
rect 2018 2542 2034 2567
rect 2087 2542 2110 2567
rect 2156 2542 2186 2567
rect 1949 2533 1984 2542
rect 2018 2533 2053 2542
rect 2087 2533 2122 2542
rect 2156 2533 2191 2542
rect 2225 2533 2259 2567
rect 2296 2542 2327 2567
rect 2372 2542 2395 2567
rect 2448 2542 2463 2567
rect 2524 2542 2531 2567
rect 2293 2533 2327 2542
rect 2361 2533 2395 2542
rect 2429 2533 2463 2542
rect 2497 2533 2531 2542
rect 2599 2567 2640 2576
rect 2674 2567 2715 2576
rect 2749 2567 2790 2576
rect 2824 2567 2865 2576
rect 2899 2567 2940 2576
rect 2974 2567 3015 2576
rect 3049 2567 3090 2576
rect 2565 2533 2599 2542
rect 2633 2542 2640 2567
rect 2701 2542 2715 2567
rect 2769 2542 2790 2567
rect 2837 2542 2865 2567
rect 2633 2533 2667 2542
rect 2701 2533 2735 2542
rect 2769 2533 2803 2542
rect 2837 2533 2871 2542
rect 2905 2533 2939 2567
rect 2974 2542 3007 2567
rect 3049 2542 3075 2567
rect 3124 2542 3133 2576
rect 2973 2533 3007 2542
rect 3041 2533 3075 2542
rect 3109 2533 3133 2542
rect 25812 2033 27880 2034
rect 25812 1999 25846 2033
rect 25880 2019 25917 2033
rect 25951 2019 25988 2033
rect 26022 2019 26059 2033
rect 26093 2019 26130 2033
rect 26164 2019 26201 2033
rect 26235 2019 26272 2033
rect 26306 2019 26342 2033
rect 26376 2019 26412 2033
rect 26446 2019 26482 2033
rect 26516 2019 26552 2033
rect 26586 2019 26622 2033
rect 25889 1999 25917 2019
rect 25962 1999 25988 2019
rect 26035 1999 26059 2019
rect 26108 1999 26130 2019
rect 26181 1999 26201 2019
rect 26254 1999 26272 2019
rect 26327 1999 26342 2019
rect 26400 1999 26412 2019
rect 26473 1999 26482 2019
rect 26546 1999 26552 2019
rect 26619 1999 26622 2019
rect 26656 2019 26692 2033
rect 26656 1999 26658 2019
rect 25812 1985 25855 1999
rect 25889 1985 25928 1999
rect 25962 1985 26001 1999
rect 26035 1985 26074 1999
rect 26108 1985 26147 1999
rect 26181 1985 26220 1999
rect 26254 1985 26293 1999
rect 26327 1985 26366 1999
rect 26400 1985 26439 1999
rect 26473 1985 26512 1999
rect 26546 1985 26585 1999
rect 26619 1985 26658 1999
rect 26726 2019 26762 2033
rect 26796 2019 26832 2033
rect 26866 2019 26902 2033
rect 26936 2019 26972 2033
rect 27006 2019 27042 2033
rect 27076 2019 27112 2033
rect 27146 2019 27182 2033
rect 27216 2019 27252 2033
rect 27286 2019 27322 2033
rect 27356 2019 27392 2033
rect 27426 2019 27462 2033
rect 27496 2019 27532 2033
rect 27566 2019 27602 2033
rect 27636 2019 27672 2033
rect 26726 1999 26731 2019
rect 26796 1999 26804 2019
rect 26866 1999 26877 2019
rect 26936 1999 26950 2019
rect 27006 1999 27022 2019
rect 27076 1999 27094 2019
rect 27146 1999 27166 2019
rect 27216 1999 27238 2019
rect 27286 1999 27310 2019
rect 27356 1999 27382 2019
rect 27426 1999 27454 2019
rect 27496 1999 27526 2019
rect 27566 1999 27598 2019
rect 27636 1999 27670 2019
rect 27706 1999 27742 2033
rect 27776 1999 27812 2033
rect 27846 2019 27880 2033
rect 26692 1985 26731 1999
rect 26765 1985 26804 1999
rect 26838 1985 26877 1999
rect 26911 1985 26950 1999
rect 26984 1985 27022 1999
rect 27056 1985 27094 1999
rect 27128 1985 27166 1999
rect 27200 1985 27238 1999
rect 27272 1985 27310 1999
rect 27344 1985 27382 1999
rect 27416 1985 27454 1999
rect 27488 1985 27526 1999
rect 27560 1985 27598 1999
rect 27632 1985 27670 1999
rect 27704 1985 27742 1999
rect 27776 1985 27814 1999
rect 27848 1985 27880 2019
rect 25812 1947 27880 1985
rect 25812 1913 25846 1947
rect 25880 1939 25917 1947
rect 25951 1939 25988 1947
rect 26022 1939 26059 1947
rect 26093 1939 26130 1947
rect 26164 1939 26201 1947
rect 26235 1939 26272 1947
rect 26306 1939 26342 1947
rect 26376 1939 26412 1947
rect 26446 1939 26482 1947
rect 26516 1939 26552 1947
rect 26586 1939 26622 1947
rect 25889 1913 25917 1939
rect 25962 1913 25988 1939
rect 26035 1913 26059 1939
rect 26108 1913 26130 1939
rect 26181 1913 26201 1939
rect 26254 1913 26272 1939
rect 26327 1913 26342 1939
rect 26400 1913 26412 1939
rect 26473 1913 26482 1939
rect 26546 1913 26552 1939
rect 26619 1913 26622 1939
rect 26656 1939 26692 1947
rect 26656 1913 26658 1939
rect 25812 1905 25855 1913
rect 25889 1905 25928 1913
rect 25962 1905 26001 1913
rect 26035 1905 26074 1913
rect 26108 1905 26147 1913
rect 26181 1905 26220 1913
rect 26254 1905 26293 1913
rect 26327 1905 26366 1913
rect 26400 1905 26439 1913
rect 26473 1905 26512 1913
rect 26546 1905 26585 1913
rect 26619 1905 26658 1913
rect 26726 1939 26762 1947
rect 26796 1939 26832 1947
rect 26866 1939 26902 1947
rect 26936 1939 26972 1947
rect 27006 1939 27042 1947
rect 27076 1939 27112 1947
rect 27146 1939 27182 1947
rect 27216 1939 27252 1947
rect 27286 1939 27322 1947
rect 27356 1939 27392 1947
rect 27426 1939 27462 1947
rect 27496 1939 27532 1947
rect 27566 1939 27602 1947
rect 27636 1939 27672 1947
rect 26726 1913 26731 1939
rect 26796 1913 26804 1939
rect 26866 1913 26877 1939
rect 26936 1913 26950 1939
rect 27006 1913 27022 1939
rect 27076 1913 27094 1939
rect 27146 1913 27166 1939
rect 27216 1913 27238 1939
rect 27286 1913 27310 1939
rect 27356 1913 27382 1939
rect 27426 1913 27454 1939
rect 27496 1913 27526 1939
rect 27566 1913 27598 1939
rect 27636 1913 27670 1939
rect 27706 1913 27742 1947
rect 27776 1913 27812 1947
rect 27846 1939 27880 1947
rect 26692 1905 26731 1913
rect 26765 1905 26804 1913
rect 26838 1905 26877 1913
rect 26911 1905 26950 1913
rect 26984 1905 27022 1913
rect 27056 1905 27094 1913
rect 27128 1905 27166 1913
rect 27200 1905 27238 1913
rect 27272 1905 27310 1913
rect 27344 1905 27382 1913
rect 27416 1905 27454 1913
rect 27488 1905 27526 1913
rect 27560 1905 27598 1913
rect 27632 1905 27670 1913
rect 27704 1905 27742 1913
rect 27776 1905 27814 1913
rect 27848 1905 27880 1939
rect 25812 1861 27880 1905
rect 25812 1827 25846 1861
rect 25880 1859 25917 1861
rect 25951 1859 25988 1861
rect 26022 1859 26059 1861
rect 26093 1859 26130 1861
rect 26164 1859 26201 1861
rect 26235 1859 26272 1861
rect 26306 1859 26342 1861
rect 26376 1859 26412 1861
rect 26446 1859 26482 1861
rect 26516 1859 26552 1861
rect 26586 1859 26622 1861
rect 25889 1827 25917 1859
rect 25962 1827 25988 1859
rect 26035 1827 26059 1859
rect 26108 1827 26130 1859
rect 26181 1827 26201 1859
rect 26254 1827 26272 1859
rect 26327 1827 26342 1859
rect 26400 1827 26412 1859
rect 26473 1827 26482 1859
rect 26546 1827 26552 1859
rect 26619 1827 26622 1859
rect 26656 1859 26692 1861
rect 26656 1827 26658 1859
rect 25812 1825 25855 1827
rect 25889 1825 25928 1827
rect 25962 1825 26001 1827
rect 26035 1825 26074 1827
rect 26108 1825 26147 1827
rect 26181 1825 26220 1827
rect 26254 1825 26293 1827
rect 26327 1825 26366 1827
rect 26400 1825 26439 1827
rect 26473 1825 26512 1827
rect 26546 1825 26585 1827
rect 26619 1825 26658 1827
rect 26726 1859 26762 1861
rect 26796 1859 26832 1861
rect 26866 1859 26902 1861
rect 26936 1859 26972 1861
rect 27006 1859 27042 1861
rect 27076 1859 27112 1861
rect 27146 1859 27182 1861
rect 27216 1859 27252 1861
rect 27286 1859 27322 1861
rect 27356 1859 27392 1861
rect 27426 1859 27462 1861
rect 27496 1859 27532 1861
rect 27566 1859 27602 1861
rect 27636 1859 27672 1861
rect 26726 1827 26731 1859
rect 26796 1827 26804 1859
rect 26866 1827 26877 1859
rect 26936 1827 26950 1859
rect 27006 1827 27022 1859
rect 27076 1827 27094 1859
rect 27146 1827 27166 1859
rect 27216 1827 27238 1859
rect 27286 1827 27310 1859
rect 27356 1827 27382 1859
rect 27426 1827 27454 1859
rect 27496 1827 27526 1859
rect 27566 1827 27598 1859
rect 27636 1827 27670 1859
rect 27706 1827 27742 1861
rect 27776 1827 27812 1861
rect 27846 1859 27880 1861
rect 26692 1825 26731 1827
rect 26765 1825 26804 1827
rect 26838 1825 26877 1827
rect 26911 1825 26950 1827
rect 26984 1825 27022 1827
rect 27056 1825 27094 1827
rect 27128 1825 27166 1827
rect 27200 1825 27238 1827
rect 27272 1825 27310 1827
rect 27344 1825 27382 1827
rect 27416 1825 27454 1827
rect 27488 1825 27526 1827
rect 27560 1825 27598 1827
rect 27632 1825 27670 1827
rect 27704 1825 27742 1827
rect 27776 1825 27814 1827
rect 27848 1825 27880 1859
rect 25812 1779 27880 1825
rect 25812 1775 25855 1779
rect 25889 1775 25928 1779
rect 25962 1775 26001 1779
rect 26035 1775 26074 1779
rect 26108 1775 26147 1779
rect 26181 1775 26220 1779
rect 26254 1775 26293 1779
rect 26327 1775 26366 1779
rect 26400 1775 26439 1779
rect 26473 1775 26512 1779
rect 26546 1775 26585 1779
rect 26619 1775 26658 1779
rect 25812 1741 25846 1775
rect 25889 1745 25917 1775
rect 25962 1745 25988 1775
rect 26035 1745 26059 1775
rect 26108 1745 26130 1775
rect 26181 1745 26201 1775
rect 26254 1745 26272 1775
rect 26327 1745 26342 1775
rect 26400 1745 26412 1775
rect 26473 1745 26482 1775
rect 26546 1745 26552 1775
rect 26619 1745 26622 1775
rect 25880 1741 25917 1745
rect 25951 1741 25988 1745
rect 26022 1741 26059 1745
rect 26093 1741 26130 1745
rect 26164 1741 26201 1745
rect 26235 1741 26272 1745
rect 26306 1741 26342 1745
rect 26376 1741 26412 1745
rect 26446 1741 26482 1745
rect 26516 1741 26552 1745
rect 26586 1741 26622 1745
rect 26656 1745 26658 1775
rect 26692 1775 26731 1779
rect 26765 1775 26804 1779
rect 26838 1775 26877 1779
rect 26911 1775 26950 1779
rect 26984 1775 27022 1779
rect 27056 1775 27094 1779
rect 27128 1775 27166 1779
rect 27200 1775 27238 1779
rect 27272 1775 27310 1779
rect 27344 1775 27382 1779
rect 27416 1775 27454 1779
rect 27488 1775 27526 1779
rect 27560 1775 27598 1779
rect 27632 1775 27670 1779
rect 27704 1775 27742 1779
rect 27776 1775 27814 1779
rect 26656 1741 26692 1745
rect 26726 1745 26731 1775
rect 26796 1745 26804 1775
rect 26866 1745 26877 1775
rect 26936 1745 26950 1775
rect 27006 1745 27022 1775
rect 27076 1745 27094 1775
rect 27146 1745 27166 1775
rect 27216 1745 27238 1775
rect 27286 1745 27310 1775
rect 27356 1745 27382 1775
rect 27426 1745 27454 1775
rect 27496 1745 27526 1775
rect 27566 1745 27598 1775
rect 27636 1745 27670 1775
rect 26726 1741 26762 1745
rect 26796 1741 26832 1745
rect 26866 1741 26902 1745
rect 26936 1741 26972 1745
rect 27006 1741 27042 1745
rect 27076 1741 27112 1745
rect 27146 1741 27182 1745
rect 27216 1741 27252 1745
rect 27286 1741 27322 1745
rect 27356 1741 27392 1745
rect 27426 1741 27462 1745
rect 27496 1741 27532 1745
rect 27566 1741 27602 1745
rect 27636 1741 27672 1745
rect 27706 1741 27742 1775
rect 27776 1741 27812 1775
rect 27848 1745 27880 1779
rect 27846 1741 27880 1745
rect 25812 1740 27880 1741
rect 25823 1739 27880 1740
<< viali >>
rect 92 39900 126 39912
rect 92 39878 110 39900
rect 110 39878 126 39900
rect 174 39900 208 39912
rect 174 39878 198 39900
rect 198 39878 208 39900
rect 92 39831 126 39840
rect 92 39806 110 39831
rect 110 39806 126 39831
rect 174 39831 208 39840
rect 174 39806 198 39831
rect 198 39806 208 39831
rect 92 39762 126 39768
rect 92 39734 110 39762
rect 110 39734 126 39762
rect 174 39762 208 39768
rect 174 39734 198 39762
rect 198 39734 208 39762
rect 92 39693 126 39696
rect 92 39662 110 39693
rect 110 39662 126 39693
rect 174 39693 208 39696
rect 174 39662 198 39693
rect 198 39662 208 39693
rect 92 39590 110 39624
rect 110 39590 126 39624
rect 174 39590 198 39624
rect 198 39590 208 39624
rect 92 39521 110 39552
rect 110 39521 126 39552
rect 92 39518 126 39521
rect 174 39521 198 39552
rect 198 39521 208 39552
rect 174 39518 208 39521
rect 92 39452 110 39480
rect 110 39452 126 39480
rect 92 39446 126 39452
rect 174 39452 198 39480
rect 198 39452 208 39480
rect 174 39446 208 39452
rect 92 39383 110 39408
rect 110 39383 126 39408
rect 92 39374 126 39383
rect 174 39383 198 39408
rect 198 39383 208 39408
rect 174 39374 208 39383
rect 92 39314 110 39336
rect 110 39314 126 39336
rect 92 39302 126 39314
rect 174 39314 198 39336
rect 198 39314 208 39336
rect 174 39302 208 39314
rect 92 39245 110 39264
rect 110 39245 126 39264
rect 92 39230 126 39245
rect 174 39245 198 39264
rect 198 39245 208 39264
rect 174 39230 208 39245
rect 92 39175 110 39192
rect 110 39175 126 39192
rect 92 39158 126 39175
rect 174 39175 198 39192
rect 198 39175 208 39192
rect 174 39158 208 39175
rect 92 39105 110 39120
rect 110 39105 126 39120
rect 92 39086 126 39105
rect 174 39105 198 39120
rect 198 39105 208 39120
rect 174 39086 208 39105
rect 92 39035 110 39048
rect 110 39035 126 39048
rect 92 39014 126 39035
rect 174 39035 198 39048
rect 198 39035 208 39048
rect 174 39014 208 39035
rect 92 38965 110 38976
rect 110 38965 126 38976
rect 92 38942 126 38965
rect 174 38965 198 38976
rect 198 38965 208 38976
rect 174 38942 208 38965
rect 92 38895 110 38904
rect 110 38895 126 38904
rect 92 38870 126 38895
rect 174 38895 198 38904
rect 198 38895 208 38904
rect 174 38870 208 38895
rect 92 38825 110 38832
rect 110 38825 126 38832
rect 92 38798 126 38825
rect 174 38825 198 38832
rect 198 38825 208 38832
rect 174 38798 208 38825
rect 92 38755 110 38760
rect 110 38755 126 38760
rect 92 38726 126 38755
rect 174 38755 198 38760
rect 198 38755 208 38760
rect 174 38726 208 38755
rect 92 38685 110 38688
rect 110 38685 126 38688
rect 92 38654 126 38685
rect 174 38685 198 38688
rect 198 38685 208 38688
rect 174 38654 208 38685
rect 92 38615 110 38616
rect 110 38615 126 38616
rect 92 38582 126 38615
rect 174 38615 198 38616
rect 198 38615 208 38616
rect 174 38582 208 38615
rect 92 38510 126 38544
rect 174 38510 208 38544
rect 92 38439 126 38472
rect 92 38438 110 38439
rect 110 38438 126 38439
rect 174 38439 208 38472
rect 174 38438 198 38439
rect 198 38438 208 38439
rect 92 38369 126 38400
rect 92 38366 110 38369
rect 110 38366 126 38369
rect 174 38369 208 38400
rect 174 38366 198 38369
rect 198 38366 208 38369
rect 92 38299 126 38328
rect 92 38294 110 38299
rect 110 38294 126 38299
rect 174 38299 208 38328
rect 174 38294 198 38299
rect 198 38294 208 38299
rect 92 38229 126 38256
rect 92 38222 110 38229
rect 110 38222 126 38229
rect 174 38229 208 38256
rect 174 38222 198 38229
rect 198 38222 208 38229
rect 92 38159 126 38184
rect 92 38150 110 38159
rect 110 38150 126 38159
rect 174 38159 208 38184
rect 174 38150 198 38159
rect 198 38150 208 38159
rect 92 38089 126 38111
rect 92 38077 110 38089
rect 110 38077 126 38089
rect 174 38089 208 38111
rect 174 38077 198 38089
rect 198 38077 208 38089
rect 92 38004 126 38038
rect 174 38004 208 38038
rect 209 37770 243 37804
rect 291 37770 325 37804
rect 209 37698 243 37732
rect 291 37698 325 37732
rect 209 37626 243 37660
rect 291 37626 325 37660
rect 209 37554 243 37588
rect 291 37554 325 37588
rect 209 37484 243 37516
rect 291 37484 325 37516
rect 209 37482 219 37484
rect 219 37482 243 37484
rect 291 37482 305 37484
rect 305 37482 325 37484
rect 209 37415 243 37444
rect 291 37415 325 37444
rect 209 37410 219 37415
rect 219 37410 243 37415
rect 291 37410 305 37415
rect 305 37410 325 37415
rect 209 37346 243 37372
rect 291 37346 325 37372
rect 209 37338 219 37346
rect 219 37338 243 37346
rect 291 37338 305 37346
rect 305 37338 325 37346
rect 209 37277 243 37300
rect 291 37277 325 37300
rect 209 37266 219 37277
rect 219 37266 243 37277
rect 291 37266 305 37277
rect 305 37266 325 37277
rect 209 37208 243 37228
rect 291 37208 325 37228
rect 209 37194 219 37208
rect 219 37194 243 37208
rect 291 37194 305 37208
rect 305 37194 325 37208
rect 209 37139 243 37156
rect 291 37139 325 37156
rect 209 37122 219 37139
rect 219 37122 243 37139
rect 291 37122 305 37139
rect 305 37122 325 37139
rect 209 37070 243 37084
rect 291 37070 325 37084
rect 209 37050 219 37070
rect 219 37050 243 37070
rect 291 37050 305 37070
rect 305 37050 325 37070
rect 209 37001 243 37012
rect 291 37001 325 37012
rect 209 36978 219 37001
rect 219 36978 243 37001
rect 291 36978 305 37001
rect 305 36978 325 37001
rect 209 36932 243 36940
rect 291 36932 325 36940
rect 209 36906 219 36932
rect 219 36906 243 36932
rect 291 36906 305 36932
rect 305 36906 325 36932
rect 209 36863 243 36868
rect 291 36863 325 36868
rect 209 36834 219 36863
rect 219 36834 243 36863
rect 291 36834 305 36863
rect 305 36834 325 36863
rect 209 36794 243 36796
rect 291 36794 325 36796
rect 209 36762 219 36794
rect 219 36762 243 36794
rect 291 36762 305 36794
rect 305 36762 325 36794
rect 209 36691 219 36724
rect 219 36691 243 36724
rect 291 36691 305 36724
rect 305 36691 325 36724
rect 209 36690 243 36691
rect 291 36690 325 36691
rect 209 36621 219 36652
rect 219 36621 243 36652
rect 291 36621 305 36652
rect 305 36621 325 36652
rect 209 36618 243 36621
rect 291 36618 325 36621
rect 209 36551 219 36580
rect 219 36551 243 36580
rect 291 36551 305 36580
rect 305 36551 325 36580
rect 209 36546 243 36551
rect 291 36546 325 36551
rect 209 36481 219 36508
rect 219 36481 243 36508
rect 291 36481 305 36508
rect 305 36481 325 36508
rect 209 36474 243 36481
rect 291 36474 325 36481
rect 209 36411 219 36436
rect 219 36411 243 36436
rect 291 36411 305 36436
rect 305 36411 325 36436
rect 209 36402 243 36411
rect 291 36402 325 36411
rect 209 36341 219 36364
rect 219 36341 243 36364
rect 291 36341 305 36364
rect 305 36341 325 36364
rect 209 36330 243 36341
rect 291 36330 325 36341
rect 209 36271 219 36292
rect 219 36271 243 36292
rect 291 36271 305 36292
rect 305 36271 325 36292
rect 209 36258 243 36271
rect 291 36258 325 36271
rect 209 36201 219 36220
rect 219 36201 243 36220
rect 291 36201 305 36220
rect 305 36201 325 36220
rect 209 36186 243 36201
rect 291 36186 325 36201
rect 209 36131 219 36148
rect 219 36131 243 36148
rect 291 36131 305 36148
rect 305 36131 325 36148
rect 209 36114 243 36131
rect 291 36114 325 36131
rect 209 36061 219 36076
rect 219 36061 243 36076
rect 291 36061 305 36076
rect 305 36061 325 36076
rect 209 36042 243 36061
rect 291 36042 325 36061
rect 209 35991 219 36004
rect 219 35991 243 36004
rect 291 35991 305 36004
rect 305 35991 325 36004
rect 209 35970 243 35991
rect 291 35970 325 35991
rect 209 35898 243 35932
rect 291 35898 325 35932
rect 209 35826 243 35860
rect 291 35857 312 35860
rect 312 35857 325 35860
rect 291 35826 325 35857
rect 209 35754 243 35788
rect 291 35755 325 35788
rect 291 35754 312 35755
rect 312 35754 325 35755
rect 209 35682 243 35716
rect 291 35687 325 35716
rect 291 35682 312 35687
rect 312 35682 325 35687
rect 22829 36361 22863 36384
rect 22911 36361 22945 36384
rect 22993 36361 23027 36384
rect 23075 36361 23109 36384
rect 23157 36361 23191 36384
rect 23239 36361 23273 36384
rect 22829 36350 22861 36361
rect 22861 36350 22863 36361
rect 22911 36350 22931 36361
rect 22931 36350 22945 36361
rect 22993 36350 23001 36361
rect 23001 36350 23027 36361
rect 23075 36350 23107 36361
rect 23107 36350 23109 36361
rect 23157 36350 23177 36361
rect 23177 36350 23191 36361
rect 23239 36350 23247 36361
rect 23247 36350 23273 36361
rect 22829 36293 22863 36312
rect 22911 36293 22945 36312
rect 22993 36293 23027 36312
rect 23075 36293 23109 36312
rect 23157 36293 23191 36312
rect 23239 36293 23273 36312
rect 22829 36278 22861 36293
rect 22861 36278 22863 36293
rect 22911 36278 22931 36293
rect 22931 36278 22945 36293
rect 22993 36278 23001 36293
rect 23001 36278 23027 36293
rect 23075 36278 23107 36293
rect 23107 36278 23109 36293
rect 23157 36278 23177 36293
rect 23177 36278 23191 36293
rect 23239 36278 23247 36293
rect 23247 36278 23273 36293
rect 22829 36225 22863 36240
rect 22911 36225 22945 36240
rect 22993 36225 23027 36240
rect 23075 36225 23109 36240
rect 23157 36225 23191 36240
rect 23239 36225 23273 36240
rect 22829 36206 22861 36225
rect 22861 36206 22863 36225
rect 22911 36206 22931 36225
rect 22931 36206 22945 36225
rect 22993 36206 23001 36225
rect 23001 36206 23027 36225
rect 23075 36206 23107 36225
rect 23107 36206 23109 36225
rect 23157 36206 23177 36225
rect 23177 36206 23191 36225
rect 23239 36206 23247 36225
rect 23247 36206 23273 36225
rect 22829 36157 22863 36168
rect 22911 36157 22945 36168
rect 22993 36157 23027 36168
rect 23075 36157 23109 36168
rect 23157 36157 23191 36168
rect 23239 36157 23273 36168
rect 22829 36134 22861 36157
rect 22861 36134 22863 36157
rect 22911 36134 22931 36157
rect 22931 36134 22945 36157
rect 22993 36134 23001 36157
rect 23001 36134 23027 36157
rect 23075 36134 23107 36157
rect 23107 36134 23109 36157
rect 23157 36134 23177 36157
rect 23177 36134 23191 36157
rect 23239 36134 23247 36157
rect 23247 36134 23273 36157
rect 22829 36089 22863 36096
rect 22911 36089 22945 36096
rect 22993 36089 23027 36096
rect 23075 36089 23109 36096
rect 23157 36089 23191 36096
rect 23239 36089 23273 36096
rect 22829 36062 22861 36089
rect 22861 36062 22863 36089
rect 22911 36062 22931 36089
rect 22931 36062 22945 36089
rect 22993 36062 23001 36089
rect 23001 36062 23027 36089
rect 23075 36062 23107 36089
rect 23107 36062 23109 36089
rect 23157 36062 23177 36089
rect 23177 36062 23191 36089
rect 23239 36062 23247 36089
rect 23247 36062 23273 36089
rect 22829 36021 22863 36024
rect 22911 36021 22945 36024
rect 22993 36021 23027 36024
rect 23075 36021 23109 36024
rect 23157 36021 23191 36024
rect 23239 36021 23273 36024
rect 22829 35990 22861 36021
rect 22861 35990 22863 36021
rect 22911 35990 22931 36021
rect 22931 35990 22945 36021
rect 22993 35990 23001 36021
rect 23001 35990 23027 36021
rect 23075 35990 23107 36021
rect 23107 35990 23109 36021
rect 23157 35990 23177 36021
rect 23177 35990 23191 36021
rect 23239 35990 23247 36021
rect 23247 35990 23273 36021
rect 22829 35919 22861 35952
rect 22861 35919 22863 35952
rect 22911 35919 22931 35952
rect 22931 35919 22945 35952
rect 22993 35919 23001 35952
rect 23001 35919 23027 35952
rect 23075 35919 23107 35952
rect 23107 35919 23109 35952
rect 23157 35919 23177 35952
rect 23177 35919 23191 35952
rect 23239 35919 23247 35952
rect 23247 35919 23273 35952
rect 22829 35918 22863 35919
rect 22911 35918 22945 35919
rect 22993 35918 23027 35919
rect 23075 35918 23109 35919
rect 23157 35918 23191 35919
rect 23239 35918 23273 35919
rect 22829 35851 22861 35880
rect 22861 35851 22863 35880
rect 22911 35851 22931 35880
rect 22931 35851 22945 35880
rect 22993 35851 23001 35880
rect 23001 35851 23027 35880
rect 23075 35851 23107 35880
rect 23107 35851 23109 35880
rect 23157 35851 23177 35880
rect 23177 35851 23191 35880
rect 23239 35851 23247 35880
rect 23247 35851 23273 35880
rect 22829 35846 22863 35851
rect 22911 35846 22945 35851
rect 22993 35846 23027 35851
rect 23075 35846 23109 35851
rect 23157 35846 23191 35851
rect 23239 35846 23273 35851
rect 22829 35783 22861 35808
rect 22861 35783 22863 35808
rect 22911 35783 22931 35808
rect 22931 35783 22945 35808
rect 22993 35783 23001 35808
rect 23001 35783 23027 35808
rect 23075 35783 23107 35808
rect 23107 35783 23109 35808
rect 23157 35783 23177 35808
rect 23177 35783 23191 35808
rect 23239 35783 23247 35808
rect 23247 35783 23273 35808
rect 22829 35774 22863 35783
rect 22911 35774 22945 35783
rect 22993 35774 23027 35783
rect 23075 35774 23109 35783
rect 23157 35774 23191 35783
rect 23239 35774 23273 35783
rect 22829 35715 22861 35736
rect 22861 35715 22863 35736
rect 22911 35715 22931 35736
rect 22931 35715 22945 35736
rect 22993 35715 23001 35736
rect 23001 35715 23027 35736
rect 23075 35715 23107 35736
rect 23107 35715 23109 35736
rect 23157 35715 23177 35736
rect 23177 35715 23191 35736
rect 23239 35715 23247 35736
rect 23247 35715 23273 35736
rect 22829 35702 22863 35715
rect 22911 35702 22945 35715
rect 22993 35702 23027 35715
rect 23075 35702 23109 35715
rect 23157 35702 23191 35715
rect 23239 35702 23273 35715
rect 209 35610 243 35644
rect 291 35619 325 35644
rect 291 35610 312 35619
rect 312 35610 325 35619
rect 209 35538 243 35572
rect 291 35551 325 35572
rect 291 35538 312 35551
rect 312 35538 325 35551
rect 209 35466 243 35500
rect 291 35483 325 35500
rect 291 35466 312 35483
rect 312 35466 325 35483
rect 209 35393 243 35427
rect 291 35415 325 35427
rect 291 35393 312 35415
rect 312 35393 325 35415
rect 209 35320 243 35354
rect 291 35347 325 35354
rect 291 35320 312 35347
rect 312 35320 325 35347
rect 209 35247 243 35281
rect 291 35279 325 35281
rect 291 35247 312 35279
rect 312 35247 325 35279
rect 209 35174 243 35208
rect 291 35177 312 35208
rect 312 35177 325 35208
rect 291 35174 325 35177
rect 209 35101 243 35135
rect 291 35109 312 35135
rect 312 35109 325 35135
rect 291 35101 325 35109
rect 209 35028 243 35062
rect 291 35041 312 35062
rect 312 35041 325 35062
rect 291 35028 325 35041
rect 209 34955 243 34989
rect 291 34972 312 34989
rect 312 34972 325 34989
rect 291 34955 325 34972
rect 209 34882 243 34916
rect 291 34903 312 34916
rect 312 34903 325 34916
rect 291 34882 325 34903
rect 209 34809 243 34843
rect 291 34834 312 34843
rect 312 34834 325 34843
rect 291 34809 325 34834
rect 209 34736 243 34770
rect 291 34765 312 34770
rect 312 34765 325 34770
rect 291 34736 325 34765
rect 209 34663 243 34697
rect 291 34696 312 34697
rect 312 34696 325 34697
rect 291 34663 325 34696
rect 209 34590 243 34624
rect 291 34592 325 34624
rect 291 34590 312 34592
rect 312 34590 325 34592
rect 209 34517 243 34551
rect 291 34523 325 34551
rect 291 34517 312 34523
rect 312 34517 325 34523
rect 209 34444 243 34478
rect 291 34454 325 34478
rect 291 34444 312 34454
rect 312 34444 325 34454
rect 209 34371 243 34405
rect 291 34385 325 34405
rect 291 34371 312 34385
rect 312 34371 325 34385
rect 209 34298 243 34332
rect 291 34316 325 34332
rect 291 34298 312 34316
rect 312 34298 325 34316
rect 209 34225 243 34259
rect 291 34247 325 34259
rect 291 34225 312 34247
rect 312 34225 325 34247
rect 209 34152 243 34186
rect 291 34178 325 34186
rect 291 34152 312 34178
rect 312 34152 325 34178
rect 209 34079 243 34113
rect 291 34109 325 34113
rect 291 34079 312 34109
rect 312 34079 325 34109
rect 209 34006 243 34040
rect 291 34006 312 34040
rect 312 34006 325 34040
rect 209 33933 243 33967
rect 291 33937 312 33967
rect 312 33937 325 33967
rect 291 33933 325 33937
rect 209 33860 243 33894
rect 291 33868 312 33894
rect 312 33868 325 33894
rect 291 33860 325 33868
rect 209 33787 243 33821
rect 291 33799 312 33821
rect 312 33799 325 33821
rect 291 33787 325 33799
rect 209 33714 243 33748
rect 291 33730 312 33748
rect 312 33730 325 33748
rect 291 33714 325 33730
rect 209 33641 243 33675
rect 291 33661 312 33675
rect 312 33661 325 33675
rect 291 33641 325 33661
rect 209 33568 243 33602
rect 291 33592 312 33602
rect 312 33592 325 33602
rect 291 33568 325 33592
rect 209 33495 243 33529
rect 291 33523 312 33529
rect 312 33523 325 33529
rect 291 33495 325 33523
rect 209 33422 243 33456
rect 291 33454 312 33456
rect 312 33454 325 33456
rect 291 33422 325 33454
rect 209 33349 243 33383
rect 291 33350 325 33383
rect 291 33349 312 33350
rect 312 33349 325 33350
rect 22829 35647 22861 35664
rect 22861 35647 22863 35664
rect 22911 35647 22931 35664
rect 22931 35647 22945 35664
rect 22993 35647 23001 35664
rect 23001 35647 23027 35664
rect 23075 35647 23107 35664
rect 23107 35647 23109 35664
rect 23157 35647 23177 35664
rect 23177 35647 23191 35664
rect 23239 35647 23247 35664
rect 23247 35647 23273 35664
rect 22829 35630 22863 35647
rect 22911 35630 22945 35647
rect 22993 35630 23027 35647
rect 23075 35630 23109 35647
rect 23157 35630 23191 35647
rect 23239 35630 23273 35647
rect 22829 35579 22861 35592
rect 22861 35579 22863 35592
rect 22911 35579 22931 35592
rect 22931 35579 22945 35592
rect 22993 35579 23001 35592
rect 23001 35579 23027 35592
rect 23075 35579 23107 35592
rect 23107 35579 23109 35592
rect 23157 35579 23177 35592
rect 23177 35579 23191 35592
rect 23239 35579 23247 35592
rect 23247 35579 23273 35592
rect 22829 35558 22863 35579
rect 22911 35558 22945 35579
rect 22993 35558 23027 35579
rect 23075 35558 23109 35579
rect 23157 35558 23191 35579
rect 23239 35558 23273 35579
rect 22829 35511 22861 35520
rect 22861 35511 22863 35520
rect 22911 35511 22931 35520
rect 22931 35511 22945 35520
rect 22993 35511 23001 35520
rect 23001 35511 23027 35520
rect 23075 35511 23107 35520
rect 23107 35511 23109 35520
rect 23157 35511 23177 35520
rect 23177 35511 23191 35520
rect 23239 35511 23247 35520
rect 23247 35511 23273 35520
rect 22829 35486 22863 35511
rect 22911 35486 22945 35511
rect 22993 35486 23027 35511
rect 23075 35486 23109 35511
rect 23157 35486 23191 35511
rect 23239 35486 23273 35511
rect 22829 35443 22861 35448
rect 22861 35443 22863 35448
rect 22911 35443 22931 35448
rect 22931 35443 22945 35448
rect 22993 35443 23001 35448
rect 23001 35443 23027 35448
rect 23075 35443 23107 35448
rect 23107 35443 23109 35448
rect 23157 35443 23177 35448
rect 23177 35443 23191 35448
rect 23239 35443 23247 35448
rect 23247 35443 23273 35448
rect 22829 35414 22863 35443
rect 22911 35414 22945 35443
rect 22993 35414 23027 35443
rect 23075 35414 23109 35443
rect 23157 35414 23191 35443
rect 23239 35414 23273 35443
rect 22829 35375 22861 35376
rect 22861 35375 22863 35376
rect 22911 35375 22931 35376
rect 22931 35375 22945 35376
rect 22993 35375 23001 35376
rect 23001 35375 23027 35376
rect 23075 35375 23107 35376
rect 23107 35375 23109 35376
rect 23157 35375 23177 35376
rect 23177 35375 23191 35376
rect 23239 35375 23247 35376
rect 23247 35375 23273 35376
rect 22829 35342 22863 35375
rect 22911 35342 22945 35375
rect 22993 35342 23027 35375
rect 23075 35342 23109 35375
rect 23157 35342 23191 35375
rect 23239 35342 23273 35375
rect 22829 35273 22863 35304
rect 22911 35273 22945 35304
rect 22993 35273 23027 35304
rect 23075 35273 23109 35304
rect 23157 35273 23191 35304
rect 23239 35273 23273 35304
rect 22829 35270 22861 35273
rect 22861 35270 22863 35273
rect 22911 35270 22931 35273
rect 22931 35270 22945 35273
rect 22993 35270 23001 35273
rect 23001 35270 23027 35273
rect 23075 35270 23107 35273
rect 23107 35270 23109 35273
rect 23157 35270 23177 35273
rect 23177 35270 23191 35273
rect 23239 35270 23247 35273
rect 23247 35270 23273 35273
rect 22829 35205 22863 35232
rect 22911 35205 22945 35232
rect 22993 35205 23027 35232
rect 23075 35205 23109 35232
rect 23157 35205 23191 35232
rect 23239 35205 23273 35232
rect 22829 35198 22861 35205
rect 22861 35198 22863 35205
rect 22911 35198 22931 35205
rect 22931 35198 22945 35205
rect 22993 35198 23001 35205
rect 23001 35198 23027 35205
rect 23075 35198 23107 35205
rect 23107 35198 23109 35205
rect 23157 35198 23177 35205
rect 23177 35198 23191 35205
rect 23239 35198 23247 35205
rect 23247 35198 23273 35205
rect 22829 35137 22863 35160
rect 22911 35137 22945 35160
rect 22993 35137 23027 35160
rect 23075 35137 23109 35160
rect 23157 35137 23191 35160
rect 23239 35137 23273 35160
rect 22829 35126 22861 35137
rect 22861 35126 22863 35137
rect 22911 35126 22931 35137
rect 22931 35126 22945 35137
rect 22993 35126 23001 35137
rect 23001 35126 23027 35137
rect 23075 35126 23107 35137
rect 23107 35126 23109 35137
rect 23157 35126 23177 35137
rect 23177 35126 23191 35137
rect 23239 35126 23247 35137
rect 23247 35126 23273 35137
rect 22829 35069 22863 35088
rect 22911 35069 22945 35088
rect 22993 35069 23027 35088
rect 23075 35069 23109 35088
rect 23157 35069 23191 35088
rect 23239 35069 23273 35088
rect 22829 35054 22861 35069
rect 22861 35054 22863 35069
rect 22911 35054 22931 35069
rect 22931 35054 22945 35069
rect 22993 35054 23001 35069
rect 23001 35054 23027 35069
rect 23075 35054 23107 35069
rect 23107 35054 23109 35069
rect 23157 35054 23177 35069
rect 23177 35054 23191 35069
rect 23239 35054 23247 35069
rect 23247 35054 23273 35069
rect 22829 35001 22863 35016
rect 22911 35001 22945 35016
rect 22993 35001 23027 35016
rect 23075 35001 23109 35016
rect 23157 35001 23191 35016
rect 23239 35001 23273 35016
rect 22829 34982 22861 35001
rect 22861 34982 22863 35001
rect 22911 34982 22931 35001
rect 22931 34982 22945 35001
rect 22993 34982 23001 35001
rect 23001 34982 23027 35001
rect 23075 34982 23107 35001
rect 23107 34982 23109 35001
rect 23157 34982 23177 35001
rect 23177 34982 23191 35001
rect 23239 34982 23247 35001
rect 23247 34982 23273 35001
rect 22829 34933 22863 34944
rect 22911 34933 22945 34944
rect 22993 34933 23027 34944
rect 23075 34933 23109 34944
rect 23157 34933 23191 34944
rect 23239 34933 23273 34944
rect 22829 34910 22861 34933
rect 22861 34910 22863 34933
rect 22911 34910 22931 34933
rect 22931 34910 22945 34933
rect 22993 34910 23001 34933
rect 23001 34910 23027 34933
rect 23075 34910 23107 34933
rect 23107 34910 23109 34933
rect 23157 34910 23177 34933
rect 23177 34910 23191 34933
rect 23239 34910 23247 34933
rect 23247 34910 23273 34933
rect 22829 34865 22863 34872
rect 22911 34865 22945 34872
rect 22993 34865 23027 34872
rect 23075 34865 23109 34872
rect 23157 34865 23191 34872
rect 23239 34865 23273 34872
rect 22829 34838 22861 34865
rect 22861 34838 22863 34865
rect 22911 34838 22931 34865
rect 22931 34838 22945 34865
rect 22993 34838 23001 34865
rect 23001 34838 23027 34865
rect 23075 34838 23107 34865
rect 23107 34838 23109 34865
rect 23157 34838 23177 34865
rect 23177 34838 23191 34865
rect 23239 34838 23247 34865
rect 23247 34838 23273 34865
rect 22829 34797 22863 34800
rect 22911 34797 22945 34800
rect 22993 34797 23027 34800
rect 23075 34797 23109 34800
rect 23157 34797 23191 34800
rect 23239 34797 23273 34800
rect 22829 34766 22861 34797
rect 22861 34766 22863 34797
rect 22911 34766 22931 34797
rect 22931 34766 22945 34797
rect 22993 34766 23001 34797
rect 23001 34766 23027 34797
rect 23075 34766 23107 34797
rect 23107 34766 23109 34797
rect 23157 34766 23177 34797
rect 23177 34766 23191 34797
rect 23239 34766 23247 34797
rect 23247 34766 23273 34797
rect 22829 34695 22861 34728
rect 22861 34695 22863 34728
rect 22911 34695 22931 34728
rect 22931 34695 22945 34728
rect 22993 34695 23001 34728
rect 23001 34695 23027 34728
rect 23075 34695 23107 34728
rect 23107 34695 23109 34728
rect 23157 34695 23177 34728
rect 23177 34695 23191 34728
rect 23239 34695 23247 34728
rect 23247 34695 23273 34728
rect 22829 34694 22863 34695
rect 22911 34694 22945 34695
rect 22993 34694 23027 34695
rect 23075 34694 23109 34695
rect 23157 34694 23191 34695
rect 23239 34694 23273 34695
rect 22829 34627 22861 34656
rect 22861 34627 22863 34656
rect 22911 34627 22931 34656
rect 22931 34627 22945 34656
rect 22993 34627 23001 34656
rect 23001 34627 23027 34656
rect 23075 34627 23107 34656
rect 23107 34627 23109 34656
rect 23157 34627 23177 34656
rect 23177 34627 23191 34656
rect 23239 34627 23247 34656
rect 23247 34627 23273 34656
rect 22829 34622 22863 34627
rect 22911 34622 22945 34627
rect 22993 34622 23027 34627
rect 23075 34622 23109 34627
rect 23157 34622 23191 34627
rect 23239 34622 23273 34627
rect 22829 34559 22861 34584
rect 22861 34559 22863 34584
rect 22911 34559 22931 34584
rect 22931 34559 22945 34584
rect 22993 34559 23001 34584
rect 23001 34559 23027 34584
rect 23075 34559 23107 34584
rect 23107 34559 23109 34584
rect 23157 34559 23177 34584
rect 23177 34559 23191 34584
rect 23239 34559 23247 34584
rect 23247 34559 23273 34584
rect 22829 34550 22863 34559
rect 22911 34550 22945 34559
rect 22993 34550 23027 34559
rect 23075 34550 23109 34559
rect 23157 34550 23191 34559
rect 23239 34550 23273 34559
rect 22829 34491 22861 34512
rect 22861 34491 22863 34512
rect 22911 34491 22931 34512
rect 22931 34491 22945 34512
rect 22993 34491 23001 34512
rect 23001 34491 23027 34512
rect 23075 34491 23107 34512
rect 23107 34491 23109 34512
rect 23157 34491 23177 34512
rect 23177 34491 23191 34512
rect 23239 34491 23247 34512
rect 23247 34491 23273 34512
rect 22829 34478 22863 34491
rect 22911 34478 22945 34491
rect 22993 34478 23027 34491
rect 23075 34478 23109 34491
rect 23157 34478 23191 34491
rect 23239 34478 23273 34491
rect 22829 34423 22861 34440
rect 22861 34423 22863 34440
rect 22911 34423 22931 34440
rect 22931 34423 22945 34440
rect 22993 34423 23001 34440
rect 23001 34423 23027 34440
rect 23075 34423 23107 34440
rect 23107 34423 23109 34440
rect 23157 34423 23177 34440
rect 23177 34423 23191 34440
rect 23239 34423 23247 34440
rect 23247 34423 23273 34440
rect 22829 34406 22863 34423
rect 22911 34406 22945 34423
rect 22993 34406 23027 34423
rect 23075 34406 23109 34423
rect 23157 34406 23191 34423
rect 23239 34406 23273 34423
rect 22829 34355 22861 34368
rect 22861 34355 22863 34368
rect 22911 34355 22931 34368
rect 22931 34355 22945 34368
rect 22993 34355 23001 34368
rect 23001 34355 23027 34368
rect 23075 34355 23107 34368
rect 23107 34355 23109 34368
rect 23157 34355 23177 34368
rect 23177 34355 23191 34368
rect 23239 34355 23247 34368
rect 23247 34355 23273 34368
rect 22829 34334 22863 34355
rect 22911 34334 22945 34355
rect 22993 34334 23027 34355
rect 23075 34334 23109 34355
rect 23157 34334 23191 34355
rect 23239 34334 23273 34355
rect 22829 34287 22861 34295
rect 22861 34287 22863 34295
rect 22911 34287 22931 34295
rect 22931 34287 22945 34295
rect 22993 34287 23001 34295
rect 23001 34287 23027 34295
rect 23075 34287 23107 34295
rect 23107 34287 23109 34295
rect 23157 34287 23177 34295
rect 23177 34287 23191 34295
rect 23239 34287 23247 34295
rect 23247 34287 23273 34295
rect 22829 34261 22863 34287
rect 22911 34261 22945 34287
rect 22993 34261 23027 34287
rect 23075 34261 23109 34287
rect 23157 34261 23191 34287
rect 23239 34261 23273 34287
rect 22829 34219 22861 34222
rect 22861 34219 22863 34222
rect 22911 34219 22931 34222
rect 22931 34219 22945 34222
rect 22993 34219 23001 34222
rect 23001 34219 23027 34222
rect 23075 34219 23107 34222
rect 23107 34219 23109 34222
rect 23157 34219 23177 34222
rect 23177 34219 23191 34222
rect 23239 34219 23247 34222
rect 23247 34219 23273 34222
rect 22829 34188 22863 34219
rect 22911 34188 22945 34219
rect 22993 34188 23027 34219
rect 23075 34188 23109 34219
rect 23157 34188 23191 34219
rect 23239 34188 23273 34219
rect 22829 34117 22863 34149
rect 22911 34117 22945 34149
rect 22993 34117 23027 34149
rect 23075 34117 23109 34149
rect 23157 34117 23191 34149
rect 23239 34117 23273 34149
rect 22829 34115 22861 34117
rect 22861 34115 22863 34117
rect 22911 34115 22931 34117
rect 22931 34115 22945 34117
rect 22993 34115 23001 34117
rect 23001 34115 23027 34117
rect 23075 34115 23107 34117
rect 23107 34115 23109 34117
rect 23157 34115 23177 34117
rect 23177 34115 23191 34117
rect 23239 34115 23247 34117
rect 23247 34115 23273 34117
rect 22829 34049 22863 34076
rect 22911 34049 22945 34076
rect 22993 34049 23027 34076
rect 23075 34049 23109 34076
rect 23157 34049 23191 34076
rect 23239 34049 23273 34076
rect 22829 34042 22861 34049
rect 22861 34042 22863 34049
rect 22911 34042 22931 34049
rect 22931 34042 22945 34049
rect 22993 34042 23001 34049
rect 23001 34042 23027 34049
rect 23075 34042 23107 34049
rect 23107 34042 23109 34049
rect 23157 34042 23177 34049
rect 23177 34042 23191 34049
rect 23239 34042 23247 34049
rect 23247 34042 23273 34049
rect 22829 33981 22863 34003
rect 22911 33981 22945 34003
rect 22993 33981 23027 34003
rect 23075 33981 23109 34003
rect 23157 33981 23191 34003
rect 23239 33981 23273 34003
rect 22829 33969 22861 33981
rect 22861 33969 22863 33981
rect 22911 33969 22931 33981
rect 22931 33969 22945 33981
rect 22993 33969 23001 33981
rect 23001 33969 23027 33981
rect 23075 33969 23107 33981
rect 23107 33969 23109 33981
rect 23157 33969 23177 33981
rect 23177 33969 23191 33981
rect 23239 33969 23247 33981
rect 23247 33969 23273 33981
rect 22829 33913 22863 33930
rect 22911 33913 22945 33930
rect 22993 33913 23027 33930
rect 23075 33913 23109 33930
rect 23157 33913 23191 33930
rect 23239 33913 23273 33930
rect 22829 33896 22861 33913
rect 22861 33896 22863 33913
rect 22911 33896 22931 33913
rect 22931 33896 22945 33913
rect 22993 33896 23001 33913
rect 23001 33896 23027 33913
rect 23075 33896 23107 33913
rect 23107 33896 23109 33913
rect 23157 33896 23177 33913
rect 23177 33896 23191 33913
rect 23239 33896 23247 33913
rect 23247 33896 23273 33913
rect 22829 33845 22863 33857
rect 22911 33845 22945 33857
rect 22993 33845 23027 33857
rect 23075 33845 23109 33857
rect 23157 33845 23191 33857
rect 23239 33845 23273 33857
rect 22829 33823 22861 33845
rect 22861 33823 22863 33845
rect 22911 33823 22931 33845
rect 22931 33823 22945 33845
rect 22993 33823 23001 33845
rect 23001 33823 23027 33845
rect 23075 33823 23107 33845
rect 23107 33823 23109 33845
rect 23157 33823 23177 33845
rect 23177 33823 23191 33845
rect 23239 33823 23247 33845
rect 23247 33823 23273 33845
rect 22829 33777 22863 33784
rect 22911 33777 22945 33784
rect 22993 33777 23027 33784
rect 23075 33777 23109 33784
rect 23157 33777 23191 33784
rect 23239 33777 23273 33784
rect 22829 33750 22861 33777
rect 22861 33750 22863 33777
rect 22911 33750 22931 33777
rect 22931 33750 22945 33777
rect 22993 33750 23001 33777
rect 23001 33750 23027 33777
rect 23075 33750 23107 33777
rect 23107 33750 23109 33777
rect 23157 33750 23177 33777
rect 23177 33750 23191 33777
rect 23239 33750 23247 33777
rect 23247 33750 23273 33777
rect 22829 33709 22863 33711
rect 22911 33709 22945 33711
rect 22993 33709 23027 33711
rect 23075 33709 23109 33711
rect 23157 33709 23191 33711
rect 23239 33709 23273 33711
rect 22829 33677 22861 33709
rect 22861 33677 22863 33709
rect 22911 33677 22931 33709
rect 22931 33677 22945 33709
rect 22993 33677 23001 33709
rect 23001 33677 23027 33709
rect 23075 33677 23107 33709
rect 23107 33677 23109 33709
rect 23157 33677 23177 33709
rect 23177 33677 23191 33709
rect 23239 33677 23247 33709
rect 23247 33677 23273 33709
rect 22829 33607 22861 33638
rect 22861 33607 22863 33638
rect 22911 33607 22931 33638
rect 22931 33607 22945 33638
rect 22993 33607 23001 33638
rect 23001 33607 23027 33638
rect 23075 33607 23107 33638
rect 23107 33607 23109 33638
rect 23157 33607 23177 33638
rect 23177 33607 23191 33638
rect 23239 33607 23247 33638
rect 23247 33607 23273 33638
rect 22829 33604 22863 33607
rect 22911 33604 22945 33607
rect 22993 33604 23027 33607
rect 23075 33604 23109 33607
rect 23157 33604 23191 33607
rect 23239 33604 23273 33607
rect 22829 33539 22861 33565
rect 22861 33539 22863 33565
rect 22911 33539 22931 33565
rect 22931 33539 22945 33565
rect 22993 33539 23001 33565
rect 23001 33539 23027 33565
rect 23075 33539 23107 33565
rect 23107 33539 23109 33565
rect 23157 33539 23177 33565
rect 23177 33539 23191 33565
rect 23239 33539 23247 33565
rect 23247 33539 23273 33565
rect 22829 33531 22863 33539
rect 22911 33531 22945 33539
rect 22993 33531 23027 33539
rect 23075 33531 23109 33539
rect 23157 33531 23191 33539
rect 23239 33531 23273 33539
rect 22829 33471 22861 33492
rect 22861 33471 22863 33492
rect 22911 33471 22931 33492
rect 22931 33471 22945 33492
rect 22993 33471 23001 33492
rect 23001 33471 23027 33492
rect 23075 33471 23107 33492
rect 23107 33471 23109 33492
rect 23157 33471 23177 33492
rect 23177 33471 23191 33492
rect 23239 33471 23247 33492
rect 23247 33471 23273 33492
rect 22829 33458 22863 33471
rect 22911 33458 22945 33471
rect 22993 33458 23027 33471
rect 23075 33458 23109 33471
rect 23157 33458 23191 33471
rect 23239 33458 23273 33471
rect 22829 33403 22861 33419
rect 22861 33403 22863 33419
rect 22911 33403 22931 33419
rect 22931 33403 22945 33419
rect 22993 33403 23001 33419
rect 23001 33403 23027 33419
rect 23075 33403 23107 33419
rect 23107 33403 23109 33419
rect 23157 33403 23177 33419
rect 23177 33403 23191 33419
rect 23239 33403 23247 33419
rect 23247 33403 23273 33419
rect 22829 33385 22863 33403
rect 22911 33385 22945 33403
rect 22993 33385 23027 33403
rect 23075 33385 23109 33403
rect 23157 33385 23191 33403
rect 23239 33385 23273 33403
rect 22829 33335 22861 33346
rect 22861 33335 22863 33346
rect 22911 33335 22931 33346
rect 22931 33335 22945 33346
rect 22993 33335 23001 33346
rect 23001 33335 23027 33346
rect 23075 33335 23107 33346
rect 23107 33335 23109 33346
rect 23157 33335 23177 33346
rect 23177 33335 23191 33346
rect 23239 33335 23247 33346
rect 23247 33335 23273 33346
rect 209 33276 243 33310
rect 291 33281 325 33310
rect 291 33276 312 33281
rect 312 33276 325 33281
rect 209 33203 243 33237
rect 291 33212 325 33237
rect 291 33203 312 33212
rect 312 33203 325 33212
rect 209 33130 243 33164
rect 291 33143 325 33164
rect 291 33130 312 33143
rect 312 33130 325 33143
rect 209 33057 243 33091
rect 291 33074 325 33091
rect 291 33057 312 33074
rect 312 33057 325 33074
rect 209 32984 243 33018
rect 291 33005 325 33018
rect 291 32984 312 33005
rect 312 32984 325 33005
rect 209 32911 243 32945
rect 291 32936 325 32945
rect 291 32911 312 32936
rect 312 32911 325 32936
rect 209 32838 243 32872
rect 291 32867 325 32872
rect 291 32838 312 32867
rect 312 32838 325 32867
rect 209 32765 243 32799
rect 291 32798 325 32799
rect 291 32765 312 32798
rect 312 32765 325 32798
rect 209 32692 243 32726
rect 291 32695 312 32726
rect 312 32695 325 32726
rect 291 32692 325 32695
rect 209 32619 243 32653
rect 291 32626 312 32653
rect 312 32626 325 32653
rect 291 32619 325 32626
rect 209 32546 243 32580
rect 291 32557 312 32580
rect 312 32557 325 32580
rect 291 32546 325 32557
rect 209 32473 243 32507
rect 291 32488 312 32507
rect 312 32488 325 32507
rect 291 32473 325 32488
rect 209 32400 243 32434
rect 291 32419 312 32434
rect 312 32419 325 32434
rect 291 32400 325 32419
rect 209 32327 243 32361
rect 291 32350 312 32361
rect 312 32350 325 32361
rect 291 32327 325 32350
rect 18022 33307 18056 33328
rect 18108 33307 18142 33328
rect 18194 33307 18228 33328
rect 18280 33307 18314 33328
rect 18022 33294 18025 33307
rect 18025 33294 18056 33307
rect 18108 33294 18135 33307
rect 18135 33294 18142 33307
rect 18194 33294 18211 33307
rect 18211 33294 18228 33307
rect 18280 33294 18287 33307
rect 18287 33294 18314 33307
rect 18366 33294 18400 33328
rect 18022 33239 18056 33256
rect 18108 33239 18142 33256
rect 18194 33239 18228 33256
rect 18280 33239 18314 33256
rect 18022 33222 18025 33239
rect 18025 33222 18056 33239
rect 18108 33222 18135 33239
rect 18135 33222 18142 33239
rect 18194 33222 18211 33239
rect 18211 33222 18228 33239
rect 18280 33222 18287 33239
rect 18287 33222 18314 33239
rect 18366 33222 18400 33256
rect 18022 33171 18056 33184
rect 18108 33171 18142 33184
rect 18194 33171 18228 33184
rect 18280 33171 18314 33184
rect 18022 33150 18025 33171
rect 18025 33150 18056 33171
rect 18108 33150 18135 33171
rect 18135 33150 18142 33171
rect 18194 33150 18211 33171
rect 18211 33150 18228 33171
rect 18280 33150 18287 33171
rect 18287 33150 18314 33171
rect 18366 33150 18400 33184
rect 18022 33103 18056 33112
rect 18108 33103 18142 33112
rect 18194 33103 18228 33112
rect 18280 33103 18314 33112
rect 18022 33078 18025 33103
rect 18025 33078 18056 33103
rect 18108 33078 18135 33103
rect 18135 33078 18142 33103
rect 18194 33078 18211 33103
rect 18211 33078 18228 33103
rect 18280 33078 18287 33103
rect 18287 33078 18314 33103
rect 18366 33078 18400 33112
rect 18022 33035 18056 33040
rect 18108 33035 18142 33040
rect 18194 33035 18228 33040
rect 18280 33035 18314 33040
rect 18022 33006 18025 33035
rect 18025 33006 18056 33035
rect 18108 33006 18135 33035
rect 18135 33006 18142 33035
rect 18194 33006 18211 33035
rect 18211 33006 18228 33035
rect 18280 33006 18287 33035
rect 18287 33006 18314 33035
rect 18366 33006 18400 33040
rect 18022 32967 18056 32968
rect 18108 32967 18142 32968
rect 18194 32967 18228 32968
rect 18280 32967 18314 32968
rect 18022 32934 18025 32967
rect 18025 32934 18056 32967
rect 18108 32934 18135 32967
rect 18135 32934 18142 32967
rect 18194 32934 18211 32967
rect 18211 32934 18228 32967
rect 18280 32934 18287 32967
rect 18287 32934 18314 32967
rect 18366 32934 18400 32968
rect 18022 32865 18025 32896
rect 18025 32865 18056 32896
rect 18108 32865 18135 32896
rect 18135 32865 18142 32896
rect 18194 32865 18211 32896
rect 18211 32865 18228 32896
rect 18280 32865 18287 32896
rect 18287 32865 18314 32896
rect 18022 32862 18056 32865
rect 18108 32862 18142 32865
rect 18194 32862 18228 32865
rect 18280 32862 18314 32865
rect 18366 32862 18400 32896
rect 18022 32797 18025 32824
rect 18025 32797 18056 32824
rect 18108 32797 18135 32824
rect 18135 32797 18142 32824
rect 18194 32797 18211 32824
rect 18211 32797 18228 32824
rect 18280 32797 18287 32824
rect 18287 32797 18314 32824
rect 18022 32790 18056 32797
rect 18108 32790 18142 32797
rect 18194 32790 18228 32797
rect 18280 32790 18314 32797
rect 18366 32790 18400 32824
rect 18022 32729 18025 32752
rect 18025 32729 18056 32752
rect 18108 32729 18135 32752
rect 18135 32729 18142 32752
rect 18194 32729 18211 32752
rect 18211 32729 18228 32752
rect 18280 32729 18287 32752
rect 18287 32729 18314 32752
rect 18022 32718 18056 32729
rect 18108 32718 18142 32729
rect 18194 32718 18228 32729
rect 18280 32718 18314 32729
rect 18366 32718 18400 32752
rect 18022 32661 18025 32680
rect 18025 32661 18056 32680
rect 18108 32661 18135 32680
rect 18135 32661 18142 32680
rect 18194 32661 18211 32680
rect 18211 32661 18228 32680
rect 18280 32661 18287 32680
rect 18287 32661 18314 32680
rect 18022 32646 18056 32661
rect 18108 32646 18142 32661
rect 18194 32646 18228 32661
rect 18280 32646 18314 32661
rect 18366 32646 18400 32680
rect 18022 32593 18025 32608
rect 18025 32593 18056 32608
rect 18108 32593 18135 32608
rect 18135 32593 18142 32608
rect 18194 32593 18211 32608
rect 18211 32593 18228 32608
rect 18280 32593 18287 32608
rect 18287 32593 18314 32608
rect 18022 32574 18056 32593
rect 18108 32574 18142 32593
rect 18194 32574 18228 32593
rect 18280 32574 18314 32593
rect 18366 32574 18400 32608
rect 18022 32525 18025 32536
rect 18025 32525 18056 32536
rect 18108 32525 18135 32536
rect 18135 32525 18142 32536
rect 18194 32525 18211 32536
rect 18211 32525 18228 32536
rect 18280 32525 18287 32536
rect 18287 32525 18314 32536
rect 18022 32502 18056 32525
rect 18108 32502 18142 32525
rect 18194 32502 18228 32525
rect 18280 32502 18314 32525
rect 18366 32502 18400 32536
rect 18022 32457 18025 32464
rect 18025 32457 18056 32464
rect 18108 32457 18135 32464
rect 18135 32457 18142 32464
rect 18194 32457 18211 32464
rect 18211 32457 18228 32464
rect 18280 32457 18287 32464
rect 18287 32457 18314 32464
rect 18022 32430 18056 32457
rect 18108 32430 18142 32457
rect 18194 32430 18228 32457
rect 18280 32430 18314 32457
rect 18366 32430 18400 32464
rect 18022 32389 18025 32392
rect 18025 32389 18056 32392
rect 18108 32389 18135 32392
rect 18135 32389 18142 32392
rect 18194 32389 18211 32392
rect 18211 32389 18228 32392
rect 18280 32389 18287 32392
rect 18287 32389 18314 32392
rect 18022 32358 18056 32389
rect 18108 32358 18142 32389
rect 18194 32358 18228 32389
rect 18280 32358 18314 32389
rect 18366 32358 18400 32392
rect 209 32254 243 32288
rect 291 32281 312 32288
rect 312 32281 325 32288
rect 291 32254 325 32281
rect 209 32181 243 32215
rect 291 32212 312 32215
rect 312 32212 325 32215
rect 291 32181 325 32212
rect 209 32108 243 32142
rect 291 32108 325 32142
rect 218 32030 252 32064
rect 218 31958 252 31992
rect 218 31886 252 31920
rect 218 31814 252 31848
rect 218 31742 252 31776
rect 18022 32287 18056 32320
rect 18108 32287 18142 32320
rect 18194 32287 18228 32320
rect 18280 32287 18314 32320
rect 18022 32286 18025 32287
rect 18025 32286 18056 32287
rect 18108 32286 18135 32287
rect 18135 32286 18142 32287
rect 18194 32286 18211 32287
rect 18211 32286 18228 32287
rect 18280 32286 18287 32287
rect 18287 32286 18314 32287
rect 18366 32286 18400 32320
rect 18022 32219 18056 32248
rect 18108 32219 18142 32248
rect 18194 32219 18228 32248
rect 18280 32219 18314 32248
rect 18022 32214 18025 32219
rect 18025 32214 18056 32219
rect 18108 32214 18135 32219
rect 18135 32214 18142 32219
rect 18194 32214 18211 32219
rect 18211 32214 18228 32219
rect 18280 32214 18287 32219
rect 18287 32214 18314 32219
rect 18366 32214 18400 32248
rect 18022 32151 18056 32176
rect 18108 32151 18142 32176
rect 18194 32151 18228 32176
rect 18280 32151 18314 32176
rect 18022 32142 18025 32151
rect 18025 32142 18056 32151
rect 18108 32142 18135 32151
rect 18135 32142 18142 32151
rect 18194 32142 18211 32151
rect 18211 32142 18228 32151
rect 18280 32142 18287 32151
rect 18287 32142 18314 32151
rect 18366 32142 18400 32176
rect 18022 32083 18056 32104
rect 18108 32083 18142 32104
rect 18194 32083 18228 32104
rect 18280 32083 18314 32104
rect 18022 32070 18025 32083
rect 18025 32070 18056 32083
rect 18108 32070 18135 32083
rect 18135 32070 18142 32083
rect 18194 32070 18211 32083
rect 18211 32070 18228 32083
rect 18280 32070 18287 32083
rect 18287 32070 18314 32083
rect 18366 32070 18400 32104
rect 18022 32015 18056 32032
rect 18108 32015 18142 32032
rect 18194 32015 18228 32032
rect 18280 32015 18314 32032
rect 18022 31998 18025 32015
rect 18025 31998 18056 32015
rect 18108 31998 18135 32015
rect 18135 31998 18142 32015
rect 18194 31998 18211 32015
rect 18211 31998 18228 32015
rect 18280 31998 18287 32015
rect 18287 31998 18314 32015
rect 18366 31998 18400 32032
rect 18022 31947 18056 31960
rect 18108 31947 18142 31960
rect 18194 31947 18228 31960
rect 18280 31947 18314 31960
rect 18022 31926 18025 31947
rect 18025 31926 18056 31947
rect 18108 31926 18135 31947
rect 18135 31926 18142 31947
rect 18194 31926 18211 31947
rect 18211 31926 18228 31947
rect 18280 31926 18287 31947
rect 18287 31926 18314 31947
rect 18366 31926 18400 31960
rect 18022 31879 18056 31888
rect 18108 31879 18142 31888
rect 18194 31879 18228 31888
rect 18280 31879 18314 31888
rect 18022 31854 18025 31879
rect 18025 31854 18056 31879
rect 18108 31854 18135 31879
rect 18135 31854 18142 31879
rect 18194 31854 18211 31879
rect 18211 31854 18228 31879
rect 18280 31854 18287 31879
rect 18287 31854 18314 31879
rect 18366 31854 18400 31888
rect 18022 31811 18056 31816
rect 18108 31811 18142 31816
rect 18194 31811 18228 31816
rect 18280 31811 18314 31816
rect 18022 31782 18025 31811
rect 18025 31782 18056 31811
rect 18108 31782 18135 31811
rect 18135 31782 18142 31811
rect 18194 31782 18211 31811
rect 18211 31782 18228 31811
rect 18280 31782 18287 31811
rect 18287 31782 18314 31811
rect 18366 31782 18400 31816
rect 18022 31743 18056 31744
rect 18108 31743 18142 31744
rect 18194 31743 18228 31744
rect 18280 31743 18314 31744
rect 18022 31710 18025 31743
rect 18025 31710 18056 31743
rect 18108 31710 18135 31743
rect 18135 31710 18142 31743
rect 18194 31710 18211 31743
rect 18211 31710 18228 31743
rect 18280 31710 18287 31743
rect 18287 31710 18314 31743
rect 18366 31710 18400 31744
rect 218 31670 252 31704
rect 218 31598 252 31632
rect 218 31526 252 31560
rect 218 31454 252 31488
rect 218 31382 252 31416
rect 218 31310 252 31344
rect 218 31238 252 31272
rect 218 31166 252 31200
rect 218 31094 252 31128
rect 218 31022 252 31056
rect 218 30950 252 30984
rect 218 30878 252 30912
rect 218 30806 252 30840
rect 218 30734 252 30768
rect 218 30662 252 30696
rect 218 30590 252 30624
rect 218 30518 252 30552
rect 218 30446 252 30480
rect 218 30374 252 30408
rect 218 30302 252 30336
rect 218 30230 252 30264
rect 218 30158 252 30192
rect 218 30086 252 30120
rect 218 30014 252 30048
rect 218 29942 252 29976
rect 218 29870 252 29904
rect 218 29798 252 29832
rect 218 29726 252 29760
rect 218 29654 252 29688
rect 218 29582 252 29616
rect 218 29510 252 29544
rect 218 29438 252 29472
rect 218 29366 252 29400
rect 218 29294 252 29328
rect 218 29222 252 29256
rect 218 29150 252 29184
rect 218 29078 252 29112
rect 218 29006 252 29040
rect 218 28934 252 28968
rect 218 28862 252 28896
rect 218 28790 252 28824
rect 218 28718 252 28752
rect 218 28646 252 28680
rect 218 28574 252 28608
rect 218 28501 252 28535
rect 218 28428 252 28462
rect 218 28355 252 28389
rect 218 28282 252 28316
rect 218 28209 252 28243
rect 218 28136 252 28170
rect 218 28063 252 28097
rect 218 27990 252 28024
rect 218 27917 252 27951
rect 218 27844 252 27878
rect 218 27771 252 27805
rect 218 27698 252 27732
rect 218 27625 252 27659
rect 218 27552 252 27586
rect 218 27479 252 27513
rect 218 27406 252 27440
rect 218 27333 252 27367
rect 218 27260 252 27294
rect 218 27187 252 27221
rect 218 27114 252 27148
rect 218 27041 252 27075
rect 218 26968 252 27002
rect 218 26895 252 26929
rect 218 26822 252 26856
rect 218 26749 252 26783
rect 218 26676 252 26710
rect 218 26603 252 26637
rect 218 26530 252 26564
rect 218 26457 252 26491
rect 218 26384 252 26418
rect 218 26311 252 26345
rect 218 26238 252 26272
rect 218 26165 252 26199
rect 218 26092 252 26126
rect 218 26019 252 26053
rect 218 25946 252 25980
rect 218 25873 252 25907
rect 218 25800 252 25834
rect 218 25727 252 25761
rect 218 25654 252 25688
rect 218 25581 252 25615
rect 218 25508 252 25542
rect 218 25435 252 25469
rect 218 25362 252 25396
rect 218 25289 252 25323
rect 218 25216 252 25250
rect 218 25143 252 25177
rect 218 25070 252 25104
rect 218 24997 252 25031
rect 218 24924 252 24958
rect 218 24851 252 24885
rect 218 24778 252 24812
rect 218 24705 252 24739
rect 218 24632 252 24666
rect 218 24559 252 24593
rect 218 24486 252 24520
rect 218 24413 252 24447
rect 218 24340 252 24374
rect 218 24267 252 24301
rect 218 24194 252 24228
rect 218 24121 252 24155
rect 218 24048 252 24082
rect 218 23975 252 24009
rect 218 23902 252 23936
rect 218 23829 252 23863
rect 18022 31641 18025 31672
rect 18025 31641 18056 31672
rect 18108 31641 18135 31672
rect 18135 31641 18142 31672
rect 18194 31641 18211 31672
rect 18211 31641 18228 31672
rect 18280 31641 18287 31672
rect 18287 31641 18314 31672
rect 18022 31638 18056 31641
rect 18108 31638 18142 31641
rect 18194 31638 18228 31641
rect 18280 31638 18314 31641
rect 18366 31638 18400 31672
rect 18022 31573 18025 31600
rect 18025 31573 18056 31600
rect 18108 31573 18135 31600
rect 18135 31573 18142 31600
rect 18194 31573 18211 31600
rect 18211 31573 18228 31600
rect 18280 31573 18287 31600
rect 18287 31573 18314 31600
rect 18022 31566 18056 31573
rect 18108 31566 18142 31573
rect 18194 31566 18228 31573
rect 18280 31566 18314 31573
rect 18366 31566 18400 31600
rect 18022 31505 18025 31528
rect 18025 31505 18056 31528
rect 18108 31505 18135 31528
rect 18135 31505 18142 31528
rect 18194 31505 18211 31528
rect 18211 31505 18228 31528
rect 18280 31505 18287 31528
rect 18287 31505 18314 31528
rect 18022 31494 18056 31505
rect 18108 31494 18142 31505
rect 18194 31494 18228 31505
rect 18280 31494 18314 31505
rect 18366 31494 18400 31528
rect 18022 31437 18025 31456
rect 18025 31437 18056 31456
rect 18108 31437 18135 31456
rect 18135 31437 18142 31456
rect 18194 31437 18211 31456
rect 18211 31437 18228 31456
rect 18280 31437 18287 31456
rect 18287 31437 18314 31456
rect 18022 31422 18056 31437
rect 18108 31422 18142 31437
rect 18194 31422 18228 31437
rect 18280 31422 18314 31437
rect 18366 31422 18400 31456
rect 18022 31369 18025 31384
rect 18025 31369 18056 31384
rect 18108 31369 18135 31384
rect 18135 31369 18142 31384
rect 18194 31369 18211 31384
rect 18211 31369 18228 31384
rect 18280 31369 18287 31384
rect 18287 31369 18314 31384
rect 18022 31350 18056 31369
rect 18108 31350 18142 31369
rect 18194 31350 18228 31369
rect 18280 31350 18314 31369
rect 18366 31350 18400 31384
rect 18022 31301 18025 31312
rect 18025 31301 18056 31312
rect 18108 31301 18135 31312
rect 18135 31301 18142 31312
rect 18194 31301 18211 31312
rect 18211 31301 18228 31312
rect 18280 31301 18287 31312
rect 18287 31301 18314 31312
rect 18022 31278 18056 31301
rect 18108 31278 18142 31301
rect 18194 31278 18228 31301
rect 18280 31278 18314 31301
rect 18366 31278 18400 31312
rect 18022 31233 18025 31240
rect 18025 31233 18056 31240
rect 18108 31233 18135 31240
rect 18135 31233 18142 31240
rect 18194 31233 18211 31240
rect 18211 31233 18228 31240
rect 18280 31233 18287 31240
rect 18287 31233 18314 31240
rect 18022 31206 18056 31233
rect 18108 31206 18142 31233
rect 18194 31206 18228 31233
rect 18280 31206 18314 31233
rect 18366 31206 18400 31240
rect 18022 31165 18025 31168
rect 18025 31165 18056 31168
rect 18108 31165 18135 31168
rect 18135 31165 18142 31168
rect 18194 31165 18211 31168
rect 18211 31165 18228 31168
rect 18280 31165 18287 31168
rect 18287 31165 18314 31168
rect 18022 31134 18056 31165
rect 18108 31134 18142 31165
rect 18194 31134 18228 31165
rect 18280 31134 18314 31165
rect 18366 31134 18400 31168
rect 18022 31063 18056 31096
rect 18108 31063 18142 31096
rect 18194 31063 18228 31096
rect 18280 31063 18314 31096
rect 18022 31062 18025 31063
rect 18025 31062 18056 31063
rect 18108 31062 18135 31063
rect 18135 31062 18142 31063
rect 18194 31062 18211 31063
rect 18211 31062 18228 31063
rect 18280 31062 18287 31063
rect 18287 31062 18314 31063
rect 18366 31062 18400 31096
rect 18022 30995 18056 31024
rect 18108 30995 18142 31024
rect 18194 30995 18228 31024
rect 18280 30995 18314 31024
rect 18022 30990 18025 30995
rect 18025 30990 18056 30995
rect 18108 30990 18135 30995
rect 18135 30990 18142 30995
rect 18194 30990 18211 30995
rect 18211 30990 18228 30995
rect 18280 30990 18287 30995
rect 18287 30990 18314 30995
rect 18366 30990 18400 31024
rect 18022 30927 18056 30952
rect 18108 30927 18142 30952
rect 18194 30927 18228 30952
rect 18280 30927 18314 30952
rect 18022 30918 18025 30927
rect 18025 30918 18056 30927
rect 18108 30918 18135 30927
rect 18135 30918 18142 30927
rect 18194 30918 18211 30927
rect 18211 30918 18228 30927
rect 18280 30918 18287 30927
rect 18287 30918 18314 30927
rect 18366 30918 18400 30952
rect 18022 30859 18056 30880
rect 18108 30859 18142 30880
rect 18194 30859 18228 30880
rect 18280 30859 18314 30880
rect 18022 30846 18025 30859
rect 18025 30846 18056 30859
rect 18108 30846 18135 30859
rect 18135 30846 18142 30859
rect 18194 30846 18211 30859
rect 18211 30846 18228 30859
rect 18280 30846 18287 30859
rect 18287 30846 18314 30859
rect 18366 30846 18400 30880
rect 18022 30791 18056 30808
rect 18108 30791 18142 30808
rect 18194 30791 18228 30808
rect 18280 30791 18314 30808
rect 18022 30774 18025 30791
rect 18025 30774 18056 30791
rect 18108 30774 18135 30791
rect 18135 30774 18142 30791
rect 18194 30774 18211 30791
rect 18211 30774 18228 30791
rect 18280 30774 18287 30791
rect 18287 30774 18314 30791
rect 18366 30774 18400 30808
rect 18022 30723 18056 30736
rect 18108 30723 18142 30736
rect 18194 30723 18228 30736
rect 18280 30723 18314 30736
rect 18022 30702 18025 30723
rect 18025 30702 18056 30723
rect 18108 30702 18135 30723
rect 18135 30702 18142 30723
rect 18194 30702 18211 30723
rect 18211 30702 18228 30723
rect 18280 30702 18287 30723
rect 18287 30702 18314 30723
rect 18366 30702 18400 30736
rect 22829 33312 22863 33335
rect 22911 33312 22945 33335
rect 22993 33312 23027 33335
rect 23075 33312 23109 33335
rect 23157 33312 23191 33335
rect 23239 33312 23273 33335
rect 22829 33267 22861 33273
rect 22861 33267 22863 33273
rect 22911 33267 22931 33273
rect 22931 33267 22945 33273
rect 22993 33267 23001 33273
rect 23001 33267 23027 33273
rect 23075 33267 23107 33273
rect 23107 33267 23109 33273
rect 23157 33267 23177 33273
rect 23177 33267 23191 33273
rect 23239 33267 23247 33273
rect 23247 33267 23273 33273
rect 22829 33239 22863 33267
rect 22911 33239 22945 33267
rect 22993 33239 23027 33267
rect 23075 33239 23109 33267
rect 23157 33239 23191 33267
rect 23239 33239 23273 33267
rect 22829 33199 22861 33200
rect 22861 33199 22863 33200
rect 22911 33199 22931 33200
rect 22931 33199 22945 33200
rect 22993 33199 23001 33200
rect 23001 33199 23027 33200
rect 23075 33199 23107 33200
rect 23107 33199 23109 33200
rect 23157 33199 23177 33200
rect 23177 33199 23191 33200
rect 23239 33199 23247 33200
rect 23247 33199 23273 33200
rect 22829 33166 22863 33199
rect 22911 33166 22945 33199
rect 22993 33166 23027 33199
rect 23075 33166 23109 33199
rect 23157 33166 23191 33199
rect 23239 33166 23273 33199
rect 22829 33097 22863 33127
rect 22911 33097 22945 33127
rect 22993 33097 23027 33127
rect 23075 33097 23109 33127
rect 23157 33097 23191 33127
rect 23239 33097 23273 33127
rect 22829 33093 22861 33097
rect 22861 33093 22863 33097
rect 22911 33093 22931 33097
rect 22931 33093 22945 33097
rect 22993 33093 23001 33097
rect 23001 33093 23027 33097
rect 23075 33093 23107 33097
rect 23107 33093 23109 33097
rect 23157 33093 23177 33097
rect 23177 33093 23191 33097
rect 23239 33093 23247 33097
rect 23247 33093 23273 33097
rect 22829 33029 22863 33054
rect 22911 33029 22945 33054
rect 22993 33029 23027 33054
rect 23075 33029 23109 33054
rect 23157 33029 23191 33054
rect 23239 33029 23273 33054
rect 22829 33020 22861 33029
rect 22861 33020 22863 33029
rect 22911 33020 22931 33029
rect 22931 33020 22945 33029
rect 22993 33020 23001 33029
rect 23001 33020 23027 33029
rect 23075 33020 23107 33029
rect 23107 33020 23109 33029
rect 23157 33020 23177 33029
rect 23177 33020 23191 33029
rect 23239 33020 23247 33029
rect 23247 33020 23273 33029
rect 22829 32961 22863 32981
rect 22911 32961 22945 32981
rect 22993 32961 23027 32981
rect 23075 32961 23109 32981
rect 23157 32961 23191 32981
rect 23239 32961 23273 32981
rect 22829 32947 22861 32961
rect 22861 32947 22863 32961
rect 22911 32947 22931 32961
rect 22931 32947 22945 32961
rect 22993 32947 23001 32961
rect 23001 32947 23027 32961
rect 23075 32947 23107 32961
rect 23107 32947 23109 32961
rect 23157 32947 23177 32961
rect 23177 32947 23191 32961
rect 23239 32947 23247 32961
rect 23247 32947 23273 32961
rect 22829 32893 22863 32908
rect 22911 32893 22945 32908
rect 22993 32893 23027 32908
rect 23075 32893 23109 32908
rect 23157 32893 23191 32908
rect 23239 32893 23273 32908
rect 22829 32874 22861 32893
rect 22861 32874 22863 32893
rect 22911 32874 22931 32893
rect 22931 32874 22945 32893
rect 22993 32874 23001 32893
rect 23001 32874 23027 32893
rect 23075 32874 23107 32893
rect 23107 32874 23109 32893
rect 23157 32874 23177 32893
rect 23177 32874 23191 32893
rect 23239 32874 23247 32893
rect 23247 32874 23273 32893
rect 22829 32825 22863 32835
rect 22911 32825 22945 32835
rect 22993 32825 23027 32835
rect 23075 32825 23109 32835
rect 23157 32825 23191 32835
rect 23239 32825 23273 32835
rect 22829 32801 22861 32825
rect 22861 32801 22863 32825
rect 22911 32801 22931 32825
rect 22931 32801 22945 32825
rect 22993 32801 23001 32825
rect 23001 32801 23027 32825
rect 23075 32801 23107 32825
rect 23107 32801 23109 32825
rect 23157 32801 23177 32825
rect 23177 32801 23191 32825
rect 23239 32801 23247 32825
rect 23247 32801 23273 32825
rect 22829 32757 22863 32762
rect 22911 32757 22945 32762
rect 22993 32757 23027 32762
rect 23075 32757 23109 32762
rect 23157 32757 23191 32762
rect 23239 32757 23273 32762
rect 22829 32728 22861 32757
rect 22861 32728 22863 32757
rect 22911 32728 22931 32757
rect 22931 32728 22945 32757
rect 22993 32728 23001 32757
rect 23001 32728 23027 32757
rect 23075 32728 23107 32757
rect 23107 32728 23109 32757
rect 23157 32728 23177 32757
rect 23177 32728 23191 32757
rect 23239 32728 23247 32757
rect 23247 32728 23273 32757
rect 22829 32655 22861 32689
rect 22861 32655 22863 32689
rect 22911 32655 22931 32689
rect 22931 32655 22945 32689
rect 22993 32655 23001 32689
rect 23001 32655 23027 32689
rect 23075 32655 23107 32689
rect 23107 32655 23109 32689
rect 23157 32655 23177 32689
rect 23177 32655 23191 32689
rect 23239 32655 23247 32689
rect 23247 32655 23273 32689
rect 22829 32587 22861 32616
rect 22861 32587 22863 32616
rect 22911 32587 22931 32616
rect 22931 32587 22945 32616
rect 22993 32587 23001 32616
rect 23001 32587 23027 32616
rect 23075 32587 23107 32616
rect 23107 32587 23109 32616
rect 23157 32587 23177 32616
rect 23177 32587 23191 32616
rect 23239 32587 23247 32616
rect 23247 32587 23273 32616
rect 22829 32582 22863 32587
rect 22911 32582 22945 32587
rect 22993 32582 23027 32587
rect 23075 32582 23109 32587
rect 23157 32582 23191 32587
rect 23239 32582 23273 32587
rect 22829 32519 22861 32543
rect 22861 32519 22863 32543
rect 22911 32519 22931 32543
rect 22931 32519 22945 32543
rect 22993 32519 23001 32543
rect 23001 32519 23027 32543
rect 23075 32519 23107 32543
rect 23107 32519 23109 32543
rect 23157 32519 23177 32543
rect 23177 32519 23191 32543
rect 23239 32519 23247 32543
rect 23247 32519 23273 32543
rect 22829 32509 22863 32519
rect 22911 32509 22945 32519
rect 22993 32509 23027 32519
rect 23075 32509 23109 32519
rect 23157 32509 23191 32519
rect 23239 32509 23273 32519
rect 22829 32451 22861 32470
rect 22861 32451 22863 32470
rect 22911 32451 22931 32470
rect 22931 32451 22945 32470
rect 22993 32451 23001 32470
rect 23001 32451 23027 32470
rect 23075 32451 23107 32470
rect 23107 32451 23109 32470
rect 23157 32451 23177 32470
rect 23177 32451 23191 32470
rect 23239 32451 23247 32470
rect 23247 32451 23273 32470
rect 22829 32436 22863 32451
rect 22911 32436 22945 32451
rect 22993 32436 23027 32451
rect 23075 32436 23109 32451
rect 23157 32436 23191 32451
rect 23239 32436 23273 32451
rect 22829 32383 22861 32397
rect 22861 32383 22863 32397
rect 22911 32383 22931 32397
rect 22931 32383 22945 32397
rect 22993 32383 23001 32397
rect 23001 32383 23027 32397
rect 23075 32383 23107 32397
rect 23107 32383 23109 32397
rect 23157 32383 23177 32397
rect 23177 32383 23191 32397
rect 23239 32383 23247 32397
rect 23247 32383 23273 32397
rect 22829 32363 22863 32383
rect 22911 32363 22945 32383
rect 22993 32363 23027 32383
rect 23075 32363 23109 32383
rect 23157 32363 23191 32383
rect 23239 32363 23273 32383
rect 22829 32315 22861 32324
rect 22861 32315 22863 32324
rect 22911 32315 22931 32324
rect 22931 32315 22945 32324
rect 22993 32315 23001 32324
rect 23001 32315 23027 32324
rect 23075 32315 23107 32324
rect 23107 32315 23109 32324
rect 23157 32315 23177 32324
rect 23177 32315 23191 32324
rect 23239 32315 23247 32324
rect 23247 32315 23273 32324
rect 22829 32290 22863 32315
rect 22911 32290 22945 32315
rect 22993 32290 23027 32315
rect 23075 32290 23109 32315
rect 23157 32290 23191 32315
rect 23239 32290 23273 32315
rect 22829 32247 22861 32251
rect 22861 32247 22863 32251
rect 22911 32247 22931 32251
rect 22931 32247 22945 32251
rect 22993 32247 23001 32251
rect 23001 32247 23027 32251
rect 23075 32247 23107 32251
rect 23107 32247 23109 32251
rect 23157 32247 23177 32251
rect 23177 32247 23191 32251
rect 23239 32247 23247 32251
rect 23247 32247 23273 32251
rect 22829 32217 22863 32247
rect 22911 32217 22945 32247
rect 22993 32217 23027 32247
rect 23075 32217 23109 32247
rect 23157 32217 23191 32247
rect 23239 32217 23273 32247
rect 22829 32145 22863 32178
rect 22911 32145 22945 32178
rect 22993 32145 23027 32178
rect 23075 32145 23109 32178
rect 23157 32145 23191 32178
rect 23239 32145 23273 32178
rect 22829 32144 22861 32145
rect 22861 32144 22863 32145
rect 22911 32144 22931 32145
rect 22931 32144 22945 32145
rect 22993 32144 23001 32145
rect 23001 32144 23027 32145
rect 23075 32144 23107 32145
rect 23107 32144 23109 32145
rect 23157 32144 23177 32145
rect 23177 32144 23191 32145
rect 23239 32144 23247 32145
rect 23247 32144 23273 32145
rect 22829 32077 22863 32105
rect 22911 32077 22945 32105
rect 22993 32077 23027 32105
rect 23075 32077 23109 32105
rect 23157 32077 23191 32105
rect 23239 32077 23273 32105
rect 22829 32071 22861 32077
rect 22861 32071 22863 32077
rect 22911 32071 22931 32077
rect 22931 32071 22945 32077
rect 22993 32071 23001 32077
rect 23001 32071 23027 32077
rect 23075 32071 23107 32077
rect 23107 32071 23109 32077
rect 23157 32071 23177 32077
rect 23177 32071 23191 32077
rect 23239 32071 23247 32077
rect 23247 32071 23273 32077
rect 22829 32009 22863 32032
rect 22911 32009 22945 32032
rect 22993 32009 23027 32032
rect 23075 32009 23109 32032
rect 23157 32009 23191 32032
rect 23239 32009 23273 32032
rect 22829 31998 22861 32009
rect 22861 31998 22863 32009
rect 22911 31998 22931 32009
rect 22931 31998 22945 32009
rect 22993 31998 23001 32009
rect 23001 31998 23027 32009
rect 23075 31998 23107 32009
rect 23107 31998 23109 32009
rect 23157 31998 23177 32009
rect 23177 31998 23191 32009
rect 23239 31998 23247 32009
rect 23247 31998 23273 32009
rect 22829 31941 22863 31959
rect 22911 31941 22945 31959
rect 22993 31941 23027 31959
rect 23075 31941 23109 31959
rect 23157 31941 23191 31959
rect 23239 31941 23273 31959
rect 22829 31925 22861 31941
rect 22861 31925 22863 31941
rect 22911 31925 22931 31941
rect 22931 31925 22945 31941
rect 22993 31925 23001 31941
rect 23001 31925 23027 31941
rect 23075 31925 23107 31941
rect 23107 31925 23109 31941
rect 23157 31925 23177 31941
rect 23177 31925 23191 31941
rect 23239 31925 23247 31941
rect 23247 31925 23273 31941
rect 22829 31873 22863 31886
rect 22911 31873 22945 31886
rect 22993 31873 23027 31886
rect 23075 31873 23109 31886
rect 23157 31873 23191 31886
rect 23239 31873 23273 31886
rect 22829 31852 22861 31873
rect 22861 31852 22863 31873
rect 22911 31852 22931 31873
rect 22931 31852 22945 31873
rect 22993 31852 23001 31873
rect 23001 31852 23027 31873
rect 23075 31852 23107 31873
rect 23107 31852 23109 31873
rect 23157 31852 23177 31873
rect 23177 31852 23191 31873
rect 23239 31852 23247 31873
rect 23247 31852 23273 31873
rect 22829 31805 22863 31813
rect 22911 31805 22945 31813
rect 22993 31805 23027 31813
rect 23075 31805 23109 31813
rect 23157 31805 23191 31813
rect 23239 31805 23273 31813
rect 22829 31779 22861 31805
rect 22861 31779 22863 31805
rect 22911 31779 22931 31805
rect 22931 31779 22945 31805
rect 22993 31779 23001 31805
rect 23001 31779 23027 31805
rect 23075 31779 23107 31805
rect 23107 31779 23109 31805
rect 23157 31779 23177 31805
rect 23177 31779 23191 31805
rect 23239 31779 23247 31805
rect 23247 31779 23273 31805
rect 22829 31737 22863 31740
rect 22911 31737 22945 31740
rect 22993 31737 23027 31740
rect 23075 31737 23109 31740
rect 23157 31737 23191 31740
rect 23239 31737 23273 31740
rect 22829 31706 22861 31737
rect 22861 31706 22863 31737
rect 22911 31706 22931 31737
rect 22931 31706 22945 31737
rect 22993 31706 23001 31737
rect 23001 31706 23027 31737
rect 23075 31706 23107 31737
rect 23107 31706 23109 31737
rect 23157 31706 23177 31737
rect 23177 31706 23191 31737
rect 23239 31706 23247 31737
rect 23247 31706 23273 31737
rect 22830 31635 22861 31642
rect 22861 31635 22864 31642
rect 22830 31608 22864 31635
rect 22932 31608 22966 31642
rect 23034 31635 23037 31642
rect 23037 31635 23068 31642
rect 23034 31608 23068 31635
rect 22830 31567 22861 31568
rect 22861 31567 22864 31568
rect 22830 31534 22864 31567
rect 22932 31534 22966 31568
rect 23034 31567 23037 31568
rect 23037 31567 23068 31568
rect 23034 31534 23068 31567
rect 22830 31465 22864 31494
rect 22830 31460 22861 31465
rect 22861 31460 22864 31465
rect 22932 31460 22966 31494
rect 23034 31465 23068 31494
rect 23034 31460 23037 31465
rect 23037 31460 23068 31465
rect 22830 31397 22864 31420
rect 22830 31386 22861 31397
rect 22861 31386 22864 31397
rect 22932 31386 22966 31420
rect 23034 31397 23068 31420
rect 23034 31386 23037 31397
rect 23037 31386 23068 31397
rect 22830 31329 22864 31346
rect 22830 31312 22861 31329
rect 22861 31312 22864 31329
rect 22932 31312 22966 31346
rect 23034 31329 23068 31346
rect 23034 31312 23037 31329
rect 23037 31312 23068 31329
rect 22830 31261 22864 31271
rect 22830 31237 22861 31261
rect 22861 31237 22864 31261
rect 22932 31237 22966 31271
rect 23034 31261 23068 31271
rect 23034 31237 23037 31261
rect 23037 31237 23068 31261
rect 22830 31193 22864 31196
rect 22830 31162 22861 31193
rect 22861 31162 22864 31193
rect 22932 31162 22966 31196
rect 23034 31193 23068 31196
rect 23034 31162 23037 31193
rect 23037 31162 23068 31193
rect 22830 31091 22861 31121
rect 22861 31091 22864 31121
rect 22830 31087 22864 31091
rect 22932 31087 22966 31121
rect 23034 31091 23037 31121
rect 23037 31091 23068 31121
rect 23034 31087 23068 31091
rect 22830 31023 22861 31046
rect 22861 31023 22864 31046
rect 22830 31012 22864 31023
rect 22932 31012 22966 31046
rect 23034 31023 23037 31046
rect 23037 31023 23068 31046
rect 23034 31012 23068 31023
rect 22830 30955 22861 30971
rect 22861 30955 22864 30971
rect 22830 30937 22864 30955
rect 22932 30937 22966 30971
rect 23034 30955 23037 30971
rect 23037 30955 23068 30971
rect 23034 30937 23068 30955
rect 22830 30887 22861 30896
rect 22861 30887 22864 30896
rect 22830 30862 22864 30887
rect 22932 30862 22966 30896
rect 23034 30887 23037 30896
rect 23037 30887 23068 30896
rect 23034 30862 23068 30887
rect 22830 30819 22861 30821
rect 22861 30819 22864 30821
rect 22830 30787 22864 30819
rect 22932 30787 22966 30821
rect 23034 30819 23037 30821
rect 23037 30819 23068 30821
rect 23034 30787 23068 30819
rect 22830 30717 22864 30746
rect 18022 30655 18056 30664
rect 18108 30655 18142 30664
rect 18194 30655 18228 30664
rect 18280 30655 18314 30664
rect 18022 30630 18025 30655
rect 18025 30630 18056 30655
rect 18108 30630 18135 30655
rect 18135 30630 18142 30655
rect 18194 30630 18211 30655
rect 18211 30630 18228 30655
rect 18280 30630 18287 30655
rect 18287 30630 18314 30655
rect 18366 30630 18400 30664
rect 18022 30587 18056 30592
rect 18108 30587 18142 30592
rect 18194 30587 18228 30592
rect 18280 30587 18314 30592
rect 18022 30558 18025 30587
rect 18025 30558 18056 30587
rect 18108 30558 18135 30587
rect 18135 30558 18142 30587
rect 18194 30558 18211 30587
rect 18211 30558 18228 30587
rect 18280 30558 18287 30587
rect 18287 30558 18314 30587
rect 18366 30558 18400 30592
rect 18022 30519 18056 30520
rect 18108 30519 18142 30520
rect 18194 30519 18228 30520
rect 18280 30519 18314 30520
rect 18022 30486 18025 30519
rect 18025 30486 18056 30519
rect 18108 30486 18135 30519
rect 18135 30486 18142 30519
rect 18194 30486 18211 30519
rect 18211 30486 18228 30519
rect 18280 30486 18287 30519
rect 18287 30486 18314 30519
rect 18366 30486 18400 30520
rect 18022 30417 18025 30448
rect 18025 30417 18056 30448
rect 18108 30417 18135 30448
rect 18135 30417 18142 30448
rect 18194 30417 18211 30448
rect 18211 30417 18228 30448
rect 18280 30417 18287 30448
rect 18287 30417 18314 30448
rect 18022 30414 18056 30417
rect 18108 30414 18142 30417
rect 18194 30414 18228 30417
rect 18280 30414 18314 30417
rect 18366 30414 18400 30448
rect 18022 30349 18025 30376
rect 18025 30349 18056 30376
rect 18108 30349 18135 30376
rect 18135 30349 18142 30376
rect 18194 30349 18211 30376
rect 18211 30349 18228 30376
rect 18280 30349 18287 30376
rect 18287 30349 18314 30376
rect 18022 30342 18056 30349
rect 18108 30342 18142 30349
rect 18194 30342 18228 30349
rect 18280 30342 18314 30349
rect 18366 30342 18400 30376
rect 18022 30281 18025 30304
rect 18025 30281 18056 30304
rect 18108 30281 18135 30304
rect 18135 30281 18142 30304
rect 18194 30281 18211 30304
rect 18211 30281 18228 30304
rect 18280 30281 18287 30304
rect 18287 30281 18314 30304
rect 18022 30270 18056 30281
rect 18108 30270 18142 30281
rect 18194 30270 18228 30281
rect 18280 30270 18314 30281
rect 18366 30270 18400 30304
rect 18022 30213 18025 30232
rect 18025 30213 18056 30232
rect 18108 30213 18135 30232
rect 18135 30213 18142 30232
rect 18194 30213 18211 30232
rect 18211 30213 18228 30232
rect 18280 30213 18287 30232
rect 18287 30213 18314 30232
rect 18022 30198 18056 30213
rect 18108 30198 18142 30213
rect 18194 30198 18228 30213
rect 18280 30198 18314 30213
rect 18366 30198 18400 30232
rect 18022 30145 18025 30160
rect 18025 30145 18056 30160
rect 18108 30145 18135 30160
rect 18135 30145 18142 30160
rect 18194 30145 18211 30160
rect 18211 30145 18228 30160
rect 18280 30145 18287 30160
rect 18287 30145 18314 30160
rect 18022 30126 18056 30145
rect 18108 30126 18142 30145
rect 18194 30126 18228 30145
rect 18280 30126 18314 30145
rect 18366 30126 18400 30160
rect 18022 30077 18025 30088
rect 18025 30077 18056 30088
rect 18108 30077 18135 30088
rect 18135 30077 18142 30088
rect 18194 30077 18211 30088
rect 18211 30077 18228 30088
rect 18280 30077 18287 30088
rect 18287 30077 18314 30088
rect 18022 30054 18056 30077
rect 18108 30054 18142 30077
rect 18194 30054 18228 30077
rect 18280 30054 18314 30077
rect 18366 30054 18400 30088
rect 18022 30009 18025 30016
rect 18025 30009 18056 30016
rect 18108 30009 18135 30016
rect 18135 30009 18142 30016
rect 18194 30009 18211 30016
rect 18211 30009 18228 30016
rect 18280 30009 18287 30016
rect 18287 30009 18314 30016
rect 18022 29982 18056 30009
rect 18108 29982 18142 30009
rect 18194 29982 18228 30009
rect 18280 29982 18314 30009
rect 18366 29982 18400 30016
rect 18022 29941 18025 29944
rect 18025 29941 18056 29944
rect 18108 29941 18135 29944
rect 18135 29941 18142 29944
rect 18194 29941 18211 29944
rect 18211 29941 18228 29944
rect 18280 29941 18287 29944
rect 18287 29941 18314 29944
rect 18022 29910 18056 29941
rect 18108 29910 18142 29941
rect 18194 29910 18228 29941
rect 18280 29910 18314 29941
rect 18366 29910 18400 29944
rect 18022 29839 18056 29872
rect 18108 29839 18142 29872
rect 18194 29839 18228 29872
rect 18280 29839 18314 29872
rect 18022 29838 18025 29839
rect 18025 29838 18056 29839
rect 18108 29838 18135 29839
rect 18135 29838 18142 29839
rect 18194 29838 18211 29839
rect 18211 29838 18228 29839
rect 18280 29838 18287 29839
rect 18287 29838 18314 29839
rect 18366 29838 18400 29872
rect 18022 29771 18056 29800
rect 18108 29771 18142 29800
rect 18194 29771 18228 29800
rect 18280 29771 18314 29800
rect 18022 29766 18025 29771
rect 18025 29766 18056 29771
rect 18108 29766 18135 29771
rect 18135 29766 18142 29771
rect 18194 29766 18211 29771
rect 18211 29766 18228 29771
rect 18280 29766 18287 29771
rect 18287 29766 18314 29771
rect 18366 29766 18400 29800
rect 18022 29703 18056 29728
rect 18108 29703 18142 29728
rect 18194 29703 18228 29728
rect 18280 29703 18314 29728
rect 18022 29694 18025 29703
rect 18025 29694 18056 29703
rect 18108 29694 18135 29703
rect 18135 29694 18142 29703
rect 18194 29694 18211 29703
rect 18211 29694 18228 29703
rect 18280 29694 18287 29703
rect 18287 29694 18314 29703
rect 18366 29694 18400 29728
rect 18022 29635 18056 29656
rect 18108 29635 18142 29656
rect 18194 29635 18228 29656
rect 18280 29635 18314 29656
rect 18022 29622 18025 29635
rect 18025 29622 18056 29635
rect 18108 29622 18135 29635
rect 18135 29622 18142 29635
rect 18194 29622 18211 29635
rect 18211 29622 18228 29635
rect 18280 29622 18287 29635
rect 18287 29622 18314 29635
rect 18366 29622 18400 29656
rect 18022 29567 18056 29584
rect 18108 29567 18142 29584
rect 18194 29567 18228 29584
rect 18280 29567 18314 29584
rect 18022 29550 18025 29567
rect 18025 29550 18056 29567
rect 18108 29550 18135 29567
rect 18135 29550 18142 29567
rect 18194 29550 18211 29567
rect 18211 29550 18228 29567
rect 18280 29550 18287 29567
rect 18287 29550 18314 29567
rect 18366 29550 18400 29584
rect 18022 29499 18056 29512
rect 18108 29499 18142 29512
rect 18194 29499 18228 29512
rect 18280 29499 18314 29512
rect 18022 29478 18025 29499
rect 18025 29478 18056 29499
rect 18108 29478 18135 29499
rect 18135 29478 18142 29499
rect 18194 29478 18211 29499
rect 18211 29478 18228 29499
rect 18280 29478 18287 29499
rect 18287 29478 18314 29499
rect 18366 29478 18400 29512
rect 18022 29431 18056 29440
rect 18108 29431 18142 29440
rect 18194 29431 18228 29440
rect 18280 29431 18314 29440
rect 18022 29406 18025 29431
rect 18025 29406 18056 29431
rect 18108 29406 18135 29431
rect 18135 29406 18142 29431
rect 18194 29406 18211 29431
rect 18211 29406 18228 29431
rect 18280 29406 18287 29431
rect 18287 29406 18314 29431
rect 18366 29406 18400 29440
rect 18022 29363 18056 29368
rect 18108 29363 18142 29368
rect 18194 29363 18228 29368
rect 18280 29363 18314 29368
rect 18022 29334 18025 29363
rect 18025 29334 18056 29363
rect 18108 29334 18135 29363
rect 18135 29334 18142 29363
rect 18194 29334 18211 29363
rect 18211 29334 18228 29363
rect 18280 29334 18287 29363
rect 18287 29334 18314 29363
rect 18366 29334 18400 29368
rect 18022 29295 18056 29296
rect 18108 29295 18142 29296
rect 18194 29295 18228 29296
rect 18280 29295 18314 29296
rect 18022 29262 18025 29295
rect 18025 29262 18056 29295
rect 18108 29262 18135 29295
rect 18135 29262 18142 29295
rect 18194 29262 18211 29295
rect 18211 29262 18228 29295
rect 18280 29262 18287 29295
rect 18287 29262 18314 29295
rect 18366 29262 18400 29296
rect 18022 29193 18025 29224
rect 18025 29193 18056 29224
rect 18108 29193 18135 29224
rect 18135 29193 18142 29224
rect 18194 29193 18211 29224
rect 18211 29193 18228 29224
rect 18280 29193 18287 29224
rect 18287 29193 18314 29224
rect 18022 29190 18056 29193
rect 18108 29190 18142 29193
rect 18194 29190 18228 29193
rect 18280 29190 18314 29193
rect 18366 29190 18400 29224
rect 18022 29125 18025 29152
rect 18025 29125 18056 29152
rect 18108 29125 18135 29152
rect 18135 29125 18142 29152
rect 18194 29125 18211 29152
rect 18211 29125 18228 29152
rect 18280 29125 18287 29152
rect 18287 29125 18314 29152
rect 18022 29118 18056 29125
rect 18108 29118 18142 29125
rect 18194 29118 18228 29125
rect 18280 29118 18314 29125
rect 18366 29118 18400 29152
rect 18022 29057 18025 29080
rect 18025 29057 18056 29080
rect 18108 29057 18135 29080
rect 18135 29057 18142 29080
rect 18194 29057 18211 29080
rect 18211 29057 18228 29080
rect 18280 29057 18287 29080
rect 18287 29057 18314 29080
rect 18022 29046 18056 29057
rect 18108 29046 18142 29057
rect 18194 29046 18228 29057
rect 18280 29046 18314 29057
rect 18366 29046 18400 29080
rect 18022 28989 18025 29008
rect 18025 28989 18056 29008
rect 18108 28989 18135 29008
rect 18135 28989 18142 29008
rect 18194 28989 18211 29008
rect 18211 28989 18228 29008
rect 18280 28989 18287 29008
rect 18287 28989 18314 29008
rect 18022 28974 18056 28989
rect 18108 28974 18142 28989
rect 18194 28974 18228 28989
rect 18280 28974 18314 28989
rect 18366 28974 18400 29008
rect 18022 28921 18025 28936
rect 18025 28921 18056 28936
rect 18108 28921 18135 28936
rect 18135 28921 18142 28936
rect 18194 28921 18211 28936
rect 18211 28921 18228 28936
rect 18280 28921 18287 28936
rect 18287 28921 18314 28936
rect 18022 28902 18056 28921
rect 18108 28902 18142 28921
rect 18194 28902 18228 28921
rect 18280 28902 18314 28921
rect 18366 28902 18400 28936
rect 18022 28853 18025 28864
rect 18025 28853 18056 28864
rect 18108 28853 18135 28864
rect 18135 28853 18142 28864
rect 18194 28853 18211 28864
rect 18211 28853 18228 28864
rect 18280 28853 18287 28864
rect 18287 28853 18314 28864
rect 18022 28830 18056 28853
rect 18108 28830 18142 28853
rect 18194 28830 18228 28853
rect 18280 28830 18314 28853
rect 18366 28830 18400 28864
rect 18022 28785 18025 28792
rect 18025 28785 18056 28792
rect 18108 28785 18135 28792
rect 18135 28785 18142 28792
rect 18194 28785 18211 28792
rect 18211 28785 18228 28792
rect 18280 28785 18287 28792
rect 18287 28785 18314 28792
rect 18022 28758 18056 28785
rect 18108 28758 18142 28785
rect 18194 28758 18228 28785
rect 18280 28758 18314 28785
rect 18366 28758 18400 28792
rect 18022 28717 18025 28720
rect 18025 28717 18056 28720
rect 18108 28717 18135 28720
rect 18135 28717 18142 28720
rect 18194 28717 18211 28720
rect 18211 28717 18228 28720
rect 18280 28717 18287 28720
rect 18287 28717 18314 28720
rect 18022 28686 18056 28717
rect 18108 28686 18142 28717
rect 18194 28686 18228 28717
rect 18280 28686 18314 28717
rect 18366 28686 18400 28720
rect 18022 28615 18056 28648
rect 18108 28615 18142 28648
rect 18194 28615 18228 28648
rect 18280 28615 18314 28648
rect 18022 28614 18025 28615
rect 18025 28614 18056 28615
rect 18108 28614 18135 28615
rect 18135 28614 18142 28615
rect 18194 28614 18211 28615
rect 18211 28614 18228 28615
rect 18280 28614 18287 28615
rect 18287 28614 18314 28615
rect 18366 28614 18400 28648
rect 18022 28547 18056 28576
rect 18108 28547 18142 28576
rect 18194 28547 18228 28576
rect 18280 28547 18314 28576
rect 18022 28542 18025 28547
rect 18025 28542 18056 28547
rect 18108 28542 18135 28547
rect 18135 28542 18142 28547
rect 18194 28542 18211 28547
rect 18211 28542 18228 28547
rect 18280 28542 18287 28547
rect 18287 28542 18314 28547
rect 18366 28542 18400 28576
rect 18022 28479 18056 28504
rect 18108 28479 18142 28504
rect 18194 28479 18228 28504
rect 18280 28479 18314 28504
rect 18022 28470 18025 28479
rect 18025 28470 18056 28479
rect 18108 28470 18135 28479
rect 18135 28470 18142 28479
rect 18194 28470 18211 28479
rect 18211 28470 18228 28479
rect 18280 28470 18287 28479
rect 18287 28470 18314 28479
rect 18366 28470 18400 28504
rect 18022 28411 18056 28432
rect 18108 28411 18142 28432
rect 18194 28411 18228 28432
rect 18280 28411 18314 28432
rect 18022 28398 18025 28411
rect 18025 28398 18056 28411
rect 18108 28398 18135 28411
rect 18135 28398 18142 28411
rect 18194 28398 18211 28411
rect 18211 28398 18228 28411
rect 18280 28398 18287 28411
rect 18287 28398 18314 28411
rect 18366 28398 18400 28432
rect 18022 28343 18056 28360
rect 18108 28343 18142 28360
rect 18194 28343 18228 28360
rect 18280 28343 18314 28360
rect 18022 28326 18025 28343
rect 18025 28326 18056 28343
rect 18108 28326 18135 28343
rect 18135 28326 18142 28343
rect 18194 28326 18211 28343
rect 18211 28326 18228 28343
rect 18280 28326 18287 28343
rect 18287 28326 18314 28343
rect 18366 28326 18400 28360
rect 18022 28275 18056 28288
rect 18108 28275 18142 28288
rect 18194 28275 18228 28288
rect 18280 28275 18314 28288
rect 18022 28254 18025 28275
rect 18025 28254 18056 28275
rect 18108 28254 18135 28275
rect 18135 28254 18142 28275
rect 18194 28254 18211 28275
rect 18211 28254 18228 28275
rect 18280 28254 18287 28275
rect 18287 28254 18314 28275
rect 18366 28254 18400 28288
rect 18022 28207 18056 28216
rect 18108 28207 18142 28216
rect 18194 28207 18228 28216
rect 18280 28207 18314 28216
rect 18022 28182 18025 28207
rect 18025 28182 18056 28207
rect 18108 28182 18135 28207
rect 18135 28182 18142 28207
rect 18194 28182 18211 28207
rect 18211 28182 18228 28207
rect 18280 28182 18287 28207
rect 18287 28182 18314 28207
rect 18366 28182 18400 28216
rect 18022 28139 18056 28144
rect 18108 28139 18142 28144
rect 18194 28139 18228 28144
rect 18280 28139 18314 28144
rect 18022 28110 18025 28139
rect 18025 28110 18056 28139
rect 18108 28110 18135 28139
rect 18135 28110 18142 28139
rect 18194 28110 18211 28139
rect 18211 28110 18228 28139
rect 18280 28110 18287 28139
rect 18287 28110 18314 28139
rect 18366 28110 18400 28144
rect 18022 28071 18056 28072
rect 18108 28071 18142 28072
rect 18194 28071 18228 28072
rect 18280 28071 18314 28072
rect 18022 28038 18025 28071
rect 18025 28038 18056 28071
rect 18108 28038 18135 28071
rect 18135 28038 18142 28071
rect 18194 28038 18211 28071
rect 18211 28038 18228 28071
rect 18280 28038 18287 28071
rect 18287 28038 18314 28071
rect 18366 28038 18400 28072
rect 18022 27969 18025 28000
rect 18025 27969 18056 28000
rect 18108 27969 18135 28000
rect 18135 27969 18142 28000
rect 18194 27969 18211 28000
rect 18211 27969 18228 28000
rect 18280 27969 18287 28000
rect 18287 27969 18314 28000
rect 18022 27966 18056 27969
rect 18108 27966 18142 27969
rect 18194 27966 18228 27969
rect 18280 27966 18314 27969
rect 18366 27966 18400 28000
rect 18022 27901 18025 27928
rect 18025 27901 18056 27928
rect 18108 27901 18135 27928
rect 18135 27901 18142 27928
rect 18194 27901 18211 27928
rect 18211 27901 18228 27928
rect 18280 27901 18287 27928
rect 18287 27901 18314 27928
rect 18022 27894 18056 27901
rect 18108 27894 18142 27901
rect 18194 27894 18228 27901
rect 18280 27894 18314 27901
rect 18366 27894 18400 27928
rect 18022 27833 18025 27856
rect 18025 27833 18056 27856
rect 18108 27833 18135 27856
rect 18135 27833 18142 27856
rect 18194 27833 18211 27856
rect 18211 27833 18228 27856
rect 18280 27833 18287 27856
rect 18287 27833 18314 27856
rect 18022 27822 18056 27833
rect 18108 27822 18142 27833
rect 18194 27822 18228 27833
rect 18280 27822 18314 27833
rect 18366 27822 18400 27856
rect 18022 27765 18025 27784
rect 18025 27765 18056 27784
rect 18108 27765 18135 27784
rect 18135 27765 18142 27784
rect 18194 27765 18211 27784
rect 18211 27765 18228 27784
rect 18280 27765 18287 27784
rect 18287 27765 18314 27784
rect 18022 27750 18056 27765
rect 18108 27750 18142 27765
rect 18194 27750 18228 27765
rect 18280 27750 18314 27765
rect 18366 27750 18400 27784
rect 18022 27697 18025 27712
rect 18025 27697 18056 27712
rect 18108 27697 18135 27712
rect 18135 27697 18142 27712
rect 18194 27697 18211 27712
rect 18211 27697 18228 27712
rect 18280 27697 18287 27712
rect 18287 27697 18314 27712
rect 18022 27678 18056 27697
rect 18108 27678 18142 27697
rect 18194 27678 18228 27697
rect 18280 27678 18314 27697
rect 18366 27678 18400 27712
rect 18022 27629 18025 27640
rect 18025 27629 18056 27640
rect 18108 27629 18135 27640
rect 18135 27629 18142 27640
rect 18194 27629 18211 27640
rect 18211 27629 18228 27640
rect 18280 27629 18287 27640
rect 18287 27629 18314 27640
rect 18022 27606 18056 27629
rect 18108 27606 18142 27629
rect 18194 27606 18228 27629
rect 18280 27606 18314 27629
rect 18366 27606 18400 27640
rect 18022 27561 18025 27568
rect 18025 27561 18056 27568
rect 18108 27561 18135 27568
rect 18135 27561 18142 27568
rect 18194 27561 18211 27568
rect 18211 27561 18228 27568
rect 18280 27561 18287 27568
rect 18287 27561 18314 27568
rect 18022 27534 18056 27561
rect 18108 27534 18142 27561
rect 18194 27534 18228 27561
rect 18280 27534 18314 27561
rect 18366 27534 18400 27568
rect 18022 27493 18025 27496
rect 18025 27493 18056 27496
rect 18108 27493 18135 27496
rect 18135 27493 18142 27496
rect 18194 27493 18211 27496
rect 18211 27493 18228 27496
rect 18280 27493 18287 27496
rect 18287 27493 18314 27496
rect 18022 27462 18056 27493
rect 18108 27462 18142 27493
rect 18194 27462 18228 27493
rect 18280 27462 18314 27493
rect 18366 27462 18400 27496
rect 18022 27391 18056 27424
rect 18108 27391 18142 27424
rect 18194 27391 18228 27424
rect 18280 27391 18314 27424
rect 18022 27390 18025 27391
rect 18025 27390 18056 27391
rect 18108 27390 18135 27391
rect 18135 27390 18142 27391
rect 18194 27390 18211 27391
rect 18211 27390 18228 27391
rect 18280 27390 18287 27391
rect 18287 27390 18314 27391
rect 18366 27390 18400 27424
rect 18022 27323 18056 27352
rect 18108 27323 18142 27352
rect 18194 27323 18228 27352
rect 18280 27323 18314 27352
rect 18022 27318 18025 27323
rect 18025 27318 18056 27323
rect 18108 27318 18135 27323
rect 18135 27318 18142 27323
rect 18194 27318 18211 27323
rect 18211 27318 18228 27323
rect 18280 27318 18287 27323
rect 18287 27318 18314 27323
rect 18366 27318 18400 27352
rect 18022 27255 18056 27280
rect 18108 27255 18142 27280
rect 18194 27255 18228 27280
rect 18280 27255 18314 27280
rect 18022 27246 18025 27255
rect 18025 27246 18056 27255
rect 18108 27246 18135 27255
rect 18135 27246 18142 27255
rect 18194 27246 18211 27255
rect 18211 27246 18228 27255
rect 18280 27246 18287 27255
rect 18287 27246 18314 27255
rect 18366 27246 18400 27280
rect 18022 27187 18056 27208
rect 18108 27187 18142 27208
rect 18194 27187 18228 27208
rect 18280 27187 18314 27208
rect 18022 27174 18025 27187
rect 18025 27174 18056 27187
rect 18108 27174 18135 27187
rect 18135 27174 18142 27187
rect 18194 27174 18211 27187
rect 18211 27174 18228 27187
rect 18280 27174 18287 27187
rect 18287 27174 18314 27187
rect 18366 27174 18400 27208
rect 1470 27010 1504 27015
rect 1544 27010 1578 27015
rect 1618 27010 1652 27015
rect 1692 27010 1726 27015
rect 1395 26976 1397 27006
rect 1397 26976 1429 27006
rect 1470 26981 1499 27010
rect 1499 26981 1504 27010
rect 1544 26981 1567 27010
rect 1567 26981 1578 27010
rect 1618 26981 1635 27010
rect 1635 26981 1652 27010
rect 1692 26981 1703 27010
rect 1703 26981 1726 27010
rect 1395 26972 1429 26976
rect 1470 26941 1504 26943
rect 1544 26941 1578 26943
rect 1618 26941 1652 26943
rect 1692 26941 1726 26943
rect 1395 26907 1397 26932
rect 1397 26907 1429 26932
rect 1470 26909 1499 26941
rect 1499 26909 1504 26941
rect 1544 26909 1567 26941
rect 1567 26909 1578 26941
rect 1618 26909 1635 26941
rect 1635 26909 1652 26941
rect 1692 26909 1703 26941
rect 1703 26909 1726 26941
rect 1395 26898 1429 26907
rect 1395 26838 1397 26858
rect 1397 26838 1429 26858
rect 1470 26838 1499 26871
rect 1499 26838 1504 26871
rect 1544 26838 1567 26871
rect 1567 26838 1578 26871
rect 1618 26838 1635 26871
rect 1635 26838 1652 26871
rect 1692 26838 1703 26871
rect 1703 26838 1726 26871
rect 1395 26824 1429 26838
rect 1470 26837 1504 26838
rect 1544 26837 1578 26838
rect 1618 26837 1652 26838
rect 1692 26837 1726 26838
rect 1395 26769 1397 26784
rect 1397 26769 1429 26784
rect 1470 26769 1499 26799
rect 1499 26769 1504 26799
rect 1544 26769 1567 26799
rect 1567 26769 1578 26799
rect 1618 26769 1635 26799
rect 1635 26769 1652 26799
rect 1692 26769 1703 26799
rect 1703 26769 1726 26799
rect 1395 26750 1429 26769
rect 1470 26765 1504 26769
rect 1544 26765 1578 26769
rect 1618 26765 1652 26769
rect 1692 26765 1726 26769
rect 1395 26700 1397 26710
rect 1397 26700 1429 26710
rect 1470 26700 1499 26727
rect 1499 26700 1504 26727
rect 1544 26700 1567 26727
rect 1567 26700 1578 26727
rect 1618 26700 1635 26727
rect 1635 26700 1652 26727
rect 1692 26700 1703 26727
rect 1703 26700 1726 26727
rect 1395 26676 1429 26700
rect 1470 26693 1504 26700
rect 1544 26693 1578 26700
rect 1618 26693 1652 26700
rect 1692 26693 1726 26700
rect 1395 26631 1397 26636
rect 1397 26631 1429 26636
rect 1470 26631 1499 26655
rect 1499 26631 1504 26655
rect 1544 26631 1567 26655
rect 1567 26631 1578 26655
rect 1618 26631 1635 26655
rect 1635 26631 1652 26655
rect 1692 26631 1703 26655
rect 1703 26631 1726 26655
rect 1395 26602 1429 26631
rect 1470 26621 1504 26631
rect 1544 26621 1578 26631
rect 1618 26621 1652 26631
rect 1692 26621 1726 26631
rect 1470 26562 1499 26583
rect 1499 26562 1504 26583
rect 1544 26562 1567 26583
rect 1567 26562 1578 26583
rect 1618 26562 1635 26583
rect 1635 26562 1652 26583
rect 1692 26562 1703 26583
rect 1703 26562 1726 26583
rect 1395 26528 1429 26562
rect 1470 26549 1504 26562
rect 1544 26549 1578 26562
rect 1618 26549 1652 26562
rect 1692 26549 1726 26562
rect 1470 26493 1499 26511
rect 1499 26493 1504 26511
rect 1544 26493 1567 26511
rect 1567 26493 1578 26511
rect 1618 26493 1635 26511
rect 1635 26493 1652 26511
rect 1692 26493 1703 26511
rect 1703 26493 1726 26511
rect 1395 26458 1429 26488
rect 1470 26477 1504 26493
rect 1544 26477 1578 26493
rect 1618 26477 1652 26493
rect 1692 26477 1726 26493
rect 1395 26454 1397 26458
rect 1397 26454 1429 26458
rect 1470 26424 1499 26439
rect 1499 26424 1504 26439
rect 1544 26424 1567 26439
rect 1567 26424 1578 26439
rect 1618 26424 1635 26439
rect 1635 26424 1652 26439
rect 1692 26424 1703 26439
rect 1703 26424 1726 26439
rect 1395 26389 1429 26414
rect 1470 26405 1504 26424
rect 1544 26405 1578 26424
rect 1618 26405 1652 26424
rect 1692 26405 1726 26424
rect 1395 26380 1397 26389
rect 1397 26380 1429 26389
rect 1470 26355 1499 26367
rect 1499 26355 1504 26367
rect 1544 26355 1567 26367
rect 1567 26355 1578 26367
rect 1618 26355 1635 26367
rect 1635 26355 1652 26367
rect 1692 26355 1703 26367
rect 1703 26355 1726 26367
rect 1395 26320 1429 26340
rect 1470 26333 1504 26355
rect 1544 26333 1578 26355
rect 1618 26333 1652 26355
rect 1692 26333 1726 26355
rect 1395 26306 1397 26320
rect 1397 26306 1429 26320
rect 1470 26286 1499 26295
rect 1499 26286 1504 26295
rect 1544 26286 1567 26295
rect 1567 26286 1578 26295
rect 1618 26286 1635 26295
rect 1635 26286 1652 26295
rect 1692 26286 1703 26295
rect 1703 26286 1726 26295
rect 1395 26251 1429 26266
rect 1470 26261 1504 26286
rect 1544 26261 1578 26286
rect 1618 26261 1652 26286
rect 1692 26261 1726 26286
rect 1395 26232 1397 26251
rect 1397 26232 1429 26251
rect 1470 26217 1499 26223
rect 1499 26217 1504 26223
rect 1544 26217 1567 26223
rect 1567 26217 1578 26223
rect 1618 26217 1635 26223
rect 1635 26217 1652 26223
rect 1692 26217 1703 26223
rect 1703 26217 1726 26223
rect 1395 26182 1429 26193
rect 1470 26189 1504 26217
rect 1544 26189 1578 26217
rect 1618 26189 1652 26217
rect 1692 26189 1726 26217
rect 1395 26159 1397 26182
rect 1397 26159 1429 26182
rect 1470 26148 1499 26151
rect 1499 26148 1504 26151
rect 1544 26148 1567 26151
rect 1567 26148 1578 26151
rect 1618 26148 1635 26151
rect 1635 26148 1652 26151
rect 1692 26148 1703 26151
rect 1703 26148 1726 26151
rect 1395 26113 1429 26120
rect 1470 26117 1504 26148
rect 1544 26117 1578 26148
rect 1618 26117 1652 26148
rect 1692 26117 1726 26148
rect 1395 26086 1397 26113
rect 1397 26086 1429 26113
rect 1395 26044 1429 26047
rect 1470 26045 1504 26079
rect 1544 26045 1578 26079
rect 1618 26045 1652 26079
rect 1692 26045 1726 26079
rect 1395 26013 1397 26044
rect 1397 26013 1429 26044
rect 1470 25975 1504 26007
rect 1544 25975 1578 26007
rect 1618 25975 1652 26007
rect 1692 25975 1726 26007
rect 1395 25941 1397 25974
rect 1397 25941 1429 25974
rect 1470 25973 1499 25975
rect 1499 25973 1504 25975
rect 1544 25973 1567 25975
rect 1567 25973 1578 25975
rect 1618 25973 1635 25975
rect 1635 25973 1652 25975
rect 1692 25973 1703 25975
rect 1703 25973 1726 25975
rect 1395 25940 1429 25941
rect 1470 25906 1504 25935
rect 1544 25906 1578 25935
rect 1618 25906 1652 25935
rect 1692 25906 1726 25935
rect 1395 25872 1397 25901
rect 1397 25872 1429 25901
rect 1470 25901 1499 25906
rect 1499 25901 1504 25906
rect 1544 25901 1567 25906
rect 1567 25901 1578 25906
rect 1618 25901 1635 25906
rect 1635 25901 1652 25906
rect 1692 25901 1703 25906
rect 1703 25901 1726 25906
rect 1395 25867 1429 25872
rect 1470 25837 1504 25863
rect 1544 25837 1578 25863
rect 1618 25837 1652 25863
rect 1692 25837 1726 25863
rect 1395 25803 1397 25828
rect 1397 25803 1429 25828
rect 1470 25829 1499 25837
rect 1499 25829 1504 25837
rect 1544 25829 1567 25837
rect 1567 25829 1578 25837
rect 1618 25829 1635 25837
rect 1635 25829 1652 25837
rect 1692 25829 1703 25837
rect 1703 25829 1726 25837
rect 1395 25794 1429 25803
rect 1470 25768 1504 25791
rect 1544 25768 1578 25791
rect 1618 25768 1652 25791
rect 1692 25768 1726 25791
rect 1395 25734 1397 25755
rect 1397 25734 1429 25755
rect 1470 25757 1499 25768
rect 1499 25757 1504 25768
rect 1544 25757 1567 25768
rect 1567 25757 1578 25768
rect 1618 25757 1635 25768
rect 1635 25757 1652 25768
rect 1692 25757 1703 25768
rect 1703 25757 1726 25768
rect 1395 25721 1429 25734
rect 1470 25699 1504 25719
rect 1544 25699 1578 25719
rect 1618 25699 1652 25719
rect 1692 25699 1726 25719
rect 1395 25665 1397 25682
rect 1397 25665 1429 25682
rect 1470 25685 1499 25699
rect 1499 25685 1504 25699
rect 1544 25685 1567 25699
rect 1567 25685 1578 25699
rect 1618 25685 1635 25699
rect 1635 25685 1652 25699
rect 1692 25685 1703 25699
rect 1703 25685 1726 25699
rect 1395 25648 1429 25665
rect 1470 25630 1504 25647
rect 1544 25630 1578 25647
rect 1618 25630 1652 25647
rect 1692 25630 1726 25647
rect 1395 25596 1397 25609
rect 1397 25596 1429 25609
rect 1470 25613 1499 25630
rect 1499 25613 1504 25630
rect 1544 25613 1567 25630
rect 1567 25613 1578 25630
rect 1618 25613 1635 25630
rect 1635 25613 1652 25630
rect 1692 25613 1703 25630
rect 1703 25613 1726 25630
rect 1395 25575 1429 25596
rect 1470 25561 1504 25575
rect 1544 25561 1578 25575
rect 1618 25561 1652 25575
rect 1692 25561 1726 25575
rect 1470 25541 1499 25561
rect 1499 25541 1504 25561
rect 1544 25541 1567 25561
rect 1567 25541 1578 25561
rect 1618 25541 1635 25561
rect 1635 25541 1652 25561
rect 1692 25541 1703 25561
rect 1703 25541 1726 25561
rect 1470 25492 1504 25502
rect 1544 25492 1578 25502
rect 1618 25492 1652 25502
rect 1692 25492 1726 25502
rect 1470 25468 1499 25492
rect 1499 25468 1504 25492
rect 1544 25468 1567 25492
rect 1567 25468 1578 25492
rect 1618 25468 1635 25492
rect 1635 25468 1652 25492
rect 1692 25468 1703 25492
rect 1703 25468 1726 25492
rect 1470 25423 1504 25429
rect 1544 25423 1578 25429
rect 1618 25423 1652 25429
rect 1692 25423 1726 25429
rect 1470 25395 1499 25423
rect 1499 25395 1504 25423
rect 1544 25395 1567 25423
rect 1567 25395 1578 25423
rect 1618 25395 1635 25423
rect 1635 25395 1652 25423
rect 1692 25395 1703 25423
rect 1703 25395 1726 25423
rect 1470 25354 1504 25356
rect 1544 25354 1578 25356
rect 1618 25354 1652 25356
rect 1692 25354 1726 25356
rect 1470 25322 1499 25354
rect 1499 25322 1504 25354
rect 1544 25322 1567 25354
rect 1567 25322 1578 25354
rect 1618 25322 1635 25354
rect 1635 25322 1652 25354
rect 1692 25322 1703 25354
rect 1703 25322 1726 25354
rect 1059 25182 1091 25209
rect 1091 25182 1093 25209
rect 1133 25182 1159 25209
rect 1159 25182 1167 25209
rect 1207 25182 1227 25209
rect 1227 25182 1241 25209
rect 1281 25182 1295 25209
rect 1295 25182 1315 25209
rect 1355 25182 1363 25209
rect 1363 25182 1389 25209
rect 1429 25182 1431 25209
rect 1431 25182 1463 25209
rect 1503 25182 1533 25209
rect 1533 25182 1537 25209
rect 1577 25182 1601 25209
rect 1601 25182 1611 25209
rect 1651 25182 1669 25209
rect 1669 25182 1685 25209
rect 1059 25175 1093 25182
rect 1133 25175 1167 25182
rect 1207 25175 1241 25182
rect 1281 25175 1315 25182
rect 1355 25175 1389 25182
rect 1429 25175 1463 25182
rect 1503 25175 1537 25182
rect 1577 25175 1611 25182
rect 1651 25175 1685 25182
rect 1059 25113 1091 25134
rect 1091 25113 1093 25134
rect 1133 25113 1159 25134
rect 1159 25113 1167 25134
rect 1207 25113 1227 25134
rect 1227 25113 1241 25134
rect 1281 25113 1295 25134
rect 1295 25113 1315 25134
rect 1355 25113 1363 25134
rect 1363 25113 1389 25134
rect 1429 25113 1431 25134
rect 1431 25113 1463 25134
rect 1503 25113 1533 25134
rect 1533 25113 1537 25134
rect 1577 25113 1601 25134
rect 1601 25113 1611 25134
rect 1651 25113 1669 25134
rect 1669 25113 1685 25134
rect 1059 25100 1093 25113
rect 1133 25100 1167 25113
rect 1207 25100 1241 25113
rect 1281 25100 1315 25113
rect 1355 25100 1389 25113
rect 1429 25100 1463 25113
rect 1503 25100 1537 25113
rect 1577 25100 1611 25113
rect 1651 25100 1685 25113
rect 1059 25043 1091 25059
rect 1091 25043 1093 25059
rect 1133 25043 1159 25059
rect 1159 25043 1167 25059
rect 1207 25043 1227 25059
rect 1227 25043 1241 25059
rect 1281 25043 1295 25059
rect 1295 25043 1315 25059
rect 1355 25043 1363 25059
rect 1363 25043 1389 25059
rect 1429 25043 1431 25059
rect 1431 25043 1463 25059
rect 1503 25043 1533 25059
rect 1533 25043 1537 25059
rect 1577 25043 1601 25059
rect 1601 25043 1611 25059
rect 1651 25043 1669 25059
rect 1669 25043 1685 25059
rect 1059 25025 1093 25043
rect 1133 25025 1167 25043
rect 1207 25025 1241 25043
rect 1281 25025 1315 25043
rect 1355 25025 1389 25043
rect 1429 25025 1463 25043
rect 1503 25025 1537 25043
rect 1577 25025 1611 25043
rect 1651 25025 1685 25043
rect 1059 24973 1091 24984
rect 1091 24973 1093 24984
rect 1133 24973 1159 24984
rect 1159 24973 1167 24984
rect 1207 24973 1227 24984
rect 1227 24973 1241 24984
rect 1281 24973 1295 24984
rect 1295 24973 1315 24984
rect 1355 24973 1363 24984
rect 1363 24973 1389 24984
rect 1429 24973 1431 24984
rect 1431 24973 1463 24984
rect 1503 24973 1533 24984
rect 1533 24973 1537 24984
rect 1577 24973 1601 24984
rect 1601 24973 1611 24984
rect 1651 24973 1669 24984
rect 1669 24973 1685 24984
rect 1059 24950 1093 24973
rect 1133 24950 1167 24973
rect 1207 24950 1241 24973
rect 1281 24950 1315 24973
rect 1355 24950 1389 24973
rect 1429 24950 1463 24973
rect 1503 24950 1537 24973
rect 1577 24950 1611 24973
rect 1651 24950 1685 24973
rect 1059 24903 1091 24909
rect 1091 24903 1093 24909
rect 1133 24903 1159 24909
rect 1159 24903 1167 24909
rect 1207 24903 1227 24909
rect 1227 24903 1241 24909
rect 1281 24903 1295 24909
rect 1295 24903 1315 24909
rect 1355 24903 1363 24909
rect 1363 24903 1389 24909
rect 1429 24903 1431 24909
rect 1431 24903 1463 24909
rect 1503 24903 1533 24909
rect 1533 24903 1537 24909
rect 1577 24903 1601 24909
rect 1601 24903 1611 24909
rect 1651 24903 1669 24909
rect 1669 24903 1685 24909
rect 1059 24875 1093 24903
rect 1133 24875 1167 24903
rect 1207 24875 1241 24903
rect 1281 24875 1315 24903
rect 1355 24875 1389 24903
rect 1429 24875 1463 24903
rect 1503 24875 1537 24903
rect 1577 24875 1611 24903
rect 1651 24875 1685 24903
rect 1059 24833 1091 24834
rect 1091 24833 1093 24834
rect 1133 24833 1159 24834
rect 1159 24833 1167 24834
rect 1207 24833 1227 24834
rect 1227 24833 1241 24834
rect 1281 24833 1295 24834
rect 1295 24833 1315 24834
rect 1355 24833 1363 24834
rect 1363 24833 1389 24834
rect 1429 24833 1431 24834
rect 1431 24833 1463 24834
rect 1503 24833 1533 24834
rect 1533 24833 1537 24834
rect 1577 24833 1601 24834
rect 1601 24833 1611 24834
rect 1651 24833 1669 24834
rect 1669 24833 1685 24834
rect 1059 24800 1093 24833
rect 1133 24800 1167 24833
rect 1207 24800 1241 24833
rect 1281 24800 1315 24833
rect 1355 24800 1389 24833
rect 1429 24800 1463 24833
rect 1503 24800 1537 24833
rect 1577 24800 1611 24833
rect 1651 24800 1685 24833
rect 1059 24727 1093 24759
rect 1133 24727 1167 24759
rect 1207 24727 1241 24759
rect 1281 24727 1315 24759
rect 1355 24727 1389 24759
rect 1429 24727 1463 24759
rect 1503 24727 1537 24759
rect 1577 24727 1611 24759
rect 1651 24727 1685 24759
rect 1059 24725 1091 24727
rect 1091 24725 1093 24727
rect 1133 24725 1159 24727
rect 1159 24725 1167 24727
rect 1207 24725 1227 24727
rect 1227 24725 1241 24727
rect 1281 24725 1295 24727
rect 1295 24725 1315 24727
rect 1355 24725 1363 24727
rect 1363 24725 1389 24727
rect 1429 24725 1431 24727
rect 1431 24725 1463 24727
rect 1503 24725 1533 24727
rect 1533 24725 1537 24727
rect 1577 24725 1601 24727
rect 1601 24725 1611 24727
rect 1651 24725 1669 24727
rect 1669 24725 1685 24727
rect 1059 24657 1093 24684
rect 1133 24657 1167 24684
rect 1207 24657 1241 24684
rect 1281 24657 1315 24684
rect 1355 24657 1389 24684
rect 1429 24657 1463 24684
rect 1503 24657 1537 24684
rect 1577 24657 1611 24684
rect 1651 24657 1685 24684
rect 1059 24650 1091 24657
rect 1091 24650 1093 24657
rect 1133 24650 1159 24657
rect 1159 24650 1167 24657
rect 1207 24650 1227 24657
rect 1227 24650 1241 24657
rect 1281 24650 1295 24657
rect 1295 24650 1315 24657
rect 1355 24650 1363 24657
rect 1363 24650 1389 24657
rect 1429 24650 1431 24657
rect 1431 24650 1463 24657
rect 1503 24650 1533 24657
rect 1533 24650 1537 24657
rect 1577 24650 1601 24657
rect 1601 24650 1611 24657
rect 1651 24650 1669 24657
rect 1669 24650 1685 24657
rect 1059 24587 1093 24609
rect 1133 24587 1167 24609
rect 1207 24587 1241 24609
rect 1281 24587 1315 24609
rect 1355 24587 1389 24609
rect 1429 24587 1463 24609
rect 1503 24587 1537 24609
rect 1577 24587 1611 24609
rect 1651 24587 1685 24609
rect 1059 24575 1091 24587
rect 1091 24575 1093 24587
rect 1133 24575 1159 24587
rect 1159 24575 1167 24587
rect 1207 24575 1227 24587
rect 1227 24575 1241 24587
rect 1281 24575 1295 24587
rect 1295 24575 1315 24587
rect 1355 24575 1363 24587
rect 1363 24575 1389 24587
rect 1429 24575 1431 24587
rect 1431 24575 1463 24587
rect 1503 24575 1533 24587
rect 1533 24575 1537 24587
rect 1577 24575 1601 24587
rect 1601 24575 1611 24587
rect 1651 24575 1669 24587
rect 1669 24575 1685 24587
rect 1059 24517 1093 24533
rect 1133 24517 1167 24533
rect 1207 24517 1241 24533
rect 1281 24517 1315 24533
rect 1355 24517 1389 24533
rect 1429 24517 1463 24533
rect 1503 24517 1537 24533
rect 1577 24517 1611 24533
rect 1651 24517 1685 24533
rect 1059 24499 1091 24517
rect 1091 24499 1093 24517
rect 1133 24499 1159 24517
rect 1159 24499 1167 24517
rect 1207 24499 1227 24517
rect 1227 24499 1241 24517
rect 1281 24499 1295 24517
rect 1295 24499 1315 24517
rect 1355 24499 1363 24517
rect 1363 24499 1389 24517
rect 1429 24499 1431 24517
rect 1431 24499 1463 24517
rect 1503 24499 1533 24517
rect 1533 24499 1537 24517
rect 1577 24499 1601 24517
rect 1601 24499 1611 24517
rect 1651 24499 1669 24517
rect 1669 24499 1685 24517
rect 1059 24447 1093 24457
rect 1133 24447 1167 24457
rect 1207 24447 1241 24457
rect 1281 24447 1315 24457
rect 1355 24447 1389 24457
rect 1429 24447 1463 24457
rect 1503 24447 1537 24457
rect 1577 24447 1611 24457
rect 1651 24447 1685 24457
rect 1059 24423 1091 24447
rect 1091 24423 1093 24447
rect 1133 24423 1159 24447
rect 1159 24423 1167 24447
rect 1207 24423 1227 24447
rect 1227 24423 1241 24447
rect 1281 24423 1295 24447
rect 1295 24423 1315 24447
rect 1355 24423 1363 24447
rect 1363 24423 1389 24447
rect 1429 24423 1431 24447
rect 1431 24423 1463 24447
rect 1503 24423 1533 24447
rect 1533 24423 1537 24447
rect 1577 24423 1601 24447
rect 1601 24423 1611 24447
rect 1651 24423 1669 24447
rect 1669 24423 1685 24447
rect 1059 24377 1093 24381
rect 1133 24377 1167 24381
rect 1207 24377 1241 24381
rect 1281 24377 1315 24381
rect 1355 24377 1389 24381
rect 1429 24377 1463 24381
rect 1503 24377 1537 24381
rect 1577 24377 1611 24381
rect 1651 24377 1685 24381
rect 1059 24347 1091 24377
rect 1091 24347 1093 24377
rect 1133 24347 1159 24377
rect 1159 24347 1167 24377
rect 1207 24347 1227 24377
rect 1227 24347 1241 24377
rect 1281 24347 1295 24377
rect 1295 24347 1315 24377
rect 1355 24347 1363 24377
rect 1363 24347 1389 24377
rect 1429 24347 1431 24377
rect 1431 24347 1463 24377
rect 1503 24347 1533 24377
rect 1533 24347 1537 24377
rect 1577 24347 1601 24377
rect 1601 24347 1611 24377
rect 1651 24347 1669 24377
rect 1669 24347 1685 24377
rect 1059 24273 1091 24305
rect 1091 24273 1093 24305
rect 1133 24273 1159 24305
rect 1159 24273 1167 24305
rect 1207 24273 1227 24305
rect 1227 24273 1241 24305
rect 1281 24273 1295 24305
rect 1295 24273 1315 24305
rect 1355 24273 1363 24305
rect 1363 24273 1389 24305
rect 1429 24273 1431 24305
rect 1431 24273 1463 24305
rect 1503 24273 1533 24305
rect 1533 24273 1537 24305
rect 1577 24273 1601 24305
rect 1601 24273 1611 24305
rect 1651 24273 1669 24305
rect 1669 24273 1685 24305
rect 1059 24271 1093 24273
rect 1133 24271 1167 24273
rect 1207 24271 1241 24273
rect 1281 24271 1315 24273
rect 1355 24271 1389 24273
rect 1429 24271 1463 24273
rect 1503 24271 1537 24273
rect 1577 24271 1611 24273
rect 1651 24271 1685 24273
rect 1059 24203 1091 24229
rect 1091 24203 1093 24229
rect 1133 24203 1159 24229
rect 1159 24203 1167 24229
rect 1207 24203 1227 24229
rect 1227 24203 1241 24229
rect 1281 24203 1295 24229
rect 1295 24203 1315 24229
rect 1355 24203 1363 24229
rect 1363 24203 1389 24229
rect 1429 24203 1431 24229
rect 1431 24203 1463 24229
rect 1503 24203 1533 24229
rect 1533 24203 1537 24229
rect 1577 24203 1601 24229
rect 1601 24203 1611 24229
rect 1651 24203 1669 24229
rect 1669 24203 1685 24229
rect 1059 24195 1093 24203
rect 1133 24195 1167 24203
rect 1207 24195 1241 24203
rect 1281 24195 1315 24203
rect 1355 24195 1389 24203
rect 1429 24195 1463 24203
rect 1503 24195 1537 24203
rect 1577 24195 1611 24203
rect 1651 24195 1685 24203
rect 1059 24133 1091 24153
rect 1091 24133 1093 24153
rect 1133 24133 1159 24153
rect 1159 24133 1167 24153
rect 1207 24133 1227 24153
rect 1227 24133 1241 24153
rect 1281 24133 1295 24153
rect 1295 24133 1315 24153
rect 1355 24133 1363 24153
rect 1363 24133 1389 24153
rect 1429 24133 1431 24153
rect 1431 24133 1463 24153
rect 1503 24133 1533 24153
rect 1533 24133 1537 24153
rect 1577 24133 1601 24153
rect 1601 24133 1611 24153
rect 1651 24133 1669 24153
rect 1669 24133 1685 24153
rect 1059 24119 1093 24133
rect 1133 24119 1167 24133
rect 1207 24119 1241 24133
rect 1281 24119 1315 24133
rect 1355 24119 1389 24133
rect 1429 24119 1463 24133
rect 1503 24119 1537 24133
rect 1577 24119 1611 24133
rect 1651 24119 1685 24133
rect 1059 24063 1091 24077
rect 1091 24063 1093 24077
rect 1133 24063 1159 24077
rect 1159 24063 1167 24077
rect 1207 24063 1227 24077
rect 1227 24063 1241 24077
rect 1281 24063 1295 24077
rect 1295 24063 1315 24077
rect 1355 24063 1363 24077
rect 1363 24063 1389 24077
rect 1429 24063 1431 24077
rect 1431 24063 1463 24077
rect 1503 24063 1533 24077
rect 1533 24063 1537 24077
rect 1577 24063 1601 24077
rect 1601 24063 1611 24077
rect 1651 24063 1669 24077
rect 1669 24063 1685 24077
rect 1059 24043 1093 24063
rect 1133 24043 1167 24063
rect 1207 24043 1241 24063
rect 1281 24043 1315 24063
rect 1355 24043 1389 24063
rect 1429 24043 1463 24063
rect 1503 24043 1537 24063
rect 1577 24043 1611 24063
rect 1651 24043 1685 24063
rect 1059 23993 1091 24001
rect 1091 23993 1093 24001
rect 1133 23993 1159 24001
rect 1159 23993 1167 24001
rect 1207 23993 1227 24001
rect 1227 23993 1241 24001
rect 1281 23993 1295 24001
rect 1295 23993 1315 24001
rect 1355 23993 1363 24001
rect 1363 23993 1389 24001
rect 1429 23993 1431 24001
rect 1431 23993 1463 24001
rect 1503 23993 1533 24001
rect 1533 23993 1537 24001
rect 1577 23993 1601 24001
rect 1601 23993 1611 24001
rect 1651 23993 1669 24001
rect 1669 23993 1685 24001
rect 1059 23967 1093 23993
rect 1133 23967 1167 23993
rect 1207 23967 1241 23993
rect 1281 23967 1315 23993
rect 1355 23967 1389 23993
rect 1429 23967 1463 23993
rect 1503 23967 1537 23993
rect 1577 23967 1611 23993
rect 1651 23967 1685 23993
rect 1059 23923 1091 23925
rect 1091 23923 1093 23925
rect 1133 23923 1159 23925
rect 1159 23923 1167 23925
rect 1207 23923 1227 23925
rect 1227 23923 1241 23925
rect 1281 23923 1295 23925
rect 1295 23923 1315 23925
rect 1355 23923 1363 23925
rect 1363 23923 1389 23925
rect 1429 23923 1431 23925
rect 1431 23923 1463 23925
rect 1503 23923 1533 23925
rect 1533 23923 1537 23925
rect 1577 23923 1601 23925
rect 1601 23923 1611 23925
rect 1651 23923 1669 23925
rect 1669 23923 1685 23925
rect 1059 23891 1093 23923
rect 1133 23891 1167 23923
rect 1207 23891 1241 23923
rect 1281 23891 1315 23923
rect 1355 23891 1389 23923
rect 1429 23891 1463 23923
rect 1503 23891 1537 23923
rect 1577 23891 1611 23923
rect 1651 23891 1685 23923
rect 1059 23815 1093 23849
rect 1133 23815 1167 23849
rect 1207 23815 1241 23849
rect 1281 23815 1315 23849
rect 1355 23815 1389 23849
rect 1429 23815 1463 23849
rect 1503 23815 1537 23849
rect 1577 23815 1611 23849
rect 1651 23815 1685 23849
rect 212 23690 246 23724
rect 288 23719 314 23724
rect 314 23719 322 23724
rect 364 23719 384 23724
rect 384 23719 398 23724
rect 440 23719 454 23724
rect 454 23719 474 23724
rect 288 23690 322 23719
rect 364 23690 398 23719
rect 440 23690 474 23719
rect 513 23683 547 23703
rect 590 23683 624 23703
rect 667 23683 701 23703
rect 744 23683 778 23703
rect 821 23683 855 23703
rect 898 23683 932 23703
rect 975 23683 1009 23703
rect 1052 23683 1086 23703
rect 1129 23683 1163 23703
rect 1206 23683 1240 23703
rect 1283 23683 1317 23703
rect 1360 23683 1394 23703
rect 1437 23683 1471 23703
rect 513 23669 524 23683
rect 524 23669 547 23683
rect 590 23669 594 23683
rect 594 23669 624 23683
rect 212 23618 246 23652
rect 288 23649 314 23652
rect 314 23649 322 23652
rect 364 23649 384 23652
rect 384 23649 398 23652
rect 440 23649 454 23652
rect 454 23649 474 23652
rect 667 23669 698 23683
rect 698 23669 701 23683
rect 744 23669 768 23683
rect 768 23669 778 23683
rect 821 23669 838 23683
rect 838 23669 855 23683
rect 898 23669 908 23683
rect 908 23669 932 23683
rect 975 23669 978 23683
rect 978 23669 1009 23683
rect 1052 23669 1084 23683
rect 1084 23669 1086 23683
rect 1129 23669 1154 23683
rect 1154 23669 1163 23683
rect 1206 23669 1224 23683
rect 1224 23669 1240 23683
rect 1283 23669 1294 23683
rect 1294 23669 1317 23683
rect 1360 23669 1364 23683
rect 1364 23669 1394 23683
rect 1437 23669 1468 23683
rect 1468 23669 1471 23683
rect 288 23618 322 23649
rect 364 23618 398 23649
rect 440 23618 474 23649
rect 513 23613 547 23623
rect 590 23613 624 23623
rect 667 23613 701 23623
rect 744 23613 778 23623
rect 821 23613 855 23623
rect 898 23613 932 23623
rect 975 23613 1009 23623
rect 1052 23613 1086 23623
rect 1129 23613 1163 23623
rect 1206 23613 1240 23623
rect 1283 23613 1317 23623
rect 1360 23613 1394 23623
rect 1437 23613 1471 23623
rect 513 23589 524 23613
rect 524 23589 547 23613
rect 590 23589 594 23613
rect 594 23589 624 23613
rect 212 23546 246 23580
rect 288 23579 314 23580
rect 314 23579 322 23580
rect 364 23579 384 23580
rect 384 23579 398 23580
rect 440 23579 454 23580
rect 454 23579 474 23580
rect 667 23589 698 23613
rect 698 23589 701 23613
rect 744 23589 768 23613
rect 768 23589 778 23613
rect 821 23589 838 23613
rect 838 23589 855 23613
rect 898 23589 908 23613
rect 908 23589 932 23613
rect 975 23589 978 23613
rect 978 23589 1009 23613
rect 1052 23589 1084 23613
rect 1084 23589 1086 23613
rect 1129 23589 1154 23613
rect 1154 23589 1163 23613
rect 1206 23589 1224 23613
rect 1224 23589 1240 23613
rect 1283 23589 1294 23613
rect 1294 23589 1317 23613
rect 1360 23589 1364 23613
rect 1364 23589 1394 23613
rect 1437 23589 1468 23613
rect 1468 23589 1471 23613
rect 18022 27119 18056 27136
rect 18108 27119 18142 27136
rect 18194 27119 18228 27136
rect 18280 27119 18314 27136
rect 18022 27102 18025 27119
rect 18025 27102 18056 27119
rect 18108 27102 18135 27119
rect 18135 27102 18142 27119
rect 18194 27102 18211 27119
rect 18211 27102 18228 27119
rect 18280 27102 18287 27119
rect 18287 27102 18314 27119
rect 18366 27102 18400 27136
rect 18022 27051 18056 27064
rect 18108 27051 18142 27064
rect 18194 27051 18228 27064
rect 18280 27051 18314 27064
rect 18022 27030 18025 27051
rect 18025 27030 18056 27051
rect 18108 27030 18135 27051
rect 18135 27030 18142 27051
rect 18194 27030 18211 27051
rect 18211 27030 18228 27051
rect 18280 27030 18287 27051
rect 18287 27030 18314 27051
rect 18366 27030 18400 27064
rect 18022 26983 18056 26992
rect 18108 26983 18142 26992
rect 18194 26983 18228 26992
rect 18280 26983 18314 26992
rect 18022 26958 18025 26983
rect 18025 26958 18056 26983
rect 18108 26958 18135 26983
rect 18135 26958 18142 26983
rect 18194 26958 18211 26983
rect 18211 26958 18228 26983
rect 18280 26958 18287 26983
rect 18287 26958 18314 26983
rect 18366 26958 18400 26992
rect 18022 26915 18056 26920
rect 18108 26915 18142 26920
rect 18194 26915 18228 26920
rect 18280 26915 18314 26920
rect 18022 26886 18025 26915
rect 18025 26886 18056 26915
rect 18108 26886 18135 26915
rect 18135 26886 18142 26915
rect 18194 26886 18211 26915
rect 18211 26886 18228 26915
rect 18280 26886 18287 26915
rect 18287 26886 18314 26915
rect 18366 26886 18400 26920
rect 18022 26847 18056 26848
rect 18108 26847 18142 26848
rect 18194 26847 18228 26848
rect 18280 26847 18314 26848
rect 18022 26814 18025 26847
rect 18025 26814 18056 26847
rect 18108 26814 18135 26847
rect 18135 26814 18142 26847
rect 18194 26814 18211 26847
rect 18211 26814 18228 26847
rect 18280 26814 18287 26847
rect 18287 26814 18314 26847
rect 18366 26814 18400 26848
rect 18022 26745 18025 26776
rect 18025 26745 18056 26776
rect 18108 26745 18135 26776
rect 18135 26745 18142 26776
rect 18194 26745 18211 26776
rect 18211 26745 18228 26776
rect 18280 26745 18287 26776
rect 18287 26745 18314 26776
rect 18022 26742 18056 26745
rect 18108 26742 18142 26745
rect 18194 26742 18228 26745
rect 18280 26742 18314 26745
rect 18366 26742 18400 26776
rect 18022 26677 18025 26704
rect 18025 26677 18056 26704
rect 18108 26677 18135 26704
rect 18135 26677 18142 26704
rect 18194 26677 18211 26704
rect 18211 26677 18228 26704
rect 18280 26677 18287 26704
rect 18287 26677 18314 26704
rect 18022 26670 18056 26677
rect 18108 26670 18142 26677
rect 18194 26670 18228 26677
rect 18280 26670 18314 26677
rect 18366 26670 18400 26704
rect 18022 26609 18025 26632
rect 18025 26609 18056 26632
rect 18108 26609 18135 26632
rect 18135 26609 18142 26632
rect 18194 26609 18211 26632
rect 18211 26609 18228 26632
rect 18280 26609 18287 26632
rect 18287 26609 18314 26632
rect 18022 26598 18056 26609
rect 18108 26598 18142 26609
rect 18194 26598 18228 26609
rect 18280 26598 18314 26609
rect 18366 26598 18400 26632
rect 18022 26541 18025 26560
rect 18025 26541 18056 26560
rect 18108 26541 18135 26560
rect 18135 26541 18142 26560
rect 18194 26541 18211 26560
rect 18211 26541 18228 26560
rect 18280 26541 18287 26560
rect 18287 26541 18314 26560
rect 18022 26526 18056 26541
rect 18108 26526 18142 26541
rect 18194 26526 18228 26541
rect 18280 26526 18314 26541
rect 18366 26526 18400 26560
rect 18022 26473 18025 26488
rect 18025 26473 18056 26488
rect 18108 26473 18135 26488
rect 18135 26473 18142 26488
rect 18194 26473 18211 26488
rect 18211 26473 18228 26488
rect 18280 26473 18287 26488
rect 18287 26473 18314 26488
rect 18022 26454 18056 26473
rect 18108 26454 18142 26473
rect 18194 26454 18228 26473
rect 18280 26454 18314 26473
rect 18366 26454 18400 26488
rect 18022 26405 18025 26416
rect 18025 26405 18056 26416
rect 18108 26405 18135 26416
rect 18135 26405 18142 26416
rect 18194 26405 18211 26416
rect 18211 26405 18228 26416
rect 18280 26405 18287 26416
rect 18287 26405 18314 26416
rect 18022 26382 18056 26405
rect 18108 26382 18142 26405
rect 18194 26382 18228 26405
rect 18280 26382 18314 26405
rect 18366 26382 18400 26416
rect 18022 26337 18025 26344
rect 18025 26337 18056 26344
rect 18108 26337 18135 26344
rect 18135 26337 18142 26344
rect 18194 26337 18211 26344
rect 18211 26337 18228 26344
rect 18280 26337 18287 26344
rect 18287 26337 18314 26344
rect 18022 26310 18056 26337
rect 18108 26310 18142 26337
rect 18194 26310 18228 26337
rect 18280 26310 18314 26337
rect 18366 26310 18400 26344
rect 18022 26269 18025 26272
rect 18025 26269 18056 26272
rect 18108 26269 18135 26272
rect 18135 26269 18142 26272
rect 18194 26269 18211 26272
rect 18211 26269 18228 26272
rect 18280 26269 18287 26272
rect 18287 26269 18314 26272
rect 18022 26238 18056 26269
rect 18108 26238 18142 26269
rect 18194 26238 18228 26269
rect 18280 26238 18314 26269
rect 18366 26238 18400 26272
rect 18022 26167 18056 26200
rect 18108 26167 18142 26200
rect 18194 26167 18228 26200
rect 18280 26167 18314 26200
rect 18022 26166 18025 26167
rect 18025 26166 18056 26167
rect 18108 26166 18135 26167
rect 18135 26166 18142 26167
rect 18194 26166 18211 26167
rect 18211 26166 18228 26167
rect 18280 26166 18287 26167
rect 18287 26166 18314 26167
rect 18366 26166 18400 26200
rect 18022 26099 18056 26128
rect 18108 26099 18142 26128
rect 18194 26099 18228 26128
rect 18280 26099 18314 26128
rect 18022 26094 18025 26099
rect 18025 26094 18056 26099
rect 18108 26094 18135 26099
rect 18135 26094 18142 26099
rect 18194 26094 18211 26099
rect 18211 26094 18228 26099
rect 18280 26094 18287 26099
rect 18287 26094 18314 26099
rect 18366 26094 18400 26128
rect 18022 26031 18056 26056
rect 18108 26031 18142 26056
rect 18194 26031 18228 26056
rect 18280 26031 18314 26056
rect 18022 26022 18025 26031
rect 18025 26022 18056 26031
rect 18108 26022 18135 26031
rect 18135 26022 18142 26031
rect 18194 26022 18211 26031
rect 18211 26022 18228 26031
rect 18280 26022 18287 26031
rect 18287 26022 18314 26031
rect 18366 26022 18400 26056
rect 18022 25963 18056 25984
rect 18108 25963 18142 25984
rect 18194 25963 18228 25984
rect 18280 25963 18314 25984
rect 18022 25950 18025 25963
rect 18025 25950 18056 25963
rect 18108 25950 18135 25963
rect 18135 25950 18142 25963
rect 18194 25950 18211 25963
rect 18211 25950 18228 25963
rect 18280 25950 18287 25963
rect 18287 25950 18314 25963
rect 18366 25950 18400 25984
rect 18022 25895 18056 25912
rect 18108 25895 18142 25912
rect 18194 25895 18228 25912
rect 18280 25895 18314 25912
rect 18022 25878 18025 25895
rect 18025 25878 18056 25895
rect 18108 25878 18135 25895
rect 18135 25878 18142 25895
rect 18194 25878 18211 25895
rect 18211 25878 18228 25895
rect 18280 25878 18287 25895
rect 18287 25878 18314 25895
rect 18366 25878 18400 25912
rect 18022 25827 18056 25840
rect 18108 25827 18142 25840
rect 18194 25827 18228 25840
rect 18280 25827 18314 25840
rect 18022 25806 18025 25827
rect 18025 25806 18056 25827
rect 18108 25806 18135 25827
rect 18135 25806 18142 25827
rect 18194 25806 18211 25827
rect 18211 25806 18228 25827
rect 18280 25806 18287 25827
rect 18287 25806 18314 25827
rect 18366 25806 18400 25840
rect 18022 25759 18056 25768
rect 18108 25759 18142 25768
rect 18194 25759 18228 25768
rect 18280 25759 18314 25768
rect 18022 25734 18025 25759
rect 18025 25734 18056 25759
rect 18108 25734 18135 25759
rect 18135 25734 18142 25759
rect 18194 25734 18211 25759
rect 18211 25734 18228 25759
rect 18280 25734 18287 25759
rect 18287 25734 18314 25759
rect 18366 25734 18400 25768
rect 18022 25691 18056 25696
rect 18108 25691 18142 25696
rect 18194 25691 18228 25696
rect 18280 25691 18314 25696
rect 18022 25662 18025 25691
rect 18025 25662 18056 25691
rect 18108 25662 18135 25691
rect 18135 25662 18142 25691
rect 18194 25662 18211 25691
rect 18211 25662 18228 25691
rect 18280 25662 18287 25691
rect 18287 25662 18314 25691
rect 18366 25662 18400 25696
rect 18022 25623 18056 25624
rect 18108 25623 18142 25624
rect 18194 25623 18228 25624
rect 18280 25623 18314 25624
rect 18022 25590 18025 25623
rect 18025 25590 18056 25623
rect 18108 25590 18135 25623
rect 18135 25590 18142 25623
rect 18194 25590 18211 25623
rect 18211 25590 18228 25623
rect 18280 25590 18287 25623
rect 18287 25590 18314 25623
rect 18366 25590 18400 25624
rect 18022 25521 18025 25552
rect 18025 25521 18056 25552
rect 18108 25521 18135 25552
rect 18135 25521 18142 25552
rect 18194 25521 18211 25552
rect 18211 25521 18228 25552
rect 18280 25521 18287 25552
rect 18287 25521 18314 25552
rect 18022 25518 18056 25521
rect 18108 25518 18142 25521
rect 18194 25518 18228 25521
rect 18280 25518 18314 25521
rect 18366 25518 18400 25552
rect 18022 25453 18025 25480
rect 18025 25453 18056 25480
rect 18108 25453 18135 25480
rect 18135 25453 18142 25480
rect 18194 25453 18211 25480
rect 18211 25453 18228 25480
rect 18280 25453 18287 25480
rect 18287 25453 18314 25480
rect 18022 25446 18056 25453
rect 18108 25446 18142 25453
rect 18194 25446 18228 25453
rect 18280 25446 18314 25453
rect 18366 25446 18400 25480
rect 18022 25385 18025 25408
rect 18025 25385 18056 25408
rect 18108 25385 18135 25408
rect 18135 25385 18142 25408
rect 18194 25385 18211 25408
rect 18211 25385 18228 25408
rect 18280 25385 18287 25408
rect 18287 25385 18314 25408
rect 18022 25374 18056 25385
rect 18108 25374 18142 25385
rect 18194 25374 18228 25385
rect 18280 25374 18314 25385
rect 18366 25374 18400 25408
rect 18022 25317 18025 25336
rect 18025 25317 18056 25336
rect 18108 25317 18135 25336
rect 18135 25317 18142 25336
rect 18194 25317 18211 25336
rect 18211 25317 18228 25336
rect 18280 25317 18287 25336
rect 18287 25317 18314 25336
rect 18022 25302 18056 25317
rect 18108 25302 18142 25317
rect 18194 25302 18228 25317
rect 18280 25302 18314 25317
rect 18366 25302 18400 25336
rect 18022 25249 18025 25264
rect 18025 25249 18056 25264
rect 18108 25249 18135 25264
rect 18135 25249 18142 25264
rect 18194 25249 18211 25264
rect 18211 25249 18228 25264
rect 18280 25249 18287 25264
rect 18287 25249 18314 25264
rect 18022 25230 18056 25249
rect 18108 25230 18142 25249
rect 18194 25230 18228 25249
rect 18280 25230 18314 25249
rect 18366 25230 18400 25264
rect 18022 25180 18025 25192
rect 18025 25180 18056 25192
rect 18108 25180 18135 25192
rect 18135 25180 18142 25192
rect 18194 25180 18211 25192
rect 18211 25180 18228 25192
rect 18280 25180 18287 25192
rect 18287 25180 18314 25192
rect 18022 25158 18056 25180
rect 18108 25158 18142 25180
rect 18194 25158 18228 25180
rect 18280 25158 18314 25180
rect 18366 25158 18400 25192
rect 18022 25111 18025 25120
rect 18025 25111 18056 25120
rect 18108 25111 18135 25120
rect 18135 25111 18142 25120
rect 18194 25111 18211 25120
rect 18211 25111 18228 25120
rect 18280 25111 18287 25120
rect 18287 25111 18314 25120
rect 18022 25086 18056 25111
rect 18108 25086 18142 25111
rect 18194 25086 18228 25111
rect 18280 25086 18314 25111
rect 18366 25086 18400 25120
rect 18022 25042 18025 25048
rect 18025 25042 18056 25048
rect 18108 25042 18135 25048
rect 18135 25042 18142 25048
rect 18194 25042 18211 25048
rect 18211 25042 18228 25048
rect 18280 25042 18287 25048
rect 18287 25042 18314 25048
rect 18022 25014 18056 25042
rect 18108 25014 18142 25042
rect 18194 25014 18228 25042
rect 18280 25014 18314 25042
rect 18366 25014 18400 25048
rect 18022 24973 18025 24976
rect 18025 24973 18056 24976
rect 18108 24973 18135 24976
rect 18135 24973 18142 24976
rect 18194 24973 18211 24976
rect 18211 24973 18228 24976
rect 18280 24973 18287 24976
rect 18287 24973 18314 24976
rect 18022 24942 18056 24973
rect 18108 24942 18142 24973
rect 18194 24942 18228 24973
rect 18280 24942 18314 24973
rect 18366 24942 18400 24976
rect 18022 24870 18056 24904
rect 18108 24870 18142 24904
rect 18194 24870 18228 24904
rect 18280 24870 18314 24904
rect 18366 24870 18400 24904
rect 18022 24800 18056 24832
rect 18108 24800 18142 24832
rect 18194 24800 18228 24832
rect 18280 24800 18314 24832
rect 18022 24798 18025 24800
rect 18025 24798 18056 24800
rect 18108 24798 18135 24800
rect 18135 24798 18142 24800
rect 18194 24798 18211 24800
rect 18211 24798 18228 24800
rect 18280 24798 18287 24800
rect 18287 24798 18314 24800
rect 18366 24798 18400 24832
rect 18022 24731 18056 24760
rect 18108 24731 18142 24760
rect 18194 24731 18228 24760
rect 18280 24731 18314 24760
rect 18022 24726 18025 24731
rect 18025 24726 18056 24731
rect 18108 24726 18135 24731
rect 18135 24726 18142 24731
rect 18194 24726 18211 24731
rect 18211 24726 18228 24731
rect 18280 24726 18287 24731
rect 18287 24726 18314 24731
rect 18366 24726 18400 24760
rect 18022 24662 18056 24688
rect 18108 24662 18142 24688
rect 18194 24662 18228 24688
rect 18280 24662 18314 24688
rect 18022 24654 18025 24662
rect 18025 24654 18056 24662
rect 18108 24654 18135 24662
rect 18135 24654 18142 24662
rect 18194 24654 18211 24662
rect 18211 24654 18228 24662
rect 18280 24654 18287 24662
rect 18287 24654 18314 24662
rect 18366 24654 18400 24688
rect 18022 24593 18056 24616
rect 18108 24593 18142 24616
rect 18194 24593 18228 24616
rect 18280 24593 18314 24616
rect 18022 24582 18025 24593
rect 18025 24582 18056 24593
rect 18108 24582 18135 24593
rect 18135 24582 18142 24593
rect 18194 24582 18211 24593
rect 18211 24582 18228 24593
rect 18280 24582 18287 24593
rect 18287 24582 18314 24593
rect 18366 24582 18400 24616
rect 18022 24524 18056 24544
rect 18108 24524 18142 24544
rect 18194 24524 18228 24544
rect 18280 24524 18314 24544
rect 18022 24510 18025 24524
rect 18025 24510 18056 24524
rect 18108 24510 18135 24524
rect 18135 24510 18142 24524
rect 18194 24510 18211 24524
rect 18211 24510 18228 24524
rect 18280 24510 18287 24524
rect 18287 24510 18314 24524
rect 18366 24510 18400 24544
rect 18022 24455 18056 24472
rect 18108 24455 18142 24472
rect 18194 24455 18228 24472
rect 18280 24455 18314 24472
rect 18022 24438 18025 24455
rect 18025 24438 18056 24455
rect 18108 24438 18135 24455
rect 18135 24438 18142 24455
rect 18194 24438 18211 24455
rect 18211 24438 18228 24455
rect 18280 24438 18287 24455
rect 18287 24438 18314 24455
rect 18366 24438 18400 24472
rect 18022 24386 18056 24400
rect 18108 24386 18142 24400
rect 18194 24386 18228 24400
rect 18280 24386 18314 24400
rect 18022 24366 18025 24386
rect 18025 24366 18056 24386
rect 18108 24366 18135 24386
rect 18135 24366 18142 24386
rect 18194 24366 18211 24386
rect 18211 24366 18228 24386
rect 18280 24366 18287 24386
rect 18287 24366 18314 24386
rect 18366 24366 18400 24400
rect 18022 24317 18056 24328
rect 18108 24317 18142 24328
rect 18194 24317 18228 24328
rect 18280 24317 18314 24328
rect 18022 24294 18025 24317
rect 18025 24294 18056 24317
rect 18108 24294 18135 24317
rect 18135 24294 18142 24317
rect 18194 24294 18211 24317
rect 18211 24294 18228 24317
rect 18280 24294 18287 24317
rect 18287 24294 18314 24317
rect 18366 24294 18400 24328
rect 18022 24248 18056 24256
rect 18108 24248 18142 24256
rect 18194 24248 18228 24256
rect 18280 24248 18314 24256
rect 18022 24222 18025 24248
rect 18025 24222 18056 24248
rect 18108 24222 18135 24248
rect 18135 24222 18142 24248
rect 18194 24222 18211 24248
rect 18211 24222 18228 24248
rect 18280 24222 18287 24248
rect 18287 24222 18314 24248
rect 18366 24222 18400 24256
rect 18022 24179 18056 24184
rect 18108 24179 18142 24184
rect 18194 24179 18228 24184
rect 18280 24179 18314 24184
rect 18022 24150 18025 24179
rect 18025 24150 18056 24179
rect 18108 24150 18135 24179
rect 18135 24150 18142 24179
rect 18194 24150 18211 24179
rect 18211 24150 18228 24179
rect 18280 24150 18287 24179
rect 18287 24150 18314 24179
rect 18366 24150 18400 24184
rect 18022 24110 18056 24112
rect 18108 24110 18142 24112
rect 18194 24110 18228 24112
rect 18280 24110 18314 24112
rect 18022 24078 18025 24110
rect 18025 24078 18056 24110
rect 18108 24078 18135 24110
rect 18135 24078 18142 24110
rect 18194 24078 18211 24110
rect 18211 24078 18228 24110
rect 18280 24078 18287 24110
rect 18287 24078 18314 24110
rect 18366 24078 18400 24112
rect 18022 24007 18025 24040
rect 18025 24007 18056 24040
rect 18108 24007 18135 24040
rect 18135 24007 18142 24040
rect 18194 24007 18211 24040
rect 18211 24007 18228 24040
rect 18280 24007 18287 24040
rect 18287 24007 18314 24040
rect 18022 24006 18056 24007
rect 18108 24006 18142 24007
rect 18194 24006 18228 24007
rect 18280 24006 18314 24007
rect 18366 24006 18400 24040
rect 18022 23938 18025 23968
rect 18025 23938 18056 23968
rect 18108 23938 18135 23968
rect 18135 23938 18142 23968
rect 18194 23938 18211 23968
rect 18211 23938 18228 23968
rect 18280 23938 18287 23968
rect 18287 23938 18314 23968
rect 18022 23934 18056 23938
rect 18108 23934 18142 23938
rect 18194 23934 18228 23938
rect 18280 23934 18314 23938
rect 18366 23934 18400 23968
rect 18022 23869 18025 23896
rect 18025 23869 18056 23896
rect 18108 23869 18135 23896
rect 18135 23869 18142 23896
rect 18194 23869 18211 23896
rect 18211 23869 18228 23896
rect 18280 23869 18287 23896
rect 18287 23869 18314 23896
rect 18022 23862 18056 23869
rect 18108 23862 18142 23869
rect 18194 23862 18228 23869
rect 18280 23862 18314 23869
rect 18366 23862 18400 23896
rect 18022 23800 18025 23824
rect 18025 23800 18056 23824
rect 18108 23800 18135 23824
rect 18135 23800 18142 23824
rect 18194 23800 18211 23824
rect 18211 23800 18228 23824
rect 18280 23800 18287 23824
rect 18287 23800 18314 23824
rect 18022 23790 18056 23800
rect 18108 23790 18142 23800
rect 18194 23790 18228 23800
rect 18280 23790 18314 23800
rect 18366 23790 18400 23824
rect 18022 23731 18025 23752
rect 18025 23731 18056 23752
rect 18108 23731 18135 23752
rect 18135 23731 18142 23752
rect 18194 23731 18211 23752
rect 18211 23731 18228 23752
rect 18280 23731 18287 23752
rect 18287 23731 18314 23752
rect 18022 23718 18056 23731
rect 18108 23718 18142 23731
rect 18194 23718 18228 23731
rect 18280 23718 18314 23731
rect 18366 23718 18400 23752
rect 18022 23662 18025 23680
rect 18025 23662 18056 23680
rect 18108 23662 18135 23680
rect 18135 23662 18142 23680
rect 18194 23662 18211 23680
rect 18211 23662 18228 23680
rect 18280 23662 18287 23680
rect 18287 23662 18314 23680
rect 18022 23646 18056 23662
rect 18108 23646 18142 23662
rect 18194 23646 18228 23662
rect 18280 23646 18314 23662
rect 18366 23646 18400 23680
rect 288 23546 322 23579
rect 364 23546 398 23579
rect 440 23546 474 23579
rect 513 23509 524 23543
rect 524 23509 547 23543
rect 590 23509 594 23543
rect 594 23509 624 23543
rect 667 23509 698 23543
rect 698 23509 701 23543
rect 744 23509 768 23543
rect 768 23509 778 23543
rect 821 23509 838 23543
rect 838 23509 855 23543
rect 898 23509 908 23543
rect 908 23509 932 23543
rect 975 23509 978 23543
rect 978 23509 1009 23543
rect 1052 23509 1084 23543
rect 1084 23509 1086 23543
rect 1129 23509 1154 23543
rect 1154 23509 1163 23543
rect 1206 23509 1224 23543
rect 1224 23509 1240 23543
rect 1283 23509 1294 23543
rect 1294 23509 1317 23543
rect 1360 23509 1364 23543
rect 1364 23509 1394 23543
rect 1437 23509 1468 23543
rect 1468 23509 1471 23543
rect 212 23474 246 23508
rect 288 23474 322 23508
rect 364 23474 398 23508
rect 440 23474 474 23508
rect 18022 23593 18025 23607
rect 18025 23593 18056 23607
rect 18108 23593 18135 23607
rect 18135 23593 18142 23607
rect 18194 23593 18211 23607
rect 18211 23593 18228 23607
rect 18280 23593 18287 23607
rect 18287 23593 18314 23607
rect 18022 23573 18056 23593
rect 18108 23573 18142 23593
rect 18194 23573 18228 23593
rect 18280 23573 18314 23593
rect 18366 23573 18400 23607
rect 18022 23524 18025 23534
rect 18025 23524 18056 23534
rect 18108 23524 18135 23534
rect 18135 23524 18142 23534
rect 18194 23524 18211 23534
rect 18211 23524 18228 23534
rect 18280 23524 18287 23534
rect 18287 23524 18314 23534
rect 18022 23500 18056 23524
rect 18108 23500 18142 23524
rect 18194 23500 18228 23524
rect 18280 23500 18314 23524
rect 18366 23500 18400 23534
rect 22830 30712 22861 30717
rect 22861 30712 22864 30717
rect 22932 30712 22966 30746
rect 23034 30717 23068 30746
rect 23034 30712 23037 30717
rect 23037 30712 23068 30717
rect 22830 30649 22864 30671
rect 22830 30637 22861 30649
rect 22861 30637 22864 30649
rect 22932 30637 22966 30671
rect 23034 30649 23068 30671
rect 23034 30637 23037 30649
rect 23037 30637 23068 30649
rect 22830 30581 22864 30596
rect 22830 30562 22861 30581
rect 22861 30562 22864 30581
rect 22932 30562 22966 30596
rect 23034 30581 23068 30596
rect 23034 30562 23037 30581
rect 23037 30562 23068 30581
rect 22830 30513 22864 30521
rect 22830 30487 22861 30513
rect 22861 30487 22864 30513
rect 22932 30487 22966 30521
rect 23034 30513 23068 30521
rect 23034 30487 23037 30513
rect 23037 30487 23068 30513
rect 22830 30445 22864 30446
rect 22830 30412 22861 30445
rect 22861 30412 22864 30445
rect 22932 30412 22966 30446
rect 23034 30445 23068 30446
rect 23034 30412 23037 30445
rect 23037 30412 23068 30445
rect 22830 30343 22861 30371
rect 22861 30343 22864 30371
rect 22830 30337 22864 30343
rect 22932 30337 22966 30371
rect 23034 30343 23037 30371
rect 23037 30343 23068 30371
rect 23034 30337 23068 30343
rect 22830 30275 22861 30296
rect 22861 30275 22864 30296
rect 22830 30262 22864 30275
rect 22932 30262 22966 30296
rect 23034 30275 23037 30296
rect 23037 30275 23068 30296
rect 23034 30262 23068 30275
rect 22830 30207 22861 30221
rect 22861 30207 22864 30221
rect 22830 30187 22864 30207
rect 22932 30187 22966 30221
rect 23034 30207 23037 30221
rect 23037 30207 23068 30221
rect 23034 30187 23068 30207
rect 22830 30139 22861 30146
rect 22861 30139 22864 30146
rect 22830 30112 22864 30139
rect 22932 30112 22966 30146
rect 23034 30139 23037 30146
rect 23037 30139 23068 30146
rect 23034 30112 23068 30139
rect 22830 30037 22864 30071
rect 22932 30037 22966 30071
rect 23034 30037 23068 30071
rect 22830 29969 22864 29996
rect 22830 29962 22861 29969
rect 22861 29962 22864 29969
rect 22932 29962 22966 29996
rect 23034 29969 23068 29996
rect 23034 29962 23037 29969
rect 23037 29962 23068 29969
rect 22830 29901 22864 29921
rect 22830 29887 22861 29901
rect 22861 29887 22864 29901
rect 22932 29887 22966 29921
rect 23034 29901 23068 29921
rect 23034 29887 23037 29901
rect 23037 29887 23068 29901
rect 22830 29833 22864 29846
rect 22830 29812 22861 29833
rect 22861 29812 22864 29833
rect 22932 29812 22966 29846
rect 23034 29833 23068 29846
rect 23034 29812 23037 29833
rect 23037 29812 23068 29833
rect 22830 29765 22864 29771
rect 22830 29737 22861 29765
rect 22861 29737 22864 29765
rect 22932 29737 22966 29771
rect 23034 29765 23068 29771
rect 23034 29737 23037 29765
rect 23037 29737 23068 29765
rect 22842 29663 22861 29693
rect 22861 29663 22876 29693
rect 22842 29659 22876 29663
rect 22842 29595 22861 29621
rect 22861 29595 22876 29621
rect 22842 29587 22876 29595
rect 22842 29527 22861 29549
rect 22861 29527 22876 29549
rect 22842 29515 22876 29527
rect 22842 29459 22861 29477
rect 22861 29459 22876 29477
rect 22842 29443 22876 29459
rect 22842 29391 22861 29405
rect 22861 29391 22876 29405
rect 22842 29371 22876 29391
rect 22842 29323 22861 29333
rect 22861 29323 22876 29333
rect 22842 29299 22876 29323
rect 22842 29255 22861 29261
rect 22861 29255 22876 29261
rect 22842 29227 22876 29255
rect 22842 29187 22861 29189
rect 22861 29187 22876 29189
rect 22842 29155 22876 29187
rect 22842 29085 22876 29117
rect 22842 29083 22861 29085
rect 22861 29083 22876 29085
rect 22842 29017 22876 29045
rect 22842 29011 22861 29017
rect 22861 29011 22876 29017
rect 22842 28949 22876 28973
rect 22842 28939 22861 28949
rect 22861 28939 22876 28949
rect 22842 28881 22876 28901
rect 22842 28867 22861 28881
rect 22861 28867 22876 28881
rect 22842 28813 22876 28829
rect 22842 28795 22861 28813
rect 22861 28795 22876 28813
rect 22842 28745 22876 28757
rect 22842 28723 22861 28745
rect 22861 28723 22876 28745
rect 22842 28677 22876 28685
rect 22842 28651 22861 28677
rect 22861 28651 22876 28677
rect 22842 28609 22876 28613
rect 22842 28579 22861 28609
rect 22861 28579 22876 28609
rect 22842 28507 22861 28541
rect 22861 28507 22876 28541
rect 22842 28439 22861 28469
rect 22861 28439 22876 28469
rect 22842 28435 22876 28439
rect 22842 28371 22861 28397
rect 22861 28371 22876 28397
rect 22842 28363 22876 28371
rect 22842 28303 22861 28325
rect 22861 28303 22876 28325
rect 22842 28291 22876 28303
rect 22842 28235 22861 28253
rect 22861 28235 22876 28253
rect 22842 28219 22876 28235
rect 22842 28167 22861 28181
rect 22861 28167 22876 28181
rect 22842 28147 22876 28167
rect 22842 28099 22861 28109
rect 22861 28099 22876 28109
rect 22842 28075 22876 28099
rect 22842 28031 22861 28037
rect 22861 28031 22876 28037
rect 22842 28003 22876 28031
rect 22842 27963 22861 27965
rect 22861 27963 22876 27965
rect 22842 27931 22876 27963
rect 22842 27861 22876 27893
rect 22842 27859 22861 27861
rect 22861 27859 22876 27861
rect 22842 27793 22876 27821
rect 22842 27787 22861 27793
rect 22861 27787 22876 27793
rect 22842 27725 22876 27749
rect 22842 27715 22861 27725
rect 22861 27715 22876 27725
rect 22842 27657 22876 27677
rect 22842 27643 22861 27657
rect 22861 27643 22876 27657
rect 22842 27589 22876 27605
rect 22842 27571 22861 27589
rect 22861 27571 22876 27589
rect 22842 27521 22876 27533
rect 22842 27499 22861 27521
rect 22861 27499 22876 27521
rect 22842 27453 22876 27461
rect 22842 27427 22861 27453
rect 22861 27427 22876 27453
rect 22842 27385 22876 27389
rect 22842 27355 22861 27385
rect 22861 27355 22876 27385
rect 22842 27283 22861 27317
rect 22861 27283 22876 27317
rect 22842 27215 22861 27245
rect 22861 27215 22876 27245
rect 22842 27211 22876 27215
rect 22842 27147 22861 27173
rect 22861 27147 22876 27173
rect 22842 27139 22876 27147
rect 22842 27079 22861 27101
rect 22861 27079 22876 27101
rect 22842 27067 22876 27079
rect 22842 27011 22861 27029
rect 22861 27011 22876 27029
rect 22842 26995 22876 27011
rect 22842 26943 22861 26957
rect 22861 26943 22876 26957
rect 22842 26923 22876 26943
rect 22842 26875 22861 26885
rect 22861 26875 22876 26885
rect 22842 26851 22876 26875
rect 22842 26807 22861 26813
rect 22861 26807 22876 26813
rect 22842 26779 22876 26807
rect 22842 26739 22861 26741
rect 22861 26739 22876 26741
rect 22842 26707 22876 26739
rect 22842 26637 22876 26669
rect 22842 26635 22861 26637
rect 22861 26635 22876 26637
rect 22842 26569 22876 26597
rect 22842 26563 22861 26569
rect 22861 26563 22876 26569
rect 22842 26501 22876 26525
rect 22842 26491 22861 26501
rect 22861 26491 22876 26501
rect 22842 26433 22876 26453
rect 22842 26419 22861 26433
rect 22861 26419 22876 26433
rect 22842 26365 22876 26381
rect 22842 26347 22861 26365
rect 22861 26347 22876 26365
rect 22842 26297 22876 26309
rect 22842 26275 22861 26297
rect 22861 26275 22876 26297
rect 22842 26229 22876 26237
rect 22842 26203 22861 26229
rect 22861 26203 22876 26229
rect 22842 26161 22876 26165
rect 22842 26131 22861 26161
rect 22861 26131 22876 26161
rect 22842 26059 22861 26093
rect 22861 26059 22876 26093
rect 22842 25991 22861 26021
rect 22861 25991 22876 26021
rect 22842 25987 22876 25991
rect 22842 25923 22861 25949
rect 22861 25923 22876 25949
rect 22842 25915 22876 25923
rect 22842 25855 22861 25877
rect 22861 25855 22876 25877
rect 22842 25843 22876 25855
rect 22842 25787 22861 25805
rect 22861 25787 22876 25805
rect 22842 25771 22876 25787
rect 22842 25719 22861 25733
rect 22861 25719 22876 25733
rect 22842 25699 22876 25719
rect 22842 25651 22861 25661
rect 22861 25651 22876 25661
rect 22842 25627 22876 25651
rect 22842 25583 22861 25589
rect 22861 25583 22876 25589
rect 22842 25555 22876 25583
rect 22842 25515 22861 25517
rect 22861 25515 22876 25517
rect 22842 25483 22876 25515
rect 22842 25413 22876 25445
rect 22842 25411 22861 25413
rect 22861 25411 22876 25413
rect 22842 25345 22876 25373
rect 22842 25339 22861 25345
rect 22861 25339 22876 25345
rect 22842 25277 22876 25300
rect 22842 25266 22861 25277
rect 22861 25266 22876 25277
rect 22842 25209 22876 25227
rect 22842 25193 22861 25209
rect 22861 25193 22876 25209
rect 22842 25140 22876 25154
rect 22842 25120 22861 25140
rect 22861 25120 22876 25140
rect 22842 25071 22876 25081
rect 22842 25047 22861 25071
rect 22861 25047 22876 25071
rect 22842 25002 22876 25008
rect 22842 24974 22861 25002
rect 22861 24974 22876 25002
rect 22842 24933 22876 24935
rect 22842 24901 22861 24933
rect 22861 24901 22876 24933
rect 22842 24830 22861 24862
rect 22861 24830 22876 24862
rect 22842 24828 22876 24830
rect 22842 24761 22861 24789
rect 22861 24761 22876 24789
rect 22842 24755 22876 24761
rect 22842 24692 22861 24716
rect 22861 24692 22876 24716
rect 22842 24682 22876 24692
rect 22842 24623 22861 24643
rect 22861 24623 22876 24643
rect 22842 24609 22876 24623
rect 22842 24554 22861 24570
rect 22861 24554 22876 24570
rect 22842 24536 22876 24554
rect 22842 24485 22861 24497
rect 22861 24485 22876 24497
rect 22842 24463 22876 24485
rect 22842 24416 22861 24424
rect 22861 24416 22876 24424
rect 22842 24390 22876 24416
rect 22842 24347 22861 24351
rect 22861 24347 22876 24351
rect 22842 24317 22876 24347
rect 22842 24244 22876 24278
rect 22842 24174 22876 24205
rect 22842 24171 22861 24174
rect 22861 24171 22876 24174
rect 22842 24105 22876 24132
rect 22842 24098 22861 24105
rect 22861 24098 22876 24105
rect 22842 24036 22876 24059
rect 22842 24025 22861 24036
rect 22861 24025 22876 24036
rect 22842 23967 22876 23986
rect 22842 23952 22861 23967
rect 22861 23952 22876 23967
rect 22842 23898 22876 23913
rect 22842 23879 22861 23898
rect 22861 23879 22876 23898
rect 22842 23829 22876 23840
rect 22842 23806 22861 23829
rect 22861 23806 22876 23829
rect 22842 23760 22876 23767
rect 22842 23733 22861 23760
rect 22861 23733 22876 23760
rect 22842 23691 22876 23694
rect 22842 23660 22861 23691
rect 22861 23660 22876 23691
rect 22842 23588 22861 23621
rect 22861 23588 22876 23621
rect 22842 23587 22876 23588
rect 22842 23519 22861 23548
rect 22861 23519 22876 23548
rect 22842 23514 22876 23519
rect 513 23439 524 23463
rect 524 23439 547 23463
rect 590 23439 594 23463
rect 594 23439 624 23463
rect 667 23439 698 23463
rect 698 23439 701 23463
rect 744 23439 768 23463
rect 768 23439 778 23463
rect 821 23439 838 23463
rect 838 23439 855 23463
rect 898 23439 908 23463
rect 908 23439 932 23463
rect 975 23439 978 23463
rect 978 23439 1009 23463
rect 1052 23439 1084 23463
rect 1084 23439 1086 23463
rect 1129 23439 1154 23463
rect 1154 23439 1163 23463
rect 1206 23439 1224 23463
rect 1224 23439 1240 23463
rect 1283 23439 1294 23463
rect 1294 23439 1317 23463
rect 1360 23439 1364 23463
rect 1364 23439 1394 23463
rect 1437 23439 1468 23463
rect 1468 23439 1471 23463
rect 212 23402 246 23436
rect 288 23403 322 23436
rect 364 23403 398 23436
rect 440 23403 474 23436
rect 513 23429 547 23439
rect 590 23429 624 23439
rect 667 23429 701 23439
rect 744 23429 778 23439
rect 821 23429 855 23439
rect 898 23429 932 23439
rect 975 23429 1009 23439
rect 1052 23429 1086 23439
rect 1129 23429 1163 23439
rect 1206 23429 1240 23439
rect 1283 23429 1317 23439
rect 1360 23429 1394 23439
rect 1437 23429 1471 23439
rect 288 23402 314 23403
rect 314 23402 322 23403
rect 364 23402 384 23403
rect 384 23402 398 23403
rect 440 23402 454 23403
rect 454 23402 474 23403
rect 513 23369 524 23383
rect 524 23369 547 23383
rect 590 23369 594 23383
rect 594 23369 624 23383
rect 667 23369 698 23383
rect 698 23369 701 23383
rect 744 23369 768 23383
rect 768 23369 778 23383
rect 821 23369 838 23383
rect 838 23369 855 23383
rect 898 23369 908 23383
rect 908 23369 932 23383
rect 975 23369 978 23383
rect 978 23369 1009 23383
rect 1052 23369 1084 23383
rect 1084 23369 1086 23383
rect 1129 23369 1154 23383
rect 1154 23369 1163 23383
rect 1206 23369 1224 23383
rect 1224 23369 1240 23383
rect 1283 23369 1294 23383
rect 1294 23369 1317 23383
rect 1360 23369 1364 23383
rect 1364 23369 1394 23383
rect 1437 23369 1468 23383
rect 1468 23369 1471 23383
rect 212 23330 246 23364
rect 288 23333 322 23364
rect 364 23333 398 23364
rect 440 23333 474 23364
rect 513 23349 547 23369
rect 590 23349 624 23369
rect 667 23349 701 23369
rect 744 23349 778 23369
rect 821 23349 855 23369
rect 898 23349 932 23369
rect 975 23349 1009 23369
rect 1052 23349 1086 23369
rect 1129 23349 1163 23369
rect 1206 23349 1240 23369
rect 1283 23349 1317 23369
rect 1360 23349 1394 23369
rect 1437 23349 1471 23369
rect 288 23330 314 23333
rect 314 23330 322 23333
rect 364 23330 384 23333
rect 384 23330 398 23333
rect 440 23330 454 23333
rect 454 23330 474 23333
rect 513 23299 524 23303
rect 524 23299 547 23303
rect 590 23299 594 23303
rect 594 23299 624 23303
rect 667 23299 698 23303
rect 698 23299 701 23303
rect 744 23299 768 23303
rect 768 23299 778 23303
rect 821 23299 838 23303
rect 838 23299 855 23303
rect 898 23299 908 23303
rect 908 23299 932 23303
rect 975 23299 978 23303
rect 978 23299 1009 23303
rect 1052 23299 1084 23303
rect 1084 23299 1086 23303
rect 1129 23299 1154 23303
rect 1154 23299 1163 23303
rect 1206 23299 1224 23303
rect 1224 23299 1240 23303
rect 1283 23299 1294 23303
rect 1294 23299 1317 23303
rect 1360 23299 1364 23303
rect 1364 23299 1394 23303
rect 1437 23299 1468 23303
rect 1468 23299 1471 23303
rect 212 23258 246 23292
rect 288 23263 322 23292
rect 364 23263 398 23292
rect 440 23263 474 23292
rect 513 23269 547 23299
rect 590 23269 624 23299
rect 667 23269 701 23299
rect 744 23269 778 23299
rect 821 23269 855 23299
rect 898 23269 932 23299
rect 975 23269 1009 23299
rect 1052 23269 1086 23299
rect 1129 23269 1163 23299
rect 1206 23269 1240 23299
rect 1283 23269 1317 23299
rect 1360 23269 1394 23299
rect 1437 23269 1471 23299
rect 288 23258 314 23263
rect 314 23258 322 23263
rect 364 23258 384 23263
rect 384 23258 398 23263
rect 440 23258 454 23263
rect 454 23258 474 23263
rect 212 23186 246 23220
rect 288 23193 322 23220
rect 364 23193 398 23220
rect 440 23193 474 23220
rect 513 23193 547 23223
rect 590 23193 624 23223
rect 667 23193 701 23223
rect 744 23193 778 23223
rect 821 23193 855 23223
rect 898 23193 932 23223
rect 975 23193 1009 23223
rect 1052 23193 1086 23223
rect 1129 23193 1163 23223
rect 1206 23193 1240 23223
rect 1283 23193 1317 23223
rect 1360 23193 1394 23223
rect 1437 23193 1471 23223
rect 288 23186 314 23193
rect 314 23186 322 23193
rect 364 23186 384 23193
rect 384 23186 398 23193
rect 440 23186 454 23193
rect 454 23186 474 23193
rect 513 23189 524 23193
rect 524 23189 547 23193
rect 590 23189 594 23193
rect 594 23189 624 23193
rect 667 23189 698 23193
rect 698 23189 701 23193
rect 744 23189 768 23193
rect 768 23189 778 23193
rect 821 23189 838 23193
rect 838 23189 855 23193
rect 898 23189 908 23193
rect 908 23189 932 23193
rect 975 23189 978 23193
rect 978 23189 1009 23193
rect 1052 23189 1084 23193
rect 1084 23189 1086 23193
rect 1129 23189 1154 23193
rect 1154 23189 1163 23193
rect 1206 23189 1224 23193
rect 1224 23189 1240 23193
rect 1283 23189 1294 23193
rect 1294 23189 1317 23193
rect 1360 23189 1364 23193
rect 1364 23189 1394 23193
rect 1437 23189 1468 23193
rect 1468 23189 1471 23193
rect 22842 23450 22861 23475
rect 22861 23450 22876 23475
rect 22842 23441 22876 23450
rect 22842 23381 22861 23402
rect 22861 23381 22876 23402
rect 22842 23368 22876 23381
rect 22842 23312 22861 23329
rect 22861 23312 22876 23329
rect 22842 23295 22876 23312
rect 22842 23243 22861 23256
rect 22861 23243 22876 23256
rect 22842 23222 22876 23243
rect 212 23114 246 23148
rect 288 23123 322 23148
rect 364 23123 398 23148
rect 440 23123 474 23148
rect 288 23114 314 23123
rect 314 23114 322 23123
rect 364 23114 384 23123
rect 384 23114 398 23123
rect 440 23114 454 23123
rect 454 23114 474 23123
rect 212 23042 246 23076
rect 288 23053 322 23076
rect 364 23053 398 23076
rect 440 23053 474 23076
rect 288 23042 314 23053
rect 314 23042 322 23053
rect 364 23042 384 23053
rect 384 23042 398 23053
rect 440 23042 454 23053
rect 454 23042 474 23053
rect 212 22970 246 23004
rect 288 22983 322 23004
rect 364 22983 398 23004
rect 440 22983 474 23004
rect 288 22970 314 22983
rect 314 22970 322 22983
rect 364 22970 384 22983
rect 384 22970 398 22983
rect 440 22970 454 22983
rect 454 22970 474 22983
rect 212 22898 246 22932
rect 288 22913 322 22932
rect 364 22913 398 22932
rect 440 22913 474 22932
rect 288 22898 314 22913
rect 314 22898 322 22913
rect 364 22898 384 22913
rect 384 22898 398 22913
rect 440 22898 454 22913
rect 454 22898 474 22913
rect 212 22826 246 22860
rect 288 22843 322 22860
rect 364 22843 398 22860
rect 440 22843 474 22860
rect 288 22826 314 22843
rect 314 22826 322 22843
rect 364 22826 384 22843
rect 384 22826 398 22843
rect 440 22826 454 22843
rect 454 22826 474 22843
rect 212 22754 246 22788
rect 288 22773 322 22788
rect 364 22773 398 22788
rect 440 22773 474 22788
rect 288 22754 314 22773
rect 314 22754 322 22773
rect 364 22754 384 22773
rect 384 22754 398 22773
rect 440 22754 454 22773
rect 454 22754 474 22773
rect 212 22681 246 22715
rect 288 22702 322 22715
rect 364 22702 398 22715
rect 440 22702 474 22715
rect 288 22681 314 22702
rect 314 22681 322 22702
rect 364 22681 384 22702
rect 384 22681 398 22702
rect 440 22681 454 22702
rect 454 22681 474 22702
rect 212 22608 246 22642
rect 288 22631 322 22642
rect 364 22631 398 22642
rect 440 22631 474 22642
rect 288 22608 314 22631
rect 314 22608 322 22631
rect 364 22608 384 22631
rect 384 22608 398 22631
rect 440 22608 454 22631
rect 454 22608 474 22631
rect 212 22535 246 22569
rect 288 22560 322 22569
rect 364 22560 398 22569
rect 440 22560 474 22569
rect 288 22535 314 22560
rect 314 22535 322 22560
rect 364 22535 384 22560
rect 384 22535 398 22560
rect 440 22535 454 22560
rect 454 22535 474 22560
rect 649 22455 664 22482
rect 664 22455 683 22482
rect 729 22455 734 22482
rect 734 22455 763 22482
rect 809 22455 838 22482
rect 838 22455 843 22482
rect 889 22455 908 22482
rect 908 22455 923 22482
rect 969 22455 978 22482
rect 978 22455 1003 22482
rect 649 22448 683 22455
rect 729 22448 763 22455
rect 809 22448 843 22455
rect 889 22448 923 22455
rect 969 22448 1003 22455
rect 1049 22448 1083 22482
rect 649 22384 664 22410
rect 664 22384 683 22410
rect 729 22384 734 22410
rect 734 22384 763 22410
rect 809 22384 838 22410
rect 838 22384 843 22410
rect 889 22384 908 22410
rect 908 22384 923 22410
rect 969 22384 978 22410
rect 978 22384 1003 22410
rect 649 22376 683 22384
rect 729 22376 763 22384
rect 809 22376 843 22384
rect 889 22376 923 22384
rect 969 22376 1003 22384
rect 1049 22376 1083 22410
rect 649 22313 664 22338
rect 664 22313 683 22338
rect 729 22313 734 22338
rect 734 22313 763 22338
rect 809 22313 838 22338
rect 838 22313 843 22338
rect 889 22313 908 22338
rect 908 22313 923 22338
rect 969 22313 978 22338
rect 978 22313 1003 22338
rect 649 22304 683 22313
rect 729 22304 763 22313
rect 809 22304 843 22313
rect 889 22304 923 22313
rect 969 22304 1003 22313
rect 1049 22304 1083 22338
rect 22842 23174 22861 23183
rect 22861 23174 22876 23183
rect 22842 23149 22876 23174
rect 22842 23105 22861 23110
rect 22861 23105 22876 23110
rect 22842 23076 22876 23105
rect 22842 23036 22861 23037
rect 22861 23036 22876 23037
rect 22842 23003 22876 23036
rect 22842 22932 22876 22964
rect 22842 22930 22861 22932
rect 22861 22930 22876 22932
rect 22842 22863 22876 22891
rect 22842 22857 22861 22863
rect 22861 22857 22876 22863
rect 22842 22794 22876 22818
rect 22842 22784 22861 22794
rect 22861 22784 22876 22794
rect 22842 22725 22876 22745
rect 22842 22711 22861 22725
rect 22861 22711 22876 22725
rect 22842 22656 22876 22672
rect 22842 22638 22861 22656
rect 22861 22638 22876 22656
rect 22842 22587 22876 22599
rect 22842 22565 22861 22587
rect 22861 22565 22876 22587
rect 22842 22518 22876 22526
rect 22842 22492 22861 22518
rect 22861 22492 22876 22518
rect 22842 22449 22876 22453
rect 22842 22419 22861 22449
rect 22861 22419 22876 22449
rect 22842 22346 22861 22380
rect 22861 22346 22876 22380
rect 649 22232 683 22266
rect 729 22232 763 22266
rect 809 22232 843 22266
rect 889 22232 923 22266
rect 969 22232 1003 22266
rect 1049 22232 1083 22266
rect 649 22160 683 22194
rect 729 22160 763 22194
rect 809 22160 843 22194
rect 889 22160 923 22194
rect 969 22160 1003 22194
rect 1049 22160 1083 22194
rect 649 22088 683 22122
rect 729 22088 763 22122
rect 809 22088 843 22122
rect 889 22088 923 22122
rect 969 22088 1003 22122
rect 1049 22088 1083 22122
rect 22842 22277 22861 22307
rect 22861 22277 22876 22307
rect 22842 22273 22876 22277
rect 22842 22208 22861 22234
rect 22861 22208 22876 22234
rect 22842 22200 22876 22208
rect 22842 22139 22861 22161
rect 22861 22139 22876 22161
rect 22842 22127 22876 22139
rect 649 22016 683 22050
rect 729 22016 763 22050
rect 809 22016 843 22050
rect 889 22016 923 22050
rect 969 22016 1003 22050
rect 1049 22016 1083 22050
rect 649 21944 683 21978
rect 729 21944 763 21978
rect 809 21944 843 21978
rect 889 21944 923 21978
rect 969 21944 1003 21978
rect 1049 21944 1083 21978
rect 649 21872 683 21906
rect 729 21872 763 21906
rect 809 21872 843 21906
rect 889 21872 923 21906
rect 969 21872 1003 21906
rect 1049 21872 1083 21906
rect 649 21800 683 21834
rect 729 21800 763 21834
rect 809 21800 843 21834
rect 889 21800 923 21834
rect 969 21800 1003 21834
rect 1049 21800 1083 21834
rect 649 21728 683 21762
rect 729 21728 763 21762
rect 809 21728 843 21762
rect 889 21728 923 21762
rect 969 21728 1003 21762
rect 1049 21728 1083 21762
rect 649 21656 683 21690
rect 729 21656 763 21690
rect 809 21656 843 21690
rect 889 21656 923 21690
rect 969 21656 1003 21690
rect 1049 21656 1083 21690
rect 649 21584 683 21618
rect 729 21584 763 21618
rect 809 21584 843 21618
rect 889 21584 923 21618
rect 969 21584 1003 21618
rect 1049 21584 1083 21618
rect 649 21512 683 21546
rect 729 21512 763 21546
rect 809 21512 843 21546
rect 889 21512 923 21546
rect 969 21512 1003 21546
rect 1049 21512 1083 21546
rect 649 21440 683 21474
rect 729 21440 763 21474
rect 809 21440 843 21474
rect 889 21440 923 21474
rect 969 21440 1003 21474
rect 1049 21440 1083 21474
rect 649 21368 683 21402
rect 729 21368 763 21402
rect 809 21368 843 21402
rect 889 21368 923 21402
rect 969 21368 1003 21402
rect 1049 21368 1083 21402
rect 649 21296 683 21330
rect 729 21296 763 21330
rect 809 21296 843 21330
rect 889 21296 923 21330
rect 969 21296 1003 21330
rect 1049 21296 1083 21330
rect 649 21224 683 21258
rect 729 21224 763 21258
rect 809 21224 843 21258
rect 889 21224 923 21258
rect 969 21224 1003 21258
rect 1049 21224 1083 21258
rect 649 21152 683 21186
rect 729 21152 763 21186
rect 809 21152 843 21186
rect 889 21152 923 21186
rect 969 21152 1003 21186
rect 1049 21152 1083 21186
rect 649 21080 683 21114
rect 729 21080 763 21114
rect 809 21080 843 21114
rect 889 21080 923 21114
rect 969 21080 1003 21114
rect 1049 21080 1083 21114
rect 649 21008 683 21042
rect 729 21008 763 21042
rect 809 21008 843 21042
rect 889 21008 923 21042
rect 969 21008 1003 21042
rect 1049 21008 1083 21042
rect 649 20936 683 20970
rect 729 20936 763 20970
rect 809 20936 843 20970
rect 889 20936 923 20970
rect 969 20936 1003 20970
rect 1049 20936 1083 20970
rect 649 20864 683 20898
rect 729 20864 763 20898
rect 809 20864 843 20898
rect 889 20864 923 20898
rect 969 20864 1003 20898
rect 1049 20864 1083 20898
rect 649 20792 683 20826
rect 729 20792 763 20826
rect 809 20792 843 20826
rect 889 20792 923 20826
rect 969 20792 1003 20826
rect 1049 20792 1083 20826
rect 649 20720 683 20754
rect 729 20720 763 20754
rect 809 20720 843 20754
rect 889 20720 923 20754
rect 969 20720 1003 20754
rect 1049 20720 1083 20754
rect 649 20648 683 20682
rect 729 20648 763 20682
rect 809 20648 843 20682
rect 889 20648 923 20682
rect 969 20648 1003 20682
rect 1049 20648 1083 20682
rect 649 20576 683 20610
rect 729 20576 763 20610
rect 809 20576 843 20610
rect 889 20576 923 20610
rect 969 20576 1003 20610
rect 1049 20576 1083 20610
rect 649 20504 683 20538
rect 729 20504 763 20538
rect 809 20504 843 20538
rect 889 20504 923 20538
rect 969 20504 1003 20538
rect 1049 20504 1083 20538
rect 649 20432 683 20466
rect 729 20432 763 20466
rect 809 20432 843 20466
rect 889 20432 923 20466
rect 969 20432 1003 20466
rect 1049 20432 1083 20466
rect 2377 20516 2411 20538
rect 2453 20516 2487 20538
rect 2529 20516 2563 20538
rect 2605 20516 2639 20538
rect 2680 20516 2714 20538
rect 2755 20516 2789 20538
rect 2830 20516 2864 20538
rect 2905 20516 2939 20538
rect 2980 20516 3014 20538
rect 3055 20516 3089 20538
rect 3130 20516 3164 20538
rect 2377 20504 2401 20516
rect 2401 20504 2411 20516
rect 2453 20504 2474 20516
rect 2474 20504 2487 20516
rect 2529 20504 2547 20516
rect 2547 20504 2563 20516
rect 2605 20504 2620 20516
rect 2620 20504 2639 20516
rect 2680 20504 2693 20516
rect 2693 20504 2714 20516
rect 2755 20504 2766 20516
rect 2766 20504 2789 20516
rect 2830 20504 2839 20516
rect 2839 20504 2864 20516
rect 2905 20504 2912 20516
rect 2912 20504 2939 20516
rect 2980 20504 2984 20516
rect 2984 20504 3014 20516
rect 3055 20504 3056 20516
rect 3056 20504 3089 20516
rect 3130 20504 3162 20516
rect 3162 20504 3164 20516
rect 2377 20438 2411 20452
rect 2453 20438 2487 20452
rect 2529 20438 2563 20452
rect 2605 20438 2639 20452
rect 2680 20438 2714 20452
rect 2755 20438 2789 20452
rect 2830 20438 2864 20452
rect 2905 20438 2939 20452
rect 2980 20438 3014 20452
rect 3055 20438 3089 20452
rect 3130 20438 3164 20452
rect 2377 20418 2401 20438
rect 2401 20418 2411 20438
rect 2453 20418 2474 20438
rect 2474 20418 2487 20438
rect 2529 20418 2547 20438
rect 2547 20418 2563 20438
rect 2605 20418 2620 20438
rect 2620 20418 2639 20438
rect 2680 20418 2693 20438
rect 2693 20418 2714 20438
rect 2755 20418 2766 20438
rect 2766 20418 2789 20438
rect 2830 20418 2839 20438
rect 2839 20418 2864 20438
rect 2905 20418 2912 20438
rect 2912 20418 2939 20438
rect 2980 20418 2984 20438
rect 2984 20418 3014 20438
rect 3055 20418 3056 20438
rect 3056 20418 3089 20438
rect 3130 20418 3162 20438
rect 3162 20418 3164 20438
rect 649 20360 683 20394
rect 729 20360 763 20394
rect 809 20360 843 20394
rect 889 20360 923 20394
rect 969 20360 1003 20394
rect 1049 20360 1083 20394
rect 649 20288 683 20322
rect 729 20288 763 20322
rect 809 20288 843 20322
rect 889 20288 923 20322
rect 969 20288 1003 20322
rect 1049 20288 1083 20322
rect 649 20216 683 20250
rect 729 20216 763 20250
rect 809 20216 843 20250
rect 889 20216 923 20250
rect 969 20216 1003 20250
rect 1049 20216 1083 20250
rect 649 20144 683 20178
rect 729 20144 763 20178
rect 809 20144 843 20178
rect 889 20144 923 20178
rect 969 20144 1003 20178
rect 1049 20144 1083 20178
rect 649 20072 683 20106
rect 729 20072 763 20106
rect 809 20072 843 20106
rect 889 20072 923 20106
rect 969 20072 1003 20106
rect 1049 20072 1083 20106
rect 649 20000 683 20034
rect 729 20000 763 20034
rect 809 20000 843 20034
rect 889 20000 923 20034
rect 969 20000 1003 20034
rect 1049 20000 1083 20034
rect 26921 20405 26955 20439
rect 27003 20405 27037 20439
rect 26921 20328 26955 20362
rect 27003 20328 27037 20362
rect 26405 20226 26439 20260
rect 26481 20258 26511 20260
rect 26511 20258 26515 20260
rect 26557 20258 26581 20260
rect 26581 20258 26591 20260
rect 26633 20258 26651 20260
rect 26651 20258 26667 20260
rect 26709 20258 26721 20260
rect 26721 20258 26743 20260
rect 26785 20258 26791 20260
rect 26791 20258 26819 20260
rect 26861 20258 26895 20260
rect 26481 20226 26515 20258
rect 26557 20226 26591 20258
rect 26633 20226 26667 20258
rect 26709 20226 26743 20258
rect 26785 20226 26819 20258
rect 26861 20226 26895 20258
rect 26937 20226 26971 20260
rect 27012 20226 27046 20260
rect 26405 20142 26439 20176
rect 26481 20150 26515 20176
rect 26557 20150 26591 20176
rect 26633 20150 26667 20176
rect 26709 20150 26743 20176
rect 26785 20150 26819 20176
rect 26861 20150 26895 20176
rect 26481 20142 26511 20150
rect 26511 20142 26515 20150
rect 26557 20142 26581 20150
rect 26581 20142 26591 20150
rect 26633 20142 26651 20150
rect 26651 20142 26667 20150
rect 26709 20142 26721 20150
rect 26721 20142 26743 20150
rect 26785 20142 26791 20150
rect 26791 20142 26819 20150
rect 26861 20142 26895 20150
rect 26937 20142 26971 20176
rect 27012 20142 27046 20176
rect 26405 20058 26439 20092
rect 26481 20078 26515 20092
rect 26557 20078 26591 20092
rect 26633 20078 26667 20092
rect 26709 20078 26743 20092
rect 26785 20078 26819 20092
rect 26861 20078 26895 20092
rect 26481 20058 26511 20078
rect 26511 20058 26515 20078
rect 26557 20058 26581 20078
rect 26581 20058 26591 20078
rect 26633 20058 26651 20078
rect 26651 20058 26667 20078
rect 26709 20058 26721 20078
rect 26721 20058 26743 20078
rect 26785 20058 26791 20078
rect 26791 20058 26819 20078
rect 26861 20058 26895 20078
rect 26937 20058 26971 20092
rect 27012 20058 27046 20092
rect 649 19928 683 19962
rect 729 19928 763 19962
rect 809 19928 843 19962
rect 889 19928 923 19962
rect 969 19928 1003 19962
rect 1049 19928 1083 19962
rect 649 19856 683 19890
rect 729 19856 763 19890
rect 809 19856 843 19890
rect 889 19856 923 19890
rect 969 19856 1003 19890
rect 1049 19856 1083 19890
rect 649 19784 683 19818
rect 729 19784 763 19818
rect 809 19784 843 19818
rect 889 19784 923 19818
rect 969 19784 1003 19818
rect 1049 19784 1083 19818
rect 649 19712 683 19746
rect 729 19712 763 19746
rect 809 19712 843 19746
rect 889 19712 923 19746
rect 969 19712 1003 19746
rect 1049 19712 1083 19746
rect 649 19640 683 19674
rect 729 19640 763 19674
rect 809 19640 843 19674
rect 889 19640 923 19674
rect 969 19640 1003 19674
rect 1049 19640 1083 19674
rect 649 19568 683 19602
rect 729 19568 763 19602
rect 809 19568 843 19602
rect 889 19568 923 19602
rect 969 19568 1003 19602
rect 1049 19568 1083 19602
rect 649 19496 683 19530
rect 729 19496 763 19530
rect 809 19496 843 19530
rect 889 19496 923 19530
rect 969 19496 1003 19530
rect 1049 19496 1083 19530
rect 649 19424 683 19458
rect 729 19424 763 19458
rect 809 19424 843 19458
rect 889 19424 923 19458
rect 969 19424 1003 19458
rect 1049 19424 1083 19458
rect 649 19352 683 19386
rect 729 19352 763 19386
rect 809 19352 843 19386
rect 889 19352 923 19386
rect 969 19352 1003 19386
rect 1049 19352 1083 19386
rect 649 19280 683 19314
rect 729 19280 763 19314
rect 809 19280 843 19314
rect 889 19280 923 19314
rect 969 19280 1003 19314
rect 1049 19280 1083 19314
rect 649 19208 683 19242
rect 729 19208 763 19242
rect 809 19208 843 19242
rect 889 19208 923 19242
rect 969 19208 1003 19242
rect 1049 19208 1083 19242
rect 649 19136 683 19170
rect 729 19136 763 19170
rect 809 19136 843 19170
rect 889 19136 923 19170
rect 969 19136 1003 19170
rect 1049 19136 1083 19170
rect 649 19064 683 19098
rect 729 19064 763 19098
rect 809 19064 843 19098
rect 889 19064 923 19098
rect 969 19064 1003 19098
rect 1049 19064 1083 19098
rect 649 18992 683 19026
rect 729 18992 763 19026
rect 809 18992 843 19026
rect 889 18992 923 19026
rect 969 18992 1003 19026
rect 1049 18992 1083 19026
rect 649 18920 683 18954
rect 729 18920 763 18954
rect 809 18920 843 18954
rect 889 18920 923 18954
rect 969 18920 1003 18954
rect 1049 18920 1083 18954
rect 649 18848 683 18882
rect 729 18848 763 18882
rect 809 18848 843 18882
rect 889 18848 923 18882
rect 969 18848 1003 18882
rect 1049 18848 1083 18882
rect 649 18776 683 18810
rect 729 18776 763 18810
rect 809 18776 843 18810
rect 889 18776 923 18810
rect 969 18776 1003 18810
rect 1049 18776 1083 18810
rect 649 18704 683 18738
rect 729 18704 763 18738
rect 809 18704 843 18738
rect 889 18704 923 18738
rect 969 18704 1003 18738
rect 1049 18704 1083 18738
rect 649 18632 683 18666
rect 729 18632 763 18666
rect 809 18632 843 18666
rect 889 18632 923 18666
rect 969 18632 1003 18666
rect 1049 18632 1083 18666
rect 649 18560 683 18594
rect 729 18560 763 18594
rect 809 18560 843 18594
rect 889 18560 923 18594
rect 969 18560 1003 18594
rect 1049 18560 1083 18594
rect 649 18488 683 18522
rect 729 18488 763 18522
rect 809 18488 843 18522
rect 889 18488 923 18522
rect 969 18488 1003 18522
rect 1049 18488 1083 18522
rect 649 18416 683 18450
rect 729 18416 763 18450
rect 809 18416 843 18450
rect 889 18416 923 18450
rect 969 18416 1003 18450
rect 1049 18416 1083 18450
rect 649 18344 683 18378
rect 729 18344 763 18378
rect 809 18344 843 18378
rect 889 18344 923 18378
rect 969 18344 1003 18378
rect 1049 18344 1083 18378
rect 649 18272 683 18306
rect 729 18272 763 18306
rect 809 18272 843 18306
rect 889 18272 923 18306
rect 969 18272 1003 18306
rect 1049 18272 1083 18306
rect 649 18200 683 18234
rect 729 18200 763 18234
rect 809 18200 843 18234
rect 889 18200 923 18234
rect 969 18200 1003 18234
rect 1049 18200 1083 18234
rect 649 18128 683 18162
rect 729 18128 763 18162
rect 809 18128 843 18162
rect 889 18128 923 18162
rect 969 18128 1003 18162
rect 1049 18128 1083 18162
rect 649 18056 683 18090
rect 729 18056 763 18090
rect 809 18056 843 18090
rect 889 18056 923 18090
rect 969 18056 1003 18090
rect 1049 18056 1083 18090
rect 649 17984 683 18018
rect 729 17984 763 18018
rect 809 17984 843 18018
rect 889 17984 923 18018
rect 969 17984 1003 18018
rect 1049 17984 1083 18018
rect 649 17912 683 17946
rect 729 17912 763 17946
rect 809 17912 843 17946
rect 889 17912 923 17946
rect 969 17912 1003 17946
rect 1049 17912 1083 17946
rect 649 17840 683 17874
rect 729 17840 763 17874
rect 809 17840 843 17874
rect 889 17840 923 17874
rect 969 17840 1003 17874
rect 1049 17840 1083 17874
rect 649 17768 683 17802
rect 729 17768 763 17802
rect 809 17768 843 17802
rect 889 17768 923 17802
rect 969 17768 1003 17802
rect 1049 17768 1083 17802
rect 649 17696 683 17730
rect 729 17696 763 17730
rect 809 17696 843 17730
rect 889 17696 923 17730
rect 969 17696 1003 17730
rect 1049 17696 1083 17730
rect 649 17624 683 17658
rect 729 17624 763 17658
rect 809 17624 843 17658
rect 889 17624 923 17658
rect 969 17624 1003 17658
rect 1049 17624 1083 17658
rect 649 17552 683 17586
rect 729 17552 763 17586
rect 809 17552 843 17586
rect 889 17552 923 17586
rect 969 17552 1003 17586
rect 1049 17552 1083 17586
rect 649 17480 683 17514
rect 729 17480 763 17514
rect 809 17480 843 17514
rect 889 17480 923 17514
rect 969 17480 1003 17514
rect 1049 17480 1083 17514
rect 649 17408 683 17442
rect 729 17419 763 17442
rect 809 17419 843 17442
rect 889 17419 923 17442
rect 969 17419 1003 17442
rect 729 17408 763 17419
rect 809 17408 843 17419
rect 889 17408 923 17419
rect 969 17408 1003 17419
rect 1049 17408 1083 17442
rect 649 17336 683 17370
rect 729 17350 748 17370
rect 748 17350 763 17370
rect 809 17350 816 17370
rect 816 17350 843 17370
rect 889 17350 918 17370
rect 918 17350 923 17370
rect 969 17350 986 17370
rect 986 17350 1003 17370
rect 729 17336 763 17350
rect 809 17336 843 17350
rect 889 17336 923 17350
rect 969 17336 1003 17350
rect 1049 17336 1083 17370
rect 649 17264 683 17298
rect 729 17281 748 17298
rect 748 17281 763 17298
rect 809 17281 816 17298
rect 816 17281 843 17298
rect 889 17281 918 17298
rect 918 17281 923 17298
rect 969 17281 986 17298
rect 986 17281 1003 17298
rect 729 17264 763 17281
rect 809 17264 843 17281
rect 889 17264 923 17281
rect 969 17264 1003 17281
rect 1049 17264 1083 17298
rect 649 17192 683 17226
rect 729 17212 748 17226
rect 748 17212 763 17226
rect 809 17212 816 17226
rect 816 17212 843 17226
rect 889 17212 918 17226
rect 918 17212 923 17226
rect 969 17212 986 17226
rect 986 17212 1003 17226
rect 729 17192 763 17212
rect 809 17192 843 17212
rect 889 17192 923 17212
rect 969 17192 1003 17212
rect 1049 17192 1083 17226
rect 649 17120 683 17154
rect 729 17143 748 17154
rect 748 17143 763 17154
rect 809 17143 816 17154
rect 816 17143 843 17154
rect 889 17143 918 17154
rect 918 17143 923 17154
rect 969 17143 986 17154
rect 986 17143 1003 17154
rect 729 17120 763 17143
rect 809 17120 843 17143
rect 889 17120 923 17143
rect 969 17120 1003 17143
rect 1049 17120 1083 17154
rect 649 17048 683 17082
rect 729 17074 748 17082
rect 748 17074 763 17082
rect 809 17074 816 17082
rect 816 17074 843 17082
rect 889 17074 918 17082
rect 918 17074 923 17082
rect 969 17074 986 17082
rect 986 17074 1003 17082
rect 729 17048 763 17074
rect 809 17048 843 17074
rect 889 17048 923 17074
rect 969 17048 1003 17074
rect 1049 17048 1083 17082
rect 649 16976 683 17010
rect 729 17005 748 17010
rect 748 17005 763 17010
rect 809 17005 816 17010
rect 816 17005 843 17010
rect 889 17005 918 17010
rect 918 17005 923 17010
rect 969 17005 986 17010
rect 986 17005 1003 17010
rect 729 16976 763 17005
rect 809 16976 843 17005
rect 889 16976 923 17005
rect 969 16976 1003 17005
rect 1049 16976 1083 17010
rect 649 16903 683 16937
rect 729 16936 748 16937
rect 748 16936 763 16937
rect 809 16936 816 16937
rect 816 16936 843 16937
rect 889 16936 918 16937
rect 918 16936 923 16937
rect 969 16936 986 16937
rect 986 16936 1003 16937
rect 729 16903 763 16936
rect 809 16903 843 16936
rect 889 16903 923 16936
rect 969 16903 1003 16936
rect 1049 16903 1083 16937
rect 649 16830 683 16864
rect 729 16832 763 16864
rect 809 16832 843 16864
rect 889 16832 923 16864
rect 969 16832 1003 16864
rect 729 16830 748 16832
rect 748 16830 763 16832
rect 809 16830 816 16832
rect 816 16830 843 16832
rect 889 16830 918 16832
rect 918 16830 923 16832
rect 969 16830 986 16832
rect 986 16830 1003 16832
rect 1049 16830 1083 16864
rect 649 16757 683 16791
rect 729 16763 763 16791
rect 809 16763 843 16791
rect 889 16763 923 16791
rect 969 16763 1003 16791
rect 729 16757 748 16763
rect 748 16757 763 16763
rect 809 16757 816 16763
rect 816 16757 843 16763
rect 889 16757 918 16763
rect 918 16757 923 16763
rect 969 16757 986 16763
rect 986 16757 1003 16763
rect 1049 16757 1083 16791
rect 649 16684 683 16718
rect 729 16694 763 16718
rect 809 16694 843 16718
rect 889 16694 923 16718
rect 969 16694 1003 16718
rect 729 16684 748 16694
rect 748 16684 763 16694
rect 809 16684 816 16694
rect 816 16684 843 16694
rect 889 16684 918 16694
rect 918 16684 923 16694
rect 969 16684 986 16694
rect 986 16684 1003 16694
rect 1049 16684 1083 16718
rect 649 16611 683 16645
rect 729 16625 763 16645
rect 809 16625 843 16645
rect 889 16625 923 16645
rect 969 16625 1003 16645
rect 729 16611 748 16625
rect 748 16611 763 16625
rect 809 16611 816 16625
rect 816 16611 843 16625
rect 889 16611 918 16625
rect 918 16611 923 16625
rect 969 16611 986 16625
rect 986 16611 1003 16625
rect 1049 16611 1083 16645
rect 649 16538 683 16572
rect 729 16556 763 16572
rect 809 16556 843 16572
rect 889 16556 923 16572
rect 969 16556 1003 16572
rect 729 16538 748 16556
rect 748 16538 763 16556
rect 809 16538 816 16556
rect 816 16538 843 16556
rect 889 16538 918 16556
rect 918 16538 923 16556
rect 969 16538 986 16556
rect 986 16538 1003 16556
rect 1049 16538 1083 16572
rect 649 16465 683 16499
rect 729 16487 763 16499
rect 809 16487 843 16499
rect 889 16487 923 16499
rect 969 16487 1003 16499
rect 729 16465 748 16487
rect 748 16465 763 16487
rect 809 16465 816 16487
rect 816 16465 843 16487
rect 889 16465 918 16487
rect 918 16465 923 16487
rect 969 16465 986 16487
rect 986 16465 1003 16487
rect 1049 16465 1083 16499
rect 3417 16527 3451 16561
rect 3493 16527 3527 16561
rect 3569 16527 3603 16561
rect 3417 16449 3451 16483
rect 3493 16449 3527 16483
rect 3569 16449 3603 16483
rect 649 16392 683 16426
rect 729 16418 763 16426
rect 809 16418 843 16426
rect 889 16418 923 16426
rect 969 16418 1003 16426
rect 729 16392 748 16418
rect 748 16392 763 16418
rect 809 16392 816 16418
rect 816 16392 843 16418
rect 889 16392 918 16418
rect 918 16392 923 16418
rect 969 16392 986 16418
rect 986 16392 1003 16418
rect 1049 16392 1083 16426
rect 8038 16244 8044 16272
rect 8044 16244 8072 16272
rect 8138 16244 8162 16272
rect 8162 16244 8172 16272
rect 8238 16244 8272 16272
rect 8038 16238 8072 16244
rect 8138 16238 8172 16244
rect 8238 16238 8272 16244
rect 8038 16175 8044 16189
rect 8044 16175 8072 16189
rect 8138 16175 8162 16189
rect 8162 16175 8172 16189
rect 8238 16175 8272 16189
rect 8038 16155 8072 16175
rect 8138 16155 8172 16175
rect 8238 16155 8272 16175
rect 8038 16072 8072 16106
rect 8138 16072 8172 16106
rect 8238 16072 8272 16106
rect 8038 16002 8072 16023
rect 8138 16002 8172 16023
rect 8238 16002 8272 16023
rect 8038 15989 8044 16002
rect 8044 15989 8072 16002
rect 8138 15989 8162 16002
rect 8162 15989 8172 16002
rect 8238 15989 8272 16002
rect 8038 15933 8072 15939
rect 8138 15933 8172 15939
rect 8238 15933 8272 15939
rect 8038 15905 8044 15933
rect 8044 15905 8072 15933
rect 8138 15905 8162 15933
rect 8162 15905 8172 15933
rect 8238 15905 8272 15933
rect 8038 15830 8044 15855
rect 8044 15830 8072 15855
rect 8138 15830 8162 15855
rect 8162 15830 8172 15855
rect 8238 15830 8272 15855
rect 8038 15821 8072 15830
rect 8138 15821 8172 15830
rect 8238 15821 8272 15830
rect 235 12914 267 12940
rect 267 12914 269 12940
rect 313 12914 335 12940
rect 335 12914 347 12940
rect 391 12914 403 12940
rect 403 12914 425 12940
rect 469 12914 471 12940
rect 471 12914 503 12940
rect 547 12914 573 12940
rect 573 12914 581 12940
rect 625 12914 641 12940
rect 641 12914 659 12940
rect 235 12906 269 12914
rect 313 12906 347 12914
rect 391 12906 425 12914
rect 469 12906 503 12914
rect 547 12906 581 12914
rect 625 12906 659 12914
rect 235 12843 267 12868
rect 267 12843 269 12868
rect 313 12843 335 12868
rect 335 12843 347 12868
rect 391 12843 403 12868
rect 403 12843 425 12868
rect 469 12843 471 12868
rect 471 12843 503 12868
rect 547 12843 573 12868
rect 573 12843 581 12868
rect 625 12843 641 12868
rect 641 12843 659 12868
rect 235 12834 269 12843
rect 313 12834 347 12843
rect 391 12834 425 12843
rect 469 12834 503 12843
rect 547 12834 581 12843
rect 625 12834 659 12843
rect 235 12772 267 12796
rect 267 12772 269 12796
rect 313 12772 335 12796
rect 335 12772 347 12796
rect 391 12772 403 12796
rect 403 12772 425 12796
rect 469 12772 471 12796
rect 471 12772 503 12796
rect 547 12772 573 12796
rect 573 12772 581 12796
rect 625 12772 641 12796
rect 641 12772 659 12796
rect 235 12762 269 12772
rect 313 12762 347 12772
rect 391 12762 425 12772
rect 469 12762 503 12772
rect 547 12762 581 12772
rect 625 12762 659 12772
rect 235 12701 267 12724
rect 267 12701 269 12724
rect 313 12701 335 12724
rect 335 12701 347 12724
rect 391 12701 403 12724
rect 403 12701 425 12724
rect 469 12701 471 12724
rect 471 12701 503 12724
rect 547 12701 573 12724
rect 573 12701 581 12724
rect 625 12701 641 12724
rect 641 12701 659 12724
rect 235 12690 269 12701
rect 313 12690 347 12701
rect 391 12690 425 12701
rect 469 12690 503 12701
rect 547 12690 581 12701
rect 625 12690 659 12701
rect 235 12630 267 12652
rect 267 12630 269 12652
rect 313 12630 335 12652
rect 335 12630 347 12652
rect 391 12630 403 12652
rect 403 12630 425 12652
rect 469 12630 471 12652
rect 471 12630 503 12652
rect 547 12630 573 12652
rect 573 12630 581 12652
rect 625 12630 641 12652
rect 641 12630 659 12652
rect 235 12618 269 12630
rect 313 12618 347 12630
rect 391 12618 425 12630
rect 469 12618 503 12630
rect 547 12618 581 12630
rect 625 12618 659 12630
rect 235 12559 267 12579
rect 267 12559 269 12579
rect 313 12559 335 12579
rect 335 12559 347 12579
rect 391 12559 403 12579
rect 403 12559 425 12579
rect 469 12559 471 12579
rect 471 12559 503 12579
rect 547 12559 573 12579
rect 573 12559 581 12579
rect 625 12559 641 12579
rect 641 12559 659 12579
rect 235 12545 269 12559
rect 313 12545 347 12559
rect 391 12545 425 12559
rect 469 12545 503 12559
rect 547 12545 581 12559
rect 625 12545 659 12559
rect 235 12488 267 12506
rect 267 12488 269 12506
rect 313 12488 335 12506
rect 335 12488 347 12506
rect 391 12488 403 12506
rect 403 12488 425 12506
rect 469 12488 471 12506
rect 471 12488 503 12506
rect 547 12488 573 12506
rect 573 12488 581 12506
rect 625 12488 641 12506
rect 641 12488 659 12506
rect 235 12472 269 12488
rect 313 12472 347 12488
rect 391 12472 425 12488
rect 469 12472 503 12488
rect 547 12472 581 12488
rect 625 12472 659 12488
rect 236 12380 270 12413
rect 309 12380 343 12413
rect 382 12380 416 12413
rect 455 12380 489 12413
rect 527 12380 561 12413
rect 599 12380 633 12413
rect 671 12380 705 12413
rect 236 12379 267 12380
rect 267 12379 270 12380
rect 309 12379 335 12380
rect 335 12379 343 12380
rect 382 12379 403 12380
rect 403 12379 416 12380
rect 455 12379 471 12380
rect 471 12379 489 12380
rect 527 12379 539 12380
rect 539 12379 561 12380
rect 599 12379 607 12380
rect 607 12379 633 12380
rect 671 12379 675 12380
rect 675 12379 705 12380
rect 743 12379 777 12413
rect 815 12380 849 12413
rect 887 12380 921 12413
rect 959 12380 993 12413
rect 1031 12380 1065 12413
rect 1103 12380 1137 12413
rect 1175 12380 1209 12413
rect 815 12379 845 12380
rect 845 12379 849 12380
rect 887 12379 913 12380
rect 913 12379 921 12380
rect 959 12379 981 12380
rect 981 12379 993 12380
rect 1031 12379 1049 12380
rect 1049 12379 1065 12380
rect 1103 12379 1117 12380
rect 1117 12379 1137 12380
rect 1175 12379 1185 12380
rect 1185 12379 1209 12380
rect 236 12309 270 12339
rect 309 12309 343 12339
rect 382 12309 416 12339
rect 455 12309 489 12339
rect 527 12309 561 12339
rect 599 12309 633 12339
rect 671 12309 705 12339
rect 236 12305 267 12309
rect 267 12305 270 12309
rect 309 12305 335 12309
rect 335 12305 343 12309
rect 382 12305 403 12309
rect 403 12305 416 12309
rect 455 12305 471 12309
rect 471 12305 489 12309
rect 527 12305 539 12309
rect 539 12305 561 12309
rect 599 12305 607 12309
rect 607 12305 633 12309
rect 671 12305 675 12309
rect 675 12305 705 12309
rect 743 12305 777 12339
rect 815 12309 849 12339
rect 887 12309 921 12339
rect 959 12309 993 12339
rect 1031 12309 1065 12339
rect 1103 12309 1137 12339
rect 1175 12309 1209 12339
rect 815 12305 845 12309
rect 845 12305 849 12309
rect 887 12305 913 12309
rect 913 12305 921 12309
rect 959 12305 981 12309
rect 981 12305 993 12309
rect 1031 12305 1049 12309
rect 1049 12305 1065 12309
rect 1103 12305 1117 12309
rect 1117 12305 1137 12309
rect 1175 12305 1185 12309
rect 1185 12305 1209 12309
rect 236 12238 270 12265
rect 309 12238 343 12265
rect 382 12238 416 12265
rect 455 12238 489 12265
rect 527 12238 561 12265
rect 599 12238 633 12265
rect 671 12238 705 12265
rect 236 12231 267 12238
rect 267 12231 270 12238
rect 309 12231 335 12238
rect 335 12231 343 12238
rect 382 12231 403 12238
rect 403 12231 416 12238
rect 455 12231 471 12238
rect 471 12231 489 12238
rect 527 12231 539 12238
rect 539 12231 561 12238
rect 599 12231 607 12238
rect 607 12231 633 12238
rect 671 12231 675 12238
rect 675 12231 705 12238
rect 743 12231 777 12265
rect 815 12238 849 12265
rect 887 12238 921 12265
rect 959 12238 993 12265
rect 1031 12238 1065 12265
rect 1103 12238 1137 12265
rect 1175 12238 1209 12265
rect 815 12231 845 12238
rect 845 12231 849 12238
rect 887 12231 913 12238
rect 913 12231 921 12238
rect 959 12231 981 12238
rect 981 12231 993 12238
rect 1031 12231 1049 12238
rect 1049 12231 1065 12238
rect 1103 12231 1117 12238
rect 1117 12231 1137 12238
rect 1175 12231 1185 12238
rect 1185 12231 1209 12238
rect 236 12167 270 12191
rect 309 12167 343 12191
rect 382 12167 416 12191
rect 455 12167 489 12191
rect 527 12167 561 12191
rect 599 12167 633 12191
rect 671 12167 705 12191
rect 236 12157 267 12167
rect 267 12157 270 12167
rect 309 12157 335 12167
rect 335 12157 343 12167
rect 382 12157 403 12167
rect 403 12157 416 12167
rect 455 12157 471 12167
rect 471 12157 489 12167
rect 527 12157 539 12167
rect 539 12157 561 12167
rect 599 12157 607 12167
rect 607 12157 633 12167
rect 671 12157 675 12167
rect 675 12157 705 12167
rect 743 12157 777 12191
rect 815 12167 849 12191
rect 887 12167 921 12191
rect 959 12167 993 12191
rect 1031 12167 1065 12191
rect 1103 12167 1137 12191
rect 1175 12167 1209 12191
rect 815 12157 845 12167
rect 845 12157 849 12167
rect 887 12157 913 12167
rect 913 12157 921 12167
rect 959 12157 981 12167
rect 981 12157 993 12167
rect 1031 12157 1049 12167
rect 1049 12157 1065 12167
rect 1103 12157 1117 12167
rect 1117 12157 1137 12167
rect 1175 12157 1185 12167
rect 1185 12157 1209 12167
rect 236 12096 270 12117
rect 309 12096 343 12117
rect 382 12096 416 12117
rect 455 12096 489 12117
rect 527 12096 561 12117
rect 599 12096 633 12117
rect 671 12096 705 12117
rect 236 12083 267 12096
rect 267 12083 270 12096
rect 309 12083 335 12096
rect 335 12083 343 12096
rect 382 12083 403 12096
rect 403 12083 416 12096
rect 455 12083 471 12096
rect 471 12083 489 12096
rect 527 12083 539 12096
rect 539 12083 561 12096
rect 599 12083 607 12096
rect 607 12083 633 12096
rect 671 12083 675 12096
rect 675 12083 705 12096
rect 743 12083 777 12117
rect 815 12096 849 12117
rect 887 12096 921 12117
rect 959 12096 993 12117
rect 1031 12096 1065 12117
rect 1103 12096 1137 12117
rect 1175 12096 1209 12117
rect 815 12083 845 12096
rect 845 12083 849 12096
rect 887 12083 913 12096
rect 913 12083 921 12096
rect 959 12083 981 12096
rect 981 12083 993 12096
rect 1031 12083 1049 12096
rect 1049 12083 1065 12096
rect 1103 12083 1117 12096
rect 1117 12083 1137 12096
rect 1175 12083 1185 12096
rect 1185 12083 1209 12096
rect 236 12025 270 12043
rect 309 12025 343 12043
rect 382 12025 416 12043
rect 455 12025 489 12043
rect 527 12025 561 12043
rect 599 12025 633 12043
rect 671 12025 705 12043
rect 236 12009 267 12025
rect 267 12009 270 12025
rect 309 12009 335 12025
rect 335 12009 343 12025
rect 382 12009 403 12025
rect 403 12009 416 12025
rect 455 12009 471 12025
rect 471 12009 489 12025
rect 527 12009 539 12025
rect 539 12009 561 12025
rect 599 12009 607 12025
rect 607 12009 633 12025
rect 671 12009 675 12025
rect 675 12009 705 12025
rect 743 12009 777 12043
rect 815 12025 849 12043
rect 887 12025 921 12043
rect 959 12025 993 12043
rect 1031 12025 1065 12043
rect 1103 12025 1137 12043
rect 1175 12025 1209 12043
rect 815 12009 845 12025
rect 845 12009 849 12025
rect 887 12009 913 12025
rect 913 12009 921 12025
rect 959 12009 981 12025
rect 981 12009 993 12025
rect 1031 12009 1049 12025
rect 1049 12009 1065 12025
rect 1103 12009 1117 12025
rect 1117 12009 1137 12025
rect 1175 12009 1185 12025
rect 1185 12009 1209 12025
rect 236 11954 270 11969
rect 309 11954 343 11969
rect 382 11954 416 11969
rect 455 11954 489 11969
rect 527 11954 561 11969
rect 599 11954 633 11969
rect 671 11954 705 11969
rect 236 11935 267 11954
rect 267 11935 270 11954
rect 309 11935 335 11954
rect 335 11935 343 11954
rect 382 11935 403 11954
rect 403 11935 416 11954
rect 455 11935 471 11954
rect 471 11935 489 11954
rect 527 11935 539 11954
rect 539 11935 561 11954
rect 599 11935 607 11954
rect 607 11935 633 11954
rect 671 11935 675 11954
rect 675 11935 705 11954
rect 743 11935 777 11969
rect 815 11954 849 11969
rect 887 11954 921 11969
rect 959 11954 993 11969
rect 1031 11954 1065 11969
rect 1103 11954 1137 11969
rect 1175 11954 1209 11969
rect 815 11935 845 11954
rect 845 11935 849 11954
rect 887 11935 913 11954
rect 913 11935 921 11954
rect 959 11935 981 11954
rect 981 11935 993 11954
rect 1031 11935 1049 11954
rect 1049 11935 1065 11954
rect 1103 11935 1117 11954
rect 1117 11935 1137 11954
rect 1175 11935 1185 11954
rect 1185 11935 1209 11954
rect 236 11883 270 11895
rect 309 11883 343 11895
rect 382 11883 416 11895
rect 455 11883 489 11895
rect 527 11883 561 11895
rect 599 11883 633 11895
rect 671 11883 705 11895
rect 236 11861 267 11883
rect 267 11861 270 11883
rect 309 11861 335 11883
rect 335 11861 343 11883
rect 382 11861 403 11883
rect 403 11861 416 11883
rect 455 11861 471 11883
rect 471 11861 489 11883
rect 527 11861 539 11883
rect 539 11861 561 11883
rect 599 11861 607 11883
rect 607 11861 633 11883
rect 671 11861 675 11883
rect 675 11861 705 11883
rect 743 11861 777 11895
rect 815 11883 849 11895
rect 887 11883 921 11895
rect 959 11883 993 11895
rect 1031 11883 1065 11895
rect 1103 11883 1137 11895
rect 1175 11883 1209 11895
rect 815 11861 845 11883
rect 845 11861 849 11883
rect 887 11861 913 11883
rect 913 11861 921 11883
rect 959 11861 981 11883
rect 981 11861 993 11883
rect 1031 11861 1049 11883
rect 1049 11861 1065 11883
rect 1103 11861 1117 11883
rect 1117 11861 1137 11883
rect 1175 11861 1185 11883
rect 1185 11861 1209 11883
rect 236 11812 270 11821
rect 309 11812 343 11821
rect 382 11812 416 11821
rect 455 11812 489 11821
rect 527 11812 561 11821
rect 599 11812 633 11821
rect 671 11812 705 11821
rect 236 11787 267 11812
rect 267 11787 270 11812
rect 309 11787 335 11812
rect 335 11787 343 11812
rect 382 11787 403 11812
rect 403 11787 416 11812
rect 455 11787 471 11812
rect 471 11787 489 11812
rect 527 11787 539 11812
rect 539 11787 561 11812
rect 599 11787 607 11812
rect 607 11787 633 11812
rect 671 11787 675 11812
rect 675 11787 705 11812
rect 743 11787 777 11821
rect 815 11812 849 11821
rect 887 11812 921 11821
rect 959 11812 993 11821
rect 1031 11812 1065 11821
rect 1103 11812 1137 11821
rect 1175 11812 1209 11821
rect 815 11787 845 11812
rect 845 11787 849 11812
rect 887 11787 913 11812
rect 913 11787 921 11812
rect 959 11787 981 11812
rect 981 11787 993 11812
rect 1031 11787 1049 11812
rect 1049 11787 1065 11812
rect 1103 11787 1117 11812
rect 1117 11787 1137 11812
rect 1175 11787 1185 11812
rect 1185 11787 1209 11812
rect 236 11741 270 11747
rect 309 11741 343 11747
rect 382 11741 416 11747
rect 455 11741 489 11747
rect 527 11741 561 11747
rect 599 11741 633 11747
rect 671 11741 705 11747
rect 236 11713 267 11741
rect 267 11713 270 11741
rect 309 11713 335 11741
rect 335 11713 343 11741
rect 382 11713 403 11741
rect 403 11713 416 11741
rect 455 11713 471 11741
rect 471 11713 489 11741
rect 527 11713 539 11741
rect 539 11713 561 11741
rect 599 11713 607 11741
rect 607 11713 633 11741
rect 671 11713 675 11741
rect 675 11713 705 11741
rect 743 11713 777 11747
rect 815 11741 849 11747
rect 887 11741 921 11747
rect 959 11741 993 11747
rect 1031 11741 1065 11747
rect 1103 11741 1137 11747
rect 1175 11741 1209 11747
rect 815 11713 845 11741
rect 845 11713 849 11741
rect 887 11713 913 11741
rect 913 11713 921 11741
rect 959 11713 981 11741
rect 981 11713 993 11741
rect 1031 11713 1049 11741
rect 1049 11713 1065 11741
rect 1103 11713 1117 11741
rect 1117 11713 1137 11741
rect 1175 11713 1185 11741
rect 1185 11713 1209 11741
rect 236 11670 270 11673
rect 309 11670 343 11673
rect 382 11670 416 11673
rect 455 11670 489 11673
rect 527 11670 561 11673
rect 599 11670 633 11673
rect 671 11670 705 11673
rect 236 11639 267 11670
rect 267 11639 270 11670
rect 309 11639 335 11670
rect 335 11639 343 11670
rect 382 11639 403 11670
rect 403 11639 416 11670
rect 455 11639 471 11670
rect 471 11639 489 11670
rect 527 11639 539 11670
rect 539 11639 561 11670
rect 599 11639 607 11670
rect 607 11639 633 11670
rect 671 11639 675 11670
rect 675 11639 705 11670
rect 743 11639 777 11673
rect 815 11670 849 11673
rect 887 11670 921 11673
rect 959 11670 993 11673
rect 1031 11670 1065 11673
rect 1103 11670 1137 11673
rect 1175 11670 1209 11673
rect 815 11639 845 11670
rect 845 11639 849 11670
rect 887 11639 913 11670
rect 913 11639 921 11670
rect 959 11639 981 11670
rect 981 11639 993 11670
rect 1031 11639 1049 11670
rect 1049 11639 1065 11670
rect 1103 11639 1117 11670
rect 1117 11639 1137 11670
rect 1175 11639 1185 11670
rect 1185 11639 1209 11670
rect 6785 11694 6819 11728
rect 6859 11694 6893 11728
rect 6932 11694 6966 11728
rect 7005 11694 7039 11728
rect 7078 11694 7112 11728
rect 7151 11694 7185 11728
rect 7224 11694 7258 11728
rect 7297 11694 7331 11728
rect 7370 11694 7404 11728
rect 7443 11694 7477 11728
rect 7516 11694 7550 11728
rect 7589 11694 7623 11728
rect 7662 11694 7696 11728
rect 6785 11622 6819 11656
rect 6859 11622 6893 11656
rect 6932 11622 6966 11656
rect 7005 11622 7039 11656
rect 7078 11622 7112 11656
rect 7151 11622 7185 11656
rect 7224 11622 7258 11656
rect 7297 11622 7331 11656
rect 7370 11622 7404 11656
rect 7443 11622 7477 11656
rect 7516 11622 7550 11656
rect 7589 11622 7623 11656
rect 7662 11622 7696 11656
rect 236 11598 270 11599
rect 309 11598 343 11599
rect 382 11598 416 11599
rect 455 11598 489 11599
rect 527 11598 561 11599
rect 599 11598 633 11599
rect 671 11598 705 11599
rect 236 11565 267 11598
rect 267 11565 270 11598
rect 309 11565 335 11598
rect 335 11565 343 11598
rect 382 11565 403 11598
rect 403 11565 416 11598
rect 455 11565 471 11598
rect 471 11565 489 11598
rect 527 11565 539 11598
rect 539 11565 561 11598
rect 599 11565 607 11598
rect 607 11565 633 11598
rect 671 11565 675 11598
rect 675 11565 705 11598
rect 743 11565 777 11599
rect 815 11598 849 11599
rect 887 11598 921 11599
rect 959 11598 993 11599
rect 1031 11598 1065 11599
rect 1103 11598 1137 11599
rect 1175 11598 1209 11599
rect 815 11565 845 11598
rect 845 11565 849 11598
rect 887 11565 913 11598
rect 913 11565 921 11598
rect 959 11565 981 11598
rect 981 11565 993 11598
rect 1031 11565 1049 11598
rect 1049 11565 1065 11598
rect 1103 11565 1117 11598
rect 1117 11565 1137 11598
rect 1175 11565 1185 11598
rect 1185 11565 1209 11598
rect 236 11492 267 11525
rect 267 11492 270 11525
rect 309 11492 335 11525
rect 335 11492 343 11525
rect 382 11492 403 11525
rect 403 11492 416 11525
rect 455 11492 471 11525
rect 471 11492 489 11525
rect 527 11492 539 11525
rect 539 11492 561 11525
rect 599 11492 607 11525
rect 607 11492 633 11525
rect 671 11492 675 11525
rect 675 11492 705 11525
rect 236 11491 270 11492
rect 309 11491 343 11492
rect 382 11491 416 11492
rect 455 11491 489 11492
rect 527 11491 561 11492
rect 599 11491 633 11492
rect 671 11491 705 11492
rect 743 11491 777 11525
rect 815 11492 845 11525
rect 845 11492 849 11525
rect 887 11492 913 11525
rect 913 11492 921 11525
rect 959 11492 981 11525
rect 981 11492 993 11525
rect 1031 11492 1049 11525
rect 1049 11492 1065 11525
rect 1103 11492 1117 11525
rect 1117 11492 1137 11525
rect 1175 11492 1185 11525
rect 1185 11492 1209 11525
rect 815 11491 849 11492
rect 887 11491 921 11492
rect 959 11491 993 11492
rect 1031 11491 1065 11492
rect 1103 11491 1137 11492
rect 1175 11491 1209 11492
rect 17445 11588 17451 11617
rect 17451 11588 17479 11617
rect 17525 11588 17555 11617
rect 17555 11588 17559 11617
rect 17605 11588 17624 11617
rect 17624 11588 17639 11617
rect 17684 11588 17693 11617
rect 17693 11588 17718 11617
rect 17763 11588 17796 11617
rect 17796 11588 17797 11617
rect 17842 11588 17865 11617
rect 17865 11588 17876 11617
rect 17921 11588 17934 11617
rect 17934 11588 17955 11617
rect 18000 11588 18003 11617
rect 18003 11588 18034 11617
rect 18079 11588 18107 11617
rect 18107 11588 18113 11617
rect 18158 11588 18176 11617
rect 18176 11588 18192 11617
rect 18500 11588 18521 11615
rect 18521 11588 18534 11615
rect 18585 11588 18590 11615
rect 18590 11588 18619 11615
rect 18669 11588 18693 11615
rect 18693 11588 18703 11615
rect 18753 11588 18762 11615
rect 18762 11588 18787 11615
rect 18837 11588 18866 11615
rect 18866 11588 18871 11615
rect 18921 11588 18935 11615
rect 18935 11588 18955 11615
rect 17445 11583 17479 11588
rect 17525 11583 17559 11588
rect 17605 11583 17639 11588
rect 17684 11583 17718 11588
rect 17763 11583 17797 11588
rect 17842 11583 17876 11588
rect 17921 11583 17955 11588
rect 18000 11583 18034 11588
rect 18079 11583 18113 11588
rect 18158 11583 18192 11588
rect 18500 11581 18534 11588
rect 18585 11581 18619 11588
rect 18669 11581 18703 11588
rect 18753 11581 18787 11588
rect 18837 11581 18871 11588
rect 18921 11581 18955 11588
rect 6779 11546 6813 11579
rect 6867 11546 6901 11579
rect 6955 11546 6989 11579
rect 7043 11546 7077 11579
rect 7131 11546 7165 11579
rect 7577 11546 7611 11577
rect 7651 11546 7685 11577
rect 7725 11546 7759 11577
rect 7799 11546 7833 11577
rect 7873 11546 7907 11577
rect 7947 11546 7981 11577
rect 8021 11546 8055 11577
rect 8095 11546 8129 11577
rect 8169 11546 8203 11577
rect 8243 11546 8277 11577
rect 8317 11546 8351 11577
rect 6779 11545 6804 11546
rect 6804 11545 6813 11546
rect 6867 11545 6873 11546
rect 6873 11545 6901 11546
rect 6955 11545 6977 11546
rect 6977 11545 6989 11546
rect 7043 11545 7046 11546
rect 7046 11545 7077 11546
rect 7131 11545 7149 11546
rect 7149 11545 7165 11546
rect 7577 11543 7598 11546
rect 7598 11543 7611 11546
rect 7651 11543 7667 11546
rect 7667 11543 7685 11546
rect 7725 11543 7736 11546
rect 7736 11543 7759 11546
rect 7799 11543 7805 11546
rect 7805 11543 7833 11546
rect 7873 11543 7874 11546
rect 7874 11543 7907 11546
rect 7947 11543 7977 11546
rect 7977 11543 7981 11546
rect 8021 11543 8046 11546
rect 8046 11543 8055 11546
rect 8095 11543 8115 11546
rect 8115 11543 8129 11546
rect 8169 11543 8184 11546
rect 8184 11543 8203 11546
rect 8243 11543 8253 11546
rect 8253 11543 8277 11546
rect 8317 11543 8322 11546
rect 8322 11543 8351 11546
rect 8391 11543 8425 11577
rect 8465 11546 8499 11577
rect 8539 11546 8573 11577
rect 8613 11546 8647 11577
rect 8687 11546 8721 11577
rect 8761 11546 8795 11577
rect 8835 11546 8869 11577
rect 8909 11546 8943 11577
rect 8983 11546 9017 11577
rect 9058 11546 9092 11577
rect 9133 11546 9167 11577
rect 9208 11546 9242 11577
rect 9283 11546 9317 11577
rect 9358 11546 9392 11577
rect 9433 11546 9467 11577
rect 9508 11546 9542 11577
rect 8465 11543 8495 11546
rect 8495 11543 8499 11546
rect 8539 11543 8564 11546
rect 8564 11543 8573 11546
rect 8613 11543 8633 11546
rect 8633 11543 8647 11546
rect 8687 11543 8702 11546
rect 8702 11543 8721 11546
rect 8761 11543 8771 11546
rect 8771 11543 8795 11546
rect 8835 11543 8840 11546
rect 8840 11543 8869 11546
rect 8909 11543 8943 11546
rect 8983 11543 9012 11546
rect 9012 11543 9017 11546
rect 9058 11543 9080 11546
rect 9080 11543 9092 11546
rect 9133 11543 9148 11546
rect 9148 11543 9167 11546
rect 9208 11543 9216 11546
rect 9216 11543 9242 11546
rect 9283 11543 9284 11546
rect 9284 11543 9317 11546
rect 9358 11543 9386 11546
rect 9386 11543 9392 11546
rect 9433 11543 9454 11546
rect 9454 11543 9467 11546
rect 9508 11543 9522 11546
rect 9522 11543 9542 11546
rect 6779 11474 6813 11507
rect 6867 11474 6901 11507
rect 6955 11474 6989 11507
rect 7043 11474 7077 11507
rect 7131 11474 7165 11507
rect 7577 11474 7611 11489
rect 7651 11474 7685 11489
rect 7725 11474 7759 11489
rect 7799 11474 7833 11489
rect 7873 11474 7907 11489
rect 7947 11474 7981 11489
rect 8021 11474 8055 11489
rect 8095 11474 8129 11489
rect 8169 11474 8203 11489
rect 8243 11474 8277 11489
rect 8317 11474 8351 11489
rect 6779 11473 6804 11474
rect 6804 11473 6813 11474
rect 6867 11473 6873 11474
rect 6873 11473 6901 11474
rect 6955 11473 6977 11474
rect 6977 11473 6989 11474
rect 7043 11473 7046 11474
rect 7046 11473 7077 11474
rect 7131 11473 7149 11474
rect 7149 11473 7165 11474
rect 7577 11455 7598 11474
rect 7598 11455 7611 11474
rect 7651 11455 7667 11474
rect 7667 11455 7685 11474
rect 7725 11455 7736 11474
rect 7736 11455 7759 11474
rect 7799 11455 7805 11474
rect 7805 11455 7833 11474
rect 7873 11455 7874 11474
rect 7874 11455 7907 11474
rect 7947 11455 7977 11474
rect 7977 11455 7981 11474
rect 8021 11455 8046 11474
rect 8046 11455 8055 11474
rect 8095 11455 8115 11474
rect 8115 11455 8129 11474
rect 8169 11455 8184 11474
rect 8184 11455 8203 11474
rect 8243 11455 8253 11474
rect 8253 11455 8277 11474
rect 8317 11455 8322 11474
rect 8322 11455 8351 11474
rect 8391 11455 8425 11489
rect 8465 11474 8499 11489
rect 8539 11474 8573 11489
rect 8613 11474 8647 11489
rect 8687 11474 8721 11489
rect 8761 11474 8795 11489
rect 8835 11474 8869 11489
rect 8909 11474 8943 11489
rect 8983 11474 9017 11489
rect 9058 11474 9092 11489
rect 9133 11474 9167 11489
rect 9208 11474 9242 11489
rect 9283 11474 9317 11489
rect 9358 11474 9392 11489
rect 9433 11474 9467 11489
rect 9508 11474 9542 11489
rect 8465 11455 8495 11474
rect 8495 11455 8499 11474
rect 8539 11455 8564 11474
rect 8564 11455 8573 11474
rect 8613 11455 8633 11474
rect 8633 11455 8647 11474
rect 8687 11455 8702 11474
rect 8702 11455 8721 11474
rect 8761 11455 8771 11474
rect 8771 11455 8795 11474
rect 8835 11455 8840 11474
rect 8840 11455 8869 11474
rect 8909 11455 8943 11474
rect 8983 11455 9012 11474
rect 9012 11455 9017 11474
rect 9058 11455 9080 11474
rect 9080 11455 9092 11474
rect 9133 11455 9148 11474
rect 9148 11455 9167 11474
rect 9208 11455 9216 11474
rect 9216 11455 9242 11474
rect 9283 11455 9284 11474
rect 9284 11455 9317 11474
rect 9358 11455 9386 11474
rect 9386 11455 9392 11474
rect 9433 11455 9454 11474
rect 9454 11455 9467 11474
rect 9508 11455 9522 11474
rect 9522 11455 9542 11474
rect 17445 11520 17451 11545
rect 17451 11520 17479 11545
rect 17525 11520 17555 11545
rect 17555 11520 17559 11545
rect 17605 11520 17624 11545
rect 17624 11520 17639 11545
rect 17684 11520 17693 11545
rect 17693 11520 17718 11545
rect 17763 11520 17796 11545
rect 17796 11520 17797 11545
rect 17842 11520 17865 11545
rect 17865 11520 17876 11545
rect 17921 11520 17934 11545
rect 17934 11520 17955 11545
rect 18000 11520 18003 11545
rect 18003 11520 18034 11545
rect 18079 11520 18107 11545
rect 18107 11520 18113 11545
rect 18158 11520 18176 11545
rect 18176 11520 18192 11545
rect 18500 11520 18521 11543
rect 18521 11520 18534 11543
rect 18585 11520 18590 11543
rect 18590 11520 18619 11543
rect 18669 11520 18693 11543
rect 18693 11520 18703 11543
rect 18753 11520 18762 11543
rect 18762 11520 18787 11543
rect 18837 11520 18866 11543
rect 18866 11520 18871 11543
rect 18921 11520 18935 11543
rect 18935 11520 18955 11543
rect 17445 11511 17479 11520
rect 17525 11511 17559 11520
rect 17605 11511 17639 11520
rect 17684 11511 17718 11520
rect 17763 11511 17797 11520
rect 17842 11511 17876 11520
rect 17921 11511 17955 11520
rect 18000 11511 18034 11520
rect 18079 11511 18113 11520
rect 18158 11511 18192 11520
rect 18500 11509 18534 11520
rect 18585 11509 18619 11520
rect 18669 11509 18703 11520
rect 18753 11509 18787 11520
rect 18837 11509 18871 11520
rect 18921 11509 18955 11520
rect 17445 11452 17451 11473
rect 17451 11452 17479 11473
rect 17525 11452 17555 11473
rect 17555 11452 17559 11473
rect 17605 11452 17624 11473
rect 17624 11452 17639 11473
rect 17684 11452 17693 11473
rect 17693 11452 17718 11473
rect 17763 11452 17796 11473
rect 17796 11452 17797 11473
rect 17842 11452 17865 11473
rect 17865 11452 17876 11473
rect 17921 11452 17934 11473
rect 17934 11452 17955 11473
rect 18000 11452 18003 11473
rect 18003 11452 18034 11473
rect 18079 11452 18107 11473
rect 18107 11452 18113 11473
rect 18158 11452 18176 11473
rect 18176 11452 18192 11473
rect 18500 11452 18521 11471
rect 18521 11452 18534 11471
rect 18585 11452 18590 11471
rect 18590 11452 18619 11471
rect 18669 11452 18693 11471
rect 18693 11452 18703 11471
rect 18753 11452 18762 11471
rect 18762 11452 18787 11471
rect 18837 11452 18866 11471
rect 18866 11452 18871 11471
rect 18921 11452 18935 11471
rect 18935 11452 18955 11471
rect 10456 11441 10490 11452
rect 10529 11441 10563 11452
rect 10602 11441 10636 11452
rect 10675 11441 10709 11452
rect 10748 11441 10782 11452
rect 10821 11441 10855 11452
rect 10893 11441 10927 11452
rect 10965 11441 10999 11452
rect 11037 11441 11071 11452
rect 11109 11441 11143 11452
rect 11181 11441 11215 11452
rect 11253 11441 11287 11452
rect 11325 11441 11359 11452
rect 11397 11441 11431 11452
rect 11469 11441 11503 11452
rect 11541 11441 11575 11452
rect 11613 11441 11647 11452
rect 11685 11441 11719 11452
rect 11757 11441 11791 11452
rect 11829 11441 11863 11452
rect 11901 11441 11935 11452
rect 11973 11441 12007 11452
rect 12045 11441 12079 11452
rect 12117 11441 12151 11452
rect 12189 11441 12223 11452
rect 12261 11441 12295 11452
rect 12333 11441 12367 11452
rect 6779 11402 6813 11435
rect 6867 11402 6901 11435
rect 6955 11402 6989 11435
rect 7043 11402 7077 11435
rect 7131 11402 7165 11435
rect 10456 11418 10473 11441
rect 10473 11418 10490 11441
rect 10529 11418 10542 11441
rect 10542 11418 10563 11441
rect 10602 11418 10611 11441
rect 10611 11418 10636 11441
rect 10675 11418 10680 11441
rect 10680 11418 10709 11441
rect 10748 11418 10749 11441
rect 10749 11418 10782 11441
rect 10821 11418 10852 11441
rect 10852 11418 10855 11441
rect 10893 11418 10921 11441
rect 10921 11418 10927 11441
rect 10965 11418 10990 11441
rect 10990 11418 10999 11441
rect 11037 11418 11059 11441
rect 11059 11418 11071 11441
rect 11109 11418 11128 11441
rect 11128 11418 11143 11441
rect 11181 11418 11197 11441
rect 11197 11418 11215 11441
rect 11253 11418 11266 11441
rect 11266 11418 11287 11441
rect 11325 11418 11335 11441
rect 11335 11418 11359 11441
rect 11397 11418 11404 11441
rect 11404 11418 11431 11441
rect 11469 11418 11473 11441
rect 11473 11418 11503 11441
rect 11541 11418 11542 11441
rect 11542 11418 11575 11441
rect 11613 11418 11646 11441
rect 11646 11418 11647 11441
rect 11685 11418 11715 11441
rect 11715 11418 11719 11441
rect 11757 11418 11784 11441
rect 11784 11418 11791 11441
rect 11829 11418 11853 11441
rect 11853 11418 11863 11441
rect 11901 11418 11922 11441
rect 11922 11418 11935 11441
rect 11973 11418 11991 11441
rect 11991 11418 12007 11441
rect 12045 11418 12060 11441
rect 12060 11418 12079 11441
rect 12117 11418 12129 11441
rect 12129 11418 12151 11441
rect 12189 11418 12198 11441
rect 12198 11418 12223 11441
rect 12261 11418 12267 11441
rect 12267 11418 12295 11441
rect 12333 11418 12336 11441
rect 12336 11418 12367 11441
rect 13411 11418 13445 11452
rect 13485 11418 13519 11452
rect 13559 11418 13593 11452
rect 13633 11418 13667 11452
rect 13707 11418 13741 11452
rect 13781 11418 13815 11452
rect 13855 11418 13889 11452
rect 13929 11418 13963 11452
rect 14003 11418 14037 11452
rect 14077 11418 14111 11452
rect 14151 11418 14185 11452
rect 14225 11418 14259 11452
rect 14299 11418 14333 11452
rect 14372 11418 14406 11452
rect 14445 11418 14479 11452
rect 14518 11418 14552 11452
rect 14591 11418 14625 11452
rect 14664 11418 14698 11452
rect 14737 11418 14771 11452
rect 14810 11418 14844 11452
rect 14883 11418 14917 11452
rect 14956 11418 14990 11452
rect 15029 11418 15063 11452
rect 15102 11418 15136 11452
rect 15175 11418 15209 11452
rect 15248 11418 15282 11452
rect 15321 11418 15355 11452
rect 15394 11418 15428 11452
rect 15467 11418 15501 11452
rect 15540 11418 15574 11452
rect 15613 11418 15647 11452
rect 17445 11439 17479 11452
rect 17525 11439 17559 11452
rect 17605 11439 17639 11452
rect 17684 11439 17718 11452
rect 17763 11439 17797 11452
rect 17842 11439 17876 11452
rect 17921 11439 17955 11452
rect 18000 11439 18034 11452
rect 18079 11439 18113 11452
rect 18158 11439 18192 11452
rect 18500 11437 18534 11452
rect 18585 11437 18619 11452
rect 18669 11437 18703 11452
rect 18753 11437 18787 11452
rect 18837 11437 18871 11452
rect 18921 11437 18955 11452
rect 6779 11401 6804 11402
rect 6804 11401 6813 11402
rect 6867 11401 6873 11402
rect 6873 11401 6901 11402
rect 6955 11401 6977 11402
rect 6977 11401 6989 11402
rect 7043 11401 7046 11402
rect 7046 11401 7077 11402
rect 7131 11401 7149 11402
rect 7149 11401 7165 11402
rect 7577 11368 7598 11401
rect 7598 11368 7611 11401
rect 7651 11368 7667 11401
rect 7667 11368 7685 11401
rect 7725 11368 7736 11401
rect 7736 11368 7759 11401
rect 7799 11368 7805 11401
rect 7805 11368 7833 11401
rect 7873 11368 7874 11401
rect 7874 11368 7907 11401
rect 7947 11368 7977 11401
rect 7977 11368 7981 11401
rect 8021 11368 8046 11401
rect 8046 11368 8055 11401
rect 8095 11368 8115 11401
rect 8115 11368 8129 11401
rect 8169 11368 8184 11401
rect 8184 11368 8203 11401
rect 8243 11368 8253 11401
rect 8253 11368 8277 11401
rect 8317 11368 8322 11401
rect 8322 11368 8351 11401
rect 7577 11367 7611 11368
rect 7651 11367 7685 11368
rect 7725 11367 7759 11368
rect 7799 11367 7833 11368
rect 7873 11367 7907 11368
rect 7947 11367 7981 11368
rect 8021 11367 8055 11368
rect 8095 11367 8129 11368
rect 8169 11367 8203 11368
rect 8243 11367 8277 11368
rect 8317 11367 8351 11368
rect 8391 11367 8425 11401
rect 8465 11368 8495 11401
rect 8495 11368 8499 11401
rect 8539 11368 8564 11401
rect 8564 11368 8573 11401
rect 8613 11368 8633 11401
rect 8633 11368 8647 11401
rect 8687 11368 8702 11401
rect 8702 11368 8721 11401
rect 8761 11368 8771 11401
rect 8771 11368 8795 11401
rect 8835 11368 8840 11401
rect 8840 11368 8869 11401
rect 8909 11368 8943 11401
rect 8983 11368 9012 11401
rect 9012 11368 9017 11401
rect 9058 11368 9080 11401
rect 9080 11368 9092 11401
rect 9133 11368 9148 11401
rect 9148 11368 9167 11401
rect 9208 11368 9216 11401
rect 9216 11368 9242 11401
rect 9283 11368 9284 11401
rect 9284 11368 9317 11401
rect 9358 11368 9386 11401
rect 9386 11368 9392 11401
rect 9433 11368 9454 11401
rect 9454 11368 9467 11401
rect 9508 11368 9522 11401
rect 9522 11368 9542 11401
rect 17445 11384 17451 11401
rect 17451 11384 17479 11401
rect 17525 11384 17555 11401
rect 17555 11384 17559 11401
rect 17605 11384 17624 11401
rect 17624 11384 17639 11401
rect 17684 11384 17693 11401
rect 17693 11384 17718 11401
rect 17763 11384 17796 11401
rect 17796 11384 17797 11401
rect 17842 11384 17865 11401
rect 17865 11384 17876 11401
rect 17921 11384 17934 11401
rect 17934 11384 17955 11401
rect 18000 11384 18003 11401
rect 18003 11384 18034 11401
rect 18079 11384 18107 11401
rect 18107 11384 18113 11401
rect 18158 11384 18176 11401
rect 18176 11384 18192 11401
rect 18500 11384 18521 11399
rect 18521 11384 18534 11399
rect 18585 11384 18590 11399
rect 18590 11384 18619 11399
rect 18669 11384 18693 11399
rect 18693 11384 18703 11399
rect 18753 11384 18762 11399
rect 18762 11384 18787 11399
rect 18837 11384 18866 11399
rect 18866 11384 18871 11399
rect 18921 11384 18935 11399
rect 18935 11384 18955 11399
rect 8465 11367 8499 11368
rect 8539 11367 8573 11368
rect 8613 11367 8647 11368
rect 8687 11367 8721 11368
rect 8761 11367 8795 11368
rect 8835 11367 8869 11368
rect 8909 11367 8943 11368
rect 8983 11367 9017 11368
rect 9058 11367 9092 11368
rect 9133 11367 9167 11368
rect 9208 11367 9242 11368
rect 9283 11367 9317 11368
rect 9358 11367 9392 11368
rect 9433 11367 9467 11368
rect 9508 11367 9542 11368
rect 17445 11367 17479 11384
rect 17525 11367 17559 11384
rect 17605 11367 17639 11384
rect 17684 11367 17718 11384
rect 17763 11367 17797 11384
rect 17842 11367 17876 11384
rect 17921 11367 17955 11384
rect 18000 11367 18034 11384
rect 18079 11367 18113 11384
rect 18158 11367 18192 11384
rect 18500 11365 18534 11384
rect 18585 11365 18619 11384
rect 18669 11365 18703 11384
rect 18753 11365 18787 11384
rect 18837 11365 18871 11384
rect 18921 11365 18955 11384
rect 6779 11330 6813 11363
rect 6867 11330 6901 11363
rect 6955 11330 6989 11363
rect 7043 11330 7077 11363
rect 7131 11330 7165 11363
rect 6779 11329 6804 11330
rect 6804 11329 6813 11330
rect 6867 11329 6873 11330
rect 6873 11329 6901 11330
rect 6955 11329 6977 11330
rect 6977 11329 6989 11330
rect 7043 11329 7046 11330
rect 7046 11329 7077 11330
rect 7131 11329 7149 11330
rect 7149 11329 7165 11330
rect 7577 11296 7598 11313
rect 7598 11296 7611 11313
rect 7651 11296 7667 11313
rect 7667 11296 7685 11313
rect 7725 11296 7736 11313
rect 7736 11296 7759 11313
rect 7799 11296 7805 11313
rect 7805 11296 7833 11313
rect 7873 11296 7874 11313
rect 7874 11296 7907 11313
rect 7947 11296 7977 11313
rect 7977 11296 7981 11313
rect 8021 11296 8046 11313
rect 8046 11296 8055 11313
rect 8095 11296 8115 11313
rect 8115 11296 8129 11313
rect 8169 11296 8184 11313
rect 8184 11296 8203 11313
rect 8243 11296 8253 11313
rect 8253 11296 8277 11313
rect 8317 11296 8322 11313
rect 8322 11296 8351 11313
rect 6779 11258 6813 11291
rect 6867 11258 6901 11291
rect 6955 11258 6989 11291
rect 7043 11258 7077 11291
rect 7131 11258 7165 11291
rect 7577 11279 7611 11296
rect 7651 11279 7685 11296
rect 7725 11279 7759 11296
rect 7799 11279 7833 11296
rect 7873 11279 7907 11296
rect 7947 11279 7981 11296
rect 8021 11279 8055 11296
rect 8095 11279 8129 11296
rect 8169 11279 8203 11296
rect 8243 11279 8277 11296
rect 8317 11279 8351 11296
rect 8391 11279 8425 11313
rect 8465 11296 8495 11313
rect 8495 11296 8499 11313
rect 8539 11296 8564 11313
rect 8564 11296 8573 11313
rect 8613 11296 8633 11313
rect 8633 11296 8647 11313
rect 8687 11296 8702 11313
rect 8702 11296 8721 11313
rect 8761 11296 8771 11313
rect 8771 11296 8795 11313
rect 8835 11296 8840 11313
rect 8840 11296 8869 11313
rect 8909 11296 8943 11313
rect 8983 11296 9012 11313
rect 9012 11296 9017 11313
rect 9058 11296 9080 11313
rect 9080 11296 9092 11313
rect 9133 11296 9148 11313
rect 9148 11296 9167 11313
rect 9208 11296 9216 11313
rect 9216 11296 9242 11313
rect 9283 11296 9284 11313
rect 9284 11296 9317 11313
rect 9358 11296 9386 11313
rect 9386 11296 9392 11313
rect 9433 11296 9454 11313
rect 9454 11296 9467 11313
rect 9508 11296 9522 11313
rect 9522 11296 9542 11313
rect 10456 11304 10490 11338
rect 10529 11304 10563 11338
rect 10602 11304 10636 11338
rect 10675 11304 10709 11338
rect 10748 11304 10782 11338
rect 10821 11304 10855 11338
rect 10893 11304 10927 11338
rect 10965 11304 10999 11338
rect 11037 11304 11071 11338
rect 11109 11304 11143 11338
rect 11181 11304 11215 11338
rect 11253 11304 11287 11338
rect 11325 11304 11359 11338
rect 11397 11304 11431 11338
rect 11469 11304 11503 11338
rect 11541 11304 11575 11338
rect 11613 11304 11647 11338
rect 11685 11304 11719 11338
rect 11757 11304 11791 11338
rect 11829 11304 11863 11338
rect 11901 11304 11935 11338
rect 11973 11304 12007 11338
rect 12045 11304 12079 11338
rect 12117 11304 12151 11338
rect 12189 11304 12223 11338
rect 12261 11304 12295 11338
rect 12333 11304 12367 11338
rect 13411 11304 13445 11338
rect 13485 11304 13519 11338
rect 13559 11304 13593 11338
rect 13633 11304 13667 11338
rect 13707 11304 13741 11338
rect 13781 11304 13815 11338
rect 13855 11304 13889 11338
rect 13929 11304 13963 11338
rect 14003 11304 14037 11338
rect 14077 11304 14111 11338
rect 14151 11304 14185 11338
rect 14225 11304 14259 11338
rect 14299 11304 14333 11338
rect 14372 11304 14406 11338
rect 14445 11304 14479 11338
rect 14518 11304 14552 11338
rect 14591 11304 14625 11338
rect 14664 11304 14698 11338
rect 14737 11304 14771 11338
rect 14810 11304 14844 11338
rect 14883 11304 14917 11338
rect 14956 11304 14990 11338
rect 15029 11304 15063 11338
rect 15102 11304 15136 11338
rect 15175 11304 15209 11338
rect 15248 11304 15282 11338
rect 15321 11304 15355 11338
rect 15394 11304 15428 11338
rect 15467 11304 15501 11338
rect 15540 11304 15574 11338
rect 15613 11304 15647 11338
rect 17445 11316 17478 11329
rect 17478 11316 17479 11329
rect 17525 11316 17546 11329
rect 17546 11316 17559 11329
rect 17605 11316 17614 11329
rect 17614 11316 17639 11329
rect 17684 11316 17716 11329
rect 17716 11316 17718 11329
rect 17763 11316 17784 11329
rect 17784 11316 17797 11329
rect 17842 11316 17852 11329
rect 17852 11316 17876 11329
rect 17921 11316 17954 11329
rect 17954 11316 17955 11329
rect 18000 11316 18022 11329
rect 18022 11316 18034 11329
rect 18079 11316 18090 11329
rect 18090 11316 18113 11329
rect 18158 11316 18192 11329
rect 18500 11316 18532 11327
rect 18532 11316 18534 11327
rect 18585 11316 18600 11327
rect 18600 11316 18619 11327
rect 18669 11316 18702 11327
rect 18702 11316 18703 11327
rect 18753 11316 18770 11327
rect 18770 11316 18787 11327
rect 18837 11316 18838 11327
rect 18838 11316 18871 11327
rect 18921 11316 18940 11327
rect 18940 11316 18955 11327
rect 8465 11279 8499 11296
rect 8539 11279 8573 11296
rect 8613 11279 8647 11296
rect 8687 11279 8721 11296
rect 8761 11279 8795 11296
rect 8835 11279 8869 11296
rect 8909 11279 8943 11296
rect 8983 11279 9017 11296
rect 9058 11279 9092 11296
rect 9133 11279 9167 11296
rect 9208 11279 9242 11296
rect 9283 11279 9317 11296
rect 9358 11279 9392 11296
rect 9433 11279 9467 11296
rect 9508 11279 9542 11296
rect 6779 11257 6804 11258
rect 6804 11257 6813 11258
rect 6867 11257 6873 11258
rect 6873 11257 6901 11258
rect 6955 11257 6977 11258
rect 6977 11257 6989 11258
rect 7043 11257 7046 11258
rect 7046 11257 7077 11258
rect 7131 11257 7149 11258
rect 7149 11257 7165 11258
rect 7577 11224 7598 11225
rect 7598 11224 7611 11225
rect 7651 11224 7667 11225
rect 7667 11224 7685 11225
rect 7725 11224 7736 11225
rect 7736 11224 7759 11225
rect 7799 11224 7805 11225
rect 7805 11224 7833 11225
rect 7873 11224 7874 11225
rect 7874 11224 7907 11225
rect 7947 11224 7977 11225
rect 7977 11224 7981 11225
rect 8021 11224 8046 11225
rect 8046 11224 8055 11225
rect 8095 11224 8115 11225
rect 8115 11224 8129 11225
rect 8169 11224 8184 11225
rect 8184 11224 8203 11225
rect 8243 11224 8253 11225
rect 8253 11224 8277 11225
rect 8317 11224 8322 11225
rect 8322 11224 8351 11225
rect 6779 11186 6813 11219
rect 6867 11186 6901 11219
rect 6955 11186 6989 11219
rect 7043 11186 7077 11219
rect 7131 11186 7165 11219
rect 7577 11191 7611 11224
rect 7651 11191 7685 11224
rect 7725 11191 7759 11224
rect 7799 11191 7833 11224
rect 7873 11191 7907 11224
rect 7947 11191 7981 11224
rect 8021 11191 8055 11224
rect 8095 11191 8129 11224
rect 8169 11191 8203 11224
rect 8243 11191 8277 11224
rect 8317 11191 8351 11224
rect 8391 11191 8425 11225
rect 8465 11224 8495 11225
rect 8495 11224 8499 11225
rect 8539 11224 8564 11225
rect 8564 11224 8573 11225
rect 8613 11224 8633 11225
rect 8633 11224 8647 11225
rect 8687 11224 8702 11225
rect 8702 11224 8721 11225
rect 8761 11224 8771 11225
rect 8771 11224 8795 11225
rect 8835 11224 8840 11225
rect 8840 11224 8869 11225
rect 8909 11224 8943 11225
rect 8983 11224 9012 11225
rect 9012 11224 9017 11225
rect 9058 11224 9080 11225
rect 9080 11224 9092 11225
rect 9133 11224 9148 11225
rect 9148 11224 9167 11225
rect 9208 11224 9216 11225
rect 9216 11224 9242 11225
rect 9283 11224 9284 11225
rect 9284 11224 9317 11225
rect 9358 11224 9386 11225
rect 9386 11224 9392 11225
rect 9433 11224 9454 11225
rect 9454 11224 9467 11225
rect 9508 11224 9522 11225
rect 9522 11224 9542 11225
rect 17445 11295 17479 11316
rect 17525 11295 17559 11316
rect 17605 11295 17639 11316
rect 17684 11295 17718 11316
rect 17763 11295 17797 11316
rect 17842 11295 17876 11316
rect 17921 11295 17955 11316
rect 18000 11295 18034 11316
rect 18079 11295 18113 11316
rect 18158 11295 18192 11316
rect 18500 11293 18534 11316
rect 18585 11293 18619 11316
rect 18669 11293 18703 11316
rect 18753 11293 18787 11316
rect 18837 11293 18871 11316
rect 18921 11293 18955 11316
rect 17445 11244 17478 11257
rect 17478 11244 17479 11257
rect 17525 11244 17546 11257
rect 17546 11244 17559 11257
rect 17605 11244 17614 11257
rect 17614 11244 17639 11257
rect 17684 11244 17716 11257
rect 17716 11244 17718 11257
rect 17763 11244 17784 11257
rect 17784 11244 17797 11257
rect 17842 11244 17852 11257
rect 17852 11244 17876 11257
rect 17921 11244 17954 11257
rect 17954 11244 17955 11257
rect 18000 11244 18022 11257
rect 18022 11244 18034 11257
rect 18079 11244 18090 11257
rect 18090 11244 18113 11257
rect 18158 11244 18192 11257
rect 18500 11244 18532 11255
rect 18532 11244 18534 11255
rect 18585 11244 18600 11255
rect 18600 11244 18619 11255
rect 18669 11244 18702 11255
rect 18702 11244 18703 11255
rect 18753 11244 18770 11255
rect 18770 11244 18787 11255
rect 18837 11244 18838 11255
rect 18838 11244 18871 11255
rect 18921 11244 18940 11255
rect 18940 11244 18955 11255
rect 8465 11191 8499 11224
rect 8539 11191 8573 11224
rect 8613 11191 8647 11224
rect 8687 11191 8721 11224
rect 8761 11191 8795 11224
rect 8835 11191 8869 11224
rect 8909 11191 8943 11224
rect 8983 11191 9017 11224
rect 9058 11191 9092 11224
rect 9133 11191 9167 11224
rect 9208 11191 9242 11224
rect 9283 11191 9317 11224
rect 9358 11191 9392 11224
rect 9433 11191 9467 11224
rect 9508 11191 9542 11224
rect 6779 11185 6804 11186
rect 6804 11185 6813 11186
rect 6867 11185 6873 11186
rect 6873 11185 6901 11186
rect 6955 11185 6977 11186
rect 6977 11185 6989 11186
rect 7043 11185 7046 11186
rect 7046 11185 7077 11186
rect 7131 11185 7149 11186
rect 7149 11185 7165 11186
rect 17445 11223 17479 11244
rect 17525 11223 17559 11244
rect 17605 11223 17639 11244
rect 17684 11223 17718 11244
rect 17763 11223 17797 11244
rect 17842 11223 17876 11244
rect 17921 11223 17955 11244
rect 18000 11223 18034 11244
rect 18079 11223 18113 11244
rect 18158 11223 18192 11244
rect 18500 11221 18534 11244
rect 18585 11221 18619 11244
rect 18669 11221 18703 11244
rect 18753 11221 18787 11244
rect 18837 11221 18871 11244
rect 18921 11221 18955 11244
rect 17445 11172 17478 11185
rect 17478 11172 17479 11185
rect 17525 11172 17546 11185
rect 17546 11172 17559 11185
rect 17605 11172 17614 11185
rect 17614 11172 17639 11185
rect 17684 11172 17716 11185
rect 17716 11172 17718 11185
rect 17763 11172 17784 11185
rect 17784 11172 17797 11185
rect 17842 11172 17852 11185
rect 17852 11172 17876 11185
rect 17921 11172 17954 11185
rect 17954 11172 17955 11185
rect 18000 11172 18022 11185
rect 18022 11172 18034 11185
rect 18079 11172 18090 11185
rect 18090 11172 18113 11185
rect 18158 11172 18192 11185
rect 18500 11172 18532 11183
rect 18532 11172 18534 11183
rect 18585 11172 18600 11183
rect 18600 11172 18619 11183
rect 18669 11172 18702 11183
rect 18702 11172 18703 11183
rect 18753 11172 18770 11183
rect 18770 11172 18787 11183
rect 18837 11172 18838 11183
rect 18838 11172 18871 11183
rect 18921 11172 18940 11183
rect 18940 11172 18955 11183
rect 17445 11151 17479 11172
rect 17525 11151 17559 11172
rect 17605 11151 17639 11172
rect 17684 11151 17718 11172
rect 17763 11151 17797 11172
rect 17842 11151 17876 11172
rect 17921 11151 17955 11172
rect 18000 11151 18034 11172
rect 18079 11151 18113 11172
rect 18158 11151 18192 11172
rect 18500 11149 18534 11172
rect 18585 11149 18619 11172
rect 18669 11149 18703 11172
rect 18753 11149 18787 11172
rect 18837 11149 18871 11172
rect 18921 11149 18955 11172
rect 6779 11113 6813 11147
rect 6867 11113 6901 11147
rect 6955 11113 6989 11147
rect 7043 11113 7077 11147
rect 7131 11113 7165 11147
rect 6779 11072 6813 11075
rect 6779 11041 6785 11072
rect 6785 11041 6813 11072
rect 6867 11041 6901 11075
rect 6955 11072 6989 11075
rect 7043 11072 7077 11075
rect 7131 11072 7165 11075
rect 6955 11041 6979 11072
rect 6979 11041 6989 11072
rect 7043 11041 7055 11072
rect 7055 11041 7077 11072
rect 7131 11041 7165 11072
rect 6779 10970 6785 11002
rect 6785 10970 6813 11002
rect 6779 10968 6813 10970
rect 6867 10968 6901 11002
rect 6955 10970 6979 11002
rect 6979 10970 6989 11002
rect 7043 10970 7055 11002
rect 7055 10970 7077 11002
rect 7131 10970 7165 11002
rect 6955 10968 6989 10970
rect 7043 10968 7077 10970
rect 7131 10968 7165 10970
rect 6779 10902 6785 10929
rect 6785 10902 6813 10929
rect 6779 10895 6813 10902
rect 6867 10895 6901 10929
rect 6955 10902 6979 10929
rect 6979 10902 6989 10929
rect 7043 10902 7055 10929
rect 7055 10902 7077 10929
rect 7131 10902 7165 10929
rect 6955 10895 6989 10902
rect 7043 10895 7077 10902
rect 7131 10895 7165 10902
rect 6779 10834 6785 10856
rect 6785 10834 6813 10856
rect 6779 10822 6813 10834
rect 6867 10822 6901 10856
rect 6955 10834 6979 10856
rect 6979 10834 6989 10856
rect 7043 10834 7055 10856
rect 7055 10834 7077 10856
rect 7131 10834 7165 10856
rect 6955 10822 6989 10834
rect 7043 10822 7077 10834
rect 7131 10822 7165 10834
rect 6779 10766 6785 10783
rect 6785 10766 6813 10783
rect 6779 10749 6813 10766
rect 6867 10749 6901 10783
rect 6955 10766 6979 10783
rect 6979 10766 6989 10783
rect 7043 10766 7055 10783
rect 7055 10766 7077 10783
rect 7131 10766 7165 10783
rect 6955 10749 6989 10766
rect 7043 10749 7077 10766
rect 7131 10749 7165 10766
rect 7155 10664 7189 10696
rect 7155 10662 7165 10664
rect 7165 10662 7189 10664
rect 7155 10596 7189 10620
rect 7155 10586 7165 10596
rect 7165 10586 7189 10596
rect 7155 10528 7189 10544
rect 7155 10510 7165 10528
rect 7165 10510 7189 10528
rect 7155 10460 7189 10468
rect 7155 10434 7165 10460
rect 7165 10434 7189 10460
rect 7155 10358 7165 10392
rect 7165 10358 7189 10392
rect 7155 10290 7165 10316
rect 7165 10290 7189 10316
rect 7155 10282 7189 10290
rect 19581 11283 19615 11317
rect 19581 11208 19615 11242
rect 19581 11133 19615 11167
rect 19581 11057 19615 11091
rect 10072 10653 10106 10687
rect 10178 10653 10212 10687
rect 10072 10581 10106 10615
rect 10178 10581 10212 10615
rect 10072 10509 10106 10543
rect 10178 10509 10212 10543
rect 10072 10437 10106 10471
rect 10178 10437 10212 10471
rect 10072 10365 10106 10399
rect 10178 10365 10212 10399
rect 10072 10293 10106 10327
rect 10178 10293 10212 10327
rect 7155 10222 7165 10240
rect 7165 10222 7189 10240
rect 7266 10227 7300 10261
rect 7155 10206 7189 10222
rect 7155 10154 7165 10164
rect 7165 10154 7189 10164
rect 7266 10155 7300 10189
rect 7155 10130 7189 10154
rect 7155 10086 7165 10088
rect 7165 10086 7189 10088
rect 7155 10054 7189 10086
rect 7266 10083 7300 10117
rect 7155 9984 7189 10012
rect 7266 10011 7300 10045
rect 7155 9978 7165 9984
rect 7165 9978 7189 9984
rect 7266 9939 7300 9973
rect 7155 9916 7189 9935
rect 7155 9901 7165 9916
rect 7165 9901 7189 9916
rect 7266 9867 7300 9901
rect 7155 9848 7189 9858
rect 7155 9824 7165 9848
rect 7165 9824 7189 9848
rect 7266 9795 7300 9829
rect 7155 9780 7189 9781
rect 7155 9747 7165 9780
rect 7165 9747 7189 9780
rect 7266 9723 7300 9757
rect 7155 9678 7165 9704
rect 7165 9678 7189 9704
rect 19581 11002 19582 11015
rect 19582 11002 19615 11015
rect 19581 10981 19615 11002
rect 19581 10933 19615 10939
rect 19581 10905 19582 10933
rect 19582 10905 19615 10933
rect 19581 10830 19615 10863
rect 19581 10829 19582 10830
rect 19582 10829 19615 10830
rect 19581 10753 19615 10787
rect 19581 10693 19582 10711
rect 19582 10693 19615 10711
rect 19581 10677 19615 10693
rect 19581 10623 19615 10635
rect 19581 10601 19582 10623
rect 19582 10601 19615 10623
rect 19581 10525 19615 10559
rect 19581 10449 19615 10483
rect 19581 10381 19582 10407
rect 19582 10381 19615 10407
rect 19581 10373 19615 10381
rect 19581 10311 19615 10331
rect 19581 10297 19582 10311
rect 19582 10297 19615 10311
rect 10072 10221 10083 10255
rect 10083 10221 10106 10255
rect 10178 10221 10185 10255
rect 10185 10221 10212 10255
rect 10072 10152 10083 10183
rect 10083 10152 10106 10183
rect 10178 10152 10185 10183
rect 10185 10152 10212 10183
rect 10072 10149 10106 10152
rect 10178 10149 10212 10152
rect 10072 10083 10083 10111
rect 10083 10083 10106 10111
rect 10178 10083 10185 10111
rect 10185 10083 10212 10111
rect 10072 10077 10106 10083
rect 10178 10077 10212 10083
rect 10072 10014 10083 10039
rect 10083 10014 10106 10039
rect 10178 10014 10185 10039
rect 10185 10014 10212 10039
rect 10072 10005 10106 10014
rect 10178 10005 10212 10014
rect 10072 9945 10083 9967
rect 10083 9945 10106 9967
rect 10178 9945 10185 9967
rect 10185 9945 10212 9967
rect 10072 9933 10106 9945
rect 10178 9933 10212 9945
rect 10072 9876 10083 9895
rect 10083 9876 10106 9895
rect 10178 9876 10185 9895
rect 10185 9876 10212 9895
rect 10072 9861 10106 9876
rect 10178 9861 10212 9876
rect 10072 9807 10083 9823
rect 10083 9807 10106 9823
rect 10178 9807 10185 9823
rect 10185 9807 10212 9823
rect 10072 9789 10106 9807
rect 10178 9789 10212 9807
rect 10072 9738 10083 9751
rect 10083 9738 10106 9751
rect 10178 9738 10185 9751
rect 10185 9738 10212 9751
rect 10072 9717 10106 9738
rect 10178 9717 10212 9738
rect 7155 9670 7189 9678
rect 7266 9651 7300 9685
rect 7360 9665 7394 9699
rect 7435 9665 7469 9699
rect 7510 9665 7544 9699
rect 7585 9665 7619 9699
rect 7660 9665 7694 9699
rect 7735 9665 7769 9699
rect 7810 9665 7844 9699
rect 7885 9665 7919 9699
rect 7960 9665 7994 9699
rect 8035 9665 8069 9699
rect 8110 9665 8144 9699
rect 8185 9665 8219 9699
rect 8260 9665 8294 9699
rect 8335 9665 8369 9699
rect 8410 9665 8444 9699
rect 8485 9665 8519 9699
rect 8559 9665 8593 9699
rect 8633 9665 8667 9699
rect 8707 9665 8741 9699
rect 8781 9665 8815 9699
rect 8855 9665 8889 9699
rect 8929 9665 8963 9699
rect 9003 9665 9037 9699
rect 9077 9665 9111 9699
rect 9151 9665 9185 9699
rect 10072 9669 10083 9678
rect 10083 9669 10106 9678
rect 10178 9669 10185 9678
rect 10185 9669 10212 9678
rect 7155 9610 7165 9627
rect 7165 9610 7189 9627
rect 7155 9593 7189 9610
rect 7266 9579 7300 9613
rect 10072 9644 10106 9669
rect 10178 9644 10212 9669
rect 10072 9600 10083 9605
rect 10083 9600 10106 9605
rect 10178 9600 10185 9605
rect 10185 9600 10212 9605
rect 8333 9588 8367 9592
rect 8406 9588 8440 9592
rect 8479 9588 8513 9592
rect 8553 9588 8587 9592
rect 8627 9588 8661 9592
rect 7883 9554 7884 9582
rect 7884 9554 7917 9582
rect 8011 9554 8022 9582
rect 8022 9554 8045 9582
rect 8333 9558 8365 9588
rect 8365 9558 8367 9588
rect 8406 9558 8433 9588
rect 8433 9558 8440 9588
rect 8479 9558 8501 9588
rect 8501 9558 8513 9588
rect 8553 9558 8569 9588
rect 8569 9558 8587 9588
rect 8627 9558 8637 9588
rect 8637 9558 8661 9588
rect 9057 9554 9079 9582
rect 9079 9554 9091 9582
rect 9185 9554 9215 9582
rect 9215 9554 9219 9582
rect 10072 9571 10106 9600
rect 10178 9571 10212 9600
rect 7883 9548 7917 9554
rect 8011 9548 8045 9554
rect 9057 9548 9091 9554
rect 9185 9548 9219 9554
rect 7266 9507 7300 9541
rect 10072 9531 10083 9532
rect 10083 9531 10106 9532
rect 19581 10221 19615 10255
rect 19581 10173 19582 10179
rect 19582 10173 19615 10179
rect 16708 10148 16733 10154
rect 16733 10148 16742 10154
rect 16781 10148 16801 10154
rect 16801 10148 16815 10154
rect 16708 10120 16742 10148
rect 16781 10120 16815 10148
rect 16854 10120 16888 10154
rect 16708 10075 16733 10082
rect 16733 10075 16742 10082
rect 16781 10075 16801 10082
rect 16801 10075 16815 10082
rect 16708 10048 16742 10075
rect 16781 10048 16815 10075
rect 16854 10048 16888 10082
rect 19581 10145 19615 10173
rect 19581 10069 19582 10103
rect 19582 10069 19615 10103
rect 19581 9999 19615 10027
rect 19581 9993 19582 9999
rect 19582 9993 19615 9999
rect 19581 9917 19615 9951
rect 26272 10302 26306 10332
rect 26348 10302 26382 10332
rect 26424 10302 26458 10332
rect 26500 10302 26534 10332
rect 26576 10302 26610 10332
rect 26652 10302 26686 10332
rect 26727 10302 26761 10332
rect 26802 10302 26836 10332
rect 26877 10302 26911 10332
rect 26272 10298 26277 10302
rect 26277 10298 26306 10302
rect 26348 10298 26382 10302
rect 26424 10298 26453 10302
rect 26453 10298 26458 10302
rect 26500 10298 26524 10302
rect 26524 10298 26534 10302
rect 26576 10298 26595 10302
rect 26595 10298 26610 10302
rect 26652 10298 26666 10302
rect 26666 10298 26686 10302
rect 26727 10298 26737 10302
rect 26737 10298 26761 10302
rect 26802 10298 26808 10302
rect 26808 10298 26836 10302
rect 26877 10298 26879 10302
rect 26879 10298 26911 10302
rect 26952 10298 26986 10332
rect 27027 10302 27061 10332
rect 27102 10302 27136 10332
rect 27177 10302 27211 10332
rect 27252 10302 27286 10332
rect 27327 10302 27361 10332
rect 27402 10302 27436 10332
rect 27501 10307 27535 10341
rect 27573 10312 27581 10341
rect 27581 10312 27607 10341
rect 27645 10312 27649 10341
rect 27649 10312 27679 10341
rect 27573 10307 27607 10312
rect 27645 10307 27679 10312
rect 27717 10307 27751 10341
rect 27789 10312 27819 10341
rect 27819 10312 27823 10341
rect 27789 10307 27823 10312
rect 27861 10307 27895 10341
rect 27027 10298 27056 10302
rect 27056 10298 27061 10302
rect 27102 10298 27126 10302
rect 27126 10298 27136 10302
rect 27177 10298 27196 10302
rect 27196 10298 27211 10302
rect 27252 10298 27266 10302
rect 27266 10298 27286 10302
rect 27327 10298 27336 10302
rect 27336 10298 27361 10302
rect 27402 10298 27406 10302
rect 27406 10298 27436 10302
rect 26272 10234 26306 10260
rect 26348 10234 26382 10260
rect 26424 10234 26458 10260
rect 26500 10234 26534 10260
rect 26576 10234 26610 10260
rect 26652 10234 26686 10260
rect 26727 10234 26761 10260
rect 26802 10234 26836 10260
rect 26877 10234 26911 10260
rect 26272 10226 26277 10234
rect 26277 10226 26306 10234
rect 26348 10226 26382 10234
rect 26424 10226 26453 10234
rect 26453 10226 26458 10234
rect 26500 10226 26524 10234
rect 26524 10226 26534 10234
rect 26576 10226 26595 10234
rect 26595 10226 26610 10234
rect 26652 10226 26666 10234
rect 26666 10226 26686 10234
rect 26727 10226 26737 10234
rect 26737 10226 26761 10234
rect 26802 10226 26808 10234
rect 26808 10226 26836 10234
rect 26877 10226 26879 10234
rect 26879 10226 26911 10234
rect 26952 10226 26986 10260
rect 27027 10234 27061 10260
rect 27102 10234 27136 10260
rect 27177 10234 27211 10260
rect 27252 10234 27286 10260
rect 27327 10234 27361 10260
rect 27402 10234 27436 10260
rect 27501 10234 27535 10268
rect 27573 10243 27581 10268
rect 27581 10243 27607 10268
rect 27645 10243 27649 10268
rect 27649 10243 27679 10268
rect 27573 10234 27607 10243
rect 27645 10234 27679 10243
rect 27717 10234 27751 10268
rect 27789 10243 27819 10268
rect 27819 10243 27823 10268
rect 27789 10234 27823 10243
rect 27861 10234 27895 10268
rect 27027 10226 27056 10234
rect 27056 10226 27061 10234
rect 27102 10226 27126 10234
rect 27126 10226 27136 10234
rect 27177 10226 27196 10234
rect 27196 10226 27211 10234
rect 27252 10226 27266 10234
rect 27266 10226 27286 10234
rect 27327 10226 27336 10234
rect 27336 10226 27361 10234
rect 27402 10226 27406 10234
rect 27406 10226 27436 10234
rect 26272 10166 26306 10188
rect 26348 10166 26382 10188
rect 26424 10166 26458 10188
rect 26500 10166 26534 10188
rect 26576 10166 26610 10188
rect 26652 10166 26686 10188
rect 26727 10166 26761 10188
rect 26802 10166 26836 10188
rect 26877 10166 26911 10188
rect 26272 10154 26277 10166
rect 26277 10154 26306 10166
rect 26348 10154 26382 10166
rect 26424 10154 26453 10166
rect 26453 10154 26458 10166
rect 26500 10154 26524 10166
rect 26524 10154 26534 10166
rect 26576 10154 26595 10166
rect 26595 10154 26610 10166
rect 26652 10154 26666 10166
rect 26666 10154 26686 10166
rect 26727 10154 26737 10166
rect 26737 10154 26761 10166
rect 26802 10154 26808 10166
rect 26808 10154 26836 10166
rect 26877 10154 26879 10166
rect 26879 10154 26911 10166
rect 26952 10154 26986 10188
rect 27027 10166 27061 10188
rect 27102 10166 27136 10188
rect 27177 10166 27211 10188
rect 27252 10166 27286 10188
rect 27327 10166 27361 10188
rect 27402 10166 27436 10188
rect 27027 10154 27056 10166
rect 27056 10154 27061 10166
rect 27102 10154 27126 10166
rect 27126 10154 27136 10166
rect 27177 10154 27196 10166
rect 27196 10154 27211 10166
rect 27252 10154 27266 10166
rect 27266 10154 27286 10166
rect 27327 10154 27336 10166
rect 27336 10154 27361 10166
rect 27402 10154 27406 10166
rect 27406 10154 27436 10166
rect 27501 10161 27535 10195
rect 27573 10174 27581 10195
rect 27581 10174 27607 10195
rect 27645 10174 27649 10195
rect 27649 10174 27679 10195
rect 27573 10161 27607 10174
rect 27645 10161 27679 10174
rect 27717 10161 27751 10195
rect 27789 10174 27819 10195
rect 27819 10174 27823 10195
rect 27789 10161 27823 10174
rect 27861 10161 27895 10195
rect 26272 10098 26306 10116
rect 26348 10098 26382 10116
rect 26424 10098 26458 10116
rect 26500 10098 26534 10116
rect 26576 10098 26610 10116
rect 26652 10098 26686 10116
rect 26727 10098 26761 10116
rect 26802 10098 26836 10116
rect 26877 10098 26911 10116
rect 26272 10082 26277 10098
rect 26277 10082 26306 10098
rect 26348 10082 26382 10098
rect 26424 10082 26453 10098
rect 26453 10082 26458 10098
rect 26500 10082 26524 10098
rect 26524 10082 26534 10098
rect 26576 10082 26595 10098
rect 26595 10082 26610 10098
rect 26652 10082 26666 10098
rect 26666 10082 26686 10098
rect 26727 10082 26737 10098
rect 26737 10082 26761 10098
rect 26802 10082 26808 10098
rect 26808 10082 26836 10098
rect 26877 10082 26879 10098
rect 26879 10082 26911 10098
rect 26952 10082 26986 10116
rect 27027 10098 27061 10116
rect 27102 10098 27136 10116
rect 27177 10098 27211 10116
rect 27252 10098 27286 10116
rect 27327 10098 27361 10116
rect 27402 10098 27436 10116
rect 27027 10082 27056 10098
rect 27056 10082 27061 10098
rect 27102 10082 27126 10098
rect 27126 10082 27136 10098
rect 27177 10082 27196 10098
rect 27196 10082 27211 10098
rect 27252 10082 27266 10098
rect 27266 10082 27286 10098
rect 27327 10082 27336 10098
rect 27336 10082 27361 10098
rect 27402 10082 27406 10098
rect 27406 10082 27436 10098
rect 27501 10088 27535 10122
rect 27573 10105 27581 10122
rect 27581 10105 27607 10122
rect 27645 10105 27649 10122
rect 27649 10105 27679 10122
rect 27573 10088 27607 10105
rect 27645 10088 27679 10105
rect 27717 10088 27751 10122
rect 27789 10105 27819 10122
rect 27819 10105 27823 10122
rect 27789 10088 27823 10105
rect 27861 10088 27895 10122
rect 26272 10030 26306 10044
rect 26348 10030 26382 10044
rect 26424 10030 26458 10044
rect 26500 10030 26534 10044
rect 26576 10030 26610 10044
rect 26652 10030 26686 10044
rect 26727 10030 26761 10044
rect 26802 10030 26836 10044
rect 26877 10030 26911 10044
rect 26272 10010 26277 10030
rect 26277 10010 26306 10030
rect 26348 10010 26382 10030
rect 26424 10010 26453 10030
rect 26453 10010 26458 10030
rect 26500 10010 26524 10030
rect 26524 10010 26534 10030
rect 26576 10010 26595 10030
rect 26595 10010 26610 10030
rect 26652 10010 26666 10030
rect 26666 10010 26686 10030
rect 26727 10010 26737 10030
rect 26737 10010 26761 10030
rect 26802 10010 26808 10030
rect 26808 10010 26836 10030
rect 26877 10010 26879 10030
rect 26879 10010 26911 10030
rect 26952 10010 26986 10044
rect 27027 10030 27061 10044
rect 27102 10030 27136 10044
rect 27177 10030 27211 10044
rect 27252 10030 27286 10044
rect 27327 10030 27361 10044
rect 27402 10030 27436 10044
rect 27027 10010 27056 10030
rect 27056 10010 27061 10030
rect 27102 10010 27126 10030
rect 27126 10010 27136 10030
rect 27177 10010 27196 10030
rect 27196 10010 27211 10030
rect 27252 10010 27266 10030
rect 27266 10010 27286 10030
rect 27327 10010 27336 10030
rect 27336 10010 27361 10030
rect 27402 10010 27406 10030
rect 27406 10010 27436 10030
rect 27501 10015 27535 10049
rect 27573 10036 27581 10049
rect 27581 10036 27607 10049
rect 27645 10036 27649 10049
rect 27649 10036 27679 10049
rect 27573 10015 27607 10036
rect 27645 10015 27679 10036
rect 27717 10015 27751 10049
rect 27789 10036 27819 10049
rect 27819 10036 27823 10049
rect 27789 10015 27823 10036
rect 27861 10015 27895 10049
rect 26272 9962 26306 9972
rect 26348 9962 26382 9972
rect 26424 9962 26458 9972
rect 26500 9962 26534 9972
rect 26576 9962 26610 9972
rect 26652 9962 26686 9972
rect 26727 9962 26761 9972
rect 26802 9962 26836 9972
rect 26877 9962 26911 9972
rect 26272 9938 26277 9962
rect 26277 9938 26306 9962
rect 26348 9938 26382 9962
rect 26424 9938 26453 9962
rect 26453 9938 26458 9962
rect 26500 9938 26524 9962
rect 26524 9938 26534 9962
rect 26576 9938 26595 9962
rect 26595 9938 26610 9962
rect 26652 9938 26666 9962
rect 26666 9938 26686 9962
rect 26727 9938 26737 9962
rect 26737 9938 26761 9962
rect 26802 9938 26808 9962
rect 26808 9938 26836 9962
rect 26877 9938 26879 9962
rect 26879 9938 26911 9962
rect 26952 9938 26986 9972
rect 27027 9962 27061 9972
rect 27102 9962 27136 9972
rect 27177 9962 27211 9972
rect 27252 9962 27286 9972
rect 27327 9962 27361 9972
rect 27402 9962 27436 9972
rect 27027 9938 27056 9962
rect 27056 9938 27061 9962
rect 27102 9938 27126 9962
rect 27126 9938 27136 9962
rect 27177 9938 27196 9962
rect 27196 9938 27211 9962
rect 27252 9938 27266 9962
rect 27266 9938 27286 9962
rect 27327 9938 27336 9962
rect 27336 9938 27361 9962
rect 27402 9938 27406 9962
rect 27406 9938 27436 9962
rect 27501 9942 27535 9976
rect 27573 9967 27581 9976
rect 27581 9967 27607 9976
rect 27645 9967 27649 9976
rect 27649 9967 27679 9976
rect 27573 9942 27607 9967
rect 27645 9942 27679 9967
rect 27717 9942 27751 9976
rect 27789 9967 27819 9976
rect 27819 9967 27823 9976
rect 27789 9942 27823 9967
rect 27861 9942 27895 9976
rect 26272 9894 26306 9900
rect 26348 9894 26382 9900
rect 26424 9894 26458 9900
rect 26500 9894 26534 9900
rect 26576 9894 26610 9900
rect 26652 9894 26686 9900
rect 26727 9894 26761 9900
rect 26802 9894 26836 9900
rect 26877 9894 26911 9900
rect 26272 9866 26277 9894
rect 26277 9866 26306 9894
rect 26348 9866 26382 9894
rect 26424 9866 26453 9894
rect 26453 9866 26458 9894
rect 26500 9866 26524 9894
rect 26524 9866 26534 9894
rect 26576 9866 26595 9894
rect 26595 9866 26610 9894
rect 26652 9866 26666 9894
rect 26666 9866 26686 9894
rect 26727 9866 26737 9894
rect 26737 9866 26761 9894
rect 26802 9866 26808 9894
rect 26808 9866 26836 9894
rect 26877 9866 26879 9894
rect 26879 9866 26911 9894
rect 26952 9866 26986 9900
rect 27027 9894 27061 9900
rect 27102 9894 27136 9900
rect 27177 9894 27211 9900
rect 27252 9894 27286 9900
rect 27327 9894 27361 9900
rect 27402 9894 27436 9900
rect 27027 9866 27056 9894
rect 27056 9866 27061 9894
rect 27102 9866 27126 9894
rect 27126 9866 27136 9894
rect 27177 9866 27196 9894
rect 27196 9866 27211 9894
rect 27252 9866 27266 9894
rect 27266 9866 27286 9894
rect 27327 9866 27336 9894
rect 27336 9866 27361 9894
rect 27402 9866 27406 9894
rect 27406 9866 27436 9894
rect 27501 9868 27535 9902
rect 27573 9898 27581 9902
rect 27581 9898 27607 9902
rect 27645 9898 27649 9902
rect 27649 9898 27679 9902
rect 27573 9868 27607 9898
rect 27645 9868 27679 9898
rect 27717 9868 27751 9902
rect 27789 9898 27819 9902
rect 27819 9898 27823 9902
rect 27789 9868 27823 9898
rect 27861 9868 27895 9902
rect 27501 9794 27535 9828
rect 27573 9794 27607 9828
rect 27645 9794 27679 9828
rect 27717 9794 27751 9828
rect 27789 9794 27823 9828
rect 27861 9794 27895 9828
rect 27501 9720 27535 9754
rect 27573 9724 27607 9754
rect 27645 9724 27679 9754
rect 27573 9720 27581 9724
rect 27581 9720 27607 9724
rect 27645 9720 27649 9724
rect 27649 9720 27679 9724
rect 27717 9720 27751 9754
rect 27789 9724 27823 9754
rect 27789 9720 27819 9724
rect 27819 9720 27823 9724
rect 27861 9720 27895 9754
rect 27501 9646 27535 9680
rect 27573 9654 27607 9680
rect 27645 9654 27679 9680
rect 27573 9646 27581 9654
rect 27581 9646 27607 9654
rect 27645 9646 27649 9654
rect 27649 9646 27679 9654
rect 27717 9646 27751 9680
rect 27789 9654 27823 9680
rect 27789 9646 27819 9654
rect 27819 9646 27823 9654
rect 27861 9646 27895 9680
rect 27501 9572 27535 9606
rect 27573 9584 27607 9606
rect 27645 9584 27679 9606
rect 27573 9572 27581 9584
rect 27581 9572 27607 9584
rect 27645 9572 27649 9584
rect 27649 9572 27679 9584
rect 27717 9572 27751 9606
rect 27789 9584 27823 9606
rect 27789 9572 27819 9584
rect 27819 9572 27823 9584
rect 27861 9572 27895 9606
rect 10178 9531 10185 9532
rect 10185 9531 10212 9532
rect 7883 9496 7917 9510
rect 8011 9496 8045 9510
rect 8333 9496 8367 9520
rect 8406 9496 8440 9520
rect 8479 9496 8513 9520
rect 8553 9496 8587 9520
rect 8627 9496 8661 9520
rect 9057 9496 9091 9508
rect 9185 9496 9219 9508
rect 10072 9498 10106 9531
rect 10178 9498 10212 9531
rect 7266 9435 7300 9469
rect 7883 9476 7884 9496
rect 7884 9476 7917 9496
rect 8011 9476 8022 9496
rect 8022 9476 8045 9496
rect 8333 9486 8365 9496
rect 8365 9486 8367 9496
rect 8406 9486 8433 9496
rect 8433 9486 8440 9496
rect 8479 9486 8501 9496
rect 8501 9486 8513 9496
rect 8553 9486 8569 9496
rect 8569 9486 8587 9496
rect 8627 9486 8637 9496
rect 8637 9486 8661 9496
rect 9057 9474 9079 9496
rect 9079 9474 9091 9496
rect 9185 9474 9215 9496
rect 9215 9474 9219 9496
rect 7883 9404 7917 9438
rect 8011 9404 8045 9438
rect 9057 9404 9091 9434
rect 9185 9404 9219 9434
rect 10072 9427 10106 9459
rect 10178 9427 10212 9459
rect 10072 9425 10083 9427
rect 10083 9425 10106 9427
rect 7266 9363 7300 9397
rect 9057 9400 9079 9404
rect 9079 9400 9091 9404
rect 9185 9400 9215 9404
rect 9215 9400 9219 9404
rect 10178 9425 10185 9427
rect 10185 9425 10212 9427
rect 27501 9498 27535 9532
rect 27573 9514 27607 9532
rect 27645 9514 27679 9532
rect 27573 9498 27581 9514
rect 27581 9498 27607 9514
rect 27645 9498 27649 9514
rect 27649 9498 27679 9514
rect 27717 9498 27751 9532
rect 27789 9514 27823 9532
rect 27789 9498 27819 9514
rect 27819 9498 27823 9514
rect 27861 9498 27895 9532
rect 7266 9290 7300 9324
rect 7028 9236 7062 9250
rect 7028 9216 7055 9236
rect 7055 9216 7062 9236
rect 7266 9217 7300 9251
rect 7028 9168 7062 9177
rect 7028 9143 7055 9168
rect 7055 9143 7062 9168
rect 7266 9144 7300 9178
rect 7028 9100 7062 9103
rect 7028 9069 7055 9100
rect 7055 9069 7062 9100
rect 7266 9071 7300 9105
rect 7028 8998 7055 9029
rect 7055 8998 7062 9029
rect 7266 8998 7300 9032
rect 7028 8995 7062 8998
rect 7028 8930 7055 8955
rect 7055 8930 7062 8955
rect 7028 8921 7062 8930
rect 7266 8925 7300 8959
rect 6931 8862 6937 8876
rect 6937 8862 6965 8876
rect 7051 8862 7055 8876
rect 7055 8862 7085 8876
rect 6931 8842 6965 8862
rect 7051 8842 7085 8862
rect 7266 8852 7300 8886
rect 6931 8760 6965 8792
rect 7051 8760 7085 8792
rect 7266 8779 7300 8813
rect 6931 8758 6937 8760
rect 6937 8758 6965 8760
rect 7051 8758 7055 8760
rect 7055 8758 7085 8760
rect 6931 8692 6965 8708
rect 7051 8692 7085 8708
rect 7266 8706 7300 8740
rect 6931 8674 6937 8692
rect 6937 8674 6965 8692
rect 7051 8674 7055 8692
rect 7055 8674 7085 8692
rect 7266 8633 7300 8667
rect 6931 8590 6937 8624
rect 6937 8590 6965 8624
rect 7051 8590 7055 8624
rect 7055 8590 7085 8624
rect 6749 8555 6783 8584
rect 6851 8555 6885 8584
rect 7266 8560 7300 8594
rect 6749 8550 6751 8555
rect 6751 8550 6783 8555
rect 6851 8550 6861 8555
rect 6861 8550 6885 8555
rect 6931 8521 6937 8540
rect 6937 8521 6965 8540
rect 7051 8521 7055 8540
rect 7055 8521 7085 8540
rect 6931 8506 6965 8521
rect 7051 8506 7085 8521
rect 6749 8471 6783 8505
rect 6851 8471 6885 8505
rect 6749 8392 6783 8426
rect 6851 8392 6885 8426
rect 6749 8313 6783 8347
rect 6851 8313 6885 8347
rect 7266 8487 7300 8521
rect 27501 9424 27535 9458
rect 27573 9444 27607 9458
rect 27645 9444 27679 9458
rect 27573 9424 27581 9444
rect 27581 9424 27607 9444
rect 27645 9424 27649 9444
rect 27649 9424 27679 9444
rect 27717 9424 27751 9458
rect 27789 9444 27823 9458
rect 27789 9424 27819 9444
rect 27819 9424 27823 9444
rect 27861 9424 27895 9458
rect 27501 9350 27535 9384
rect 27573 9374 27607 9384
rect 27645 9374 27679 9384
rect 27573 9350 27581 9374
rect 27581 9350 27607 9374
rect 27645 9350 27649 9374
rect 27649 9350 27679 9374
rect 27717 9350 27751 9384
rect 27789 9374 27823 9384
rect 27789 9350 27819 9374
rect 27819 9350 27823 9374
rect 27861 9350 27895 9384
rect 27501 9276 27535 9310
rect 27573 9304 27607 9310
rect 27645 9304 27679 9310
rect 27573 9276 27581 9304
rect 27581 9276 27607 9304
rect 27645 9276 27649 9304
rect 27649 9276 27679 9304
rect 27717 9276 27751 9310
rect 27789 9304 27823 9310
rect 27789 9276 27819 9304
rect 27819 9276 27823 9304
rect 27861 9276 27895 9310
rect 27501 9202 27535 9236
rect 27573 9234 27607 9236
rect 27645 9234 27679 9236
rect 27573 9202 27581 9234
rect 27581 9202 27607 9234
rect 27645 9202 27649 9234
rect 27649 9202 27679 9234
rect 27717 9202 27751 9236
rect 27789 9234 27823 9236
rect 27789 9202 27819 9234
rect 27819 9202 27823 9234
rect 27861 9202 27895 9236
rect 27501 9128 27535 9162
rect 27573 9130 27581 9162
rect 27581 9130 27607 9162
rect 27645 9130 27649 9162
rect 27649 9130 27679 9162
rect 27573 9128 27607 9130
rect 27645 9128 27679 9130
rect 27717 9128 27751 9162
rect 27789 9130 27819 9162
rect 27819 9130 27823 9162
rect 27789 9128 27823 9130
rect 27861 9128 27895 9162
rect 27501 9054 27535 9088
rect 27573 9060 27581 9088
rect 27581 9060 27607 9088
rect 27645 9060 27649 9088
rect 27649 9060 27679 9088
rect 27573 9054 27607 9060
rect 27645 9054 27679 9060
rect 27717 9054 27751 9088
rect 27789 9060 27819 9088
rect 27819 9060 27823 9088
rect 27789 9054 27823 9060
rect 27861 9054 27895 9088
rect 27501 8980 27535 9014
rect 27573 8990 27581 9014
rect 27581 8990 27607 9014
rect 27645 8990 27649 9014
rect 27649 8990 27679 9014
rect 27573 8980 27607 8990
rect 27645 8980 27679 8990
rect 27717 8980 27751 9014
rect 27789 8990 27819 9014
rect 27819 8990 27823 9014
rect 27789 8980 27823 8990
rect 27861 8980 27895 9014
rect 27501 8906 27535 8940
rect 27573 8920 27581 8940
rect 27581 8920 27607 8940
rect 27645 8920 27649 8940
rect 27649 8920 27679 8940
rect 27573 8906 27607 8920
rect 27645 8906 27679 8920
rect 27717 8906 27751 8940
rect 27789 8920 27819 8940
rect 27819 8920 27823 8940
rect 27789 8906 27823 8920
rect 27861 8906 27895 8940
rect 27501 8832 27535 8866
rect 27573 8850 27581 8866
rect 27581 8850 27607 8866
rect 27645 8850 27649 8866
rect 27649 8850 27679 8866
rect 27573 8832 27607 8850
rect 27645 8832 27679 8850
rect 27717 8832 27751 8866
rect 27789 8850 27819 8866
rect 27819 8850 27823 8866
rect 27789 8832 27823 8850
rect 27861 8832 27895 8866
rect 27501 8758 27535 8792
rect 27573 8780 27581 8792
rect 27581 8780 27607 8792
rect 27645 8780 27649 8792
rect 27649 8780 27679 8792
rect 27573 8758 27607 8780
rect 27645 8758 27679 8780
rect 27717 8758 27751 8792
rect 27789 8780 27819 8792
rect 27819 8780 27823 8792
rect 27789 8758 27823 8780
rect 27861 8758 27895 8792
rect 27501 8684 27535 8718
rect 27573 8710 27581 8718
rect 27581 8710 27607 8718
rect 27645 8710 27649 8718
rect 27649 8710 27679 8718
rect 27573 8684 27607 8710
rect 27645 8684 27679 8710
rect 27717 8684 27751 8718
rect 27789 8710 27819 8718
rect 27819 8710 27823 8718
rect 27789 8684 27823 8710
rect 27861 8684 27895 8718
rect 27501 8610 27535 8644
rect 27573 8640 27581 8644
rect 27581 8640 27607 8644
rect 27645 8640 27649 8644
rect 27649 8640 27679 8644
rect 27573 8610 27607 8640
rect 27645 8610 27679 8640
rect 27717 8610 27751 8644
rect 27789 8640 27819 8644
rect 27819 8640 27823 8644
rect 27789 8610 27823 8640
rect 27861 8610 27895 8644
rect 7266 8414 7300 8448
rect 7266 8341 7300 8375
rect 27272 8361 27306 8395
rect 27344 8361 27378 8395
rect 27416 8361 27450 8395
rect 27488 8361 27522 8395
rect 27560 8361 27594 8395
rect 27632 8361 27666 8395
rect 27704 8361 27738 8395
rect 27776 8361 27810 8395
rect 27848 8361 27882 8395
rect 27920 8361 27954 8395
rect 15709 8302 15743 8336
rect 15782 8302 15816 8336
rect 15855 8302 15889 8336
rect 15928 8302 15962 8336
rect 16000 8302 16034 8336
rect 16072 8302 16106 8336
rect 16144 8302 16178 8336
rect 16216 8302 16250 8336
rect 16288 8302 16322 8336
rect 16360 8302 16394 8336
rect 16432 8302 16466 8336
rect 16504 8302 16538 8336
rect 16576 8302 16610 8336
rect 7266 8268 7300 8302
rect 27272 8283 27306 8315
rect 27344 8283 27378 8315
rect 27416 8283 27450 8315
rect 27488 8283 27522 8315
rect 27560 8283 27594 8315
rect 27632 8283 27666 8315
rect 27704 8283 27738 8315
rect 27776 8283 27810 8315
rect 27272 8281 27304 8283
rect 27304 8281 27306 8283
rect 27344 8281 27372 8283
rect 27372 8281 27378 8283
rect 27416 8281 27440 8283
rect 27440 8281 27450 8283
rect 27488 8281 27508 8283
rect 27508 8281 27522 8283
rect 27560 8281 27576 8283
rect 27576 8281 27594 8283
rect 27632 8281 27644 8283
rect 27644 8281 27666 8283
rect 27704 8281 27712 8283
rect 27712 8281 27738 8283
rect 27776 8281 27780 8283
rect 27780 8281 27810 8283
rect 179 8052 213 8068
rect 257 8052 291 8068
rect 335 8052 369 8068
rect 413 8052 447 8068
rect 179 8034 209 8052
rect 209 8034 213 8052
rect 257 8034 279 8052
rect 279 8034 291 8052
rect 335 8034 349 8052
rect 349 8034 369 8052
rect 413 8034 419 8052
rect 419 8034 447 8052
rect 491 8034 525 8068
rect 569 8052 603 8068
rect 647 8052 681 8068
rect 725 8052 759 8068
rect 803 8052 837 8068
rect 569 8034 595 8052
rect 595 8034 603 8052
rect 647 8034 665 8052
rect 665 8034 681 8052
rect 725 8034 735 8052
rect 735 8034 759 8052
rect 803 8034 805 8052
rect 805 8034 837 8052
rect 179 7984 213 7996
rect 257 7984 291 7996
rect 335 7984 369 7996
rect 413 7984 447 7996
rect 179 7962 209 7984
rect 209 7962 213 7984
rect 257 7962 279 7984
rect 279 7962 291 7984
rect 335 7962 349 7984
rect 349 7962 369 7984
rect 413 7962 419 7984
rect 419 7962 447 7984
rect 491 7962 525 7996
rect 569 7984 603 7996
rect 647 7984 681 7996
rect 725 7984 759 7996
rect 803 7984 837 7996
rect 569 7962 595 7984
rect 595 7962 603 7984
rect 647 7962 665 7984
rect 665 7962 681 7984
rect 725 7962 735 7984
rect 735 7962 759 7984
rect 803 7962 805 7984
rect 805 7962 837 7984
rect 179 7915 213 7924
rect 257 7915 291 7924
rect 335 7915 369 7924
rect 413 7915 447 7924
rect 179 7890 209 7915
rect 209 7890 213 7915
rect 257 7890 279 7915
rect 279 7890 291 7915
rect 335 7890 349 7915
rect 349 7890 369 7915
rect 413 7890 419 7915
rect 419 7890 447 7915
rect 491 7890 525 7924
rect 569 7915 603 7924
rect 647 7915 681 7924
rect 725 7915 759 7924
rect 803 7915 837 7924
rect 569 7890 595 7915
rect 595 7890 603 7915
rect 647 7890 665 7915
rect 665 7890 681 7915
rect 725 7890 735 7915
rect 735 7890 759 7915
rect 803 7890 805 7915
rect 805 7890 837 7915
rect 179 7846 213 7852
rect 257 7846 291 7852
rect 335 7846 369 7852
rect 413 7846 447 7852
rect 179 7818 209 7846
rect 209 7818 213 7846
rect 257 7818 279 7846
rect 279 7818 291 7846
rect 335 7818 349 7846
rect 349 7818 369 7846
rect 413 7818 419 7846
rect 419 7818 447 7846
rect 491 7818 525 7852
rect 569 7846 603 7852
rect 647 7846 681 7852
rect 725 7846 759 7852
rect 803 7846 837 7852
rect 569 7818 595 7846
rect 595 7818 603 7846
rect 647 7818 665 7846
rect 665 7818 681 7846
rect 725 7818 735 7846
rect 735 7818 759 7846
rect 803 7818 805 7846
rect 805 7818 837 7846
rect 179 7777 213 7780
rect 257 7777 291 7780
rect 335 7777 369 7780
rect 413 7777 447 7780
rect 179 7746 209 7777
rect 209 7746 213 7777
rect 257 7746 279 7777
rect 279 7746 291 7777
rect 335 7746 349 7777
rect 349 7746 369 7777
rect 413 7746 419 7777
rect 419 7746 447 7777
rect 491 7746 525 7780
rect 569 7777 603 7780
rect 647 7777 681 7780
rect 725 7777 759 7780
rect 803 7777 837 7780
rect 569 7746 595 7777
rect 595 7746 603 7777
rect 647 7746 665 7777
rect 665 7746 681 7777
rect 725 7746 735 7777
rect 735 7746 759 7777
rect 803 7746 805 7777
rect 805 7746 837 7777
rect 179 7674 209 7707
rect 209 7674 213 7707
rect 257 7674 279 7707
rect 279 7674 291 7707
rect 335 7674 349 7707
rect 349 7674 369 7707
rect 413 7674 419 7707
rect 419 7674 447 7707
rect 179 7673 213 7674
rect 257 7673 291 7674
rect 335 7673 369 7674
rect 413 7673 447 7674
rect 491 7673 525 7707
rect 569 7674 595 7707
rect 595 7674 603 7707
rect 647 7674 665 7707
rect 665 7674 681 7707
rect 725 7674 735 7707
rect 735 7674 759 7707
rect 803 7674 805 7707
rect 805 7674 837 7707
rect 569 7673 603 7674
rect 647 7673 681 7674
rect 725 7673 759 7674
rect 803 7673 837 7674
rect 179 7605 209 7634
rect 209 7605 213 7634
rect 257 7605 279 7634
rect 279 7605 291 7634
rect 335 7605 349 7634
rect 349 7605 369 7634
rect 413 7605 419 7634
rect 419 7605 447 7634
rect 179 7600 213 7605
rect 257 7600 291 7605
rect 335 7600 369 7605
rect 413 7600 447 7605
rect 491 7600 525 7634
rect 569 7605 595 7634
rect 595 7605 603 7634
rect 647 7605 665 7634
rect 665 7605 681 7634
rect 725 7605 735 7634
rect 735 7605 759 7634
rect 803 7605 805 7634
rect 805 7605 837 7634
rect 569 7600 603 7605
rect 647 7600 681 7605
rect 725 7600 759 7605
rect 803 7600 837 7605
rect 179 7536 209 7561
rect 209 7536 213 7561
rect 257 7536 279 7561
rect 279 7536 291 7561
rect 335 7536 349 7561
rect 349 7536 369 7561
rect 413 7536 419 7561
rect 419 7536 447 7561
rect 179 7527 213 7536
rect 257 7527 291 7536
rect 335 7527 369 7536
rect 413 7527 447 7536
rect 491 7527 525 7561
rect 569 7536 595 7561
rect 595 7536 603 7561
rect 647 7536 665 7561
rect 665 7536 681 7561
rect 725 7536 735 7561
rect 735 7536 759 7561
rect 803 7536 805 7561
rect 805 7536 837 7561
rect 569 7527 603 7536
rect 647 7527 681 7536
rect 725 7527 759 7536
rect 803 7527 837 7536
rect 179 7467 209 7488
rect 209 7467 213 7488
rect 257 7467 279 7488
rect 279 7467 291 7488
rect 335 7467 349 7488
rect 349 7467 369 7488
rect 413 7467 419 7488
rect 419 7467 447 7488
rect 179 7454 213 7467
rect 257 7454 291 7467
rect 335 7454 369 7467
rect 413 7454 447 7467
rect 491 7454 525 7488
rect 569 7467 595 7488
rect 595 7467 603 7488
rect 647 7467 665 7488
rect 665 7467 681 7488
rect 725 7467 735 7488
rect 735 7467 759 7488
rect 803 7467 805 7488
rect 805 7467 837 7488
rect 569 7454 603 7467
rect 647 7454 681 7467
rect 725 7454 759 7467
rect 803 7454 837 7467
rect 179 7398 209 7415
rect 209 7398 213 7415
rect 257 7398 279 7415
rect 279 7398 291 7415
rect 335 7398 349 7415
rect 349 7398 369 7415
rect 413 7398 419 7415
rect 419 7398 447 7415
rect 179 7381 213 7398
rect 257 7381 291 7398
rect 335 7381 369 7398
rect 413 7381 447 7398
rect 491 7381 525 7415
rect 569 7398 595 7415
rect 595 7398 603 7415
rect 647 7398 665 7415
rect 665 7398 681 7415
rect 725 7398 735 7415
rect 735 7398 759 7415
rect 803 7398 805 7415
rect 805 7398 837 7415
rect 569 7381 603 7398
rect 647 7381 681 7398
rect 725 7381 759 7398
rect 803 7381 837 7398
rect 179 7329 209 7342
rect 209 7329 213 7342
rect 257 7329 279 7342
rect 279 7329 291 7342
rect 335 7329 349 7342
rect 349 7329 369 7342
rect 413 7329 419 7342
rect 419 7329 447 7342
rect 179 7308 213 7329
rect 257 7308 291 7329
rect 335 7308 369 7329
rect 413 7308 447 7329
rect 491 7308 525 7342
rect 569 7329 595 7342
rect 595 7329 603 7342
rect 647 7329 665 7342
rect 665 7329 681 7342
rect 725 7329 735 7342
rect 735 7329 759 7342
rect 803 7329 805 7342
rect 805 7329 837 7342
rect 569 7308 603 7329
rect 647 7308 681 7329
rect 725 7308 759 7329
rect 803 7308 837 7329
rect 179 7260 209 7269
rect 209 7260 213 7269
rect 257 7260 279 7269
rect 279 7260 291 7269
rect 335 7260 349 7269
rect 349 7260 369 7269
rect 413 7260 419 7269
rect 419 7260 447 7269
rect 179 7235 213 7260
rect 257 7235 291 7260
rect 335 7235 369 7260
rect 413 7235 447 7260
rect 491 7235 525 7269
rect 569 7260 595 7269
rect 595 7260 603 7269
rect 647 7260 665 7269
rect 665 7260 681 7269
rect 725 7260 735 7269
rect 735 7260 759 7269
rect 803 7260 805 7269
rect 805 7260 837 7269
rect 7091 8187 7125 8212
rect 7091 8178 7122 8187
rect 7122 8178 7125 8187
rect 7205 8187 7239 8212
rect 7205 8178 7212 8187
rect 7212 8178 7239 8187
rect 7091 8048 7125 8080
rect 7091 8046 7122 8048
rect 7122 8046 7125 8048
rect 7205 8048 7239 8080
rect 7205 8046 7212 8048
rect 7212 8046 7239 8048
rect 27848 8281 27882 8315
rect 27920 8281 27954 8315
rect 27272 8212 27306 8235
rect 27344 8212 27378 8235
rect 27416 8212 27450 8235
rect 27488 8212 27522 8235
rect 27560 8212 27594 8235
rect 27632 8212 27666 8235
rect 27704 8212 27738 8235
rect 27776 8212 27810 8235
rect 27272 8201 27304 8212
rect 27304 8201 27306 8212
rect 27344 8201 27372 8212
rect 27372 8201 27378 8212
rect 27416 8201 27440 8212
rect 27440 8201 27450 8212
rect 27488 8201 27508 8212
rect 27508 8201 27522 8212
rect 27560 8201 27576 8212
rect 27576 8201 27594 8212
rect 27632 8201 27644 8212
rect 27644 8201 27666 8212
rect 27704 8201 27712 8212
rect 27712 8201 27738 8212
rect 27776 8201 27780 8212
rect 27780 8201 27810 8212
rect 27848 8201 27882 8235
rect 27920 8201 27954 8235
rect 27272 8141 27306 8155
rect 27344 8141 27378 8155
rect 27416 8141 27450 8155
rect 27488 8141 27522 8155
rect 27560 8141 27594 8155
rect 27632 8141 27666 8155
rect 27704 8141 27738 8155
rect 27776 8141 27810 8155
rect 27272 8121 27304 8141
rect 27304 8121 27306 8141
rect 27344 8121 27372 8141
rect 27372 8121 27378 8141
rect 27416 8121 27440 8141
rect 27440 8121 27450 8141
rect 27488 8121 27508 8141
rect 27508 8121 27522 8141
rect 27560 8121 27576 8141
rect 27576 8121 27594 8141
rect 27632 8121 27644 8141
rect 27644 8121 27666 8141
rect 27704 8121 27712 8141
rect 27712 8121 27738 8141
rect 27776 8121 27780 8141
rect 27780 8121 27810 8141
rect 27848 8121 27882 8155
rect 27920 8121 27954 8155
rect 27272 8070 27306 8074
rect 27344 8070 27378 8074
rect 27416 8070 27450 8074
rect 27488 8070 27522 8074
rect 27560 8070 27594 8074
rect 27632 8070 27666 8074
rect 27704 8070 27738 8074
rect 27776 8070 27810 8074
rect 27272 8040 27304 8070
rect 27304 8040 27306 8070
rect 27344 8040 27372 8070
rect 27372 8040 27378 8070
rect 27416 8040 27440 8070
rect 27440 8040 27450 8070
rect 27488 8040 27508 8070
rect 27508 8040 27522 8070
rect 27560 8040 27576 8070
rect 27576 8040 27594 8070
rect 27632 8040 27644 8070
rect 27644 8040 27666 8070
rect 27704 8040 27712 8070
rect 27712 8040 27738 8070
rect 27776 8040 27780 8070
rect 27780 8040 27810 8070
rect 27848 8040 27882 8074
rect 27920 8040 27954 8074
rect 27272 7965 27304 7993
rect 27304 7965 27306 7993
rect 27344 7965 27372 7993
rect 27372 7965 27378 7993
rect 27416 7965 27440 7993
rect 27440 7965 27450 7993
rect 27488 7965 27508 7993
rect 27508 7965 27522 7993
rect 27560 7965 27576 7993
rect 27576 7965 27594 7993
rect 27632 7965 27644 7993
rect 27644 7965 27666 7993
rect 27704 7965 27712 7993
rect 27712 7965 27738 7993
rect 27776 7965 27780 7993
rect 27780 7965 27810 7993
rect 27272 7959 27306 7965
rect 27344 7959 27378 7965
rect 27416 7959 27450 7965
rect 27488 7959 27522 7965
rect 27560 7959 27594 7965
rect 27632 7959 27666 7965
rect 27704 7959 27738 7965
rect 27776 7959 27810 7965
rect 27848 7959 27882 7993
rect 27920 7959 27954 7993
rect 27272 7894 27304 7912
rect 27304 7894 27306 7912
rect 27344 7894 27372 7912
rect 27372 7894 27378 7912
rect 27416 7894 27440 7912
rect 27440 7894 27450 7912
rect 27488 7894 27508 7912
rect 27508 7894 27522 7912
rect 27560 7894 27576 7912
rect 27576 7894 27594 7912
rect 27632 7894 27644 7912
rect 27644 7894 27666 7912
rect 27704 7894 27712 7912
rect 27712 7894 27738 7912
rect 27776 7894 27780 7912
rect 27780 7894 27810 7912
rect 27272 7878 27306 7894
rect 27344 7878 27378 7894
rect 27416 7878 27450 7894
rect 27488 7878 27522 7894
rect 27560 7878 27594 7894
rect 27632 7878 27666 7894
rect 27704 7878 27738 7894
rect 27776 7878 27810 7894
rect 27848 7878 27882 7912
rect 27920 7878 27954 7912
rect 27272 7823 27304 7831
rect 27304 7823 27306 7831
rect 27344 7823 27372 7831
rect 27372 7823 27378 7831
rect 27416 7823 27440 7831
rect 27440 7823 27450 7831
rect 27488 7823 27508 7831
rect 27508 7823 27522 7831
rect 27560 7823 27576 7831
rect 27576 7823 27594 7831
rect 27632 7823 27644 7831
rect 27644 7823 27666 7831
rect 27704 7823 27712 7831
rect 27712 7823 27738 7831
rect 27776 7823 27780 7831
rect 27780 7823 27810 7831
rect 27272 7797 27306 7823
rect 27344 7797 27378 7823
rect 27416 7797 27450 7823
rect 27488 7797 27522 7823
rect 27560 7797 27594 7823
rect 27632 7797 27666 7823
rect 27704 7797 27738 7823
rect 27776 7797 27810 7823
rect 27848 7797 27882 7831
rect 27920 7797 27954 7831
rect 27272 7716 27306 7750
rect 27344 7716 27378 7750
rect 27416 7716 27450 7750
rect 27488 7716 27522 7750
rect 27560 7716 27594 7750
rect 27632 7716 27666 7750
rect 27704 7716 27738 7750
rect 27776 7716 27810 7750
rect 27848 7716 27882 7750
rect 27920 7716 27954 7750
rect 569 7235 603 7260
rect 647 7235 681 7260
rect 725 7235 759 7260
rect 803 7235 837 7260
rect 179 7191 209 7196
rect 209 7191 213 7196
rect 257 7191 279 7196
rect 279 7191 291 7196
rect 335 7191 349 7196
rect 349 7191 369 7196
rect 413 7191 419 7196
rect 419 7191 447 7196
rect 179 7162 213 7191
rect 257 7162 291 7191
rect 335 7162 369 7191
rect 413 7162 447 7191
rect 491 7162 525 7196
rect 569 7191 595 7196
rect 595 7191 603 7196
rect 647 7191 665 7196
rect 665 7191 681 7196
rect 725 7191 735 7196
rect 735 7191 759 7196
rect 803 7191 805 7196
rect 805 7191 837 7196
rect 569 7162 603 7191
rect 647 7162 681 7191
rect 725 7162 759 7191
rect 803 7162 837 7191
rect 179 7122 209 7123
rect 209 7122 213 7123
rect 257 7122 279 7123
rect 279 7122 291 7123
rect 335 7122 349 7123
rect 349 7122 369 7123
rect 413 7122 419 7123
rect 419 7122 447 7123
rect 179 7089 213 7122
rect 257 7089 291 7122
rect 335 7089 369 7122
rect 413 7089 447 7122
rect 491 7089 525 7123
rect 569 7122 595 7123
rect 595 7122 603 7123
rect 647 7122 665 7123
rect 665 7122 681 7123
rect 725 7122 735 7123
rect 735 7122 759 7123
rect 803 7122 805 7123
rect 805 7122 837 7123
rect 569 7089 603 7122
rect 647 7089 681 7122
rect 725 7089 759 7122
rect 803 7089 837 7122
rect 179 7018 213 7050
rect 257 7018 291 7050
rect 335 7018 369 7050
rect 413 7018 447 7050
rect 179 7016 209 7018
rect 209 7016 213 7018
rect 257 7016 279 7018
rect 279 7016 291 7018
rect 335 7016 349 7018
rect 349 7016 369 7018
rect 413 7016 419 7018
rect 419 7016 447 7018
rect 491 7016 525 7050
rect 569 7018 603 7050
rect 647 7018 681 7050
rect 725 7018 759 7050
rect 803 7018 837 7050
rect 569 7016 595 7018
rect 595 7016 603 7018
rect 647 7016 665 7018
rect 665 7016 681 7018
rect 725 7016 735 7018
rect 735 7016 759 7018
rect 803 7016 805 7018
rect 805 7016 837 7018
rect 179 6949 213 6977
rect 257 6949 291 6977
rect 335 6949 369 6977
rect 413 6949 447 6977
rect 179 6943 209 6949
rect 209 6943 213 6949
rect 257 6943 279 6949
rect 279 6943 291 6949
rect 335 6943 349 6949
rect 349 6943 369 6949
rect 413 6943 419 6949
rect 419 6943 447 6949
rect 491 6943 525 6977
rect 569 6949 603 6977
rect 647 6949 681 6977
rect 725 6949 759 6977
rect 803 6949 837 6977
rect 569 6943 595 6949
rect 595 6943 603 6949
rect 647 6943 665 6949
rect 665 6943 681 6949
rect 725 6943 735 6949
rect 735 6943 759 6949
rect 803 6943 805 6949
rect 805 6943 837 6949
rect 14263 7013 14441 7058
rect 14763 7013 15085 7058
rect 14263 6979 14296 7013
rect 14296 6979 14334 7013
rect 14334 6979 14368 7013
rect 14368 6979 14406 7013
rect 14406 6979 14440 7013
rect 14440 6979 14441 7013
rect 14763 6979 14766 7013
rect 14766 6979 14800 7013
rect 14800 6979 14838 7013
rect 14838 6979 14872 7013
rect 14872 6979 14910 7013
rect 14910 6979 14944 7013
rect 14944 6979 14982 7013
rect 14982 6979 15016 7013
rect 15016 6979 15054 7013
rect 15054 6979 15085 7013
rect 14263 6940 14441 6979
rect 14763 6940 15085 6979
rect 179 6880 213 6904
rect 257 6880 291 6904
rect 335 6880 369 6904
rect 413 6880 447 6904
rect 179 6870 209 6880
rect 209 6870 213 6880
rect 257 6870 279 6880
rect 279 6870 291 6880
rect 335 6870 349 6880
rect 349 6870 369 6880
rect 413 6870 419 6880
rect 419 6870 447 6880
rect 491 6870 525 6904
rect 569 6880 603 6904
rect 647 6880 681 6904
rect 725 6880 759 6904
rect 803 6880 837 6904
rect 569 6870 595 6880
rect 595 6870 603 6880
rect 647 6870 665 6880
rect 665 6870 681 6880
rect 725 6870 735 6880
rect 735 6870 759 6880
rect 803 6870 805 6880
rect 805 6870 837 6880
rect 179 6811 213 6831
rect 257 6811 291 6831
rect 335 6811 369 6831
rect 413 6811 447 6831
rect 179 6797 209 6811
rect 209 6797 213 6811
rect 257 6797 279 6811
rect 279 6797 291 6811
rect 335 6797 349 6811
rect 349 6797 369 6811
rect 413 6797 419 6811
rect 419 6797 447 6811
rect 491 6797 525 6831
rect 569 6811 603 6831
rect 647 6811 681 6831
rect 725 6811 759 6831
rect 803 6811 837 6831
rect 569 6797 595 6811
rect 595 6797 603 6811
rect 647 6797 665 6811
rect 665 6797 681 6811
rect 725 6797 735 6811
rect 735 6797 759 6811
rect 803 6797 805 6811
rect 805 6797 837 6811
rect 179 6742 213 6758
rect 257 6742 291 6758
rect 335 6742 369 6758
rect 413 6742 447 6758
rect 179 6724 209 6742
rect 209 6724 213 6742
rect 257 6724 279 6742
rect 279 6724 291 6742
rect 335 6724 349 6742
rect 349 6724 369 6742
rect 413 6724 419 6742
rect 419 6724 447 6742
rect 491 6724 525 6758
rect 569 6742 603 6758
rect 647 6742 681 6758
rect 725 6742 759 6758
rect 803 6742 837 6758
rect 569 6724 595 6742
rect 595 6724 603 6742
rect 647 6724 665 6742
rect 665 6724 681 6742
rect 725 6724 735 6742
rect 735 6724 759 6742
rect 803 6724 805 6742
rect 805 6724 837 6742
rect 179 6673 213 6685
rect 257 6673 291 6685
rect 335 6673 369 6685
rect 413 6673 447 6685
rect 179 6651 209 6673
rect 209 6651 213 6673
rect 257 6651 279 6673
rect 279 6651 291 6673
rect 335 6651 349 6673
rect 349 6651 369 6673
rect 413 6651 419 6673
rect 419 6651 447 6673
rect 491 6651 525 6685
rect 569 6673 603 6685
rect 647 6673 681 6685
rect 725 6673 759 6685
rect 803 6673 837 6685
rect 569 6651 595 6673
rect 595 6651 603 6673
rect 647 6651 665 6673
rect 665 6651 681 6673
rect 725 6651 735 6673
rect 735 6651 759 6673
rect 803 6651 805 6673
rect 805 6651 837 6673
rect 179 6604 213 6612
rect 257 6604 291 6612
rect 335 6604 369 6612
rect 413 6604 447 6612
rect 179 6578 209 6604
rect 209 6578 213 6604
rect 257 6578 279 6604
rect 279 6578 291 6604
rect 335 6578 349 6604
rect 349 6578 369 6604
rect 413 6578 419 6604
rect 419 6578 447 6604
rect 491 6578 525 6612
rect 569 6604 603 6612
rect 647 6604 681 6612
rect 725 6604 759 6612
rect 803 6604 837 6612
rect 569 6578 595 6604
rect 595 6578 603 6604
rect 647 6578 665 6604
rect 665 6578 681 6604
rect 725 6578 735 6604
rect 735 6578 759 6604
rect 803 6578 805 6604
rect 805 6578 837 6604
rect 179 6535 213 6539
rect 257 6535 291 6539
rect 335 6535 369 6539
rect 413 6535 447 6539
rect 179 6505 209 6535
rect 209 6505 213 6535
rect 257 6505 279 6535
rect 279 6505 291 6535
rect 335 6505 349 6535
rect 349 6505 369 6535
rect 413 6505 419 6535
rect 419 6505 447 6535
rect 491 6505 525 6539
rect 569 6535 603 6539
rect 647 6535 681 6539
rect 725 6535 759 6539
rect 803 6535 837 6539
rect 569 6505 595 6535
rect 595 6505 603 6535
rect 647 6505 665 6535
rect 665 6505 681 6535
rect 725 6505 735 6535
rect 735 6505 759 6535
rect 803 6505 805 6535
rect 805 6505 837 6535
rect 179 6432 209 6466
rect 209 6432 213 6466
rect 257 6432 279 6466
rect 279 6432 291 6466
rect 335 6432 349 6466
rect 349 6432 369 6466
rect 413 6432 419 6466
rect 419 6432 447 6466
rect 491 6432 525 6466
rect 569 6432 595 6466
rect 595 6432 603 6466
rect 647 6432 665 6466
rect 665 6432 681 6466
rect 725 6432 735 6466
rect 735 6432 759 6466
rect 803 6432 805 6466
rect 805 6432 837 6466
rect 179 6363 209 6393
rect 209 6363 213 6393
rect 257 6363 279 6393
rect 279 6363 291 6393
rect 335 6363 349 6393
rect 349 6363 369 6393
rect 413 6363 419 6393
rect 419 6363 447 6393
rect 179 6359 213 6363
rect 257 6359 291 6363
rect 335 6359 369 6363
rect 413 6359 447 6363
rect 491 6359 525 6393
rect 569 6363 595 6393
rect 595 6363 603 6393
rect 647 6363 665 6393
rect 665 6363 681 6393
rect 725 6363 735 6393
rect 735 6363 759 6393
rect 803 6363 805 6393
rect 805 6363 837 6393
rect 569 6359 603 6363
rect 647 6359 681 6363
rect 725 6359 759 6363
rect 803 6359 837 6363
rect 179 6294 209 6320
rect 209 6294 213 6320
rect 257 6294 279 6320
rect 279 6294 291 6320
rect 335 6294 349 6320
rect 349 6294 369 6320
rect 413 6294 419 6320
rect 419 6294 447 6320
rect 179 6286 213 6294
rect 257 6286 291 6294
rect 335 6286 369 6294
rect 413 6286 447 6294
rect 491 6286 525 6320
rect 569 6294 595 6320
rect 595 6294 603 6320
rect 647 6294 665 6320
rect 665 6294 681 6320
rect 725 6294 735 6320
rect 735 6294 759 6320
rect 803 6294 805 6320
rect 805 6294 837 6320
rect 569 6286 603 6294
rect 647 6286 681 6294
rect 725 6286 759 6294
rect 803 6286 837 6294
rect 14263 6906 14296 6940
rect 14296 6906 14334 6940
rect 14334 6906 14368 6940
rect 14368 6906 14406 6940
rect 14406 6906 14440 6940
rect 14440 6906 14441 6940
rect 14763 6906 14766 6940
rect 14766 6906 14800 6940
rect 14800 6906 14838 6940
rect 14838 6906 14872 6940
rect 14872 6906 14910 6940
rect 14910 6906 14944 6940
rect 14944 6906 14982 6940
rect 14982 6906 15016 6940
rect 15016 6906 15054 6940
rect 15054 6906 15085 6940
rect 14263 6866 14441 6906
rect 14763 6866 15085 6906
rect 13187 6815 13192 6828
rect 13192 6815 13221 6828
rect 13260 6815 13261 6828
rect 13261 6815 13294 6828
rect 13333 6815 13364 6828
rect 13364 6815 13367 6828
rect 13406 6815 13433 6828
rect 13433 6815 13440 6828
rect 13479 6815 13501 6828
rect 13501 6815 13513 6828
rect 13552 6815 13569 6828
rect 13569 6815 13586 6828
rect 13624 6815 13637 6828
rect 13637 6815 13658 6828
rect 13696 6815 13705 6828
rect 13705 6815 13730 6828
rect 13768 6815 13773 6828
rect 13773 6815 13802 6828
rect 13840 6815 13841 6828
rect 13841 6815 13874 6828
rect 13912 6815 13943 6828
rect 13943 6815 13946 6828
rect 14263 6832 14296 6866
rect 14296 6832 14334 6866
rect 14334 6832 14368 6866
rect 14368 6832 14406 6866
rect 14406 6832 14440 6866
rect 14440 6832 14441 6866
rect 14763 6832 14766 6866
rect 14766 6832 14800 6866
rect 14800 6832 14838 6866
rect 14838 6832 14872 6866
rect 14872 6832 14910 6866
rect 14910 6832 14944 6866
rect 14944 6832 14982 6866
rect 14982 6832 15016 6866
rect 15016 6832 15054 6866
rect 15054 6832 15085 6866
rect 13187 6794 13221 6815
rect 13260 6794 13294 6815
rect 13333 6794 13367 6815
rect 13406 6794 13440 6815
rect 13479 6794 13513 6815
rect 13552 6794 13586 6815
rect 13624 6794 13658 6815
rect 13696 6794 13730 6815
rect 13768 6794 13802 6815
rect 13840 6794 13874 6815
rect 13912 6794 13946 6815
rect 14263 6792 14441 6832
rect 14763 6792 15085 6832
rect 13187 6741 13192 6750
rect 13192 6741 13221 6750
rect 13260 6741 13261 6750
rect 13261 6741 13294 6750
rect 13333 6741 13364 6750
rect 13364 6741 13367 6750
rect 13406 6741 13433 6750
rect 13433 6741 13440 6750
rect 13479 6741 13501 6750
rect 13501 6741 13513 6750
rect 13552 6741 13569 6750
rect 13569 6741 13586 6750
rect 13624 6741 13637 6750
rect 13637 6741 13658 6750
rect 13696 6741 13705 6750
rect 13705 6741 13730 6750
rect 13768 6741 13773 6750
rect 13773 6741 13802 6750
rect 13840 6741 13841 6750
rect 13841 6741 13874 6750
rect 13912 6741 13943 6750
rect 13943 6741 13946 6750
rect 14263 6758 14296 6792
rect 14296 6758 14334 6792
rect 14334 6758 14368 6792
rect 14368 6758 14406 6792
rect 14406 6758 14440 6792
rect 14440 6758 14441 6792
rect 14763 6758 14766 6792
rect 14766 6758 14800 6792
rect 14800 6758 14838 6792
rect 14838 6758 14872 6792
rect 14872 6758 14910 6792
rect 14910 6758 14944 6792
rect 14944 6758 14982 6792
rect 14982 6758 15016 6792
rect 15016 6758 15054 6792
rect 15054 6758 15085 6792
rect 13187 6716 13221 6741
rect 13260 6716 13294 6741
rect 13333 6716 13367 6741
rect 13406 6716 13440 6741
rect 13479 6716 13513 6741
rect 13552 6716 13586 6741
rect 13624 6716 13658 6741
rect 13696 6716 13730 6741
rect 13768 6716 13802 6741
rect 13840 6716 13874 6741
rect 13912 6716 13946 6741
rect 14263 6718 14441 6758
rect 14763 6718 15085 6758
rect 13187 6667 13192 6672
rect 13192 6667 13221 6672
rect 13260 6667 13261 6672
rect 13261 6667 13294 6672
rect 13333 6667 13364 6672
rect 13364 6667 13367 6672
rect 13406 6667 13433 6672
rect 13433 6667 13440 6672
rect 13479 6667 13501 6672
rect 13501 6667 13513 6672
rect 13552 6667 13569 6672
rect 13569 6667 13586 6672
rect 13624 6667 13637 6672
rect 13637 6667 13658 6672
rect 13696 6667 13705 6672
rect 13705 6667 13730 6672
rect 13768 6667 13773 6672
rect 13773 6667 13802 6672
rect 13840 6667 13841 6672
rect 13841 6667 13874 6672
rect 13912 6667 13943 6672
rect 13943 6667 13946 6672
rect 14263 6684 14296 6718
rect 14296 6684 14334 6718
rect 14334 6684 14368 6718
rect 14368 6684 14406 6718
rect 14406 6684 14440 6718
rect 14440 6684 14441 6718
rect 14763 6684 14766 6718
rect 14766 6684 14800 6718
rect 14800 6684 14838 6718
rect 14838 6684 14872 6718
rect 14872 6684 14910 6718
rect 14910 6684 14944 6718
rect 14944 6684 14982 6718
rect 14982 6684 15016 6718
rect 15016 6684 15054 6718
rect 15054 6684 15085 6718
rect 13187 6638 13221 6667
rect 13260 6638 13294 6667
rect 13333 6638 13367 6667
rect 13406 6638 13440 6667
rect 13479 6638 13513 6667
rect 13552 6638 13586 6667
rect 13624 6638 13658 6667
rect 13696 6638 13730 6667
rect 13768 6638 13802 6667
rect 13840 6638 13874 6667
rect 13912 6638 13946 6667
rect 14263 6644 14441 6684
rect 14763 6644 15085 6684
rect 13187 6593 13192 6594
rect 13192 6593 13221 6594
rect 13260 6593 13261 6594
rect 13261 6593 13294 6594
rect 13333 6593 13364 6594
rect 13364 6593 13367 6594
rect 13406 6593 13433 6594
rect 13433 6593 13440 6594
rect 13479 6593 13501 6594
rect 13501 6593 13513 6594
rect 13552 6593 13569 6594
rect 13569 6593 13586 6594
rect 13624 6593 13637 6594
rect 13637 6593 13658 6594
rect 13696 6593 13705 6594
rect 13705 6593 13730 6594
rect 13768 6593 13773 6594
rect 13773 6593 13802 6594
rect 13840 6593 13841 6594
rect 13841 6593 13874 6594
rect 13912 6593 13943 6594
rect 13943 6593 13946 6594
rect 14263 6610 14296 6644
rect 14296 6610 14334 6644
rect 14334 6610 14368 6644
rect 14368 6610 14406 6644
rect 14406 6610 14440 6644
rect 14440 6610 14441 6644
rect 14763 6610 14766 6644
rect 14766 6610 14800 6644
rect 14800 6610 14838 6644
rect 14838 6610 14872 6644
rect 14872 6610 14910 6644
rect 14910 6610 14944 6644
rect 14944 6610 14982 6644
rect 14982 6610 15016 6644
rect 15016 6610 15054 6644
rect 15054 6610 15085 6644
rect 13187 6560 13221 6593
rect 13260 6560 13294 6593
rect 13333 6560 13367 6593
rect 13406 6560 13440 6593
rect 13479 6560 13513 6593
rect 13552 6560 13586 6593
rect 13624 6560 13658 6593
rect 13696 6560 13730 6593
rect 13768 6560 13802 6593
rect 13840 6560 13874 6593
rect 13912 6560 13946 6593
rect 14263 6570 14441 6610
rect 14763 6570 15085 6610
rect 14263 6536 14296 6570
rect 14296 6536 14334 6570
rect 14334 6536 14368 6570
rect 14368 6536 14406 6570
rect 14406 6536 14440 6570
rect 14440 6536 14441 6570
rect 14763 6536 14766 6570
rect 14766 6536 14800 6570
rect 14800 6536 14838 6570
rect 14838 6536 14872 6570
rect 14872 6536 14910 6570
rect 14910 6536 14944 6570
rect 14944 6536 14982 6570
rect 14982 6536 15016 6570
rect 15016 6536 15054 6570
rect 15054 6536 15085 6570
rect 13187 6482 13221 6516
rect 13260 6482 13294 6516
rect 13333 6482 13367 6516
rect 13406 6482 13440 6516
rect 13479 6482 13513 6516
rect 13552 6482 13586 6516
rect 13624 6482 13658 6516
rect 13696 6482 13730 6516
rect 13768 6482 13802 6516
rect 13840 6482 13874 6516
rect 13912 6482 13946 6516
rect 14263 6496 14441 6536
rect 14763 6496 15085 6536
rect 14263 6462 14296 6496
rect 14296 6462 14334 6496
rect 14334 6462 14368 6496
rect 14368 6462 14406 6496
rect 14406 6462 14440 6496
rect 14440 6462 14441 6496
rect 14763 6462 14766 6496
rect 14766 6462 14800 6496
rect 14800 6462 14838 6496
rect 14838 6462 14872 6496
rect 14872 6462 14910 6496
rect 14910 6462 14944 6496
rect 14944 6462 14982 6496
rect 14982 6462 15016 6496
rect 15016 6462 15054 6496
rect 15054 6462 15085 6496
rect 14263 6448 14441 6462
rect 14763 6448 15085 6462
rect 13187 6405 13221 6438
rect 13260 6405 13294 6438
rect 13333 6405 13367 6438
rect 13406 6405 13440 6438
rect 13479 6405 13513 6438
rect 13552 6405 13586 6438
rect 13624 6405 13658 6438
rect 13696 6405 13730 6438
rect 13768 6405 13802 6438
rect 13840 6405 13874 6438
rect 13912 6405 13946 6438
rect 13187 6404 13192 6405
rect 13192 6404 13221 6405
rect 13260 6404 13261 6405
rect 13261 6404 13294 6405
rect 13333 6404 13364 6405
rect 13364 6404 13367 6405
rect 13406 6404 13433 6405
rect 13433 6404 13440 6405
rect 13479 6404 13501 6405
rect 13501 6404 13513 6405
rect 13552 6404 13569 6405
rect 13569 6404 13586 6405
rect 13624 6404 13637 6405
rect 13637 6404 13658 6405
rect 13696 6404 13705 6405
rect 13705 6404 13730 6405
rect 13768 6404 13773 6405
rect 13773 6404 13802 6405
rect 13840 6404 13841 6405
rect 13841 6404 13874 6405
rect 13912 6404 13943 6405
rect 13943 6404 13946 6405
rect 14263 6388 14296 6409
rect 14296 6388 14297 6409
rect 14335 6388 14368 6409
rect 14368 6388 14369 6409
rect 14407 6388 14440 6409
rect 14440 6388 14441 6409
rect 14763 6388 14766 6409
rect 14766 6388 14797 6409
rect 14835 6388 14838 6409
rect 14838 6388 14869 6409
rect 14907 6388 14910 6409
rect 14910 6388 14941 6409
rect 14979 6388 14982 6409
rect 14982 6388 15013 6409
rect 15051 6388 15054 6409
rect 15054 6388 15085 6409
rect 14263 6375 14297 6388
rect 14335 6375 14369 6388
rect 14407 6375 14441 6388
rect 14763 6375 14797 6388
rect 14835 6375 14869 6388
rect 14907 6375 14941 6388
rect 14979 6375 15013 6388
rect 15051 6375 15085 6388
rect 13187 6331 13221 6360
rect 13260 6331 13294 6360
rect 13333 6331 13367 6360
rect 13406 6331 13440 6360
rect 13479 6331 13513 6360
rect 13552 6331 13586 6360
rect 13624 6331 13658 6360
rect 13696 6331 13730 6360
rect 13768 6331 13802 6360
rect 13840 6331 13874 6360
rect 13912 6331 13946 6360
rect 13187 6326 13192 6331
rect 13192 6326 13221 6331
rect 13260 6326 13261 6331
rect 13261 6326 13294 6331
rect 13333 6326 13364 6331
rect 13364 6326 13367 6331
rect 13406 6326 13433 6331
rect 13433 6326 13440 6331
rect 13479 6326 13501 6331
rect 13501 6326 13513 6331
rect 13552 6326 13569 6331
rect 13569 6326 13586 6331
rect 13624 6326 13637 6331
rect 13637 6326 13658 6331
rect 13696 6326 13705 6331
rect 13705 6326 13730 6331
rect 13768 6326 13773 6331
rect 13773 6326 13802 6331
rect 13840 6326 13841 6331
rect 13841 6326 13874 6331
rect 13912 6326 13943 6331
rect 13943 6326 13946 6331
rect 14263 6314 14296 6336
rect 14296 6314 14297 6336
rect 14335 6314 14368 6336
rect 14368 6314 14369 6336
rect 14407 6314 14440 6336
rect 14440 6314 14441 6336
rect 14763 6314 14766 6336
rect 14766 6314 14797 6336
rect 14835 6314 14838 6336
rect 14838 6314 14869 6336
rect 14907 6314 14910 6336
rect 14910 6314 14941 6336
rect 14979 6314 14982 6336
rect 14982 6314 15013 6336
rect 15051 6314 15054 6336
rect 15054 6314 15085 6336
rect 14263 6302 14297 6314
rect 14335 6302 14369 6314
rect 14407 6302 14441 6314
rect 14763 6302 14797 6314
rect 14835 6302 14869 6314
rect 14907 6302 14941 6314
rect 14979 6302 15013 6314
rect 15051 6302 15085 6314
rect 179 6225 209 6247
rect 209 6225 213 6247
rect 257 6225 279 6247
rect 279 6225 291 6247
rect 335 6225 349 6247
rect 349 6225 369 6247
rect 413 6225 419 6247
rect 419 6225 447 6247
rect 179 6213 213 6225
rect 257 6213 291 6225
rect 335 6213 369 6225
rect 413 6213 447 6225
rect 491 6213 525 6247
rect 569 6225 595 6247
rect 595 6225 603 6247
rect 647 6225 665 6247
rect 665 6225 681 6247
rect 725 6225 735 6247
rect 735 6225 759 6247
rect 803 6225 805 6247
rect 805 6225 837 6247
rect 569 6213 603 6225
rect 647 6213 681 6225
rect 725 6213 759 6225
rect 803 6213 837 6225
rect 173 6125 351 6166
rect 173 6091 203 6125
rect 203 6091 245 6125
rect 245 6091 279 6125
rect 279 6091 321 6125
rect 321 6091 351 6125
rect 173 6056 351 6091
rect 173 6022 203 6056
rect 203 6022 245 6056
rect 245 6022 279 6056
rect 279 6022 321 6056
rect 321 6022 351 6056
rect 173 5987 351 6022
rect 173 5953 203 5987
rect 203 5953 245 5987
rect 245 5953 279 5987
rect 279 5953 321 5987
rect 321 5953 351 5987
rect 173 5918 351 5953
rect 173 5884 203 5918
rect 203 5884 245 5918
rect 245 5884 279 5918
rect 279 5884 321 5918
rect 321 5884 351 5918
rect 173 5849 351 5884
rect 173 5815 203 5849
rect 203 5815 245 5849
rect 245 5815 279 5849
rect 279 5815 321 5849
rect 321 5815 351 5849
rect 173 5780 351 5815
rect 173 5746 203 5780
rect 203 5746 245 5780
rect 245 5746 279 5780
rect 279 5746 321 5780
rect 321 5746 351 5780
rect 173 5711 351 5746
rect 173 5677 203 5711
rect 203 5677 245 5711
rect 245 5677 279 5711
rect 279 5677 321 5711
rect 321 5677 351 5711
rect 173 5642 351 5677
rect 173 5608 203 5642
rect 203 5608 245 5642
rect 245 5608 279 5642
rect 279 5608 321 5642
rect 321 5608 351 5642
rect 173 5573 351 5608
rect 173 5539 203 5573
rect 203 5539 245 5573
rect 245 5539 279 5573
rect 279 5539 321 5573
rect 321 5539 351 5573
rect 173 5504 351 5539
rect 173 5470 203 5504
rect 203 5470 245 5504
rect 245 5470 279 5504
rect 279 5470 321 5504
rect 321 5470 351 5504
rect 173 5435 351 5470
rect 173 5401 203 5435
rect 203 5401 245 5435
rect 245 5401 279 5435
rect 279 5401 321 5435
rect 321 5401 351 5435
rect 173 5366 351 5401
rect 173 5332 203 5366
rect 203 5332 245 5366
rect 245 5332 279 5366
rect 279 5332 321 5366
rect 321 5332 351 5366
rect 173 5297 351 5332
rect 173 5263 203 5297
rect 203 5263 245 5297
rect 245 5263 279 5297
rect 279 5263 321 5297
rect 321 5263 351 5297
rect 173 5228 351 5263
rect 173 5194 203 5228
rect 203 5194 245 5228
rect 245 5194 279 5228
rect 279 5194 321 5228
rect 321 5194 351 5228
rect 173 5159 351 5194
rect 173 5125 203 5159
rect 203 5125 245 5159
rect 245 5125 279 5159
rect 279 5125 321 5159
rect 321 5125 351 5159
rect 173 5124 351 5125
rect 173 5056 203 5085
rect 203 5056 207 5085
rect 173 5051 207 5056
rect 245 5056 279 5085
rect 245 5051 279 5056
rect 317 5056 321 5085
rect 321 5056 351 5085
rect 317 5051 351 5056
rect 173 4987 203 5012
rect 203 4987 207 5012
rect 173 4978 207 4987
rect 245 4987 279 5012
rect 245 4978 279 4987
rect 317 4987 321 5012
rect 321 4987 351 5012
rect 317 4978 351 4987
rect 176 4124 210 4146
rect 254 4124 288 4146
rect 176 4112 203 4124
rect 203 4112 210 4124
rect 254 4112 279 4124
rect 279 4112 288 4124
rect 176 4055 210 4074
rect 254 4055 288 4074
rect 176 4040 203 4055
rect 203 4040 210 4055
rect 254 4040 279 4055
rect 279 4040 288 4055
rect 176 3986 210 4002
rect 254 3986 288 4002
rect 176 3968 203 3986
rect 203 3968 210 3986
rect 254 3968 279 3986
rect 279 3968 288 3986
rect 176 3917 210 3930
rect 254 3917 288 3930
rect 176 3896 203 3917
rect 203 3896 210 3917
rect 254 3896 279 3917
rect 279 3896 288 3917
rect 176 3848 210 3858
rect 254 3848 288 3858
rect 176 3824 203 3848
rect 203 3824 210 3848
rect 254 3824 279 3848
rect 279 3824 288 3848
rect 176 3779 210 3786
rect 254 3779 288 3786
rect 176 3752 203 3779
rect 203 3752 210 3779
rect 254 3752 279 3779
rect 279 3752 288 3779
rect 176 3710 210 3714
rect 254 3710 288 3714
rect 176 3680 203 3710
rect 203 3680 210 3710
rect 254 3680 279 3710
rect 279 3680 288 3710
rect 176 3641 210 3642
rect 254 3641 288 3642
rect 176 3608 203 3641
rect 203 3608 210 3641
rect 254 3608 279 3641
rect 279 3608 288 3641
rect 176 3537 203 3570
rect 203 3537 210 3570
rect 254 3537 279 3570
rect 279 3537 288 3570
rect 176 3536 210 3537
rect 254 3536 288 3537
rect 176 3467 203 3497
rect 203 3467 210 3497
rect 254 3467 279 3497
rect 279 3467 288 3497
rect 176 3463 210 3467
rect 254 3463 288 3467
rect 176 3397 203 3424
rect 203 3397 210 3424
rect 254 3397 279 3424
rect 279 3397 288 3424
rect 176 3390 210 3397
rect 254 3390 288 3397
rect 176 3327 203 3351
rect 203 3327 210 3351
rect 254 3327 279 3351
rect 279 3327 288 3351
rect 176 3317 210 3327
rect 254 3317 288 3327
rect 176 3257 203 3278
rect 203 3257 210 3278
rect 254 3257 279 3278
rect 279 3257 288 3278
rect 176 3244 210 3257
rect 254 3244 288 3257
rect 176 3187 203 3205
rect 203 3187 210 3205
rect 254 3187 279 3205
rect 279 3187 288 3205
rect 176 3171 210 3187
rect 254 3171 288 3187
rect 176 3117 203 3132
rect 203 3117 210 3132
rect 254 3117 279 3132
rect 279 3117 288 3132
rect 176 3098 210 3117
rect 254 3098 288 3117
rect 1356 3603 1390 3637
rect 1436 3603 1470 3637
rect 1516 3603 1550 3637
rect 1596 3603 1630 3637
rect 1676 3603 1710 3637
rect 1755 3603 1789 3637
rect 1834 3603 1868 3637
rect 1913 3603 1947 3637
rect 1992 3603 2026 3637
rect 2071 3603 2105 3637
rect 1356 3527 1390 3561
rect 1436 3527 1470 3561
rect 1516 3527 1550 3561
rect 1596 3527 1630 3561
rect 1676 3527 1710 3561
rect 1755 3527 1789 3561
rect 1834 3527 1868 3561
rect 1913 3527 1947 3561
rect 1992 3527 2026 3561
rect 2071 3527 2105 3561
rect 1356 3451 1390 3485
rect 1436 3451 1470 3485
rect 1516 3451 1550 3485
rect 1596 3451 1630 3485
rect 1676 3451 1710 3485
rect 1755 3451 1789 3485
rect 1834 3451 1868 3485
rect 1913 3451 1947 3485
rect 1992 3451 2026 3485
rect 2071 3451 2105 3485
rect 176 3047 203 3059
rect 203 3047 210 3059
rect 254 3047 279 3059
rect 279 3047 288 3059
rect 176 3025 210 3047
rect 254 3025 288 3047
rect 176 2977 203 2986
rect 203 2977 210 2986
rect 254 2977 279 2986
rect 279 2977 288 2986
rect 341 2977 355 3000
rect 355 2977 375 3000
rect 415 2979 444 3000
rect 444 2979 449 3000
rect 489 2979 515 3000
rect 515 2979 523 3000
rect 563 2979 586 3000
rect 586 2979 597 3000
rect 637 2979 657 3000
rect 657 2979 671 3000
rect 711 2979 728 3000
rect 728 2979 745 3000
rect 785 2979 799 3000
rect 799 2979 819 3000
rect 859 2979 869 3000
rect 869 2979 893 3000
rect 933 2979 939 3000
rect 939 2979 967 3000
rect 1006 2979 1009 3000
rect 1009 2979 1040 3000
rect 176 2952 210 2977
rect 254 2952 288 2977
rect 341 2966 375 2977
rect 415 2966 449 2979
rect 489 2966 523 2979
rect 563 2966 597 2979
rect 637 2966 671 2979
rect 711 2966 745 2979
rect 785 2966 819 2979
rect 859 2966 893 2979
rect 933 2966 967 2979
rect 1006 2966 1040 2979
rect 2700 2977 2701 3011
rect 2701 2977 2734 3011
rect 2778 2977 2803 3011
rect 2803 2977 2812 3011
rect 2856 2977 2871 3011
rect 2871 2977 2890 3011
rect 2934 2977 2939 3011
rect 2939 2977 2968 3011
rect 3012 2977 3041 3011
rect 3041 2977 3046 3011
rect 3090 2977 3109 3011
rect 3109 2977 3124 3011
rect 2700 2903 2701 2935
rect 2701 2903 2734 2935
rect 2778 2903 2803 2935
rect 2803 2903 2812 2935
rect 2856 2903 2871 2935
rect 2871 2903 2890 2935
rect 2934 2903 2939 2935
rect 2939 2903 2968 2935
rect 3012 2903 3041 2935
rect 3041 2903 3046 2935
rect 3090 2903 3109 2935
rect 3109 2903 3124 2935
rect 2700 2901 2734 2903
rect 2778 2901 2812 2903
rect 2856 2901 2890 2903
rect 2934 2901 2968 2903
rect 3012 2901 3046 2903
rect 3090 2901 3124 2903
rect 341 2837 355 2866
rect 355 2837 375 2866
rect 415 2865 449 2866
rect 489 2865 523 2866
rect 563 2865 597 2866
rect 637 2865 671 2866
rect 711 2865 745 2866
rect 785 2865 819 2866
rect 859 2865 893 2866
rect 933 2865 967 2866
rect 1006 2865 1040 2866
rect 341 2832 375 2837
rect 415 2832 444 2865
rect 444 2832 449 2865
rect 489 2832 515 2865
rect 515 2832 523 2865
rect 563 2832 586 2865
rect 586 2832 597 2865
rect 637 2832 657 2865
rect 657 2832 671 2865
rect 711 2832 728 2865
rect 728 2832 745 2865
rect 785 2832 799 2865
rect 799 2832 819 2865
rect 859 2832 869 2865
rect 869 2832 893 2865
rect 933 2832 939 2865
rect 939 2832 967 2865
rect 1006 2832 1009 2865
rect 1009 2832 1040 2865
rect 2700 2829 2701 2859
rect 2701 2829 2734 2859
rect 2778 2829 2803 2859
rect 2803 2829 2812 2859
rect 2856 2829 2871 2859
rect 2871 2829 2890 2859
rect 2934 2829 2939 2859
rect 2939 2829 2968 2859
rect 3012 2829 3041 2859
rect 3041 2829 3046 2859
rect 3090 2829 3109 2859
rect 3109 2829 3124 2859
rect 2700 2825 2734 2829
rect 2778 2825 2812 2829
rect 2856 2825 2890 2829
rect 2934 2825 2968 2829
rect 3012 2825 3046 2829
rect 3090 2825 3124 2829
rect 2700 2755 2701 2783
rect 2701 2755 2734 2783
rect 2778 2755 2803 2783
rect 2803 2755 2812 2783
rect 2856 2755 2871 2783
rect 2871 2755 2890 2783
rect 2934 2755 2939 2783
rect 2939 2755 2968 2783
rect 3012 2755 3041 2783
rect 3041 2755 3046 2783
rect 3090 2755 3109 2783
rect 3109 2755 3124 2783
rect 2700 2749 2734 2755
rect 2778 2749 2812 2755
rect 2856 2749 2890 2755
rect 2934 2749 2968 2755
rect 3012 2749 3046 2755
rect 3090 2749 3124 2755
rect 1958 2681 1984 2686
rect 1984 2681 1992 2686
rect 2034 2681 2053 2686
rect 2053 2681 2068 2686
rect 2110 2681 2122 2686
rect 2122 2681 2144 2686
rect 2186 2681 2191 2686
rect 2191 2681 2220 2686
rect 2262 2681 2293 2686
rect 2293 2681 2296 2686
rect 2338 2681 2361 2686
rect 2361 2681 2372 2686
rect 2414 2681 2429 2686
rect 2429 2681 2448 2686
rect 2490 2681 2497 2686
rect 2497 2681 2524 2686
rect 1958 2652 1992 2681
rect 2034 2652 2068 2681
rect 2110 2652 2144 2681
rect 2186 2652 2220 2681
rect 2262 2652 2296 2681
rect 2338 2652 2372 2681
rect 2414 2652 2448 2681
rect 2490 2652 2524 2681
rect 2565 2652 2599 2686
rect 2640 2681 2667 2686
rect 2667 2681 2674 2686
rect 2715 2681 2735 2686
rect 2735 2681 2749 2686
rect 2790 2681 2803 2686
rect 2803 2681 2824 2686
rect 2865 2681 2871 2686
rect 2871 2681 2899 2686
rect 2940 2681 2973 2686
rect 2973 2681 2974 2686
rect 3015 2681 3041 2686
rect 3041 2681 3049 2686
rect 3090 2681 3109 2686
rect 3109 2681 3124 2686
rect 2640 2652 2674 2681
rect 2715 2652 2749 2681
rect 2790 2652 2824 2681
rect 2865 2652 2899 2681
rect 2940 2652 2974 2681
rect 3015 2652 3049 2681
rect 3090 2652 3124 2681
rect 1958 2567 1992 2576
rect 2034 2567 2068 2576
rect 2110 2567 2144 2576
rect 2186 2567 2220 2576
rect 2262 2567 2296 2576
rect 2338 2567 2372 2576
rect 2414 2567 2448 2576
rect 2490 2567 2524 2576
rect 1958 2542 1984 2567
rect 1984 2542 1992 2567
rect 2034 2542 2053 2567
rect 2053 2542 2068 2567
rect 2110 2542 2122 2567
rect 2122 2542 2144 2567
rect 2186 2542 2191 2567
rect 2191 2542 2220 2567
rect 2262 2542 2293 2567
rect 2293 2542 2296 2567
rect 2338 2542 2361 2567
rect 2361 2542 2372 2567
rect 2414 2542 2429 2567
rect 2429 2542 2448 2567
rect 2490 2542 2497 2567
rect 2497 2542 2524 2567
rect 2565 2542 2599 2576
rect 2640 2567 2674 2576
rect 2715 2567 2749 2576
rect 2790 2567 2824 2576
rect 2865 2567 2899 2576
rect 2940 2567 2974 2576
rect 3015 2567 3049 2576
rect 3090 2567 3124 2576
rect 2640 2542 2667 2567
rect 2667 2542 2674 2567
rect 2715 2542 2735 2567
rect 2735 2542 2749 2567
rect 2790 2542 2803 2567
rect 2803 2542 2824 2567
rect 2865 2542 2871 2567
rect 2871 2542 2899 2567
rect 2940 2542 2973 2567
rect 2973 2542 2974 2567
rect 3015 2542 3041 2567
rect 3041 2542 3049 2567
rect 3090 2542 3109 2567
rect 3109 2542 3124 2567
rect 25855 1999 25880 2019
rect 25880 1999 25889 2019
rect 25928 1999 25951 2019
rect 25951 1999 25962 2019
rect 26001 1999 26022 2019
rect 26022 1999 26035 2019
rect 26074 1999 26093 2019
rect 26093 1999 26108 2019
rect 26147 1999 26164 2019
rect 26164 1999 26181 2019
rect 26220 1999 26235 2019
rect 26235 1999 26254 2019
rect 26293 1999 26306 2019
rect 26306 1999 26327 2019
rect 26366 1999 26376 2019
rect 26376 1999 26400 2019
rect 26439 1999 26446 2019
rect 26446 1999 26473 2019
rect 26512 1999 26516 2019
rect 26516 1999 26546 2019
rect 26585 1999 26586 2019
rect 26586 1999 26619 2019
rect 25855 1985 25889 1999
rect 25928 1985 25962 1999
rect 26001 1985 26035 1999
rect 26074 1985 26108 1999
rect 26147 1985 26181 1999
rect 26220 1985 26254 1999
rect 26293 1985 26327 1999
rect 26366 1985 26400 1999
rect 26439 1985 26473 1999
rect 26512 1985 26546 1999
rect 26585 1985 26619 1999
rect 26658 1985 26692 2019
rect 26731 1999 26762 2019
rect 26762 1999 26765 2019
rect 26804 1999 26832 2019
rect 26832 1999 26838 2019
rect 26877 1999 26902 2019
rect 26902 1999 26911 2019
rect 26950 1999 26972 2019
rect 26972 1999 26984 2019
rect 27022 1999 27042 2019
rect 27042 1999 27056 2019
rect 27094 1999 27112 2019
rect 27112 1999 27128 2019
rect 27166 1999 27182 2019
rect 27182 1999 27200 2019
rect 27238 1999 27252 2019
rect 27252 1999 27272 2019
rect 27310 1999 27322 2019
rect 27322 1999 27344 2019
rect 27382 1999 27392 2019
rect 27392 1999 27416 2019
rect 27454 1999 27462 2019
rect 27462 1999 27488 2019
rect 27526 1999 27532 2019
rect 27532 1999 27560 2019
rect 27598 1999 27602 2019
rect 27602 1999 27632 2019
rect 27670 1999 27672 2019
rect 27672 1999 27704 2019
rect 27742 1999 27776 2019
rect 27814 1999 27846 2019
rect 27846 1999 27848 2019
rect 26731 1985 26765 1999
rect 26804 1985 26838 1999
rect 26877 1985 26911 1999
rect 26950 1985 26984 1999
rect 27022 1985 27056 1999
rect 27094 1985 27128 1999
rect 27166 1985 27200 1999
rect 27238 1985 27272 1999
rect 27310 1985 27344 1999
rect 27382 1985 27416 1999
rect 27454 1985 27488 1999
rect 27526 1985 27560 1999
rect 27598 1985 27632 1999
rect 27670 1985 27704 1999
rect 27742 1985 27776 1999
rect 27814 1985 27848 1999
rect 25855 1913 25880 1939
rect 25880 1913 25889 1939
rect 25928 1913 25951 1939
rect 25951 1913 25962 1939
rect 26001 1913 26022 1939
rect 26022 1913 26035 1939
rect 26074 1913 26093 1939
rect 26093 1913 26108 1939
rect 26147 1913 26164 1939
rect 26164 1913 26181 1939
rect 26220 1913 26235 1939
rect 26235 1913 26254 1939
rect 26293 1913 26306 1939
rect 26306 1913 26327 1939
rect 26366 1913 26376 1939
rect 26376 1913 26400 1939
rect 26439 1913 26446 1939
rect 26446 1913 26473 1939
rect 26512 1913 26516 1939
rect 26516 1913 26546 1939
rect 26585 1913 26586 1939
rect 26586 1913 26619 1939
rect 25855 1905 25889 1913
rect 25928 1905 25962 1913
rect 26001 1905 26035 1913
rect 26074 1905 26108 1913
rect 26147 1905 26181 1913
rect 26220 1905 26254 1913
rect 26293 1905 26327 1913
rect 26366 1905 26400 1913
rect 26439 1905 26473 1913
rect 26512 1905 26546 1913
rect 26585 1905 26619 1913
rect 26658 1905 26692 1939
rect 26731 1913 26762 1939
rect 26762 1913 26765 1939
rect 26804 1913 26832 1939
rect 26832 1913 26838 1939
rect 26877 1913 26902 1939
rect 26902 1913 26911 1939
rect 26950 1913 26972 1939
rect 26972 1913 26984 1939
rect 27022 1913 27042 1939
rect 27042 1913 27056 1939
rect 27094 1913 27112 1939
rect 27112 1913 27128 1939
rect 27166 1913 27182 1939
rect 27182 1913 27200 1939
rect 27238 1913 27252 1939
rect 27252 1913 27272 1939
rect 27310 1913 27322 1939
rect 27322 1913 27344 1939
rect 27382 1913 27392 1939
rect 27392 1913 27416 1939
rect 27454 1913 27462 1939
rect 27462 1913 27488 1939
rect 27526 1913 27532 1939
rect 27532 1913 27560 1939
rect 27598 1913 27602 1939
rect 27602 1913 27632 1939
rect 27670 1913 27672 1939
rect 27672 1913 27704 1939
rect 27742 1913 27776 1939
rect 27814 1913 27846 1939
rect 27846 1913 27848 1939
rect 26731 1905 26765 1913
rect 26804 1905 26838 1913
rect 26877 1905 26911 1913
rect 26950 1905 26984 1913
rect 27022 1905 27056 1913
rect 27094 1905 27128 1913
rect 27166 1905 27200 1913
rect 27238 1905 27272 1913
rect 27310 1905 27344 1913
rect 27382 1905 27416 1913
rect 27454 1905 27488 1913
rect 27526 1905 27560 1913
rect 27598 1905 27632 1913
rect 27670 1905 27704 1913
rect 27742 1905 27776 1913
rect 27814 1905 27848 1913
rect 25855 1827 25880 1859
rect 25880 1827 25889 1859
rect 25928 1827 25951 1859
rect 25951 1827 25962 1859
rect 26001 1827 26022 1859
rect 26022 1827 26035 1859
rect 26074 1827 26093 1859
rect 26093 1827 26108 1859
rect 26147 1827 26164 1859
rect 26164 1827 26181 1859
rect 26220 1827 26235 1859
rect 26235 1827 26254 1859
rect 26293 1827 26306 1859
rect 26306 1827 26327 1859
rect 26366 1827 26376 1859
rect 26376 1827 26400 1859
rect 26439 1827 26446 1859
rect 26446 1827 26473 1859
rect 26512 1827 26516 1859
rect 26516 1827 26546 1859
rect 26585 1827 26586 1859
rect 26586 1827 26619 1859
rect 25855 1825 25889 1827
rect 25928 1825 25962 1827
rect 26001 1825 26035 1827
rect 26074 1825 26108 1827
rect 26147 1825 26181 1827
rect 26220 1825 26254 1827
rect 26293 1825 26327 1827
rect 26366 1825 26400 1827
rect 26439 1825 26473 1827
rect 26512 1825 26546 1827
rect 26585 1825 26619 1827
rect 26658 1825 26692 1859
rect 26731 1827 26762 1859
rect 26762 1827 26765 1859
rect 26804 1827 26832 1859
rect 26832 1827 26838 1859
rect 26877 1827 26902 1859
rect 26902 1827 26911 1859
rect 26950 1827 26972 1859
rect 26972 1827 26984 1859
rect 27022 1827 27042 1859
rect 27042 1827 27056 1859
rect 27094 1827 27112 1859
rect 27112 1827 27128 1859
rect 27166 1827 27182 1859
rect 27182 1827 27200 1859
rect 27238 1827 27252 1859
rect 27252 1827 27272 1859
rect 27310 1827 27322 1859
rect 27322 1827 27344 1859
rect 27382 1827 27392 1859
rect 27392 1827 27416 1859
rect 27454 1827 27462 1859
rect 27462 1827 27488 1859
rect 27526 1827 27532 1859
rect 27532 1827 27560 1859
rect 27598 1827 27602 1859
rect 27602 1827 27632 1859
rect 27670 1827 27672 1859
rect 27672 1827 27704 1859
rect 27742 1827 27776 1859
rect 27814 1827 27846 1859
rect 27846 1827 27848 1859
rect 26731 1825 26765 1827
rect 26804 1825 26838 1827
rect 26877 1825 26911 1827
rect 26950 1825 26984 1827
rect 27022 1825 27056 1827
rect 27094 1825 27128 1827
rect 27166 1825 27200 1827
rect 27238 1825 27272 1827
rect 27310 1825 27344 1827
rect 27382 1825 27416 1827
rect 27454 1825 27488 1827
rect 27526 1825 27560 1827
rect 27598 1825 27632 1827
rect 27670 1825 27704 1827
rect 27742 1825 27776 1827
rect 27814 1825 27848 1827
rect 25855 1775 25889 1779
rect 25928 1775 25962 1779
rect 26001 1775 26035 1779
rect 26074 1775 26108 1779
rect 26147 1775 26181 1779
rect 26220 1775 26254 1779
rect 26293 1775 26327 1779
rect 26366 1775 26400 1779
rect 26439 1775 26473 1779
rect 26512 1775 26546 1779
rect 26585 1775 26619 1779
rect 25855 1745 25880 1775
rect 25880 1745 25889 1775
rect 25928 1745 25951 1775
rect 25951 1745 25962 1775
rect 26001 1745 26022 1775
rect 26022 1745 26035 1775
rect 26074 1745 26093 1775
rect 26093 1745 26108 1775
rect 26147 1745 26164 1775
rect 26164 1745 26181 1775
rect 26220 1745 26235 1775
rect 26235 1745 26254 1775
rect 26293 1745 26306 1775
rect 26306 1745 26327 1775
rect 26366 1745 26376 1775
rect 26376 1745 26400 1775
rect 26439 1745 26446 1775
rect 26446 1745 26473 1775
rect 26512 1745 26516 1775
rect 26516 1745 26546 1775
rect 26585 1745 26586 1775
rect 26586 1745 26619 1775
rect 26658 1745 26692 1779
rect 26731 1775 26765 1779
rect 26804 1775 26838 1779
rect 26877 1775 26911 1779
rect 26950 1775 26984 1779
rect 27022 1775 27056 1779
rect 27094 1775 27128 1779
rect 27166 1775 27200 1779
rect 27238 1775 27272 1779
rect 27310 1775 27344 1779
rect 27382 1775 27416 1779
rect 27454 1775 27488 1779
rect 27526 1775 27560 1779
rect 27598 1775 27632 1779
rect 27670 1775 27704 1779
rect 27742 1775 27776 1779
rect 27814 1775 27848 1779
rect 26731 1745 26762 1775
rect 26762 1745 26765 1775
rect 26804 1745 26832 1775
rect 26832 1745 26838 1775
rect 26877 1745 26902 1775
rect 26902 1745 26911 1775
rect 26950 1745 26972 1775
rect 26972 1745 26984 1775
rect 27022 1745 27042 1775
rect 27042 1745 27056 1775
rect 27094 1745 27112 1775
rect 27112 1745 27128 1775
rect 27166 1745 27182 1775
rect 27182 1745 27200 1775
rect 27238 1745 27252 1775
rect 27252 1745 27272 1775
rect 27310 1745 27322 1775
rect 27322 1745 27344 1775
rect 27382 1745 27392 1775
rect 27392 1745 27416 1775
rect 27454 1745 27462 1775
rect 27462 1745 27488 1775
rect 27526 1745 27532 1775
rect 27532 1745 27560 1775
rect 27598 1745 27602 1775
rect 27602 1745 27632 1775
rect 27670 1745 27672 1775
rect 27672 1745 27704 1775
rect 27742 1745 27776 1775
rect 27814 1745 27846 1775
rect 27846 1745 27848 1775
<< metal1 >>
rect 86 39912 214 39924
rect 86 39878 92 39912
rect 126 39878 174 39912
rect 208 39878 214 39912
rect 86 39840 214 39878
rect 86 39806 92 39840
rect 126 39806 174 39840
rect 208 39806 214 39840
rect 86 39768 214 39806
rect 86 39734 92 39768
rect 126 39734 174 39768
rect 208 39734 214 39768
rect 86 39696 214 39734
rect 86 39662 92 39696
rect 126 39662 174 39696
rect 208 39662 214 39696
rect 86 39624 214 39662
rect 86 39590 92 39624
rect 126 39590 174 39624
rect 208 39590 214 39624
rect 86 39552 214 39590
rect 86 39518 92 39552
rect 126 39518 174 39552
rect 208 39518 214 39552
rect 86 39480 214 39518
rect 86 39446 92 39480
rect 126 39446 174 39480
rect 208 39446 214 39480
rect 86 39408 214 39446
rect 86 39374 92 39408
rect 126 39374 174 39408
rect 208 39374 214 39408
rect 86 39336 214 39374
rect 86 39302 92 39336
rect 126 39302 174 39336
rect 208 39302 214 39336
rect 86 39264 214 39302
rect 86 39230 92 39264
rect 126 39230 174 39264
rect 208 39230 214 39264
rect 86 39192 214 39230
rect 86 39158 92 39192
rect 126 39158 174 39192
rect 208 39158 214 39192
rect 86 39120 214 39158
rect 86 39086 92 39120
rect 126 39086 174 39120
rect 208 39086 214 39120
rect 86 39048 214 39086
rect 86 39014 92 39048
rect 126 39014 174 39048
rect 208 39014 214 39048
rect 86 38976 214 39014
rect 86 38942 92 38976
rect 126 38942 174 38976
rect 208 38942 214 38976
rect 86 38904 214 38942
rect 86 38870 92 38904
rect 126 38870 174 38904
rect 208 38870 214 38904
rect 86 38832 214 38870
rect 86 38798 92 38832
rect 126 38798 174 38832
rect 208 38798 214 38832
rect 86 38760 214 38798
rect 86 38726 92 38760
rect 126 38726 174 38760
rect 208 38726 214 38760
rect 86 38688 214 38726
rect 86 38654 92 38688
rect 126 38654 174 38688
rect 208 38654 214 38688
rect 86 38616 214 38654
rect 86 38582 92 38616
rect 126 38582 174 38616
rect 208 38582 214 38616
rect 86 38544 214 38582
rect 86 38510 92 38544
rect 126 38510 174 38544
rect 208 38510 214 38544
rect 86 38472 214 38510
rect 86 38438 92 38472
rect 126 38438 174 38472
rect 208 38438 214 38472
rect 86 38400 214 38438
rect 86 38366 92 38400
rect 126 38366 174 38400
rect 208 38366 214 38400
rect 86 38328 214 38366
rect 86 38294 92 38328
rect 126 38294 174 38328
rect 208 38294 214 38328
rect 86 38256 214 38294
rect 86 38222 92 38256
rect 126 38222 174 38256
rect 208 38222 214 38256
rect 86 38184 214 38222
rect 86 38150 92 38184
rect 126 38150 174 38184
rect 208 38150 214 38184
rect 86 38111 214 38150
rect 86 38077 92 38111
rect 126 38077 174 38111
rect 208 38077 214 38111
rect 86 38038 214 38077
rect 86 38004 92 38038
rect 126 38004 174 38038
rect 208 38004 214 38038
rect 86 37842 214 38004
tri 86 37836 92 37842 ne
rect 92 37836 214 37842
tri 214 37836 285 37907 sw
tri 92 37804 124 37836 ne
rect 124 37804 331 37836
tri 124 37770 158 37804 ne
rect 158 37770 209 37804
rect 243 37770 291 37804
rect 325 37770 331 37804
tri 158 37732 196 37770 ne
rect 196 37732 331 37770
tri 196 37725 203 37732 ne
rect 203 37698 209 37732
rect 243 37698 291 37732
rect 325 37698 331 37732
rect 203 37660 331 37698
rect 203 37626 209 37660
rect 243 37626 291 37660
rect 325 37626 331 37660
rect 203 37588 331 37626
rect 203 37554 209 37588
rect 243 37554 291 37588
rect 325 37554 331 37588
rect 203 37516 331 37554
rect 203 37482 209 37516
rect 243 37482 291 37516
rect 325 37482 331 37516
rect 203 37444 331 37482
rect 203 37410 209 37444
rect 243 37410 291 37444
rect 325 37410 331 37444
rect 203 37372 331 37410
rect 203 37338 209 37372
rect 243 37338 291 37372
rect 325 37338 331 37372
rect 203 37300 331 37338
rect 203 37266 209 37300
rect 243 37266 291 37300
rect 325 37266 331 37300
rect 203 37228 331 37266
rect 203 37194 209 37228
rect 243 37194 291 37228
rect 325 37194 331 37228
rect 203 37156 331 37194
rect 203 37122 209 37156
rect 243 37122 291 37156
rect 325 37122 331 37156
rect 203 37084 331 37122
rect 203 37050 209 37084
rect 243 37050 291 37084
rect 325 37050 331 37084
rect 203 37012 331 37050
rect 203 36978 209 37012
rect 243 36978 291 37012
rect 325 36978 331 37012
rect 203 36940 331 36978
rect 203 36906 209 36940
rect 243 36906 291 36940
rect 325 36906 331 36940
rect 203 36868 331 36906
rect 203 36834 209 36868
rect 243 36834 291 36868
rect 325 36834 331 36868
rect 203 36796 331 36834
rect 203 36762 209 36796
rect 243 36762 291 36796
rect 325 36762 331 36796
rect 203 36724 331 36762
rect 203 36690 209 36724
rect 243 36690 291 36724
rect 325 36690 331 36724
rect 203 36652 331 36690
rect 203 36618 209 36652
rect 243 36618 291 36652
rect 325 36618 331 36652
rect 203 36580 331 36618
rect 203 36546 209 36580
rect 243 36546 291 36580
rect 325 36546 331 36580
rect 203 36508 331 36546
rect 17645 36836 17763 36842
rect 17697 36784 17711 36836
rect 17645 36758 17763 36784
rect 17697 36706 17711 36758
rect 17645 36679 17763 36706
rect 17697 36627 17711 36679
rect 17645 36600 17763 36627
rect 17697 36548 17711 36600
rect 17645 36542 17763 36548
rect 203 36474 209 36508
rect 243 36474 291 36508
rect 325 36474 331 36508
rect 203 36436 331 36474
rect 203 36402 209 36436
rect 243 36402 291 36436
rect 325 36402 331 36436
rect 203 36364 331 36402
rect 203 36330 209 36364
rect 243 36330 291 36364
rect 325 36330 331 36364
rect 203 36292 331 36330
rect 203 36258 209 36292
rect 243 36258 291 36292
rect 325 36258 331 36292
rect 203 36220 331 36258
rect 203 36186 209 36220
rect 243 36186 291 36220
rect 325 36186 331 36220
tri 22680 36416 22750 36486 sw
rect 22680 36384 23279 36416
rect 22680 36350 22829 36384
rect 22863 36350 22911 36384
rect 22945 36350 22993 36384
rect 23027 36350 23075 36384
rect 23109 36350 23157 36384
rect 23191 36350 23239 36384
rect 23273 36350 23279 36384
rect 22680 36312 23279 36350
rect 22680 36278 22829 36312
rect 22863 36278 22911 36312
rect 22945 36278 22993 36312
rect 23027 36278 23075 36312
rect 23109 36278 23157 36312
rect 23191 36278 23239 36312
rect 23273 36278 23279 36312
rect 22680 36240 23279 36278
rect 22680 36210 22829 36240
tri 22744 36206 22748 36210 ne
rect 22748 36206 22829 36210
rect 22863 36206 22911 36240
rect 22945 36206 22993 36240
rect 23027 36206 23075 36240
rect 23109 36206 23157 36240
rect 23191 36206 23239 36240
rect 23273 36206 23279 36240
rect 203 36148 331 36186
tri 22748 36168 22786 36206 ne
rect 22786 36168 23279 36206
rect 203 36114 209 36148
rect 243 36114 291 36148
rect 325 36114 331 36148
tri 22786 36134 22820 36168 ne
rect 22820 36134 22829 36168
rect 22863 36134 22911 36168
rect 22945 36134 22993 36168
rect 23027 36134 23075 36168
rect 23109 36134 23157 36168
rect 23191 36134 23239 36168
rect 23273 36134 23279 36168
tri 22820 36131 22823 36134 ne
rect 203 36076 331 36114
rect 203 36042 209 36076
rect 243 36042 291 36076
rect 325 36042 331 36076
rect 203 36004 331 36042
rect 203 35970 209 36004
rect 243 35970 291 36004
rect 325 35970 331 36004
rect 203 35932 331 35970
rect 203 35898 209 35932
rect 243 35898 291 35932
rect 325 35898 331 35932
rect 203 35860 331 35898
rect 203 35826 209 35860
rect 243 35826 291 35860
rect 325 35826 331 35860
rect 203 35788 331 35826
rect 203 35754 209 35788
rect 243 35754 291 35788
rect 325 35754 331 35788
rect 203 35716 331 35754
rect 203 35682 209 35716
rect 243 35682 291 35716
rect 325 35682 331 35716
rect 203 35644 331 35682
rect 203 35610 209 35644
rect 243 35610 291 35644
rect 325 35610 331 35644
rect 203 35572 331 35610
rect 203 35538 209 35572
rect 243 35538 291 35572
rect 325 35538 331 35572
rect 203 35500 331 35538
rect 203 35466 209 35500
rect 243 35466 291 35500
rect 325 35466 331 35500
rect 203 35427 331 35466
rect 203 35393 209 35427
rect 243 35393 291 35427
rect 325 35393 331 35427
rect 203 35354 331 35393
rect 203 35320 209 35354
rect 243 35320 291 35354
rect 325 35320 331 35354
rect 203 35281 331 35320
rect 203 35247 209 35281
rect 243 35247 291 35281
rect 325 35247 331 35281
rect 203 35208 331 35247
rect 203 35174 209 35208
rect 243 35174 291 35208
rect 325 35174 331 35208
rect 203 35135 331 35174
rect 203 35101 209 35135
rect 243 35101 291 35135
rect 325 35101 331 35135
rect 203 35062 331 35101
rect 203 35028 209 35062
rect 243 35028 291 35062
rect 325 35028 331 35062
rect 203 34989 331 35028
rect 203 34955 209 34989
rect 243 34955 291 34989
rect 325 34955 331 34989
rect 203 34916 331 34955
rect 203 34882 209 34916
rect 243 34882 291 34916
rect 325 34882 331 34916
rect 203 34843 331 34882
rect 203 34809 209 34843
rect 243 34809 291 34843
rect 325 34809 331 34843
rect 203 34770 331 34809
rect 203 34736 209 34770
rect 243 34736 291 34770
rect 325 34736 331 34770
rect 203 34697 331 34736
rect 203 34663 209 34697
rect 243 34663 291 34697
rect 325 34663 331 34697
rect 203 34624 331 34663
rect 203 34590 209 34624
rect 243 34590 291 34624
rect 325 34590 331 34624
rect 203 34551 331 34590
rect 203 34517 209 34551
rect 243 34517 291 34551
rect 325 34517 331 34551
rect 203 34478 331 34517
rect 203 34444 209 34478
rect 243 34444 291 34478
rect 325 34444 331 34478
rect 203 34405 331 34444
rect 203 34371 209 34405
rect 243 34371 291 34405
rect 325 34371 331 34405
rect 203 34332 331 34371
rect 203 34298 209 34332
rect 243 34298 291 34332
rect 325 34298 331 34332
rect 203 34259 331 34298
rect 203 34225 209 34259
rect 243 34225 291 34259
rect 325 34225 331 34259
rect 203 34186 331 34225
rect 203 34152 209 34186
rect 243 34152 291 34186
rect 325 34152 331 34186
rect 203 34113 331 34152
rect 203 34079 209 34113
rect 243 34079 291 34113
rect 325 34079 331 34113
rect 203 34040 331 34079
rect 203 34006 209 34040
rect 243 34006 291 34040
rect 325 34006 331 34040
rect 203 33967 331 34006
rect 203 33933 209 33967
rect 243 33933 291 33967
rect 325 33933 331 33967
rect 203 33894 331 33933
rect 203 33860 209 33894
rect 243 33860 291 33894
rect 325 33860 331 33894
rect 203 33821 331 33860
rect 203 33787 209 33821
rect 243 33787 291 33821
rect 325 33787 331 33821
rect 203 33748 331 33787
rect 203 33714 209 33748
rect 243 33714 291 33748
rect 325 33714 331 33748
rect 203 33675 331 33714
rect 203 33641 209 33675
rect 243 33641 291 33675
rect 325 33641 331 33675
rect 203 33602 331 33641
rect 203 33568 209 33602
rect 243 33568 291 33602
rect 325 33568 331 33602
rect 203 33529 331 33568
rect 203 33495 209 33529
rect 243 33495 291 33529
rect 325 33495 331 33529
rect 203 33456 331 33495
rect 203 33422 209 33456
rect 243 33422 291 33456
rect 325 33422 331 33456
rect 203 33383 331 33422
rect 203 33349 209 33383
rect 243 33349 291 33383
rect 325 33349 331 33383
rect 203 33310 331 33349
rect 22823 36096 23279 36134
rect 22823 36062 22829 36096
rect 22863 36062 22911 36096
rect 22945 36062 22993 36096
rect 23027 36062 23075 36096
rect 23109 36062 23157 36096
rect 23191 36062 23239 36096
rect 23273 36062 23279 36096
rect 22823 36024 23279 36062
rect 22823 35990 22829 36024
rect 22863 35990 22911 36024
rect 22945 35990 22993 36024
rect 23027 35990 23075 36024
rect 23109 35990 23157 36024
rect 23191 35990 23239 36024
rect 23273 35990 23279 36024
rect 22823 35952 23279 35990
rect 22823 35918 22829 35952
rect 22863 35918 22911 35952
rect 22945 35918 22993 35952
rect 23027 35918 23075 35952
rect 23109 35918 23157 35952
rect 23191 35918 23239 35952
rect 23273 35918 23279 35952
rect 22823 35880 23279 35918
rect 22823 35846 22829 35880
rect 22863 35846 22911 35880
rect 22945 35846 22993 35880
rect 23027 35846 23075 35880
rect 23109 35846 23157 35880
rect 23191 35846 23239 35880
rect 23273 35846 23279 35880
rect 22823 35808 23279 35846
rect 22823 35774 22829 35808
rect 22863 35774 22911 35808
rect 22945 35774 22993 35808
rect 23027 35774 23075 35808
rect 23109 35774 23157 35808
rect 23191 35774 23239 35808
rect 23273 35774 23279 35808
rect 22823 35736 23279 35774
rect 22823 35702 22829 35736
rect 22863 35702 22911 35736
rect 22945 35702 22993 35736
rect 23027 35702 23075 35736
rect 23109 35702 23157 35736
rect 23191 35702 23239 35736
rect 23273 35702 23279 35736
rect 22823 35664 23279 35702
rect 22823 35630 22829 35664
rect 22863 35630 22911 35664
rect 22945 35630 22993 35664
rect 23027 35630 23075 35664
rect 23109 35630 23157 35664
rect 23191 35630 23239 35664
rect 23273 35630 23279 35664
rect 22823 35592 23279 35630
rect 22823 35558 22829 35592
rect 22863 35558 22911 35592
rect 22945 35558 22993 35592
rect 23027 35558 23075 35592
rect 23109 35558 23157 35592
rect 23191 35558 23239 35592
rect 23273 35558 23279 35592
rect 22823 35520 23279 35558
rect 22823 35486 22829 35520
rect 22863 35486 22911 35520
rect 22945 35486 22993 35520
rect 23027 35486 23075 35520
rect 23109 35486 23157 35520
rect 23191 35486 23239 35520
rect 23273 35486 23279 35520
rect 22823 35448 23279 35486
rect 22823 35414 22829 35448
rect 22863 35414 22911 35448
rect 22945 35414 22993 35448
rect 23027 35414 23075 35448
rect 23109 35414 23157 35448
rect 23191 35414 23239 35448
rect 23273 35414 23279 35448
rect 22823 35376 23279 35414
rect 22823 35342 22829 35376
rect 22863 35342 22911 35376
rect 22945 35342 22993 35376
rect 23027 35342 23075 35376
rect 23109 35342 23157 35376
rect 23191 35342 23239 35376
rect 23273 35342 23279 35376
rect 22823 35304 23279 35342
rect 22823 35270 22829 35304
rect 22863 35270 22911 35304
rect 22945 35270 22993 35304
rect 23027 35270 23075 35304
rect 23109 35270 23157 35304
rect 23191 35270 23239 35304
rect 23273 35270 23279 35304
rect 22823 35232 23279 35270
rect 22823 35198 22829 35232
rect 22863 35198 22911 35232
rect 22945 35198 22993 35232
rect 23027 35198 23075 35232
rect 23109 35198 23157 35232
rect 23191 35198 23239 35232
rect 23273 35198 23279 35232
rect 22823 35160 23279 35198
rect 22823 35126 22829 35160
rect 22863 35126 22911 35160
rect 22945 35126 22993 35160
rect 23027 35126 23075 35160
rect 23109 35126 23157 35160
rect 23191 35126 23239 35160
rect 23273 35126 23279 35160
rect 22823 35088 23279 35126
rect 22823 35054 22829 35088
rect 22863 35054 22911 35088
rect 22945 35054 22993 35088
rect 23027 35054 23075 35088
rect 23109 35054 23157 35088
rect 23191 35054 23239 35088
rect 23273 35054 23279 35088
rect 22823 35016 23279 35054
rect 22823 34982 22829 35016
rect 22863 34982 22911 35016
rect 22945 34982 22993 35016
rect 23027 34982 23075 35016
rect 23109 34982 23157 35016
rect 23191 34982 23239 35016
rect 23273 34982 23279 35016
rect 22823 34944 23279 34982
rect 22823 34910 22829 34944
rect 22863 34910 22911 34944
rect 22945 34910 22993 34944
rect 23027 34910 23075 34944
rect 23109 34910 23157 34944
rect 23191 34910 23239 34944
rect 23273 34910 23279 34944
rect 22823 34872 23279 34910
rect 22823 34838 22829 34872
rect 22863 34838 22911 34872
rect 22945 34838 22993 34872
rect 23027 34838 23075 34872
rect 23109 34838 23157 34872
rect 23191 34838 23239 34872
rect 23273 34838 23279 34872
rect 22823 34800 23279 34838
rect 22823 34766 22829 34800
rect 22863 34766 22911 34800
rect 22945 34766 22993 34800
rect 23027 34766 23075 34800
rect 23109 34766 23157 34800
rect 23191 34766 23239 34800
rect 23273 34766 23279 34800
rect 22823 34728 23279 34766
rect 22823 34694 22829 34728
rect 22863 34694 22911 34728
rect 22945 34694 22993 34728
rect 23027 34694 23075 34728
rect 23109 34694 23157 34728
rect 23191 34694 23239 34728
rect 23273 34694 23279 34728
rect 22823 34656 23279 34694
rect 22823 34622 22829 34656
rect 22863 34622 22911 34656
rect 22945 34622 22993 34656
rect 23027 34622 23075 34656
rect 23109 34622 23157 34656
rect 23191 34622 23239 34656
rect 23273 34622 23279 34656
rect 22823 34584 23279 34622
rect 22823 34550 22829 34584
rect 22863 34550 22911 34584
rect 22945 34550 22993 34584
rect 23027 34550 23075 34584
rect 23109 34550 23157 34584
rect 23191 34550 23239 34584
rect 23273 34550 23279 34584
rect 22823 34512 23279 34550
rect 22823 34478 22829 34512
rect 22863 34478 22911 34512
rect 22945 34478 22993 34512
rect 23027 34478 23075 34512
rect 23109 34478 23157 34512
rect 23191 34478 23239 34512
rect 23273 34478 23279 34512
rect 22823 34440 23279 34478
rect 22823 34406 22829 34440
rect 22863 34406 22911 34440
rect 22945 34406 22993 34440
rect 23027 34406 23075 34440
rect 23109 34406 23157 34440
rect 23191 34406 23239 34440
rect 23273 34406 23279 34440
rect 22823 34368 23279 34406
rect 22823 34334 22829 34368
rect 22863 34334 22911 34368
rect 22945 34334 22993 34368
rect 23027 34334 23075 34368
rect 23109 34334 23157 34368
rect 23191 34334 23239 34368
rect 23273 34334 23279 34368
rect 22823 34295 23279 34334
rect 22823 34261 22829 34295
rect 22863 34261 22911 34295
rect 22945 34261 22993 34295
rect 23027 34261 23075 34295
rect 23109 34261 23157 34295
rect 23191 34261 23239 34295
rect 23273 34261 23279 34295
rect 22823 34222 23279 34261
rect 22823 34188 22829 34222
rect 22863 34188 22911 34222
rect 22945 34188 22993 34222
rect 23027 34188 23075 34222
rect 23109 34188 23157 34222
rect 23191 34188 23239 34222
rect 23273 34188 23279 34222
rect 22823 34149 23279 34188
rect 22823 34115 22829 34149
rect 22863 34115 22911 34149
rect 22945 34115 22993 34149
rect 23027 34115 23075 34149
rect 23109 34115 23157 34149
rect 23191 34115 23239 34149
rect 23273 34115 23279 34149
rect 22823 34076 23279 34115
rect 22823 34042 22829 34076
rect 22863 34042 22911 34076
rect 22945 34042 22993 34076
rect 23027 34042 23075 34076
rect 23109 34042 23157 34076
rect 23191 34042 23239 34076
rect 23273 34042 23279 34076
rect 22823 34003 23279 34042
rect 22823 33969 22829 34003
rect 22863 33969 22911 34003
rect 22945 33969 22993 34003
rect 23027 33969 23075 34003
rect 23109 33969 23157 34003
rect 23191 33969 23239 34003
rect 23273 33969 23279 34003
rect 22823 33930 23279 33969
rect 22823 33896 22829 33930
rect 22863 33896 22911 33930
rect 22945 33896 22993 33930
rect 23027 33896 23075 33930
rect 23109 33896 23157 33930
rect 23191 33896 23239 33930
rect 23273 33896 23279 33930
rect 22823 33857 23279 33896
rect 22823 33823 22829 33857
rect 22863 33823 22911 33857
rect 22945 33823 22993 33857
rect 23027 33823 23075 33857
rect 23109 33823 23157 33857
rect 23191 33823 23239 33857
rect 23273 33823 23279 33857
rect 22823 33784 23279 33823
rect 22823 33750 22829 33784
rect 22863 33750 22911 33784
rect 22945 33750 22993 33784
rect 23027 33750 23075 33784
rect 23109 33750 23157 33784
rect 23191 33750 23239 33784
rect 23273 33750 23279 33784
rect 22823 33711 23279 33750
rect 22823 33677 22829 33711
rect 22863 33677 22911 33711
rect 22945 33677 22993 33711
rect 23027 33677 23075 33711
rect 23109 33677 23157 33711
rect 23191 33677 23239 33711
rect 23273 33677 23279 33711
rect 22823 33638 23279 33677
rect 22823 33604 22829 33638
rect 22863 33604 22911 33638
rect 22945 33604 22993 33638
rect 23027 33604 23075 33638
rect 23109 33604 23157 33638
rect 23191 33604 23239 33638
rect 23273 33604 23279 33638
rect 22823 33565 23279 33604
rect 22823 33531 22829 33565
rect 22863 33531 22911 33565
rect 22945 33531 22993 33565
rect 23027 33531 23075 33565
rect 23109 33531 23157 33565
rect 23191 33531 23239 33565
rect 23273 33531 23279 33565
rect 22823 33492 23279 33531
rect 22823 33458 22829 33492
rect 22863 33458 22911 33492
rect 22945 33458 22993 33492
rect 23027 33458 23075 33492
rect 23109 33458 23157 33492
rect 23191 33458 23239 33492
rect 23273 33458 23279 33492
rect 22823 33419 23279 33458
rect 22823 33385 22829 33419
rect 22863 33385 22911 33419
rect 22945 33385 22993 33419
rect 23027 33385 23075 33419
rect 23109 33385 23157 33419
rect 23191 33385 23239 33419
rect 23273 33385 23279 33419
rect 22823 33346 23279 33385
rect 203 33276 209 33310
rect 243 33276 291 33310
rect 325 33276 331 33310
rect 203 33237 331 33276
rect 203 33203 209 33237
rect 243 33203 291 33237
rect 325 33203 331 33237
rect 203 33164 331 33203
rect 203 33130 209 33164
rect 243 33130 291 33164
rect 325 33130 331 33164
rect 203 33091 331 33130
rect 203 33057 209 33091
rect 243 33057 291 33091
rect 325 33057 331 33091
rect 203 33018 331 33057
rect 203 32984 209 33018
rect 243 32984 291 33018
rect 325 32984 331 33018
rect 203 32945 331 32984
rect 203 32911 209 32945
rect 243 32911 291 32945
rect 325 32911 331 32945
rect 203 32872 331 32911
rect 203 32838 209 32872
rect 243 32838 291 32872
rect 325 32838 331 32872
rect 203 32799 331 32838
rect 203 32765 209 32799
rect 243 32765 291 32799
rect 325 32765 331 32799
rect 203 32726 331 32765
rect 203 32692 209 32726
rect 243 32692 291 32726
rect 325 32692 331 32726
rect 203 32653 331 32692
rect 203 32619 209 32653
rect 243 32619 291 32653
rect 325 32619 331 32653
rect 203 32580 331 32619
rect 203 32546 209 32580
rect 243 32546 291 32580
rect 325 32546 331 32580
rect 203 32507 331 32546
rect 203 32473 209 32507
rect 243 32473 291 32507
rect 325 32473 331 32507
rect 203 32434 331 32473
rect 203 32400 209 32434
rect 243 32400 291 32434
rect 325 32400 331 32434
rect 203 32361 331 32400
rect 203 32327 209 32361
rect 243 32327 291 32361
rect 325 32327 331 32361
rect 203 32288 331 32327
rect 203 32254 209 32288
rect 243 32254 291 32288
rect 325 32254 331 32288
rect 203 32215 331 32254
rect 203 32181 209 32215
rect 243 32181 291 32215
rect 325 32181 331 32215
rect 203 32142 331 32181
rect 203 32108 209 32142
rect 243 32108 291 32142
rect 325 32108 331 32142
rect 203 32070 331 32108
rect 18015 33328 18407 33340
rect 18015 33294 18022 33328
rect 18056 33294 18108 33328
rect 18142 33294 18194 33328
rect 18228 33294 18280 33328
rect 18314 33294 18366 33328
rect 18400 33294 18407 33328
rect 18015 33256 18407 33294
rect 18015 33222 18022 33256
rect 18056 33222 18108 33256
rect 18142 33222 18194 33256
rect 18228 33222 18280 33256
rect 18314 33222 18366 33256
rect 18400 33222 18407 33256
rect 18015 33184 18407 33222
rect 18015 33150 18022 33184
rect 18056 33150 18108 33184
rect 18142 33150 18194 33184
rect 18228 33150 18280 33184
rect 18314 33150 18366 33184
rect 18400 33150 18407 33184
rect 18015 33112 18407 33150
rect 18015 33078 18022 33112
rect 18056 33078 18108 33112
rect 18142 33078 18194 33112
rect 18228 33078 18280 33112
rect 18314 33078 18366 33112
rect 18400 33078 18407 33112
rect 18015 33040 18407 33078
rect 18015 33006 18022 33040
rect 18056 33006 18108 33040
rect 18142 33006 18194 33040
rect 18228 33006 18280 33040
rect 18314 33006 18366 33040
rect 18400 33006 18407 33040
rect 18015 32968 18407 33006
rect 18015 32934 18022 32968
rect 18056 32934 18108 32968
rect 18142 32934 18194 32968
rect 18228 32934 18280 32968
rect 18314 32934 18366 32968
rect 18400 32934 18407 32968
rect 18015 32896 18407 32934
rect 18015 32862 18022 32896
rect 18056 32862 18108 32896
rect 18142 32862 18194 32896
rect 18228 32862 18280 32896
rect 18314 32862 18366 32896
rect 18400 32862 18407 32896
rect 18015 32824 18407 32862
rect 18015 32818 18022 32824
rect 18056 32818 18108 32824
rect 18142 32818 18194 32824
rect 18015 32766 18018 32818
rect 18070 32790 18108 32818
rect 18180 32790 18194 32818
rect 18228 32790 18280 32824
rect 18314 32790 18366 32824
rect 18400 32790 18407 32824
rect 18070 32766 18128 32790
rect 18180 32766 18407 32790
rect 18015 32752 18407 32766
rect 18015 32751 18022 32752
rect 18056 32751 18108 32752
rect 18142 32751 18194 32752
rect 18015 32699 18018 32751
rect 18070 32718 18108 32751
rect 18180 32718 18194 32751
rect 18228 32718 18280 32752
rect 18314 32718 18366 32752
rect 18400 32718 18407 32752
rect 18070 32699 18128 32718
rect 18180 32699 18407 32718
rect 18015 32684 18407 32699
rect 18015 32632 18018 32684
rect 18070 32680 18128 32684
rect 18180 32680 18407 32684
rect 18070 32646 18108 32680
rect 18180 32646 18194 32680
rect 18228 32646 18280 32680
rect 18314 32646 18366 32680
rect 18400 32646 18407 32680
rect 18070 32632 18128 32646
rect 18180 32632 18407 32646
rect 18015 32617 18407 32632
rect 18015 32565 18018 32617
rect 18070 32608 18128 32617
rect 18180 32608 18407 32617
rect 18070 32574 18108 32608
rect 18180 32574 18194 32608
rect 18228 32574 18280 32608
rect 18314 32574 18366 32608
rect 18400 32574 18407 32608
rect 18070 32565 18128 32574
rect 18180 32565 18407 32574
rect 18015 32550 18407 32565
rect 18015 32498 18018 32550
rect 18070 32536 18128 32550
rect 18180 32536 18407 32550
rect 18070 32502 18108 32536
rect 18180 32502 18194 32536
rect 18228 32502 18280 32536
rect 18314 32502 18366 32536
rect 18400 32502 18407 32536
rect 18070 32498 18128 32502
rect 18180 32498 18407 32502
rect 18015 32482 18407 32498
rect 18015 32430 18018 32482
rect 18070 32464 18128 32482
rect 18180 32464 18407 32482
rect 18070 32430 18108 32464
rect 18180 32430 18194 32464
rect 18228 32430 18280 32464
rect 18314 32430 18366 32464
rect 18400 32430 18407 32464
rect 18015 32414 18407 32430
rect 18015 32362 18018 32414
rect 18070 32392 18128 32414
rect 18180 32392 18407 32414
rect 18070 32362 18108 32392
rect 18180 32362 18194 32392
rect 18015 32358 18022 32362
rect 18056 32358 18108 32362
rect 18142 32358 18194 32362
rect 18228 32358 18280 32392
rect 18314 32358 18366 32392
rect 18400 32358 18407 32392
rect 18015 32346 18407 32358
rect 18015 32294 18018 32346
rect 18070 32320 18128 32346
rect 18180 32320 18407 32346
rect 18070 32294 18108 32320
rect 18180 32294 18194 32320
rect 18015 32286 18022 32294
rect 18056 32286 18108 32294
rect 18142 32286 18194 32294
rect 18228 32286 18280 32320
rect 18314 32286 18366 32320
rect 18400 32286 18407 32320
rect 18015 32278 18407 32286
rect 18015 32226 18018 32278
rect 18070 32248 18128 32278
rect 18180 32248 18407 32278
rect 18070 32226 18108 32248
rect 18180 32226 18194 32248
rect 18015 32214 18022 32226
rect 18056 32214 18108 32226
rect 18142 32214 18194 32226
rect 18228 32214 18280 32248
rect 18314 32214 18366 32248
rect 18400 32214 18407 32248
rect 18015 32210 18407 32214
rect 18015 32158 18018 32210
rect 18070 32176 18128 32210
rect 18180 32176 18407 32210
rect 18070 32158 18108 32176
rect 18180 32158 18194 32176
rect 18015 32142 18022 32158
rect 18056 32142 18108 32158
rect 18142 32142 18194 32158
rect 18228 32142 18280 32176
rect 18314 32142 18366 32176
rect 18400 32142 18407 32176
rect 18015 32090 18018 32142
rect 18070 32104 18128 32142
rect 18180 32104 18407 32142
rect 18070 32090 18108 32104
rect 18180 32090 18194 32104
tri 331 32070 337 32076 sw
rect 18015 32074 18022 32090
rect 18056 32074 18108 32090
rect 18142 32074 18194 32090
rect 203 32064 337 32070
rect 203 32030 218 32064
rect 252 32034 337 32064
tri 337 32034 373 32070 sw
rect 252 32030 373 32034
rect 203 31992 373 32030
rect 203 31985 218 31992
tri 203 31977 211 31985 ne
rect 211 31958 218 31985
rect 252 31958 373 31992
rect 211 31920 373 31958
rect 211 31886 218 31920
rect 252 31886 373 31920
rect 211 31848 373 31886
rect 211 31814 218 31848
rect 252 31814 373 31848
rect 211 31776 373 31814
rect 211 31742 218 31776
rect 252 31742 373 31776
rect 211 31704 373 31742
rect 211 31670 218 31704
rect 252 31670 373 31704
rect 211 31632 373 31670
rect 211 31598 218 31632
rect 252 31598 373 31632
rect 211 31560 373 31598
rect 211 31526 218 31560
rect 252 31526 373 31560
rect 211 31488 373 31526
rect 211 31454 218 31488
rect 252 31454 373 31488
rect 211 31416 373 31454
rect 211 31382 218 31416
rect 252 31382 373 31416
rect 211 31344 373 31382
rect 211 31310 218 31344
rect 252 31310 373 31344
rect 211 31272 373 31310
rect 211 31238 218 31272
rect 252 31238 373 31272
rect 211 31200 373 31238
rect 18015 32022 18018 32074
rect 18070 32070 18108 32074
rect 18180 32070 18194 32074
rect 18228 32070 18280 32104
rect 18314 32070 18366 32104
rect 18400 32070 18407 32104
rect 18070 32032 18128 32070
rect 18180 32032 18407 32070
rect 18070 32022 18108 32032
rect 18180 32022 18194 32032
rect 18015 31998 18022 32022
rect 18056 31998 18108 32022
rect 18142 31998 18194 32022
rect 18228 31998 18280 32032
rect 18314 31998 18366 32032
rect 18400 31998 18407 32032
rect 18015 31960 18407 31998
rect 18015 31926 18022 31960
rect 18056 31926 18108 31960
rect 18142 31926 18194 31960
rect 18228 31926 18280 31960
rect 18314 31926 18366 31960
rect 18400 31926 18407 31960
rect 18015 31888 18407 31926
rect 18015 31854 18022 31888
rect 18056 31854 18108 31888
rect 18142 31854 18194 31888
rect 18228 31854 18280 31888
rect 18314 31854 18366 31888
rect 18400 31854 18407 31888
rect 18015 31816 18407 31854
rect 18015 31782 18022 31816
rect 18056 31782 18108 31816
rect 18142 31782 18194 31816
rect 18228 31782 18280 31816
rect 18314 31782 18366 31816
rect 18400 31782 18407 31816
rect 18015 31744 18407 31782
rect 18015 31710 18022 31744
rect 18056 31710 18108 31744
rect 18142 31710 18194 31744
rect 18228 31710 18280 31744
rect 18314 31710 18366 31744
rect 18400 31710 18407 31744
rect 18015 31672 18407 31710
rect 18015 31638 18022 31672
rect 18056 31638 18108 31672
rect 18142 31638 18194 31672
rect 18228 31638 18280 31672
rect 18314 31638 18366 31672
rect 18400 31638 18407 31672
rect 18015 31600 18407 31638
rect 18015 31566 18022 31600
rect 18056 31566 18108 31600
rect 18142 31566 18194 31600
rect 18228 31566 18280 31600
rect 18314 31566 18366 31600
rect 18400 31566 18407 31600
rect 18015 31528 18407 31566
rect 18015 31494 18022 31528
rect 18056 31494 18108 31528
rect 18142 31494 18194 31528
rect 18228 31494 18280 31528
rect 18314 31494 18366 31528
rect 18400 31494 18407 31528
rect 18015 31456 18407 31494
rect 18015 31422 18022 31456
rect 18056 31422 18108 31456
rect 18142 31422 18194 31456
rect 18228 31422 18280 31456
rect 18314 31422 18366 31456
rect 18400 31422 18407 31456
rect 18015 31384 18407 31422
rect 18015 31350 18022 31384
rect 18056 31350 18108 31384
rect 18142 31350 18194 31384
rect 18228 31350 18280 31384
rect 18314 31350 18366 31384
rect 18400 31350 18407 31384
rect 18015 31312 18407 31350
rect 18015 31278 18022 31312
rect 18056 31278 18108 31312
rect 18142 31278 18194 31312
rect 18228 31278 18280 31312
rect 18314 31278 18366 31312
rect 18400 31278 18407 31312
rect 18015 31240 18407 31278
rect 18015 31206 18022 31240
rect 18056 31206 18108 31240
rect 18142 31206 18194 31240
rect 18228 31206 18280 31240
rect 18314 31206 18366 31240
rect 18400 31206 18407 31240
rect 211 31195 218 31200
rect 252 31195 373 31200
rect 211 31143 215 31195
rect 267 31143 313 31195
rect 365 31143 373 31195
rect 211 31128 373 31143
rect 211 31076 215 31128
rect 267 31076 313 31128
rect 365 31076 373 31128
rect 211 31061 373 31076
rect 211 31009 215 31061
rect 267 31009 313 31061
rect 365 31009 373 31061
rect 211 30984 373 31009
rect 959 31195 1011 31201
rect 959 31128 1011 31143
rect 959 31061 1011 31076
rect 959 31003 1011 31009
rect 18015 31168 18407 31206
rect 18015 31134 18022 31168
rect 18056 31134 18108 31168
rect 18142 31134 18194 31168
rect 18228 31134 18280 31168
rect 18314 31134 18366 31168
rect 18400 31134 18407 31168
rect 18015 31096 18407 31134
rect 18015 31062 18022 31096
rect 18056 31062 18108 31096
rect 18142 31062 18194 31096
rect 18228 31062 18280 31096
rect 18314 31062 18366 31096
rect 18400 31062 18407 31096
rect 18015 31024 18407 31062
rect 211 30950 218 30984
rect 252 30950 373 30984
rect 211 30912 373 30950
rect 211 30878 218 30912
rect 252 30878 373 30912
rect 211 30840 373 30878
rect 211 30806 218 30840
rect 252 30806 373 30840
rect 211 30768 373 30806
rect 211 30734 218 30768
rect 252 30734 373 30768
rect 211 30696 373 30734
rect 211 30662 218 30696
rect 252 30662 373 30696
rect 211 30624 373 30662
rect 211 30590 218 30624
rect 252 30590 373 30624
rect 211 30552 373 30590
rect 211 30518 218 30552
rect 252 30518 373 30552
rect 211 30480 373 30518
rect 211 30446 218 30480
rect 252 30446 373 30480
rect 211 30408 373 30446
rect 211 30374 218 30408
rect 252 30374 373 30408
rect 211 30336 373 30374
rect 211 30302 218 30336
rect 252 30302 373 30336
rect 211 30264 373 30302
rect 211 30230 218 30264
rect 252 30230 373 30264
rect 211 30192 373 30230
rect 211 30158 218 30192
rect 252 30158 373 30192
rect 211 30120 373 30158
rect 211 30086 218 30120
rect 252 30086 373 30120
rect 211 30048 373 30086
rect 211 30014 218 30048
rect 252 30014 373 30048
rect 211 29976 373 30014
rect 211 29942 218 29976
rect 252 29942 373 29976
rect 211 29904 373 29942
rect 211 29870 218 29904
rect 252 29870 373 29904
rect 211 29832 373 29870
rect 211 29798 218 29832
rect 252 29798 373 29832
rect 211 29760 373 29798
rect 211 29726 218 29760
rect 252 29726 373 29760
rect 211 29688 373 29726
rect 211 29654 218 29688
rect 252 29654 373 29688
rect 211 29616 373 29654
rect 211 29582 218 29616
rect 252 29582 373 29616
rect 211 29544 373 29582
rect 211 29510 218 29544
rect 252 29510 373 29544
rect 211 29472 373 29510
rect 211 29438 218 29472
rect 252 29438 373 29472
rect 211 29400 373 29438
rect 211 29366 218 29400
rect 252 29366 373 29400
rect 211 29328 373 29366
rect 211 29294 218 29328
rect 252 29294 373 29328
rect 211 29256 373 29294
rect 211 29222 218 29256
rect 252 29222 373 29256
rect 211 29184 373 29222
rect 211 29150 218 29184
rect 252 29150 373 29184
rect 211 29112 373 29150
rect 211 29078 218 29112
rect 252 29078 373 29112
rect 211 29040 373 29078
rect 211 29006 218 29040
rect 252 29006 373 29040
rect 211 28968 373 29006
rect 211 28934 218 28968
rect 252 28934 373 28968
rect 211 28896 373 28934
rect 211 28862 218 28896
rect 252 28862 373 28896
rect 211 28824 373 28862
rect 211 28790 218 28824
rect 252 28790 373 28824
rect 211 28752 373 28790
rect 211 28718 218 28752
rect 252 28718 373 28752
rect 211 28680 373 28718
rect 211 28646 218 28680
rect 252 28646 373 28680
rect 211 28608 373 28646
rect 211 28574 218 28608
rect 252 28574 373 28608
rect 211 28535 373 28574
rect 211 28501 218 28535
rect 252 28501 373 28535
rect 211 28462 373 28501
rect 211 28428 218 28462
rect 252 28428 373 28462
rect 211 28389 373 28428
rect 211 28355 218 28389
rect 252 28355 373 28389
rect 211 28316 373 28355
rect 211 28282 218 28316
rect 252 28282 373 28316
rect 211 28243 373 28282
rect 211 28209 218 28243
rect 252 28209 373 28243
rect 211 28170 373 28209
rect 211 28136 218 28170
rect 252 28136 373 28170
rect 211 28097 373 28136
rect 211 28063 218 28097
rect 252 28063 373 28097
rect 211 28024 373 28063
rect 211 27990 218 28024
rect 252 27990 373 28024
rect 211 27951 373 27990
rect 211 27917 218 27951
rect 252 27917 373 27951
rect 211 27878 373 27917
rect 211 27844 218 27878
rect 252 27844 373 27878
rect 211 27805 373 27844
rect 211 27771 218 27805
rect 252 27771 373 27805
rect 211 27732 373 27771
rect 211 27698 218 27732
rect 252 27698 373 27732
rect 211 27659 373 27698
rect 211 27625 218 27659
rect 252 27625 373 27659
rect 211 27586 373 27625
rect 211 27552 218 27586
rect 252 27552 373 27586
rect 211 27513 373 27552
rect 211 27479 218 27513
rect 252 27479 373 27513
rect 211 27440 373 27479
rect 211 27406 218 27440
rect 252 27406 373 27440
rect 211 27367 373 27406
rect 211 27333 218 27367
rect 252 27333 373 27367
rect 211 27294 373 27333
rect 211 27260 218 27294
rect 252 27260 373 27294
rect 211 27221 373 27260
rect 211 27187 218 27221
rect 252 27187 373 27221
rect 211 27148 373 27187
rect 211 27114 218 27148
rect 252 27114 373 27148
rect 211 27075 373 27114
rect 211 27041 218 27075
rect 252 27041 373 27075
rect 211 27002 373 27041
rect 18015 30990 18022 31024
rect 18056 30990 18108 31024
rect 18142 30990 18194 31024
rect 18228 30990 18280 31024
rect 18314 30990 18366 31024
rect 18400 30990 18407 31024
rect 18015 30952 18407 30990
rect 18015 30918 18022 30952
rect 18056 30918 18108 30952
rect 18142 30918 18194 30952
rect 18228 30918 18280 30952
rect 18314 30918 18366 30952
rect 18400 30918 18407 30952
rect 18015 30880 18407 30918
rect 18015 30846 18022 30880
rect 18056 30846 18108 30880
rect 18142 30846 18194 30880
rect 18228 30846 18280 30880
rect 18314 30846 18366 30880
rect 18400 30846 18407 30880
rect 18015 30808 18407 30846
rect 18015 30774 18022 30808
rect 18056 30774 18108 30808
rect 18142 30774 18194 30808
rect 18228 30774 18280 30808
rect 18314 30774 18366 30808
rect 18400 30774 18407 30808
rect 18015 30736 18407 30774
rect 18015 30702 18022 30736
rect 18056 30702 18108 30736
rect 18142 30702 18194 30736
rect 18228 30702 18280 30736
rect 18314 30702 18366 30736
rect 18400 30702 18407 30736
rect 18015 30664 18407 30702
rect 18015 30630 18022 30664
rect 18056 30630 18108 30664
rect 18142 30630 18194 30664
rect 18228 30630 18280 30664
rect 18314 30630 18366 30664
rect 18400 30630 18407 30664
rect 18015 30592 18407 30630
rect 18015 30558 18022 30592
rect 18056 30558 18108 30592
rect 18142 30558 18194 30592
rect 18228 30558 18280 30592
rect 18314 30558 18366 30592
rect 18400 30558 18407 30592
rect 18015 30520 18407 30558
rect 18015 30486 18022 30520
rect 18056 30486 18108 30520
rect 18142 30486 18194 30520
rect 18228 30486 18280 30520
rect 18314 30486 18366 30520
rect 18400 30486 18407 30520
rect 18015 30448 18407 30486
rect 18015 30414 18022 30448
rect 18056 30414 18108 30448
rect 18142 30414 18194 30448
rect 18228 30414 18280 30448
rect 18314 30414 18366 30448
rect 18400 30414 18407 30448
rect 18015 30376 18407 30414
rect 18015 30342 18022 30376
rect 18056 30342 18108 30376
rect 18142 30342 18194 30376
rect 18228 30342 18280 30376
rect 18314 30342 18366 30376
rect 18400 30342 18407 30376
rect 18015 30304 18407 30342
rect 18015 30270 18022 30304
rect 18056 30270 18108 30304
rect 18142 30270 18194 30304
rect 18228 30270 18280 30304
rect 18314 30270 18366 30304
rect 18400 30270 18407 30304
rect 18015 30232 18407 30270
rect 18015 30198 18022 30232
rect 18056 30198 18108 30232
rect 18142 30198 18194 30232
rect 18228 30198 18280 30232
rect 18314 30198 18366 30232
rect 18400 30198 18407 30232
rect 18015 30160 18407 30198
rect 18015 30126 18022 30160
rect 18056 30126 18108 30160
rect 18142 30126 18194 30160
rect 18228 30126 18280 30160
rect 18314 30126 18366 30160
rect 18400 30126 18407 30160
rect 18015 30088 18407 30126
rect 18015 30054 18022 30088
rect 18056 30054 18108 30088
rect 18142 30054 18194 30088
rect 18228 30054 18280 30088
rect 18314 30054 18366 30088
rect 18400 30054 18407 30088
rect 18015 30016 18407 30054
rect 18015 29982 18022 30016
rect 18056 29982 18108 30016
rect 18142 29982 18194 30016
rect 18228 29982 18280 30016
rect 18314 29982 18366 30016
rect 18400 29982 18407 30016
rect 18015 29944 18407 29982
rect 18015 29910 18022 29944
rect 18056 29910 18108 29944
rect 18142 29910 18194 29944
rect 18228 29910 18280 29944
rect 18314 29910 18366 29944
rect 18400 29910 18407 29944
rect 18015 29872 18407 29910
rect 18015 29838 18022 29872
rect 18056 29838 18108 29872
rect 18142 29838 18194 29872
rect 18228 29838 18280 29872
rect 18314 29838 18366 29872
rect 18400 29838 18407 29872
rect 18015 29800 18407 29838
rect 18015 29766 18022 29800
rect 18056 29766 18108 29800
rect 18142 29766 18194 29800
rect 18228 29766 18280 29800
rect 18314 29766 18366 29800
rect 18400 29766 18407 29800
rect 18015 29728 18407 29766
rect 18015 29694 18022 29728
rect 18056 29694 18108 29728
rect 18142 29694 18194 29728
rect 18228 29694 18280 29728
rect 18314 29694 18366 29728
rect 18400 29694 18407 29728
rect 18015 29656 18407 29694
rect 18015 29622 18022 29656
rect 18056 29622 18108 29656
rect 18142 29622 18194 29656
rect 18228 29622 18280 29656
rect 18314 29622 18366 29656
rect 18400 29622 18407 29656
rect 18015 29584 18407 29622
rect 18015 29550 18022 29584
rect 18056 29550 18108 29584
rect 18142 29550 18194 29584
rect 18228 29550 18280 29584
rect 18314 29550 18366 29584
rect 18400 29550 18407 29584
rect 18015 29512 18407 29550
rect 18015 29478 18022 29512
rect 18056 29478 18108 29512
rect 18142 29478 18194 29512
rect 18228 29478 18280 29512
rect 18314 29478 18366 29512
rect 18400 29478 18407 29512
rect 18015 29440 18407 29478
rect 18015 29406 18022 29440
rect 18056 29406 18108 29440
rect 18142 29406 18194 29440
rect 18228 29406 18280 29440
rect 18314 29406 18366 29440
rect 18400 29406 18407 29440
rect 18015 29368 18407 29406
rect 18015 29334 18022 29368
rect 18056 29334 18108 29368
rect 18142 29334 18194 29368
rect 18228 29334 18280 29368
rect 18314 29334 18366 29368
rect 18400 29334 18407 29368
rect 18015 29296 18407 29334
rect 18015 29262 18022 29296
rect 18056 29262 18108 29296
rect 18142 29262 18194 29296
rect 18228 29262 18280 29296
rect 18314 29262 18366 29296
rect 18400 29262 18407 29296
rect 18015 29224 18407 29262
rect 18015 29190 18022 29224
rect 18056 29190 18108 29224
rect 18142 29190 18194 29224
rect 18228 29190 18280 29224
rect 18314 29190 18366 29224
rect 18400 29190 18407 29224
rect 18015 29152 18407 29190
rect 18015 29118 18022 29152
rect 18056 29118 18108 29152
rect 18142 29118 18194 29152
rect 18228 29118 18280 29152
rect 18314 29118 18366 29152
rect 18400 29118 18407 29152
rect 18015 29080 18407 29118
rect 18015 29046 18022 29080
rect 18056 29046 18108 29080
rect 18142 29046 18194 29080
rect 18228 29046 18280 29080
rect 18314 29046 18366 29080
rect 18400 29046 18407 29080
rect 18015 29008 18407 29046
rect 18015 28974 18022 29008
rect 18056 28974 18108 29008
rect 18142 28974 18194 29008
rect 18228 28974 18280 29008
rect 18314 28974 18366 29008
rect 18400 28974 18407 29008
rect 18015 28936 18407 28974
rect 18015 28902 18022 28936
rect 18056 28902 18108 28936
rect 18142 28902 18194 28936
rect 18228 28902 18280 28936
rect 18314 28902 18366 28936
rect 18400 28902 18407 28936
rect 18015 28864 18407 28902
rect 18015 28830 18022 28864
rect 18056 28830 18108 28864
rect 18142 28830 18194 28864
rect 18228 28830 18280 28864
rect 18314 28830 18366 28864
rect 18400 28830 18407 28864
rect 18015 28792 18407 28830
rect 18015 28758 18022 28792
rect 18056 28758 18108 28792
rect 18142 28758 18194 28792
rect 18228 28758 18280 28792
rect 18314 28758 18366 28792
rect 18400 28758 18407 28792
rect 18015 28720 18407 28758
rect 18015 28686 18022 28720
rect 18056 28686 18108 28720
rect 18142 28686 18194 28720
rect 18228 28686 18280 28720
rect 18314 28686 18366 28720
rect 18400 28686 18407 28720
rect 18015 28648 18407 28686
rect 18015 28614 18022 28648
rect 18056 28614 18108 28648
rect 18142 28614 18194 28648
rect 18228 28614 18280 28648
rect 18314 28614 18366 28648
rect 18400 28614 18407 28648
rect 18015 28576 18407 28614
rect 18015 28542 18022 28576
rect 18056 28542 18108 28576
rect 18142 28542 18194 28576
rect 18228 28542 18280 28576
rect 18314 28542 18366 28576
rect 18400 28542 18407 28576
rect 18015 28504 18407 28542
rect 18015 28470 18022 28504
rect 18056 28470 18108 28504
rect 18142 28470 18194 28504
rect 18228 28470 18280 28504
rect 18314 28470 18366 28504
rect 18400 28470 18407 28504
rect 18015 28432 18407 28470
rect 18015 28398 18022 28432
rect 18056 28398 18108 28432
rect 18142 28398 18194 28432
rect 18228 28398 18280 28432
rect 18314 28398 18366 28432
rect 18400 28398 18407 28432
rect 18015 28360 18407 28398
rect 18015 28326 18022 28360
rect 18056 28326 18108 28360
rect 18142 28326 18194 28360
rect 18228 28326 18280 28360
rect 18314 28326 18366 28360
rect 18400 28326 18407 28360
rect 18015 28288 18407 28326
rect 18015 28254 18022 28288
rect 18056 28254 18108 28288
rect 18142 28254 18194 28288
rect 18228 28254 18280 28288
rect 18314 28254 18366 28288
rect 18400 28254 18407 28288
rect 18015 28216 18407 28254
rect 18015 28182 18022 28216
rect 18056 28182 18108 28216
rect 18142 28182 18194 28216
rect 18228 28182 18280 28216
rect 18314 28182 18366 28216
rect 18400 28182 18407 28216
rect 18015 28144 18407 28182
rect 18015 28110 18022 28144
rect 18056 28110 18108 28144
rect 18142 28110 18194 28144
rect 18228 28110 18280 28144
rect 18314 28110 18366 28144
rect 18400 28110 18407 28144
rect 18015 28072 18407 28110
rect 18015 28038 18022 28072
rect 18056 28038 18108 28072
rect 18142 28038 18194 28072
rect 18228 28038 18280 28072
rect 18314 28038 18366 28072
rect 18400 28038 18407 28072
rect 18015 28000 18407 28038
rect 18015 27966 18022 28000
rect 18056 27966 18108 28000
rect 18142 27966 18194 28000
rect 18228 27966 18280 28000
rect 18314 27966 18366 28000
rect 18400 27966 18407 28000
rect 18015 27928 18407 27966
rect 18015 27894 18022 27928
rect 18056 27894 18108 27928
rect 18142 27894 18194 27928
rect 18228 27894 18280 27928
rect 18314 27894 18366 27928
rect 18400 27894 18407 27928
rect 18015 27856 18407 27894
rect 18015 27822 18022 27856
rect 18056 27822 18108 27856
rect 18142 27822 18194 27856
rect 18228 27822 18280 27856
rect 18314 27822 18366 27856
rect 18400 27822 18407 27856
rect 18015 27784 18407 27822
rect 18015 27750 18022 27784
rect 18056 27750 18108 27784
rect 18142 27750 18194 27784
rect 18228 27750 18280 27784
rect 18314 27750 18366 27784
rect 18400 27750 18407 27784
rect 18015 27712 18407 27750
rect 18015 27678 18022 27712
rect 18056 27678 18108 27712
rect 18142 27678 18194 27712
rect 18228 27678 18280 27712
rect 18314 27678 18366 27712
rect 18400 27678 18407 27712
rect 18015 27640 18407 27678
rect 18015 27606 18022 27640
rect 18056 27606 18108 27640
rect 18142 27606 18194 27640
rect 18228 27606 18280 27640
rect 18314 27606 18366 27640
rect 18400 27606 18407 27640
rect 18015 27568 18407 27606
rect 18015 27534 18022 27568
rect 18056 27534 18108 27568
rect 18142 27534 18194 27568
rect 18228 27534 18280 27568
rect 18314 27534 18366 27568
rect 18400 27534 18407 27568
rect 18015 27496 18407 27534
rect 18015 27462 18022 27496
rect 18056 27462 18108 27496
rect 18142 27462 18194 27496
rect 18228 27462 18280 27496
rect 18314 27462 18366 27496
rect 18400 27462 18407 27496
rect 18015 27424 18407 27462
rect 18015 27390 18022 27424
rect 18056 27390 18108 27424
rect 18142 27390 18194 27424
rect 18228 27390 18280 27424
rect 18314 27390 18366 27424
rect 18400 27390 18407 27424
rect 18015 27352 18407 27390
rect 18015 27318 18022 27352
rect 18056 27318 18108 27352
rect 18142 27318 18194 27352
rect 18228 27318 18280 27352
rect 18314 27318 18366 27352
rect 18400 27318 18407 27352
rect 18015 27280 18407 27318
rect 18015 27246 18022 27280
rect 18056 27246 18108 27280
rect 18142 27246 18194 27280
rect 18228 27246 18280 27280
rect 18314 27246 18366 27280
rect 18400 27246 18407 27280
rect 18015 27208 18407 27246
rect 18015 27174 18022 27208
rect 18056 27174 18108 27208
rect 18142 27174 18194 27208
rect 18228 27174 18280 27208
rect 18314 27174 18366 27208
rect 18400 27174 18407 27208
rect 18015 27136 18407 27174
rect 18015 27102 18022 27136
rect 18056 27102 18108 27136
rect 18142 27102 18194 27136
rect 18228 27102 18280 27136
rect 18314 27102 18366 27136
rect 18400 27102 18407 27136
rect 18015 27064 18407 27102
rect 18015 27030 18022 27064
rect 18056 27030 18108 27064
rect 18142 27030 18194 27064
rect 18228 27030 18280 27064
rect 18314 27030 18366 27064
rect 18400 27030 18407 27064
rect 211 26968 218 27002
rect 252 26968 373 27002
rect 211 26929 373 26968
rect 211 26895 218 26929
rect 252 26895 373 26929
rect 211 26856 373 26895
rect 211 26822 218 26856
rect 252 26822 373 26856
rect 211 26783 373 26822
rect 211 26749 218 26783
rect 252 26749 373 26783
rect 211 26710 373 26749
rect 211 26676 218 26710
rect 252 26676 373 26710
rect 211 26637 373 26676
rect 211 26603 218 26637
rect 252 26603 373 26637
rect 211 26564 373 26603
rect 211 26530 218 26564
rect 252 26530 373 26564
rect 211 26491 373 26530
rect 211 26457 218 26491
rect 252 26457 373 26491
rect 211 26418 373 26457
rect 211 26384 218 26418
rect 252 26384 373 26418
rect 211 26345 373 26384
rect 211 26311 218 26345
rect 252 26311 373 26345
rect 211 26272 373 26311
rect 211 26238 218 26272
rect 252 26238 373 26272
rect 211 26199 373 26238
rect 211 26165 218 26199
rect 252 26165 373 26199
rect 211 26126 373 26165
rect 211 26092 218 26126
rect 252 26092 373 26126
rect 211 26053 373 26092
rect 211 26019 218 26053
rect 252 26019 373 26053
rect 211 25980 373 26019
rect 211 25946 218 25980
rect 252 25946 373 25980
rect 211 25907 373 25946
rect 211 25873 218 25907
rect 252 25873 373 25907
rect 211 25834 373 25873
rect 211 25800 218 25834
rect 252 25800 373 25834
rect 211 25761 373 25800
rect 211 25727 218 25761
rect 252 25727 373 25761
rect 211 25688 373 25727
rect 211 25654 218 25688
rect 252 25654 373 25688
rect 211 25615 373 25654
rect 211 25581 218 25615
rect 252 25581 373 25615
rect 211 25542 373 25581
rect 211 25508 218 25542
rect 252 25508 373 25542
rect 1367 27015 1734 27027
rect 1367 27006 1470 27015
rect 1367 26972 1395 27006
rect 1429 26981 1470 27006
rect 1504 26981 1544 27015
rect 1578 26981 1618 27015
rect 1652 26981 1692 27015
rect 1726 26981 1734 27015
rect 1429 26972 1734 26981
rect 1367 26943 1734 26972
rect 1367 26932 1470 26943
rect 1367 26898 1395 26932
rect 1429 26909 1470 26932
rect 1504 26909 1544 26943
rect 1578 26909 1618 26943
rect 1652 26909 1692 26943
rect 1726 26909 1734 26943
rect 1429 26898 1734 26909
rect 1367 26871 1734 26898
rect 1367 26858 1470 26871
rect 1367 26824 1395 26858
rect 1429 26837 1470 26858
rect 1504 26837 1544 26871
rect 1578 26837 1618 26871
rect 1652 26837 1692 26871
rect 1726 26837 1734 26871
rect 1429 26824 1734 26837
rect 1367 26799 1734 26824
rect 1367 26784 1470 26799
rect 1367 26750 1395 26784
rect 1429 26765 1470 26784
rect 1504 26765 1544 26799
rect 1578 26765 1618 26799
rect 1652 26765 1692 26799
rect 1726 26765 1734 26799
rect 1429 26750 1734 26765
rect 1367 26727 1734 26750
rect 1367 26710 1470 26727
rect 1367 26676 1395 26710
rect 1429 26693 1470 26710
rect 1504 26693 1544 26727
rect 1578 26693 1618 26727
rect 1652 26693 1692 26727
rect 1726 26693 1734 26727
rect 1429 26676 1734 26693
rect 1367 26655 1734 26676
rect 1367 26636 1470 26655
rect 1367 26602 1395 26636
rect 1429 26621 1470 26636
rect 1504 26621 1544 26655
rect 1578 26621 1618 26655
rect 1652 26621 1692 26655
rect 1726 26621 1734 26655
rect 1429 26602 1734 26621
rect 1367 26583 1734 26602
rect 1367 26562 1470 26583
rect 1367 26528 1395 26562
rect 1429 26549 1470 26562
rect 1504 26549 1544 26583
rect 1578 26549 1618 26583
rect 1652 26549 1692 26583
rect 1726 26549 1734 26583
rect 1429 26528 1734 26549
rect 1367 26511 1734 26528
rect 1367 26488 1470 26511
rect 1367 26454 1395 26488
rect 1429 26477 1470 26488
rect 1504 26477 1544 26511
rect 1578 26477 1618 26511
rect 1652 26477 1692 26511
rect 1726 26477 1734 26511
rect 1429 26454 1734 26477
rect 1367 26439 1734 26454
rect 1367 26414 1470 26439
rect 1367 26380 1395 26414
rect 1429 26405 1470 26414
rect 1504 26405 1544 26439
rect 1578 26405 1618 26439
rect 1652 26405 1692 26439
rect 1726 26405 1734 26439
rect 1429 26380 1734 26405
rect 1367 26367 1734 26380
rect 1367 26340 1470 26367
rect 1367 26306 1395 26340
rect 1429 26333 1470 26340
rect 1504 26333 1544 26367
rect 1578 26333 1618 26367
rect 1652 26333 1692 26367
rect 1726 26333 1734 26367
rect 1429 26306 1734 26333
rect 1367 26295 1734 26306
rect 1367 26266 1470 26295
rect 1367 26232 1395 26266
rect 1429 26261 1470 26266
rect 1504 26261 1544 26295
rect 1578 26261 1618 26295
rect 1652 26261 1692 26295
rect 1726 26261 1734 26295
rect 1429 26232 1734 26261
rect 1367 26223 1734 26232
rect 1367 26193 1470 26223
rect 1367 26159 1395 26193
rect 1429 26189 1470 26193
rect 1504 26189 1544 26223
rect 1578 26189 1618 26223
rect 1652 26189 1692 26223
rect 1726 26189 1734 26223
rect 1429 26159 1734 26189
rect 1367 26151 1734 26159
rect 1367 26120 1470 26151
rect 1367 26086 1395 26120
rect 1429 26117 1470 26120
rect 1504 26117 1544 26151
rect 1578 26117 1618 26151
rect 1652 26117 1692 26151
rect 1726 26117 1734 26151
rect 1429 26086 1734 26117
rect 1367 26079 1734 26086
rect 1367 26047 1470 26079
rect 1367 26013 1395 26047
rect 1429 26045 1470 26047
rect 1504 26045 1544 26079
rect 1578 26045 1618 26079
rect 1652 26045 1692 26079
rect 1726 26045 1734 26079
rect 1429 26013 1734 26045
rect 1367 26007 1734 26013
rect 1367 25974 1470 26007
rect 1367 25940 1395 25974
rect 1429 25973 1470 25974
rect 1504 25973 1544 26007
rect 1578 25973 1618 26007
rect 1652 25973 1692 26007
rect 1726 25973 1734 26007
rect 1429 25940 1734 25973
rect 1367 25935 1734 25940
rect 1367 25901 1470 25935
rect 1504 25901 1544 25935
rect 1578 25901 1618 25935
rect 1652 25901 1692 25935
rect 1726 25901 1734 25935
rect 1367 25867 1395 25901
rect 1429 25867 1734 25901
rect 1367 25863 1734 25867
rect 1367 25829 1470 25863
rect 1504 25829 1544 25863
rect 1578 25829 1618 25863
rect 1652 25829 1692 25863
rect 1726 25829 1734 25863
rect 1367 25828 1734 25829
rect 1367 25794 1395 25828
rect 1429 25794 1734 25828
rect 1367 25791 1734 25794
rect 1367 25757 1470 25791
rect 1504 25757 1544 25791
rect 1578 25757 1618 25791
rect 1652 25757 1692 25791
rect 1726 25757 1734 25791
rect 1367 25755 1734 25757
rect 1367 25721 1395 25755
rect 1429 25721 1734 25755
rect 1367 25719 1734 25721
rect 1367 25685 1470 25719
rect 1504 25685 1544 25719
rect 1578 25685 1618 25719
rect 1652 25685 1692 25719
rect 1726 25685 1734 25719
rect 1367 25682 1734 25685
rect 1367 25648 1395 25682
rect 1429 25648 1734 25682
rect 1367 25647 1734 25648
rect 1367 25613 1470 25647
rect 1504 25613 1544 25647
rect 1578 25613 1618 25647
rect 1652 25613 1692 25647
rect 1726 25613 1734 25647
rect 1367 25609 1734 25613
rect 1367 25575 1395 25609
rect 1429 25575 1734 25609
rect 1367 25563 1470 25575
tri 1367 25541 1389 25563 ne
rect 1389 25541 1470 25563
rect 1504 25541 1544 25575
rect 1578 25541 1618 25575
rect 1652 25541 1692 25575
rect 1726 25541 1734 25575
tri 1389 25518 1412 25541 ne
rect 1412 25518 1734 25541
tri 1412 25517 1413 25518 ne
rect 1413 25517 1734 25518
rect 211 25469 373 25508
tri 1413 25502 1428 25517 ne
rect 1428 25502 1734 25517
rect 211 25435 218 25469
rect 252 25435 373 25469
tri 1428 25468 1462 25502 ne
rect 1462 25468 1470 25502
rect 1504 25468 1544 25502
rect 1578 25468 1618 25502
rect 1652 25468 1692 25502
rect 1726 25468 1734 25502
rect 211 25396 373 25435
rect 211 25362 218 25396
rect 252 25362 373 25396
rect 211 25323 373 25362
rect 211 25289 218 25323
rect 252 25289 373 25323
rect 1462 25429 1734 25468
rect 1462 25395 1470 25429
rect 1504 25395 1544 25429
rect 1578 25395 1618 25429
rect 1652 25395 1692 25429
rect 1726 25395 1734 25429
rect 1462 25356 1734 25395
rect 1462 25322 1470 25356
rect 1504 25322 1544 25356
rect 1578 25322 1618 25356
rect 1652 25322 1692 25356
rect 1726 25322 1734 25356
tri 1460 25310 1462 25312 se
rect 1462 25310 1734 25322
rect 18015 26992 18407 27030
rect 18015 26958 18022 26992
rect 18056 26958 18108 26992
rect 18142 26958 18194 26992
rect 18228 26958 18280 26992
rect 18314 26958 18366 26992
rect 18400 26958 18407 26992
rect 18015 26920 18407 26958
rect 18015 26886 18022 26920
rect 18056 26886 18108 26920
rect 18142 26886 18194 26920
rect 18228 26886 18280 26920
rect 18314 26886 18366 26920
rect 18400 26886 18407 26920
rect 18015 26848 18407 26886
rect 18015 26814 18022 26848
rect 18056 26814 18108 26848
rect 18142 26814 18194 26848
rect 18228 26814 18280 26848
rect 18314 26814 18366 26848
rect 18400 26814 18407 26848
rect 18015 26776 18407 26814
rect 18015 26742 18022 26776
rect 18056 26742 18108 26776
rect 18142 26742 18194 26776
rect 18228 26742 18280 26776
rect 18314 26742 18366 26776
rect 18400 26742 18407 26776
rect 18015 26704 18407 26742
rect 18015 26670 18022 26704
rect 18056 26670 18108 26704
rect 18142 26670 18194 26704
rect 18228 26670 18280 26704
rect 18314 26670 18366 26704
rect 18400 26670 18407 26704
rect 18015 26632 18407 26670
rect 18015 26598 18022 26632
rect 18056 26598 18108 26632
rect 18142 26598 18194 26632
rect 18228 26598 18280 26632
rect 18314 26598 18366 26632
rect 18400 26598 18407 26632
rect 18015 26560 18407 26598
rect 18015 26526 18022 26560
rect 18056 26526 18108 26560
rect 18142 26526 18194 26560
rect 18228 26526 18280 26560
rect 18314 26526 18366 26560
rect 18400 26526 18407 26560
rect 18015 26488 18407 26526
rect 18015 26454 18022 26488
rect 18056 26454 18108 26488
rect 18142 26454 18194 26488
rect 18228 26454 18280 26488
rect 18314 26454 18366 26488
rect 18400 26454 18407 26488
rect 18015 26416 18407 26454
rect 18015 26382 18022 26416
rect 18056 26382 18108 26416
rect 18142 26382 18194 26416
rect 18228 26382 18280 26416
rect 18314 26382 18366 26416
rect 18400 26382 18407 26416
rect 18015 26344 18407 26382
rect 18015 26310 18022 26344
rect 18056 26310 18108 26344
rect 18142 26310 18194 26344
rect 18228 26310 18280 26344
rect 18314 26310 18366 26344
rect 18400 26310 18407 26344
rect 18015 26272 18407 26310
rect 18015 26238 18022 26272
rect 18056 26238 18108 26272
rect 18142 26238 18194 26272
rect 18228 26238 18280 26272
rect 18314 26238 18366 26272
rect 18400 26238 18407 26272
rect 18015 26200 18407 26238
rect 18015 26166 18022 26200
rect 18056 26166 18108 26200
rect 18142 26166 18194 26200
rect 18228 26166 18280 26200
rect 18314 26166 18366 26200
rect 18400 26166 18407 26200
rect 18015 26128 18407 26166
rect 18015 26094 18022 26128
rect 18056 26094 18108 26128
rect 18142 26094 18194 26128
rect 18228 26094 18280 26128
rect 18314 26094 18366 26128
rect 18400 26094 18407 26128
rect 18015 26056 18407 26094
rect 18015 26022 18022 26056
rect 18056 26022 18108 26056
rect 18142 26022 18194 26056
rect 18228 26022 18280 26056
rect 18314 26022 18366 26056
rect 18400 26022 18407 26056
rect 18015 25984 18407 26022
rect 18015 25950 18022 25984
rect 18056 25950 18108 25984
rect 18142 25950 18194 25984
rect 18228 25950 18280 25984
rect 18314 25950 18366 25984
rect 18400 25950 18407 25984
rect 18015 25912 18407 25950
rect 18015 25878 18022 25912
rect 18056 25878 18108 25912
rect 18142 25878 18194 25912
rect 18228 25878 18280 25912
rect 18314 25878 18366 25912
rect 18400 25878 18407 25912
rect 18015 25840 18407 25878
rect 18015 25806 18022 25840
rect 18056 25806 18108 25840
rect 18142 25806 18194 25840
rect 18228 25806 18280 25840
rect 18314 25806 18366 25840
rect 18400 25806 18407 25840
rect 18015 25768 18407 25806
rect 18015 25734 18022 25768
rect 18056 25734 18108 25768
rect 18142 25734 18194 25768
rect 18228 25734 18280 25768
rect 18314 25734 18366 25768
rect 18400 25734 18407 25768
rect 18015 25696 18407 25734
rect 18015 25662 18022 25696
rect 18056 25662 18108 25696
rect 18142 25662 18194 25696
rect 18228 25662 18280 25696
rect 18314 25662 18366 25696
rect 18400 25662 18407 25696
rect 18015 25624 18407 25662
rect 18015 25590 18022 25624
rect 18056 25590 18108 25624
rect 18142 25590 18194 25624
rect 18228 25590 18280 25624
rect 18314 25590 18366 25624
rect 18400 25590 18407 25624
rect 18015 25552 18407 25590
rect 18015 25518 18022 25552
rect 18056 25518 18108 25552
rect 18142 25518 18194 25552
rect 18228 25518 18280 25552
rect 18314 25518 18366 25552
rect 18400 25518 18407 25552
rect 18015 25480 18407 25518
rect 18015 25446 18022 25480
rect 18056 25446 18108 25480
rect 18142 25446 18194 25480
rect 18228 25446 18280 25480
rect 18314 25446 18366 25480
rect 18400 25446 18407 25480
rect 18015 25408 18407 25446
rect 18015 25374 18022 25408
rect 18056 25374 18108 25408
rect 18142 25374 18194 25408
rect 18228 25374 18280 25408
rect 18314 25374 18366 25408
rect 18400 25374 18407 25408
rect 18015 25336 18407 25374
tri 1452 25302 1460 25310 se
rect 1460 25302 1728 25310
tri 1450 25300 1452 25302 se
rect 1452 25300 1728 25302
rect 211 25250 373 25289
tri 1416 25266 1450 25300 se
rect 1450 25266 1728 25300
tri 1414 25264 1416 25266 se
rect 1416 25264 1728 25266
rect 211 25216 218 25250
rect 252 25216 373 25250
tri 1391 25241 1414 25264 se
rect 1414 25241 1728 25264
rect 211 25177 373 25216
rect 211 25143 218 25177
rect 252 25143 373 25177
rect 211 25104 373 25143
rect 211 25070 218 25104
rect 252 25070 373 25104
rect 211 25031 373 25070
rect 211 24997 218 25031
rect 252 24997 373 25031
rect 211 24958 373 24997
rect 211 24924 218 24958
rect 252 24924 373 24958
rect 211 24885 373 24924
rect 211 24851 218 24885
rect 252 24851 373 24885
rect 211 24812 373 24851
rect 211 24778 218 24812
rect 252 24778 373 24812
rect 211 24739 373 24778
rect 211 24705 218 24739
rect 252 24705 373 24739
rect 211 24666 373 24705
rect 211 24632 218 24666
rect 252 24632 373 24666
rect 211 24593 373 24632
rect 211 24559 218 24593
rect 252 24559 373 24593
rect 211 24520 373 24559
rect 211 24486 218 24520
rect 252 24486 373 24520
rect 211 24447 373 24486
rect 211 24413 218 24447
rect 252 24413 373 24447
rect 211 24374 373 24413
rect 211 24340 218 24374
rect 252 24340 373 24374
rect 211 24301 373 24340
rect 211 24267 218 24301
rect 252 24267 373 24301
rect 211 24228 373 24267
rect 211 24194 218 24228
rect 252 24194 373 24228
rect 211 24155 373 24194
rect 211 24121 218 24155
rect 252 24121 373 24155
rect 211 24082 373 24121
rect 211 24048 218 24082
rect 252 24048 373 24082
rect 211 24009 373 24048
rect 211 23975 218 24009
rect 252 23975 373 24009
rect 211 23936 373 23975
rect 211 23902 218 23936
rect 252 23902 373 23936
rect 211 23863 373 23902
rect 211 23829 218 23863
rect 252 23831 373 23863
rect 1005 25209 1728 25241
rect 1005 25175 1059 25209
rect 1093 25175 1133 25209
rect 1167 25175 1207 25209
rect 1241 25175 1281 25209
rect 1315 25175 1355 25209
rect 1389 25175 1429 25209
rect 1463 25175 1503 25209
rect 1537 25175 1577 25209
rect 1611 25175 1651 25209
rect 1685 25175 1728 25209
rect 1005 25134 1728 25175
rect 1005 25100 1059 25134
rect 1093 25100 1133 25134
rect 1167 25100 1207 25134
rect 1241 25100 1281 25134
rect 1315 25100 1355 25134
rect 1389 25100 1429 25134
rect 1463 25100 1503 25134
rect 1537 25100 1577 25134
rect 1611 25100 1651 25134
rect 1685 25100 1728 25134
rect 1005 25059 1728 25100
rect 1005 25025 1059 25059
rect 1093 25025 1133 25059
rect 1167 25025 1207 25059
rect 1241 25025 1281 25059
rect 1315 25025 1355 25059
rect 1389 25025 1429 25059
rect 1463 25025 1503 25059
rect 1537 25025 1577 25059
rect 1611 25025 1651 25059
rect 1685 25025 1728 25059
rect 1005 24984 1728 25025
rect 1005 24950 1059 24984
rect 1093 24950 1133 24984
rect 1167 24950 1207 24984
rect 1241 24950 1281 24984
rect 1315 24950 1355 24984
rect 1389 24950 1429 24984
rect 1463 24950 1503 24984
rect 1537 24950 1577 24984
rect 1611 24950 1651 24984
rect 1685 24950 1728 24984
rect 1005 24909 1728 24950
rect 1005 24875 1059 24909
rect 1093 24875 1133 24909
rect 1167 24875 1207 24909
rect 1241 24875 1281 24909
rect 1315 24875 1355 24909
rect 1389 24875 1429 24909
rect 1463 24875 1503 24909
rect 1537 24875 1577 24909
rect 1611 24875 1651 24909
rect 1685 24875 1728 24909
rect 1005 24834 1728 24875
rect 1005 24800 1059 24834
rect 1093 24800 1133 24834
rect 1167 24800 1207 24834
rect 1241 24800 1281 24834
rect 1315 24800 1355 24834
rect 1389 24800 1429 24834
rect 1463 24800 1503 24834
rect 1537 24800 1577 24834
rect 1611 24800 1651 24834
rect 1685 24800 1728 24834
rect 1005 24759 1728 24800
rect 1005 24725 1059 24759
rect 1093 24725 1133 24759
rect 1167 24725 1207 24759
rect 1241 24725 1281 24759
rect 1315 24725 1355 24759
rect 1389 24725 1429 24759
rect 1463 24725 1503 24759
rect 1537 24725 1577 24759
rect 1611 24725 1651 24759
rect 1685 24725 1728 24759
rect 1005 24684 1728 24725
rect 1005 24650 1059 24684
rect 1093 24650 1133 24684
rect 1167 24650 1207 24684
rect 1241 24650 1281 24684
rect 1315 24650 1355 24684
rect 1389 24650 1429 24684
rect 1463 24650 1503 24684
rect 1537 24650 1577 24684
rect 1611 24650 1651 24684
rect 1685 24650 1728 24684
rect 1005 24609 1728 24650
rect 1005 24575 1059 24609
rect 1093 24575 1133 24609
rect 1167 24575 1207 24609
rect 1241 24575 1281 24609
rect 1315 24575 1355 24609
rect 1389 24575 1429 24609
rect 1463 24575 1503 24609
rect 1537 24575 1577 24609
rect 1611 24575 1651 24609
rect 1685 24575 1728 24609
rect 1005 24533 1728 24575
rect 1005 24499 1059 24533
rect 1093 24499 1133 24533
rect 1167 24499 1207 24533
rect 1241 24499 1281 24533
rect 1315 24499 1355 24533
rect 1389 24499 1429 24533
rect 1463 24499 1503 24533
rect 1537 24499 1577 24533
rect 1611 24499 1651 24533
rect 1685 24499 1728 24533
rect 1005 24457 1728 24499
rect 1005 24423 1059 24457
rect 1093 24423 1133 24457
rect 1167 24423 1207 24457
rect 1241 24423 1281 24457
rect 1315 24423 1355 24457
rect 1389 24423 1429 24457
rect 1463 24423 1503 24457
rect 1537 24423 1577 24457
rect 1611 24423 1651 24457
rect 1685 24423 1728 24457
rect 1005 24381 1728 24423
rect 1005 24347 1059 24381
rect 1093 24347 1133 24381
rect 1167 24347 1207 24381
rect 1241 24347 1281 24381
rect 1315 24347 1355 24381
rect 1389 24347 1429 24381
rect 1463 24347 1503 24381
rect 1537 24347 1577 24381
rect 1611 24347 1651 24381
rect 1685 24347 1728 24381
rect 1005 24305 1728 24347
rect 1005 24271 1059 24305
rect 1093 24271 1133 24305
rect 1167 24271 1207 24305
rect 1241 24271 1281 24305
rect 1315 24271 1355 24305
rect 1389 24271 1429 24305
rect 1463 24271 1503 24305
rect 1537 24271 1577 24305
rect 1611 24271 1651 24305
rect 1685 24271 1728 24305
rect 1005 24229 1728 24271
rect 1005 24195 1059 24229
rect 1093 24195 1133 24229
rect 1167 24195 1207 24229
rect 1241 24195 1281 24229
rect 1315 24195 1355 24229
rect 1389 24195 1429 24229
rect 1463 24195 1503 24229
rect 1537 24195 1577 24229
rect 1611 24195 1651 24229
rect 1685 24195 1728 24229
rect 1005 24153 1728 24195
rect 1005 24119 1059 24153
rect 1093 24119 1133 24153
rect 1167 24119 1207 24153
rect 1241 24119 1281 24153
rect 1315 24119 1355 24153
rect 1389 24119 1429 24153
rect 1463 24119 1503 24153
rect 1537 24119 1577 24153
rect 1611 24119 1651 24153
rect 1685 24119 1728 24153
rect 1005 24077 1728 24119
rect 1005 24043 1059 24077
rect 1093 24043 1133 24077
rect 1167 24043 1207 24077
rect 1241 24043 1281 24077
rect 1315 24043 1355 24077
rect 1389 24043 1429 24077
rect 1463 24043 1503 24077
rect 1537 24043 1577 24077
rect 1611 24043 1651 24077
rect 1685 24043 1728 24077
rect 1005 24001 1728 24043
rect 1005 23967 1059 24001
rect 1093 23967 1133 24001
rect 1167 23967 1207 24001
rect 1241 23967 1281 24001
rect 1315 23967 1355 24001
rect 1389 23967 1429 24001
rect 1463 23967 1503 24001
rect 1537 23967 1577 24001
rect 1611 23967 1651 24001
rect 1685 23967 1728 24001
rect 1005 23925 1728 23967
rect 1005 23891 1059 23925
rect 1093 23891 1133 23925
rect 1167 23891 1207 23925
rect 1241 23891 1281 23925
rect 1315 23891 1355 23925
rect 1389 23891 1429 23925
rect 1463 23891 1503 23925
rect 1537 23891 1577 23925
rect 1611 23891 1651 23925
rect 1685 23891 1728 23925
rect 1005 23849 1728 23891
rect 1005 23831 1059 23849
rect 252 23829 1059 23831
rect 211 23815 1059 23829
rect 1093 23815 1133 23849
rect 1167 23815 1207 23849
rect 1241 23815 1281 23849
rect 1315 23815 1355 23849
rect 1389 23815 1429 23849
rect 1463 23815 1503 23849
rect 1537 23815 1577 23849
rect 1611 23815 1651 23849
rect 1685 23815 1728 23849
rect 211 23783 1728 23815
rect 18015 25302 18022 25336
rect 18056 25302 18108 25336
rect 18142 25302 18194 25336
rect 18228 25302 18280 25336
rect 18314 25302 18366 25336
rect 18400 25302 18407 25336
rect 18015 25264 18407 25302
rect 18015 25230 18022 25264
rect 18056 25230 18108 25264
rect 18142 25230 18194 25264
rect 18228 25230 18280 25264
rect 18314 25230 18366 25264
rect 18400 25230 18407 25264
rect 18015 25192 18407 25230
rect 18015 25158 18022 25192
rect 18056 25158 18108 25192
rect 18142 25158 18194 25192
rect 18228 25158 18280 25192
rect 18314 25158 18366 25192
rect 18400 25158 18407 25192
rect 18015 25120 18407 25158
rect 18015 25086 18022 25120
rect 18056 25086 18108 25120
rect 18142 25086 18194 25120
rect 18228 25086 18280 25120
rect 18314 25086 18366 25120
rect 18400 25086 18407 25120
rect 18015 25048 18407 25086
rect 18015 25014 18022 25048
rect 18056 25014 18108 25048
rect 18142 25014 18194 25048
rect 18228 25014 18280 25048
rect 18314 25014 18366 25048
rect 18400 25014 18407 25048
rect 18015 24976 18407 25014
rect 18015 24942 18022 24976
rect 18056 24942 18108 24976
rect 18142 24942 18194 24976
rect 18228 24942 18280 24976
rect 18314 24942 18366 24976
rect 18400 24942 18407 24976
rect 18015 24904 18407 24942
rect 18015 24870 18022 24904
rect 18056 24870 18108 24904
rect 18142 24870 18194 24904
rect 18228 24870 18280 24904
rect 18314 24870 18366 24904
rect 18400 24870 18407 24904
rect 18015 24832 18407 24870
rect 18015 24798 18022 24832
rect 18056 24798 18108 24832
rect 18142 24798 18194 24832
rect 18228 24798 18280 24832
rect 18314 24798 18366 24832
rect 18400 24798 18407 24832
rect 18015 24760 18407 24798
rect 18015 24726 18022 24760
rect 18056 24726 18108 24760
rect 18142 24726 18194 24760
rect 18228 24726 18280 24760
rect 18314 24726 18366 24760
rect 18400 24726 18407 24760
rect 18015 24688 18407 24726
rect 18015 24654 18022 24688
rect 18056 24654 18108 24688
rect 18142 24654 18194 24688
rect 18228 24654 18280 24688
rect 18314 24654 18366 24688
rect 18400 24654 18407 24688
rect 18015 24616 18407 24654
rect 18015 24582 18022 24616
rect 18056 24582 18108 24616
rect 18142 24582 18194 24616
rect 18228 24582 18280 24616
rect 18314 24582 18366 24616
rect 18400 24582 18407 24616
rect 18015 24544 18407 24582
rect 18015 24510 18022 24544
rect 18056 24510 18108 24544
rect 18142 24510 18194 24544
rect 18228 24510 18280 24544
rect 18314 24510 18366 24544
rect 18400 24510 18407 24544
rect 18015 24472 18407 24510
rect 18015 24438 18022 24472
rect 18056 24438 18108 24472
rect 18142 24438 18194 24472
rect 18228 24438 18280 24472
rect 18314 24438 18366 24472
rect 18400 24438 18407 24472
rect 18015 24400 18407 24438
rect 18015 24366 18022 24400
rect 18056 24366 18108 24400
rect 18142 24366 18194 24400
rect 18228 24366 18280 24400
rect 18314 24366 18366 24400
rect 18400 24366 18407 24400
rect 18015 24328 18407 24366
rect 18015 24294 18022 24328
rect 18056 24294 18108 24328
rect 18142 24294 18194 24328
rect 18228 24294 18280 24328
rect 18314 24294 18366 24328
rect 18400 24294 18407 24328
rect 18015 24256 18407 24294
rect 18015 24222 18022 24256
rect 18056 24222 18108 24256
rect 18142 24222 18194 24256
rect 18228 24222 18280 24256
rect 18314 24222 18366 24256
rect 18400 24222 18407 24256
rect 18015 24184 18407 24222
rect 18015 24150 18022 24184
rect 18056 24150 18108 24184
rect 18142 24150 18194 24184
rect 18228 24150 18280 24184
rect 18314 24150 18366 24184
rect 18400 24150 18407 24184
rect 18015 24112 18407 24150
rect 18015 24078 18022 24112
rect 18056 24078 18108 24112
rect 18142 24078 18194 24112
rect 18228 24078 18280 24112
rect 18314 24078 18366 24112
rect 18400 24078 18407 24112
rect 18015 24040 18407 24078
rect 18015 24006 18022 24040
rect 18056 24006 18108 24040
rect 18142 24006 18194 24040
rect 18228 24006 18280 24040
rect 18314 24006 18366 24040
rect 18400 24006 18407 24040
rect 18015 23968 18407 24006
rect 18015 23934 18022 23968
rect 18056 23934 18108 23968
rect 18142 23934 18194 23968
rect 18228 23934 18280 23968
rect 18314 23934 18366 23968
rect 18400 23934 18407 23968
rect 18015 23896 18407 23934
rect 18015 23862 18022 23896
rect 18056 23862 18108 23896
rect 18142 23862 18194 23896
rect 18228 23862 18280 23896
rect 18314 23862 18366 23896
rect 18400 23862 18407 23896
rect 18015 23824 18407 23862
rect 18015 23790 18022 23824
rect 18056 23790 18108 23824
rect 18142 23790 18194 23824
rect 18228 23790 18280 23824
rect 18314 23790 18366 23824
rect 18400 23790 18407 23824
rect 211 23736 1646 23783
rect 205 23724 1646 23736
rect 205 23690 212 23724
rect 246 23690 288 23724
rect 322 23690 364 23724
rect 398 23690 440 23724
rect 474 23703 1646 23724
rect 474 23690 513 23703
rect 205 23669 513 23690
rect 547 23669 590 23703
rect 624 23669 667 23703
rect 701 23669 744 23703
rect 778 23669 821 23703
rect 855 23669 898 23703
rect 932 23669 975 23703
rect 1009 23669 1052 23703
rect 1086 23669 1129 23703
rect 1163 23669 1206 23703
rect 1240 23669 1283 23703
rect 1317 23669 1360 23703
rect 1394 23669 1437 23703
rect 1471 23669 1646 23703
rect 205 23652 1646 23669
rect 205 23618 212 23652
rect 246 23618 288 23652
rect 322 23618 364 23652
rect 398 23618 440 23652
rect 474 23623 1646 23652
rect 474 23618 513 23623
rect 205 23589 513 23618
rect 547 23589 590 23623
rect 624 23589 667 23623
rect 701 23589 744 23623
rect 778 23589 821 23623
rect 855 23589 898 23623
rect 932 23589 975 23623
rect 1009 23589 1052 23623
rect 1086 23589 1129 23623
rect 1163 23589 1206 23623
rect 1240 23589 1283 23623
rect 1317 23589 1360 23623
rect 1394 23589 1437 23623
rect 1471 23607 1646 23623
rect 18015 23752 18407 23790
rect 18015 23718 18022 23752
rect 18056 23718 18108 23752
rect 18142 23718 18194 23752
rect 18228 23718 18280 23752
rect 18314 23718 18366 23752
rect 18400 23718 18407 23752
rect 18015 23680 18407 23718
rect 18015 23646 18022 23680
rect 18056 23646 18108 23680
rect 18142 23646 18194 23680
rect 18228 23646 18280 23680
rect 18314 23646 18366 23680
rect 18400 23646 18407 23680
rect 18015 23607 18407 23646
rect 1471 23589 1505 23607
rect 205 23580 1505 23589
rect 205 23546 212 23580
rect 246 23546 288 23580
rect 322 23546 364 23580
rect 398 23546 440 23580
rect 474 23546 1505 23580
rect 205 23543 1505 23546
rect 205 23509 513 23543
rect 547 23509 590 23543
rect 624 23509 667 23543
rect 701 23509 744 23543
rect 778 23509 821 23543
rect 855 23509 898 23543
rect 932 23509 975 23543
rect 1009 23509 1052 23543
rect 1086 23509 1129 23543
rect 1163 23509 1206 23543
rect 1240 23509 1283 23543
rect 1317 23509 1360 23543
rect 1394 23509 1437 23543
rect 1471 23509 1505 23543
rect 205 23508 1505 23509
rect 205 23474 212 23508
rect 246 23474 288 23508
rect 322 23474 364 23508
rect 398 23474 440 23508
rect 474 23474 1505 23508
rect 18015 23573 18022 23607
rect 18056 23573 18108 23607
rect 18142 23573 18194 23607
rect 18228 23573 18280 23607
rect 18314 23573 18366 23607
rect 18400 23573 18407 23607
rect 18015 23534 18407 23573
rect 18015 23500 18022 23534
rect 18056 23500 18108 23534
rect 18142 23500 18194 23534
rect 18228 23500 18280 23534
rect 18314 23500 18366 23534
rect 18400 23500 18407 23534
rect 18015 23488 18407 23500
rect 22823 33312 22829 33346
rect 22863 33312 22911 33346
rect 22945 33312 22993 33346
rect 23027 33312 23075 33346
rect 23109 33312 23157 33346
rect 23191 33312 23239 33346
rect 23273 33312 23279 33346
rect 22823 33273 23279 33312
rect 22823 33239 22829 33273
rect 22863 33239 22911 33273
rect 22945 33239 22993 33273
rect 23027 33239 23075 33273
rect 23109 33239 23157 33273
rect 23191 33239 23239 33273
rect 23273 33239 23279 33273
rect 22823 33200 23279 33239
rect 22823 33166 22829 33200
rect 22863 33166 22911 33200
rect 22945 33166 22993 33200
rect 23027 33166 23075 33200
rect 23109 33166 23157 33200
rect 23191 33166 23239 33200
rect 23273 33166 23279 33200
rect 22823 33127 23279 33166
rect 22823 33093 22829 33127
rect 22863 33093 22911 33127
rect 22945 33093 22993 33127
rect 23027 33093 23075 33127
rect 23109 33093 23157 33127
rect 23191 33093 23239 33127
rect 23273 33093 23279 33127
rect 22823 33054 23279 33093
rect 22823 33020 22829 33054
rect 22863 33020 22911 33054
rect 22945 33020 22993 33054
rect 23027 33020 23075 33054
rect 23109 33020 23157 33054
rect 23191 33020 23239 33054
rect 23273 33020 23279 33054
rect 22823 32981 23279 33020
rect 22823 32947 22829 32981
rect 22863 32947 22911 32981
rect 22945 32947 22993 32981
rect 23027 32947 23075 32981
rect 23109 32947 23157 32981
rect 23191 32947 23239 32981
rect 23273 32947 23279 32981
rect 22823 32908 23279 32947
rect 22823 32874 22829 32908
rect 22863 32874 22911 32908
rect 22945 32874 22993 32908
rect 23027 32874 23075 32908
rect 23109 32874 23157 32908
rect 23191 32874 23239 32908
rect 23273 32874 23279 32908
rect 22823 32835 23279 32874
rect 22823 32801 22829 32835
rect 22863 32801 22911 32835
rect 22945 32801 22993 32835
rect 23027 32801 23075 32835
rect 23109 32801 23157 32835
rect 23191 32801 23239 32835
rect 23273 32801 23279 32835
rect 22823 32762 23279 32801
rect 22823 32728 22829 32762
rect 22863 32728 22911 32762
rect 22945 32728 22993 32762
rect 23027 32728 23075 32762
rect 23109 32728 23157 32762
rect 23191 32728 23239 32762
rect 23273 32728 23279 32762
rect 22823 32689 23279 32728
rect 22823 32655 22829 32689
rect 22863 32655 22911 32689
rect 22945 32655 22993 32689
rect 23027 32655 23075 32689
rect 23109 32655 23157 32689
rect 23191 32655 23239 32689
rect 23273 32655 23279 32689
rect 22823 32616 23279 32655
rect 22823 32582 22829 32616
rect 22863 32582 22911 32616
rect 22945 32582 22993 32616
rect 23027 32582 23075 32616
rect 23109 32582 23157 32616
rect 23191 32582 23239 32616
rect 23273 32582 23279 32616
rect 22823 32543 23279 32582
rect 22823 32509 22829 32543
rect 22863 32509 22911 32543
rect 22945 32509 22993 32543
rect 23027 32509 23075 32543
rect 23109 32509 23157 32543
rect 23191 32509 23239 32543
rect 23273 32509 23279 32543
rect 22823 32470 23279 32509
rect 22823 32436 22829 32470
rect 22863 32436 22911 32470
rect 22945 32436 22993 32470
rect 23027 32436 23075 32470
rect 23109 32436 23157 32470
rect 23191 32436 23239 32470
rect 23273 32436 23279 32470
rect 22823 32397 23279 32436
rect 22823 32363 22829 32397
rect 22863 32363 22911 32397
rect 22945 32363 22993 32397
rect 23027 32363 23075 32397
rect 23109 32363 23157 32397
rect 23191 32363 23239 32397
rect 23273 32363 23279 32397
rect 22823 32324 23279 32363
rect 22823 32290 22829 32324
rect 22863 32290 22911 32324
rect 22945 32290 22993 32324
rect 23027 32290 23075 32324
rect 23109 32290 23157 32324
rect 23191 32290 23239 32324
rect 23273 32290 23279 32324
rect 22823 32251 23279 32290
rect 22823 32217 22829 32251
rect 22863 32217 22911 32251
rect 22945 32217 22993 32251
rect 23027 32217 23075 32251
rect 23109 32217 23157 32251
rect 23191 32217 23239 32251
rect 23273 32217 23279 32251
rect 22823 32178 23279 32217
rect 22823 32144 22829 32178
rect 22863 32144 22911 32178
rect 22945 32144 22993 32178
rect 23027 32144 23075 32178
rect 23109 32144 23157 32178
rect 23191 32144 23239 32178
rect 23273 32144 23279 32178
rect 22823 32105 23279 32144
rect 22823 32071 22829 32105
rect 22863 32071 22911 32105
rect 22945 32071 22993 32105
rect 23027 32071 23075 32105
rect 23109 32071 23157 32105
rect 23191 32071 23239 32105
rect 23273 32071 23279 32105
rect 22823 32032 23279 32071
rect 22823 31998 22829 32032
rect 22863 31998 22911 32032
rect 22945 31998 22993 32032
rect 23027 31998 23075 32032
rect 23109 31998 23157 32032
rect 23191 31998 23239 32032
rect 23273 31998 23279 32032
rect 22823 31959 23279 31998
rect 22823 31925 22829 31959
rect 22863 31925 22911 31959
rect 22945 31925 22993 31959
rect 23027 31925 23075 31959
rect 23109 31925 23157 31959
rect 23191 31925 23239 31959
rect 23273 31925 23279 31959
rect 22823 31886 23279 31925
rect 22823 31852 22829 31886
rect 22863 31852 22911 31886
rect 22945 31852 22993 31886
rect 23027 31852 23075 31886
rect 23109 31852 23157 31886
rect 23191 31852 23239 31886
rect 23273 31852 23279 31886
rect 22823 31813 23279 31852
rect 22823 31779 22829 31813
rect 22863 31779 22911 31813
rect 22945 31779 22993 31813
rect 23027 31779 23075 31813
rect 23109 31779 23157 31813
rect 23191 31779 23239 31813
rect 23273 31779 23279 31813
rect 22823 31740 23279 31779
rect 22823 31706 22829 31740
rect 22863 31706 22911 31740
rect 22945 31706 22993 31740
rect 23027 31706 23075 31740
rect 23109 31706 23157 31740
rect 23191 31706 23239 31740
rect 23273 31706 23279 31740
rect 22823 31674 23279 31706
rect 22823 31642 23075 31674
rect 22823 31608 22830 31642
rect 22864 31608 22932 31642
rect 22966 31608 23034 31642
rect 23068 31608 23075 31642
rect 22823 31568 23075 31608
rect 22823 31534 22830 31568
rect 22864 31534 22932 31568
rect 22966 31534 23034 31568
rect 23068 31534 23075 31568
rect 22823 31494 23075 31534
rect 22823 31460 22830 31494
rect 22864 31460 22932 31494
rect 22966 31460 23034 31494
rect 23068 31460 23075 31494
rect 22823 31420 23075 31460
rect 22823 31386 22830 31420
rect 22864 31386 22932 31420
rect 22966 31386 23034 31420
rect 23068 31386 23075 31420
rect 22823 31346 23075 31386
rect 22823 31312 22830 31346
rect 22864 31312 22932 31346
rect 22966 31312 23034 31346
rect 23068 31312 23075 31346
rect 22823 31271 23075 31312
rect 22823 31237 22830 31271
rect 22864 31237 22932 31271
rect 22966 31237 23034 31271
rect 23068 31237 23075 31271
rect 22823 31196 23075 31237
rect 22823 31162 22830 31196
rect 22864 31162 22932 31196
rect 22966 31162 23034 31196
rect 23068 31162 23075 31196
rect 22823 31121 23075 31162
rect 22823 31087 22830 31121
rect 22864 31087 22932 31121
rect 22966 31087 23034 31121
rect 23068 31087 23075 31121
rect 22823 31046 23075 31087
rect 22823 31012 22830 31046
rect 22864 31012 22932 31046
rect 22966 31012 23034 31046
rect 23068 31012 23075 31046
rect 22823 30971 23075 31012
rect 22823 30937 22830 30971
rect 22864 30937 22932 30971
rect 22966 30937 23034 30971
rect 23068 30937 23075 30971
rect 22823 30896 23075 30937
rect 22823 30862 22830 30896
rect 22864 30862 22932 30896
rect 22966 30862 23034 30896
rect 23068 30862 23075 30896
rect 22823 30821 23075 30862
rect 22823 30787 22830 30821
rect 22864 30787 22932 30821
rect 22966 30787 23034 30821
rect 23068 30787 23075 30821
rect 22823 30746 23075 30787
rect 22823 30712 22830 30746
rect 22864 30712 22932 30746
rect 22966 30712 23034 30746
rect 23068 30712 23075 30746
rect 22823 30671 23075 30712
rect 22823 30637 22830 30671
rect 22864 30637 22932 30671
rect 22966 30637 23034 30671
rect 23068 30637 23075 30671
rect 22823 30596 23075 30637
rect 22823 30562 22830 30596
rect 22864 30562 22932 30596
rect 22966 30562 23034 30596
rect 23068 30562 23075 30596
rect 22823 30521 23075 30562
rect 22823 30487 22830 30521
rect 22864 30487 22932 30521
rect 22966 30487 23034 30521
rect 23068 30487 23075 30521
rect 22823 30446 23075 30487
rect 22823 30412 22830 30446
rect 22864 30412 22932 30446
rect 22966 30412 23034 30446
rect 23068 30412 23075 30446
rect 22823 30371 23075 30412
rect 22823 30337 22830 30371
rect 22864 30337 22932 30371
rect 22966 30337 23034 30371
rect 23068 30337 23075 30371
rect 22823 30296 23075 30337
rect 22823 30262 22830 30296
rect 22864 30262 22932 30296
rect 22966 30262 23034 30296
rect 23068 30262 23075 30296
rect 22823 30221 23075 30262
rect 22823 30187 22830 30221
rect 22864 30187 22932 30221
rect 22966 30187 23034 30221
rect 23068 30187 23075 30221
rect 22823 30146 23075 30187
rect 22823 30112 22830 30146
rect 22864 30112 22932 30146
rect 22966 30112 23034 30146
rect 23068 30112 23075 30146
rect 22823 30071 23075 30112
rect 22823 30037 22830 30071
rect 22864 30037 22932 30071
rect 22966 30037 23034 30071
rect 23068 30037 23075 30071
rect 22823 29996 23075 30037
rect 22823 29962 22830 29996
rect 22864 29962 22932 29996
rect 22966 29962 23034 29996
rect 23068 29962 23075 29996
rect 22823 29921 23075 29962
rect 22823 29887 22830 29921
rect 22864 29887 22932 29921
rect 22966 29887 23034 29921
rect 23068 29887 23075 29921
rect 22823 29846 23075 29887
rect 22823 29812 22830 29846
rect 22864 29812 22932 29846
rect 22966 29812 23034 29846
rect 23068 29812 23075 29846
rect 22823 29771 23075 29812
rect 22823 29737 22830 29771
rect 22864 29737 22932 29771
rect 22966 29737 23034 29771
rect 23068 29737 23075 29771
rect 22823 29705 23075 29737
rect 22823 29693 22895 29705
rect 22823 29659 22842 29693
rect 22876 29659 22895 29693
rect 22823 29621 22895 29659
rect 22823 29587 22842 29621
rect 22876 29587 22895 29621
rect 22823 29549 22895 29587
rect 22823 29515 22842 29549
rect 22876 29515 22895 29549
rect 22823 29477 22895 29515
rect 22823 29443 22842 29477
rect 22876 29443 22895 29477
rect 22823 29405 22895 29443
rect 22823 29371 22842 29405
rect 22876 29371 22895 29405
rect 22823 29333 22895 29371
rect 22823 29299 22842 29333
rect 22876 29299 22895 29333
rect 22823 29261 22895 29299
rect 22823 29227 22842 29261
rect 22876 29227 22895 29261
rect 22823 29189 22895 29227
rect 22823 29155 22842 29189
rect 22876 29155 22895 29189
rect 22823 29117 22895 29155
rect 22823 29083 22842 29117
rect 22876 29083 22895 29117
rect 22823 29045 22895 29083
rect 22823 29011 22842 29045
rect 22876 29011 22895 29045
rect 22823 28973 22895 29011
rect 22823 28939 22842 28973
rect 22876 28939 22895 28973
rect 22823 28901 22895 28939
rect 22823 28867 22842 28901
rect 22876 28867 22895 28901
rect 22823 28829 22895 28867
rect 22823 28795 22842 28829
rect 22876 28795 22895 28829
rect 22823 28757 22895 28795
rect 22823 28723 22842 28757
rect 22876 28723 22895 28757
rect 22823 28685 22895 28723
rect 22823 28651 22842 28685
rect 22876 28651 22895 28685
rect 22823 28613 22895 28651
rect 22823 28579 22842 28613
rect 22876 28579 22895 28613
rect 22823 28541 22895 28579
rect 22823 28507 22842 28541
rect 22876 28507 22895 28541
rect 22823 28469 22895 28507
rect 22823 28435 22842 28469
rect 22876 28435 22895 28469
rect 22823 28397 22895 28435
rect 22823 28363 22842 28397
rect 22876 28363 22895 28397
rect 22823 28325 22895 28363
rect 22823 28291 22842 28325
rect 22876 28291 22895 28325
rect 22823 28253 22895 28291
rect 22823 28219 22842 28253
rect 22876 28219 22895 28253
rect 22823 28181 22895 28219
rect 22823 28147 22842 28181
rect 22876 28147 22895 28181
rect 22823 28109 22895 28147
rect 22823 28075 22842 28109
rect 22876 28075 22895 28109
rect 22823 28037 22895 28075
rect 22823 28003 22842 28037
rect 22876 28003 22895 28037
rect 22823 27965 22895 28003
rect 22823 27931 22842 27965
rect 22876 27931 22895 27965
rect 22823 27893 22895 27931
rect 22823 27859 22842 27893
rect 22876 27859 22895 27893
rect 22823 27821 22895 27859
rect 22823 27787 22842 27821
rect 22876 27787 22895 27821
rect 22823 27749 22895 27787
rect 22823 27715 22842 27749
rect 22876 27715 22895 27749
rect 22823 27677 22895 27715
rect 22823 27643 22842 27677
rect 22876 27643 22895 27677
rect 22823 27605 22895 27643
rect 22823 27571 22842 27605
rect 22876 27571 22895 27605
rect 22823 27533 22895 27571
rect 22823 27499 22842 27533
rect 22876 27499 22895 27533
rect 22823 27461 22895 27499
rect 22823 27427 22842 27461
rect 22876 27427 22895 27461
rect 22823 27389 22895 27427
rect 22823 27355 22842 27389
rect 22876 27355 22895 27389
rect 22823 27317 22895 27355
rect 22823 27283 22842 27317
rect 22876 27283 22895 27317
rect 22823 27245 22895 27283
rect 22823 27211 22842 27245
rect 22876 27211 22895 27245
rect 22823 27173 22895 27211
rect 22823 27139 22842 27173
rect 22876 27139 22895 27173
rect 22823 27101 22895 27139
rect 22823 27067 22842 27101
rect 22876 27067 22895 27101
rect 22823 27029 22895 27067
rect 22823 26995 22842 27029
rect 22876 26995 22895 27029
rect 22823 26957 22895 26995
rect 22823 26923 22842 26957
rect 22876 26923 22895 26957
rect 22823 26885 22895 26923
rect 22823 26851 22842 26885
rect 22876 26851 22895 26885
rect 22823 26813 22895 26851
rect 22823 26779 22842 26813
rect 22876 26779 22895 26813
rect 22823 26741 22895 26779
rect 22823 26707 22842 26741
rect 22876 26707 22895 26741
rect 22823 26669 22895 26707
rect 22823 26635 22842 26669
rect 22876 26635 22895 26669
rect 22823 26597 22895 26635
rect 22823 26563 22842 26597
rect 22876 26563 22895 26597
rect 22823 26525 22895 26563
rect 22823 26491 22842 26525
rect 22876 26491 22895 26525
rect 22823 26453 22895 26491
rect 22823 26419 22842 26453
rect 22876 26419 22895 26453
rect 22823 26381 22895 26419
rect 22823 26347 22842 26381
rect 22876 26347 22895 26381
rect 22823 26309 22895 26347
rect 22823 26275 22842 26309
rect 22876 26275 22895 26309
rect 22823 26237 22895 26275
rect 22823 26203 22842 26237
rect 22876 26203 22895 26237
rect 22823 26165 22895 26203
rect 22823 26131 22842 26165
rect 22876 26131 22895 26165
rect 22823 26093 22895 26131
rect 22823 26059 22842 26093
rect 22876 26059 22895 26093
rect 22823 26021 22895 26059
rect 22823 25987 22842 26021
rect 22876 25987 22895 26021
rect 22823 25949 22895 25987
rect 22823 25915 22842 25949
rect 22876 25915 22895 25949
rect 22823 25877 22895 25915
rect 22823 25843 22842 25877
rect 22876 25843 22895 25877
rect 22823 25805 22895 25843
rect 22823 25771 22842 25805
rect 22876 25771 22895 25805
rect 22823 25733 22895 25771
rect 22823 25699 22842 25733
rect 22876 25699 22895 25733
rect 22823 25661 22895 25699
rect 22823 25627 22842 25661
rect 22876 25627 22895 25661
rect 22823 25589 22895 25627
rect 22823 25555 22842 25589
rect 22876 25555 22895 25589
rect 22823 25517 22895 25555
rect 22823 25483 22842 25517
rect 22876 25483 22895 25517
rect 22823 25445 22895 25483
rect 22823 25411 22842 25445
rect 22876 25411 22895 25445
rect 22823 25373 22895 25411
rect 22823 25339 22842 25373
rect 22876 25339 22895 25373
rect 22823 25300 22895 25339
rect 22823 25266 22842 25300
rect 22876 25266 22895 25300
rect 22823 25227 22895 25266
rect 22823 25193 22842 25227
rect 22876 25193 22895 25227
rect 22823 25154 22895 25193
rect 22823 25120 22842 25154
rect 22876 25120 22895 25154
rect 22823 25081 22895 25120
rect 22823 25047 22842 25081
rect 22876 25047 22895 25081
rect 22823 25008 22895 25047
rect 22823 24974 22842 25008
rect 22876 24974 22895 25008
rect 22823 24935 22895 24974
rect 22823 24901 22842 24935
rect 22876 24901 22895 24935
rect 22823 24862 22895 24901
rect 22823 24828 22842 24862
rect 22876 24828 22895 24862
rect 22823 24789 22895 24828
rect 22823 24755 22842 24789
rect 22876 24755 22895 24789
rect 22823 24716 22895 24755
rect 22823 24682 22842 24716
rect 22876 24682 22895 24716
rect 22823 24643 22895 24682
rect 22823 24609 22842 24643
rect 22876 24609 22895 24643
rect 22823 24570 22895 24609
rect 22823 24536 22842 24570
rect 22876 24536 22895 24570
rect 22823 24497 22895 24536
rect 22823 24463 22842 24497
rect 22876 24463 22895 24497
rect 22823 24424 22895 24463
rect 22823 24390 22842 24424
rect 22876 24390 22895 24424
rect 22823 24351 22895 24390
rect 22823 24317 22842 24351
rect 22876 24317 22895 24351
rect 22823 24278 22895 24317
rect 22823 24244 22842 24278
rect 22876 24244 22895 24278
rect 22823 24205 22895 24244
rect 22823 24171 22842 24205
rect 22876 24171 22895 24205
rect 22823 24132 22895 24171
rect 22823 24098 22842 24132
rect 22876 24098 22895 24132
rect 22823 24059 22895 24098
rect 22823 24025 22842 24059
rect 22876 24025 22895 24059
rect 22823 23986 22895 24025
rect 22823 23952 22842 23986
rect 22876 23952 22895 23986
rect 22823 23913 22895 23952
rect 22823 23879 22842 23913
rect 22876 23879 22895 23913
rect 22823 23840 22895 23879
rect 22823 23806 22842 23840
rect 22876 23806 22895 23840
rect 22823 23767 22895 23806
rect 22823 23733 22842 23767
rect 22876 23733 22895 23767
rect 22823 23694 22895 23733
rect 22823 23660 22842 23694
rect 22876 23660 22895 23694
rect 22823 23621 22895 23660
rect 22823 23587 22842 23621
rect 22876 23587 22895 23621
rect 22823 23548 22895 23587
rect 22823 23514 22842 23548
rect 22876 23514 22895 23548
rect 205 23463 1505 23474
rect 205 23436 513 23463
rect 205 23402 212 23436
rect 246 23402 288 23436
rect 322 23402 364 23436
rect 398 23402 440 23436
rect 474 23429 513 23436
rect 547 23429 590 23463
rect 624 23429 667 23463
rect 701 23429 744 23463
rect 778 23429 821 23463
rect 855 23429 898 23463
rect 932 23429 975 23463
rect 1009 23429 1052 23463
rect 1086 23429 1129 23463
rect 1163 23429 1206 23463
rect 1240 23429 1283 23463
rect 1317 23429 1360 23463
rect 1394 23429 1437 23463
rect 1471 23429 1505 23463
rect 474 23402 1505 23429
rect 205 23383 1505 23402
rect 205 23364 513 23383
rect 205 23330 212 23364
rect 246 23330 288 23364
rect 322 23330 364 23364
rect 398 23330 440 23364
rect 474 23349 513 23364
rect 547 23349 590 23383
rect 624 23349 667 23383
rect 701 23349 744 23383
rect 778 23349 821 23383
rect 855 23349 898 23383
rect 932 23349 975 23383
rect 1009 23349 1052 23383
rect 1086 23349 1129 23383
rect 1163 23349 1206 23383
rect 1240 23349 1283 23383
rect 1317 23349 1360 23383
rect 1394 23349 1437 23383
rect 1471 23349 1505 23383
rect 474 23330 1505 23349
rect 205 23303 1505 23330
rect 205 23292 513 23303
rect 205 23258 212 23292
rect 246 23258 288 23292
rect 322 23258 364 23292
rect 398 23258 440 23292
rect 474 23269 513 23292
rect 547 23269 590 23303
rect 624 23269 667 23303
rect 701 23269 744 23303
rect 778 23269 821 23303
rect 855 23269 898 23303
rect 932 23269 975 23303
rect 1009 23269 1052 23303
rect 1086 23269 1129 23303
rect 1163 23269 1206 23303
rect 1240 23269 1283 23303
rect 1317 23269 1360 23303
rect 1394 23269 1437 23303
rect 1471 23269 1505 23303
rect 474 23258 1505 23269
rect 205 23223 1505 23258
rect 205 23220 513 23223
rect 205 23186 212 23220
rect 246 23186 288 23220
rect 322 23186 364 23220
rect 398 23186 440 23220
rect 474 23189 513 23220
rect 547 23189 590 23223
rect 624 23189 667 23223
rect 701 23189 744 23223
rect 778 23189 821 23223
rect 855 23189 898 23223
rect 932 23189 975 23223
rect 1009 23189 1052 23223
rect 1086 23189 1129 23223
rect 1163 23189 1206 23223
rect 1240 23189 1283 23223
rect 1317 23189 1360 23223
rect 1394 23189 1437 23223
rect 1471 23189 1505 23223
rect 474 23186 1505 23189
rect 205 23182 1505 23186
rect 22823 23475 22895 23514
rect 22823 23441 22842 23475
rect 22876 23441 22895 23475
rect 22823 23402 22895 23441
rect 22823 23368 22842 23402
rect 22876 23368 22895 23402
rect 22823 23329 22895 23368
rect 22823 23295 22842 23329
rect 22876 23295 22895 23329
rect 22823 23256 22895 23295
rect 22823 23241 22842 23256
rect 22876 23241 22895 23256
rect 22823 23189 22833 23241
rect 22885 23189 22895 23241
rect 22823 23183 22895 23189
rect 205 23180 1503 23182
rect 205 23148 481 23180
rect 205 23114 212 23148
rect 246 23114 288 23148
rect 322 23114 364 23148
rect 398 23114 440 23148
rect 474 23114 481 23148
rect 205 23076 481 23114
rect 205 23042 212 23076
rect 246 23042 288 23076
rect 322 23042 364 23076
rect 398 23042 440 23076
rect 474 23042 481 23076
rect 205 23004 481 23042
rect 205 22970 212 23004
rect 246 22970 288 23004
rect 322 22970 364 23004
rect 398 22970 440 23004
rect 474 22970 481 23004
rect 205 22932 481 22970
rect 205 22898 212 22932
rect 246 22898 288 22932
rect 322 22898 364 22932
rect 398 22898 440 22932
rect 474 22898 481 22932
rect 205 22860 481 22898
rect 205 22826 212 22860
rect 246 22826 288 22860
rect 322 22826 364 22860
rect 398 22826 440 22860
rect 474 22826 481 22860
rect 205 22788 481 22826
rect 205 22754 212 22788
rect 246 22754 288 22788
rect 322 22754 364 22788
rect 398 22754 440 22788
rect 474 22754 481 22788
rect 205 22715 481 22754
rect 205 22681 212 22715
rect 246 22681 288 22715
rect 322 22681 364 22715
rect 398 22681 440 22715
rect 474 22681 481 22715
rect 205 22642 481 22681
rect 205 22608 212 22642
rect 246 22608 288 22642
rect 322 22608 364 22642
rect 398 22608 440 22642
rect 474 22608 481 22642
rect 205 22569 481 22608
rect 205 22535 212 22569
rect 246 22535 288 22569
rect 322 22535 364 22569
rect 398 22535 440 22569
rect 474 22535 481 22569
rect 205 22523 481 22535
rect 22823 23176 22842 23183
rect 22876 23176 22895 23183
rect 22823 23124 22833 23176
rect 22885 23124 22895 23176
rect 22823 23111 22895 23124
rect 22823 23059 22833 23111
rect 22885 23059 22895 23111
rect 22823 23045 22895 23059
rect 22823 22993 22833 23045
rect 22885 22993 22895 23045
rect 22823 22964 22895 22993
rect 23768 23241 23948 23247
rect 23820 23189 23832 23241
rect 23884 23189 23896 23241
rect 23768 23143 23948 23189
rect 23820 23091 23832 23143
rect 23884 23091 23896 23143
rect 23768 23045 23948 23091
rect 23820 22993 23832 23045
rect 23884 22993 23896 23045
rect 23768 22987 23948 22993
rect 22823 22930 22842 22964
rect 22876 22930 22895 22964
rect 22823 22891 22895 22930
rect 22823 22857 22842 22891
rect 22876 22857 22895 22891
rect 22823 22818 22895 22857
rect 22823 22784 22842 22818
rect 22876 22784 22895 22818
rect 22823 22745 22895 22784
rect 22823 22711 22842 22745
rect 22876 22711 22895 22745
rect 22823 22672 22895 22711
rect 22823 22638 22842 22672
rect 22876 22638 22895 22672
rect 22823 22599 22895 22638
rect 22823 22565 22842 22599
rect 22876 22565 22895 22599
rect 22823 22526 22895 22565
rect 643 22482 1089 22494
rect 643 22448 649 22482
rect 683 22448 729 22482
rect 763 22448 809 22482
rect 843 22448 889 22482
rect 923 22448 969 22482
rect 1003 22448 1049 22482
rect 1083 22448 1089 22482
rect 643 22410 1089 22448
rect 643 22376 649 22410
rect 683 22376 729 22410
rect 763 22376 809 22410
rect 843 22376 889 22410
rect 923 22376 969 22410
rect 1003 22376 1049 22410
rect 1083 22376 1089 22410
rect 643 22338 1089 22376
rect 643 22304 649 22338
rect 683 22304 729 22338
rect 763 22304 809 22338
rect 843 22304 889 22338
rect 923 22304 969 22338
rect 1003 22304 1049 22338
rect 1083 22304 1089 22338
rect 643 22266 1089 22304
rect 643 22232 649 22266
rect 683 22232 729 22266
rect 763 22232 809 22266
rect 843 22232 889 22266
rect 923 22232 969 22266
rect 1003 22232 1049 22266
rect 1083 22232 1089 22266
rect 643 22194 1089 22232
rect 643 22160 649 22194
rect 683 22160 729 22194
rect 763 22160 809 22194
rect 843 22160 889 22194
rect 923 22160 969 22194
rect 1003 22160 1049 22194
rect 1083 22160 1089 22194
rect 643 22122 1089 22160
rect 643 22088 649 22122
rect 683 22088 729 22122
rect 763 22088 809 22122
rect 843 22088 889 22122
rect 923 22088 969 22122
rect 1003 22088 1049 22122
rect 1083 22088 1089 22122
rect 22823 22492 22842 22526
rect 22876 22492 22895 22526
rect 22823 22453 22895 22492
rect 22823 22419 22842 22453
rect 22876 22419 22895 22453
rect 22823 22380 22895 22419
rect 22823 22346 22842 22380
rect 22876 22346 22895 22380
rect 22823 22307 22895 22346
rect 22823 22273 22842 22307
rect 22876 22273 22895 22307
rect 22823 22234 22895 22273
rect 22823 22200 22842 22234
rect 22876 22200 22895 22234
rect 22823 22161 22895 22200
rect 22823 22127 22842 22161
rect 22876 22127 22895 22161
rect 22823 22115 22895 22127
rect 643 22050 1089 22088
rect 643 22016 649 22050
rect 683 22016 729 22050
rect 763 22016 809 22050
rect 843 22016 889 22050
rect 923 22016 969 22050
rect 1003 22016 1049 22050
rect 1083 22016 1089 22050
rect 643 21978 1089 22016
rect 643 21944 649 21978
rect 683 21944 729 21978
rect 763 21944 809 21978
rect 843 21944 889 21978
rect 923 21944 969 21978
rect 1003 21944 1049 21978
rect 1083 21944 1089 21978
rect 643 21906 1089 21944
rect 643 21872 649 21906
rect 683 21872 729 21906
rect 763 21872 809 21906
rect 843 21872 889 21906
rect 923 21872 969 21906
rect 1003 21872 1049 21906
rect 1083 21872 1089 21906
rect 643 21834 1089 21872
rect 643 21800 649 21834
rect 683 21800 729 21834
rect 763 21800 809 21834
rect 843 21800 889 21834
rect 923 21800 969 21834
rect 1003 21800 1049 21834
rect 1083 21800 1089 21834
rect 643 21762 1089 21800
rect 643 21728 649 21762
rect 683 21728 729 21762
rect 763 21728 809 21762
rect 843 21728 889 21762
rect 923 21728 969 21762
rect 1003 21728 1049 21762
rect 1083 21728 1089 21762
rect 643 21690 1089 21728
rect 643 21656 649 21690
rect 683 21656 729 21690
rect 763 21656 809 21690
rect 843 21656 889 21690
rect 923 21656 969 21690
rect 1003 21656 1049 21690
rect 1083 21656 1089 21690
rect 643 21618 1089 21656
rect 643 21584 649 21618
rect 683 21584 729 21618
rect 763 21584 809 21618
rect 843 21584 889 21618
rect 923 21584 969 21618
rect 1003 21584 1049 21618
rect 1083 21584 1089 21618
rect 643 21546 1089 21584
rect 643 21512 649 21546
rect 683 21512 729 21546
rect 763 21512 809 21546
rect 843 21512 889 21546
rect 923 21512 969 21546
rect 1003 21512 1049 21546
rect 1083 21512 1089 21546
rect 643 21474 1089 21512
rect 643 21440 649 21474
rect 683 21440 729 21474
rect 763 21440 809 21474
rect 843 21440 889 21474
rect 923 21440 969 21474
rect 1003 21440 1049 21474
rect 1083 21440 1089 21474
rect 643 21402 1089 21440
rect 643 21368 649 21402
rect 683 21368 729 21402
rect 763 21368 809 21402
rect 843 21368 889 21402
rect 923 21368 969 21402
rect 1003 21368 1049 21402
rect 1083 21368 1089 21402
rect 643 21330 1089 21368
rect 643 21296 649 21330
rect 683 21296 729 21330
rect 763 21296 809 21330
rect 843 21296 889 21330
rect 923 21296 969 21330
rect 1003 21296 1049 21330
rect 1083 21296 1089 21330
rect 643 21258 1089 21296
rect 643 21224 649 21258
rect 683 21224 729 21258
rect 763 21224 809 21258
rect 843 21224 889 21258
rect 923 21224 969 21258
rect 1003 21224 1049 21258
rect 1083 21224 1089 21258
rect 643 21186 1089 21224
rect 643 21152 649 21186
rect 683 21152 729 21186
rect 763 21152 809 21186
rect 843 21152 889 21186
rect 923 21152 969 21186
rect 1003 21152 1049 21186
rect 1083 21152 1089 21186
rect 643 21114 1089 21152
rect 643 21080 649 21114
rect 683 21080 729 21114
rect 763 21080 809 21114
rect 843 21080 889 21114
rect 923 21080 969 21114
rect 1003 21080 1049 21114
rect 1083 21080 1089 21114
rect 643 21042 1089 21080
rect 643 21008 649 21042
rect 683 21008 729 21042
rect 763 21008 809 21042
rect 843 21008 889 21042
rect 923 21008 969 21042
rect 1003 21008 1049 21042
rect 1083 21008 1089 21042
rect 643 20970 1089 21008
rect 643 20936 649 20970
rect 683 20936 729 20970
rect 763 20936 809 20970
rect 843 20936 889 20970
rect 923 20936 969 20970
rect 1003 20936 1049 20970
rect 1083 20936 1089 20970
rect 643 20898 1089 20936
rect 643 20864 649 20898
rect 683 20864 729 20898
rect 763 20864 809 20898
rect 843 20864 889 20898
rect 923 20864 969 20898
rect 1003 20864 1049 20898
rect 1083 20864 1089 20898
rect 643 20826 1089 20864
rect 643 20792 649 20826
rect 683 20792 729 20826
rect 763 20792 809 20826
rect 843 20792 889 20826
rect 923 20792 969 20826
rect 1003 20792 1049 20826
rect 1083 20792 1089 20826
rect 643 20754 1089 20792
rect 643 20720 649 20754
rect 683 20720 729 20754
rect 763 20720 809 20754
rect 843 20720 889 20754
rect 923 20720 969 20754
rect 1003 20720 1049 20754
rect 1083 20720 1089 20754
rect 643 20682 1089 20720
rect 643 20648 649 20682
rect 683 20648 729 20682
rect 763 20648 809 20682
rect 843 20648 889 20682
rect 923 20648 969 20682
rect 1003 20648 1049 20682
rect 1083 20648 1089 20682
rect 643 20610 1089 20648
rect 643 20576 649 20610
rect 683 20576 729 20610
rect 763 20576 809 20610
rect 843 20576 889 20610
rect 923 20576 969 20610
rect 1003 20576 1049 20610
rect 1083 20576 1089 20610
rect 643 20538 1089 20576
rect 643 20504 649 20538
rect 683 20504 729 20538
rect 763 20504 809 20538
rect 843 20504 889 20538
rect 923 20504 969 20538
rect 1003 20504 1049 20538
rect 1083 20504 1089 20538
rect 643 20466 1089 20504
rect 643 20432 649 20466
rect 683 20432 729 20466
rect 763 20432 809 20466
rect 843 20432 889 20466
rect 923 20432 969 20466
rect 1003 20432 1049 20466
rect 1083 20432 1089 20466
rect 643 20394 1089 20432
rect 643 20360 649 20394
rect 683 20360 729 20394
rect 763 20360 809 20394
rect 843 20360 889 20394
rect 923 20360 969 20394
rect 1003 20360 1049 20394
rect 1083 20360 1089 20394
rect 643 20322 1089 20360
tri 2345 20578 2366 20599 sw
rect 2345 20544 2366 20578
tri 2366 20544 2400 20578 sw
tri 27051 20544 27085 20578 se
rect 2345 20538 3196 20544
rect 2345 20504 2377 20538
rect 2411 20504 2453 20538
rect 2487 20504 2529 20538
rect 2563 20504 2605 20538
rect 2639 20504 2680 20538
rect 2714 20504 2755 20538
rect 2789 20504 2830 20538
rect 2864 20504 2905 20538
rect 2939 20504 2980 20538
rect 3014 20504 3055 20538
rect 3089 20504 3130 20538
rect 3164 20504 3196 20538
rect 2345 20452 3196 20504
tri 26978 20471 27051 20544 se
rect 27051 20471 27085 20544
rect 2345 20418 2377 20452
rect 2411 20418 2453 20452
rect 2487 20418 2529 20452
rect 2563 20418 2605 20452
rect 2639 20418 2680 20452
rect 2714 20418 2755 20452
rect 2789 20418 2830 20452
rect 2864 20418 2905 20452
rect 2939 20418 2980 20452
rect 3014 20418 3055 20452
rect 3089 20418 3130 20452
rect 3164 20418 3196 20452
rect 2345 20412 3196 20418
rect 26915 20439 27085 20471
rect 2345 20405 2393 20412
tri 2393 20405 2400 20412 nw
rect 26915 20405 26921 20439
rect 26955 20405 27003 20439
rect 27037 20405 27085 20439
rect 2345 20362 2350 20405
tri 2350 20362 2393 20405 nw
rect 26915 20362 27085 20405
tri 2345 20357 2350 20362 nw
rect 26915 20337 26921 20362
tri 26905 20328 26914 20337 se
rect 26914 20328 26921 20337
rect 26955 20328 27003 20362
rect 27037 20328 27085 20362
rect 643 20288 649 20322
rect 683 20288 729 20322
rect 763 20288 809 20322
rect 843 20288 889 20322
rect 923 20288 969 20322
rect 1003 20288 1049 20322
rect 1083 20288 1089 20322
rect 643 20250 1089 20288
tri 26844 20267 26905 20328 se
rect 26905 20267 27085 20328
rect 643 20216 649 20250
rect 683 20216 729 20250
rect 763 20216 809 20250
rect 843 20216 889 20250
rect 923 20216 969 20250
rect 1003 20216 1049 20250
rect 1083 20216 1089 20250
rect 643 20178 1089 20216
rect 643 20144 649 20178
rect 683 20144 729 20178
rect 763 20144 809 20178
rect 843 20144 889 20178
rect 923 20144 969 20178
rect 1003 20144 1049 20178
rect 1083 20144 1089 20178
rect 643 20106 1089 20144
rect 643 20072 649 20106
rect 683 20072 729 20106
rect 763 20072 809 20106
rect 843 20072 889 20106
rect 923 20072 969 20106
rect 1003 20072 1049 20106
rect 1083 20072 1089 20106
rect 643 20034 1089 20072
rect 26373 20260 27085 20267
rect 26373 20226 26405 20260
rect 26439 20226 26481 20260
rect 26515 20226 26557 20260
rect 26591 20226 26633 20260
rect 26667 20226 26709 20260
rect 26743 20226 26785 20260
rect 26819 20226 26861 20260
rect 26895 20226 26937 20260
rect 26971 20226 27012 20260
rect 27046 20247 27085 20260
rect 27046 20226 27083 20247
rect 26373 20176 27083 20226
rect 26373 20142 26405 20176
rect 26439 20142 26481 20176
rect 26515 20142 26557 20176
rect 26591 20142 26633 20176
rect 26667 20142 26709 20176
rect 26743 20142 26785 20176
rect 26819 20142 26861 20176
rect 26895 20142 26937 20176
rect 26971 20142 27012 20176
rect 27046 20142 27083 20176
rect 26373 20092 27083 20142
rect 26373 20058 26405 20092
rect 26439 20058 26481 20092
rect 26515 20058 26557 20092
rect 26591 20058 26633 20092
rect 26667 20058 26709 20092
rect 26743 20058 26785 20092
rect 26819 20058 26861 20092
rect 26895 20058 26937 20092
rect 26971 20058 27012 20092
rect 27046 20058 27083 20092
rect 26373 20051 27083 20058
rect 26843 20050 27083 20051
rect 643 20000 649 20034
rect 683 20000 729 20034
rect 763 20000 809 20034
rect 843 20000 889 20034
rect 923 20000 969 20034
rect 1003 20000 1049 20034
rect 1083 20000 1089 20034
rect 643 19962 1089 20000
tri 26968 19968 27050 20050 ne
rect 643 19928 649 19962
rect 683 19928 729 19962
rect 763 19928 809 19962
rect 843 19928 889 19962
rect 923 19928 969 19962
rect 1003 19928 1049 19962
rect 1083 19928 1089 19962
rect 643 19890 1089 19928
rect 643 19856 649 19890
rect 683 19856 729 19890
rect 763 19856 809 19890
rect 843 19856 889 19890
rect 923 19856 969 19890
rect 1003 19856 1049 19890
rect 1083 19856 1089 19890
rect 27050 19884 27083 20050
rect 643 19818 1089 19856
rect 643 19784 649 19818
rect 683 19784 729 19818
rect 763 19784 809 19818
rect 843 19784 889 19818
rect 923 19784 969 19818
rect 1003 19784 1049 19818
rect 1083 19784 1089 19818
rect 643 19746 1089 19784
rect 643 19712 649 19746
rect 683 19712 729 19746
rect 763 19712 809 19746
rect 843 19712 889 19746
rect 923 19712 969 19746
rect 1003 19712 1049 19746
rect 1083 19712 1089 19746
rect 643 19674 1089 19712
rect 643 19640 649 19674
rect 683 19640 729 19674
rect 763 19640 809 19674
rect 843 19640 889 19674
rect 923 19640 969 19674
rect 1003 19640 1049 19674
rect 1083 19640 1089 19674
rect 643 19602 1089 19640
rect 643 19568 649 19602
rect 683 19568 729 19602
rect 763 19568 809 19602
rect 843 19568 889 19602
rect 923 19568 969 19602
rect 1003 19568 1049 19602
rect 1083 19568 1089 19602
rect 643 19530 1089 19568
rect 643 19496 649 19530
rect 683 19496 729 19530
rect 763 19496 809 19530
rect 843 19496 889 19530
rect 923 19496 969 19530
rect 1003 19496 1049 19530
rect 1083 19496 1089 19530
rect 643 19458 1089 19496
rect 643 19424 649 19458
rect 683 19424 729 19458
rect 763 19424 809 19458
rect 843 19424 889 19458
rect 923 19424 969 19458
rect 1003 19424 1049 19458
rect 1083 19424 1089 19458
rect 643 19386 1089 19424
rect 643 19352 649 19386
rect 683 19352 729 19386
rect 763 19352 809 19386
rect 843 19352 889 19386
rect 923 19352 969 19386
rect 1003 19352 1049 19386
rect 1083 19352 1089 19386
rect 643 19314 1089 19352
rect 643 19280 649 19314
rect 683 19280 729 19314
rect 763 19280 809 19314
rect 843 19280 889 19314
rect 923 19280 969 19314
rect 1003 19280 1049 19314
rect 1083 19280 1089 19314
rect 643 19242 1089 19280
rect 643 19208 649 19242
rect 683 19208 729 19242
rect 763 19208 809 19242
rect 843 19208 889 19242
rect 923 19208 969 19242
rect 1003 19208 1049 19242
rect 1083 19208 1089 19242
rect 643 19170 1089 19208
rect 643 19136 649 19170
rect 683 19136 729 19170
rect 763 19136 809 19170
rect 843 19136 889 19170
rect 923 19136 969 19170
rect 1003 19136 1049 19170
rect 1083 19136 1089 19170
rect 643 19098 1089 19136
rect 643 19064 649 19098
rect 683 19064 729 19098
rect 763 19064 809 19098
rect 843 19064 889 19098
rect 923 19064 969 19098
rect 1003 19064 1049 19098
rect 1083 19064 1089 19098
rect 643 19026 1089 19064
rect 643 18992 649 19026
rect 683 18992 729 19026
rect 763 18992 809 19026
rect 843 18992 889 19026
rect 923 18992 969 19026
rect 1003 18992 1049 19026
rect 1083 18992 1089 19026
rect 643 18954 1089 18992
rect 643 18920 649 18954
rect 683 18920 729 18954
rect 763 18920 809 18954
rect 843 18920 889 18954
rect 923 18920 969 18954
rect 1003 18920 1049 18954
rect 1083 18920 1089 18954
rect 643 18882 1089 18920
rect 643 18848 649 18882
rect 683 18848 729 18882
rect 763 18848 809 18882
rect 843 18848 889 18882
rect 923 18848 969 18882
rect 1003 18848 1049 18882
rect 1083 18848 1089 18882
rect 643 18810 1089 18848
rect 643 18776 649 18810
rect 683 18776 729 18810
rect 763 18776 809 18810
rect 843 18776 889 18810
rect 923 18776 969 18810
rect 1003 18776 1049 18810
rect 1083 18776 1089 18810
rect 643 18738 1089 18776
rect 643 18704 649 18738
rect 683 18704 729 18738
rect 763 18704 809 18738
rect 843 18704 889 18738
rect 923 18704 969 18738
rect 1003 18704 1049 18738
rect 1083 18704 1089 18738
rect 643 18666 1089 18704
rect 643 18632 649 18666
rect 683 18632 729 18666
rect 763 18632 809 18666
rect 843 18632 889 18666
rect 923 18632 969 18666
rect 1003 18632 1049 18666
rect 1083 18632 1089 18666
rect 643 18594 1089 18632
rect 643 18560 649 18594
rect 683 18560 729 18594
rect 763 18560 809 18594
rect 843 18560 889 18594
rect 923 18560 969 18594
rect 1003 18560 1049 18594
rect 1083 18560 1089 18594
rect 643 18522 1089 18560
rect 643 18488 649 18522
rect 683 18488 729 18522
rect 763 18488 809 18522
rect 843 18488 889 18522
rect 923 18488 969 18522
rect 1003 18488 1049 18522
rect 1083 18488 1089 18522
rect 643 18450 1089 18488
rect 643 18416 649 18450
rect 683 18416 729 18450
rect 763 18416 809 18450
rect 843 18416 889 18450
rect 923 18416 969 18450
rect 1003 18416 1049 18450
rect 1083 18416 1089 18450
rect 643 18378 1089 18416
rect 643 18344 649 18378
rect 683 18344 729 18378
rect 763 18344 809 18378
rect 843 18344 889 18378
rect 923 18344 969 18378
rect 1003 18344 1049 18378
rect 1083 18344 1089 18378
rect 643 18306 1089 18344
rect 643 18272 649 18306
rect 683 18272 729 18306
rect 763 18272 809 18306
rect 843 18272 889 18306
rect 923 18272 969 18306
rect 1003 18272 1049 18306
rect 1083 18272 1089 18306
rect 643 18234 1089 18272
rect 643 18200 649 18234
rect 683 18200 729 18234
rect 763 18200 809 18234
rect 843 18200 889 18234
rect 923 18200 969 18234
rect 1003 18200 1049 18234
rect 1083 18200 1089 18234
rect 643 18162 1089 18200
rect 643 18128 649 18162
rect 683 18128 729 18162
rect 763 18128 809 18162
rect 843 18128 889 18162
rect 923 18128 969 18162
rect 1003 18128 1049 18162
rect 1083 18128 1089 18162
rect 643 18090 1089 18128
rect 643 18056 649 18090
rect 683 18056 729 18090
rect 763 18056 809 18090
rect 843 18056 889 18090
rect 923 18056 969 18090
rect 1003 18056 1049 18090
rect 1083 18056 1089 18090
rect 643 18018 1089 18056
rect 643 17984 649 18018
rect 683 17984 729 18018
rect 763 17984 809 18018
rect 843 17984 889 18018
rect 923 17984 969 18018
rect 1003 17984 1049 18018
rect 1083 17984 1089 18018
rect 643 17946 1089 17984
rect 643 17912 649 17946
rect 683 17912 729 17946
rect 763 17912 809 17946
rect 843 17912 889 17946
rect 923 17912 969 17946
rect 1003 17912 1049 17946
rect 1083 17912 1089 17946
rect 643 17874 1089 17912
rect 643 17840 649 17874
rect 683 17840 729 17874
rect 763 17840 809 17874
rect 843 17840 889 17874
rect 923 17840 969 17874
rect 1003 17840 1049 17874
rect 1083 17840 1089 17874
rect 643 17802 1089 17840
rect 643 17768 649 17802
rect 683 17768 729 17802
rect 763 17768 809 17802
rect 843 17768 889 17802
rect 923 17768 969 17802
rect 1003 17768 1049 17802
rect 1083 17768 1089 17802
rect 643 17730 1089 17768
rect 643 17696 649 17730
rect 683 17696 729 17730
rect 763 17696 809 17730
rect 843 17696 889 17730
rect 923 17696 969 17730
rect 1003 17696 1049 17730
rect 1083 17696 1089 17730
rect 643 17658 1089 17696
rect 643 17624 649 17658
rect 683 17624 729 17658
rect 763 17624 809 17658
rect 843 17624 889 17658
rect 923 17624 969 17658
rect 1003 17624 1049 17658
rect 1083 17624 1089 17658
rect 643 17586 1089 17624
rect 643 17552 649 17586
rect 683 17552 729 17586
rect 763 17552 809 17586
rect 843 17552 889 17586
rect 923 17552 969 17586
rect 1003 17552 1049 17586
rect 1083 17552 1089 17586
rect 643 17514 1089 17552
rect 643 17480 649 17514
rect 683 17480 729 17514
rect 763 17480 809 17514
rect 843 17480 889 17514
rect 923 17480 969 17514
rect 1003 17480 1049 17514
rect 1083 17480 1089 17514
rect 643 17442 1089 17480
rect 643 17408 649 17442
rect 683 17408 729 17442
rect 763 17408 809 17442
rect 843 17408 889 17442
rect 923 17408 969 17442
rect 1003 17408 1049 17442
rect 1083 17408 1089 17442
rect 643 17370 1089 17408
rect 643 17336 649 17370
rect 683 17336 729 17370
rect 763 17336 809 17370
rect 843 17336 889 17370
rect 923 17336 969 17370
rect 1003 17336 1049 17370
rect 1083 17336 1089 17370
rect 643 17298 1089 17336
rect 643 17264 649 17298
rect 683 17264 729 17298
rect 763 17264 809 17298
rect 843 17264 889 17298
rect 923 17264 969 17298
rect 1003 17264 1049 17298
rect 1083 17264 1089 17298
rect 643 17226 1089 17264
rect 643 17192 649 17226
rect 683 17192 729 17226
rect 763 17192 809 17226
rect 843 17192 889 17226
rect 923 17192 969 17226
rect 1003 17192 1049 17226
rect 1083 17192 1089 17226
rect 643 17154 1089 17192
rect 643 17120 649 17154
rect 683 17120 729 17154
rect 763 17120 809 17154
rect 843 17120 889 17154
rect 923 17120 969 17154
rect 1003 17120 1049 17154
rect 1083 17120 1089 17154
rect 643 17082 1089 17120
rect 643 17048 649 17082
rect 683 17048 729 17082
rect 763 17048 809 17082
rect 843 17048 889 17082
rect 923 17048 969 17082
rect 1003 17048 1049 17082
rect 1083 17048 1089 17082
rect 643 17010 1089 17048
rect 643 16976 649 17010
rect 683 16976 729 17010
rect 763 16976 809 17010
rect 843 16976 889 17010
rect 923 16976 969 17010
rect 1003 16976 1049 17010
rect 1083 16976 1089 17010
rect 643 16937 1089 16976
rect 643 16903 649 16937
rect 683 16903 729 16937
rect 763 16903 809 16937
rect 843 16903 889 16937
rect 923 16903 969 16937
rect 1003 16903 1049 16937
rect 1083 16903 1089 16937
rect 643 16864 1089 16903
rect 643 16830 649 16864
rect 683 16830 729 16864
rect 763 16830 809 16864
rect 843 16830 889 16864
rect 923 16830 969 16864
rect 1003 16830 1049 16864
rect 1083 16830 1089 16864
rect 643 16791 1089 16830
rect 643 16757 649 16791
rect 683 16757 729 16791
rect 763 16757 809 16791
rect 843 16757 889 16791
rect 923 16757 969 16791
rect 1003 16757 1049 16791
rect 1083 16757 1089 16791
rect 643 16718 1089 16757
rect 643 16684 649 16718
rect 683 16684 729 16718
rect 763 16684 809 16718
rect 843 16684 889 16718
rect 923 16684 969 16718
rect 1003 16684 1049 16718
rect 1083 16684 1089 16718
rect 643 16645 1089 16684
rect 643 16611 649 16645
rect 683 16611 729 16645
rect 763 16611 809 16645
rect 843 16611 889 16645
rect 923 16611 969 16645
rect 1003 16611 1049 16645
rect 1083 16611 1089 16645
rect 643 16572 1089 16611
rect 643 16538 649 16572
rect 683 16538 729 16572
rect 763 16538 809 16572
rect 843 16538 889 16572
rect 923 16538 969 16572
rect 1003 16538 1049 16572
rect 1083 16538 1089 16572
rect 643 16499 1089 16538
rect 643 16465 649 16499
rect 683 16465 729 16499
rect 763 16465 809 16499
rect 843 16465 889 16499
rect 923 16465 969 16499
rect 1003 16465 1049 16499
rect 1083 16465 1089 16499
rect 643 16426 1089 16465
rect 643 16392 649 16426
rect 683 16392 729 16426
rect 763 16392 809 16426
rect 843 16392 889 16426
rect 923 16392 969 16426
rect 1003 16392 1049 16426
rect 1083 16392 1089 16426
rect 3405 16561 3615 16596
rect 3405 16527 3417 16561
rect 3451 16527 3493 16561
rect 3527 16527 3569 16561
rect 3603 16527 3615 16561
rect 3405 16483 3615 16527
rect 3405 16449 3417 16483
rect 3451 16449 3493 16483
rect 3527 16449 3569 16483
rect 3603 16449 3615 16483
rect 3405 16425 3615 16449
rect 643 16380 1089 16392
rect 8032 16272 8278 16284
rect 8032 16238 8038 16272
rect 8072 16238 8138 16272
rect 8172 16238 8238 16272
rect 8272 16238 8278 16272
rect 8032 16189 8278 16238
rect 8032 16155 8038 16189
rect 8072 16155 8138 16189
rect 8172 16155 8238 16189
rect 8272 16155 8278 16189
rect 8032 16106 8278 16155
rect 8032 16072 8038 16106
rect 8072 16072 8138 16106
rect 8172 16072 8238 16106
rect 8272 16072 8278 16106
rect 8032 16023 8278 16072
rect 8032 15989 8038 16023
rect 8072 15989 8138 16023
rect 8172 15989 8238 16023
rect 8272 15989 8278 16023
rect 8032 15939 8278 15989
rect 8032 15905 8038 15939
rect 8072 15905 8138 15939
rect 8172 15905 8238 15939
rect 8272 15905 8278 15939
rect 8032 15855 8278 15905
rect 8032 15821 8038 15855
rect 8072 15821 8138 15855
rect 8172 15821 8238 15855
rect 8272 15821 8278 15855
rect 8032 15809 8278 15821
rect 224 12940 666 12972
rect 224 12906 235 12940
rect 269 12906 313 12940
rect 347 12906 391 12940
rect 425 12906 469 12940
rect 503 12906 547 12940
rect 581 12906 625 12940
rect 659 12906 666 12940
rect 224 12868 666 12906
rect 224 12834 235 12868
rect 269 12834 313 12868
rect 347 12834 391 12868
rect 425 12834 469 12868
rect 503 12834 547 12868
rect 581 12834 625 12868
rect 659 12834 666 12868
rect 224 12796 666 12834
rect 224 12762 235 12796
rect 269 12762 313 12796
rect 347 12762 391 12796
rect 425 12762 469 12796
rect 503 12762 547 12796
rect 581 12762 625 12796
rect 659 12762 666 12796
rect 224 12724 666 12762
rect 224 12690 235 12724
rect 269 12690 313 12724
rect 347 12690 391 12724
rect 425 12690 469 12724
rect 503 12690 547 12724
rect 581 12690 625 12724
rect 659 12690 666 12724
rect 224 12652 666 12690
rect 224 12618 235 12652
rect 269 12618 313 12652
rect 347 12618 391 12652
rect 425 12618 469 12652
rect 503 12618 547 12652
rect 581 12618 625 12652
rect 659 12618 666 12652
rect 224 12579 666 12618
rect 224 12545 235 12579
rect 269 12545 313 12579
rect 347 12545 391 12579
rect 425 12545 469 12579
rect 503 12545 547 12579
rect 581 12545 625 12579
rect 659 12545 666 12579
rect 224 12506 666 12545
rect 224 12472 235 12506
rect 269 12472 313 12506
rect 347 12472 391 12506
rect 425 12472 469 12506
rect 503 12472 547 12506
rect 581 12472 625 12506
rect 659 12472 666 12506
rect 224 12421 666 12472
rect 224 12413 1221 12421
rect 224 12379 236 12413
rect 270 12379 309 12413
rect 343 12379 382 12413
rect 416 12379 455 12413
rect 489 12379 527 12413
rect 561 12379 599 12413
rect 633 12379 671 12413
rect 705 12379 743 12413
rect 777 12379 815 12413
rect 849 12379 887 12413
rect 921 12379 959 12413
rect 993 12379 1031 12413
rect 1065 12379 1103 12413
rect 1137 12379 1175 12413
rect 1209 12379 1221 12413
rect 224 12339 1221 12379
rect 224 12305 236 12339
rect 270 12305 309 12339
rect 343 12305 382 12339
rect 416 12305 455 12339
rect 489 12305 527 12339
rect 561 12305 599 12339
rect 633 12305 671 12339
rect 705 12305 743 12339
rect 777 12305 815 12339
rect 849 12305 887 12339
rect 921 12305 959 12339
rect 993 12305 1031 12339
rect 1065 12305 1103 12339
rect 1137 12305 1175 12339
rect 1209 12305 1221 12339
rect 224 12265 1221 12305
rect 224 12231 236 12265
rect 270 12231 309 12265
rect 343 12231 382 12265
rect 416 12231 455 12265
rect 489 12231 527 12265
rect 561 12231 599 12265
rect 633 12231 671 12265
rect 705 12231 743 12265
rect 777 12231 815 12265
rect 849 12231 887 12265
rect 921 12231 959 12265
rect 993 12231 1031 12265
rect 1065 12231 1103 12265
rect 1137 12231 1175 12265
rect 1209 12231 1221 12265
rect 224 12191 1221 12231
rect 224 12157 236 12191
rect 270 12157 309 12191
rect 343 12157 382 12191
rect 416 12157 455 12191
rect 489 12157 527 12191
rect 561 12157 599 12191
rect 633 12157 671 12191
rect 705 12157 743 12191
rect 777 12157 815 12191
rect 849 12157 887 12191
rect 921 12157 959 12191
rect 993 12157 1031 12191
rect 1065 12157 1103 12191
rect 1137 12157 1175 12191
rect 1209 12157 1221 12191
rect 224 12117 1221 12157
rect 224 12083 236 12117
rect 270 12083 309 12117
rect 343 12083 382 12117
rect 416 12083 455 12117
rect 489 12083 527 12117
rect 561 12083 599 12117
rect 633 12083 671 12117
rect 705 12083 743 12117
rect 777 12083 815 12117
rect 849 12083 887 12117
rect 921 12083 959 12117
rect 993 12083 1031 12117
rect 1065 12083 1103 12117
rect 1137 12083 1175 12117
rect 1209 12083 1221 12117
rect 224 12043 1221 12083
rect 224 12009 236 12043
rect 270 12009 309 12043
rect 343 12009 382 12043
rect 416 12009 455 12043
rect 489 12009 527 12043
rect 561 12009 599 12043
rect 633 12009 671 12043
rect 705 12009 743 12043
rect 777 12009 815 12043
rect 849 12009 887 12043
rect 921 12009 959 12043
rect 993 12009 1031 12043
rect 1065 12009 1103 12043
rect 1137 12009 1175 12043
rect 1209 12009 1221 12043
rect 224 11969 1221 12009
rect 224 11935 236 11969
rect 270 11935 309 11969
rect 343 11935 382 11969
rect 416 11935 455 11969
rect 489 11935 527 11969
rect 561 11935 599 11969
rect 633 11935 671 11969
rect 705 11935 743 11969
rect 777 11935 815 11969
rect 849 11935 887 11969
rect 921 11935 959 11969
rect 993 11935 1031 11969
rect 1065 11935 1103 11969
rect 1137 11935 1175 11969
rect 1209 11935 1221 11969
rect 224 11895 1221 11935
rect 224 11861 236 11895
rect 270 11861 309 11895
rect 343 11861 382 11895
rect 416 11861 455 11895
rect 489 11861 527 11895
rect 561 11861 599 11895
rect 633 11861 671 11895
rect 705 11861 743 11895
rect 777 11861 815 11895
rect 849 11861 887 11895
rect 921 11861 959 11895
rect 993 11861 1031 11895
rect 1065 11861 1103 11895
rect 1137 11861 1175 11895
rect 1209 11861 1221 11895
rect 224 11821 1221 11861
rect 224 11787 236 11821
rect 270 11787 309 11821
rect 343 11787 382 11821
rect 416 11787 455 11821
rect 489 11787 527 11821
rect 561 11787 599 11821
rect 633 11787 671 11821
rect 705 11787 743 11821
rect 777 11787 815 11821
rect 849 11787 887 11821
rect 921 11787 959 11821
rect 993 11787 1031 11821
rect 1065 11787 1103 11821
rect 1137 11787 1175 11821
rect 1209 11787 1221 11821
rect 224 11747 1221 11787
rect 224 11713 236 11747
rect 270 11713 309 11747
rect 343 11713 382 11747
rect 416 11713 455 11747
rect 489 11713 527 11747
rect 561 11713 599 11747
rect 633 11713 671 11747
rect 705 11713 743 11747
rect 777 11713 815 11747
rect 849 11713 887 11747
rect 921 11713 959 11747
rect 993 11713 1031 11747
rect 1065 11713 1103 11747
rect 1137 11713 1175 11747
rect 1209 11713 1221 11747
rect 224 11673 1221 11713
rect 224 11639 236 11673
rect 270 11639 309 11673
rect 343 11639 382 11673
rect 416 11639 455 11673
rect 489 11639 527 11673
rect 561 11639 599 11673
rect 633 11639 671 11673
rect 705 11639 743 11673
rect 777 11639 815 11673
rect 849 11639 887 11673
rect 921 11639 959 11673
rect 993 11639 1031 11673
rect 1065 11639 1103 11673
rect 1137 11639 1175 11673
rect 1209 11639 1221 11673
rect 224 11622 1221 11639
rect 6773 11728 7708 11734
rect 6773 11694 6785 11728
rect 6819 11694 6859 11728
rect 6893 11694 6932 11728
rect 6966 11694 7005 11728
rect 7039 11694 7078 11728
rect 7112 11694 7151 11728
rect 7185 11694 7224 11728
rect 7258 11694 7297 11728
rect 7331 11694 7370 11728
rect 7404 11694 7443 11728
rect 7477 11694 7516 11728
rect 7550 11694 7589 11728
rect 7623 11694 7662 11728
rect 7696 11723 7708 11728
rect 7696 11694 7710 11723
rect 6773 11656 7710 11694
tri 1221 11622 1235 11636 sw
rect 6773 11622 6785 11656
rect 6819 11622 6859 11656
rect 6893 11622 6932 11656
rect 6966 11622 7005 11656
rect 7039 11622 7078 11656
rect 7112 11622 7151 11656
rect 7185 11622 7224 11656
rect 7258 11622 7297 11656
rect 7331 11622 7370 11656
rect 7404 11622 7443 11656
rect 7477 11622 7516 11656
rect 7550 11622 7589 11656
rect 7623 11622 7662 11656
rect 7696 11622 7710 11656
rect 224 11617 1235 11622
tri 1235 11617 1240 11622 sw
rect 6773 11617 7710 11622
tri 7710 11617 7816 11723 sw
rect 17433 11617 18204 11623
rect 224 11599 1240 11617
rect 224 11565 236 11599
rect 270 11565 309 11599
rect 343 11565 382 11599
rect 416 11565 455 11599
rect 489 11565 527 11599
rect 561 11565 599 11599
rect 633 11565 671 11599
rect 705 11565 743 11599
rect 777 11565 815 11599
rect 849 11565 887 11599
rect 921 11565 959 11599
rect 993 11565 1031 11599
rect 1065 11565 1103 11599
rect 1137 11565 1175 11599
rect 1209 11583 1240 11599
tri 1240 11583 1274 11617 sw
rect 6773 11616 7816 11617
tri 7816 11616 7817 11617 sw
rect 6773 11604 7817 11616
rect 1209 11581 1274 11583
tri 1274 11581 1276 11583 sw
rect 1209 11579 1276 11581
tri 1276 11579 1278 11581 sw
rect 6773 11579 7173 11604
tri 7489 11583 7510 11604 ne
rect 7510 11583 7817 11604
tri 7817 11583 7850 11616 sw
rect 17433 11583 17445 11617
rect 17479 11583 17525 11617
rect 17559 11583 17605 11617
rect 17639 11583 17684 11617
rect 17718 11583 17763 11617
rect 17797 11583 17842 11617
rect 17876 11583 17921 11617
rect 17955 11583 18000 11617
rect 18034 11583 18079 11617
rect 18113 11583 18158 11617
rect 18192 11583 18204 11617
tri 7510 11581 7512 11583 ne
rect 7512 11581 9554 11583
rect 1209 11565 1278 11579
rect 224 11559 1278 11565
tri 1278 11559 1298 11579 sw
rect 224 11545 1298 11559
tri 1298 11545 1312 11559 sw
tri 1930 11545 1944 11559 se
rect 1944 11553 2064 11559
rect 224 11543 1312 11545
tri 1312 11543 1314 11545 sw
tri 1928 11543 1930 11545 se
rect 1930 11543 1944 11545
rect 224 11533 1314 11543
tri 1314 11533 1324 11543 sw
tri 1918 11533 1928 11543 se
rect 1928 11533 1944 11543
rect 224 11525 1944 11533
rect 224 11491 236 11525
rect 270 11491 309 11525
rect 343 11491 382 11525
rect 416 11491 455 11525
rect 489 11491 527 11525
rect 561 11491 599 11525
rect 633 11491 671 11525
rect 705 11491 743 11525
rect 777 11491 815 11525
rect 849 11491 887 11525
rect 921 11491 959 11525
rect 993 11491 1031 11525
rect 1065 11491 1103 11525
rect 1137 11491 1175 11525
rect 1209 11501 1944 11525
rect 1996 11501 2012 11553
rect 1209 11491 2064 11501
rect 224 11485 2064 11491
rect 224 11483 1944 11485
tri 861 11473 871 11483 ne
rect 871 11473 1944 11483
tri 871 11455 889 11473 ne
rect 889 11455 1944 11473
tri 889 11452 892 11455 ne
rect 892 11452 1944 11455
tri 892 11435 909 11452 ne
rect 909 11435 1944 11452
tri 909 11401 943 11435 ne
rect 943 11433 1944 11435
rect 1996 11433 2012 11485
rect 943 11417 2064 11433
rect 943 11401 1944 11417
tri 943 11367 977 11401 ne
rect 977 11367 1944 11401
tri 977 11365 979 11367 ne
rect 979 11365 1944 11367
rect 1996 11365 2012 11417
tri 979 11363 981 11365 ne
rect 981 11363 2064 11365
tri 981 11358 986 11363 ne
rect 986 11358 2064 11363
tri 1876 11329 1905 11358 ne
rect 1905 11348 2064 11358
rect 1905 11329 1944 11348
tri 1905 11313 1921 11329 ne
rect 1921 11313 1944 11329
tri 1921 11291 1943 11313 ne
rect 1943 11296 1944 11313
rect 1996 11296 2012 11348
rect 1943 11291 2064 11296
tri 1943 11290 1944 11291 ne
rect 1944 11290 2064 11291
rect 6773 11545 6779 11579
rect 6813 11545 6867 11579
rect 6901 11545 6955 11579
rect 6989 11545 7043 11579
rect 7077 11545 7131 11579
rect 7165 11545 7173 11579
tri 7512 11577 7516 11581 ne
rect 7516 11577 9554 11581
rect 6773 11507 7173 11545
tri 7516 11543 7550 11577 ne
rect 7550 11543 7577 11577
rect 7611 11543 7651 11577
rect 7685 11543 7725 11577
rect 7759 11543 7799 11577
rect 7833 11543 7873 11577
rect 7907 11543 7947 11577
rect 7981 11543 8021 11577
rect 8055 11543 8095 11577
rect 8129 11543 8169 11577
rect 8203 11543 8243 11577
rect 8277 11543 8317 11577
rect 8351 11543 8391 11577
rect 8425 11543 8465 11577
rect 8499 11543 8539 11577
rect 8573 11543 8613 11577
rect 8647 11543 8687 11577
rect 8721 11543 8761 11577
rect 8795 11543 8835 11577
rect 8869 11543 8909 11577
rect 8943 11543 8983 11577
rect 9017 11543 9058 11577
rect 9092 11543 9133 11577
rect 9167 11543 9208 11577
rect 9242 11543 9283 11577
rect 9317 11543 9358 11577
rect 9392 11543 9433 11577
rect 9467 11543 9508 11577
rect 9542 11543 9554 11577
tri 7550 11528 7565 11543 ne
rect 6773 11473 6779 11507
rect 6813 11473 6867 11507
rect 6901 11473 6955 11507
rect 6989 11473 7043 11507
rect 7077 11473 7131 11507
rect 7165 11473 7173 11507
rect 6773 11435 7173 11473
rect 6773 11401 6779 11435
rect 6813 11401 6867 11435
rect 6901 11401 6955 11435
rect 6989 11401 7043 11435
rect 7077 11401 7131 11435
rect 7165 11401 7173 11435
rect 6773 11363 7173 11401
rect 6773 11329 6779 11363
rect 6813 11329 6867 11363
rect 6901 11329 6955 11363
rect 6989 11329 7043 11363
rect 7077 11329 7131 11363
rect 7165 11329 7173 11363
rect 6773 11291 7173 11329
rect 6773 11257 6779 11291
rect 6813 11257 6867 11291
rect 6901 11257 6955 11291
rect 6989 11257 7043 11291
rect 7077 11257 7131 11291
rect 7165 11257 7173 11291
rect 6773 11219 7173 11257
rect 6773 11185 6779 11219
rect 6813 11185 6867 11219
rect 6901 11185 6955 11219
rect 6989 11185 7043 11219
rect 7077 11185 7131 11219
rect 7165 11185 7173 11219
rect 7565 11489 9554 11543
rect 7565 11455 7577 11489
rect 7611 11455 7651 11489
rect 7685 11455 7725 11489
rect 7759 11455 7799 11489
rect 7833 11455 7873 11489
rect 7907 11455 7947 11489
rect 7981 11455 8021 11489
rect 8055 11455 8095 11489
rect 8129 11455 8169 11489
rect 8203 11455 8243 11489
rect 8277 11455 8317 11489
rect 8351 11455 8391 11489
rect 8425 11455 8465 11489
rect 8499 11455 8539 11489
rect 8573 11455 8613 11489
rect 8647 11455 8687 11489
rect 8721 11455 8761 11489
rect 8795 11455 8835 11489
rect 8869 11455 8909 11489
rect 8943 11455 8983 11489
rect 9017 11455 9058 11489
rect 9092 11455 9133 11489
rect 9167 11455 9208 11489
rect 9242 11455 9283 11489
rect 9317 11455 9358 11489
rect 9392 11455 9433 11489
rect 9467 11455 9508 11489
rect 9542 11455 9554 11489
rect 17433 11545 18204 11583
rect 17433 11511 17445 11545
rect 17479 11511 17525 11545
rect 17559 11511 17605 11545
rect 17639 11511 17684 11545
rect 17718 11511 17763 11545
rect 17797 11511 17842 11545
rect 17876 11511 17921 11545
rect 17955 11511 18000 11545
rect 18034 11511 18079 11545
rect 18113 11511 18158 11545
rect 18192 11511 18204 11545
rect 17433 11473 18204 11511
rect 7565 11401 9554 11455
rect 7565 11367 7577 11401
rect 7611 11367 7651 11401
rect 7685 11367 7725 11401
rect 7759 11367 7799 11401
rect 7833 11367 7873 11401
rect 7907 11367 7947 11401
rect 7981 11367 8021 11401
rect 8055 11367 8095 11401
rect 8129 11367 8169 11401
rect 8203 11367 8243 11401
rect 8277 11367 8317 11401
rect 8351 11367 8391 11401
rect 8425 11367 8465 11401
rect 8499 11367 8539 11401
rect 8573 11367 8613 11401
rect 8647 11367 8687 11401
rect 8721 11367 8761 11401
rect 8795 11367 8835 11401
rect 8869 11367 8909 11401
rect 8943 11367 8983 11401
rect 9017 11367 9058 11401
rect 9092 11367 9133 11401
rect 9167 11367 9208 11401
rect 9242 11367 9283 11401
rect 9317 11367 9358 11401
rect 9392 11367 9433 11401
rect 9467 11367 9508 11401
rect 9542 11367 9554 11401
rect 7565 11313 9554 11367
rect 7565 11279 7577 11313
rect 7611 11279 7651 11313
rect 7685 11279 7725 11313
rect 7759 11279 7799 11313
rect 7833 11279 7873 11313
rect 7907 11279 7947 11313
rect 7981 11279 8021 11313
rect 8055 11279 8095 11313
rect 8129 11279 8169 11313
rect 8203 11279 8243 11313
rect 8277 11279 8317 11313
rect 8351 11279 8391 11313
rect 8425 11279 8465 11313
rect 8499 11279 8539 11313
rect 8573 11279 8613 11313
rect 8647 11279 8687 11313
rect 8721 11279 8761 11313
rect 8795 11279 8835 11313
rect 8869 11279 8909 11313
rect 8943 11279 8983 11313
rect 9017 11279 9058 11313
rect 9092 11279 9133 11313
rect 9167 11279 9208 11313
rect 9242 11279 9283 11313
rect 9317 11279 9358 11313
rect 9392 11279 9433 11313
rect 9467 11279 9508 11313
rect 9542 11279 9554 11313
rect 10444 11452 12379 11458
rect 10444 11418 10456 11452
rect 10490 11418 10529 11452
rect 10563 11418 10602 11452
rect 10636 11418 10675 11452
rect 10709 11418 10748 11452
rect 10782 11418 10821 11452
rect 10855 11418 10893 11452
rect 10927 11418 10965 11452
rect 10999 11418 11037 11452
rect 11071 11418 11109 11452
rect 11143 11418 11181 11452
rect 11215 11418 11253 11452
rect 11287 11418 11325 11452
rect 11359 11418 11397 11452
rect 11431 11418 11469 11452
rect 11503 11418 11541 11452
rect 11575 11418 11613 11452
rect 11647 11418 11685 11452
rect 11719 11418 11757 11452
rect 11791 11418 11829 11452
rect 11863 11418 11901 11452
rect 11935 11418 11973 11452
rect 12007 11418 12045 11452
rect 12079 11418 12117 11452
rect 12151 11418 12189 11452
rect 12223 11418 12261 11452
rect 12295 11418 12333 11452
rect 12367 11418 12379 11452
rect 10444 11367 12379 11418
rect 13399 11452 15659 11458
rect 13399 11418 13411 11452
rect 13445 11418 13485 11452
rect 13519 11418 13559 11452
rect 13593 11418 13633 11452
rect 13667 11418 13707 11452
rect 13741 11418 13781 11452
rect 13815 11418 13855 11452
rect 13889 11418 13929 11452
rect 13963 11418 14003 11452
rect 14037 11418 14077 11452
rect 14111 11418 14151 11452
rect 14185 11418 14225 11452
rect 14259 11418 14299 11452
rect 14333 11418 14372 11452
rect 14406 11418 14445 11452
rect 14479 11418 14518 11452
rect 14552 11418 14591 11452
rect 14625 11418 14664 11452
rect 14698 11418 14737 11452
rect 14771 11418 14810 11452
rect 14844 11418 14883 11452
rect 14917 11418 14956 11452
rect 14990 11418 15029 11452
rect 15063 11418 15102 11452
rect 15136 11418 15175 11452
rect 15209 11418 15248 11452
rect 15282 11418 15321 11452
rect 15355 11418 15394 11452
rect 15428 11418 15467 11452
rect 15501 11418 15540 11452
rect 15574 11418 15613 11452
rect 15647 11418 15659 11452
tri 12379 11367 12390 11378 sw
rect 10444 11365 12390 11367
tri 12390 11365 12392 11367 sw
rect 10444 11347 12392 11365
tri 12392 11347 12410 11365 sw
rect 10444 11338 12410 11347
tri 12410 11338 12419 11347 sw
tri 13390 11338 13399 11347 se
rect 13399 11338 15659 11418
rect 10444 11304 10456 11338
rect 10490 11304 10529 11338
rect 10563 11304 10602 11338
rect 10636 11304 10675 11338
rect 10709 11304 10748 11338
rect 10782 11304 10821 11338
rect 10855 11304 10893 11338
rect 10927 11304 10965 11338
rect 10999 11304 11037 11338
rect 11071 11304 11109 11338
rect 11143 11304 11181 11338
rect 11215 11304 11253 11338
rect 11287 11304 11325 11338
rect 11359 11304 11397 11338
rect 11431 11304 11469 11338
rect 11503 11304 11541 11338
rect 11575 11304 11613 11338
rect 11647 11304 11685 11338
rect 11719 11304 11757 11338
rect 11791 11304 11829 11338
rect 11863 11304 11901 11338
rect 11935 11304 11973 11338
rect 12007 11304 12045 11338
rect 12079 11304 12117 11338
rect 12151 11304 12189 11338
rect 12223 11304 12261 11338
rect 12295 11304 12333 11338
rect 12367 11304 12419 11338
tri 12419 11304 12453 11338 sw
tri 13356 11304 13390 11338 se
rect 13390 11304 13411 11338
rect 13445 11304 13485 11338
rect 13519 11304 13559 11338
rect 13593 11304 13633 11338
rect 13667 11304 13707 11338
rect 13741 11304 13781 11338
rect 13815 11304 13855 11338
rect 13889 11304 13929 11338
rect 13963 11304 14003 11338
rect 14037 11304 14077 11338
rect 14111 11304 14151 11338
rect 14185 11304 14225 11338
rect 14259 11304 14299 11338
rect 14333 11304 14372 11338
rect 14406 11304 14445 11338
rect 14479 11304 14518 11338
rect 14552 11304 14591 11338
rect 14625 11304 14664 11338
rect 14698 11304 14737 11338
rect 14771 11304 14810 11338
rect 14844 11304 14883 11338
rect 14917 11304 14956 11338
rect 14990 11304 15029 11338
rect 15063 11304 15102 11338
rect 15136 11304 15175 11338
rect 15209 11304 15248 11338
rect 15282 11304 15321 11338
rect 15355 11304 15394 11338
rect 15428 11304 15467 11338
rect 15501 11304 15540 11338
rect 15574 11304 15613 11338
rect 15647 11304 15659 11338
rect 10444 11297 12453 11304
tri 12453 11297 12460 11304 sw
tri 13349 11297 13356 11304 se
rect 13356 11298 15659 11304
rect 17433 11439 17445 11473
rect 17479 11439 17525 11473
rect 17559 11439 17605 11473
rect 17639 11439 17684 11473
rect 17718 11439 17763 11473
rect 17797 11439 17842 11473
rect 17876 11439 17921 11473
rect 17955 11439 18000 11473
rect 18034 11439 18079 11473
rect 18113 11439 18158 11473
rect 18192 11439 18204 11473
rect 17433 11401 18204 11439
rect 17433 11367 17445 11401
rect 17479 11367 17525 11401
rect 17559 11367 17605 11401
rect 17639 11367 17684 11401
rect 17718 11367 17763 11401
rect 17797 11367 17842 11401
rect 17876 11367 17921 11401
rect 17955 11367 18000 11401
rect 18034 11367 18079 11401
rect 18113 11367 18158 11401
rect 18192 11367 18204 11401
rect 17433 11329 18204 11367
rect 13356 11297 14190 11298
tri 14190 11297 14191 11298 nw
tri 14934 11297 14935 11298 ne
rect 14935 11297 15052 11298
rect 10444 11295 12460 11297
tri 12460 11295 12462 11297 sw
rect 13131 11295 14188 11297
tri 14188 11295 14190 11297 nw
tri 14935 11295 14937 11297 ne
rect 14937 11295 15052 11297
tri 15052 11295 15055 11298 nw
rect 17433 11295 17445 11329
rect 17479 11295 17525 11329
rect 17559 11295 17605 11329
rect 17639 11295 17684 11329
rect 17718 11295 17763 11329
rect 17797 11295 17842 11329
rect 17876 11295 17921 11329
rect 17955 11295 18000 11329
rect 18034 11295 18079 11329
rect 18113 11295 18158 11329
rect 18192 11295 18204 11329
rect 10444 11293 12462 11295
tri 12462 11293 12464 11295 sw
rect 13131 11293 14186 11295
tri 14186 11293 14188 11295 nw
tri 14937 11293 14939 11295 ne
rect 14939 11293 15050 11295
tri 15050 11293 15052 11295 nw
rect 10444 11286 12464 11293
tri 12464 11286 12471 11293 sw
rect 7565 11225 9554 11279
rect 7565 11191 7577 11225
rect 7611 11191 7651 11225
rect 7685 11191 7725 11225
rect 7759 11191 7799 11225
rect 7833 11191 7873 11225
rect 7907 11191 7947 11225
rect 7981 11191 8021 11225
rect 8055 11191 8095 11225
rect 8129 11191 8169 11225
rect 8203 11191 8243 11225
rect 8277 11191 8317 11225
rect 8351 11191 8391 11225
rect 8425 11191 8465 11225
rect 8499 11191 8539 11225
rect 8573 11191 8613 11225
rect 8647 11191 8687 11225
rect 8721 11191 8761 11225
rect 8795 11191 8835 11225
rect 8869 11191 8909 11225
rect 8943 11191 8983 11225
rect 9017 11191 9058 11225
rect 9092 11191 9133 11225
rect 9167 11191 9208 11225
rect 9242 11191 9283 11225
rect 9317 11191 9358 11225
rect 9392 11191 9433 11225
rect 9467 11191 9508 11225
rect 9542 11191 9554 11225
rect 13131 11283 14176 11293
tri 14176 11283 14186 11293 nw
tri 14939 11283 14949 11293 ne
rect 14949 11283 15040 11293
tri 15040 11283 15050 11293 nw
rect 13131 11257 14150 11283
tri 14150 11257 14176 11283 nw
tri 14949 11266 14966 11283 ne
rect 14966 11266 15023 11283
tri 15023 11266 15040 11283 nw
rect 17433 11257 18204 11295
rect 13131 11223 14116 11257
tri 14116 11223 14150 11257 nw
rect 17433 11223 17445 11257
rect 17479 11223 17525 11257
rect 17559 11223 17605 11257
rect 17639 11223 17684 11257
rect 17718 11223 17763 11257
rect 17797 11223 17842 11257
rect 17876 11223 17921 11257
rect 17955 11252 18000 11257
rect 18034 11252 18079 11257
rect 18113 11252 18158 11257
rect 18192 11252 18204 11257
rect 18068 11223 18079 11252
rect 13131 11221 14114 11223
tri 14114 11221 14116 11223 nw
rect 13131 11208 14101 11221
tri 14101 11208 14114 11221 nw
rect 13131 11199 14092 11208
tri 14092 11199 14101 11208 nw
rect 17433 11200 17950 11223
rect 18002 11200 18016 11223
rect 18068 11200 18081 11223
rect 18133 11200 18146 11252
rect 18198 11200 18204 11252
rect 7565 11185 9554 11191
rect 17433 11185 18204 11200
rect 6773 11147 7173 11185
rect 6773 11113 6779 11147
rect 6813 11113 6867 11147
rect 6901 11113 6955 11147
rect 6989 11113 7043 11147
rect 7077 11113 7131 11147
rect 7165 11113 7173 11147
rect 17433 11151 17445 11185
rect 17479 11151 17525 11185
rect 17559 11151 17605 11185
rect 17639 11151 17684 11185
rect 17718 11151 17763 11185
rect 17797 11151 17842 11185
rect 17876 11151 17921 11185
rect 17955 11151 18000 11185
rect 18034 11151 18079 11185
rect 18113 11151 18158 11185
rect 18192 11151 18204 11185
rect 17433 11145 18204 11151
rect 18488 11615 18967 11621
rect 18488 11581 18500 11615
rect 18534 11581 18585 11615
rect 18619 11581 18669 11615
rect 18703 11581 18753 11615
rect 18787 11581 18837 11615
rect 18871 11581 18921 11615
rect 18955 11581 18967 11615
rect 18488 11543 18967 11581
rect 18488 11509 18500 11543
rect 18534 11509 18585 11543
rect 18619 11509 18669 11543
rect 18703 11509 18753 11543
rect 18787 11509 18837 11543
rect 18871 11509 18921 11543
rect 18955 11509 18967 11543
rect 18488 11471 18967 11509
rect 18488 11437 18500 11471
rect 18534 11437 18585 11471
rect 18619 11437 18669 11471
rect 18703 11437 18753 11471
rect 18787 11437 18837 11471
rect 18871 11437 18921 11471
rect 18955 11437 18967 11471
rect 18488 11399 18967 11437
rect 18488 11365 18500 11399
rect 18534 11365 18585 11399
rect 18619 11365 18669 11399
rect 18703 11365 18753 11399
rect 18787 11365 18837 11399
rect 18871 11365 18921 11399
rect 18955 11365 18967 11399
rect 18488 11327 18967 11365
rect 18488 11293 18500 11327
rect 18534 11293 18585 11327
rect 18619 11293 18669 11327
rect 18703 11293 18753 11327
rect 18787 11293 18837 11327
rect 18871 11293 18921 11327
rect 18955 11293 18967 11327
rect 18488 11255 18967 11293
rect 19552 11384 19751 11503
rect 19552 11317 19644 11384
tri 19544 11283 19552 11291 se
rect 19552 11283 19581 11317
rect 19615 11283 19644 11317
tri 19527 11266 19544 11283 se
rect 19544 11266 19644 11283
rect 18488 11252 18500 11255
rect 18534 11252 18585 11255
rect 18619 11252 18669 11255
rect 18703 11252 18753 11255
rect 18488 11200 18494 11252
rect 18546 11200 18560 11252
rect 18619 11221 18625 11252
rect 18742 11221 18753 11252
rect 18787 11221 18837 11255
rect 18871 11221 18921 11255
rect 18955 11221 18967 11255
tri 19513 11252 19527 11266 se
rect 19527 11252 19644 11266
rect 18612 11200 18625 11221
rect 18677 11200 18690 11221
rect 18742 11200 18967 11221
rect 19211 11200 19217 11252
rect 19269 11200 19283 11252
rect 19335 11200 19348 11252
rect 19400 11200 19413 11252
rect 19465 11242 19644 11252
rect 19465 11208 19581 11242
rect 19615 11208 19644 11242
rect 19465 11200 19644 11208
rect 18488 11183 18967 11200
tri 19514 11199 19515 11200 ne
rect 19515 11199 19644 11200
tri 19515 11185 19529 11199 ne
rect 19529 11185 19644 11199
rect 18488 11149 18500 11183
rect 18534 11149 18585 11183
rect 18619 11149 18669 11183
rect 18703 11149 18753 11183
rect 18787 11149 18837 11183
rect 18871 11149 18921 11183
rect 18955 11149 18967 11183
tri 19529 11167 19547 11185 ne
rect 19547 11167 19644 11185
tri 19547 11162 19552 11167 ne
rect 18488 11143 18967 11149
rect 6773 11075 7173 11113
rect 6773 11041 6779 11075
rect 6813 11041 6867 11075
rect 6901 11041 6955 11075
rect 6989 11041 7043 11075
rect 7077 11041 7131 11075
rect 7165 11041 7173 11075
rect 6773 11002 7173 11041
rect 6773 10968 6779 11002
rect 6813 10968 6867 11002
rect 6901 10968 6955 11002
rect 6989 10968 7043 11002
rect 7077 10968 7131 11002
rect 7165 10968 7173 11002
rect 6773 10929 7173 10968
rect 6773 10895 6779 10929
rect 6813 10895 6867 10929
rect 6901 10895 6955 10929
rect 6989 10895 7043 10929
rect 7077 10895 7131 10929
rect 7165 10895 7173 10929
rect 6773 10856 7173 10895
rect 6773 10822 6779 10856
rect 6813 10822 6867 10856
rect 6901 10822 6955 10856
rect 6989 10822 7043 10856
rect 7077 10822 7131 10856
rect 7165 10822 7173 10856
rect 6773 10787 7173 10822
rect 19552 11133 19581 11167
rect 19615 11133 19644 11167
rect 19552 11091 19644 11133
rect 19552 11057 19581 11091
rect 19615 11057 19644 11091
rect 19552 11015 19644 11057
rect 19552 10981 19581 11015
rect 19615 10981 19644 11015
rect 19552 10939 19644 10981
rect 19552 10905 19581 10939
rect 19615 10905 19644 10939
rect 19552 10863 19644 10905
rect 19552 10829 19581 10863
rect 19615 10829 19644 10863
tri 7173 10787 7203 10817 sw
rect 19552 10787 19644 10829
rect 6773 10783 7203 10787
rect 6773 10749 6779 10783
rect 6813 10749 6867 10783
rect 6901 10749 6955 10783
rect 6989 10749 7043 10783
rect 7077 10749 7131 10783
rect 7165 10763 7203 10783
tri 7203 10763 7227 10787 sw
rect 7165 10749 7227 10763
rect 6773 10737 7227 10749
tri 7065 10711 7091 10737 ne
rect 7091 10711 7227 10737
tri 7091 10699 7103 10711 ne
rect 7103 10699 7227 10711
rect 19552 10753 19581 10787
rect 19615 10753 19644 10787
rect 19552 10711 19644 10753
tri 7103 10696 7106 10699 ne
rect 7106 10696 7227 10699
tri 7106 10662 7140 10696 ne
rect 7140 10662 7155 10696
rect 7189 10662 7227 10696
tri 7140 10653 7149 10662 ne
rect 7149 10620 7227 10662
rect 7149 10586 7155 10620
rect 7189 10586 7227 10620
rect 7149 10544 7227 10586
rect 7149 10510 7155 10544
rect 7189 10510 7227 10544
rect 7149 10468 7227 10510
rect 7149 10434 7155 10468
rect 7189 10434 7227 10468
rect 7149 10392 7227 10434
rect 7149 10358 7155 10392
rect 7189 10365 7227 10392
rect 10066 10687 10218 10699
rect 10066 10653 10072 10687
rect 10106 10653 10178 10687
rect 10212 10653 10218 10687
rect 10066 10615 10218 10653
rect 10066 10581 10072 10615
rect 10106 10581 10178 10615
rect 10212 10581 10218 10615
rect 10066 10543 10218 10581
rect 10066 10509 10072 10543
rect 10106 10509 10178 10543
rect 10212 10509 10218 10543
rect 10066 10471 10218 10509
rect 10066 10437 10072 10471
rect 10106 10437 10178 10471
rect 10212 10437 10218 10471
rect 10066 10399 10218 10437
tri 7227 10365 7233 10371 sw
rect 10066 10365 10072 10399
rect 10106 10365 10178 10399
rect 10212 10365 10218 10399
rect 7189 10358 7233 10365
rect 7149 10341 7233 10358
tri 7233 10341 7257 10365 sw
rect 7149 10332 7257 10341
tri 7257 10332 7266 10341 sw
rect 7149 10331 7266 10332
tri 7266 10331 7267 10332 sw
rect 7149 10327 7267 10331
tri 7267 10327 7271 10331 sw
rect 10066 10327 10218 10365
rect 7149 10316 7271 10327
rect 7149 10282 7155 10316
rect 7189 10293 7271 10316
tri 7271 10293 7305 10327 sw
rect 10066 10293 10072 10327
rect 10106 10293 10178 10327
rect 10212 10293 10218 10327
rect 7189 10282 7305 10293
rect 7149 10273 7305 10282
tri 7305 10273 7325 10293 sw
rect 7149 10261 7329 10273
rect 7149 10240 7266 10261
rect 7149 10206 7155 10240
rect 7189 10227 7266 10240
rect 7300 10227 7329 10261
rect 7189 10206 7329 10227
rect 7149 10189 7329 10206
rect 7149 10164 7266 10189
rect 7149 10130 7155 10164
rect 7189 10155 7266 10164
rect 7300 10155 7329 10189
rect 7189 10130 7329 10155
rect 7149 10117 7329 10130
rect 7149 10088 7266 10117
rect 7149 10054 7155 10088
rect 7189 10083 7266 10088
rect 7300 10083 7329 10117
rect 7189 10054 7329 10083
rect 7149 10045 7329 10054
rect 7149 10012 7266 10045
rect 7149 9978 7155 10012
rect 7189 10011 7266 10012
rect 7300 10011 7329 10045
rect 7189 9978 7329 10011
rect 7149 9973 7329 9978
rect 7149 9939 7266 9973
rect 7300 9939 7329 9973
rect 7149 9935 7329 9939
rect 7149 9901 7155 9935
rect 7189 9901 7329 9935
rect 7149 9867 7266 9901
rect 7300 9867 7329 9901
rect 7149 9858 7329 9867
rect 7149 9824 7155 9858
rect 7189 9829 7329 9858
rect 7189 9824 7266 9829
rect 7149 9795 7266 9824
rect 7300 9795 7329 9829
rect 7149 9781 7329 9795
rect 7149 9747 7155 9781
rect 7189 9757 7329 9781
rect 7189 9747 7266 9757
rect 7149 9723 7266 9747
rect 7300 9751 7329 9757
rect 10066 10255 10218 10293
rect 10066 10221 10072 10255
rect 10106 10221 10178 10255
rect 10212 10221 10218 10255
rect 10066 10183 10218 10221
rect 10066 10149 10072 10183
rect 10106 10149 10178 10183
rect 10212 10149 10218 10183
rect 19552 10677 19581 10711
rect 19615 10677 19644 10711
rect 19552 10635 19644 10677
rect 19552 10601 19581 10635
rect 19615 10601 19644 10635
rect 19552 10559 19644 10601
rect 19552 10525 19581 10559
rect 19615 10525 19644 10559
rect 19552 10483 19644 10525
rect 19552 10449 19581 10483
rect 19615 10449 19644 10483
rect 19552 10407 19644 10449
rect 19552 10373 19581 10407
rect 19615 10373 19644 10407
rect 19552 10331 19644 10373
rect 19552 10297 19581 10331
rect 19615 10297 19644 10331
rect 19552 10255 19644 10297
rect 19552 10221 19581 10255
rect 19615 10221 19644 10255
rect 19552 10179 19644 10221
rect 10066 10111 10218 10149
rect 10066 10077 10072 10111
rect 10106 10077 10178 10111
rect 10212 10077 10218 10111
rect 10066 10039 10218 10077
rect 10066 10005 10072 10039
rect 10106 10005 10178 10039
rect 10212 10005 10218 10039
rect 16696 10154 16901 10160
rect 16696 10120 16708 10154
rect 16742 10120 16781 10154
rect 16888 10120 16901 10154
rect 16696 10102 16811 10120
rect 16863 10102 16901 10120
rect 16696 10090 16901 10102
rect 16696 10082 16811 10090
rect 16863 10082 16901 10090
rect 16696 10048 16708 10082
rect 16742 10048 16781 10082
rect 16888 10048 16901 10082
rect 16696 10038 16811 10048
rect 16863 10038 16901 10048
rect 16696 10032 16901 10038
rect 19552 10145 19581 10179
rect 19615 10145 19644 10179
rect 19552 10103 19644 10145
rect 26260 10341 27974 10353
rect 26260 10332 27501 10341
rect 26260 10298 26272 10332
rect 26306 10298 26348 10332
rect 26382 10298 26424 10332
rect 26458 10298 26500 10332
rect 26534 10298 26576 10332
rect 26610 10298 26652 10332
rect 26686 10298 26727 10332
rect 26761 10298 26802 10332
rect 26836 10298 26877 10332
rect 26911 10298 26952 10332
rect 26986 10298 27027 10332
rect 27061 10298 27102 10332
rect 27136 10298 27177 10332
rect 27211 10298 27252 10332
rect 27286 10298 27327 10332
rect 27361 10298 27402 10332
rect 27436 10331 27501 10332
rect 27535 10331 27573 10341
rect 27607 10331 27645 10341
rect 27679 10331 27717 10341
rect 27751 10331 27789 10341
rect 27436 10298 27498 10331
rect 27823 10307 27861 10341
rect 27895 10307 27974 10341
rect 26260 10260 27498 10298
rect 27806 10268 27974 10307
rect 26260 10226 26272 10260
rect 26306 10226 26348 10260
rect 26382 10226 26424 10260
rect 26458 10226 26500 10260
rect 26534 10226 26576 10260
rect 26610 10226 26652 10260
rect 26686 10226 26727 10260
rect 26761 10226 26802 10260
rect 26836 10226 26877 10260
rect 26911 10226 26952 10260
rect 26986 10226 27027 10260
rect 27061 10226 27102 10260
rect 27136 10226 27177 10260
rect 27211 10226 27252 10260
rect 27286 10226 27327 10260
rect 27361 10226 27402 10260
rect 27436 10226 27498 10260
rect 27823 10234 27861 10268
rect 27895 10234 27974 10268
rect 26260 10188 27498 10226
rect 27806 10195 27974 10234
rect 26260 10154 26272 10188
rect 26306 10154 26348 10188
rect 26382 10154 26424 10188
rect 26458 10154 26500 10188
rect 26534 10154 26576 10188
rect 26610 10154 26652 10188
rect 26686 10154 26727 10188
rect 26761 10154 26802 10188
rect 26836 10154 26877 10188
rect 26911 10154 26952 10188
rect 26986 10154 27027 10188
rect 27061 10154 27102 10188
rect 27136 10154 27177 10188
rect 27211 10154 27252 10188
rect 27286 10154 27327 10188
rect 27361 10154 27402 10188
rect 27436 10154 27498 10188
rect 27823 10161 27861 10195
rect 27895 10161 27974 10195
rect 26260 10116 27498 10154
rect 27806 10122 27974 10161
rect 19552 10069 19581 10103
rect 19615 10069 19644 10103
tri 26227 10082 26260 10115 se
rect 26260 10082 26272 10116
rect 26306 10082 26348 10116
rect 26382 10082 26424 10116
rect 26458 10082 26500 10116
rect 26534 10082 26576 10116
rect 26610 10082 26652 10116
rect 26686 10082 26727 10116
rect 26761 10082 26802 10116
rect 26836 10082 26877 10116
rect 26911 10082 26952 10116
rect 26986 10082 27027 10116
rect 27061 10082 27102 10116
rect 27136 10082 27177 10116
rect 27211 10082 27252 10116
rect 27286 10082 27327 10116
rect 27361 10082 27402 10116
rect 27436 10082 27498 10116
rect 27823 10088 27861 10122
rect 27895 10088 27974 10122
rect 10066 9967 10218 10005
rect 10066 9933 10072 9967
rect 10106 9933 10178 9967
rect 10212 9933 10218 9967
rect 10066 9895 10218 9933
rect 19552 10027 19644 10069
tri 26194 10049 26227 10082 se
rect 26227 10049 27498 10082
rect 27806 10049 27974 10088
tri 26189 10044 26194 10049 se
rect 26194 10044 27498 10049
rect 19552 9993 19581 10027
rect 19615 9993 19644 10027
tri 26155 10010 26189 10044 se
rect 26189 10010 26272 10044
rect 26306 10010 26348 10044
rect 26382 10010 26424 10044
rect 26458 10010 26500 10044
rect 26534 10010 26576 10044
rect 26610 10010 26652 10044
rect 26686 10010 26727 10044
rect 26761 10010 26802 10044
rect 26836 10010 26877 10044
rect 26911 10010 26952 10044
rect 26986 10010 27027 10044
rect 27061 10010 27102 10044
rect 27136 10010 27177 10044
rect 27211 10010 27252 10044
rect 27286 10010 27327 10044
rect 27361 10010 27402 10044
rect 27436 10010 27498 10044
rect 27823 10015 27861 10049
rect 27895 10015 27974 10049
rect 19552 9951 19644 9993
tri 26121 9976 26155 10010 se
rect 26155 9976 27498 10010
rect 27806 9976 27974 10015
tri 26117 9972 26121 9976 se
rect 26121 9972 27498 9976
rect 19552 9917 19581 9951
rect 19615 9917 19644 9951
tri 26083 9938 26117 9972 se
rect 26117 9938 26272 9972
rect 26306 9938 26348 9972
rect 26382 9938 26424 9972
rect 26458 9938 26500 9972
rect 26534 9938 26576 9972
rect 26610 9938 26652 9972
rect 26686 9938 26727 9972
rect 26761 9938 26802 9972
rect 26836 9938 26877 9972
rect 26911 9938 26952 9972
rect 26986 9938 27027 9972
rect 27061 9938 27102 9972
rect 27136 9938 27177 9972
rect 27211 9938 27252 9972
rect 27286 9938 27327 9972
rect 27361 9938 27402 9972
rect 27436 9938 27498 9972
rect 27823 9942 27861 9976
rect 27895 9942 27974 9976
rect 19552 9905 19644 9917
tri 26050 9905 26083 9938 se
rect 26083 9905 27498 9938
tri 26047 9902 26050 9905 se
rect 26050 9902 27498 9905
rect 27806 9902 27974 9942
tri 26045 9900 26047 9902 se
rect 26047 9900 27498 9902
rect 10066 9861 10072 9895
rect 10106 9861 10178 9895
rect 10212 9861 10218 9895
tri 26028 9883 26045 9900 se
rect 26045 9883 26272 9900
rect 10066 9828 10218 9861
rect 25277 9866 26272 9883
rect 26306 9866 26348 9900
rect 26382 9866 26424 9900
rect 26458 9866 26500 9900
rect 26534 9866 26576 9900
rect 26610 9866 26652 9900
rect 26686 9866 26727 9900
rect 26761 9866 26802 9900
rect 26836 9866 26877 9900
rect 26911 9866 26952 9900
rect 26986 9866 27027 9900
rect 27061 9866 27102 9900
rect 27136 9866 27177 9900
rect 27211 9866 27252 9900
rect 27286 9866 27327 9900
rect 27361 9866 27402 9900
rect 27436 9866 27498 9900
rect 27823 9868 27861 9902
rect 27895 9868 27974 9902
rect 25277 9860 27498 9866
rect 25277 9858 26423 9860
tri 26423 9858 26425 9860 nw
tri 10218 9828 10248 9858 sw
rect 25277 9828 26393 9858
tri 26393 9828 26423 9858 nw
rect 10066 9823 10248 9828
rect 10066 9789 10072 9823
rect 10106 9789 10178 9823
rect 10212 9803 10248 9823
tri 10248 9803 10273 9828 sw
rect 25277 9803 26368 9828
tri 26368 9803 26393 9828 nw
rect 10212 9789 10444 9803
tri 7329 9751 7331 9753 sw
rect 10066 9751 10444 9789
rect 25277 9794 26359 9803
tri 26359 9794 26368 9803 nw
rect 25277 9766 26331 9794
tri 26331 9766 26359 9794 nw
rect 7300 9723 7331 9751
rect 7149 9717 7331 9723
tri 7331 9717 7365 9751 sw
rect 10066 9717 10072 9751
rect 10106 9717 10178 9751
rect 10212 9717 10444 9751
rect 7149 9705 7365 9717
tri 7365 9705 7377 9717 sw
rect 7149 9704 9197 9705
rect 7149 9670 7155 9704
rect 7189 9699 9197 9704
rect 7189 9685 7360 9699
rect 7189 9670 7266 9685
rect 7149 9651 7266 9670
rect 7300 9665 7360 9685
rect 7394 9665 7435 9699
rect 7469 9665 7510 9699
rect 7544 9665 7585 9699
rect 7619 9665 7660 9699
rect 7694 9665 7735 9699
rect 7769 9665 7810 9699
rect 7844 9665 7885 9699
rect 7919 9665 7960 9699
rect 7994 9665 8035 9699
rect 8069 9665 8110 9699
rect 8144 9665 8185 9699
rect 8219 9665 8260 9699
rect 8294 9665 8335 9699
rect 8369 9665 8410 9699
rect 8444 9665 8485 9699
rect 8519 9665 8559 9699
rect 8593 9665 8633 9699
rect 8667 9665 8707 9699
rect 8741 9665 8781 9699
rect 8815 9665 8855 9699
rect 8889 9665 8929 9699
rect 8963 9665 9003 9699
rect 9037 9665 9077 9699
rect 9111 9665 9151 9699
rect 9185 9665 9197 9699
rect 7300 9659 9197 9665
rect 7300 9651 7362 9659
rect 7149 9644 7362 9651
tri 7362 9644 7377 9659 nw
tri 7853 9644 7868 9659 ne
rect 7868 9644 8062 9659
tri 8062 9644 8077 9659 nw
tri 8297 9644 8312 9659 ne
rect 8312 9644 8684 9659
tri 8684 9644 8699 9659 nw
tri 9027 9644 9042 9659 ne
rect 9042 9644 9197 9659
rect 7149 9635 7353 9644
tri 7353 9635 7362 9644 nw
tri 7868 9635 7877 9644 ne
rect 7877 9635 8053 9644
tri 8053 9635 8062 9644 nw
tri 8312 9635 8321 9644 ne
rect 8321 9635 8675 9644
tri 8675 9635 8684 9644 nw
tri 9042 9635 9051 9644 ne
rect 7149 9627 7329 9635
rect 7149 9593 7155 9627
rect 7189 9613 7329 9627
rect 7189 9593 7266 9613
rect 7149 9581 7266 9593
tri 7192 9579 7194 9581 ne
rect 7194 9579 7266 9581
rect 7300 9579 7329 9613
tri 7329 9611 7353 9635 nw
tri 7194 9548 7225 9579 ne
rect 7225 9548 7329 9579
tri 7225 9541 7232 9548 ne
rect 7232 9541 7329 9548
tri 7232 9536 7237 9541 ne
rect 7237 9507 7266 9541
rect 7300 9507 7329 9541
rect 7237 9469 7329 9507
rect 7237 9435 7266 9469
rect 7300 9435 7329 9469
rect 7237 9397 7329 9435
rect 7237 9363 7266 9397
rect 7300 9363 7329 9397
rect 7877 9582 8051 9635
tri 8051 9633 8053 9635 nw
rect 7877 9548 7883 9582
rect 7917 9548 8011 9582
rect 8045 9548 8051 9582
rect 7877 9510 8051 9548
rect 7877 9476 7883 9510
rect 7917 9476 8011 9510
rect 8045 9476 8051 9510
rect 8321 9592 8673 9635
tri 8673 9633 8675 9635 nw
rect 8321 9558 8333 9592
rect 8367 9558 8406 9592
rect 8440 9558 8479 9592
rect 8513 9558 8553 9592
rect 8587 9558 8627 9592
rect 8661 9558 8673 9592
rect 8321 9520 8673 9558
rect 8321 9486 8333 9520
rect 8367 9486 8406 9520
rect 8440 9486 8479 9520
rect 8513 9486 8553 9520
rect 8587 9486 8627 9520
rect 8661 9486 8673 9520
rect 8321 9480 8673 9486
rect 9051 9606 9197 9644
rect 10066 9678 10444 9717
rect 10066 9644 10072 9678
rect 10106 9644 10178 9678
rect 10212 9659 10444 9678
rect 10212 9646 10281 9659
tri 10281 9646 10294 9659 nw
rect 10212 9644 10267 9646
rect 10066 9632 10267 9644
tri 10267 9632 10281 9646 nw
tri 9197 9606 9223 9632 sw
rect 10066 9606 10241 9632
tri 10241 9606 10267 9632 nw
rect 9051 9605 9223 9606
tri 9223 9605 9224 9606 sw
rect 10066 9605 10218 9606
rect 9051 9604 9224 9605
tri 9224 9604 9225 9605 sw
rect 9051 9582 9225 9604
rect 9051 9548 9057 9582
rect 9091 9548 9185 9582
rect 9219 9548 9225 9582
rect 9051 9508 9225 9548
rect 7877 9438 8051 9476
rect 7877 9404 7883 9438
rect 7917 9404 8011 9438
rect 8045 9404 8051 9438
rect 7877 9392 8051 9404
rect 9051 9474 9057 9508
rect 9091 9474 9185 9508
rect 9219 9474 9225 9508
rect 9051 9434 9225 9474
rect 9051 9400 9057 9434
rect 9091 9400 9185 9434
rect 9219 9400 9225 9434
rect 10066 9571 10072 9605
rect 10106 9571 10178 9605
rect 10212 9571 10218 9605
tri 10218 9583 10241 9606 nw
rect 10066 9532 10218 9571
rect 10066 9498 10072 9532
rect 10106 9498 10178 9532
rect 10212 9498 10218 9532
rect 10066 9459 10218 9498
rect 10066 9425 10072 9459
rect 10106 9425 10178 9459
rect 10212 9425 10218 9459
rect 10066 9413 10218 9425
rect 9051 9388 9225 9400
rect 7237 9324 7329 9363
rect 7237 9290 7266 9324
rect 7300 9290 7329 9324
rect 6999 9250 7091 9262
rect 6999 9216 7028 9250
rect 7062 9216 7091 9250
rect 6999 9177 7091 9216
rect 6999 9143 7028 9177
rect 7062 9143 7091 9177
rect 6999 9103 7091 9143
rect 6999 9069 7028 9103
rect 7062 9069 7091 9103
rect 6999 9029 7091 9069
rect 6999 8995 7028 9029
rect 7062 8995 7091 9029
rect 6999 8955 7091 8995
rect 6999 8921 7028 8955
rect 7062 8921 7091 8955
rect 6999 8888 7091 8921
rect 6925 8876 7091 8888
rect 6925 8842 6931 8876
rect 6965 8842 7051 8876
rect 7085 8842 7091 8876
rect 6925 8792 7091 8842
rect 6925 8758 6931 8792
rect 6965 8758 7051 8792
rect 7085 8758 7091 8792
rect 6925 8708 7091 8758
rect 6925 8674 6931 8708
rect 6965 8674 7051 8708
rect 7085 8674 7091 8708
tri 6894 8633 6925 8664 se
rect 6925 8633 7091 8674
tri 6885 8624 6894 8633 se
rect 6894 8624 7091 8633
tri 6878 8617 6885 8624 se
rect 6885 8617 6931 8624
rect 6743 8590 6931 8617
rect 6965 8590 7051 8624
rect 7085 8590 7091 8624
rect 6743 8584 7091 8590
rect 6743 8550 6749 8584
rect 6783 8550 6851 8584
rect 6885 8550 7091 8584
rect 6743 8540 7091 8550
rect 6743 8506 6931 8540
rect 6965 8506 7051 8540
rect 7085 8506 7091 8540
rect 6743 8505 7091 8506
rect 6743 8471 6749 8505
rect 6783 8471 6851 8505
rect 6885 8493 7091 8505
rect 6885 8487 7085 8493
tri 7085 8487 7091 8493 nw
rect 7237 9251 7329 9290
rect 7237 9217 7266 9251
rect 7300 9217 7329 9251
rect 7237 9178 7329 9217
rect 7237 9144 7266 9178
rect 7300 9144 7329 9178
rect 7237 9105 7329 9144
rect 7237 9071 7266 9105
rect 7300 9071 7329 9105
rect 7237 9032 7329 9071
rect 7237 8998 7266 9032
rect 7300 8998 7329 9032
rect 7237 8959 7329 8998
rect 7237 8925 7266 8959
rect 7300 8925 7329 8959
rect 7237 8886 7329 8925
rect 7237 8852 7266 8886
rect 7300 8852 7329 8886
rect 7237 8813 7329 8852
rect 7237 8779 7266 8813
rect 7300 8779 7329 8813
rect 7237 8740 7329 8779
rect 7237 8706 7266 8740
rect 7300 8706 7329 8740
rect 7237 8667 7329 8706
rect 7237 8633 7266 8667
rect 7300 8633 7329 8667
rect 7237 8594 7329 8633
rect 27494 9319 27498 9860
rect 27806 9828 27974 9868
rect 27823 9794 27861 9828
rect 27895 9794 27974 9828
rect 27806 9754 27974 9794
rect 27823 9720 27861 9754
rect 27895 9720 27974 9754
rect 27806 9680 27974 9720
rect 27823 9646 27861 9680
rect 27895 9646 27974 9680
rect 27806 9606 27974 9646
rect 27823 9572 27861 9606
rect 27895 9572 27974 9606
rect 27806 9532 27974 9572
rect 27823 9498 27861 9532
rect 27895 9498 27974 9532
rect 27806 9458 27974 9498
rect 27823 9424 27861 9458
rect 27895 9424 27974 9458
rect 27806 9384 27974 9424
rect 27823 9350 27861 9384
rect 27895 9350 27974 9384
rect 27806 9319 27974 9350
rect 27494 9310 27974 9319
rect 27494 9306 27501 9310
rect 27535 9306 27573 9310
rect 27607 9306 27645 9310
rect 27679 9306 27717 9310
rect 27751 9306 27789 9310
rect 27494 9254 27498 9306
rect 27550 9254 27562 9306
rect 27614 9254 27626 9306
rect 27679 9276 27690 9306
rect 27751 9276 27754 9306
rect 27823 9276 27861 9310
rect 27895 9276 27974 9310
rect 27678 9254 27690 9276
rect 27742 9254 27754 9276
rect 27806 9254 27974 9276
rect 27494 9241 27974 9254
rect 27494 9189 27498 9241
rect 27550 9189 27562 9241
rect 27614 9189 27626 9241
rect 27678 9236 27690 9241
rect 27742 9236 27754 9241
rect 27806 9236 27974 9241
rect 27679 9202 27690 9236
rect 27751 9202 27754 9236
rect 27823 9202 27861 9236
rect 27895 9202 27974 9236
rect 27678 9189 27690 9202
rect 27742 9189 27754 9202
rect 27806 9189 27974 9202
rect 27494 9176 27974 9189
rect 27494 9124 27498 9176
rect 27550 9124 27562 9176
rect 27614 9124 27626 9176
rect 27678 9162 27690 9176
rect 27742 9162 27754 9176
rect 27806 9162 27974 9176
rect 27679 9128 27690 9162
rect 27751 9128 27754 9162
rect 27823 9128 27861 9162
rect 27895 9128 27974 9162
rect 27678 9124 27690 9128
rect 27742 9124 27754 9128
rect 27806 9124 27974 9128
rect 27494 9111 27974 9124
rect 27494 9059 27498 9111
rect 27550 9059 27562 9111
rect 27614 9059 27626 9111
rect 27678 9088 27690 9111
rect 27742 9088 27754 9111
rect 27806 9088 27974 9111
rect 27679 9059 27690 9088
rect 27751 9059 27754 9088
rect 27494 9054 27501 9059
rect 27535 9054 27573 9059
rect 27607 9054 27645 9059
rect 27679 9054 27717 9059
rect 27751 9054 27789 9059
rect 27823 9054 27861 9088
rect 27895 9054 27974 9088
rect 27494 9046 27974 9054
rect 27494 8994 27498 9046
rect 27550 8994 27562 9046
rect 27614 8994 27626 9046
rect 27678 9014 27690 9046
rect 27742 9014 27754 9046
rect 27806 9014 27974 9046
rect 27679 8994 27690 9014
rect 27751 8994 27754 9014
rect 27494 8981 27501 8994
rect 27535 8981 27573 8994
rect 27607 8981 27645 8994
rect 27679 8981 27717 8994
rect 27751 8981 27789 8994
rect 27494 8929 27498 8981
rect 27550 8929 27562 8981
rect 27614 8929 27626 8981
rect 27679 8980 27690 8981
rect 27751 8980 27754 8981
rect 27823 8980 27861 9014
rect 27895 8980 27974 9014
rect 27678 8940 27690 8980
rect 27742 8940 27754 8980
rect 27806 8940 27974 8980
rect 27679 8929 27690 8940
rect 27751 8929 27754 8940
rect 27494 8916 27501 8929
rect 27535 8916 27573 8929
rect 27607 8916 27645 8929
rect 27679 8916 27717 8929
rect 27751 8916 27789 8929
rect 27494 8864 27498 8916
rect 27550 8864 27562 8916
rect 27614 8864 27626 8916
rect 27679 8906 27690 8916
rect 27751 8906 27754 8916
rect 27823 8906 27861 8940
rect 27895 8906 27974 8940
rect 27678 8866 27690 8906
rect 27742 8866 27754 8906
rect 27806 8866 27974 8906
rect 27679 8864 27690 8866
rect 27751 8864 27754 8866
rect 27494 8851 27501 8864
rect 27535 8851 27573 8864
rect 27607 8851 27645 8864
rect 27679 8851 27717 8864
rect 27751 8851 27789 8864
rect 27494 8799 27498 8851
rect 27550 8799 27562 8851
rect 27614 8799 27626 8851
rect 27679 8832 27690 8851
rect 27751 8832 27754 8851
rect 27823 8832 27861 8866
rect 27895 8832 27974 8866
rect 27678 8799 27690 8832
rect 27742 8799 27754 8832
rect 27806 8799 27974 8832
rect 27494 8792 27974 8799
rect 27494 8786 27501 8792
rect 27535 8786 27573 8792
rect 27607 8786 27645 8792
rect 27679 8786 27717 8792
rect 27751 8786 27789 8792
rect 27494 8734 27498 8786
rect 27550 8734 27562 8786
rect 27614 8734 27626 8786
rect 27679 8758 27690 8786
rect 27751 8758 27754 8786
rect 27823 8758 27861 8792
rect 27895 8758 27974 8792
rect 27678 8734 27690 8758
rect 27742 8734 27754 8758
rect 27806 8734 27974 8758
rect 27494 8721 27974 8734
rect 27494 8669 27498 8721
rect 27550 8669 27562 8721
rect 27614 8669 27626 8721
rect 27678 8718 27690 8721
rect 27742 8718 27754 8721
rect 27806 8718 27974 8721
rect 27679 8684 27690 8718
rect 27751 8684 27754 8718
rect 27823 8684 27861 8718
rect 27895 8684 27974 8718
rect 27678 8669 27690 8684
rect 27742 8669 27754 8684
rect 27806 8669 27974 8684
rect 27494 8656 27974 8669
rect 27494 8604 27498 8656
rect 27550 8604 27562 8656
rect 27614 8604 27626 8656
rect 27678 8644 27690 8656
rect 27742 8644 27754 8656
rect 27806 8644 27974 8656
rect 27679 8610 27690 8644
rect 27751 8610 27754 8644
rect 27823 8610 27861 8644
rect 27895 8610 27974 8644
rect 27678 8604 27690 8610
rect 27742 8604 27754 8610
rect 27806 8604 27974 8610
rect 27494 8594 27974 8604
rect 7237 8560 7266 8594
rect 7300 8560 7329 8594
rect 7237 8521 7329 8560
rect 7237 8487 7266 8521
rect 7300 8487 7329 8521
rect 6885 8471 7046 8487
rect 6743 8448 7046 8471
tri 7046 8448 7085 8487 nw
rect 7237 8448 7329 8487
rect 6743 8426 7012 8448
rect 6743 8392 6749 8426
rect 6783 8392 6851 8426
rect 6885 8414 7012 8426
tri 7012 8414 7046 8448 nw
rect 7237 8414 7266 8448
rect 7300 8414 7329 8448
rect 6885 8395 6993 8414
tri 6993 8395 7012 8414 nw
rect 6885 8392 6979 8395
rect 6743 8347 6979 8392
tri 6979 8381 6993 8395 nw
rect 6743 8313 6749 8347
rect 6783 8313 6851 8347
rect 6885 8313 6979 8347
tri 672 8268 679 8275 se
rect 679 8268 945 8275
tri 639 8235 672 8268 se
rect 672 8235 945 8268
tri 616 8212 639 8235 se
rect 639 8212 945 8235
tri 582 8178 616 8212 se
rect 616 8178 945 8212
tri 559 8155 582 8178 se
rect 582 8155 945 8178
tri 539 8135 559 8155 se
rect 559 8135 945 8155
rect 6743 8268 6979 8313
rect 7237 8375 7329 8414
rect 27828 8407 27974 8594
rect 7237 8341 7266 8375
rect 7300 8341 7329 8375
rect 27266 8395 27974 8407
rect 27266 8361 27272 8395
rect 27306 8361 27344 8395
rect 27378 8361 27416 8395
rect 27450 8361 27488 8395
rect 27522 8361 27560 8395
rect 27594 8361 27632 8395
rect 27666 8361 27704 8395
rect 27738 8361 27776 8395
rect 27810 8361 27848 8395
rect 27882 8361 27920 8395
rect 27954 8361 27974 8395
rect 7237 8302 7329 8341
tri 6979 8268 6985 8274 sw
rect 7237 8268 7266 8302
rect 7300 8268 7329 8302
rect 15697 8336 16622 8342
rect 15697 8302 15709 8336
rect 15743 8302 15782 8336
rect 15816 8302 15855 8336
rect 15889 8302 15928 8336
rect 15962 8302 16000 8336
rect 16034 8302 16072 8336
rect 16106 8302 16144 8336
rect 16178 8302 16216 8336
rect 16250 8302 16288 8336
rect 16322 8302 16360 8336
rect 16394 8302 16432 8336
rect 16466 8302 16504 8336
rect 16538 8302 16576 8336
rect 16610 8302 16622 8336
rect 15697 8296 16622 8302
rect 27266 8315 27974 8361
rect 6743 8262 6985 8268
tri 6985 8262 6991 8268 sw
rect 6743 8256 6991 8262
tri 6991 8256 6997 8262 sw
tri 7231 8256 7237 8262 se
rect 7237 8256 7329 8268
rect 6743 8235 6997 8256
tri 6997 8235 7018 8256 sw
tri 7210 8235 7231 8256 se
rect 7231 8235 7329 8256
rect 6743 8224 7018 8235
tri 7018 8224 7029 8235 sw
tri 7199 8224 7210 8235 se
rect 7210 8224 7329 8235
rect 6743 8212 7329 8224
rect 6743 8178 7091 8212
rect 7125 8178 7205 8212
rect 7239 8178 7329 8212
rect 6743 8135 7329 8178
rect 27266 8281 27272 8315
rect 27306 8281 27344 8315
rect 27378 8281 27416 8315
rect 27450 8281 27488 8315
rect 27522 8281 27560 8315
rect 27594 8281 27632 8315
rect 27666 8281 27704 8315
rect 27738 8281 27776 8315
rect 27810 8281 27848 8315
rect 27882 8281 27920 8315
rect 27954 8281 27974 8315
rect 27266 8235 27974 8281
rect 27266 8201 27272 8235
rect 27306 8201 27344 8235
rect 27378 8201 27416 8235
rect 27450 8201 27488 8235
rect 27522 8201 27560 8235
rect 27594 8201 27632 8235
rect 27666 8201 27704 8235
rect 27738 8201 27776 8235
rect 27810 8201 27848 8235
rect 27882 8201 27920 8235
rect 27954 8201 27974 8235
rect 27266 8155 27974 8201
tri 525 8121 539 8135 se
rect 539 8121 945 8135
tri 484 8080 525 8121 se
rect 525 8080 945 8121
rect 166 8068 945 8080
rect 166 8034 179 8068
rect 213 8034 257 8068
rect 291 8034 335 8068
rect 369 8034 413 8068
rect 447 8034 491 8068
rect 525 8034 569 8068
rect 603 8034 647 8068
rect 681 8034 725 8068
rect 759 8034 803 8068
rect 837 8034 945 8068
rect 7085 8080 7245 8135
rect 7085 8046 7091 8080
rect 7125 8046 7205 8080
rect 7239 8046 7245 8080
rect 7085 8034 7245 8046
rect 27266 8121 27272 8155
rect 27306 8121 27344 8155
rect 27378 8121 27416 8155
rect 27450 8121 27488 8155
rect 27522 8121 27560 8155
rect 27594 8121 27632 8155
rect 27666 8121 27704 8155
rect 27738 8121 27776 8155
rect 27810 8121 27848 8155
rect 27882 8121 27920 8155
rect 27954 8121 27974 8155
rect 27266 8074 27974 8121
rect 27266 8040 27272 8074
rect 27306 8040 27344 8074
rect 27378 8040 27416 8074
rect 27450 8040 27488 8074
rect 27522 8040 27560 8074
rect 27594 8040 27632 8074
rect 27666 8040 27704 8074
rect 27738 8040 27776 8074
rect 27810 8040 27848 8074
rect 27882 8040 27920 8074
rect 27954 8040 27974 8074
rect 166 7996 945 8034
rect 166 7962 179 7996
rect 213 7962 257 7996
rect 291 7962 335 7996
rect 369 7962 413 7996
rect 447 7962 491 7996
rect 525 7962 569 7996
rect 603 7962 647 7996
rect 681 7962 725 7996
rect 759 7962 803 7996
rect 837 7962 945 7996
rect 166 7924 945 7962
rect 166 7890 179 7924
rect 213 7890 257 7924
rect 291 7890 335 7924
rect 369 7890 413 7924
rect 447 7890 491 7924
rect 525 7890 569 7924
rect 603 7890 647 7924
rect 681 7890 725 7924
rect 759 7890 803 7924
rect 837 7890 945 7924
rect 166 7852 945 7890
rect 166 7818 179 7852
rect 213 7818 257 7852
rect 291 7818 335 7852
rect 369 7818 413 7852
rect 447 7818 491 7852
rect 525 7818 569 7852
rect 603 7818 647 7852
rect 681 7818 725 7852
rect 759 7818 803 7852
rect 837 7827 945 7852
rect 27266 7993 27974 8040
rect 27266 7959 27272 7993
rect 27306 7959 27344 7993
rect 27378 7959 27416 7993
rect 27450 7959 27488 7993
rect 27522 7959 27560 7993
rect 27594 7959 27632 7993
rect 27666 7959 27704 7993
rect 27738 7959 27776 7993
rect 27810 7959 27848 7993
rect 27882 7959 27920 7993
rect 27954 7959 27974 7993
rect 27266 7912 27974 7959
rect 27266 7878 27272 7912
rect 27306 7878 27344 7912
rect 27378 7878 27416 7912
rect 27450 7878 27488 7912
rect 27522 7878 27560 7912
rect 27594 7878 27632 7912
rect 27666 7878 27704 7912
rect 27738 7878 27776 7912
rect 27810 7878 27848 7912
rect 27882 7878 27920 7912
rect 27954 7878 27974 7912
rect 27266 7831 27974 7878
rect 837 7818 961 7827
rect 166 7797 961 7818
tri 961 7797 991 7827 nw
rect 27266 7797 27272 7831
rect 27306 7797 27344 7831
rect 27378 7797 27416 7831
rect 27450 7797 27488 7831
rect 27522 7797 27560 7831
rect 27594 7797 27632 7831
rect 27666 7797 27704 7831
rect 27738 7797 27776 7831
rect 27810 7797 27848 7831
rect 27882 7797 27920 7831
rect 27954 7797 27974 7831
rect 166 7780 914 7797
rect 166 7746 179 7780
rect 213 7746 257 7780
rect 291 7746 335 7780
rect 369 7746 413 7780
rect 447 7746 491 7780
rect 525 7746 569 7780
rect 603 7746 647 7780
rect 681 7746 725 7780
rect 759 7746 803 7780
rect 837 7750 914 7780
tri 914 7750 961 7797 nw
rect 27266 7750 27974 7797
rect 837 7746 880 7750
rect 166 7716 880 7746
tri 880 7716 914 7750 nw
rect 27266 7716 27272 7750
rect 27306 7716 27344 7750
rect 27378 7716 27416 7750
rect 27450 7716 27488 7750
rect 27522 7716 27560 7750
rect 27594 7716 27632 7750
rect 27666 7716 27704 7750
rect 27738 7716 27776 7750
rect 27810 7716 27848 7750
rect 27882 7716 27920 7750
rect 27954 7716 27974 7750
rect 166 7707 868 7716
rect 166 7673 179 7707
rect 213 7673 257 7707
rect 291 7673 335 7707
rect 369 7673 413 7707
rect 447 7673 491 7707
rect 525 7673 569 7707
rect 603 7673 647 7707
rect 681 7673 725 7707
rect 759 7673 803 7707
rect 837 7704 868 7707
tri 868 7704 880 7716 nw
rect 27266 7704 27974 7716
rect 837 7673 850 7704
tri 850 7686 868 7704 nw
rect 166 7634 850 7673
rect 166 7600 179 7634
rect 213 7600 257 7634
rect 291 7600 335 7634
rect 369 7600 413 7634
rect 447 7600 491 7634
rect 525 7600 569 7634
rect 603 7600 647 7634
rect 681 7600 725 7634
rect 759 7600 803 7634
rect 837 7600 850 7634
rect 166 7561 850 7600
rect 166 7527 179 7561
rect 213 7527 257 7561
rect 291 7527 335 7561
rect 369 7527 413 7561
rect 447 7527 491 7561
rect 525 7527 569 7561
rect 603 7527 647 7561
rect 681 7527 725 7561
rect 759 7527 803 7561
rect 837 7527 850 7561
rect 166 7488 850 7527
rect 166 7454 179 7488
rect 213 7454 257 7488
rect 291 7454 335 7488
rect 369 7454 413 7488
rect 447 7454 491 7488
rect 525 7454 569 7488
rect 603 7454 647 7488
rect 681 7454 725 7488
rect 759 7454 803 7488
rect 837 7454 850 7488
rect 166 7415 850 7454
rect 166 7381 179 7415
rect 213 7381 257 7415
rect 291 7381 335 7415
rect 369 7381 413 7415
rect 447 7381 491 7415
rect 525 7381 569 7415
rect 603 7381 647 7415
rect 681 7381 725 7415
rect 759 7381 803 7415
rect 837 7381 850 7415
rect 166 7342 850 7381
rect 166 7308 179 7342
rect 213 7308 257 7342
rect 291 7308 335 7342
rect 369 7308 413 7342
rect 447 7308 491 7342
rect 525 7308 569 7342
rect 603 7308 647 7342
rect 681 7308 725 7342
rect 759 7308 803 7342
rect 837 7308 850 7342
rect 166 7269 850 7308
rect 166 7235 179 7269
rect 213 7235 257 7269
rect 291 7235 335 7269
rect 369 7235 413 7269
rect 447 7235 491 7269
rect 525 7235 569 7269
rect 603 7235 647 7269
rect 681 7235 725 7269
rect 759 7235 803 7269
rect 837 7235 850 7269
rect 166 7196 850 7235
rect 166 7162 179 7196
rect 213 7162 257 7196
rect 291 7162 335 7196
rect 369 7162 413 7196
rect 447 7162 491 7196
rect 525 7162 569 7196
rect 603 7162 647 7196
rect 681 7162 725 7196
rect 759 7162 803 7196
rect 837 7162 850 7196
rect 166 7123 850 7162
rect 166 7089 179 7123
rect 213 7089 257 7123
rect 291 7089 335 7123
rect 369 7089 413 7123
rect 447 7089 491 7123
rect 525 7089 569 7123
rect 603 7089 647 7123
rect 681 7089 725 7123
rect 759 7089 803 7123
rect 837 7089 850 7123
rect 166 7050 850 7089
rect 166 7016 179 7050
rect 213 7016 257 7050
rect 291 7016 335 7050
rect 369 7016 413 7050
rect 447 7016 491 7050
rect 525 7016 569 7050
rect 603 7016 647 7050
rect 681 7016 725 7050
rect 759 7016 803 7050
rect 837 7016 850 7050
rect 166 6977 850 7016
rect 166 6943 179 6977
rect 213 6943 257 6977
rect 291 6943 335 6977
rect 369 6943 413 6977
rect 447 6943 491 6977
rect 525 6943 569 6977
rect 603 6943 647 6977
rect 681 6943 725 6977
rect 759 6943 803 6977
rect 837 6943 850 6977
rect 166 6904 850 6943
rect 166 6870 179 6904
rect 213 6870 257 6904
rect 291 6870 335 6904
rect 369 6870 413 6904
rect 447 6870 491 6904
rect 525 6870 569 6904
rect 603 6870 647 6904
rect 681 6870 725 6904
rect 759 6870 803 6904
rect 837 6870 850 6904
rect 166 6831 850 6870
rect 13555 7296 13956 7302
rect 13555 7244 13565 7296
rect 13617 7244 13631 7296
rect 13683 7244 13697 7296
rect 13749 7244 13763 7296
rect 13815 7244 13828 7296
rect 13880 7244 13893 7296
rect 13945 7244 13956 7296
rect 13555 7210 13956 7244
rect 13555 7158 13565 7210
rect 13617 7158 13631 7210
rect 13683 7158 13697 7210
rect 13749 7158 13763 7210
rect 13815 7158 13828 7210
rect 13880 7158 13893 7210
rect 13945 7158 13956 7210
rect 13555 6837 13956 7158
rect 14877 7298 15086 7299
rect 14877 7246 14883 7298
rect 14935 7246 14956 7298
rect 15008 7246 15028 7298
rect 15080 7246 15086 7298
rect 14877 7210 15086 7246
rect 14877 7158 14883 7210
rect 14935 7158 14956 7210
rect 15008 7158 15028 7210
rect 15080 7158 15086 7210
rect 14877 7070 15086 7158
rect 14257 7058 14447 7070
rect 166 6797 179 6831
rect 213 6797 257 6831
rect 291 6797 335 6831
rect 369 6797 413 6831
rect 447 6797 491 6831
rect 525 6797 569 6831
rect 603 6797 647 6831
rect 681 6797 725 6831
rect 759 6797 803 6831
rect 837 6797 850 6831
rect 166 6758 850 6797
rect 166 6724 179 6758
rect 213 6724 257 6758
rect 291 6724 335 6758
rect 369 6724 413 6758
rect 447 6724 491 6758
rect 525 6724 569 6758
rect 603 6724 647 6758
rect 681 6724 725 6758
rect 759 6724 803 6758
rect 837 6724 850 6758
rect 166 6685 850 6724
rect 166 6651 179 6685
rect 213 6651 257 6685
rect 291 6651 335 6685
rect 369 6651 413 6685
rect 447 6651 491 6685
rect 525 6651 569 6685
rect 603 6651 647 6685
rect 681 6651 725 6685
rect 759 6651 803 6685
rect 837 6651 850 6685
rect 166 6612 850 6651
rect 166 6578 179 6612
rect 213 6578 257 6612
rect 291 6578 335 6612
rect 369 6578 413 6612
rect 447 6578 491 6612
rect 525 6578 569 6612
rect 603 6578 647 6612
rect 681 6578 725 6612
rect 759 6578 803 6612
rect 837 6578 850 6612
rect 166 6539 850 6578
rect 166 6505 179 6539
rect 213 6505 257 6539
rect 291 6505 335 6539
rect 369 6505 413 6539
rect 447 6505 491 6539
rect 525 6505 569 6539
rect 603 6505 647 6539
rect 681 6505 725 6539
rect 759 6505 803 6539
rect 837 6505 850 6539
rect 166 6466 850 6505
rect 166 6432 179 6466
rect 213 6432 257 6466
rect 291 6432 335 6466
rect 369 6432 413 6466
rect 447 6432 491 6466
rect 525 6432 569 6466
rect 603 6432 647 6466
rect 681 6432 725 6466
rect 759 6432 803 6466
rect 837 6432 850 6466
rect 166 6393 850 6432
rect 166 6359 179 6393
rect 213 6359 257 6393
rect 291 6359 335 6393
rect 369 6359 413 6393
rect 447 6359 491 6393
rect 525 6359 569 6393
rect 603 6359 647 6393
rect 681 6359 725 6393
rect 759 6359 803 6393
rect 837 6359 850 6393
rect 166 6320 850 6359
rect 166 6286 179 6320
rect 213 6286 257 6320
rect 291 6286 335 6320
rect 369 6286 413 6320
rect 447 6286 491 6320
rect 525 6286 569 6320
rect 603 6286 647 6320
rect 681 6286 725 6320
rect 759 6286 803 6320
rect 837 6286 850 6320
rect 13175 6828 13958 6837
rect 13175 6794 13187 6828
rect 13221 6794 13260 6828
rect 13294 6794 13333 6828
rect 13367 6794 13406 6828
rect 13440 6794 13479 6828
rect 13513 6794 13552 6828
rect 13586 6794 13624 6828
rect 13658 6794 13696 6828
rect 13730 6794 13768 6828
rect 13802 6794 13840 6828
rect 13874 6794 13912 6828
rect 13946 6794 13958 6828
rect 13175 6750 13958 6794
rect 13175 6716 13187 6750
rect 13221 6716 13260 6750
rect 13294 6716 13333 6750
rect 13367 6716 13406 6750
rect 13440 6716 13479 6750
rect 13513 6716 13552 6750
rect 13586 6716 13624 6750
rect 13658 6716 13696 6750
rect 13730 6716 13768 6750
rect 13802 6716 13840 6750
rect 13874 6716 13912 6750
rect 13946 6716 13958 6750
rect 13175 6672 13958 6716
rect 13175 6638 13187 6672
rect 13221 6638 13260 6672
rect 13294 6638 13333 6672
rect 13367 6638 13406 6672
rect 13440 6638 13479 6672
rect 13513 6638 13552 6672
rect 13586 6638 13624 6672
rect 13658 6638 13696 6672
rect 13730 6638 13768 6672
rect 13802 6638 13840 6672
rect 13874 6638 13912 6672
rect 13946 6638 13958 6672
rect 13175 6594 13958 6638
rect 13175 6560 13187 6594
rect 13221 6560 13260 6594
rect 13294 6560 13333 6594
rect 13367 6560 13406 6594
rect 13440 6560 13479 6594
rect 13513 6560 13552 6594
rect 13586 6560 13624 6594
rect 13658 6560 13696 6594
rect 13730 6560 13768 6594
rect 13802 6560 13840 6594
rect 13874 6560 13912 6594
rect 13946 6560 13958 6594
rect 13175 6516 13958 6560
rect 13175 6482 13187 6516
rect 13221 6482 13260 6516
rect 13294 6482 13333 6516
rect 13367 6482 13406 6516
rect 13440 6482 13479 6516
rect 13513 6482 13552 6516
rect 13586 6482 13624 6516
rect 13658 6482 13696 6516
rect 13730 6482 13768 6516
rect 13802 6482 13840 6516
rect 13874 6482 13912 6516
rect 13946 6482 13958 6516
rect 13175 6438 13958 6482
rect 13175 6404 13187 6438
rect 13221 6404 13260 6438
rect 13294 6404 13333 6438
rect 13367 6404 13406 6438
rect 13440 6404 13479 6438
rect 13513 6404 13552 6438
rect 13586 6404 13624 6438
rect 13658 6404 13696 6438
rect 13730 6404 13768 6438
rect 13802 6404 13840 6438
rect 13874 6404 13912 6438
rect 13946 6404 13958 6438
rect 13175 6360 13958 6404
rect 13175 6326 13187 6360
rect 13221 6326 13260 6360
rect 13294 6326 13333 6360
rect 13367 6326 13406 6360
rect 13440 6326 13479 6360
rect 13513 6326 13552 6360
rect 13586 6326 13624 6360
rect 13658 6326 13696 6360
rect 13730 6326 13768 6360
rect 13802 6326 13840 6360
rect 13874 6326 13912 6360
rect 13946 6326 13958 6360
rect 13175 6317 13958 6326
rect 166 6247 850 6286
rect 166 6213 179 6247
rect 213 6213 257 6247
rect 291 6213 335 6247
rect 369 6213 413 6247
rect 447 6213 491 6247
rect 525 6213 569 6247
rect 603 6213 647 6247
rect 681 6213 725 6247
rect 759 6213 803 6247
rect 837 6213 850 6247
rect 13569 6282 13958 6317
rect 14257 6448 14263 7058
rect 14441 6448 14447 7058
rect 14257 6409 14447 6448
rect 14257 6375 14263 6409
rect 14297 6375 14335 6409
rect 14369 6375 14407 6409
rect 14441 6375 14447 6409
rect 14257 6350 14447 6375
rect 14757 7058 15091 7070
rect 14757 6448 14763 7058
rect 15085 6448 15091 7058
rect 14757 6409 15091 6448
rect 14757 6375 14763 6409
rect 14797 6375 14835 6409
rect 14869 6375 14907 6409
rect 14941 6375 14979 6409
rect 15013 6375 15051 6409
rect 15085 6375 15091 6409
rect 14757 6350 15091 6375
rect 14257 6336 15091 6350
rect 14257 6302 14263 6336
rect 14297 6302 14335 6336
rect 14369 6302 14407 6336
rect 14441 6302 14763 6336
rect 14797 6302 14835 6336
rect 14869 6302 14907 6336
rect 14941 6302 14979 6336
rect 15013 6302 15051 6336
rect 15085 6302 15091 6336
rect 14257 6290 15091 6302
rect 14257 6282 15086 6290
rect 13569 6224 15086 6282
rect 166 6166 850 6213
rect 166 5124 173 6166
rect 351 5930 850 6166
rect 351 5124 359 5930
tri 359 5829 460 5930 nw
rect 166 5085 359 5124
tri 141 5051 166 5076 se
rect 166 5051 173 5085
rect 207 5051 245 5085
rect 279 5051 317 5085
rect 351 5051 359 5085
tri 102 5012 141 5051 se
rect 141 5012 359 5051
tri 83 4993 102 5012 se
rect 102 4993 173 5012
rect 83 4978 173 4993
rect 207 4978 245 5012
rect 279 4978 317 5012
rect 351 4978 359 5012
rect 83 4964 359 4978
rect 83 4391 148 4964
tri 148 4753 359 4964 nw
tri 148 4391 166 4409 sw
rect 83 4343 166 4391
tri 83 4260 166 4343 ne
tri 166 4260 297 4391 sw
rect 2103 4320 2239 4326
rect 2155 4268 2187 4320
rect 166 4247 297 4260
tri 297 4247 310 4260 sw
rect 2103 4252 2239 4268
rect 166 4146 1143 4247
rect 166 4112 176 4146
rect 210 4112 254 4146
rect 288 4119 1143 4146
rect 2155 4200 2187 4252
rect 2103 4183 2239 4200
rect 2155 4131 2187 4183
rect 2103 4125 2239 4131
rect 288 4118 1046 4119
rect 288 4112 309 4118
rect 166 4074 309 4112
rect 166 4040 176 4074
rect 210 4040 254 4074
rect 288 4040 309 4074
rect 166 4002 309 4040
rect 166 3968 176 4002
rect 210 3968 254 4002
rect 288 3968 309 4002
tri 309 3986 441 4118 nw
rect 166 3930 309 3968
rect 166 3896 176 3930
rect 210 3896 254 3930
rect 288 3896 309 3930
rect 166 3858 309 3896
rect 166 3824 176 3858
rect 210 3824 254 3858
rect 288 3824 309 3858
rect 166 3786 309 3824
rect 166 3752 176 3786
rect 210 3752 254 3786
rect 288 3752 309 3786
rect 166 3714 309 3752
rect 166 3680 176 3714
rect 210 3680 254 3714
rect 288 3680 309 3714
rect 166 3642 309 3680
rect 166 3608 176 3642
rect 210 3608 254 3642
rect 288 3608 309 3642
rect 166 3570 309 3608
rect 166 3536 176 3570
rect 210 3536 254 3570
rect 288 3536 309 3570
rect 166 3497 309 3536
rect 166 3463 176 3497
rect 210 3463 254 3497
rect 288 3463 309 3497
rect 166 3424 309 3463
rect 1344 3638 2239 3644
rect 1344 3637 2103 3638
rect 1344 3603 1356 3637
rect 1390 3603 1436 3637
rect 1470 3603 1516 3637
rect 1550 3603 1596 3637
rect 1630 3603 1676 3637
rect 1710 3603 1755 3637
rect 1789 3603 1834 3637
rect 1868 3603 1913 3637
rect 1947 3603 1992 3637
rect 2026 3603 2071 3637
rect 1344 3586 2103 3603
rect 2155 3586 2187 3638
rect 1344 3570 2239 3586
rect 1344 3561 2103 3570
rect 1344 3527 1356 3561
rect 1390 3527 1436 3561
rect 1470 3527 1516 3561
rect 1550 3527 1596 3561
rect 1630 3527 1676 3561
rect 1710 3527 1755 3561
rect 1789 3527 1834 3561
rect 1868 3527 1913 3561
rect 1947 3527 1992 3561
rect 2026 3527 2071 3561
rect 1344 3518 2103 3527
rect 2155 3518 2187 3570
rect 1344 3502 2239 3518
rect 1344 3485 2103 3502
rect 1344 3451 1356 3485
rect 1390 3451 1436 3485
rect 1470 3451 1516 3485
rect 1550 3451 1596 3485
rect 1630 3451 1676 3485
rect 1710 3451 1755 3485
rect 1789 3451 1834 3485
rect 1868 3451 1913 3485
rect 1947 3451 1992 3485
rect 2026 3451 2071 3485
rect 1344 3450 2103 3451
rect 2155 3450 2187 3502
rect 1344 3444 2239 3450
rect 166 3390 176 3424
rect 210 3390 254 3424
rect 288 3390 309 3424
rect 166 3351 309 3390
rect 166 3317 176 3351
rect 210 3317 254 3351
rect 288 3317 309 3351
rect 166 3278 309 3317
rect 166 3244 176 3278
rect 210 3244 254 3278
rect 288 3244 309 3278
rect 166 3205 309 3244
rect 166 3171 176 3205
rect 210 3171 254 3205
rect 288 3171 309 3205
rect 166 3132 309 3171
rect 166 3098 176 3132
rect 210 3098 254 3132
rect 288 3098 309 3132
rect 166 3059 309 3098
rect 166 3025 176 3059
rect 210 3025 254 3059
rect 288 3025 309 3059
rect 26768 3197 26774 3249
rect 26826 3197 26849 3249
rect 26901 3197 26924 3249
rect 26976 3197 26998 3249
rect 27050 3197 27072 3249
rect 27124 3197 27146 3249
rect 27198 3197 27204 3249
rect 26768 3173 27204 3197
rect 26768 3121 26774 3173
rect 26826 3121 26849 3173
rect 26901 3121 26924 3173
rect 26976 3121 26998 3173
rect 27050 3121 27072 3173
rect 27124 3121 27146 3173
rect 27198 3121 27204 3173
rect 26768 3097 27204 3121
rect 26768 3045 26774 3097
rect 26826 3045 26849 3097
rect 26901 3045 26924 3097
rect 26976 3045 26998 3097
rect 27050 3045 27072 3097
rect 27124 3045 27146 3097
rect 27198 3045 27204 3097
rect 166 3006 309 3025
rect 2688 3011 3136 3018
rect 166 3000 1072 3006
rect 166 2986 341 3000
rect 166 2952 176 2986
rect 210 2952 254 2986
rect 288 2966 341 2986
rect 375 2966 415 3000
rect 449 2966 489 3000
rect 523 2966 563 3000
rect 597 2966 637 3000
rect 671 2966 711 3000
rect 745 2966 785 3000
rect 819 2966 859 3000
rect 893 2966 933 3000
rect 967 2966 1006 3000
rect 1040 2966 1072 3000
rect 288 2952 1072 2966
rect 166 2934 1072 2952
tri 167 2901 200 2934 ne
rect 200 2901 1072 2934
tri 200 2866 235 2901 ne
rect 235 2866 1072 2901
tri 235 2832 269 2866 ne
rect 269 2832 341 2866
rect 375 2832 415 2866
rect 449 2832 489 2866
rect 523 2832 563 2866
rect 597 2832 637 2866
rect 671 2832 711 2866
rect 745 2832 785 2866
rect 819 2832 859 2866
rect 893 2832 933 2866
rect 967 2832 1006 2866
rect 1040 2832 1072 2866
tri 269 2826 275 2832 ne
rect 275 2826 1072 2832
rect 2688 2977 2700 3011
rect 2734 2977 2778 3011
rect 2812 2977 2856 3011
rect 2890 2977 2934 3011
rect 2968 2977 3012 3011
rect 3046 2977 3090 3011
rect 3124 2977 3136 3011
rect 2688 2935 3136 2977
rect 2688 2901 2700 2935
rect 2734 2901 2778 2935
rect 2812 2901 2856 2935
rect 2890 2901 2934 2935
rect 2968 2901 3012 2935
rect 3046 2901 3090 2935
rect 3124 2901 3136 2935
rect 2688 2859 3136 2901
rect 2688 2825 2700 2859
rect 2734 2825 2778 2859
rect 2812 2825 2856 2859
rect 2890 2825 2934 2859
rect 2968 2825 3012 2859
rect 3046 2825 3090 2859
rect 3124 2825 3136 2859
rect 2688 2783 3136 2825
rect 2688 2749 2700 2783
rect 2734 2749 2778 2783
rect 2812 2749 2856 2783
rect 2890 2749 2934 2783
rect 2968 2749 3012 2783
rect 3046 2749 3090 2783
rect 3124 2749 3136 2783
tri 2638 2692 2688 2742 se
rect 2688 2692 3136 2749
rect 1946 2686 3136 2692
rect 1946 2652 1958 2686
rect 1992 2652 2034 2686
rect 2068 2652 2103 2686
rect 2155 2652 2186 2686
rect 2239 2652 2262 2686
rect 2296 2652 2338 2686
rect 2372 2652 2414 2686
rect 2448 2652 2490 2686
rect 2524 2652 2565 2686
rect 2599 2652 2640 2686
rect 2674 2652 2715 2686
rect 2749 2652 2790 2686
rect 2824 2652 2865 2686
rect 2899 2652 2940 2686
rect 2974 2652 3015 2686
rect 3049 2652 3090 2686
rect 3124 2652 3136 2686
rect 1946 2634 2103 2652
rect 2155 2634 2187 2652
rect 2239 2634 3136 2652
rect 1946 2594 3136 2634
rect 1946 2576 2103 2594
rect 2155 2576 2187 2594
rect 2239 2576 3136 2594
rect 1946 2542 1958 2576
rect 1992 2542 2034 2576
rect 2068 2542 2103 2576
rect 2155 2542 2186 2576
rect 2239 2542 2262 2576
rect 2296 2542 2338 2576
rect 2372 2542 2414 2576
rect 2448 2542 2490 2576
rect 2524 2542 2565 2576
rect 2599 2542 2640 2576
rect 2674 2542 2715 2576
rect 2749 2542 2790 2576
rect 2824 2542 2865 2576
rect 2899 2542 2940 2576
rect 2974 2542 3015 2576
rect 3049 2542 3090 2576
rect 3124 2542 3136 2576
rect 1946 2536 3136 2542
rect 26309 2025 26766 2026
rect 25823 2019 26774 2025
rect 26826 2019 26849 2025
rect 26901 2019 26924 2025
rect 26976 2019 26998 2025
rect 27050 2019 27072 2025
rect 27124 2019 27146 2025
rect 27198 2019 27880 2025
rect 25823 1985 25855 2019
rect 25889 1985 25928 2019
rect 25962 1985 26001 2019
rect 26035 1985 26074 2019
rect 26108 1985 26147 2019
rect 26181 1985 26220 2019
rect 26254 1985 26293 2019
rect 26327 1985 26366 2019
rect 26400 1985 26439 2019
rect 26473 1985 26512 2019
rect 26546 1985 26585 2019
rect 26619 1985 26658 2019
rect 26692 1985 26731 2019
rect 26765 1985 26774 2019
rect 26838 1985 26849 2019
rect 26911 1985 26924 2019
rect 26984 1985 26998 2019
rect 27056 1985 27072 2019
rect 27128 1985 27146 2019
rect 27200 1985 27238 2019
rect 27272 1985 27310 2019
rect 27344 1985 27382 2019
rect 27416 1985 27454 2019
rect 27488 1985 27526 2019
rect 27560 1985 27598 2019
rect 27632 1985 27670 2019
rect 27704 1985 27742 2019
rect 27776 1985 27814 2019
rect 27848 1985 27880 2019
rect 25823 1973 26774 1985
rect 26826 1973 26849 1985
rect 26901 1973 26924 1985
rect 26976 1973 26998 1985
rect 27050 1973 27072 1985
rect 27124 1973 27146 1985
rect 27198 1973 27880 1985
rect 25823 1961 27880 1973
rect 25823 1939 26774 1961
rect 26826 1939 26849 1961
rect 26901 1939 26924 1961
rect 26976 1939 26998 1961
rect 27050 1939 27072 1961
rect 27124 1939 27146 1961
rect 27198 1939 27880 1961
rect 25823 1905 25855 1939
rect 25889 1905 25928 1939
rect 25962 1905 26001 1939
rect 26035 1905 26074 1939
rect 26108 1905 26147 1939
rect 26181 1905 26220 1939
rect 26254 1905 26293 1939
rect 26327 1905 26366 1939
rect 26400 1905 26439 1939
rect 26473 1905 26512 1939
rect 26546 1905 26585 1939
rect 26619 1905 26658 1939
rect 26692 1905 26731 1939
rect 26765 1909 26774 1939
rect 26838 1909 26849 1939
rect 26911 1909 26924 1939
rect 26984 1909 26998 1939
rect 27056 1909 27072 1939
rect 27128 1909 27146 1939
rect 26765 1905 26804 1909
rect 26838 1905 26877 1909
rect 26911 1905 26950 1909
rect 26984 1905 27022 1909
rect 27056 1905 27094 1909
rect 27128 1905 27166 1909
rect 27200 1905 27238 1939
rect 27272 1905 27310 1939
rect 27344 1905 27382 1939
rect 27416 1905 27454 1939
rect 27488 1905 27526 1939
rect 27560 1905 27598 1939
rect 27632 1905 27670 1939
rect 27704 1905 27742 1939
rect 27776 1905 27814 1939
rect 27848 1905 27880 1939
rect 25823 1859 27880 1905
rect 25823 1825 25855 1859
rect 25889 1825 25928 1859
rect 25962 1825 26001 1859
rect 26035 1825 26074 1859
rect 26108 1825 26147 1859
rect 26181 1825 26220 1859
rect 26254 1825 26293 1859
rect 26327 1825 26366 1859
rect 26400 1825 26439 1859
rect 26473 1825 26512 1859
rect 26546 1825 26585 1859
rect 26619 1825 26658 1859
rect 26692 1825 26731 1859
rect 26765 1825 26804 1859
rect 26838 1825 26877 1859
rect 26911 1825 26950 1859
rect 26984 1825 27022 1859
rect 27056 1825 27094 1859
rect 27128 1825 27166 1859
rect 27200 1825 27238 1859
rect 27272 1825 27310 1859
rect 27344 1825 27382 1859
rect 27416 1825 27454 1859
rect 27488 1825 27526 1859
rect 27560 1825 27598 1859
rect 27632 1825 27670 1859
rect 27704 1825 27742 1859
rect 27776 1825 27814 1859
rect 27848 1825 27880 1859
rect 25823 1779 27880 1825
rect 25823 1745 25855 1779
rect 25889 1745 25928 1779
rect 25962 1745 26001 1779
rect 26035 1745 26074 1779
rect 26108 1745 26147 1779
rect 26181 1745 26220 1779
rect 26254 1745 26293 1779
rect 26327 1745 26366 1779
rect 26400 1745 26439 1779
rect 26473 1745 26512 1779
rect 26546 1745 26585 1779
rect 26619 1745 26658 1779
rect 26692 1745 26731 1779
rect 26765 1745 26804 1779
rect 26838 1745 26877 1779
rect 26911 1745 26950 1779
rect 26984 1745 27022 1779
rect 27056 1745 27094 1779
rect 27128 1745 27166 1779
rect 27200 1745 27238 1779
rect 27272 1745 27310 1779
rect 27344 1745 27382 1779
rect 27416 1745 27454 1779
rect 27488 1745 27526 1779
rect 27560 1745 27598 1779
rect 27632 1745 27670 1779
rect 27704 1745 27742 1779
rect 27776 1745 27814 1779
rect 27848 1745 27880 1779
rect 25823 1739 27880 1745
rect 26309 1591 26766 1739
<< via1 >>
rect 17645 36784 17697 36836
rect 17711 36784 17763 36836
rect 17645 36706 17697 36758
rect 17711 36706 17763 36758
rect 17645 36627 17697 36679
rect 17711 36627 17763 36679
rect 17645 36548 17697 36600
rect 17711 36548 17763 36600
rect 18018 32790 18022 32818
rect 18022 32790 18056 32818
rect 18056 32790 18070 32818
rect 18128 32790 18142 32818
rect 18142 32790 18180 32818
rect 18018 32766 18070 32790
rect 18128 32766 18180 32790
rect 18018 32718 18022 32751
rect 18022 32718 18056 32751
rect 18056 32718 18070 32751
rect 18128 32718 18142 32751
rect 18142 32718 18180 32751
rect 18018 32699 18070 32718
rect 18128 32699 18180 32718
rect 18018 32680 18070 32684
rect 18128 32680 18180 32684
rect 18018 32646 18022 32680
rect 18022 32646 18056 32680
rect 18056 32646 18070 32680
rect 18128 32646 18142 32680
rect 18142 32646 18180 32680
rect 18018 32632 18070 32646
rect 18128 32632 18180 32646
rect 18018 32608 18070 32617
rect 18128 32608 18180 32617
rect 18018 32574 18022 32608
rect 18022 32574 18056 32608
rect 18056 32574 18070 32608
rect 18128 32574 18142 32608
rect 18142 32574 18180 32608
rect 18018 32565 18070 32574
rect 18128 32565 18180 32574
rect 18018 32536 18070 32550
rect 18128 32536 18180 32550
rect 18018 32502 18022 32536
rect 18022 32502 18056 32536
rect 18056 32502 18070 32536
rect 18128 32502 18142 32536
rect 18142 32502 18180 32536
rect 18018 32498 18070 32502
rect 18128 32498 18180 32502
rect 18018 32464 18070 32482
rect 18128 32464 18180 32482
rect 18018 32430 18022 32464
rect 18022 32430 18056 32464
rect 18056 32430 18070 32464
rect 18128 32430 18142 32464
rect 18142 32430 18180 32464
rect 18018 32392 18070 32414
rect 18128 32392 18180 32414
rect 18018 32362 18022 32392
rect 18022 32362 18056 32392
rect 18056 32362 18070 32392
rect 18128 32362 18142 32392
rect 18142 32362 18180 32392
rect 18018 32320 18070 32346
rect 18128 32320 18180 32346
rect 18018 32294 18022 32320
rect 18022 32294 18056 32320
rect 18056 32294 18070 32320
rect 18128 32294 18142 32320
rect 18142 32294 18180 32320
rect 18018 32248 18070 32278
rect 18128 32248 18180 32278
rect 18018 32226 18022 32248
rect 18022 32226 18056 32248
rect 18056 32226 18070 32248
rect 18128 32226 18142 32248
rect 18142 32226 18180 32248
rect 18018 32176 18070 32210
rect 18128 32176 18180 32210
rect 18018 32158 18022 32176
rect 18022 32158 18056 32176
rect 18056 32158 18070 32176
rect 18128 32158 18142 32176
rect 18142 32158 18180 32176
rect 18018 32104 18070 32142
rect 18128 32104 18180 32142
rect 18018 32090 18022 32104
rect 18022 32090 18056 32104
rect 18056 32090 18070 32104
rect 18128 32090 18142 32104
rect 18142 32090 18180 32104
rect 18018 32070 18022 32074
rect 18022 32070 18056 32074
rect 18056 32070 18070 32074
rect 18128 32070 18142 32074
rect 18142 32070 18180 32074
rect 18018 32032 18070 32070
rect 18128 32032 18180 32070
rect 18018 32022 18022 32032
rect 18022 32022 18056 32032
rect 18056 32022 18070 32032
rect 18128 32022 18142 32032
rect 18142 32022 18180 32032
rect 215 31166 218 31195
rect 218 31166 252 31195
rect 252 31166 267 31195
rect 215 31143 267 31166
rect 313 31143 365 31195
rect 215 31094 218 31128
rect 218 31094 252 31128
rect 252 31094 267 31128
rect 215 31076 267 31094
rect 313 31076 365 31128
rect 215 31056 267 31061
rect 215 31022 218 31056
rect 218 31022 252 31056
rect 252 31022 267 31056
rect 215 31009 267 31022
rect 313 31009 365 31061
rect 959 31143 1011 31195
rect 959 31076 1011 31128
rect 959 31009 1011 31061
rect 22833 23222 22842 23241
rect 22842 23222 22876 23241
rect 22876 23222 22885 23241
rect 22833 23189 22885 23222
rect 22833 23149 22842 23176
rect 22842 23149 22876 23176
rect 22876 23149 22885 23176
rect 22833 23124 22885 23149
rect 22833 23110 22885 23111
rect 22833 23076 22842 23110
rect 22842 23076 22876 23110
rect 22876 23076 22885 23110
rect 22833 23059 22885 23076
rect 22833 23037 22885 23045
rect 22833 23003 22842 23037
rect 22842 23003 22876 23037
rect 22876 23003 22885 23037
rect 22833 22993 22885 23003
rect 23768 23189 23820 23241
rect 23832 23189 23884 23241
rect 23896 23189 23948 23241
rect 23768 23091 23820 23143
rect 23832 23091 23884 23143
rect 23896 23091 23948 23143
rect 23768 22993 23820 23045
rect 23832 22993 23884 23045
rect 23896 22993 23948 23045
rect 1944 11501 1996 11553
rect 2012 11501 2064 11553
rect 1944 11433 1996 11485
rect 2012 11433 2064 11485
rect 1944 11365 1996 11417
rect 2012 11365 2064 11417
rect 1944 11296 1996 11348
rect 2012 11296 2064 11348
rect 17950 11223 17955 11252
rect 17955 11223 18000 11252
rect 18000 11223 18002 11252
rect 18016 11223 18034 11252
rect 18034 11223 18068 11252
rect 18081 11223 18113 11252
rect 18113 11223 18133 11252
rect 17950 11200 18002 11223
rect 18016 11200 18068 11223
rect 18081 11200 18133 11223
rect 18146 11223 18158 11252
rect 18158 11223 18192 11252
rect 18192 11223 18198 11252
rect 18146 11200 18198 11223
rect 18494 11221 18500 11252
rect 18500 11221 18534 11252
rect 18534 11221 18546 11252
rect 18494 11200 18546 11221
rect 18560 11221 18585 11252
rect 18585 11221 18612 11252
rect 18625 11221 18669 11252
rect 18669 11221 18677 11252
rect 18690 11221 18703 11252
rect 18703 11221 18742 11252
rect 18560 11200 18612 11221
rect 18625 11200 18677 11221
rect 18690 11200 18742 11221
rect 19217 11200 19269 11252
rect 19283 11200 19335 11252
rect 19348 11200 19400 11252
rect 19413 11200 19465 11252
rect 16811 10120 16815 10154
rect 16815 10120 16854 10154
rect 16854 10120 16863 10154
rect 16811 10102 16863 10120
rect 16811 10082 16863 10090
rect 16811 10048 16815 10082
rect 16815 10048 16854 10082
rect 16854 10048 16863 10082
rect 16811 10038 16863 10048
rect 27498 10307 27501 10331
rect 27501 10307 27535 10331
rect 27535 10307 27573 10331
rect 27573 10307 27607 10331
rect 27607 10307 27645 10331
rect 27645 10307 27679 10331
rect 27679 10307 27717 10331
rect 27717 10307 27751 10331
rect 27751 10307 27789 10331
rect 27789 10307 27806 10331
rect 27498 10268 27806 10307
rect 27498 10234 27501 10268
rect 27501 10234 27535 10268
rect 27535 10234 27573 10268
rect 27573 10234 27607 10268
rect 27607 10234 27645 10268
rect 27645 10234 27679 10268
rect 27679 10234 27717 10268
rect 27717 10234 27751 10268
rect 27751 10234 27789 10268
rect 27789 10234 27806 10268
rect 27498 10195 27806 10234
rect 27498 10161 27501 10195
rect 27501 10161 27535 10195
rect 27535 10161 27573 10195
rect 27573 10161 27607 10195
rect 27607 10161 27645 10195
rect 27645 10161 27679 10195
rect 27679 10161 27717 10195
rect 27717 10161 27751 10195
rect 27751 10161 27789 10195
rect 27789 10161 27806 10195
rect 27498 10122 27806 10161
rect 27498 10088 27501 10122
rect 27501 10088 27535 10122
rect 27535 10088 27573 10122
rect 27573 10088 27607 10122
rect 27607 10088 27645 10122
rect 27645 10088 27679 10122
rect 27679 10088 27717 10122
rect 27717 10088 27751 10122
rect 27751 10088 27789 10122
rect 27789 10088 27806 10122
rect 27498 10049 27806 10088
rect 27498 10015 27501 10049
rect 27501 10015 27535 10049
rect 27535 10015 27573 10049
rect 27573 10015 27607 10049
rect 27607 10015 27645 10049
rect 27645 10015 27679 10049
rect 27679 10015 27717 10049
rect 27717 10015 27751 10049
rect 27751 10015 27789 10049
rect 27789 10015 27806 10049
rect 27498 9976 27806 10015
rect 27498 9942 27501 9976
rect 27501 9942 27535 9976
rect 27535 9942 27573 9976
rect 27573 9942 27607 9976
rect 27607 9942 27645 9976
rect 27645 9942 27679 9976
rect 27679 9942 27717 9976
rect 27717 9942 27751 9976
rect 27751 9942 27789 9976
rect 27789 9942 27806 9976
rect 27498 9902 27806 9942
rect 27498 9868 27501 9902
rect 27501 9868 27535 9902
rect 27535 9868 27573 9902
rect 27573 9868 27607 9902
rect 27607 9868 27645 9902
rect 27645 9868 27679 9902
rect 27679 9868 27717 9902
rect 27717 9868 27751 9902
rect 27751 9868 27789 9902
rect 27789 9868 27806 9902
rect 27498 9828 27806 9868
rect 27498 9794 27501 9828
rect 27501 9794 27535 9828
rect 27535 9794 27573 9828
rect 27573 9794 27607 9828
rect 27607 9794 27645 9828
rect 27645 9794 27679 9828
rect 27679 9794 27717 9828
rect 27717 9794 27751 9828
rect 27751 9794 27789 9828
rect 27789 9794 27806 9828
rect 27498 9754 27806 9794
rect 27498 9720 27501 9754
rect 27501 9720 27535 9754
rect 27535 9720 27573 9754
rect 27573 9720 27607 9754
rect 27607 9720 27645 9754
rect 27645 9720 27679 9754
rect 27679 9720 27717 9754
rect 27717 9720 27751 9754
rect 27751 9720 27789 9754
rect 27789 9720 27806 9754
rect 27498 9680 27806 9720
rect 27498 9646 27501 9680
rect 27501 9646 27535 9680
rect 27535 9646 27573 9680
rect 27573 9646 27607 9680
rect 27607 9646 27645 9680
rect 27645 9646 27679 9680
rect 27679 9646 27717 9680
rect 27717 9646 27751 9680
rect 27751 9646 27789 9680
rect 27789 9646 27806 9680
rect 27498 9606 27806 9646
rect 27498 9572 27501 9606
rect 27501 9572 27535 9606
rect 27535 9572 27573 9606
rect 27573 9572 27607 9606
rect 27607 9572 27645 9606
rect 27645 9572 27679 9606
rect 27679 9572 27717 9606
rect 27717 9572 27751 9606
rect 27751 9572 27789 9606
rect 27789 9572 27806 9606
rect 27498 9532 27806 9572
rect 27498 9498 27501 9532
rect 27501 9498 27535 9532
rect 27535 9498 27573 9532
rect 27573 9498 27607 9532
rect 27607 9498 27645 9532
rect 27645 9498 27679 9532
rect 27679 9498 27717 9532
rect 27717 9498 27751 9532
rect 27751 9498 27789 9532
rect 27789 9498 27806 9532
rect 27498 9458 27806 9498
rect 27498 9424 27501 9458
rect 27501 9424 27535 9458
rect 27535 9424 27573 9458
rect 27573 9424 27607 9458
rect 27607 9424 27645 9458
rect 27645 9424 27679 9458
rect 27679 9424 27717 9458
rect 27717 9424 27751 9458
rect 27751 9424 27789 9458
rect 27789 9424 27806 9458
rect 27498 9384 27806 9424
rect 27498 9350 27501 9384
rect 27501 9350 27535 9384
rect 27535 9350 27573 9384
rect 27573 9350 27607 9384
rect 27607 9350 27645 9384
rect 27645 9350 27679 9384
rect 27679 9350 27717 9384
rect 27717 9350 27751 9384
rect 27751 9350 27789 9384
rect 27789 9350 27806 9384
rect 27498 9319 27806 9350
rect 27498 9276 27501 9306
rect 27501 9276 27535 9306
rect 27535 9276 27550 9306
rect 27498 9254 27550 9276
rect 27562 9276 27573 9306
rect 27573 9276 27607 9306
rect 27607 9276 27614 9306
rect 27562 9254 27614 9276
rect 27626 9276 27645 9306
rect 27645 9276 27678 9306
rect 27690 9276 27717 9306
rect 27717 9276 27742 9306
rect 27754 9276 27789 9306
rect 27789 9276 27806 9306
rect 27626 9254 27678 9276
rect 27690 9254 27742 9276
rect 27754 9254 27806 9276
rect 27498 9236 27550 9241
rect 27498 9202 27501 9236
rect 27501 9202 27535 9236
rect 27535 9202 27550 9236
rect 27498 9189 27550 9202
rect 27562 9236 27614 9241
rect 27562 9202 27573 9236
rect 27573 9202 27607 9236
rect 27607 9202 27614 9236
rect 27562 9189 27614 9202
rect 27626 9236 27678 9241
rect 27690 9236 27742 9241
rect 27754 9236 27806 9241
rect 27626 9202 27645 9236
rect 27645 9202 27678 9236
rect 27690 9202 27717 9236
rect 27717 9202 27742 9236
rect 27754 9202 27789 9236
rect 27789 9202 27806 9236
rect 27626 9189 27678 9202
rect 27690 9189 27742 9202
rect 27754 9189 27806 9202
rect 27498 9162 27550 9176
rect 27498 9128 27501 9162
rect 27501 9128 27535 9162
rect 27535 9128 27550 9162
rect 27498 9124 27550 9128
rect 27562 9162 27614 9176
rect 27562 9128 27573 9162
rect 27573 9128 27607 9162
rect 27607 9128 27614 9162
rect 27562 9124 27614 9128
rect 27626 9162 27678 9176
rect 27690 9162 27742 9176
rect 27754 9162 27806 9176
rect 27626 9128 27645 9162
rect 27645 9128 27678 9162
rect 27690 9128 27717 9162
rect 27717 9128 27742 9162
rect 27754 9128 27789 9162
rect 27789 9128 27806 9162
rect 27626 9124 27678 9128
rect 27690 9124 27742 9128
rect 27754 9124 27806 9128
rect 27498 9088 27550 9111
rect 27498 9059 27501 9088
rect 27501 9059 27535 9088
rect 27535 9059 27550 9088
rect 27562 9088 27614 9111
rect 27562 9059 27573 9088
rect 27573 9059 27607 9088
rect 27607 9059 27614 9088
rect 27626 9088 27678 9111
rect 27690 9088 27742 9111
rect 27754 9088 27806 9111
rect 27626 9059 27645 9088
rect 27645 9059 27678 9088
rect 27690 9059 27717 9088
rect 27717 9059 27742 9088
rect 27754 9059 27789 9088
rect 27789 9059 27806 9088
rect 27498 9014 27550 9046
rect 27498 8994 27501 9014
rect 27501 8994 27535 9014
rect 27535 8994 27550 9014
rect 27562 9014 27614 9046
rect 27562 8994 27573 9014
rect 27573 8994 27607 9014
rect 27607 8994 27614 9014
rect 27626 9014 27678 9046
rect 27690 9014 27742 9046
rect 27754 9014 27806 9046
rect 27626 8994 27645 9014
rect 27645 8994 27678 9014
rect 27690 8994 27717 9014
rect 27717 8994 27742 9014
rect 27754 8994 27789 9014
rect 27789 8994 27806 9014
rect 27498 8980 27501 8981
rect 27501 8980 27535 8981
rect 27535 8980 27550 8981
rect 27498 8940 27550 8980
rect 27498 8929 27501 8940
rect 27501 8929 27535 8940
rect 27535 8929 27550 8940
rect 27562 8980 27573 8981
rect 27573 8980 27607 8981
rect 27607 8980 27614 8981
rect 27562 8940 27614 8980
rect 27562 8929 27573 8940
rect 27573 8929 27607 8940
rect 27607 8929 27614 8940
rect 27626 8980 27645 8981
rect 27645 8980 27678 8981
rect 27690 8980 27717 8981
rect 27717 8980 27742 8981
rect 27754 8980 27789 8981
rect 27789 8980 27806 8981
rect 27626 8940 27678 8980
rect 27690 8940 27742 8980
rect 27754 8940 27806 8980
rect 27626 8929 27645 8940
rect 27645 8929 27678 8940
rect 27690 8929 27717 8940
rect 27717 8929 27742 8940
rect 27754 8929 27789 8940
rect 27789 8929 27806 8940
rect 27498 8906 27501 8916
rect 27501 8906 27535 8916
rect 27535 8906 27550 8916
rect 27498 8866 27550 8906
rect 27498 8864 27501 8866
rect 27501 8864 27535 8866
rect 27535 8864 27550 8866
rect 27562 8906 27573 8916
rect 27573 8906 27607 8916
rect 27607 8906 27614 8916
rect 27562 8866 27614 8906
rect 27562 8864 27573 8866
rect 27573 8864 27607 8866
rect 27607 8864 27614 8866
rect 27626 8906 27645 8916
rect 27645 8906 27678 8916
rect 27690 8906 27717 8916
rect 27717 8906 27742 8916
rect 27754 8906 27789 8916
rect 27789 8906 27806 8916
rect 27626 8866 27678 8906
rect 27690 8866 27742 8906
rect 27754 8866 27806 8906
rect 27626 8864 27645 8866
rect 27645 8864 27678 8866
rect 27690 8864 27717 8866
rect 27717 8864 27742 8866
rect 27754 8864 27789 8866
rect 27789 8864 27806 8866
rect 27498 8832 27501 8851
rect 27501 8832 27535 8851
rect 27535 8832 27550 8851
rect 27498 8799 27550 8832
rect 27562 8832 27573 8851
rect 27573 8832 27607 8851
rect 27607 8832 27614 8851
rect 27562 8799 27614 8832
rect 27626 8832 27645 8851
rect 27645 8832 27678 8851
rect 27690 8832 27717 8851
rect 27717 8832 27742 8851
rect 27754 8832 27789 8851
rect 27789 8832 27806 8851
rect 27626 8799 27678 8832
rect 27690 8799 27742 8832
rect 27754 8799 27806 8832
rect 27498 8758 27501 8786
rect 27501 8758 27535 8786
rect 27535 8758 27550 8786
rect 27498 8734 27550 8758
rect 27562 8758 27573 8786
rect 27573 8758 27607 8786
rect 27607 8758 27614 8786
rect 27562 8734 27614 8758
rect 27626 8758 27645 8786
rect 27645 8758 27678 8786
rect 27690 8758 27717 8786
rect 27717 8758 27742 8786
rect 27754 8758 27789 8786
rect 27789 8758 27806 8786
rect 27626 8734 27678 8758
rect 27690 8734 27742 8758
rect 27754 8734 27806 8758
rect 27498 8718 27550 8721
rect 27498 8684 27501 8718
rect 27501 8684 27535 8718
rect 27535 8684 27550 8718
rect 27498 8669 27550 8684
rect 27562 8718 27614 8721
rect 27562 8684 27573 8718
rect 27573 8684 27607 8718
rect 27607 8684 27614 8718
rect 27562 8669 27614 8684
rect 27626 8718 27678 8721
rect 27690 8718 27742 8721
rect 27754 8718 27806 8721
rect 27626 8684 27645 8718
rect 27645 8684 27678 8718
rect 27690 8684 27717 8718
rect 27717 8684 27742 8718
rect 27754 8684 27789 8718
rect 27789 8684 27806 8718
rect 27626 8669 27678 8684
rect 27690 8669 27742 8684
rect 27754 8669 27806 8684
rect 27498 8644 27550 8656
rect 27498 8610 27501 8644
rect 27501 8610 27535 8644
rect 27535 8610 27550 8644
rect 27498 8604 27550 8610
rect 27562 8644 27614 8656
rect 27562 8610 27573 8644
rect 27573 8610 27607 8644
rect 27607 8610 27614 8644
rect 27562 8604 27614 8610
rect 27626 8644 27678 8656
rect 27690 8644 27742 8656
rect 27754 8644 27806 8656
rect 27626 8610 27645 8644
rect 27645 8610 27678 8644
rect 27690 8610 27717 8644
rect 27717 8610 27742 8644
rect 27754 8610 27789 8644
rect 27789 8610 27806 8644
rect 27626 8604 27678 8610
rect 27690 8604 27742 8610
rect 27754 8604 27806 8610
rect 13565 7244 13617 7296
rect 13631 7244 13683 7296
rect 13697 7244 13749 7296
rect 13763 7244 13815 7296
rect 13828 7244 13880 7296
rect 13893 7244 13945 7296
rect 13565 7158 13617 7210
rect 13631 7158 13683 7210
rect 13697 7158 13749 7210
rect 13763 7158 13815 7210
rect 13828 7158 13880 7210
rect 13893 7158 13945 7210
rect 14883 7246 14935 7298
rect 14956 7246 15008 7298
rect 15028 7246 15080 7298
rect 14883 7158 14935 7210
rect 14956 7158 15008 7210
rect 15028 7158 15080 7210
rect 2103 4268 2155 4320
rect 2187 4268 2239 4320
rect 2103 4200 2155 4252
rect 2187 4200 2239 4252
rect 2103 4131 2155 4183
rect 2187 4131 2239 4183
rect 2103 3637 2155 3638
rect 2103 3603 2105 3637
rect 2105 3603 2155 3637
rect 2103 3586 2155 3603
rect 2187 3586 2239 3638
rect 2103 3561 2155 3570
rect 2103 3527 2105 3561
rect 2105 3527 2155 3561
rect 2103 3518 2155 3527
rect 2187 3518 2239 3570
rect 2103 3485 2155 3502
rect 2103 3451 2105 3485
rect 2105 3451 2155 3485
rect 2103 3450 2155 3451
rect 2187 3450 2239 3502
rect 26774 3197 26826 3249
rect 26849 3197 26901 3249
rect 26924 3197 26976 3249
rect 26998 3197 27050 3249
rect 27072 3197 27124 3249
rect 27146 3197 27198 3249
rect 26774 3121 26826 3173
rect 26849 3121 26901 3173
rect 26924 3121 26976 3173
rect 26998 3121 27050 3173
rect 27072 3121 27124 3173
rect 27146 3121 27198 3173
rect 26774 3045 26826 3097
rect 26849 3045 26901 3097
rect 26924 3045 26976 3097
rect 26998 3045 27050 3097
rect 27072 3045 27124 3097
rect 27146 3045 27198 3097
rect 2103 2652 2110 2686
rect 2110 2652 2144 2686
rect 2144 2652 2155 2686
rect 2187 2652 2220 2686
rect 2220 2652 2239 2686
rect 2103 2634 2155 2652
rect 2187 2634 2239 2652
rect 2103 2576 2155 2594
rect 2187 2576 2239 2594
rect 2103 2542 2110 2576
rect 2110 2542 2144 2576
rect 2144 2542 2155 2576
rect 2187 2542 2220 2576
rect 2220 2542 2239 2576
rect 26774 2019 26826 2025
rect 26849 2019 26901 2025
rect 26924 2019 26976 2025
rect 26998 2019 27050 2025
rect 27072 2019 27124 2025
rect 27146 2019 27198 2025
rect 26774 1985 26804 2019
rect 26804 1985 26826 2019
rect 26849 1985 26877 2019
rect 26877 1985 26901 2019
rect 26924 1985 26950 2019
rect 26950 1985 26976 2019
rect 26998 1985 27022 2019
rect 27022 1985 27050 2019
rect 27072 1985 27094 2019
rect 27094 1985 27124 2019
rect 27146 1985 27166 2019
rect 27166 1985 27198 2019
rect 26774 1973 26826 1985
rect 26849 1973 26901 1985
rect 26924 1973 26976 1985
rect 26998 1973 27050 1985
rect 27072 1973 27124 1985
rect 27146 1973 27198 1985
rect 26774 1939 26826 1961
rect 26849 1939 26901 1961
rect 26924 1939 26976 1961
rect 26998 1939 27050 1961
rect 27072 1939 27124 1961
rect 27146 1939 27198 1961
rect 26774 1909 26804 1939
rect 26804 1909 26826 1939
rect 26849 1909 26877 1939
rect 26877 1909 26901 1939
rect 26924 1909 26950 1939
rect 26950 1909 26976 1939
rect 26998 1909 27022 1939
rect 27022 1909 27050 1939
rect 27072 1909 27094 1939
rect 27094 1909 27124 1939
rect 27146 1909 27166 1939
rect 27166 1909 27198 1939
<< metal2 >>
rect 17650 36842 17758 36843
rect 17645 36836 17763 36842
rect 17697 36834 17711 36836
rect 17645 36778 17676 36784
rect 17732 36778 17763 36784
rect 17645 36758 17763 36778
rect 17697 36720 17711 36758
rect 17645 36679 17676 36706
rect 17732 36679 17763 36706
rect 17697 36627 17711 36664
rect 17645 36605 17763 36627
rect 17645 36600 17676 36605
rect 17732 36600 17763 36605
rect 17697 36548 17711 36549
rect 17645 36542 17763 36548
rect 17650 36540 17758 36542
rect 17876 32818 18180 32824
rect 17876 32815 18018 32818
rect 17876 32759 17898 32815
rect 17954 32766 18018 32815
rect 18070 32766 18128 32818
rect 17954 32759 18180 32766
rect 17876 32751 18180 32759
rect 17876 32734 18018 32751
rect 17876 32678 17898 32734
rect 17954 32699 18018 32734
rect 18070 32699 18128 32751
rect 17954 32684 18180 32699
rect 17954 32678 18018 32684
rect 17876 32653 18018 32678
rect 17876 32597 17898 32653
rect 17954 32632 18018 32653
rect 18070 32632 18128 32684
rect 17954 32617 18180 32632
rect 17954 32597 18018 32617
rect 17876 32572 18018 32597
rect 17876 32516 17898 32572
rect 17954 32565 18018 32572
rect 18070 32565 18128 32617
rect 17954 32550 18180 32565
rect 17954 32516 18018 32550
rect 17876 32498 18018 32516
rect 18070 32498 18128 32550
rect 17876 32491 18180 32498
rect 17876 32435 17898 32491
rect 17954 32482 18180 32491
rect 17954 32435 18018 32482
rect 17876 32430 18018 32435
rect 18070 32430 18128 32482
rect 17876 32414 18180 32430
rect 17876 32409 18018 32414
rect 17876 32353 17898 32409
rect 17954 32362 18018 32409
rect 18070 32362 18128 32414
rect 17954 32353 18180 32362
rect 17876 32346 18180 32353
rect 17876 32327 18018 32346
rect 17876 32271 17898 32327
rect 17954 32294 18018 32327
rect 18070 32294 18128 32346
rect 17954 32278 18180 32294
rect 17954 32271 18018 32278
rect 17876 32245 18018 32271
rect 17876 32189 17898 32245
rect 17954 32226 18018 32245
rect 18070 32226 18128 32278
rect 17954 32210 18180 32226
rect 17954 32189 18018 32210
rect 17876 32163 18018 32189
rect 17876 32107 17898 32163
rect 17954 32158 18018 32163
rect 18070 32158 18128 32210
rect 17954 32142 18180 32158
rect 17954 32107 18018 32142
rect 17876 32090 18018 32107
rect 18070 32090 18128 32142
rect 17876 32081 18180 32090
rect 17876 32025 17898 32081
rect 17954 32074 18180 32081
rect 17954 32025 18018 32074
rect 17876 32022 18018 32025
rect 18070 32022 18128 32074
rect 17876 32016 18180 32022
rect 212 31195 1757 31201
rect 212 31143 215 31195
rect 267 31143 313 31195
rect 365 31143 959 31195
rect 1011 31143 1757 31195
rect 212 31128 1757 31143
rect 212 31076 215 31128
rect 267 31076 313 31128
rect 365 31076 959 31128
rect 1011 31094 1757 31128
tri 1757 31094 1864 31201 sw
rect 1011 31076 1864 31094
rect 212 31061 1864 31076
rect 212 31009 215 31061
rect 267 31009 313 31061
rect 365 31009 959 31061
rect 1011 31009 1864 31061
rect 212 31003 1864 31009
tri 1570 30932 1641 31003 ne
rect 1641 30909 1864 31003
rect 22833 23241 23948 23247
rect 22885 23189 23768 23241
rect 23820 23189 23832 23241
rect 23884 23189 23896 23241
rect 22833 23176 23948 23189
rect 22885 23143 23948 23176
rect 22885 23124 23768 23143
rect 22833 23111 23768 23124
rect 22885 23091 23768 23111
rect 23820 23091 23832 23143
rect 23884 23091 23896 23143
rect 22885 23059 23948 23091
rect 22833 23045 23948 23059
rect 22885 22993 23768 23045
rect 23820 22993 23832 23045
rect 23884 22993 23896 23045
rect 22833 22987 23948 22993
rect 1944 11553 2105 11559
rect 1996 11550 2012 11553
rect 2064 11550 2105 11553
rect 2005 11501 2012 11550
rect 1944 11494 1949 11501
rect 2005 11494 2049 11501
rect 1944 11485 2105 11494
rect 1996 11451 2012 11485
rect 2064 11451 2105 11485
rect 2005 11433 2012 11451
rect 1944 11417 1949 11433
rect 2005 11417 2049 11433
rect 2005 11395 2012 11417
rect 1996 11365 2012 11395
rect 2064 11365 2105 11395
rect 1944 11351 2105 11365
rect 1944 11348 1949 11351
rect 2005 11348 2049 11351
rect 2005 11296 2012 11348
rect 1944 11295 1949 11296
rect 2005 11295 2049 11296
rect 1944 11290 2105 11295
rect 1949 11286 2105 11290
rect 17944 11200 17950 11252
rect 18002 11200 18016 11252
rect 18068 11200 18081 11252
rect 18133 11200 18146 11252
rect 18198 11200 18494 11252
rect 18546 11200 18560 11252
rect 18612 11200 18625 11252
rect 18677 11200 18690 11252
rect 18742 11200 19217 11252
rect 19269 11200 19283 11252
rect 19335 11200 19348 11252
rect 19400 11200 19413 11252
rect 19465 11200 19471 11252
rect 27498 10331 27806 10337
rect 16811 10154 16867 10160
rect 16863 10102 16867 10154
rect 16811 10090 16867 10102
rect 16863 10038 16867 10090
rect 16811 9871 16867 10038
tri 16811 9863 16819 9871 ne
rect 16819 9863 16867 9871
tri 16867 9863 16897 9893 sw
tri 16819 9815 16867 9863 ne
rect 16867 9815 16897 9863
tri 16867 9785 16897 9815 ne
tri 16897 9785 16975 9863 sw
tri 16897 9729 16953 9785 ne
rect 16953 9729 17866 9785
rect 17922 9729 17979 9785
rect 18035 9729 18091 9785
rect 18147 9729 18156 9785
rect 27498 9306 27806 9319
rect 27550 9254 27562 9306
rect 27614 9254 27626 9306
rect 27678 9254 27690 9306
rect 27742 9254 27754 9306
rect 27498 9241 27806 9254
rect 27550 9189 27562 9241
rect 27614 9189 27626 9241
rect 27678 9189 27690 9241
rect 27742 9189 27754 9241
rect 27498 9176 27806 9189
rect 27550 9124 27562 9176
rect 27614 9124 27626 9176
rect 27678 9124 27690 9176
rect 27742 9124 27754 9176
rect 27498 9111 27806 9124
rect 27550 9059 27562 9111
rect 27614 9059 27626 9111
rect 27678 9059 27690 9111
rect 27742 9059 27754 9111
rect 27498 9046 27806 9059
rect 27550 8994 27562 9046
rect 27614 8994 27626 9046
rect 27678 8994 27690 9046
rect 27742 8994 27754 9046
rect 27498 8981 27806 8994
rect 27550 8929 27562 8981
rect 27614 8929 27626 8981
rect 27678 8929 27690 8981
rect 27742 8929 27754 8981
rect 27498 8916 27806 8929
rect 27550 8864 27562 8916
rect 27614 8864 27626 8916
rect 27678 8864 27690 8916
rect 27742 8864 27754 8916
rect 27498 8851 27806 8864
rect 27550 8799 27562 8851
rect 27614 8799 27626 8851
rect 27678 8799 27690 8851
rect 27742 8799 27754 8851
rect 27498 8786 27806 8799
rect 27550 8734 27562 8786
rect 27614 8734 27626 8786
rect 27678 8734 27690 8786
rect 27742 8734 27754 8786
rect 27498 8721 27806 8734
rect 27550 8669 27562 8721
rect 27614 8669 27626 8721
rect 27678 8669 27690 8721
rect 27742 8669 27754 8721
rect 27498 8656 27806 8669
rect 27550 8604 27562 8656
rect 27614 8604 27626 8656
rect 27678 8604 27690 8656
rect 27742 8604 27754 8656
rect 27498 8598 27806 8604
rect 13556 7298 15086 7299
rect 13556 7296 14883 7298
rect 13556 7244 13565 7296
rect 13617 7244 13631 7296
rect 13683 7244 13697 7296
rect 13749 7244 13763 7296
rect 13815 7244 13828 7296
rect 13880 7244 13893 7296
rect 13945 7256 14883 7296
rect 14935 7256 14956 7298
rect 13945 7244 14512 7256
rect 13556 7210 14512 7244
rect 13556 7158 13565 7210
rect 13617 7158 13631 7210
rect 13683 7158 13697 7210
rect 13749 7158 13763 7210
rect 13815 7158 13828 7210
rect 13880 7158 13893 7210
rect 13945 7200 14512 7210
rect 14568 7200 14617 7256
rect 14673 7200 14722 7256
rect 14778 7200 14827 7256
rect 15008 7246 15028 7298
rect 15080 7294 15086 7298
rect 15080 7256 15101 7294
rect 14883 7210 14932 7246
rect 14988 7210 15036 7246
rect 13945 7158 14883 7200
rect 14935 7158 14956 7200
rect 15008 7158 15028 7210
rect 15092 7200 15101 7256
rect 15080 7162 15101 7200
rect 15080 7158 15086 7162
rect 2103 4320 2239 4326
rect 2155 4268 2187 4320
rect 2103 4252 2239 4268
rect 2155 4200 2187 4252
rect 2103 4183 2239 4200
rect 2155 4131 2187 4183
rect 2103 3638 2239 4131
rect 2155 3586 2187 3638
rect 2103 3570 2239 3586
rect 2155 3518 2187 3570
rect 2103 3502 2239 3518
rect 2155 3450 2187 3502
rect 2103 2686 2239 3450
rect 2155 2634 2187 2686
rect 2103 2594 2239 2634
rect 2155 2542 2187 2594
rect 2103 2536 2239 2542
rect 26768 3197 26774 3249
rect 26826 3197 26849 3249
rect 26901 3197 26924 3249
rect 26976 3197 26998 3249
rect 27050 3197 27072 3249
rect 27124 3197 27146 3249
rect 27198 3197 27204 3249
rect 26768 3173 27204 3197
rect 26768 3121 26774 3173
rect 26826 3121 26849 3173
rect 26901 3121 26924 3173
rect 26976 3121 26998 3173
rect 27050 3121 27072 3173
rect 27124 3121 27146 3173
rect 27198 3121 27204 3173
rect 26768 3097 27204 3121
rect 26768 3045 26774 3097
rect 26826 3045 26849 3097
rect 26901 3045 26924 3097
rect 26976 3045 26998 3097
rect 27050 3045 27072 3097
rect 27124 3045 27146 3097
rect 27198 3045 27204 3097
rect 26768 2025 27204 3045
rect 26768 1973 26774 2025
rect 26826 1973 26849 2025
rect 26901 1973 26924 2025
rect 26976 1973 26998 2025
rect 27050 1973 27072 2025
rect 27124 1973 27146 2025
rect 27198 1973 27204 2025
rect 26768 1961 27204 1973
rect 26768 1909 26774 1961
rect 26826 1909 26849 1961
rect 26901 1909 26924 1961
rect 26976 1909 26998 1961
rect 27050 1909 27072 1961
rect 27124 1909 27146 1961
rect 27198 1909 27204 1961
<< via2 >>
rect 17676 36784 17697 36834
rect 17697 36784 17711 36834
rect 17711 36784 17732 36834
rect 17676 36778 17732 36784
rect 17676 36706 17697 36720
rect 17697 36706 17711 36720
rect 17711 36706 17732 36720
rect 17676 36679 17732 36706
rect 17676 36664 17697 36679
rect 17697 36664 17711 36679
rect 17711 36664 17732 36679
rect 17676 36600 17732 36605
rect 17676 36549 17697 36600
rect 17697 36549 17711 36600
rect 17711 36549 17732 36600
rect 17898 32759 17954 32815
rect 17898 32678 17954 32734
rect 17898 32597 17954 32653
rect 17898 32516 17954 32572
rect 17898 32435 17954 32491
rect 17898 32353 17954 32409
rect 17898 32271 17954 32327
rect 17898 32189 17954 32245
rect 17898 32107 17954 32163
rect 17898 32025 17954 32081
rect 1949 11501 1996 11550
rect 1996 11501 2005 11550
rect 2049 11501 2064 11550
rect 2064 11501 2105 11550
rect 1949 11494 2005 11501
rect 2049 11494 2105 11501
rect 1949 11433 1996 11451
rect 1996 11433 2005 11451
rect 2049 11433 2064 11451
rect 2064 11433 2105 11451
rect 1949 11417 2005 11433
rect 2049 11417 2105 11433
rect 1949 11395 1996 11417
rect 1996 11395 2005 11417
rect 2049 11395 2064 11417
rect 2064 11395 2105 11417
rect 1949 11348 2005 11351
rect 2049 11348 2105 11351
rect 1949 11296 1996 11348
rect 1996 11296 2005 11348
rect 2049 11296 2064 11348
rect 2064 11296 2105 11348
rect 1949 11295 2005 11296
rect 2049 11295 2105 11296
rect 17866 9729 17922 9785
rect 17979 9729 18035 9785
rect 18091 9729 18147 9785
rect 14512 7200 14568 7256
rect 14617 7200 14673 7256
rect 14722 7200 14778 7256
rect 14827 7200 14883 7256
rect 14932 7246 14935 7256
rect 14935 7246 14956 7256
rect 14956 7246 14988 7256
rect 15036 7246 15080 7256
rect 15080 7246 15092 7256
rect 14932 7210 14988 7246
rect 15036 7210 15092 7246
rect 14932 7200 14935 7210
rect 14935 7200 14956 7210
rect 14956 7200 14988 7210
rect 15036 7200 15080 7210
rect 15080 7200 15092 7210
<< metal3 >>
rect 17642 36834 17766 36845
rect 17642 36778 17676 36834
rect 17732 36778 17766 36834
rect 17642 36720 17766 36778
rect 17642 36664 17676 36720
rect 17732 36664 17766 36720
rect 17642 36605 17766 36664
rect 17642 36549 17676 36605
rect 17732 36549 17766 36605
tri 17592 35221 17642 35271 se
rect 17642 35221 17766 36549
tri 17525 35154 17592 35221 se
rect 17592 35154 17699 35221
tri 17699 35154 17766 35221 nw
tri 17401 35030 17525 35154 se
rect 17401 34148 17525 35030
tri 17525 34980 17699 35154 nw
tri 17401 34121 17428 34148 ne
rect 17428 34121 17525 34148
tri 17525 34121 17614 34210 sw
tri 17428 34024 17525 34121 ne
rect 17525 34024 17614 34121
tri 17525 33935 17614 34024 ne
tri 17614 33935 17800 34121 sw
tri 17614 33749 17800 33935 ne
tri 17800 33749 17986 33935 sw
tri 17800 33686 17863 33749 ne
rect 17863 32815 17986 33749
rect 17863 32759 17898 32815
rect 17954 32759 17986 32815
rect 17863 32734 17986 32759
rect 17863 32678 17898 32734
rect 17954 32678 17986 32734
rect 17863 32653 17986 32678
rect 17863 32597 17898 32653
rect 17954 32597 17986 32653
rect 17863 32572 17986 32597
rect 17863 32516 17898 32572
rect 17954 32516 17986 32572
rect 17863 32491 17986 32516
rect 17863 32435 17898 32491
rect 17954 32435 17986 32491
rect 17863 32409 17986 32435
rect 17863 32353 17898 32409
rect 17954 32353 17986 32409
rect 17863 32327 17986 32353
rect 17863 32271 17898 32327
rect 17954 32271 17986 32327
rect 17863 32245 17986 32271
rect 17863 32189 17898 32245
rect 17954 32189 17986 32245
rect 17863 32163 17986 32189
rect 17863 32107 17898 32163
rect 17954 32107 17986 32163
rect 17863 32081 17986 32107
rect 17863 32025 17898 32081
rect 17954 32025 17986 32081
rect 17863 32013 17986 32025
rect 1944 11550 2110 11555
rect 1944 11494 1949 11550
rect 2005 11494 2049 11550
rect 2105 11494 2110 11550
rect 1944 11451 2110 11494
rect 1944 11395 1949 11451
rect 2005 11395 2049 11451
rect 2105 11395 2110 11451
rect 1944 11351 2110 11395
rect 1944 11295 1949 11351
rect 2005 11295 2049 11351
rect 2105 11295 2110 11351
rect 1944 11290 2110 11295
rect 17861 9785 18152 9790
rect 17861 9729 17866 9785
rect 17922 9729 17979 9785
rect 18035 9729 18091 9785
rect 18147 9729 18152 9785
rect 17861 9724 18152 9729
rect 14507 7256 15097 7299
rect 14507 7200 14512 7256
rect 14568 7200 14617 7256
rect 14673 7200 14722 7256
rect 14778 7200 14827 7256
rect 14883 7200 14932 7256
rect 14988 7200 15036 7256
rect 15092 7200 15097 7256
rect 14507 7157 15097 7200
<< properties >>
string GDS_END 47705610
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 46641046
<< end >>
