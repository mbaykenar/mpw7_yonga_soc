magic
tech sky130B
magscale 1 2
timestamp 1662364221
<< obsli1 >>
rect 1104 2159 478860 117521
<< obsm1 >>
rect 14 824 479858 118720
<< metal2 >>
rect 18 119200 74 120000
rect 662 119200 718 120000
rect 1306 119200 1362 120000
rect 1950 119200 2006 120000
rect 2594 119200 2650 120000
rect 3882 119200 3938 120000
rect 4526 119200 4582 120000
rect 5170 119200 5226 120000
rect 5814 119200 5870 120000
rect 6458 119200 6514 120000
rect 7102 119200 7158 120000
rect 8390 119200 8446 120000
rect 9034 119200 9090 120000
rect 9678 119200 9734 120000
rect 10322 119200 10378 120000
rect 10966 119200 11022 120000
rect 12254 119200 12310 120000
rect 12898 119200 12954 120000
rect 13542 119200 13598 120000
rect 14186 119200 14242 120000
rect 14830 119200 14886 120000
rect 15474 119200 15530 120000
rect 16762 119200 16818 120000
rect 17406 119200 17462 120000
rect 18050 119200 18106 120000
rect 18694 119200 18750 120000
rect 19338 119200 19394 120000
rect 20626 119200 20682 120000
rect 21270 119200 21326 120000
rect 21914 119200 21970 120000
rect 22558 119200 22614 120000
rect 23202 119200 23258 120000
rect 23846 119200 23902 120000
rect 25134 119200 25190 120000
rect 25778 119200 25834 120000
rect 26422 119200 26478 120000
rect 27066 119200 27122 120000
rect 27710 119200 27766 120000
rect 28998 119200 29054 120000
rect 29642 119200 29698 120000
rect 30286 119200 30342 120000
rect 30930 119200 30986 120000
rect 31574 119200 31630 120000
rect 32218 119200 32274 120000
rect 33506 119200 33562 120000
rect 34150 119200 34206 120000
rect 34794 119200 34850 120000
rect 35438 119200 35494 120000
rect 36082 119200 36138 120000
rect 37370 119200 37426 120000
rect 38014 119200 38070 120000
rect 38658 119200 38714 120000
rect 39302 119200 39358 120000
rect 39946 119200 40002 120000
rect 40590 119200 40646 120000
rect 41878 119200 41934 120000
rect 42522 119200 42578 120000
rect 43166 119200 43222 120000
rect 43810 119200 43866 120000
rect 44454 119200 44510 120000
rect 45742 119200 45798 120000
rect 46386 119200 46442 120000
rect 47030 119200 47086 120000
rect 47674 119200 47730 120000
rect 48318 119200 48374 120000
rect 48962 119200 49018 120000
rect 50250 119200 50306 120000
rect 50894 119200 50950 120000
rect 51538 119200 51594 120000
rect 52182 119200 52238 120000
rect 52826 119200 52882 120000
rect 54114 119200 54170 120000
rect 54758 119200 54814 120000
rect 55402 119200 55458 120000
rect 56046 119200 56102 120000
rect 56690 119200 56746 120000
rect 57334 119200 57390 120000
rect 58622 119200 58678 120000
rect 59266 119200 59322 120000
rect 59910 119200 59966 120000
rect 60554 119200 60610 120000
rect 61198 119200 61254 120000
rect 62486 119200 62542 120000
rect 63130 119200 63186 120000
rect 63774 119200 63830 120000
rect 64418 119200 64474 120000
rect 65062 119200 65118 120000
rect 65706 119200 65762 120000
rect 66994 119200 67050 120000
rect 67638 119200 67694 120000
rect 68282 119200 68338 120000
rect 68926 119200 68982 120000
rect 69570 119200 69626 120000
rect 70214 119200 70270 120000
rect 71502 119200 71558 120000
rect 72146 119200 72202 120000
rect 72790 119200 72846 120000
rect 73434 119200 73490 120000
rect 74078 119200 74134 120000
rect 75366 119200 75422 120000
rect 76010 119200 76066 120000
rect 76654 119200 76710 120000
rect 77298 119200 77354 120000
rect 77942 119200 77998 120000
rect 78586 119200 78642 120000
rect 79874 119200 79930 120000
rect 80518 119200 80574 120000
rect 81162 119200 81218 120000
rect 81806 119200 81862 120000
rect 82450 119200 82506 120000
rect 83738 119200 83794 120000
rect 84382 119200 84438 120000
rect 85026 119200 85082 120000
rect 85670 119200 85726 120000
rect 86314 119200 86370 120000
rect 86958 119200 87014 120000
rect 88246 119200 88302 120000
rect 88890 119200 88946 120000
rect 89534 119200 89590 120000
rect 90178 119200 90234 120000
rect 90822 119200 90878 120000
rect 92110 119200 92166 120000
rect 92754 119200 92810 120000
rect 93398 119200 93454 120000
rect 94042 119200 94098 120000
rect 94686 119200 94742 120000
rect 95330 119200 95386 120000
rect 96618 119200 96674 120000
rect 97262 119200 97318 120000
rect 97906 119200 97962 120000
rect 98550 119200 98606 120000
rect 99194 119200 99250 120000
rect 100482 119200 100538 120000
rect 101126 119200 101182 120000
rect 101770 119200 101826 120000
rect 102414 119200 102470 120000
rect 103058 119200 103114 120000
rect 103702 119200 103758 120000
rect 104990 119200 105046 120000
rect 105634 119200 105690 120000
rect 106278 119200 106334 120000
rect 106922 119200 106978 120000
rect 107566 119200 107622 120000
rect 108854 119200 108910 120000
rect 109498 119200 109554 120000
rect 110142 119200 110198 120000
rect 110786 119200 110842 120000
rect 111430 119200 111486 120000
rect 112074 119200 112130 120000
rect 113362 119200 113418 120000
rect 114006 119200 114062 120000
rect 114650 119200 114706 120000
rect 115294 119200 115350 120000
rect 115938 119200 115994 120000
rect 117226 119200 117282 120000
rect 117870 119200 117926 120000
rect 118514 119200 118570 120000
rect 119158 119200 119214 120000
rect 119802 119200 119858 120000
rect 120446 119200 120502 120000
rect 121734 119200 121790 120000
rect 122378 119200 122434 120000
rect 123022 119200 123078 120000
rect 123666 119200 123722 120000
rect 124310 119200 124366 120000
rect 125598 119200 125654 120000
rect 126242 119200 126298 120000
rect 126886 119200 126942 120000
rect 127530 119200 127586 120000
rect 128174 119200 128230 120000
rect 128818 119200 128874 120000
rect 130106 119200 130162 120000
rect 130750 119200 130806 120000
rect 131394 119200 131450 120000
rect 132038 119200 132094 120000
rect 132682 119200 132738 120000
rect 133970 119200 134026 120000
rect 134614 119200 134670 120000
rect 135258 119200 135314 120000
rect 135902 119200 135958 120000
rect 136546 119200 136602 120000
rect 137190 119200 137246 120000
rect 138478 119200 138534 120000
rect 139122 119200 139178 120000
rect 139766 119200 139822 120000
rect 140410 119200 140466 120000
rect 141054 119200 141110 120000
rect 142342 119200 142398 120000
rect 142986 119200 143042 120000
rect 143630 119200 143686 120000
rect 144274 119200 144330 120000
rect 144918 119200 144974 120000
rect 145562 119200 145618 120000
rect 146850 119200 146906 120000
rect 147494 119200 147550 120000
rect 148138 119200 148194 120000
rect 148782 119200 148838 120000
rect 149426 119200 149482 120000
rect 150714 119200 150770 120000
rect 151358 119200 151414 120000
rect 152002 119200 152058 120000
rect 152646 119200 152702 120000
rect 153290 119200 153346 120000
rect 153934 119200 153990 120000
rect 155222 119200 155278 120000
rect 155866 119200 155922 120000
rect 156510 119200 156566 120000
rect 157154 119200 157210 120000
rect 157798 119200 157854 120000
rect 159086 119200 159142 120000
rect 159730 119200 159786 120000
rect 160374 119200 160430 120000
rect 161018 119200 161074 120000
rect 161662 119200 161718 120000
rect 162306 119200 162362 120000
rect 163594 119200 163650 120000
rect 164238 119200 164294 120000
rect 164882 119200 164938 120000
rect 165526 119200 165582 120000
rect 166170 119200 166226 120000
rect 166814 119200 166870 120000
rect 168102 119200 168158 120000
rect 168746 119200 168802 120000
rect 169390 119200 169446 120000
rect 170034 119200 170090 120000
rect 170678 119200 170734 120000
rect 171966 119200 172022 120000
rect 172610 119200 172666 120000
rect 173254 119200 173310 120000
rect 173898 119200 173954 120000
rect 174542 119200 174598 120000
rect 175186 119200 175242 120000
rect 176474 119200 176530 120000
rect 177118 119200 177174 120000
rect 177762 119200 177818 120000
rect 178406 119200 178462 120000
rect 179050 119200 179106 120000
rect 180338 119200 180394 120000
rect 180982 119200 181038 120000
rect 181626 119200 181682 120000
rect 182270 119200 182326 120000
rect 182914 119200 182970 120000
rect 183558 119200 183614 120000
rect 184846 119200 184902 120000
rect 185490 119200 185546 120000
rect 186134 119200 186190 120000
rect 186778 119200 186834 120000
rect 187422 119200 187478 120000
rect 188710 119200 188766 120000
rect 189354 119200 189410 120000
rect 189998 119200 190054 120000
rect 190642 119200 190698 120000
rect 191286 119200 191342 120000
rect 191930 119200 191986 120000
rect 193218 119200 193274 120000
rect 193862 119200 193918 120000
rect 194506 119200 194562 120000
rect 195150 119200 195206 120000
rect 195794 119200 195850 120000
rect 197082 119200 197138 120000
rect 197726 119200 197782 120000
rect 198370 119200 198426 120000
rect 199014 119200 199070 120000
rect 199658 119200 199714 120000
rect 200302 119200 200358 120000
rect 201590 119200 201646 120000
rect 202234 119200 202290 120000
rect 202878 119200 202934 120000
rect 203522 119200 203578 120000
rect 204166 119200 204222 120000
rect 205454 119200 205510 120000
rect 206098 119200 206154 120000
rect 206742 119200 206798 120000
rect 207386 119200 207442 120000
rect 208030 119200 208086 120000
rect 208674 119200 208730 120000
rect 209962 119200 210018 120000
rect 210606 119200 210662 120000
rect 211250 119200 211306 120000
rect 211894 119200 211950 120000
rect 212538 119200 212594 120000
rect 213826 119200 213882 120000
rect 214470 119200 214526 120000
rect 215114 119200 215170 120000
rect 215758 119200 215814 120000
rect 216402 119200 216458 120000
rect 217046 119200 217102 120000
rect 218334 119200 218390 120000
rect 218978 119200 219034 120000
rect 219622 119200 219678 120000
rect 220266 119200 220322 120000
rect 220910 119200 220966 120000
rect 222198 119200 222254 120000
rect 222842 119200 222898 120000
rect 223486 119200 223542 120000
rect 224130 119200 224186 120000
rect 224774 119200 224830 120000
rect 225418 119200 225474 120000
rect 226706 119200 226762 120000
rect 227350 119200 227406 120000
rect 227994 119200 228050 120000
rect 228638 119200 228694 120000
rect 229282 119200 229338 120000
rect 230570 119200 230626 120000
rect 231214 119200 231270 120000
rect 231858 119200 231914 120000
rect 232502 119200 232558 120000
rect 233146 119200 233202 120000
rect 233790 119200 233846 120000
rect 235078 119200 235134 120000
rect 235722 119200 235778 120000
rect 236366 119200 236422 120000
rect 237010 119200 237066 120000
rect 237654 119200 237710 120000
rect 238942 119200 238998 120000
rect 239586 119200 239642 120000
rect 240230 119200 240286 120000
rect 240874 119200 240930 120000
rect 241518 119200 241574 120000
rect 242162 119200 242218 120000
rect 243450 119200 243506 120000
rect 244094 119200 244150 120000
rect 244738 119200 244794 120000
rect 245382 119200 245438 120000
rect 246026 119200 246082 120000
rect 247314 119200 247370 120000
rect 247958 119200 248014 120000
rect 248602 119200 248658 120000
rect 249246 119200 249302 120000
rect 249890 119200 249946 120000
rect 250534 119200 250590 120000
rect 251822 119200 251878 120000
rect 252466 119200 252522 120000
rect 253110 119200 253166 120000
rect 253754 119200 253810 120000
rect 254398 119200 254454 120000
rect 255042 119200 255098 120000
rect 256330 119200 256386 120000
rect 256974 119200 257030 120000
rect 257618 119200 257674 120000
rect 258262 119200 258318 120000
rect 258906 119200 258962 120000
rect 260194 119200 260250 120000
rect 260838 119200 260894 120000
rect 261482 119200 261538 120000
rect 262126 119200 262182 120000
rect 262770 119200 262826 120000
rect 263414 119200 263470 120000
rect 264702 119200 264758 120000
rect 265346 119200 265402 120000
rect 265990 119200 266046 120000
rect 266634 119200 266690 120000
rect 267278 119200 267334 120000
rect 268566 119200 268622 120000
rect 269210 119200 269266 120000
rect 269854 119200 269910 120000
rect 270498 119200 270554 120000
rect 271142 119200 271198 120000
rect 271786 119200 271842 120000
rect 273074 119200 273130 120000
rect 273718 119200 273774 120000
rect 274362 119200 274418 120000
rect 275006 119200 275062 120000
rect 275650 119200 275706 120000
rect 276938 119200 276994 120000
rect 277582 119200 277638 120000
rect 278226 119200 278282 120000
rect 278870 119200 278926 120000
rect 279514 119200 279570 120000
rect 280158 119200 280214 120000
rect 281446 119200 281502 120000
rect 282090 119200 282146 120000
rect 282734 119200 282790 120000
rect 283378 119200 283434 120000
rect 284022 119200 284078 120000
rect 285310 119200 285366 120000
rect 285954 119200 286010 120000
rect 286598 119200 286654 120000
rect 287242 119200 287298 120000
rect 287886 119200 287942 120000
rect 288530 119200 288586 120000
rect 289818 119200 289874 120000
rect 290462 119200 290518 120000
rect 291106 119200 291162 120000
rect 291750 119200 291806 120000
rect 292394 119200 292450 120000
rect 293682 119200 293738 120000
rect 294326 119200 294382 120000
rect 294970 119200 295026 120000
rect 295614 119200 295670 120000
rect 296258 119200 296314 120000
rect 296902 119200 296958 120000
rect 298190 119200 298246 120000
rect 298834 119200 298890 120000
rect 299478 119200 299534 120000
rect 300122 119200 300178 120000
rect 300766 119200 300822 120000
rect 302054 119200 302110 120000
rect 302698 119200 302754 120000
rect 303342 119200 303398 120000
rect 303986 119200 304042 120000
rect 304630 119200 304686 120000
rect 305274 119200 305330 120000
rect 306562 119200 306618 120000
rect 307206 119200 307262 120000
rect 307850 119200 307906 120000
rect 308494 119200 308550 120000
rect 309138 119200 309194 120000
rect 310426 119200 310482 120000
rect 311070 119200 311126 120000
rect 311714 119200 311770 120000
rect 312358 119200 312414 120000
rect 313002 119200 313058 120000
rect 313646 119200 313702 120000
rect 314934 119200 314990 120000
rect 315578 119200 315634 120000
rect 316222 119200 316278 120000
rect 316866 119200 316922 120000
rect 317510 119200 317566 120000
rect 318798 119200 318854 120000
rect 319442 119200 319498 120000
rect 320086 119200 320142 120000
rect 320730 119200 320786 120000
rect 321374 119200 321430 120000
rect 322018 119200 322074 120000
rect 323306 119200 323362 120000
rect 323950 119200 324006 120000
rect 324594 119200 324650 120000
rect 325238 119200 325294 120000
rect 325882 119200 325938 120000
rect 327170 119200 327226 120000
rect 327814 119200 327870 120000
rect 328458 119200 328514 120000
rect 329102 119200 329158 120000
rect 329746 119200 329802 120000
rect 330390 119200 330446 120000
rect 331678 119200 331734 120000
rect 332322 119200 332378 120000
rect 332966 119200 333022 120000
rect 333610 119200 333666 120000
rect 334254 119200 334310 120000
rect 335542 119200 335598 120000
rect 336186 119200 336242 120000
rect 336830 119200 336886 120000
rect 337474 119200 337530 120000
rect 338118 119200 338174 120000
rect 338762 119200 338818 120000
rect 340050 119200 340106 120000
rect 340694 119200 340750 120000
rect 341338 119200 341394 120000
rect 341982 119200 342038 120000
rect 342626 119200 342682 120000
rect 343270 119200 343326 120000
rect 344558 119200 344614 120000
rect 345202 119200 345258 120000
rect 345846 119200 345902 120000
rect 346490 119200 346546 120000
rect 347134 119200 347190 120000
rect 348422 119200 348478 120000
rect 349066 119200 349122 120000
rect 349710 119200 349766 120000
rect 350354 119200 350410 120000
rect 350998 119200 351054 120000
rect 351642 119200 351698 120000
rect 352930 119200 352986 120000
rect 353574 119200 353630 120000
rect 354218 119200 354274 120000
rect 354862 119200 354918 120000
rect 355506 119200 355562 120000
rect 356794 119200 356850 120000
rect 357438 119200 357494 120000
rect 358082 119200 358138 120000
rect 358726 119200 358782 120000
rect 359370 119200 359426 120000
rect 360014 119200 360070 120000
rect 361302 119200 361358 120000
rect 361946 119200 362002 120000
rect 362590 119200 362646 120000
rect 363234 119200 363290 120000
rect 363878 119200 363934 120000
rect 365166 119200 365222 120000
rect 365810 119200 365866 120000
rect 366454 119200 366510 120000
rect 367098 119200 367154 120000
rect 367742 119200 367798 120000
rect 368386 119200 368442 120000
rect 369674 119200 369730 120000
rect 370318 119200 370374 120000
rect 370962 119200 371018 120000
rect 371606 119200 371662 120000
rect 372250 119200 372306 120000
rect 373538 119200 373594 120000
rect 374182 119200 374238 120000
rect 374826 119200 374882 120000
rect 375470 119200 375526 120000
rect 376114 119200 376170 120000
rect 376758 119200 376814 120000
rect 378046 119200 378102 120000
rect 378690 119200 378746 120000
rect 379334 119200 379390 120000
rect 379978 119200 380034 120000
rect 380622 119200 380678 120000
rect 381910 119200 381966 120000
rect 382554 119200 382610 120000
rect 383198 119200 383254 120000
rect 383842 119200 383898 120000
rect 384486 119200 384542 120000
rect 385130 119200 385186 120000
rect 386418 119200 386474 120000
rect 387062 119200 387118 120000
rect 387706 119200 387762 120000
rect 388350 119200 388406 120000
rect 388994 119200 389050 120000
rect 390282 119200 390338 120000
rect 390926 119200 390982 120000
rect 391570 119200 391626 120000
rect 392214 119200 392270 120000
rect 392858 119200 392914 120000
rect 393502 119200 393558 120000
rect 394790 119200 394846 120000
rect 395434 119200 395490 120000
rect 396078 119200 396134 120000
rect 396722 119200 396778 120000
rect 397366 119200 397422 120000
rect 398654 119200 398710 120000
rect 399298 119200 399354 120000
rect 399942 119200 399998 120000
rect 400586 119200 400642 120000
rect 401230 119200 401286 120000
rect 401874 119200 401930 120000
rect 403162 119200 403218 120000
rect 403806 119200 403862 120000
rect 404450 119200 404506 120000
rect 405094 119200 405150 120000
rect 405738 119200 405794 120000
rect 407026 119200 407082 120000
rect 407670 119200 407726 120000
rect 408314 119200 408370 120000
rect 408958 119200 409014 120000
rect 409602 119200 409658 120000
rect 410246 119200 410302 120000
rect 411534 119200 411590 120000
rect 412178 119200 412234 120000
rect 412822 119200 412878 120000
rect 413466 119200 413522 120000
rect 414110 119200 414166 120000
rect 415398 119200 415454 120000
rect 416042 119200 416098 120000
rect 416686 119200 416742 120000
rect 417330 119200 417386 120000
rect 417974 119200 418030 120000
rect 418618 119200 418674 120000
rect 419906 119200 419962 120000
rect 420550 119200 420606 120000
rect 421194 119200 421250 120000
rect 421838 119200 421894 120000
rect 422482 119200 422538 120000
rect 423770 119200 423826 120000
rect 424414 119200 424470 120000
rect 425058 119200 425114 120000
rect 425702 119200 425758 120000
rect 426346 119200 426402 120000
rect 426990 119200 427046 120000
rect 428278 119200 428334 120000
rect 428922 119200 428978 120000
rect 429566 119200 429622 120000
rect 430210 119200 430266 120000
rect 430854 119200 430910 120000
rect 432142 119200 432198 120000
rect 432786 119200 432842 120000
rect 433430 119200 433486 120000
rect 434074 119200 434130 120000
rect 434718 119200 434774 120000
rect 435362 119200 435418 120000
rect 436650 119200 436706 120000
rect 437294 119200 437350 120000
rect 437938 119200 437994 120000
rect 438582 119200 438638 120000
rect 439226 119200 439282 120000
rect 439870 119200 439926 120000
rect 441158 119200 441214 120000
rect 441802 119200 441858 120000
rect 442446 119200 442502 120000
rect 443090 119200 443146 120000
rect 443734 119200 443790 120000
rect 445022 119200 445078 120000
rect 445666 119200 445722 120000
rect 446310 119200 446366 120000
rect 446954 119200 447010 120000
rect 447598 119200 447654 120000
rect 448242 119200 448298 120000
rect 449530 119200 449586 120000
rect 450174 119200 450230 120000
rect 450818 119200 450874 120000
rect 451462 119200 451518 120000
rect 452106 119200 452162 120000
rect 453394 119200 453450 120000
rect 454038 119200 454094 120000
rect 454682 119200 454738 120000
rect 455326 119200 455382 120000
rect 455970 119200 456026 120000
rect 456614 119200 456670 120000
rect 457902 119200 457958 120000
rect 458546 119200 458602 120000
rect 459190 119200 459246 120000
rect 459834 119200 459890 120000
rect 460478 119200 460534 120000
rect 461766 119200 461822 120000
rect 462410 119200 462466 120000
rect 463054 119200 463110 120000
rect 463698 119200 463754 120000
rect 464342 119200 464398 120000
rect 464986 119200 465042 120000
rect 466274 119200 466330 120000
rect 466918 119200 466974 120000
rect 467562 119200 467618 120000
rect 468206 119200 468262 120000
rect 468850 119200 468906 120000
rect 470138 119200 470194 120000
rect 470782 119200 470838 120000
rect 471426 119200 471482 120000
rect 472070 119200 472126 120000
rect 472714 119200 472770 120000
rect 473358 119200 473414 120000
rect 474646 119200 474702 120000
rect 475290 119200 475346 120000
rect 475934 119200 475990 120000
rect 476578 119200 476634 120000
rect 477222 119200 477278 120000
rect 478510 119200 478566 120000
rect 479154 119200 479210 120000
rect 479798 119200 479854 120000
rect 18 0 74 800
rect 662 0 718 800
rect 1306 0 1362 800
rect 1950 0 2006 800
rect 2594 0 2650 800
rect 3238 0 3294 800
rect 4526 0 4582 800
rect 5170 0 5226 800
rect 5814 0 5870 800
rect 6458 0 6514 800
rect 7102 0 7158 800
rect 7746 0 7802 800
rect 9034 0 9090 800
rect 9678 0 9734 800
rect 10322 0 10378 800
rect 10966 0 11022 800
rect 11610 0 11666 800
rect 12898 0 12954 800
rect 13542 0 13598 800
rect 14186 0 14242 800
rect 14830 0 14886 800
rect 15474 0 15530 800
rect 16118 0 16174 800
rect 17406 0 17462 800
rect 18050 0 18106 800
rect 18694 0 18750 800
rect 19338 0 19394 800
rect 19982 0 20038 800
rect 21270 0 21326 800
rect 21914 0 21970 800
rect 22558 0 22614 800
rect 23202 0 23258 800
rect 23846 0 23902 800
rect 24490 0 24546 800
rect 25778 0 25834 800
rect 26422 0 26478 800
rect 27066 0 27122 800
rect 27710 0 27766 800
rect 28354 0 28410 800
rect 29642 0 29698 800
rect 30286 0 30342 800
rect 30930 0 30986 800
rect 31574 0 31630 800
rect 32218 0 32274 800
rect 32862 0 32918 800
rect 34150 0 34206 800
rect 34794 0 34850 800
rect 35438 0 35494 800
rect 36082 0 36138 800
rect 36726 0 36782 800
rect 38014 0 38070 800
rect 38658 0 38714 800
rect 39302 0 39358 800
rect 39946 0 40002 800
rect 40590 0 40646 800
rect 41234 0 41290 800
rect 42522 0 42578 800
rect 43166 0 43222 800
rect 43810 0 43866 800
rect 44454 0 44510 800
rect 45098 0 45154 800
rect 46386 0 46442 800
rect 47030 0 47086 800
rect 47674 0 47730 800
rect 48318 0 48374 800
rect 48962 0 49018 800
rect 49606 0 49662 800
rect 50894 0 50950 800
rect 51538 0 51594 800
rect 52182 0 52238 800
rect 52826 0 52882 800
rect 53470 0 53526 800
rect 54758 0 54814 800
rect 55402 0 55458 800
rect 56046 0 56102 800
rect 56690 0 56746 800
rect 57334 0 57390 800
rect 57978 0 58034 800
rect 59266 0 59322 800
rect 59910 0 59966 800
rect 60554 0 60610 800
rect 61198 0 61254 800
rect 61842 0 61898 800
rect 63130 0 63186 800
rect 63774 0 63830 800
rect 64418 0 64474 800
rect 65062 0 65118 800
rect 65706 0 65762 800
rect 66350 0 66406 800
rect 67638 0 67694 800
rect 68282 0 68338 800
rect 68926 0 68982 800
rect 69570 0 69626 800
rect 70214 0 70270 800
rect 71502 0 71558 800
rect 72146 0 72202 800
rect 72790 0 72846 800
rect 73434 0 73490 800
rect 74078 0 74134 800
rect 74722 0 74778 800
rect 76010 0 76066 800
rect 76654 0 76710 800
rect 77298 0 77354 800
rect 77942 0 77998 800
rect 78586 0 78642 800
rect 79874 0 79930 800
rect 80518 0 80574 800
rect 81162 0 81218 800
rect 81806 0 81862 800
rect 82450 0 82506 800
rect 83094 0 83150 800
rect 84382 0 84438 800
rect 85026 0 85082 800
rect 85670 0 85726 800
rect 86314 0 86370 800
rect 86958 0 87014 800
rect 88246 0 88302 800
rect 88890 0 88946 800
rect 89534 0 89590 800
rect 90178 0 90234 800
rect 90822 0 90878 800
rect 91466 0 91522 800
rect 92754 0 92810 800
rect 93398 0 93454 800
rect 94042 0 94098 800
rect 94686 0 94742 800
rect 95330 0 95386 800
rect 95974 0 96030 800
rect 97262 0 97318 800
rect 97906 0 97962 800
rect 98550 0 98606 800
rect 99194 0 99250 800
rect 99838 0 99894 800
rect 101126 0 101182 800
rect 101770 0 101826 800
rect 102414 0 102470 800
rect 103058 0 103114 800
rect 103702 0 103758 800
rect 104346 0 104402 800
rect 105634 0 105690 800
rect 106278 0 106334 800
rect 106922 0 106978 800
rect 107566 0 107622 800
rect 108210 0 108266 800
rect 109498 0 109554 800
rect 110142 0 110198 800
rect 110786 0 110842 800
rect 111430 0 111486 800
rect 112074 0 112130 800
rect 112718 0 112774 800
rect 114006 0 114062 800
rect 114650 0 114706 800
rect 115294 0 115350 800
rect 115938 0 115994 800
rect 116582 0 116638 800
rect 117870 0 117926 800
rect 118514 0 118570 800
rect 119158 0 119214 800
rect 119802 0 119858 800
rect 120446 0 120502 800
rect 121090 0 121146 800
rect 122378 0 122434 800
rect 123022 0 123078 800
rect 123666 0 123722 800
rect 124310 0 124366 800
rect 124954 0 125010 800
rect 126242 0 126298 800
rect 126886 0 126942 800
rect 127530 0 127586 800
rect 128174 0 128230 800
rect 128818 0 128874 800
rect 129462 0 129518 800
rect 130750 0 130806 800
rect 131394 0 131450 800
rect 132038 0 132094 800
rect 132682 0 132738 800
rect 133326 0 133382 800
rect 134614 0 134670 800
rect 135258 0 135314 800
rect 135902 0 135958 800
rect 136546 0 136602 800
rect 137190 0 137246 800
rect 137834 0 137890 800
rect 139122 0 139178 800
rect 139766 0 139822 800
rect 140410 0 140466 800
rect 141054 0 141110 800
rect 141698 0 141754 800
rect 142986 0 143042 800
rect 143630 0 143686 800
rect 144274 0 144330 800
rect 144918 0 144974 800
rect 145562 0 145618 800
rect 146206 0 146262 800
rect 147494 0 147550 800
rect 148138 0 148194 800
rect 148782 0 148838 800
rect 149426 0 149482 800
rect 150070 0 150126 800
rect 151358 0 151414 800
rect 152002 0 152058 800
rect 152646 0 152702 800
rect 153290 0 153346 800
rect 153934 0 153990 800
rect 154578 0 154634 800
rect 155866 0 155922 800
rect 156510 0 156566 800
rect 157154 0 157210 800
rect 157798 0 157854 800
rect 158442 0 158498 800
rect 159730 0 159786 800
rect 160374 0 160430 800
rect 161018 0 161074 800
rect 161662 0 161718 800
rect 162306 0 162362 800
rect 162950 0 163006 800
rect 164238 0 164294 800
rect 164882 0 164938 800
rect 165526 0 165582 800
rect 166170 0 166226 800
rect 166814 0 166870 800
rect 168102 0 168158 800
rect 168746 0 168802 800
rect 169390 0 169446 800
rect 170034 0 170090 800
rect 170678 0 170734 800
rect 171322 0 171378 800
rect 172610 0 172666 800
rect 173254 0 173310 800
rect 173898 0 173954 800
rect 174542 0 174598 800
rect 175186 0 175242 800
rect 176474 0 176530 800
rect 177118 0 177174 800
rect 177762 0 177818 800
rect 178406 0 178462 800
rect 179050 0 179106 800
rect 179694 0 179750 800
rect 180982 0 181038 800
rect 181626 0 181682 800
rect 182270 0 182326 800
rect 182914 0 182970 800
rect 183558 0 183614 800
rect 184202 0 184258 800
rect 185490 0 185546 800
rect 186134 0 186190 800
rect 186778 0 186834 800
rect 187422 0 187478 800
rect 188066 0 188122 800
rect 189354 0 189410 800
rect 189998 0 190054 800
rect 190642 0 190698 800
rect 191286 0 191342 800
rect 191930 0 191986 800
rect 192574 0 192630 800
rect 193862 0 193918 800
rect 194506 0 194562 800
rect 195150 0 195206 800
rect 195794 0 195850 800
rect 196438 0 196494 800
rect 197726 0 197782 800
rect 198370 0 198426 800
rect 199014 0 199070 800
rect 199658 0 199714 800
rect 200302 0 200358 800
rect 200946 0 201002 800
rect 202234 0 202290 800
rect 202878 0 202934 800
rect 203522 0 203578 800
rect 204166 0 204222 800
rect 204810 0 204866 800
rect 206098 0 206154 800
rect 206742 0 206798 800
rect 207386 0 207442 800
rect 208030 0 208086 800
rect 208674 0 208730 800
rect 209318 0 209374 800
rect 210606 0 210662 800
rect 211250 0 211306 800
rect 211894 0 211950 800
rect 212538 0 212594 800
rect 213182 0 213238 800
rect 214470 0 214526 800
rect 215114 0 215170 800
rect 215758 0 215814 800
rect 216402 0 216458 800
rect 217046 0 217102 800
rect 217690 0 217746 800
rect 218978 0 219034 800
rect 219622 0 219678 800
rect 220266 0 220322 800
rect 220910 0 220966 800
rect 221554 0 221610 800
rect 222842 0 222898 800
rect 223486 0 223542 800
rect 224130 0 224186 800
rect 224774 0 224830 800
rect 225418 0 225474 800
rect 226062 0 226118 800
rect 227350 0 227406 800
rect 227994 0 228050 800
rect 228638 0 228694 800
rect 229282 0 229338 800
rect 229926 0 229982 800
rect 231214 0 231270 800
rect 231858 0 231914 800
rect 232502 0 232558 800
rect 233146 0 233202 800
rect 233790 0 233846 800
rect 234434 0 234490 800
rect 235722 0 235778 800
rect 236366 0 236422 800
rect 237010 0 237066 800
rect 237654 0 237710 800
rect 238298 0 238354 800
rect 239586 0 239642 800
rect 240230 0 240286 800
rect 240874 0 240930 800
rect 241518 0 241574 800
rect 242162 0 242218 800
rect 242806 0 242862 800
rect 244094 0 244150 800
rect 244738 0 244794 800
rect 245382 0 245438 800
rect 246026 0 246082 800
rect 246670 0 246726 800
rect 247958 0 248014 800
rect 248602 0 248658 800
rect 249246 0 249302 800
rect 249890 0 249946 800
rect 250534 0 250590 800
rect 251178 0 251234 800
rect 252466 0 252522 800
rect 253110 0 253166 800
rect 253754 0 253810 800
rect 254398 0 254454 800
rect 255042 0 255098 800
rect 256330 0 256386 800
rect 256974 0 257030 800
rect 257618 0 257674 800
rect 258262 0 258318 800
rect 258906 0 258962 800
rect 259550 0 259606 800
rect 260838 0 260894 800
rect 261482 0 261538 800
rect 262126 0 262182 800
rect 262770 0 262826 800
rect 263414 0 263470 800
rect 264702 0 264758 800
rect 265346 0 265402 800
rect 265990 0 266046 800
rect 266634 0 266690 800
rect 267278 0 267334 800
rect 267922 0 267978 800
rect 269210 0 269266 800
rect 269854 0 269910 800
rect 270498 0 270554 800
rect 271142 0 271198 800
rect 271786 0 271842 800
rect 273074 0 273130 800
rect 273718 0 273774 800
rect 274362 0 274418 800
rect 275006 0 275062 800
rect 275650 0 275706 800
rect 276294 0 276350 800
rect 277582 0 277638 800
rect 278226 0 278282 800
rect 278870 0 278926 800
rect 279514 0 279570 800
rect 280158 0 280214 800
rect 280802 0 280858 800
rect 282090 0 282146 800
rect 282734 0 282790 800
rect 283378 0 283434 800
rect 284022 0 284078 800
rect 284666 0 284722 800
rect 285954 0 286010 800
rect 286598 0 286654 800
rect 287242 0 287298 800
rect 287886 0 287942 800
rect 288530 0 288586 800
rect 289174 0 289230 800
rect 290462 0 290518 800
rect 291106 0 291162 800
rect 291750 0 291806 800
rect 292394 0 292450 800
rect 293038 0 293094 800
rect 294326 0 294382 800
rect 294970 0 295026 800
rect 295614 0 295670 800
rect 296258 0 296314 800
rect 296902 0 296958 800
rect 297546 0 297602 800
rect 298834 0 298890 800
rect 299478 0 299534 800
rect 300122 0 300178 800
rect 300766 0 300822 800
rect 301410 0 301466 800
rect 302698 0 302754 800
rect 303342 0 303398 800
rect 303986 0 304042 800
rect 304630 0 304686 800
rect 305274 0 305330 800
rect 305918 0 305974 800
rect 307206 0 307262 800
rect 307850 0 307906 800
rect 308494 0 308550 800
rect 309138 0 309194 800
rect 309782 0 309838 800
rect 311070 0 311126 800
rect 311714 0 311770 800
rect 312358 0 312414 800
rect 313002 0 313058 800
rect 313646 0 313702 800
rect 314290 0 314346 800
rect 315578 0 315634 800
rect 316222 0 316278 800
rect 316866 0 316922 800
rect 317510 0 317566 800
rect 318154 0 318210 800
rect 319442 0 319498 800
rect 320086 0 320142 800
rect 320730 0 320786 800
rect 321374 0 321430 800
rect 322018 0 322074 800
rect 322662 0 322718 800
rect 323950 0 324006 800
rect 324594 0 324650 800
rect 325238 0 325294 800
rect 325882 0 325938 800
rect 326526 0 326582 800
rect 327814 0 327870 800
rect 328458 0 328514 800
rect 329102 0 329158 800
rect 329746 0 329802 800
rect 330390 0 330446 800
rect 331034 0 331090 800
rect 332322 0 332378 800
rect 332966 0 333022 800
rect 333610 0 333666 800
rect 334254 0 334310 800
rect 334898 0 334954 800
rect 336186 0 336242 800
rect 336830 0 336886 800
rect 337474 0 337530 800
rect 338118 0 338174 800
rect 338762 0 338818 800
rect 339406 0 339462 800
rect 340694 0 340750 800
rect 341338 0 341394 800
rect 341982 0 342038 800
rect 342626 0 342682 800
rect 343270 0 343326 800
rect 344558 0 344614 800
rect 345202 0 345258 800
rect 345846 0 345902 800
rect 346490 0 346546 800
rect 347134 0 347190 800
rect 347778 0 347834 800
rect 349066 0 349122 800
rect 349710 0 349766 800
rect 350354 0 350410 800
rect 350998 0 351054 800
rect 351642 0 351698 800
rect 352930 0 352986 800
rect 353574 0 353630 800
rect 354218 0 354274 800
rect 354862 0 354918 800
rect 355506 0 355562 800
rect 356150 0 356206 800
rect 357438 0 357494 800
rect 358082 0 358138 800
rect 358726 0 358782 800
rect 359370 0 359426 800
rect 360014 0 360070 800
rect 361302 0 361358 800
rect 361946 0 362002 800
rect 362590 0 362646 800
rect 363234 0 363290 800
rect 363878 0 363934 800
rect 364522 0 364578 800
rect 365810 0 365866 800
rect 366454 0 366510 800
rect 367098 0 367154 800
rect 367742 0 367798 800
rect 368386 0 368442 800
rect 369030 0 369086 800
rect 370318 0 370374 800
rect 370962 0 371018 800
rect 371606 0 371662 800
rect 372250 0 372306 800
rect 372894 0 372950 800
rect 374182 0 374238 800
rect 374826 0 374882 800
rect 375470 0 375526 800
rect 376114 0 376170 800
rect 376758 0 376814 800
rect 377402 0 377458 800
rect 378690 0 378746 800
rect 379334 0 379390 800
rect 379978 0 380034 800
rect 380622 0 380678 800
rect 381266 0 381322 800
rect 382554 0 382610 800
rect 383198 0 383254 800
rect 383842 0 383898 800
rect 384486 0 384542 800
rect 385130 0 385186 800
rect 385774 0 385830 800
rect 387062 0 387118 800
rect 387706 0 387762 800
rect 388350 0 388406 800
rect 388994 0 389050 800
rect 389638 0 389694 800
rect 390926 0 390982 800
rect 391570 0 391626 800
rect 392214 0 392270 800
rect 392858 0 392914 800
rect 393502 0 393558 800
rect 394146 0 394202 800
rect 395434 0 395490 800
rect 396078 0 396134 800
rect 396722 0 396778 800
rect 397366 0 397422 800
rect 398010 0 398066 800
rect 399298 0 399354 800
rect 399942 0 399998 800
rect 400586 0 400642 800
rect 401230 0 401286 800
rect 401874 0 401930 800
rect 402518 0 402574 800
rect 403806 0 403862 800
rect 404450 0 404506 800
rect 405094 0 405150 800
rect 405738 0 405794 800
rect 406382 0 406438 800
rect 407670 0 407726 800
rect 408314 0 408370 800
rect 408958 0 409014 800
rect 409602 0 409658 800
rect 410246 0 410302 800
rect 410890 0 410946 800
rect 412178 0 412234 800
rect 412822 0 412878 800
rect 413466 0 413522 800
rect 414110 0 414166 800
rect 414754 0 414810 800
rect 416042 0 416098 800
rect 416686 0 416742 800
rect 417330 0 417386 800
rect 417974 0 418030 800
rect 418618 0 418674 800
rect 419262 0 419318 800
rect 420550 0 420606 800
rect 421194 0 421250 800
rect 421838 0 421894 800
rect 422482 0 422538 800
rect 423126 0 423182 800
rect 424414 0 424470 800
rect 425058 0 425114 800
rect 425702 0 425758 800
rect 426346 0 426402 800
rect 426990 0 427046 800
rect 427634 0 427690 800
rect 428922 0 428978 800
rect 429566 0 429622 800
rect 430210 0 430266 800
rect 430854 0 430910 800
rect 431498 0 431554 800
rect 432786 0 432842 800
rect 433430 0 433486 800
rect 434074 0 434130 800
rect 434718 0 434774 800
rect 435362 0 435418 800
rect 436006 0 436062 800
rect 437294 0 437350 800
rect 437938 0 437994 800
rect 438582 0 438638 800
rect 439226 0 439282 800
rect 439870 0 439926 800
rect 441158 0 441214 800
rect 441802 0 441858 800
rect 442446 0 442502 800
rect 443090 0 443146 800
rect 443734 0 443790 800
rect 444378 0 444434 800
rect 445666 0 445722 800
rect 446310 0 446366 800
rect 446954 0 447010 800
rect 447598 0 447654 800
rect 448242 0 448298 800
rect 449530 0 449586 800
rect 450174 0 450230 800
rect 450818 0 450874 800
rect 451462 0 451518 800
rect 452106 0 452162 800
rect 452750 0 452806 800
rect 454038 0 454094 800
rect 454682 0 454738 800
rect 455326 0 455382 800
rect 455970 0 456026 800
rect 456614 0 456670 800
rect 457258 0 457314 800
rect 458546 0 458602 800
rect 459190 0 459246 800
rect 459834 0 459890 800
rect 460478 0 460534 800
rect 461122 0 461178 800
rect 462410 0 462466 800
rect 463054 0 463110 800
rect 463698 0 463754 800
rect 464342 0 464398 800
rect 464986 0 465042 800
rect 465630 0 465686 800
rect 466918 0 466974 800
rect 467562 0 467618 800
rect 468206 0 468262 800
rect 468850 0 468906 800
rect 469494 0 469550 800
rect 470782 0 470838 800
rect 471426 0 471482 800
rect 472070 0 472126 800
rect 472714 0 472770 800
rect 473358 0 473414 800
rect 474002 0 474058 800
rect 475290 0 475346 800
rect 475934 0 475990 800
rect 476578 0 476634 800
rect 477222 0 477278 800
rect 477866 0 477922 800
rect 479154 0 479210 800
rect 479798 0 479854 800
<< obsm2 >>
rect 130 119144 606 119785
rect 774 119144 1250 119785
rect 1418 119144 1894 119785
rect 2062 119144 2538 119785
rect 2706 119144 3826 119785
rect 3994 119144 4470 119785
rect 4638 119144 5114 119785
rect 5282 119144 5758 119785
rect 5926 119144 6402 119785
rect 6570 119144 7046 119785
rect 7214 119144 8334 119785
rect 8502 119144 8978 119785
rect 9146 119144 9622 119785
rect 9790 119144 10266 119785
rect 10434 119144 10910 119785
rect 11078 119144 12198 119785
rect 12366 119144 12842 119785
rect 13010 119144 13486 119785
rect 13654 119144 14130 119785
rect 14298 119144 14774 119785
rect 14942 119144 15418 119785
rect 15586 119144 16706 119785
rect 16874 119144 17350 119785
rect 17518 119144 17994 119785
rect 18162 119144 18638 119785
rect 18806 119144 19282 119785
rect 19450 119144 20570 119785
rect 20738 119144 21214 119785
rect 21382 119144 21858 119785
rect 22026 119144 22502 119785
rect 22670 119144 23146 119785
rect 23314 119144 23790 119785
rect 23958 119144 25078 119785
rect 25246 119144 25722 119785
rect 25890 119144 26366 119785
rect 26534 119144 27010 119785
rect 27178 119144 27654 119785
rect 27822 119144 28942 119785
rect 29110 119144 29586 119785
rect 29754 119144 30230 119785
rect 30398 119144 30874 119785
rect 31042 119144 31518 119785
rect 31686 119144 32162 119785
rect 32330 119144 33450 119785
rect 33618 119144 34094 119785
rect 34262 119144 34738 119785
rect 34906 119144 35382 119785
rect 35550 119144 36026 119785
rect 36194 119144 37314 119785
rect 37482 119144 37958 119785
rect 38126 119144 38602 119785
rect 38770 119144 39246 119785
rect 39414 119144 39890 119785
rect 40058 119144 40534 119785
rect 40702 119144 41822 119785
rect 41990 119144 42466 119785
rect 42634 119144 43110 119785
rect 43278 119144 43754 119785
rect 43922 119144 44398 119785
rect 44566 119144 45686 119785
rect 45854 119144 46330 119785
rect 46498 119144 46974 119785
rect 47142 119144 47618 119785
rect 47786 119144 48262 119785
rect 48430 119144 48906 119785
rect 49074 119144 50194 119785
rect 50362 119144 50838 119785
rect 51006 119144 51482 119785
rect 51650 119144 52126 119785
rect 52294 119144 52770 119785
rect 52938 119144 54058 119785
rect 54226 119144 54702 119785
rect 54870 119144 55346 119785
rect 55514 119144 55990 119785
rect 56158 119144 56634 119785
rect 56802 119144 57278 119785
rect 57446 119144 58566 119785
rect 58734 119144 59210 119785
rect 59378 119144 59854 119785
rect 60022 119144 60498 119785
rect 60666 119144 61142 119785
rect 61310 119144 62430 119785
rect 62598 119144 63074 119785
rect 63242 119144 63718 119785
rect 63886 119144 64362 119785
rect 64530 119144 65006 119785
rect 65174 119144 65650 119785
rect 65818 119144 66938 119785
rect 67106 119144 67582 119785
rect 67750 119144 68226 119785
rect 68394 119144 68870 119785
rect 69038 119144 69514 119785
rect 69682 119144 70158 119785
rect 70326 119144 71446 119785
rect 71614 119144 72090 119785
rect 72258 119144 72734 119785
rect 72902 119144 73378 119785
rect 73546 119144 74022 119785
rect 74190 119144 75310 119785
rect 75478 119144 75954 119785
rect 76122 119144 76598 119785
rect 76766 119144 77242 119785
rect 77410 119144 77886 119785
rect 78054 119144 78530 119785
rect 78698 119144 79818 119785
rect 79986 119144 80462 119785
rect 80630 119144 81106 119785
rect 81274 119144 81750 119785
rect 81918 119144 82394 119785
rect 82562 119144 83682 119785
rect 83850 119144 84326 119785
rect 84494 119144 84970 119785
rect 85138 119144 85614 119785
rect 85782 119144 86258 119785
rect 86426 119144 86902 119785
rect 87070 119144 88190 119785
rect 88358 119144 88834 119785
rect 89002 119144 89478 119785
rect 89646 119144 90122 119785
rect 90290 119144 90766 119785
rect 90934 119144 92054 119785
rect 92222 119144 92698 119785
rect 92866 119144 93342 119785
rect 93510 119144 93986 119785
rect 94154 119144 94630 119785
rect 94798 119144 95274 119785
rect 95442 119144 96562 119785
rect 96730 119144 97206 119785
rect 97374 119144 97850 119785
rect 98018 119144 98494 119785
rect 98662 119144 99138 119785
rect 99306 119144 100426 119785
rect 100594 119144 101070 119785
rect 101238 119144 101714 119785
rect 101882 119144 102358 119785
rect 102526 119144 103002 119785
rect 103170 119144 103646 119785
rect 103814 119144 104934 119785
rect 105102 119144 105578 119785
rect 105746 119144 106222 119785
rect 106390 119144 106866 119785
rect 107034 119144 107510 119785
rect 107678 119144 108798 119785
rect 108966 119144 109442 119785
rect 109610 119144 110086 119785
rect 110254 119144 110730 119785
rect 110898 119144 111374 119785
rect 111542 119144 112018 119785
rect 112186 119144 113306 119785
rect 113474 119144 113950 119785
rect 114118 119144 114594 119785
rect 114762 119144 115238 119785
rect 115406 119144 115882 119785
rect 116050 119144 117170 119785
rect 117338 119144 117814 119785
rect 117982 119144 118458 119785
rect 118626 119144 119102 119785
rect 119270 119144 119746 119785
rect 119914 119144 120390 119785
rect 120558 119144 121678 119785
rect 121846 119144 122322 119785
rect 122490 119144 122966 119785
rect 123134 119144 123610 119785
rect 123778 119144 124254 119785
rect 124422 119144 125542 119785
rect 125710 119144 126186 119785
rect 126354 119144 126830 119785
rect 126998 119144 127474 119785
rect 127642 119144 128118 119785
rect 128286 119144 128762 119785
rect 128930 119144 130050 119785
rect 130218 119144 130694 119785
rect 130862 119144 131338 119785
rect 131506 119144 131982 119785
rect 132150 119144 132626 119785
rect 132794 119144 133914 119785
rect 134082 119144 134558 119785
rect 134726 119144 135202 119785
rect 135370 119144 135846 119785
rect 136014 119144 136490 119785
rect 136658 119144 137134 119785
rect 137302 119144 138422 119785
rect 138590 119144 139066 119785
rect 139234 119144 139710 119785
rect 139878 119144 140354 119785
rect 140522 119144 140998 119785
rect 141166 119144 142286 119785
rect 142454 119144 142930 119785
rect 143098 119144 143574 119785
rect 143742 119144 144218 119785
rect 144386 119144 144862 119785
rect 145030 119144 145506 119785
rect 145674 119144 146794 119785
rect 146962 119144 147438 119785
rect 147606 119144 148082 119785
rect 148250 119144 148726 119785
rect 148894 119144 149370 119785
rect 149538 119144 150658 119785
rect 150826 119144 151302 119785
rect 151470 119144 151946 119785
rect 152114 119144 152590 119785
rect 152758 119144 153234 119785
rect 153402 119144 153878 119785
rect 154046 119144 155166 119785
rect 155334 119144 155810 119785
rect 155978 119144 156454 119785
rect 156622 119144 157098 119785
rect 157266 119144 157742 119785
rect 157910 119144 159030 119785
rect 159198 119144 159674 119785
rect 159842 119144 160318 119785
rect 160486 119144 160962 119785
rect 161130 119144 161606 119785
rect 161774 119144 162250 119785
rect 162418 119144 163538 119785
rect 163706 119144 164182 119785
rect 164350 119144 164826 119785
rect 164994 119144 165470 119785
rect 165638 119144 166114 119785
rect 166282 119144 166758 119785
rect 166926 119144 168046 119785
rect 168214 119144 168690 119785
rect 168858 119144 169334 119785
rect 169502 119144 169978 119785
rect 170146 119144 170622 119785
rect 170790 119144 171910 119785
rect 172078 119144 172554 119785
rect 172722 119144 173198 119785
rect 173366 119144 173842 119785
rect 174010 119144 174486 119785
rect 174654 119144 175130 119785
rect 175298 119144 176418 119785
rect 176586 119144 177062 119785
rect 177230 119144 177706 119785
rect 177874 119144 178350 119785
rect 178518 119144 178994 119785
rect 179162 119144 180282 119785
rect 180450 119144 180926 119785
rect 181094 119144 181570 119785
rect 181738 119144 182214 119785
rect 182382 119144 182858 119785
rect 183026 119144 183502 119785
rect 183670 119144 184790 119785
rect 184958 119144 185434 119785
rect 185602 119144 186078 119785
rect 186246 119144 186722 119785
rect 186890 119144 187366 119785
rect 187534 119144 188654 119785
rect 188822 119144 189298 119785
rect 189466 119144 189942 119785
rect 190110 119144 190586 119785
rect 190754 119144 191230 119785
rect 191398 119144 191874 119785
rect 192042 119144 193162 119785
rect 193330 119144 193806 119785
rect 193974 119144 194450 119785
rect 194618 119144 195094 119785
rect 195262 119144 195738 119785
rect 195906 119144 197026 119785
rect 197194 119144 197670 119785
rect 197838 119144 198314 119785
rect 198482 119144 198958 119785
rect 199126 119144 199602 119785
rect 199770 119144 200246 119785
rect 200414 119144 201534 119785
rect 201702 119144 202178 119785
rect 202346 119144 202822 119785
rect 202990 119144 203466 119785
rect 203634 119144 204110 119785
rect 204278 119144 205398 119785
rect 205566 119144 206042 119785
rect 206210 119144 206686 119785
rect 206854 119144 207330 119785
rect 207498 119144 207974 119785
rect 208142 119144 208618 119785
rect 208786 119144 209906 119785
rect 210074 119144 210550 119785
rect 210718 119144 211194 119785
rect 211362 119144 211838 119785
rect 212006 119144 212482 119785
rect 212650 119144 213770 119785
rect 213938 119144 214414 119785
rect 214582 119144 215058 119785
rect 215226 119144 215702 119785
rect 215870 119144 216346 119785
rect 216514 119144 216990 119785
rect 217158 119144 218278 119785
rect 218446 119144 218922 119785
rect 219090 119144 219566 119785
rect 219734 119144 220210 119785
rect 220378 119144 220854 119785
rect 221022 119144 222142 119785
rect 222310 119144 222786 119785
rect 222954 119144 223430 119785
rect 223598 119144 224074 119785
rect 224242 119144 224718 119785
rect 224886 119144 225362 119785
rect 225530 119144 226650 119785
rect 226818 119144 227294 119785
rect 227462 119144 227938 119785
rect 228106 119144 228582 119785
rect 228750 119144 229226 119785
rect 229394 119144 230514 119785
rect 230682 119144 231158 119785
rect 231326 119144 231802 119785
rect 231970 119144 232446 119785
rect 232614 119144 233090 119785
rect 233258 119144 233734 119785
rect 233902 119144 235022 119785
rect 235190 119144 235666 119785
rect 235834 119144 236310 119785
rect 236478 119144 236954 119785
rect 237122 119144 237598 119785
rect 237766 119144 238886 119785
rect 239054 119144 239530 119785
rect 239698 119144 240174 119785
rect 240342 119144 240818 119785
rect 240986 119144 241462 119785
rect 241630 119144 242106 119785
rect 242274 119144 243394 119785
rect 243562 119144 244038 119785
rect 244206 119144 244682 119785
rect 244850 119144 245326 119785
rect 245494 119144 245970 119785
rect 246138 119144 247258 119785
rect 247426 119144 247902 119785
rect 248070 119144 248546 119785
rect 248714 119144 249190 119785
rect 249358 119144 249834 119785
rect 250002 119144 250478 119785
rect 250646 119144 251766 119785
rect 251934 119144 252410 119785
rect 252578 119144 253054 119785
rect 253222 119144 253698 119785
rect 253866 119144 254342 119785
rect 254510 119144 254986 119785
rect 255154 119144 256274 119785
rect 256442 119144 256918 119785
rect 257086 119144 257562 119785
rect 257730 119144 258206 119785
rect 258374 119144 258850 119785
rect 259018 119144 260138 119785
rect 260306 119144 260782 119785
rect 260950 119144 261426 119785
rect 261594 119144 262070 119785
rect 262238 119144 262714 119785
rect 262882 119144 263358 119785
rect 263526 119144 264646 119785
rect 264814 119144 265290 119785
rect 265458 119144 265934 119785
rect 266102 119144 266578 119785
rect 266746 119144 267222 119785
rect 267390 119144 268510 119785
rect 268678 119144 269154 119785
rect 269322 119144 269798 119785
rect 269966 119144 270442 119785
rect 270610 119144 271086 119785
rect 271254 119144 271730 119785
rect 271898 119144 273018 119785
rect 273186 119144 273662 119785
rect 273830 119144 274306 119785
rect 274474 119144 274950 119785
rect 275118 119144 275594 119785
rect 275762 119144 276882 119785
rect 277050 119144 277526 119785
rect 277694 119144 278170 119785
rect 278338 119144 278814 119785
rect 278982 119144 279458 119785
rect 279626 119144 280102 119785
rect 280270 119144 281390 119785
rect 281558 119144 282034 119785
rect 282202 119144 282678 119785
rect 282846 119144 283322 119785
rect 283490 119144 283966 119785
rect 284134 119144 285254 119785
rect 285422 119144 285898 119785
rect 286066 119144 286542 119785
rect 286710 119144 287186 119785
rect 287354 119144 287830 119785
rect 287998 119144 288474 119785
rect 288642 119144 289762 119785
rect 289930 119144 290406 119785
rect 290574 119144 291050 119785
rect 291218 119144 291694 119785
rect 291862 119144 292338 119785
rect 292506 119144 293626 119785
rect 293794 119144 294270 119785
rect 294438 119144 294914 119785
rect 295082 119144 295558 119785
rect 295726 119144 296202 119785
rect 296370 119144 296846 119785
rect 297014 119144 298134 119785
rect 298302 119144 298778 119785
rect 298946 119144 299422 119785
rect 299590 119144 300066 119785
rect 300234 119144 300710 119785
rect 300878 119144 301998 119785
rect 302166 119144 302642 119785
rect 302810 119144 303286 119785
rect 303454 119144 303930 119785
rect 304098 119144 304574 119785
rect 304742 119144 305218 119785
rect 305386 119144 306506 119785
rect 306674 119144 307150 119785
rect 307318 119144 307794 119785
rect 307962 119144 308438 119785
rect 308606 119144 309082 119785
rect 309250 119144 310370 119785
rect 310538 119144 311014 119785
rect 311182 119144 311658 119785
rect 311826 119144 312302 119785
rect 312470 119144 312946 119785
rect 313114 119144 313590 119785
rect 313758 119144 314878 119785
rect 315046 119144 315522 119785
rect 315690 119144 316166 119785
rect 316334 119144 316810 119785
rect 316978 119144 317454 119785
rect 317622 119144 318742 119785
rect 318910 119144 319386 119785
rect 319554 119144 320030 119785
rect 320198 119144 320674 119785
rect 320842 119144 321318 119785
rect 321486 119144 321962 119785
rect 322130 119144 323250 119785
rect 323418 119144 323894 119785
rect 324062 119144 324538 119785
rect 324706 119144 325182 119785
rect 325350 119144 325826 119785
rect 325994 119144 327114 119785
rect 327282 119144 327758 119785
rect 327926 119144 328402 119785
rect 328570 119144 329046 119785
rect 329214 119144 329690 119785
rect 329858 119144 330334 119785
rect 330502 119144 331622 119785
rect 331790 119144 332266 119785
rect 332434 119144 332910 119785
rect 333078 119144 333554 119785
rect 333722 119144 334198 119785
rect 334366 119144 335486 119785
rect 335654 119144 336130 119785
rect 336298 119144 336774 119785
rect 336942 119144 337418 119785
rect 337586 119144 338062 119785
rect 338230 119144 338706 119785
rect 338874 119144 339994 119785
rect 340162 119144 340638 119785
rect 340806 119144 341282 119785
rect 341450 119144 341926 119785
rect 342094 119144 342570 119785
rect 342738 119144 343214 119785
rect 343382 119144 344502 119785
rect 344670 119144 345146 119785
rect 345314 119144 345790 119785
rect 345958 119144 346434 119785
rect 346602 119144 347078 119785
rect 347246 119144 348366 119785
rect 348534 119144 349010 119785
rect 349178 119144 349654 119785
rect 349822 119144 350298 119785
rect 350466 119144 350942 119785
rect 351110 119144 351586 119785
rect 351754 119144 352874 119785
rect 353042 119144 353518 119785
rect 353686 119144 354162 119785
rect 354330 119144 354806 119785
rect 354974 119144 355450 119785
rect 355618 119144 356738 119785
rect 356906 119144 357382 119785
rect 357550 119144 358026 119785
rect 358194 119144 358670 119785
rect 358838 119144 359314 119785
rect 359482 119144 359958 119785
rect 360126 119144 361246 119785
rect 361414 119144 361890 119785
rect 362058 119144 362534 119785
rect 362702 119144 363178 119785
rect 363346 119144 363822 119785
rect 363990 119144 365110 119785
rect 365278 119144 365754 119785
rect 365922 119144 366398 119785
rect 366566 119144 367042 119785
rect 367210 119144 367686 119785
rect 367854 119144 368330 119785
rect 368498 119144 369618 119785
rect 369786 119144 370262 119785
rect 370430 119144 370906 119785
rect 371074 119144 371550 119785
rect 371718 119144 372194 119785
rect 372362 119144 373482 119785
rect 373650 119144 374126 119785
rect 374294 119144 374770 119785
rect 374938 119144 375414 119785
rect 375582 119144 376058 119785
rect 376226 119144 376702 119785
rect 376870 119144 377990 119785
rect 378158 119144 378634 119785
rect 378802 119144 379278 119785
rect 379446 119144 379922 119785
rect 380090 119144 380566 119785
rect 380734 119144 381854 119785
rect 382022 119144 382498 119785
rect 382666 119144 383142 119785
rect 383310 119144 383786 119785
rect 383954 119144 384430 119785
rect 384598 119144 385074 119785
rect 385242 119144 386362 119785
rect 386530 119144 387006 119785
rect 387174 119144 387650 119785
rect 387818 119144 388294 119785
rect 388462 119144 388938 119785
rect 389106 119144 390226 119785
rect 390394 119144 390870 119785
rect 391038 119144 391514 119785
rect 391682 119144 392158 119785
rect 392326 119144 392802 119785
rect 392970 119144 393446 119785
rect 393614 119144 394734 119785
rect 394902 119144 395378 119785
rect 395546 119144 396022 119785
rect 396190 119144 396666 119785
rect 396834 119144 397310 119785
rect 397478 119144 398598 119785
rect 398766 119144 399242 119785
rect 399410 119144 399886 119785
rect 400054 119144 400530 119785
rect 400698 119144 401174 119785
rect 401342 119144 401818 119785
rect 401986 119144 403106 119785
rect 403274 119144 403750 119785
rect 403918 119144 404394 119785
rect 404562 119144 405038 119785
rect 405206 119144 405682 119785
rect 405850 119144 406970 119785
rect 407138 119144 407614 119785
rect 407782 119144 408258 119785
rect 408426 119144 408902 119785
rect 409070 119144 409546 119785
rect 409714 119144 410190 119785
rect 410358 119144 411478 119785
rect 411646 119144 412122 119785
rect 412290 119144 412766 119785
rect 412934 119144 413410 119785
rect 413578 119144 414054 119785
rect 414222 119144 415342 119785
rect 415510 119144 415986 119785
rect 416154 119144 416630 119785
rect 416798 119144 417274 119785
rect 417442 119144 417918 119785
rect 418086 119144 418562 119785
rect 418730 119144 419850 119785
rect 420018 119144 420494 119785
rect 420662 119144 421138 119785
rect 421306 119144 421782 119785
rect 421950 119144 422426 119785
rect 422594 119144 423714 119785
rect 423882 119144 424358 119785
rect 424526 119144 425002 119785
rect 425170 119144 425646 119785
rect 425814 119144 426290 119785
rect 426458 119144 426934 119785
rect 427102 119144 428222 119785
rect 428390 119144 428866 119785
rect 429034 119144 429510 119785
rect 429678 119144 430154 119785
rect 430322 119144 430798 119785
rect 430966 119144 432086 119785
rect 432254 119144 432730 119785
rect 432898 119144 433374 119785
rect 433542 119144 434018 119785
rect 434186 119144 434662 119785
rect 434830 119144 435306 119785
rect 435474 119144 436594 119785
rect 436762 119144 437238 119785
rect 437406 119144 437882 119785
rect 438050 119144 438526 119785
rect 438694 119144 439170 119785
rect 439338 119144 439814 119785
rect 439982 119144 441102 119785
rect 441270 119144 441746 119785
rect 441914 119144 442390 119785
rect 442558 119144 443034 119785
rect 443202 119144 443678 119785
rect 443846 119144 444966 119785
rect 445134 119144 445610 119785
rect 445778 119144 446254 119785
rect 446422 119144 446898 119785
rect 447066 119144 447542 119785
rect 447710 119144 448186 119785
rect 448354 119144 449474 119785
rect 449642 119144 450118 119785
rect 450286 119144 450762 119785
rect 450930 119144 451406 119785
rect 451574 119144 452050 119785
rect 452218 119144 453338 119785
rect 453506 119144 453982 119785
rect 454150 119144 454626 119785
rect 454794 119144 455270 119785
rect 455438 119144 455914 119785
rect 456082 119144 456558 119785
rect 456726 119144 457846 119785
rect 458014 119144 458490 119785
rect 458658 119144 459134 119785
rect 459302 119144 459778 119785
rect 459946 119144 460422 119785
rect 460590 119144 461710 119785
rect 461878 119144 462354 119785
rect 462522 119144 462998 119785
rect 463166 119144 463642 119785
rect 463810 119144 464286 119785
rect 464454 119144 464930 119785
rect 465098 119144 466218 119785
rect 466386 119144 466862 119785
rect 467030 119144 467506 119785
rect 467674 119144 468150 119785
rect 468318 119144 468794 119785
rect 468962 119144 470082 119785
rect 470250 119144 470726 119785
rect 470894 119144 471370 119785
rect 471538 119144 472014 119785
rect 472182 119144 472658 119785
rect 472826 119144 473302 119785
rect 473470 119144 474590 119785
rect 474758 119144 475234 119785
rect 475402 119144 475878 119785
rect 476046 119144 476522 119785
rect 476690 119144 477166 119785
rect 477334 119144 478454 119785
rect 478622 119144 479098 119785
rect 479266 119144 479742 119785
rect 20 856 479852 119144
rect 130 31 606 856
rect 774 31 1250 856
rect 1418 31 1894 856
rect 2062 31 2538 856
rect 2706 31 3182 856
rect 3350 31 4470 856
rect 4638 31 5114 856
rect 5282 31 5758 856
rect 5926 31 6402 856
rect 6570 31 7046 856
rect 7214 31 7690 856
rect 7858 31 8978 856
rect 9146 31 9622 856
rect 9790 31 10266 856
rect 10434 31 10910 856
rect 11078 31 11554 856
rect 11722 31 12842 856
rect 13010 31 13486 856
rect 13654 31 14130 856
rect 14298 31 14774 856
rect 14942 31 15418 856
rect 15586 31 16062 856
rect 16230 31 17350 856
rect 17518 31 17994 856
rect 18162 31 18638 856
rect 18806 31 19282 856
rect 19450 31 19926 856
rect 20094 31 21214 856
rect 21382 31 21858 856
rect 22026 31 22502 856
rect 22670 31 23146 856
rect 23314 31 23790 856
rect 23958 31 24434 856
rect 24602 31 25722 856
rect 25890 31 26366 856
rect 26534 31 27010 856
rect 27178 31 27654 856
rect 27822 31 28298 856
rect 28466 31 29586 856
rect 29754 31 30230 856
rect 30398 31 30874 856
rect 31042 31 31518 856
rect 31686 31 32162 856
rect 32330 31 32806 856
rect 32974 31 34094 856
rect 34262 31 34738 856
rect 34906 31 35382 856
rect 35550 31 36026 856
rect 36194 31 36670 856
rect 36838 31 37958 856
rect 38126 31 38602 856
rect 38770 31 39246 856
rect 39414 31 39890 856
rect 40058 31 40534 856
rect 40702 31 41178 856
rect 41346 31 42466 856
rect 42634 31 43110 856
rect 43278 31 43754 856
rect 43922 31 44398 856
rect 44566 31 45042 856
rect 45210 31 46330 856
rect 46498 31 46974 856
rect 47142 31 47618 856
rect 47786 31 48262 856
rect 48430 31 48906 856
rect 49074 31 49550 856
rect 49718 31 50838 856
rect 51006 31 51482 856
rect 51650 31 52126 856
rect 52294 31 52770 856
rect 52938 31 53414 856
rect 53582 31 54702 856
rect 54870 31 55346 856
rect 55514 31 55990 856
rect 56158 31 56634 856
rect 56802 31 57278 856
rect 57446 31 57922 856
rect 58090 31 59210 856
rect 59378 31 59854 856
rect 60022 31 60498 856
rect 60666 31 61142 856
rect 61310 31 61786 856
rect 61954 31 63074 856
rect 63242 31 63718 856
rect 63886 31 64362 856
rect 64530 31 65006 856
rect 65174 31 65650 856
rect 65818 31 66294 856
rect 66462 31 67582 856
rect 67750 31 68226 856
rect 68394 31 68870 856
rect 69038 31 69514 856
rect 69682 31 70158 856
rect 70326 31 71446 856
rect 71614 31 72090 856
rect 72258 31 72734 856
rect 72902 31 73378 856
rect 73546 31 74022 856
rect 74190 31 74666 856
rect 74834 31 75954 856
rect 76122 31 76598 856
rect 76766 31 77242 856
rect 77410 31 77886 856
rect 78054 31 78530 856
rect 78698 31 79818 856
rect 79986 31 80462 856
rect 80630 31 81106 856
rect 81274 31 81750 856
rect 81918 31 82394 856
rect 82562 31 83038 856
rect 83206 31 84326 856
rect 84494 31 84970 856
rect 85138 31 85614 856
rect 85782 31 86258 856
rect 86426 31 86902 856
rect 87070 31 88190 856
rect 88358 31 88834 856
rect 89002 31 89478 856
rect 89646 31 90122 856
rect 90290 31 90766 856
rect 90934 31 91410 856
rect 91578 31 92698 856
rect 92866 31 93342 856
rect 93510 31 93986 856
rect 94154 31 94630 856
rect 94798 31 95274 856
rect 95442 31 95918 856
rect 96086 31 97206 856
rect 97374 31 97850 856
rect 98018 31 98494 856
rect 98662 31 99138 856
rect 99306 31 99782 856
rect 99950 31 101070 856
rect 101238 31 101714 856
rect 101882 31 102358 856
rect 102526 31 103002 856
rect 103170 31 103646 856
rect 103814 31 104290 856
rect 104458 31 105578 856
rect 105746 31 106222 856
rect 106390 31 106866 856
rect 107034 31 107510 856
rect 107678 31 108154 856
rect 108322 31 109442 856
rect 109610 31 110086 856
rect 110254 31 110730 856
rect 110898 31 111374 856
rect 111542 31 112018 856
rect 112186 31 112662 856
rect 112830 31 113950 856
rect 114118 31 114594 856
rect 114762 31 115238 856
rect 115406 31 115882 856
rect 116050 31 116526 856
rect 116694 31 117814 856
rect 117982 31 118458 856
rect 118626 31 119102 856
rect 119270 31 119746 856
rect 119914 31 120390 856
rect 120558 31 121034 856
rect 121202 31 122322 856
rect 122490 31 122966 856
rect 123134 31 123610 856
rect 123778 31 124254 856
rect 124422 31 124898 856
rect 125066 31 126186 856
rect 126354 31 126830 856
rect 126998 31 127474 856
rect 127642 31 128118 856
rect 128286 31 128762 856
rect 128930 31 129406 856
rect 129574 31 130694 856
rect 130862 31 131338 856
rect 131506 31 131982 856
rect 132150 31 132626 856
rect 132794 31 133270 856
rect 133438 31 134558 856
rect 134726 31 135202 856
rect 135370 31 135846 856
rect 136014 31 136490 856
rect 136658 31 137134 856
rect 137302 31 137778 856
rect 137946 31 139066 856
rect 139234 31 139710 856
rect 139878 31 140354 856
rect 140522 31 140998 856
rect 141166 31 141642 856
rect 141810 31 142930 856
rect 143098 31 143574 856
rect 143742 31 144218 856
rect 144386 31 144862 856
rect 145030 31 145506 856
rect 145674 31 146150 856
rect 146318 31 147438 856
rect 147606 31 148082 856
rect 148250 31 148726 856
rect 148894 31 149370 856
rect 149538 31 150014 856
rect 150182 31 151302 856
rect 151470 31 151946 856
rect 152114 31 152590 856
rect 152758 31 153234 856
rect 153402 31 153878 856
rect 154046 31 154522 856
rect 154690 31 155810 856
rect 155978 31 156454 856
rect 156622 31 157098 856
rect 157266 31 157742 856
rect 157910 31 158386 856
rect 158554 31 159674 856
rect 159842 31 160318 856
rect 160486 31 160962 856
rect 161130 31 161606 856
rect 161774 31 162250 856
rect 162418 31 162894 856
rect 163062 31 164182 856
rect 164350 31 164826 856
rect 164994 31 165470 856
rect 165638 31 166114 856
rect 166282 31 166758 856
rect 166926 31 168046 856
rect 168214 31 168690 856
rect 168858 31 169334 856
rect 169502 31 169978 856
rect 170146 31 170622 856
rect 170790 31 171266 856
rect 171434 31 172554 856
rect 172722 31 173198 856
rect 173366 31 173842 856
rect 174010 31 174486 856
rect 174654 31 175130 856
rect 175298 31 176418 856
rect 176586 31 177062 856
rect 177230 31 177706 856
rect 177874 31 178350 856
rect 178518 31 178994 856
rect 179162 31 179638 856
rect 179806 31 180926 856
rect 181094 31 181570 856
rect 181738 31 182214 856
rect 182382 31 182858 856
rect 183026 31 183502 856
rect 183670 31 184146 856
rect 184314 31 185434 856
rect 185602 31 186078 856
rect 186246 31 186722 856
rect 186890 31 187366 856
rect 187534 31 188010 856
rect 188178 31 189298 856
rect 189466 31 189942 856
rect 190110 31 190586 856
rect 190754 31 191230 856
rect 191398 31 191874 856
rect 192042 31 192518 856
rect 192686 31 193806 856
rect 193974 31 194450 856
rect 194618 31 195094 856
rect 195262 31 195738 856
rect 195906 31 196382 856
rect 196550 31 197670 856
rect 197838 31 198314 856
rect 198482 31 198958 856
rect 199126 31 199602 856
rect 199770 31 200246 856
rect 200414 31 200890 856
rect 201058 31 202178 856
rect 202346 31 202822 856
rect 202990 31 203466 856
rect 203634 31 204110 856
rect 204278 31 204754 856
rect 204922 31 206042 856
rect 206210 31 206686 856
rect 206854 31 207330 856
rect 207498 31 207974 856
rect 208142 31 208618 856
rect 208786 31 209262 856
rect 209430 31 210550 856
rect 210718 31 211194 856
rect 211362 31 211838 856
rect 212006 31 212482 856
rect 212650 31 213126 856
rect 213294 31 214414 856
rect 214582 31 215058 856
rect 215226 31 215702 856
rect 215870 31 216346 856
rect 216514 31 216990 856
rect 217158 31 217634 856
rect 217802 31 218922 856
rect 219090 31 219566 856
rect 219734 31 220210 856
rect 220378 31 220854 856
rect 221022 31 221498 856
rect 221666 31 222786 856
rect 222954 31 223430 856
rect 223598 31 224074 856
rect 224242 31 224718 856
rect 224886 31 225362 856
rect 225530 31 226006 856
rect 226174 31 227294 856
rect 227462 31 227938 856
rect 228106 31 228582 856
rect 228750 31 229226 856
rect 229394 31 229870 856
rect 230038 31 231158 856
rect 231326 31 231802 856
rect 231970 31 232446 856
rect 232614 31 233090 856
rect 233258 31 233734 856
rect 233902 31 234378 856
rect 234546 31 235666 856
rect 235834 31 236310 856
rect 236478 31 236954 856
rect 237122 31 237598 856
rect 237766 31 238242 856
rect 238410 31 239530 856
rect 239698 31 240174 856
rect 240342 31 240818 856
rect 240986 31 241462 856
rect 241630 31 242106 856
rect 242274 31 242750 856
rect 242918 31 244038 856
rect 244206 31 244682 856
rect 244850 31 245326 856
rect 245494 31 245970 856
rect 246138 31 246614 856
rect 246782 31 247902 856
rect 248070 31 248546 856
rect 248714 31 249190 856
rect 249358 31 249834 856
rect 250002 31 250478 856
rect 250646 31 251122 856
rect 251290 31 252410 856
rect 252578 31 253054 856
rect 253222 31 253698 856
rect 253866 31 254342 856
rect 254510 31 254986 856
rect 255154 31 256274 856
rect 256442 31 256918 856
rect 257086 31 257562 856
rect 257730 31 258206 856
rect 258374 31 258850 856
rect 259018 31 259494 856
rect 259662 31 260782 856
rect 260950 31 261426 856
rect 261594 31 262070 856
rect 262238 31 262714 856
rect 262882 31 263358 856
rect 263526 31 264646 856
rect 264814 31 265290 856
rect 265458 31 265934 856
rect 266102 31 266578 856
rect 266746 31 267222 856
rect 267390 31 267866 856
rect 268034 31 269154 856
rect 269322 31 269798 856
rect 269966 31 270442 856
rect 270610 31 271086 856
rect 271254 31 271730 856
rect 271898 31 273018 856
rect 273186 31 273662 856
rect 273830 31 274306 856
rect 274474 31 274950 856
rect 275118 31 275594 856
rect 275762 31 276238 856
rect 276406 31 277526 856
rect 277694 31 278170 856
rect 278338 31 278814 856
rect 278982 31 279458 856
rect 279626 31 280102 856
rect 280270 31 280746 856
rect 280914 31 282034 856
rect 282202 31 282678 856
rect 282846 31 283322 856
rect 283490 31 283966 856
rect 284134 31 284610 856
rect 284778 31 285898 856
rect 286066 31 286542 856
rect 286710 31 287186 856
rect 287354 31 287830 856
rect 287998 31 288474 856
rect 288642 31 289118 856
rect 289286 31 290406 856
rect 290574 31 291050 856
rect 291218 31 291694 856
rect 291862 31 292338 856
rect 292506 31 292982 856
rect 293150 31 294270 856
rect 294438 31 294914 856
rect 295082 31 295558 856
rect 295726 31 296202 856
rect 296370 31 296846 856
rect 297014 31 297490 856
rect 297658 31 298778 856
rect 298946 31 299422 856
rect 299590 31 300066 856
rect 300234 31 300710 856
rect 300878 31 301354 856
rect 301522 31 302642 856
rect 302810 31 303286 856
rect 303454 31 303930 856
rect 304098 31 304574 856
rect 304742 31 305218 856
rect 305386 31 305862 856
rect 306030 31 307150 856
rect 307318 31 307794 856
rect 307962 31 308438 856
rect 308606 31 309082 856
rect 309250 31 309726 856
rect 309894 31 311014 856
rect 311182 31 311658 856
rect 311826 31 312302 856
rect 312470 31 312946 856
rect 313114 31 313590 856
rect 313758 31 314234 856
rect 314402 31 315522 856
rect 315690 31 316166 856
rect 316334 31 316810 856
rect 316978 31 317454 856
rect 317622 31 318098 856
rect 318266 31 319386 856
rect 319554 31 320030 856
rect 320198 31 320674 856
rect 320842 31 321318 856
rect 321486 31 321962 856
rect 322130 31 322606 856
rect 322774 31 323894 856
rect 324062 31 324538 856
rect 324706 31 325182 856
rect 325350 31 325826 856
rect 325994 31 326470 856
rect 326638 31 327758 856
rect 327926 31 328402 856
rect 328570 31 329046 856
rect 329214 31 329690 856
rect 329858 31 330334 856
rect 330502 31 330978 856
rect 331146 31 332266 856
rect 332434 31 332910 856
rect 333078 31 333554 856
rect 333722 31 334198 856
rect 334366 31 334842 856
rect 335010 31 336130 856
rect 336298 31 336774 856
rect 336942 31 337418 856
rect 337586 31 338062 856
rect 338230 31 338706 856
rect 338874 31 339350 856
rect 339518 31 340638 856
rect 340806 31 341282 856
rect 341450 31 341926 856
rect 342094 31 342570 856
rect 342738 31 343214 856
rect 343382 31 344502 856
rect 344670 31 345146 856
rect 345314 31 345790 856
rect 345958 31 346434 856
rect 346602 31 347078 856
rect 347246 31 347722 856
rect 347890 31 349010 856
rect 349178 31 349654 856
rect 349822 31 350298 856
rect 350466 31 350942 856
rect 351110 31 351586 856
rect 351754 31 352874 856
rect 353042 31 353518 856
rect 353686 31 354162 856
rect 354330 31 354806 856
rect 354974 31 355450 856
rect 355618 31 356094 856
rect 356262 31 357382 856
rect 357550 31 358026 856
rect 358194 31 358670 856
rect 358838 31 359314 856
rect 359482 31 359958 856
rect 360126 31 361246 856
rect 361414 31 361890 856
rect 362058 31 362534 856
rect 362702 31 363178 856
rect 363346 31 363822 856
rect 363990 31 364466 856
rect 364634 31 365754 856
rect 365922 31 366398 856
rect 366566 31 367042 856
rect 367210 31 367686 856
rect 367854 31 368330 856
rect 368498 31 368974 856
rect 369142 31 370262 856
rect 370430 31 370906 856
rect 371074 31 371550 856
rect 371718 31 372194 856
rect 372362 31 372838 856
rect 373006 31 374126 856
rect 374294 31 374770 856
rect 374938 31 375414 856
rect 375582 31 376058 856
rect 376226 31 376702 856
rect 376870 31 377346 856
rect 377514 31 378634 856
rect 378802 31 379278 856
rect 379446 31 379922 856
rect 380090 31 380566 856
rect 380734 31 381210 856
rect 381378 31 382498 856
rect 382666 31 383142 856
rect 383310 31 383786 856
rect 383954 31 384430 856
rect 384598 31 385074 856
rect 385242 31 385718 856
rect 385886 31 387006 856
rect 387174 31 387650 856
rect 387818 31 388294 856
rect 388462 31 388938 856
rect 389106 31 389582 856
rect 389750 31 390870 856
rect 391038 31 391514 856
rect 391682 31 392158 856
rect 392326 31 392802 856
rect 392970 31 393446 856
rect 393614 31 394090 856
rect 394258 31 395378 856
rect 395546 31 396022 856
rect 396190 31 396666 856
rect 396834 31 397310 856
rect 397478 31 397954 856
rect 398122 31 399242 856
rect 399410 31 399886 856
rect 400054 31 400530 856
rect 400698 31 401174 856
rect 401342 31 401818 856
rect 401986 31 402462 856
rect 402630 31 403750 856
rect 403918 31 404394 856
rect 404562 31 405038 856
rect 405206 31 405682 856
rect 405850 31 406326 856
rect 406494 31 407614 856
rect 407782 31 408258 856
rect 408426 31 408902 856
rect 409070 31 409546 856
rect 409714 31 410190 856
rect 410358 31 410834 856
rect 411002 31 412122 856
rect 412290 31 412766 856
rect 412934 31 413410 856
rect 413578 31 414054 856
rect 414222 31 414698 856
rect 414866 31 415986 856
rect 416154 31 416630 856
rect 416798 31 417274 856
rect 417442 31 417918 856
rect 418086 31 418562 856
rect 418730 31 419206 856
rect 419374 31 420494 856
rect 420662 31 421138 856
rect 421306 31 421782 856
rect 421950 31 422426 856
rect 422594 31 423070 856
rect 423238 31 424358 856
rect 424526 31 425002 856
rect 425170 31 425646 856
rect 425814 31 426290 856
rect 426458 31 426934 856
rect 427102 31 427578 856
rect 427746 31 428866 856
rect 429034 31 429510 856
rect 429678 31 430154 856
rect 430322 31 430798 856
rect 430966 31 431442 856
rect 431610 31 432730 856
rect 432898 31 433374 856
rect 433542 31 434018 856
rect 434186 31 434662 856
rect 434830 31 435306 856
rect 435474 31 435950 856
rect 436118 31 437238 856
rect 437406 31 437882 856
rect 438050 31 438526 856
rect 438694 31 439170 856
rect 439338 31 439814 856
rect 439982 31 441102 856
rect 441270 31 441746 856
rect 441914 31 442390 856
rect 442558 31 443034 856
rect 443202 31 443678 856
rect 443846 31 444322 856
rect 444490 31 445610 856
rect 445778 31 446254 856
rect 446422 31 446898 856
rect 447066 31 447542 856
rect 447710 31 448186 856
rect 448354 31 449474 856
rect 449642 31 450118 856
rect 450286 31 450762 856
rect 450930 31 451406 856
rect 451574 31 452050 856
rect 452218 31 452694 856
rect 452862 31 453982 856
rect 454150 31 454626 856
rect 454794 31 455270 856
rect 455438 31 455914 856
rect 456082 31 456558 856
rect 456726 31 457202 856
rect 457370 31 458490 856
rect 458658 31 459134 856
rect 459302 31 459778 856
rect 459946 31 460422 856
rect 460590 31 461066 856
rect 461234 31 462354 856
rect 462522 31 462998 856
rect 463166 31 463642 856
rect 463810 31 464286 856
rect 464454 31 464930 856
rect 465098 31 465574 856
rect 465742 31 466862 856
rect 467030 31 467506 856
rect 467674 31 468150 856
rect 468318 31 468794 856
rect 468962 31 469438 856
rect 469606 31 470726 856
rect 470894 31 471370 856
rect 471538 31 472014 856
rect 472182 31 472658 856
rect 472826 31 473302 856
rect 473470 31 473946 856
rect 474114 31 475234 856
rect 475402 31 475878 856
rect 476046 31 476522 856
rect 476690 31 477166 856
rect 477334 31 477810 856
rect 477978 31 479098 856
rect 479266 31 479742 856
<< metal3 >>
rect 479200 119688 480000 119808
rect 0 119008 800 119128
rect 479200 119008 480000 119128
rect 0 118328 800 118448
rect 479200 118328 480000 118448
rect 0 117648 800 117768
rect 0 116968 800 117088
rect 479200 116968 480000 117088
rect 0 116288 800 116408
rect 479200 116288 480000 116408
rect 0 115608 800 115728
rect 479200 115608 480000 115728
rect 479200 114928 480000 115048
rect 0 114248 800 114368
rect 479200 114248 480000 114368
rect 0 113568 800 113688
rect 0 112888 800 113008
rect 479200 112888 480000 113008
rect 0 112208 800 112328
rect 479200 112208 480000 112328
rect 0 111528 800 111648
rect 479200 111528 480000 111648
rect 479200 110848 480000 110968
rect 0 110168 800 110288
rect 479200 110168 480000 110288
rect 0 109488 800 109608
rect 479200 109488 480000 109608
rect 0 108808 800 108928
rect 0 108128 800 108248
rect 479200 108128 480000 108248
rect 0 107448 800 107568
rect 479200 107448 480000 107568
rect 0 106768 800 106888
rect 479200 106768 480000 106888
rect 479200 106088 480000 106208
rect 0 105408 800 105528
rect 479200 105408 480000 105528
rect 0 104728 800 104848
rect 0 104048 800 104168
rect 479200 104048 480000 104168
rect 0 103368 800 103488
rect 479200 103368 480000 103488
rect 0 102688 800 102808
rect 479200 102688 480000 102808
rect 479200 102008 480000 102128
rect 0 101328 800 101448
rect 479200 101328 480000 101448
rect 0 100648 800 100768
rect 479200 100648 480000 100768
rect 0 99968 800 100088
rect 0 99288 800 99408
rect 479200 99288 480000 99408
rect 0 98608 800 98728
rect 479200 98608 480000 98728
rect 0 97928 800 98048
rect 479200 97928 480000 98048
rect 479200 97248 480000 97368
rect 0 96568 800 96688
rect 479200 96568 480000 96688
rect 0 95888 800 96008
rect 0 95208 800 95328
rect 479200 95208 480000 95328
rect 0 94528 800 94648
rect 479200 94528 480000 94648
rect 0 93848 800 93968
rect 479200 93848 480000 93968
rect 0 93168 800 93288
rect 479200 93168 480000 93288
rect 479200 92488 480000 92608
rect 0 91808 800 91928
rect 479200 91808 480000 91928
rect 0 91128 800 91248
rect 0 90448 800 90568
rect 479200 90448 480000 90568
rect 0 89768 800 89888
rect 479200 89768 480000 89888
rect 0 89088 800 89208
rect 479200 89088 480000 89208
rect 479200 88408 480000 88528
rect 0 87728 800 87848
rect 479200 87728 480000 87848
rect 0 87048 800 87168
rect 0 86368 800 86488
rect 479200 86368 480000 86488
rect 0 85688 800 85808
rect 479200 85688 480000 85808
rect 0 85008 800 85128
rect 479200 85008 480000 85128
rect 0 84328 800 84448
rect 479200 84328 480000 84448
rect 479200 83648 480000 83768
rect 0 82968 800 83088
rect 479200 82968 480000 83088
rect 0 82288 800 82408
rect 0 81608 800 81728
rect 479200 81608 480000 81728
rect 0 80928 800 81048
rect 479200 80928 480000 81048
rect 0 80248 800 80368
rect 479200 80248 480000 80368
rect 479200 79568 480000 79688
rect 0 78888 800 79008
rect 479200 78888 480000 79008
rect 0 78208 800 78328
rect 0 77528 800 77648
rect 479200 77528 480000 77648
rect 0 76848 800 76968
rect 479200 76848 480000 76968
rect 0 76168 800 76288
rect 479200 76168 480000 76288
rect 0 75488 800 75608
rect 479200 75488 480000 75608
rect 479200 74808 480000 74928
rect 0 74128 800 74248
rect 479200 74128 480000 74248
rect 0 73448 800 73568
rect 0 72768 800 72888
rect 479200 72768 480000 72888
rect 0 72088 800 72208
rect 479200 72088 480000 72208
rect 0 71408 800 71528
rect 479200 71408 480000 71528
rect 479200 70728 480000 70848
rect 0 70048 800 70168
rect 479200 70048 480000 70168
rect 0 69368 800 69488
rect 479200 69368 480000 69488
rect 0 68688 800 68808
rect 0 68008 800 68128
rect 479200 68008 480000 68128
rect 0 67328 800 67448
rect 479200 67328 480000 67448
rect 0 66648 800 66768
rect 479200 66648 480000 66768
rect 479200 65968 480000 66088
rect 0 65288 800 65408
rect 479200 65288 480000 65408
rect 0 64608 800 64728
rect 0 63928 800 64048
rect 479200 63928 480000 64048
rect 0 63248 800 63368
rect 479200 63248 480000 63368
rect 0 62568 800 62688
rect 479200 62568 480000 62688
rect 479200 61888 480000 62008
rect 0 61208 800 61328
rect 479200 61208 480000 61328
rect 0 60528 800 60648
rect 479200 60528 480000 60648
rect 0 59848 800 59968
rect 0 59168 800 59288
rect 479200 59168 480000 59288
rect 0 58488 800 58608
rect 479200 58488 480000 58608
rect 0 57808 800 57928
rect 479200 57808 480000 57928
rect 479200 57128 480000 57248
rect 0 56448 800 56568
rect 479200 56448 480000 56568
rect 0 55768 800 55888
rect 0 55088 800 55208
rect 479200 55088 480000 55208
rect 0 54408 800 54528
rect 479200 54408 480000 54528
rect 0 53728 800 53848
rect 479200 53728 480000 53848
rect 479200 53048 480000 53168
rect 0 52368 800 52488
rect 479200 52368 480000 52488
rect 0 51688 800 51808
rect 479200 51688 480000 51808
rect 0 51008 800 51128
rect 0 50328 800 50448
rect 479200 50328 480000 50448
rect 0 49648 800 49768
rect 479200 49648 480000 49768
rect 0 48968 800 49088
rect 479200 48968 480000 49088
rect 479200 48288 480000 48408
rect 0 47608 800 47728
rect 479200 47608 480000 47728
rect 0 46928 800 47048
rect 0 46248 800 46368
rect 479200 46248 480000 46368
rect 0 45568 800 45688
rect 479200 45568 480000 45688
rect 0 44888 800 45008
rect 479200 44888 480000 45008
rect 479200 44208 480000 44328
rect 0 43528 800 43648
rect 479200 43528 480000 43648
rect 0 42848 800 42968
rect 479200 42848 480000 42968
rect 0 42168 800 42288
rect 0 41488 800 41608
rect 479200 41488 480000 41608
rect 0 40808 800 40928
rect 479200 40808 480000 40928
rect 0 40128 800 40248
rect 479200 40128 480000 40248
rect 479200 39448 480000 39568
rect 0 38768 800 38888
rect 479200 38768 480000 38888
rect 0 38088 800 38208
rect 0 37408 800 37528
rect 479200 37408 480000 37528
rect 0 36728 800 36848
rect 479200 36728 480000 36848
rect 0 36048 800 36168
rect 479200 36048 480000 36168
rect 479200 35368 480000 35488
rect 0 34688 800 34808
rect 479200 34688 480000 34808
rect 0 34008 800 34128
rect 479200 34008 480000 34128
rect 0 33328 800 33448
rect 0 32648 800 32768
rect 479200 32648 480000 32768
rect 0 31968 800 32088
rect 479200 31968 480000 32088
rect 0 31288 800 31408
rect 479200 31288 480000 31408
rect 479200 30608 480000 30728
rect 0 29928 800 30048
rect 479200 29928 480000 30048
rect 0 29248 800 29368
rect 0 28568 800 28688
rect 479200 28568 480000 28688
rect 0 27888 800 28008
rect 479200 27888 480000 28008
rect 0 27208 800 27328
rect 479200 27208 480000 27328
rect 479200 26528 480000 26648
rect 0 25848 800 25968
rect 479200 25848 480000 25968
rect 0 25168 800 25288
rect 479200 25168 480000 25288
rect 0 24488 800 24608
rect 0 23808 800 23928
rect 479200 23808 480000 23928
rect 0 23128 800 23248
rect 479200 23128 480000 23248
rect 0 22448 800 22568
rect 479200 22448 480000 22568
rect 479200 21768 480000 21888
rect 0 21088 800 21208
rect 479200 21088 480000 21208
rect 0 20408 800 20528
rect 0 19728 800 19848
rect 479200 19728 480000 19848
rect 0 19048 800 19168
rect 479200 19048 480000 19168
rect 0 18368 800 18488
rect 479200 18368 480000 18488
rect 479200 17688 480000 17808
rect 0 17008 800 17128
rect 479200 17008 480000 17128
rect 0 16328 800 16448
rect 479200 16328 480000 16448
rect 0 15648 800 15768
rect 0 14968 800 15088
rect 479200 14968 480000 15088
rect 0 14288 800 14408
rect 479200 14288 480000 14408
rect 0 13608 800 13728
rect 479200 13608 480000 13728
rect 479200 12928 480000 13048
rect 0 12248 800 12368
rect 479200 12248 480000 12368
rect 0 11568 800 11688
rect 0 10888 800 11008
rect 479200 10888 480000 11008
rect 0 10208 800 10328
rect 479200 10208 480000 10328
rect 0 9528 800 9648
rect 479200 9528 480000 9648
rect 479200 8848 480000 8968
rect 0 8168 800 8288
rect 479200 8168 480000 8288
rect 0 7488 800 7608
rect 479200 7488 480000 7608
rect 0 6808 800 6928
rect 0 6128 800 6248
rect 479200 6128 480000 6248
rect 0 5448 800 5568
rect 479200 5448 480000 5568
rect 0 4768 800 4888
rect 479200 4768 480000 4888
rect 479200 4088 480000 4208
rect 0 3408 800 3528
rect 479200 3408 480000 3528
rect 0 2728 800 2848
rect 0 2048 800 2168
rect 479200 2048 480000 2168
rect 0 1368 800 1488
rect 479200 1368 480000 1488
rect 0 688 800 808
rect 479200 688 480000 808
rect 479200 8 480000 128
<< obsm3 >>
rect 800 119608 479120 119781
rect 800 119208 479200 119608
rect 880 118928 479120 119208
rect 800 118528 479200 118928
rect 880 118248 479120 118528
rect 800 117848 479200 118248
rect 880 117568 479200 117848
rect 800 117168 479200 117568
rect 880 116888 479120 117168
rect 800 116488 479200 116888
rect 880 116208 479120 116488
rect 800 115808 479200 116208
rect 880 115528 479120 115808
rect 800 115128 479200 115528
rect 800 114848 479120 115128
rect 800 114448 479200 114848
rect 880 114168 479120 114448
rect 800 113768 479200 114168
rect 880 113488 479200 113768
rect 800 113088 479200 113488
rect 880 112808 479120 113088
rect 800 112408 479200 112808
rect 880 112128 479120 112408
rect 800 111728 479200 112128
rect 880 111448 479120 111728
rect 800 111048 479200 111448
rect 800 110768 479120 111048
rect 800 110368 479200 110768
rect 880 110088 479120 110368
rect 800 109688 479200 110088
rect 880 109408 479120 109688
rect 800 109008 479200 109408
rect 880 108728 479200 109008
rect 800 108328 479200 108728
rect 880 108048 479120 108328
rect 800 107648 479200 108048
rect 880 107368 479120 107648
rect 800 106968 479200 107368
rect 880 106688 479120 106968
rect 800 106288 479200 106688
rect 800 106008 479120 106288
rect 800 105608 479200 106008
rect 880 105328 479120 105608
rect 800 104928 479200 105328
rect 880 104648 479200 104928
rect 800 104248 479200 104648
rect 880 103968 479120 104248
rect 800 103568 479200 103968
rect 880 103288 479120 103568
rect 800 102888 479200 103288
rect 880 102608 479120 102888
rect 800 102208 479200 102608
rect 800 101928 479120 102208
rect 800 101528 479200 101928
rect 880 101248 479120 101528
rect 800 100848 479200 101248
rect 880 100568 479120 100848
rect 800 100168 479200 100568
rect 880 99888 479200 100168
rect 800 99488 479200 99888
rect 880 99208 479120 99488
rect 800 98808 479200 99208
rect 880 98528 479120 98808
rect 800 98128 479200 98528
rect 880 97848 479120 98128
rect 800 97448 479200 97848
rect 800 97168 479120 97448
rect 800 96768 479200 97168
rect 880 96488 479120 96768
rect 800 96088 479200 96488
rect 880 95808 479200 96088
rect 800 95408 479200 95808
rect 880 95128 479120 95408
rect 800 94728 479200 95128
rect 880 94448 479120 94728
rect 800 94048 479200 94448
rect 880 93768 479120 94048
rect 800 93368 479200 93768
rect 880 93088 479120 93368
rect 800 92688 479200 93088
rect 800 92408 479120 92688
rect 800 92008 479200 92408
rect 880 91728 479120 92008
rect 800 91328 479200 91728
rect 880 91048 479200 91328
rect 800 90648 479200 91048
rect 880 90368 479120 90648
rect 800 89968 479200 90368
rect 880 89688 479120 89968
rect 800 89288 479200 89688
rect 880 89008 479120 89288
rect 800 88608 479200 89008
rect 800 88328 479120 88608
rect 800 87928 479200 88328
rect 880 87648 479120 87928
rect 800 87248 479200 87648
rect 880 86968 479200 87248
rect 800 86568 479200 86968
rect 880 86288 479120 86568
rect 800 85888 479200 86288
rect 880 85608 479120 85888
rect 800 85208 479200 85608
rect 880 84928 479120 85208
rect 800 84528 479200 84928
rect 880 84248 479120 84528
rect 800 83848 479200 84248
rect 800 83568 479120 83848
rect 800 83168 479200 83568
rect 880 82888 479120 83168
rect 800 82488 479200 82888
rect 880 82208 479200 82488
rect 800 81808 479200 82208
rect 880 81528 479120 81808
rect 800 81128 479200 81528
rect 880 80848 479120 81128
rect 800 80448 479200 80848
rect 880 80168 479120 80448
rect 800 79768 479200 80168
rect 800 79488 479120 79768
rect 800 79088 479200 79488
rect 880 78808 479120 79088
rect 800 78408 479200 78808
rect 880 78128 479200 78408
rect 800 77728 479200 78128
rect 880 77448 479120 77728
rect 800 77048 479200 77448
rect 880 76768 479120 77048
rect 800 76368 479200 76768
rect 880 76088 479120 76368
rect 800 75688 479200 76088
rect 880 75408 479120 75688
rect 800 75008 479200 75408
rect 800 74728 479120 75008
rect 800 74328 479200 74728
rect 880 74048 479120 74328
rect 800 73648 479200 74048
rect 880 73368 479200 73648
rect 800 72968 479200 73368
rect 880 72688 479120 72968
rect 800 72288 479200 72688
rect 880 72008 479120 72288
rect 800 71608 479200 72008
rect 880 71328 479120 71608
rect 800 70928 479200 71328
rect 800 70648 479120 70928
rect 800 70248 479200 70648
rect 880 69968 479120 70248
rect 800 69568 479200 69968
rect 880 69288 479120 69568
rect 800 68888 479200 69288
rect 880 68608 479200 68888
rect 800 68208 479200 68608
rect 880 67928 479120 68208
rect 800 67528 479200 67928
rect 880 67248 479120 67528
rect 800 66848 479200 67248
rect 880 66568 479120 66848
rect 800 66168 479200 66568
rect 800 65888 479120 66168
rect 800 65488 479200 65888
rect 880 65208 479120 65488
rect 800 64808 479200 65208
rect 880 64528 479200 64808
rect 800 64128 479200 64528
rect 880 63848 479120 64128
rect 800 63448 479200 63848
rect 880 63168 479120 63448
rect 800 62768 479200 63168
rect 880 62488 479120 62768
rect 800 62088 479200 62488
rect 800 61808 479120 62088
rect 800 61408 479200 61808
rect 880 61128 479120 61408
rect 800 60728 479200 61128
rect 880 60448 479120 60728
rect 800 60048 479200 60448
rect 880 59768 479200 60048
rect 800 59368 479200 59768
rect 880 59088 479120 59368
rect 800 58688 479200 59088
rect 880 58408 479120 58688
rect 800 58008 479200 58408
rect 880 57728 479120 58008
rect 800 57328 479200 57728
rect 800 57048 479120 57328
rect 800 56648 479200 57048
rect 880 56368 479120 56648
rect 800 55968 479200 56368
rect 880 55688 479200 55968
rect 800 55288 479200 55688
rect 880 55008 479120 55288
rect 800 54608 479200 55008
rect 880 54328 479120 54608
rect 800 53928 479200 54328
rect 880 53648 479120 53928
rect 800 53248 479200 53648
rect 800 52968 479120 53248
rect 800 52568 479200 52968
rect 880 52288 479120 52568
rect 800 51888 479200 52288
rect 880 51608 479120 51888
rect 800 51208 479200 51608
rect 880 50928 479200 51208
rect 800 50528 479200 50928
rect 880 50248 479120 50528
rect 800 49848 479200 50248
rect 880 49568 479120 49848
rect 800 49168 479200 49568
rect 880 48888 479120 49168
rect 800 48488 479200 48888
rect 800 48208 479120 48488
rect 800 47808 479200 48208
rect 880 47528 479120 47808
rect 800 47128 479200 47528
rect 880 46848 479200 47128
rect 800 46448 479200 46848
rect 880 46168 479120 46448
rect 800 45768 479200 46168
rect 880 45488 479120 45768
rect 800 45088 479200 45488
rect 880 44808 479120 45088
rect 800 44408 479200 44808
rect 800 44128 479120 44408
rect 800 43728 479200 44128
rect 880 43448 479120 43728
rect 800 43048 479200 43448
rect 880 42768 479120 43048
rect 800 42368 479200 42768
rect 880 42088 479200 42368
rect 800 41688 479200 42088
rect 880 41408 479120 41688
rect 800 41008 479200 41408
rect 880 40728 479120 41008
rect 800 40328 479200 40728
rect 880 40048 479120 40328
rect 800 39648 479200 40048
rect 800 39368 479120 39648
rect 800 38968 479200 39368
rect 880 38688 479120 38968
rect 800 38288 479200 38688
rect 880 38008 479200 38288
rect 800 37608 479200 38008
rect 880 37328 479120 37608
rect 800 36928 479200 37328
rect 880 36648 479120 36928
rect 800 36248 479200 36648
rect 880 35968 479120 36248
rect 800 35568 479200 35968
rect 800 35288 479120 35568
rect 800 34888 479200 35288
rect 880 34608 479120 34888
rect 800 34208 479200 34608
rect 880 33928 479120 34208
rect 800 33528 479200 33928
rect 880 33248 479200 33528
rect 800 32848 479200 33248
rect 880 32568 479120 32848
rect 800 32168 479200 32568
rect 880 31888 479120 32168
rect 800 31488 479200 31888
rect 880 31208 479120 31488
rect 800 30808 479200 31208
rect 800 30528 479120 30808
rect 800 30128 479200 30528
rect 880 29848 479120 30128
rect 800 29448 479200 29848
rect 880 29168 479200 29448
rect 800 28768 479200 29168
rect 880 28488 479120 28768
rect 800 28088 479200 28488
rect 880 27808 479120 28088
rect 800 27408 479200 27808
rect 880 27128 479120 27408
rect 800 26728 479200 27128
rect 800 26448 479120 26728
rect 800 26048 479200 26448
rect 880 25768 479120 26048
rect 800 25368 479200 25768
rect 880 25088 479120 25368
rect 800 24688 479200 25088
rect 880 24408 479200 24688
rect 800 24008 479200 24408
rect 880 23728 479120 24008
rect 800 23328 479200 23728
rect 880 23048 479120 23328
rect 800 22648 479200 23048
rect 880 22368 479120 22648
rect 800 21968 479200 22368
rect 800 21688 479120 21968
rect 800 21288 479200 21688
rect 880 21008 479120 21288
rect 800 20608 479200 21008
rect 880 20328 479200 20608
rect 800 19928 479200 20328
rect 880 19648 479120 19928
rect 800 19248 479200 19648
rect 880 18968 479120 19248
rect 800 18568 479200 18968
rect 880 18288 479120 18568
rect 800 17888 479200 18288
rect 800 17608 479120 17888
rect 800 17208 479200 17608
rect 880 16928 479120 17208
rect 800 16528 479200 16928
rect 880 16248 479120 16528
rect 800 15848 479200 16248
rect 880 15568 479200 15848
rect 800 15168 479200 15568
rect 880 14888 479120 15168
rect 800 14488 479200 14888
rect 880 14208 479120 14488
rect 800 13808 479200 14208
rect 880 13528 479120 13808
rect 800 13128 479200 13528
rect 800 12848 479120 13128
rect 800 12448 479200 12848
rect 880 12168 479120 12448
rect 800 11768 479200 12168
rect 880 11488 479200 11768
rect 800 11088 479200 11488
rect 880 10808 479120 11088
rect 800 10408 479200 10808
rect 880 10128 479120 10408
rect 800 9728 479200 10128
rect 880 9448 479120 9728
rect 800 9048 479200 9448
rect 800 8768 479120 9048
rect 800 8368 479200 8768
rect 880 8088 479120 8368
rect 800 7688 479200 8088
rect 880 7408 479120 7688
rect 800 7008 479200 7408
rect 880 6728 479200 7008
rect 800 6328 479200 6728
rect 880 6048 479120 6328
rect 800 5648 479200 6048
rect 880 5368 479120 5648
rect 800 4968 479200 5368
rect 880 4688 479120 4968
rect 800 4288 479200 4688
rect 800 4008 479120 4288
rect 800 3608 479200 4008
rect 880 3328 479120 3608
rect 800 2928 479200 3328
rect 880 2648 479200 2928
rect 800 2248 479200 2648
rect 880 1968 479120 2248
rect 800 1568 479200 1968
rect 880 1288 479120 1568
rect 800 888 479200 1288
rect 880 608 479120 888
rect 800 208 479200 608
rect 800 35 479120 208
<< metal4 >>
rect 4208 2128 4528 117552
rect 19568 2128 19888 117552
rect 34928 2128 35248 117552
rect 50288 2128 50608 117552
rect 65648 2128 65968 117552
rect 81008 2128 81328 117552
rect 96368 2128 96688 117552
rect 111728 2128 112048 117552
rect 127088 2128 127408 117552
rect 142448 2128 142768 117552
rect 157808 2128 158128 117552
rect 173168 2128 173488 117552
rect 188528 2128 188848 117552
rect 203888 2128 204208 117552
rect 219248 2128 219568 117552
rect 234608 2128 234928 117552
rect 249968 2128 250288 117552
rect 265328 2128 265648 117552
rect 280688 2128 281008 117552
rect 296048 2128 296368 117552
rect 311408 2128 311728 117552
rect 326768 2128 327088 117552
rect 342128 2128 342448 117552
rect 357488 2128 357808 117552
rect 372848 2128 373168 117552
rect 388208 2128 388528 117552
rect 403568 2128 403888 117552
rect 418928 2128 419248 117552
rect 434288 2128 434608 117552
rect 449648 2128 449968 117552
rect 465008 2128 465328 117552
<< obsm4 >>
rect 169891 2048 173088 117333
rect 173568 2048 188448 117333
rect 188928 2048 203808 117333
rect 204288 2048 219168 117333
rect 219648 2048 234528 117333
rect 235008 2048 249888 117333
rect 250368 2048 265248 117333
rect 265728 2048 280608 117333
rect 281088 2048 295968 117333
rect 296448 2048 311328 117333
rect 311808 2048 326541 117333
rect 169891 1667 326541 2048
<< labels >>
rlabel metal2 s 390926 0 390982 800 6 clk
port 1 nsew signal input
rlabel metal2 s 226062 0 226118 800 6 m00_ar_addr[0]
port 2 nsew signal output
rlabel metal2 s 161662 119200 161718 120000 6 m00_ar_addr[10]
port 3 nsew signal output
rlabel metal2 s 128818 0 128874 800 6 m00_ar_addr[11]
port 4 nsew signal output
rlabel metal2 s 81806 119200 81862 120000 6 m00_ar_addr[12]
port 5 nsew signal output
rlabel metal2 s 343270 119200 343326 120000 6 m00_ar_addr[13]
port 6 nsew signal output
rlabel metal3 s 0 15648 800 15768 6 m00_ar_addr[14]
port 7 nsew signal output
rlabel metal2 s 170034 119200 170090 120000 6 m00_ar_addr[15]
port 8 nsew signal output
rlabel metal2 s 242162 119200 242218 120000 6 m00_ar_addr[16]
port 9 nsew signal output
rlabel metal3 s 479200 4768 480000 4888 6 m00_ar_addr[17]
port 10 nsew signal output
rlabel metal2 s 442446 0 442502 800 6 m00_ar_addr[18]
port 11 nsew signal output
rlabel metal2 s 451462 0 451518 800 6 m00_ar_addr[19]
port 12 nsew signal output
rlabel metal3 s 479200 99288 480000 99408 6 m00_ar_addr[1]
port 13 nsew signal output
rlabel metal2 s 206098 119200 206154 120000 6 m00_ar_addr[20]
port 14 nsew signal output
rlabel metal2 s 454038 0 454094 800 6 m00_ar_addr[21]
port 15 nsew signal output
rlabel metal2 s 262770 119200 262826 120000 6 m00_ar_addr[22]
port 16 nsew signal output
rlabel metal2 s 59910 119200 59966 120000 6 m00_ar_addr[23]
port 17 nsew signal output
rlabel metal2 s 356150 0 356206 800 6 m00_ar_addr[24]
port 18 nsew signal output
rlabel metal2 s 468206 0 468262 800 6 m00_ar_addr[25]
port 19 nsew signal output
rlabel metal2 s 69570 0 69626 800 6 m00_ar_addr[26]
port 20 nsew signal output
rlabel metal2 s 239586 0 239642 800 6 m00_ar_addr[27]
port 21 nsew signal output
rlabel metal2 s 340694 119200 340750 120000 6 m00_ar_addr[28]
port 22 nsew signal output
rlabel metal2 s 172610 119200 172666 120000 6 m00_ar_addr[29]
port 23 nsew signal output
rlabel metal2 s 354862 119200 354918 120000 6 m00_ar_addr[2]
port 24 nsew signal output
rlabel metal2 s 16762 119200 16818 120000 6 m00_ar_addr[30]
port 25 nsew signal output
rlabel metal2 s 1306 0 1362 800 6 m00_ar_addr[31]
port 26 nsew signal output
rlabel metal3 s 479200 25848 480000 25968 6 m00_ar_addr[3]
port 27 nsew signal output
rlabel metal3 s 0 109488 800 109608 6 m00_ar_addr[4]
port 28 nsew signal output
rlabel metal2 s 367098 0 367154 800 6 m00_ar_addr[5]
port 29 nsew signal output
rlabel metal2 s 110786 119200 110842 120000 6 m00_ar_addr[6]
port 30 nsew signal output
rlabel metal2 s 235722 119200 235778 120000 6 m00_ar_addr[7]
port 31 nsew signal output
rlabel metal2 s 199014 0 199070 800 6 m00_ar_addr[8]
port 32 nsew signal output
rlabel metal2 s 304630 0 304686 800 6 m00_ar_addr[9]
port 33 nsew signal output
rlabel metal2 s 106922 119200 106978 120000 6 m00_ar_burst[0]
port 34 nsew signal output
rlabel metal2 s 153934 0 153990 800 6 m00_ar_burst[1]
port 35 nsew signal output
rlabel metal2 s 115938 119200 115994 120000 6 m00_ar_cache[0]
port 36 nsew signal output
rlabel metal2 s 358082 119200 358138 120000 6 m00_ar_cache[1]
port 37 nsew signal output
rlabel metal2 s 132682 0 132738 800 6 m00_ar_cache[2]
port 38 nsew signal output
rlabel metal2 s 331678 119200 331734 120000 6 m00_ar_cache[3]
port 39 nsew signal output
rlabel metal3 s 0 23808 800 23928 6 m00_ar_id[0]
port 40 nsew signal output
rlabel metal2 s 278870 0 278926 800 6 m00_ar_id[10]
port 41 nsew signal output
rlabel metal2 s 355506 0 355562 800 6 m00_ar_id[11]
port 42 nsew signal output
rlabel metal3 s 479200 68008 480000 68128 6 m00_ar_id[1]
port 43 nsew signal output
rlabel metal3 s 479200 25168 480000 25288 6 m00_ar_id[2]
port 44 nsew signal output
rlabel metal2 s 101770 0 101826 800 6 m00_ar_id[3]
port 45 nsew signal output
rlabel metal3 s 479200 53048 480000 53168 6 m00_ar_id[4]
port 46 nsew signal output
rlabel metal2 s 76654 119200 76710 120000 6 m00_ar_id[5]
port 47 nsew signal output
rlabel metal3 s 479200 110168 480000 110288 6 m00_ar_id[6]
port 48 nsew signal output
rlabel metal2 s 364522 0 364578 800 6 m00_ar_id[7]
port 49 nsew signal output
rlabel metal2 s 265990 119200 266046 120000 6 m00_ar_id[8]
port 50 nsew signal output
rlabel metal3 s 479200 98608 480000 98728 6 m00_ar_id[9]
port 51 nsew signal output
rlabel metal2 s 180338 119200 180394 120000 6 m00_ar_len[0]
port 52 nsew signal output
rlabel metal2 s 222198 119200 222254 120000 6 m00_ar_len[1]
port 53 nsew signal output
rlabel metal2 s 263414 119200 263470 120000 6 m00_ar_len[2]
port 54 nsew signal output
rlabel metal2 s 191930 119200 191986 120000 6 m00_ar_len[3]
port 55 nsew signal output
rlabel metal2 s 164238 119200 164294 120000 6 m00_ar_len[4]
port 56 nsew signal output
rlabel metal3 s 0 72768 800 72888 6 m00_ar_len[5]
port 57 nsew signal output
rlabel metal2 s 351642 119200 351698 120000 6 m00_ar_len[6]
port 58 nsew signal output
rlabel metal2 s 408958 0 409014 800 6 m00_ar_len[7]
port 59 nsew signal output
rlabel metal2 s 280158 119200 280214 120000 6 m00_ar_lock
port 60 nsew signal output
rlabel metal2 s 442446 119200 442502 120000 6 m00_ar_prot[0]
port 61 nsew signal output
rlabel metal2 s 418618 0 418674 800 6 m00_ar_prot[1]
port 62 nsew signal output
rlabel metal2 s 169390 119200 169446 120000 6 m00_ar_prot[2]
port 63 nsew signal output
rlabel metal3 s 479200 12248 480000 12368 6 m00_ar_qos[0]
port 64 nsew signal output
rlabel metal2 s 258262 119200 258318 120000 6 m00_ar_qos[1]
port 65 nsew signal output
rlabel metal3 s 479200 16328 480000 16448 6 m00_ar_qos[2]
port 66 nsew signal output
rlabel metal2 s 225418 119200 225474 120000 6 m00_ar_qos[3]
port 67 nsew signal output
rlabel metal2 s 2594 0 2650 800 6 m00_ar_ready
port 68 nsew signal input
rlabel metal3 s 0 46928 800 47048 6 m00_ar_region[0]
port 69 nsew signal output
rlabel metal2 s 110786 0 110842 800 6 m00_ar_region[1]
port 70 nsew signal output
rlabel metal2 s 320730 119200 320786 120000 6 m00_ar_region[2]
port 71 nsew signal output
rlabel metal2 s 7102 119200 7158 120000 6 m00_ar_region[3]
port 72 nsew signal output
rlabel metal2 s 1306 119200 1362 120000 6 m00_ar_size[0]
port 73 nsew signal output
rlabel metal3 s 479200 76168 480000 76288 6 m00_ar_size[1]
port 74 nsew signal output
rlabel metal2 s 307206 0 307262 800 6 m00_ar_size[2]
port 75 nsew signal output
rlabel metal2 s 124310 0 124366 800 6 m00_ar_user[-1]
port 76 nsew signal output
rlabel metal2 s 170678 119200 170734 120000 6 m00_ar_user[0]
port 77 nsew signal output
rlabel metal2 s 365166 119200 365222 120000 6 m00_ar_valid
port 78 nsew signal output
rlabel metal2 s 186778 0 186834 800 6 m00_aw_addr[0]
port 79 nsew signal output
rlabel metal2 s 386418 119200 386474 120000 6 m00_aw_addr[10]
port 80 nsew signal output
rlabel metal2 s 101770 119200 101826 120000 6 m00_aw_addr[11]
port 81 nsew signal output
rlabel metal2 s 156510 0 156566 800 6 m00_aw_addr[12]
port 82 nsew signal output
rlabel metal3 s 479200 100648 480000 100768 6 m00_aw_addr[13]
port 83 nsew signal output
rlabel metal3 s 479200 8168 480000 8288 6 m00_aw_addr[14]
port 84 nsew signal output
rlabel metal2 s 191286 0 191342 800 6 m00_aw_addr[15]
port 85 nsew signal output
rlabel metal3 s 479200 44888 480000 45008 6 m00_aw_addr[16]
port 86 nsew signal output
rlabel metal2 s 432786 119200 432842 120000 6 m00_aw_addr[17]
port 87 nsew signal output
rlabel metal3 s 479200 65288 480000 65408 6 m00_aw_addr[18]
port 88 nsew signal output
rlabel metal2 s 265990 0 266046 800 6 m00_aw_addr[19]
port 89 nsew signal output
rlabel metal3 s 479200 82968 480000 83088 6 m00_aw_addr[1]
port 90 nsew signal output
rlabel metal2 s 135902 0 135958 800 6 m00_aw_addr[20]
port 91 nsew signal output
rlabel metal3 s 0 97928 800 98048 6 m00_aw_addr[21]
port 92 nsew signal output
rlabel metal2 s 249890 119200 249946 120000 6 m00_aw_addr[22]
port 93 nsew signal output
rlabel metal2 s 296258 0 296314 800 6 m00_aw_addr[23]
port 94 nsew signal output
rlabel metal2 s 204166 119200 204222 120000 6 m00_aw_addr[24]
port 95 nsew signal output
rlabel metal2 s 99194 119200 99250 120000 6 m00_aw_addr[25]
port 96 nsew signal output
rlabel metal2 s 294970 0 295026 800 6 m00_aw_addr[26]
port 97 nsew signal output
rlabel metal2 s 367742 0 367798 800 6 m00_aw_addr[27]
port 98 nsew signal output
rlabel metal3 s 479200 77528 480000 77648 6 m00_aw_addr[28]
port 99 nsew signal output
rlabel metal2 s 19338 119200 19394 120000 6 m00_aw_addr[29]
port 100 nsew signal output
rlabel metal2 s 413466 0 413522 800 6 m00_aw_addr[2]
port 101 nsew signal output
rlabel metal2 s 421194 119200 421250 120000 6 m00_aw_addr[30]
port 102 nsew signal output
rlabel metal2 s 106922 0 106978 800 6 m00_aw_addr[31]
port 103 nsew signal output
rlabel metal2 s 399942 119200 399998 120000 6 m00_aw_addr[3]
port 104 nsew signal output
rlabel metal2 s 403806 0 403862 800 6 m00_aw_addr[4]
port 105 nsew signal output
rlabel metal2 s 48962 119200 49018 120000 6 m00_aw_addr[5]
port 106 nsew signal output
rlabel metal2 s 322018 0 322074 800 6 m00_aw_addr[6]
port 107 nsew signal output
rlabel metal2 s 277582 0 277638 800 6 m00_aw_addr[7]
port 108 nsew signal output
rlabel metal2 s 199658 119200 199714 120000 6 m00_aw_addr[8]
port 109 nsew signal output
rlabel metal3 s 0 90448 800 90568 6 m00_aw_addr[9]
port 110 nsew signal output
rlabel metal2 s 283378 0 283434 800 6 m00_aw_burst[0]
port 111 nsew signal output
rlabel metal2 s 65706 0 65762 800 6 m00_aw_burst[1]
port 112 nsew signal output
rlabel metal3 s 0 14968 800 15088 6 m00_aw_cache[0]
port 113 nsew signal output
rlabel metal2 s 324594 119200 324650 120000 6 m00_aw_cache[1]
port 114 nsew signal output
rlabel metal3 s 479200 74128 480000 74248 6 m00_aw_cache[2]
port 115 nsew signal output
rlabel metal3 s 0 40128 800 40248 6 m00_aw_cache[3]
port 116 nsew signal output
rlabel metal2 s 113362 119200 113418 120000 6 m00_aw_id[0]
port 117 nsew signal output
rlabel metal2 s 320086 0 320142 800 6 m00_aw_id[10]
port 118 nsew signal output
rlabel metal3 s 0 61208 800 61328 6 m00_aw_id[11]
port 119 nsew signal output
rlabel metal2 s 187422 119200 187478 120000 6 m00_aw_id[1]
port 120 nsew signal output
rlabel metal2 s 209962 119200 210018 120000 6 m00_aw_id[2]
port 121 nsew signal output
rlabel metal2 s 36082 119200 36138 120000 6 m00_aw_id[3]
port 122 nsew signal output
rlabel metal3 s 479200 116968 480000 117088 6 m00_aw_id[4]
port 123 nsew signal output
rlabel metal2 s 92754 0 92810 800 6 m00_aw_id[5]
port 124 nsew signal output
rlabel metal2 s 312358 0 312414 800 6 m00_aw_id[6]
port 125 nsew signal output
rlabel metal2 s 370318 0 370374 800 6 m00_aw_id[7]
port 126 nsew signal output
rlabel metal2 s 18694 119200 18750 120000 6 m00_aw_id[8]
port 127 nsew signal output
rlabel metal2 s 106278 119200 106334 120000 6 m00_aw_id[9]
port 128 nsew signal output
rlabel metal2 s 274362 0 274418 800 6 m00_aw_len[0]
port 129 nsew signal output
rlabel metal2 s 446310 119200 446366 120000 6 m00_aw_len[1]
port 130 nsew signal output
rlabel metal2 s 102414 0 102470 800 6 m00_aw_len[2]
port 131 nsew signal output
rlabel metal3 s 479200 71408 480000 71528 6 m00_aw_len[3]
port 132 nsew signal output
rlabel metal2 s 115294 119200 115350 120000 6 m00_aw_len[4]
port 133 nsew signal output
rlabel metal2 s 326526 0 326582 800 6 m00_aw_len[5]
port 134 nsew signal output
rlabel metal2 s 193218 119200 193274 120000 6 m00_aw_len[6]
port 135 nsew signal output
rlabel metal2 s 185490 119200 185546 120000 6 m00_aw_len[7]
port 136 nsew signal output
rlabel metal2 s 166170 119200 166226 120000 6 m00_aw_lock
port 137 nsew signal output
rlabel metal2 s 197726 0 197782 800 6 m00_aw_prot[0]
port 138 nsew signal output
rlabel metal2 s 283378 119200 283434 120000 6 m00_aw_prot[1]
port 139 nsew signal output
rlabel metal2 s 49606 0 49662 800 6 m00_aw_prot[2]
port 140 nsew signal output
rlabel metal2 s 9034 119200 9090 120000 6 m00_aw_qos[0]
port 141 nsew signal output
rlabel metal2 s 257618 119200 257674 120000 6 m00_aw_qos[1]
port 142 nsew signal output
rlabel metal3 s 0 85008 800 85128 6 m00_aw_qos[2]
port 143 nsew signal output
rlabel metal2 s 26422 119200 26478 120000 6 m00_aw_qos[3]
port 144 nsew signal output
rlabel metal2 s 375470 119200 375526 120000 6 m00_aw_ready
port 145 nsew signal input
rlabel metal2 s 262770 0 262826 800 6 m00_aw_region[0]
port 146 nsew signal output
rlabel metal2 s 27710 0 27766 800 6 m00_aw_region[1]
port 147 nsew signal output
rlabel metal2 s 259550 0 259606 800 6 m00_aw_region[2]
port 148 nsew signal output
rlabel metal3 s 0 93168 800 93288 6 m00_aw_region[3]
port 149 nsew signal output
rlabel metal2 s 247958 119200 248014 120000 6 m00_aw_size[0]
port 150 nsew signal output
rlabel metal2 s 36082 0 36138 800 6 m00_aw_size[1]
port 151 nsew signal output
rlabel metal3 s 479200 103368 480000 103488 6 m00_aw_size[2]
port 152 nsew signal output
rlabel metal2 s 195794 0 195850 800 6 m00_aw_user[-1]
port 153 nsew signal output
rlabel metal2 s 371606 119200 371662 120000 6 m00_aw_user[0]
port 154 nsew signal output
rlabel metal2 s 406382 0 406438 800 6 m00_aw_valid
port 155 nsew signal output
rlabel metal2 s 126886 0 126942 800 6 m00_b_id[0]
port 156 nsew signal input
rlabel metal2 s 15474 0 15530 800 6 m00_b_id[10]
port 157 nsew signal input
rlabel metal2 s 345202 119200 345258 120000 6 m00_b_id[11]
port 158 nsew signal input
rlabel metal2 s 362590 0 362646 800 6 m00_b_id[1]
port 159 nsew signal input
rlabel metal2 s 417974 0 418030 800 6 m00_b_id[2]
port 160 nsew signal input
rlabel metal3 s 479200 93168 480000 93288 6 m00_b_id[3]
port 161 nsew signal input
rlabel metal2 s 72790 0 72846 800 6 m00_b_id[4]
port 162 nsew signal input
rlabel metal2 s 354218 0 354274 800 6 m00_b_id[5]
port 163 nsew signal input
rlabel metal2 s 155866 0 155922 800 6 m00_b_id[6]
port 164 nsew signal input
rlabel metal2 s 293682 119200 293738 120000 6 m00_b_id[7]
port 165 nsew signal input
rlabel metal2 s 376114 0 376170 800 6 m00_b_id[8]
port 166 nsew signal input
rlabel metal2 s 18694 0 18750 800 6 m00_b_id[9]
port 167 nsew signal input
rlabel metal2 s 64418 0 64474 800 6 m00_b_ready
port 168 nsew signal output
rlabel metal2 s 402518 0 402574 800 6 m00_b_resp[0]
port 169 nsew signal input
rlabel metal2 s 276294 0 276350 800 6 m00_b_resp[1]
port 170 nsew signal input
rlabel metal2 s 323950 0 324006 800 6 m00_b_user[-1]
port 171 nsew signal input
rlabel metal3 s 479200 89088 480000 89208 6 m00_b_user[0]
port 172 nsew signal input
rlabel metal2 s 79874 0 79930 800 6 m00_b_valid
port 173 nsew signal input
rlabel metal2 s 278226 119200 278282 120000 6 m00_r_data[0]
port 174 nsew signal input
rlabel metal2 s 250534 0 250590 800 6 m00_r_data[10]
port 175 nsew signal input
rlabel metal2 s 228638 119200 228694 120000 6 m00_r_data[11]
port 176 nsew signal input
rlabel metal2 s 447598 0 447654 800 6 m00_r_data[12]
port 177 nsew signal input
rlabel metal3 s 0 106768 800 106888 6 m00_r_data[13]
port 178 nsew signal input
rlabel metal2 s 267922 0 267978 800 6 m00_r_data[14]
port 179 nsew signal input
rlabel metal2 s 477222 119200 477278 120000 6 m00_r_data[15]
port 180 nsew signal input
rlabel metal2 s 65706 119200 65762 120000 6 m00_r_data[16]
port 181 nsew signal input
rlabel metal2 s 97906 0 97962 800 6 m00_r_data[17]
port 182 nsew signal input
rlabel metal2 s 258262 0 258318 800 6 m00_r_data[18]
port 183 nsew signal input
rlabel metal2 s 294326 0 294382 800 6 m00_r_data[19]
port 184 nsew signal input
rlabel metal3 s 0 14288 800 14408 6 m00_r_data[1]
port 185 nsew signal input
rlabel metal2 s 10966 119200 11022 120000 6 m00_r_data[20]
port 186 nsew signal input
rlabel metal3 s 479200 87728 480000 87848 6 m00_r_data[21]
port 187 nsew signal input
rlabel metal2 s 119158 0 119214 800 6 m00_r_data[22]
port 188 nsew signal input
rlabel metal2 s 155866 119200 155922 120000 6 m00_r_data[23]
port 189 nsew signal input
rlabel metal2 s 18 119200 74 120000 6 m00_r_data[24]
port 190 nsew signal input
rlabel metal3 s 479200 10208 480000 10328 6 m00_r_data[25]
port 191 nsew signal input
rlabel metal2 s 77298 0 77354 800 6 m00_r_data[26]
port 192 nsew signal input
rlabel metal2 s 216402 119200 216458 120000 6 m00_r_data[27]
port 193 nsew signal input
rlabel metal3 s 479200 8848 480000 8968 6 m00_r_data[28]
port 194 nsew signal input
rlabel metal2 s 137190 0 137246 800 6 m00_r_data[29]
port 195 nsew signal input
rlabel metal2 s 88890 119200 88946 120000 6 m00_r_data[2]
port 196 nsew signal input
rlabel metal2 s 271142 119200 271198 120000 6 m00_r_data[30]
port 197 nsew signal input
rlabel metal2 s 105634 119200 105690 120000 6 m00_r_data[31]
port 198 nsew signal input
rlabel metal2 s 35438 119200 35494 120000 6 m00_r_data[3]
port 199 nsew signal input
rlabel metal2 s 42522 119200 42578 120000 6 m00_r_data[4]
port 200 nsew signal input
rlabel metal2 s 130106 119200 130162 120000 6 m00_r_data[5]
port 201 nsew signal input
rlabel metal2 s 123666 119200 123722 120000 6 m00_r_data[6]
port 202 nsew signal input
rlabel metal2 s 336186 0 336242 800 6 m00_r_data[7]
port 203 nsew signal input
rlabel metal2 s 374826 119200 374882 120000 6 m00_r_data[8]
port 204 nsew signal input
rlabel metal2 s 134614 0 134670 800 6 m00_r_data[9]
port 205 nsew signal input
rlabel metal2 s 186778 119200 186834 120000 6 m00_r_id[0]
port 206 nsew signal input
rlabel metal3 s 479200 102008 480000 102128 6 m00_r_id[10]
port 207 nsew signal input
rlabel metal2 s 90178 0 90234 800 6 m00_r_id[11]
port 208 nsew signal input
rlabel metal2 s 97262 119200 97318 120000 6 m00_r_id[1]
port 209 nsew signal input
rlabel metal2 s 370962 119200 371018 120000 6 m00_r_id[2]
port 210 nsew signal input
rlabel metal2 s 177762 0 177818 800 6 m00_r_id[3]
port 211 nsew signal input
rlabel metal2 s 344558 119200 344614 120000 6 m00_r_id[4]
port 212 nsew signal input
rlabel metal2 s 23846 119200 23902 120000 6 m00_r_id[5]
port 213 nsew signal input
rlabel metal2 s 328458 119200 328514 120000 6 m00_r_id[6]
port 214 nsew signal input
rlabel metal2 s 358726 119200 358782 120000 6 m00_r_id[7]
port 215 nsew signal input
rlabel metal2 s 1950 0 2006 800 6 m00_r_id[8]
port 216 nsew signal input
rlabel metal2 s 85670 0 85726 800 6 m00_r_id[9]
port 217 nsew signal input
rlabel metal2 s 252466 0 252522 800 6 m00_r_last
port 218 nsew signal input
rlabel metal2 s 12898 0 12954 800 6 m00_r_ready
port 219 nsew signal output
rlabel metal2 s 305274 0 305330 800 6 m00_r_resp[0]
port 220 nsew signal input
rlabel metal2 s 399942 0 399998 800 6 m00_r_resp[1]
port 221 nsew signal input
rlabel metal2 s 340694 0 340750 800 6 m00_r_user[-1]
port 222 nsew signal input
rlabel metal3 s 0 12248 800 12368 6 m00_r_user[0]
port 223 nsew signal input
rlabel metal2 s 479154 0 479210 800 6 m00_r_valid
port 224 nsew signal input
rlabel metal2 s 48318 0 48374 800 6 m00_w_data[0]
port 225 nsew signal output
rlabel metal2 s 392214 119200 392270 120000 6 m00_w_data[10]
port 226 nsew signal output
rlabel metal2 s 468206 119200 468262 120000 6 m00_w_data[11]
port 227 nsew signal output
rlabel metal2 s 245382 0 245438 800 6 m00_w_data[12]
port 228 nsew signal output
rlabel metal2 s 40590 119200 40646 120000 6 m00_w_data[13]
port 229 nsew signal output
rlabel metal2 s 85026 0 85082 800 6 m00_w_data[14]
port 230 nsew signal output
rlabel metal3 s 0 108808 800 108928 6 m00_w_data[15]
port 231 nsew signal output
rlabel metal2 s 189354 0 189410 800 6 m00_w_data[16]
port 232 nsew signal output
rlabel metal2 s 320086 119200 320142 120000 6 m00_w_data[17]
port 233 nsew signal output
rlabel metal2 s 412178 0 412234 800 6 m00_w_data[18]
port 234 nsew signal output
rlabel metal2 s 361302 119200 361358 120000 6 m00_w_data[19]
port 235 nsew signal output
rlabel metal3 s 0 22448 800 22568 6 m00_w_data[1]
port 236 nsew signal output
rlabel metal2 s 42522 0 42578 800 6 m00_w_data[20]
port 237 nsew signal output
rlabel metal2 s 435362 0 435418 800 6 m00_w_data[21]
port 238 nsew signal output
rlabel metal2 s 73434 119200 73490 120000 6 m00_w_data[22]
port 239 nsew signal output
rlabel metal2 s 59910 0 59966 800 6 m00_w_data[23]
port 240 nsew signal output
rlabel metal3 s 479200 8 480000 128 6 m00_w_data[24]
port 241 nsew signal output
rlabel metal3 s 479200 75488 480000 75608 6 m00_w_data[25]
port 242 nsew signal output
rlabel metal2 s 401874 119200 401930 120000 6 m00_w_data[26]
port 243 nsew signal output
rlabel metal3 s 479200 119008 480000 119128 6 m00_w_data[27]
port 244 nsew signal output
rlabel metal2 s 335542 119200 335598 120000 6 m00_w_data[28]
port 245 nsew signal output
rlabel metal2 s 112718 0 112774 800 6 m00_w_data[29]
port 246 nsew signal output
rlabel metal3 s 0 118328 800 118448 6 m00_w_data[2]
port 247 nsew signal output
rlabel metal2 s 225418 0 225474 800 6 m00_w_data[30]
port 248 nsew signal output
rlabel metal3 s 0 31288 800 31408 6 m00_w_data[31]
port 249 nsew signal output
rlabel metal2 s 395434 119200 395490 120000 6 m00_w_data[3]
port 250 nsew signal output
rlabel metal2 s 308494 119200 308550 120000 6 m00_w_data[4]
port 251 nsew signal output
rlabel metal2 s 202878 0 202934 800 6 m00_w_data[5]
port 252 nsew signal output
rlabel metal2 s 454682 119200 454738 120000 6 m00_w_data[6]
port 253 nsew signal output
rlabel metal2 s 195150 0 195206 800 6 m00_w_data[7]
port 254 nsew signal output
rlabel metal2 s 407670 119200 407726 120000 6 m00_w_data[8]
port 255 nsew signal output
rlabel metal3 s 0 104048 800 104168 6 m00_w_data[9]
port 256 nsew signal output
rlabel metal3 s 479200 6128 480000 6248 6 m00_w_last
port 257 nsew signal output
rlabel metal3 s 479200 108128 480000 108248 6 m00_w_ready
port 258 nsew signal input
rlabel metal3 s 479200 70728 480000 70848 6 m00_w_strb[0]
port 259 nsew signal output
rlabel metal3 s 479200 3408 480000 3528 6 m00_w_strb[1]
port 260 nsew signal output
rlabel metal2 s 475934 0 475990 800 6 m00_w_strb[2]
port 261 nsew signal output
rlabel metal2 s 84382 119200 84438 120000 6 m00_w_strb[3]
port 262 nsew signal output
rlabel metal2 s 359370 0 359426 800 6 m00_w_user[-1]
port 263 nsew signal output
rlabel metal2 s 411534 119200 411590 120000 6 m00_w_user[0]
port 264 nsew signal output
rlabel metal2 s 155222 119200 155278 120000 6 m00_w_valid
port 265 nsew signal output
rlabel metal2 s 361946 119200 362002 120000 6 m01_ar_addr[0]
port 266 nsew signal output
rlabel metal2 s 216402 0 216458 800 6 m01_ar_addr[10]
port 267 nsew signal output
rlabel metal2 s 72146 0 72202 800 6 m01_ar_addr[11]
port 268 nsew signal output
rlabel metal2 s 15474 119200 15530 120000 6 m01_ar_addr[12]
port 269 nsew signal output
rlabel metal2 s 399298 0 399354 800 6 m01_ar_addr[13]
port 270 nsew signal output
rlabel metal2 s 439226 0 439282 800 6 m01_ar_addr[14]
port 271 nsew signal output
rlabel metal2 s 334254 0 334310 800 6 m01_ar_addr[15]
port 272 nsew signal output
rlabel metal2 s 466918 0 466974 800 6 m01_ar_addr[16]
port 273 nsew signal output
rlabel metal2 s 133970 119200 134026 120000 6 m01_ar_addr[17]
port 274 nsew signal output
rlabel metal2 s 389638 0 389694 800 6 m01_ar_addr[18]
port 275 nsew signal output
rlabel metal2 s 421838 119200 421894 120000 6 m01_ar_addr[19]
port 276 nsew signal output
rlabel metal2 s 212538 0 212594 800 6 m01_ar_addr[1]
port 277 nsew signal output
rlabel metal2 s 450174 0 450230 800 6 m01_ar_addr[20]
port 278 nsew signal output
rlabel metal2 s 437294 119200 437350 120000 6 m01_ar_addr[21]
port 279 nsew signal output
rlabel metal2 s 360014 119200 360070 120000 6 m01_ar_addr[22]
port 280 nsew signal output
rlabel metal3 s 0 10208 800 10328 6 m01_ar_addr[23]
port 281 nsew signal output
rlabel metal2 s 380622 119200 380678 120000 6 m01_ar_addr[24]
port 282 nsew signal output
rlabel metal3 s 0 63928 800 64048 6 m01_ar_addr[25]
port 283 nsew signal output
rlabel metal2 s 38658 0 38714 800 6 m01_ar_addr[26]
port 284 nsew signal output
rlabel metal2 s 436650 119200 436706 120000 6 m01_ar_addr[27]
port 285 nsew signal output
rlabel metal2 s 330390 119200 330446 120000 6 m01_ar_addr[28]
port 286 nsew signal output
rlabel metal2 s 452106 119200 452162 120000 6 m01_ar_addr[29]
port 287 nsew signal output
rlabel metal2 s 22558 0 22614 800 6 m01_ar_addr[2]
port 288 nsew signal output
rlabel metal2 s 278226 0 278282 800 6 m01_ar_addr[30]
port 289 nsew signal output
rlabel metal2 s 338118 0 338174 800 6 m01_ar_addr[31]
port 290 nsew signal output
rlabel metal2 s 349066 0 349122 800 6 m01_ar_addr[3]
port 291 nsew signal output
rlabel metal2 s 52182 119200 52238 120000 6 m01_ar_addr[4]
port 292 nsew signal output
rlabel metal3 s 0 100648 800 100768 6 m01_ar_addr[5]
port 293 nsew signal output
rlabel metal2 s 352930 119200 352986 120000 6 m01_ar_addr[6]
port 294 nsew signal output
rlabel metal2 s 258906 0 258962 800 6 m01_ar_addr[7]
port 295 nsew signal output
rlabel metal2 s 81162 119200 81218 120000 6 m01_ar_addr[8]
port 296 nsew signal output
rlabel metal2 s 119802 0 119858 800 6 m01_ar_addr[9]
port 297 nsew signal output
rlabel metal2 s 322662 0 322718 800 6 m01_ar_burst[0]
port 298 nsew signal output
rlabel metal3 s 479200 31968 480000 32088 6 m01_ar_burst[1]
port 299 nsew signal output
rlabel metal2 s 260838 119200 260894 120000 6 m01_ar_cache[0]
port 300 nsew signal output
rlabel metal2 s 90178 119200 90234 120000 6 m01_ar_cache[1]
port 301 nsew signal output
rlabel metal2 s 157154 0 157210 800 6 m01_ar_cache[2]
port 302 nsew signal output
rlabel metal2 s 341338 0 341394 800 6 m01_ar_cache[3]
port 303 nsew signal output
rlabel metal2 s 345846 0 345902 800 6 m01_ar_id[0]
port 304 nsew signal output
rlabel metal3 s 479200 9528 480000 9648 6 m01_ar_id[10]
port 305 nsew signal output
rlabel metal3 s 479200 66648 480000 66768 6 m01_ar_id[11]
port 306 nsew signal output
rlabel metal2 s 314290 0 314346 800 6 m01_ar_id[1]
port 307 nsew signal output
rlabel metal3 s 0 116968 800 117088 6 m01_ar_id[2]
port 308 nsew signal output
rlabel metal3 s 479200 50328 480000 50448 6 m01_ar_id[3]
port 309 nsew signal output
rlabel metal2 s 473358 119200 473414 120000 6 m01_ar_id[4]
port 310 nsew signal output
rlabel metal2 s 269854 119200 269910 120000 6 m01_ar_id[5]
port 311 nsew signal output
rlabel metal2 s 376114 119200 376170 120000 6 m01_ar_id[6]
port 312 nsew signal output
rlabel metal2 s 86958 0 87014 800 6 m01_ar_id[7]
port 313 nsew signal output
rlabel metal2 s 470782 0 470838 800 6 m01_ar_id[8]
port 314 nsew signal output
rlabel metal2 s 439870 0 439926 800 6 m01_ar_id[9]
port 315 nsew signal output
rlabel metal2 s 56046 0 56102 800 6 m01_ar_len[0]
port 316 nsew signal output
rlabel metal3 s 479200 101328 480000 101448 6 m01_ar_len[1]
port 317 nsew signal output
rlabel metal3 s 0 89768 800 89888 6 m01_ar_len[2]
port 318 nsew signal output
rlabel metal2 s 89534 0 89590 800 6 m01_ar_len[3]
port 319 nsew signal output
rlabel metal2 s 464986 119200 465042 120000 6 m01_ar_len[4]
port 320 nsew signal output
rlabel metal3 s 479200 79568 480000 79688 6 m01_ar_len[5]
port 321 nsew signal output
rlabel metal2 s 240874 0 240930 800 6 m01_ar_len[6]
port 322 nsew signal output
rlabel metal2 s 332966 0 333022 800 6 m01_ar_len[7]
port 323 nsew signal output
rlabel metal2 s 146206 0 146262 800 6 m01_ar_lock
port 324 nsew signal output
rlabel metal2 s 184202 0 184258 800 6 m01_ar_prot[0]
port 325 nsew signal output
rlabel metal2 s 379334 0 379390 800 6 m01_ar_prot[1]
port 326 nsew signal output
rlabel metal3 s 0 25168 800 25288 6 m01_ar_prot[2]
port 327 nsew signal output
rlabel metal3 s 0 2048 800 2168 6 m01_ar_qos[0]
port 328 nsew signal output
rlabel metal2 s 68926 0 68982 800 6 m01_ar_qos[1]
port 329 nsew signal output
rlabel metal2 s 77298 119200 77354 120000 6 m01_ar_qos[2]
port 330 nsew signal output
rlabel metal2 s 212538 119200 212594 120000 6 m01_ar_qos[3]
port 331 nsew signal output
rlabel metal3 s 479200 40808 480000 40928 6 m01_ar_ready
port 332 nsew signal input
rlabel metal2 s 353574 119200 353630 120000 6 m01_ar_region[0]
port 333 nsew signal output
rlabel metal3 s 479200 61208 480000 61328 6 m01_ar_region[1]
port 334 nsew signal output
rlabel metal2 s 144918 119200 144974 120000 6 m01_ar_region[2]
port 335 nsew signal output
rlabel metal2 s 398654 119200 398710 120000 6 m01_ar_region[3]
port 336 nsew signal output
rlabel metal2 s 128818 119200 128874 120000 6 m01_ar_size[0]
port 337 nsew signal output
rlabel metal2 s 150714 119200 150770 120000 6 m01_ar_size[1]
port 338 nsew signal output
rlabel metal3 s 0 34008 800 34128 6 m01_ar_size[2]
port 339 nsew signal output
rlabel metal2 s 425702 119200 425758 120000 6 m01_ar_user[-1]
port 340 nsew signal output
rlabel metal2 s 454682 0 454738 800 6 m01_ar_user[0]
port 341 nsew signal output
rlabel metal2 s 369674 119200 369730 120000 6 m01_ar_valid
port 342 nsew signal output
rlabel metal2 s 416686 119200 416742 120000 6 m01_aw_addr[0]
port 343 nsew signal output
rlabel metal2 s 175186 119200 175242 120000 6 m01_aw_addr[10]
port 344 nsew signal output
rlabel metal2 s 13542 119200 13598 120000 6 m01_aw_addr[11]
port 345 nsew signal output
rlabel metal2 s 86314 0 86370 800 6 m01_aw_addr[12]
port 346 nsew signal output
rlabel metal2 s 132038 0 132094 800 6 m01_aw_addr[13]
port 347 nsew signal output
rlabel metal2 s 430210 119200 430266 120000 6 m01_aw_addr[14]
port 348 nsew signal output
rlabel metal2 s 95974 0 96030 800 6 m01_aw_addr[15]
port 349 nsew signal output
rlabel metal2 s 307850 0 307906 800 6 m01_aw_addr[16]
port 350 nsew signal output
rlabel metal2 s 21914 119200 21970 120000 6 m01_aw_addr[17]
port 351 nsew signal output
rlabel metal2 s 287886 119200 287942 120000 6 m01_aw_addr[18]
port 352 nsew signal output
rlabel metal2 s 6458 119200 6514 120000 6 m01_aw_addr[19]
port 353 nsew signal output
rlabel metal2 s 143630 0 143686 800 6 m01_aw_addr[1]
port 354 nsew signal output
rlabel metal2 s 379334 119200 379390 120000 6 m01_aw_addr[20]
port 355 nsew signal output
rlabel metal2 s 148138 0 148194 800 6 m01_aw_addr[21]
port 356 nsew signal output
rlabel metal2 s 470138 119200 470194 120000 6 m01_aw_addr[22]
port 357 nsew signal output
rlabel metal2 s 7746 0 7802 800 6 m01_aw_addr[23]
port 358 nsew signal output
rlabel metal3 s 0 56448 800 56568 6 m01_aw_addr[24]
port 359 nsew signal output
rlabel metal2 s 94686 0 94742 800 6 m01_aw_addr[25]
port 360 nsew signal output
rlabel metal3 s 479200 115608 480000 115728 6 m01_aw_addr[26]
port 361 nsew signal output
rlabel metal2 s 372250 0 372306 800 6 m01_aw_addr[27]
port 362 nsew signal output
rlabel metal3 s 0 66648 800 66768 6 m01_aw_addr[28]
port 363 nsew signal output
rlabel metal2 s 75366 119200 75422 120000 6 m01_aw_addr[29]
port 364 nsew signal output
rlabel metal2 s 404450 0 404506 800 6 m01_aw_addr[2]
port 365 nsew signal output
rlabel metal2 s 27710 119200 27766 120000 6 m01_aw_addr[30]
port 366 nsew signal output
rlabel metal3 s 0 85688 800 85808 6 m01_aw_addr[31]
port 367 nsew signal output
rlabel metal2 s 374182 0 374238 800 6 m01_aw_addr[3]
port 368 nsew signal output
rlabel metal2 s 47674 0 47730 800 6 m01_aw_addr[4]
port 369 nsew signal output
rlabel metal2 s 361302 0 361358 800 6 m01_aw_addr[5]
port 370 nsew signal output
rlabel metal2 s 64418 119200 64474 120000 6 m01_aw_addr[6]
port 371 nsew signal output
rlabel metal2 s 144918 0 144974 800 6 m01_aw_addr[7]
port 372 nsew signal output
rlabel metal2 s 381910 119200 381966 120000 6 m01_aw_addr[8]
port 373 nsew signal output
rlabel metal2 s 98550 119200 98606 120000 6 m01_aw_addr[9]
port 374 nsew signal output
rlabel metal2 s 255042 0 255098 800 6 m01_aw_burst[0]
port 375 nsew signal output
rlabel metal3 s 479200 38768 480000 38888 6 m01_aw_burst[1]
port 376 nsew signal output
rlabel metal2 s 93398 119200 93454 120000 6 m01_aw_cache[0]
port 377 nsew signal output
rlabel metal3 s 0 87048 800 87168 6 m01_aw_cache[1]
port 378 nsew signal output
rlabel metal2 s 471426 0 471482 800 6 m01_aw_cache[2]
port 379 nsew signal output
rlabel metal2 s 387062 0 387118 800 6 m01_aw_cache[3]
port 380 nsew signal output
rlabel metal2 s 185490 0 185546 800 6 m01_aw_id[0]
port 381 nsew signal output
rlabel metal3 s 479200 96568 480000 96688 6 m01_aw_id[10]
port 382 nsew signal output
rlabel metal2 s 71502 119200 71558 120000 6 m01_aw_id[11]
port 383 nsew signal output
rlabel metal2 s 322018 119200 322074 120000 6 m01_aw_id[1]
port 384 nsew signal output
rlabel metal3 s 479200 49648 480000 49768 6 m01_aw_id[2]
port 385 nsew signal output
rlabel metal2 s 170678 0 170734 800 6 m01_aw_id[3]
port 386 nsew signal output
rlabel metal2 s 342626 119200 342682 120000 6 m01_aw_id[4]
port 387 nsew signal output
rlabel metal2 s 273074 119200 273130 120000 6 m01_aw_id[5]
port 388 nsew signal output
rlabel metal2 s 43166 119200 43222 120000 6 m01_aw_id[6]
port 389 nsew signal output
rlabel metal2 s 338118 119200 338174 120000 6 m01_aw_id[7]
port 390 nsew signal output
rlabel metal2 s 327814 119200 327870 120000 6 m01_aw_id[8]
port 391 nsew signal output
rlabel metal2 s 12254 119200 12310 120000 6 m01_aw_id[9]
port 392 nsew signal output
rlabel metal3 s 0 77528 800 77648 6 m01_aw_len[0]
port 393 nsew signal output
rlabel metal2 s 450818 0 450874 800 6 m01_aw_len[1]
port 394 nsew signal output
rlabel metal2 s 346490 119200 346546 120000 6 m01_aw_len[2]
port 395 nsew signal output
rlabel metal3 s 479200 57808 480000 57928 6 m01_aw_len[3]
port 396 nsew signal output
rlabel metal2 s 456614 0 456670 800 6 m01_aw_len[4]
port 397 nsew signal output
rlabel metal2 s 104346 0 104402 800 6 m01_aw_len[5]
port 398 nsew signal output
rlabel metal2 s 135258 119200 135314 120000 6 m01_aw_len[6]
port 399 nsew signal output
rlabel metal2 s 309138 119200 309194 120000 6 m01_aw_len[7]
port 400 nsew signal output
rlabel metal2 s 22558 119200 22614 120000 6 m01_aw_lock
port 401 nsew signal output
rlabel metal2 s 387706 119200 387762 120000 6 m01_aw_prot[0]
port 402 nsew signal output
rlabel metal2 s 371606 0 371662 800 6 m01_aw_prot[1]
port 403 nsew signal output
rlabel metal2 s 439870 119200 439926 120000 6 m01_aw_prot[2]
port 404 nsew signal output
rlabel metal2 s 392858 119200 392914 120000 6 m01_aw_qos[0]
port 405 nsew signal output
rlabel metal2 s 341982 119200 342038 120000 6 m01_aw_qos[1]
port 406 nsew signal output
rlabel metal2 s 152002 0 152058 800 6 m01_aw_qos[2]
port 407 nsew signal output
rlabel metal3 s 0 60528 800 60648 6 m01_aw_qos[3]
port 408 nsew signal output
rlabel metal2 s 287242 0 287298 800 6 m01_aw_ready
port 409 nsew signal input
rlabel metal2 s 339406 0 339462 800 6 m01_aw_region[0]
port 410 nsew signal output
rlabel metal2 s 479798 119200 479854 120000 6 m01_aw_region[1]
port 411 nsew signal output
rlabel metal2 s 79874 119200 79930 120000 6 m01_aw_region[2]
port 412 nsew signal output
rlabel metal2 s 231214 119200 231270 120000 6 m01_aw_region[3]
port 413 nsew signal output
rlabel metal2 s 85670 119200 85726 120000 6 m01_aw_size[0]
port 414 nsew signal output
rlabel metal2 s 271142 0 271198 800 6 m01_aw_size[1]
port 415 nsew signal output
rlabel metal2 s 223486 119200 223542 120000 6 m01_aw_size[2]
port 416 nsew signal output
rlabel metal2 s 456614 119200 456670 120000 6 m01_aw_user[-1]
port 417 nsew signal output
rlabel metal2 s 94042 0 94098 800 6 m01_aw_user[0]
port 418 nsew signal output
rlabel metal2 s 126242 0 126298 800 6 m01_aw_valid
port 419 nsew signal output
rlabel metal2 s 290462 0 290518 800 6 m01_b_id[0]
port 420 nsew signal input
rlabel metal3 s 479200 109488 480000 109608 6 m01_b_id[10]
port 421 nsew signal input
rlabel metal2 s 144274 0 144330 800 6 m01_b_id[11]
port 422 nsew signal input
rlabel metal3 s 0 47608 800 47728 6 m01_b_id[1]
port 423 nsew signal input
rlabel metal2 s 176474 0 176530 800 6 m01_b_id[2]
port 424 nsew signal input
rlabel metal2 s 112074 0 112130 800 6 m01_b_id[3]
port 425 nsew signal input
rlabel metal2 s 173254 119200 173310 120000 6 m01_b_id[4]
port 426 nsew signal input
rlabel metal3 s 479200 60528 480000 60648 6 m01_b_id[5]
port 427 nsew signal input
rlabel metal2 s 47030 119200 47086 120000 6 m01_b_id[6]
port 428 nsew signal input
rlabel metal2 s 193862 119200 193918 120000 6 m01_b_id[7]
port 429 nsew signal input
rlabel metal2 s 180982 0 181038 800 6 m01_b_id[8]
port 430 nsew signal input
rlabel metal3 s 0 48968 800 49088 6 m01_b_id[9]
port 431 nsew signal input
rlabel metal2 s 157798 119200 157854 120000 6 m01_b_ready
port 432 nsew signal output
rlabel metal2 s 446310 0 446366 800 6 m01_b_resp[0]
port 433 nsew signal input
rlabel metal3 s 0 11568 800 11688 6 m01_b_resp[1]
port 434 nsew signal input
rlabel metal2 s 407026 119200 407082 120000 6 m01_b_user[-1]
port 435 nsew signal input
rlabel metal2 s 41878 119200 41934 120000 6 m01_b_user[0]
port 436 nsew signal input
rlabel metal2 s 385130 0 385186 800 6 m01_b_valid
port 437 nsew signal input
rlabel metal3 s 0 78888 800 79008 6 m01_r_data[0]
port 438 nsew signal input
rlabel metal2 s 44454 0 44510 800 6 m01_r_data[10]
port 439 nsew signal input
rlabel metal2 s 301410 0 301466 800 6 m01_r_data[11]
port 440 nsew signal input
rlabel metal2 s 77942 119200 77998 120000 6 m01_r_data[12]
port 441 nsew signal input
rlabel metal2 s 269854 0 269910 800 6 m01_r_data[13]
port 442 nsew signal input
rlabel metal2 s 236366 0 236422 800 6 m01_r_data[14]
port 443 nsew signal input
rlabel metal3 s 0 91808 800 91928 6 m01_r_data[15]
port 444 nsew signal input
rlabel metal2 s 376758 0 376814 800 6 m01_r_data[16]
port 445 nsew signal input
rlabel metal2 s 205454 119200 205510 120000 6 m01_r_data[17]
port 446 nsew signal input
rlabel metal2 s 464986 0 465042 800 6 m01_r_data[18]
port 447 nsew signal input
rlabel metal2 s 104990 119200 105046 120000 6 m01_r_data[19]
port 448 nsew signal input
rlabel metal2 s 391570 119200 391626 120000 6 m01_r_data[1]
port 449 nsew signal input
rlabel metal2 s 307850 119200 307906 120000 6 m01_r_data[20]
port 450 nsew signal input
rlabel metal2 s 141054 119200 141110 120000 6 m01_r_data[21]
port 451 nsew signal input
rlabel metal2 s 436006 0 436062 800 6 m01_r_data[22]
port 452 nsew signal input
rlabel metal3 s 0 76168 800 76288 6 m01_r_data[23]
port 453 nsew signal input
rlabel metal2 s 240230 119200 240286 120000 6 m01_r_data[24]
port 454 nsew signal input
rlabel metal2 s 463698 119200 463754 120000 6 m01_r_data[25]
port 455 nsew signal input
rlabel metal3 s 479200 93848 480000 93968 6 m01_r_data[26]
port 456 nsew signal input
rlabel metal2 s 378046 119200 378102 120000 6 m01_r_data[27]
port 457 nsew signal input
rlabel metal3 s 0 36048 800 36168 6 m01_r_data[28]
port 458 nsew signal input
rlabel metal2 s 424414 119200 424470 120000 6 m01_r_data[29]
port 459 nsew signal input
rlabel metal2 s 315578 119200 315634 120000 6 m01_r_data[2]
port 460 nsew signal input
rlabel metal2 s 273718 119200 273774 120000 6 m01_r_data[30]
port 461 nsew signal input
rlabel metal2 s 107566 0 107622 800 6 m01_r_data[31]
port 462 nsew signal input
rlabel metal2 s 271786 119200 271842 120000 6 m01_r_data[3]
port 463 nsew signal input
rlabel metal2 s 237010 119200 237066 120000 6 m01_r_data[4]
port 464 nsew signal input
rlabel metal2 s 273074 0 273130 800 6 m01_r_data[5]
port 465 nsew signal input
rlabel metal2 s 372250 119200 372306 120000 6 m01_r_data[6]
port 466 nsew signal input
rlabel metal3 s 0 8168 800 8288 6 m01_r_data[7]
port 467 nsew signal input
rlabel metal2 s 319442 119200 319498 120000 6 m01_r_data[8]
port 468 nsew signal input
rlabel metal2 s 238298 0 238354 800 6 m01_r_data[9]
port 469 nsew signal input
rlabel metal2 s 198370 119200 198426 120000 6 m01_r_id[0]
port 470 nsew signal input
rlabel metal2 s 39946 0 40002 800 6 m01_r_id[10]
port 471 nsew signal input
rlabel metal2 s 349710 119200 349766 120000 6 m01_r_id[11]
port 472 nsew signal input
rlabel metal2 s 128174 0 128230 800 6 m01_r_id[1]
port 473 nsew signal input
rlabel metal2 s 184846 119200 184902 120000 6 m01_r_id[2]
port 474 nsew signal input
rlabel metal2 s 426346 119200 426402 120000 6 m01_r_id[3]
port 475 nsew signal input
rlabel metal2 s 441158 0 441214 800 6 m01_r_id[4]
port 476 nsew signal input
rlabel metal2 s 242806 0 242862 800 6 m01_r_id[5]
port 477 nsew signal input
rlabel metal2 s 72146 119200 72202 120000 6 m01_r_id[6]
port 478 nsew signal input
rlabel metal2 s 82450 0 82506 800 6 m01_r_id[7]
port 479 nsew signal input
rlabel metal3 s 479200 102688 480000 102808 6 m01_r_id[8]
port 480 nsew signal input
rlabel metal2 s 220910 0 220966 800 6 m01_r_id[9]
port 481 nsew signal input
rlabel metal2 s 219622 119200 219678 120000 6 m01_r_last
port 482 nsew signal input
rlabel metal2 s 349710 0 349766 800 6 m01_r_ready
port 483 nsew signal output
rlabel metal2 s 91466 0 91522 800 6 m01_r_resp[0]
port 484 nsew signal input
rlabel metal2 s 25134 119200 25190 120000 6 m01_r_resp[1]
port 485 nsew signal input
rlabel metal3 s 479200 118328 480000 118448 6 m01_r_user[-1]
port 486 nsew signal input
rlabel metal2 s 166170 0 166226 800 6 m01_r_user[0]
port 487 nsew signal input
rlabel metal2 s 88890 0 88946 800 6 m01_r_valid
port 488 nsew signal input
rlabel metal2 s 90822 0 90878 800 6 m01_w_data[0]
port 489 nsew signal output
rlabel metal3 s 0 81608 800 81728 6 m01_w_data[10]
port 490 nsew signal output
rlabel metal2 s 405094 119200 405150 120000 6 m01_w_data[11]
port 491 nsew signal output
rlabel metal2 s 472714 119200 472770 120000 6 m01_w_data[12]
port 492 nsew signal output
rlabel metal2 s 61198 119200 61254 120000 6 m01_w_data[13]
port 493 nsew signal output
rlabel metal2 s 74078 119200 74134 120000 6 m01_w_data[14]
port 494 nsew signal output
rlabel metal2 s 176474 119200 176530 120000 6 m01_w_data[15]
port 495 nsew signal output
rlabel metal2 s 63774 119200 63830 120000 6 m01_w_data[16]
port 496 nsew signal output
rlabel metal2 s 209318 0 209374 800 6 m01_w_data[17]
port 497 nsew signal output
rlabel metal3 s 0 58488 800 58608 6 m01_w_data[18]
port 498 nsew signal output
rlabel metal2 s 429566 119200 429622 120000 6 m01_w_data[19]
port 499 nsew signal output
rlabel metal2 s 278870 119200 278926 120000 6 m01_w_data[1]
port 500 nsew signal output
rlabel metal2 s 246026 119200 246082 120000 6 m01_w_data[20]
port 501 nsew signal output
rlabel metal3 s 0 82288 800 82408 6 m01_w_data[21]
port 502 nsew signal output
rlabel metal2 s 29642 119200 29698 120000 6 m01_w_data[22]
port 503 nsew signal output
rlabel metal2 s 409602 119200 409658 120000 6 m01_w_data[23]
port 504 nsew signal output
rlabel metal2 s 63130 119200 63186 120000 6 m01_w_data[24]
port 505 nsew signal output
rlabel metal2 s 241518 119200 241574 120000 6 m01_w_data[25]
port 506 nsew signal output
rlabel metal2 s 21270 0 21326 800 6 m01_w_data[26]
port 507 nsew signal output
rlabel metal2 s 4526 0 4582 800 6 m01_w_data[27]
port 508 nsew signal output
rlabel metal2 s 475290 119200 475346 120000 6 m01_w_data[28]
port 509 nsew signal output
rlabel metal3 s 479200 89768 480000 89888 6 m01_w_data[29]
port 510 nsew signal output
rlabel metal2 s 152646 119200 152702 120000 6 m01_w_data[2]
port 511 nsew signal output
rlabel metal3 s 0 113568 800 113688 6 m01_w_data[30]
port 512 nsew signal output
rlabel metal2 s 182270 0 182326 800 6 m01_w_data[31]
port 513 nsew signal output
rlabel metal2 s 23846 0 23902 800 6 m01_w_data[3]
port 514 nsew signal output
rlabel metal2 s 419906 119200 419962 120000 6 m01_w_data[4]
port 515 nsew signal output
rlabel metal2 s 222842 0 222898 800 6 m01_w_data[5]
port 516 nsew signal output
rlabel metal2 s 163594 119200 163650 120000 6 m01_w_data[6]
port 517 nsew signal output
rlabel metal3 s 0 49648 800 49768 6 m01_w_data[7]
port 518 nsew signal output
rlabel metal2 s 382554 0 382610 800 6 m01_w_data[8]
port 519 nsew signal output
rlabel metal3 s 479200 44208 480000 44328 6 m01_w_data[9]
port 520 nsew signal output
rlabel metal2 s 150070 0 150126 800 6 m01_w_last
port 521 nsew signal output
rlabel metal3 s 479200 63928 480000 64048 6 m01_w_ready
port 522 nsew signal input
rlabel metal3 s 0 94528 800 94648 6 m01_w_strb[0]
port 523 nsew signal output
rlabel metal2 s 149426 0 149482 800 6 m01_w_strb[1]
port 524 nsew signal output
rlabel metal2 s 397366 119200 397422 120000 6 m01_w_strb[2]
port 525 nsew signal output
rlabel metal2 s 345846 119200 345902 120000 6 m01_w_strb[3]
port 526 nsew signal output
rlabel metal2 s 470782 119200 470838 120000 6 m01_w_user[-1]
port 527 nsew signal output
rlabel metal2 s 132682 119200 132738 120000 6 m01_w_user[0]
port 528 nsew signal output
rlabel metal2 s 199014 119200 199070 120000 6 m01_w_valid
port 529 nsew signal output
rlabel metal2 s 313002 0 313058 800 6 m02_ar_addr[0]
port 530 nsew signal output
rlabel metal2 s 468850 0 468906 800 6 m02_ar_addr[10]
port 531 nsew signal output
rlabel metal2 s 281446 119200 281502 120000 6 m02_ar_addr[11]
port 532 nsew signal output
rlabel metal2 s 66994 119200 67050 120000 6 m02_ar_addr[12]
port 533 nsew signal output
rlabel metal2 s 12898 119200 12954 120000 6 m02_ar_addr[13]
port 534 nsew signal output
rlabel metal2 s 18050 0 18106 800 6 m02_ar_addr[14]
port 535 nsew signal output
rlabel metal2 s 349066 119200 349122 120000 6 m02_ar_addr[15]
port 536 nsew signal output
rlabel metal3 s 0 29248 800 29368 6 m02_ar_addr[16]
port 537 nsew signal output
rlabel metal3 s 479200 26528 480000 26648 6 m02_ar_addr[17]
port 538 nsew signal output
rlabel metal2 s 443090 119200 443146 120000 6 m02_ar_addr[18]
port 539 nsew signal output
rlabel metal2 s 114650 119200 114706 120000 6 m02_ar_addr[19]
port 540 nsew signal output
rlabel metal2 s 76010 119200 76066 120000 6 m02_ar_addr[1]
port 541 nsew signal output
rlabel metal3 s 479200 58488 480000 58608 6 m02_ar_addr[20]
port 542 nsew signal output
rlabel metal2 s 433430 0 433486 800 6 m02_ar_addr[21]
port 543 nsew signal output
rlabel metal2 s 459190 0 459246 800 6 m02_ar_addr[22]
port 544 nsew signal output
rlabel metal2 s 218978 119200 219034 120000 6 m02_ar_addr[23]
port 545 nsew signal output
rlabel metal2 s 172610 0 172666 800 6 m02_ar_addr[24]
port 546 nsew signal output
rlabel metal2 s 17406 119200 17462 120000 6 m02_ar_addr[25]
port 547 nsew signal output
rlabel metal2 s 384486 119200 384542 120000 6 m02_ar_addr[26]
port 548 nsew signal output
rlabel metal3 s 0 4768 800 4888 6 m02_ar_addr[27]
port 549 nsew signal output
rlabel metal2 s 67638 119200 67694 120000 6 m02_ar_addr[28]
port 550 nsew signal output
rlabel metal2 s 380622 0 380678 800 6 m02_ar_addr[29]
port 551 nsew signal output
rlabel metal2 s 359370 119200 359426 120000 6 m02_ar_addr[2]
port 552 nsew signal output
rlabel metal2 s 67638 0 67694 800 6 m02_ar_addr[30]
port 553 nsew signal output
rlabel metal2 s 114006 0 114062 800 6 m02_ar_addr[31]
port 554 nsew signal output
rlabel metal2 s 236366 119200 236422 120000 6 m02_ar_addr[3]
port 555 nsew signal output
rlabel metal2 s 254398 0 254454 800 6 m02_ar_addr[4]
port 556 nsew signal output
rlabel metal2 s 344558 0 344614 800 6 m02_ar_addr[5]
port 557 nsew signal output
rlabel metal2 s 140410 119200 140466 120000 6 m02_ar_addr[6]
port 558 nsew signal output
rlabel metal2 s 131394 0 131450 800 6 m02_ar_addr[7]
port 559 nsew signal output
rlabel metal2 s 118514 0 118570 800 6 m02_ar_addr[8]
port 560 nsew signal output
rlabel metal2 s 295614 119200 295670 120000 6 m02_ar_addr[9]
port 561 nsew signal output
rlabel metal2 s 211894 119200 211950 120000 6 m02_ar_burst[0]
port 562 nsew signal output
rlabel metal2 s 298834 0 298890 800 6 m02_ar_burst[1]
port 563 nsew signal output
rlabel metal2 s 356794 119200 356850 120000 6 m02_ar_cache[0]
port 564 nsew signal output
rlabel metal2 s 376758 119200 376814 120000 6 m02_ar_cache[1]
port 565 nsew signal output
rlabel metal2 s 37370 119200 37426 120000 6 m02_ar_cache[2]
port 566 nsew signal output
rlabel metal2 s 459190 119200 459246 120000 6 m02_ar_cache[3]
port 567 nsew signal output
rlabel metal2 s 154578 0 154634 800 6 m02_ar_id[0]
port 568 nsew signal output
rlabel metal2 s 32862 0 32918 800 6 m02_ar_id[10]
port 569 nsew signal output
rlabel metal2 s 305274 119200 305330 120000 6 m02_ar_id[11]
port 570 nsew signal output
rlabel metal3 s 0 99968 800 100088 6 m02_ar_id[1]
port 571 nsew signal output
rlabel metal2 s 99194 0 99250 800 6 m02_ar_id[2]
port 572 nsew signal output
rlabel metal2 s 177118 119200 177174 120000 6 m02_ar_id[3]
port 573 nsew signal output
rlabel metal2 s 168746 0 168802 800 6 m02_ar_id[4]
port 574 nsew signal output
rlabel metal2 s 202234 0 202290 800 6 m02_ar_id[5]
port 575 nsew signal output
rlabel metal2 s 195150 119200 195206 120000 6 m02_ar_id[6]
port 576 nsew signal output
rlabel metal2 s 390926 119200 390982 120000 6 m02_ar_id[7]
port 577 nsew signal output
rlabel metal2 s 74078 0 74134 800 6 m02_ar_id[8]
port 578 nsew signal output
rlabel metal2 s 302054 119200 302110 120000 6 m02_ar_id[9]
port 579 nsew signal output
rlabel metal2 s 21270 119200 21326 120000 6 m02_ar_len[0]
port 580 nsew signal output
rlabel metal2 s 273718 0 273774 800 6 m02_ar_len[1]
port 581 nsew signal output
rlabel metal2 s 47030 0 47086 800 6 m02_ar_len[2]
port 582 nsew signal output
rlabel metal2 s 200946 0 201002 800 6 m02_ar_len[3]
port 583 nsew signal output
rlabel metal2 s 174542 0 174598 800 6 m02_ar_len[4]
port 584 nsew signal output
rlabel metal2 s 95330 119200 95386 120000 6 m02_ar_len[5]
port 585 nsew signal output
rlabel metal2 s 24490 0 24546 800 6 m02_ar_len[6]
port 586 nsew signal output
rlabel metal2 s 423126 0 423182 800 6 m02_ar_len[7]
port 587 nsew signal output
rlabel metal2 s 427634 0 427690 800 6 m02_ar_lock
port 588 nsew signal output
rlabel metal3 s 479200 14968 480000 15088 6 m02_ar_prot[0]
port 589 nsew signal output
rlabel metal2 s 443734 119200 443790 120000 6 m02_ar_prot[1]
port 590 nsew signal output
rlabel metal2 s 119158 119200 119214 120000 6 m02_ar_prot[2]
port 591 nsew signal output
rlabel metal2 s 317510 119200 317566 120000 6 m02_ar_qos[0]
port 592 nsew signal output
rlabel metal2 s 405738 0 405794 800 6 m02_ar_qos[1]
port 593 nsew signal output
rlabel metal2 s 173254 0 173310 800 6 m02_ar_qos[2]
port 594 nsew signal output
rlabel metal2 s 263414 0 263470 800 6 m02_ar_qos[3]
port 595 nsew signal output
rlabel metal2 s 275006 119200 275062 120000 6 m02_ar_ready
port 596 nsew signal input
rlabel metal2 s 284022 0 284078 800 6 m02_ar_region[0]
port 597 nsew signal output
rlabel metal3 s 0 82968 800 83088 6 m02_ar_region[1]
port 598 nsew signal output
rlabel metal2 s 166814 119200 166870 120000 6 m02_ar_region[2]
port 599 nsew signal output
rlabel metal2 s 448242 119200 448298 120000 6 m02_ar_region[3]
port 600 nsew signal output
rlabel metal2 s 317510 0 317566 800 6 m02_ar_size[0]
port 601 nsew signal output
rlabel metal2 s 98550 0 98606 800 6 m02_ar_size[1]
port 602 nsew signal output
rlabel metal2 s 287886 0 287942 800 6 m02_ar_size[2]
port 603 nsew signal output
rlabel metal2 s 143630 119200 143686 120000 6 m02_ar_user[-1]
port 604 nsew signal output
rlabel metal3 s 0 19728 800 19848 6 m02_ar_user[0]
port 605 nsew signal output
rlabel metal3 s 0 112888 800 113008 6 m02_ar_valid
port 606 nsew signal output
rlabel metal2 s 446954 0 447010 800 6 m02_aw_addr[0]
port 607 nsew signal output
rlabel metal3 s 479200 83648 480000 83768 6 m02_aw_addr[10]
port 608 nsew signal output
rlabel metal2 s 46386 119200 46442 120000 6 m02_aw_addr[11]
port 609 nsew signal output
rlabel metal3 s 479200 47608 480000 47728 6 m02_aw_addr[12]
port 610 nsew signal output
rlabel metal3 s 0 80248 800 80368 6 m02_aw_addr[13]
port 611 nsew signal output
rlabel metal2 s 119802 119200 119858 120000 6 m02_aw_addr[14]
port 612 nsew signal output
rlabel metal2 s 472070 0 472126 800 6 m02_aw_addr[15]
port 613 nsew signal output
rlabel metal2 s 294970 119200 295026 120000 6 m02_aw_addr[16]
port 614 nsew signal output
rlabel metal2 s 39946 119200 40002 120000 6 m02_aw_addr[17]
port 615 nsew signal output
rlabel metal2 s 469494 0 469550 800 6 m02_aw_addr[18]
port 616 nsew signal output
rlabel metal2 s 417330 0 417386 800 6 m02_aw_addr[19]
port 617 nsew signal output
rlabel metal2 s 211250 119200 211306 120000 6 m02_aw_addr[1]
port 618 nsew signal output
rlabel metal2 s 1950 119200 2006 120000 6 m02_aw_addr[20]
port 619 nsew signal output
rlabel metal2 s 261482 0 261538 800 6 m02_aw_addr[21]
port 620 nsew signal output
rlabel metal2 s 148138 119200 148194 120000 6 m02_aw_addr[22]
port 621 nsew signal output
rlabel metal2 s 62486 119200 62542 120000 6 m02_aw_addr[23]
port 622 nsew signal output
rlabel metal3 s 479200 14288 480000 14408 6 m02_aw_addr[24]
port 623 nsew signal output
rlabel metal3 s 479200 85688 480000 85808 6 m02_aw_addr[25]
port 624 nsew signal output
rlabel metal2 s 340050 119200 340106 120000 6 m02_aw_addr[26]
port 625 nsew signal output
rlabel metal3 s 479200 45568 480000 45688 6 m02_aw_addr[27]
port 626 nsew signal output
rlabel metal2 s 137190 119200 137246 120000 6 m02_aw_addr[28]
port 627 nsew signal output
rlabel metal2 s 471426 119200 471482 120000 6 m02_aw_addr[29]
port 628 nsew signal output
rlabel metal2 s 414754 0 414810 800 6 m02_aw_addr[2]
port 629 nsew signal output
rlabel metal2 s 39302 0 39358 800 6 m02_aw_addr[30]
port 630 nsew signal output
rlabel metal3 s 0 44888 800 45008 6 m02_aw_addr[31]
port 631 nsew signal output
rlabel metal2 s 253754 119200 253810 120000 6 m02_aw_addr[3]
port 632 nsew signal output
rlabel metal2 s 208674 119200 208730 120000 6 m02_aw_addr[4]
port 633 nsew signal output
rlabel metal2 s 191930 0 191986 800 6 m02_aw_addr[5]
port 634 nsew signal output
rlabel metal2 s 347134 119200 347190 120000 6 m02_aw_addr[6]
port 635 nsew signal output
rlabel metal2 s 34794 119200 34850 120000 6 m02_aw_addr[7]
port 636 nsew signal output
rlabel metal2 s 282090 0 282146 800 6 m02_aw_addr[8]
port 637 nsew signal output
rlabel metal2 s 418618 119200 418674 120000 6 m02_aw_addr[9]
port 638 nsew signal output
rlabel metal3 s 479200 5448 480000 5568 6 m02_aw_burst[0]
port 639 nsew signal output
rlabel metal2 s 361946 0 362002 800 6 m02_aw_burst[1]
port 640 nsew signal output
rlabel metal3 s 0 115608 800 115728 6 m02_aw_cache[0]
port 641 nsew signal output
rlabel metal2 s 401230 0 401286 800 6 m02_aw_cache[1]
port 642 nsew signal output
rlabel metal3 s 479200 95208 480000 95328 6 m02_aw_cache[2]
port 643 nsew signal output
rlabel metal2 s 375470 0 375526 800 6 m02_aw_cache[3]
port 644 nsew signal output
rlabel metal2 s 57334 0 57390 800 6 m02_aw_id[0]
port 645 nsew signal output
rlabel metal2 s 363234 0 363290 800 6 m02_aw_id[10]
port 646 nsew signal output
rlabel metal2 s 233790 119200 233846 120000 6 m02_aw_id[11]
port 647 nsew signal output
rlabel metal2 s 280802 0 280858 800 6 m02_aw_id[1]
port 648 nsew signal output
rlabel metal2 s 405738 119200 405794 120000 6 m02_aw_id[2]
port 649 nsew signal output
rlabel metal2 s 337474 119200 337530 120000 6 m02_aw_id[3]
port 650 nsew signal output
rlabel metal3 s 0 80928 800 81048 6 m02_aw_id[4]
port 651 nsew signal output
rlabel metal2 s 159086 119200 159142 120000 6 m02_aw_id[5]
port 652 nsew signal output
rlabel metal2 s 72790 119200 72846 120000 6 m02_aw_id[6]
port 653 nsew signal output
rlabel metal3 s 0 87728 800 87848 6 m02_aw_id[7]
port 654 nsew signal output
rlabel metal2 s 54758 0 54814 800 6 m02_aw_id[8]
port 655 nsew signal output
rlabel metal2 s 55402 119200 55458 120000 6 m02_aw_id[9]
port 656 nsew signal output
rlabel metal3 s 0 51008 800 51128 6 m02_aw_len[0]
port 657 nsew signal output
rlabel metal2 s 123666 0 123722 800 6 m02_aw_len[1]
port 658 nsew signal output
rlabel metal2 s 227994 119200 228050 120000 6 m02_aw_len[2]
port 659 nsew signal output
rlabel metal3 s 0 25848 800 25968 6 m02_aw_len[3]
port 660 nsew signal output
rlabel metal2 s 294326 119200 294382 120000 6 m02_aw_len[4]
port 661 nsew signal output
rlabel metal2 s 4526 119200 4582 120000 6 m02_aw_len[5]
port 662 nsew signal output
rlabel metal2 s 391570 0 391626 800 6 m02_aw_len[6]
port 663 nsew signal output
rlabel metal2 s 242162 0 242218 800 6 m02_aw_len[7]
port 664 nsew signal output
rlabel metal3 s 479200 41488 480000 41608 6 m02_aw_lock
port 665 nsew signal output
rlabel metal2 s 188710 119200 188766 120000 6 m02_aw_prot[0]
port 666 nsew signal output
rlabel metal2 s 190642 119200 190698 120000 6 m02_aw_prot[1]
port 667 nsew signal output
rlabel metal2 s 177118 0 177174 800 6 m02_aw_prot[2]
port 668 nsew signal output
rlabel metal3 s 0 111528 800 111648 6 m02_aw_qos[0]
port 669 nsew signal output
rlabel metal2 s 194506 119200 194562 120000 6 m02_aw_qos[1]
port 670 nsew signal output
rlabel metal3 s 479200 110848 480000 110968 6 m02_aw_qos[2]
port 671 nsew signal output
rlabel metal2 s 463054 0 463110 800 6 m02_aw_qos[3]
port 672 nsew signal output
rlabel metal2 s 472070 119200 472126 120000 6 m02_aw_ready
port 673 nsew signal input
rlabel metal3 s 479200 86368 480000 86488 6 m02_aw_region[0]
port 674 nsew signal output
rlabel metal2 s 416686 0 416742 800 6 m02_aw_region[1]
port 675 nsew signal output
rlabel metal2 s 452106 0 452162 800 6 m02_aw_region[2]
port 676 nsew signal output
rlabel metal2 s 162306 119200 162362 120000 6 m02_aw_region[3]
port 677 nsew signal output
rlabel metal2 s 164882 119200 164938 120000 6 m02_aw_size[0]
port 678 nsew signal output
rlabel metal2 s 210606 119200 210662 120000 6 m02_aw_size[1]
port 679 nsew signal output
rlabel metal3 s 0 105408 800 105528 6 m02_aw_size[2]
port 680 nsew signal output
rlabel metal3 s 0 117648 800 117768 6 m02_aw_user[-1]
port 681 nsew signal output
rlabel metal2 s 120446 0 120502 800 6 m02_aw_user[0]
port 682 nsew signal output
rlabel metal2 s 447598 119200 447654 120000 6 m02_aw_valid
port 683 nsew signal output
rlabel metal2 s 332322 119200 332378 120000 6 m02_b_id[0]
port 684 nsew signal input
rlabel metal2 s 31574 119200 31630 120000 6 m02_b_id[10]
port 685 nsew signal input
rlabel metal2 s 220910 119200 220966 120000 6 m02_b_id[11]
port 686 nsew signal input
rlabel metal3 s 0 7488 800 7608 6 m02_b_id[1]
port 687 nsew signal input
rlabel metal3 s 0 40808 800 40928 6 m02_b_id[2]
port 688 nsew signal input
rlabel metal2 s 289818 119200 289874 120000 6 m02_b_id[3]
port 689 nsew signal input
rlabel metal2 s 50250 119200 50306 120000 6 m02_b_id[4]
port 690 nsew signal input
rlabel metal2 s 311714 119200 311770 120000 6 m02_b_id[5]
port 691 nsew signal input
rlabel metal3 s 479200 74808 480000 74928 6 m02_b_id[6]
port 692 nsew signal input
rlabel metal2 s 368386 0 368442 800 6 m02_b_id[7]
port 693 nsew signal input
rlabel metal2 s 227350 119200 227406 120000 6 m02_b_id[8]
port 694 nsew signal input
rlabel metal2 s 455326 119200 455382 120000 6 m02_b_id[9]
port 695 nsew signal input
rlabel metal2 s 443090 0 443146 800 6 m02_b_ready
port 696 nsew signal output
rlabel metal3 s 0 34688 800 34808 6 m02_b_resp[0]
port 697 nsew signal input
rlabel metal2 s 459834 0 459890 800 6 m02_b_resp[1]
port 698 nsew signal input
rlabel metal2 s 244094 119200 244150 120000 6 m02_b_user[-1]
port 699 nsew signal input
rlabel metal2 s 34150 119200 34206 120000 6 m02_b_user[0]
port 700 nsew signal input
rlabel metal2 s 159730 119200 159786 120000 6 m02_b_valid
port 701 nsew signal input
rlabel metal3 s 0 55768 800 55888 6 m02_r_data[0]
port 702 nsew signal input
rlabel metal2 s 76010 0 76066 800 6 m02_r_data[10]
port 703 nsew signal input
rlabel metal3 s 479200 39448 480000 39568 6 m02_r_data[11]
port 704 nsew signal input
rlabel metal2 s 449530 119200 449586 120000 6 m02_r_data[12]
port 705 nsew signal input
rlabel metal2 s 378690 0 378746 800 6 m02_r_data[13]
port 706 nsew signal input
rlabel metal2 s 188066 0 188122 800 6 m02_r_data[14]
port 707 nsew signal input
rlabel metal2 s 293038 0 293094 800 6 m02_r_data[15]
port 708 nsew signal input
rlabel metal2 s 10322 119200 10378 120000 6 m02_r_data[16]
port 709 nsew signal input
rlabel metal2 s 397366 0 397422 800 6 m02_r_data[17]
port 710 nsew signal input
rlabel metal2 s 237654 0 237710 800 6 m02_r_data[18]
port 711 nsew signal input
rlabel metal2 s 414110 119200 414166 120000 6 m02_r_data[19]
port 712 nsew signal input
rlabel metal3 s 0 98608 800 98728 6 m02_r_data[1]
port 713 nsew signal input
rlabel metal2 s 404450 119200 404506 120000 6 m02_r_data[20]
port 714 nsew signal input
rlabel metal2 s 394790 119200 394846 120000 6 m02_r_data[21]
port 715 nsew signal input
rlabel metal2 s 235078 119200 235134 120000 6 m02_r_data[22]
port 716 nsew signal input
rlabel metal2 s 260194 119200 260250 120000 6 m02_r_data[23]
port 717 nsew signal input
rlabel metal3 s 479200 28568 480000 28688 6 m02_r_data[24]
port 718 nsew signal input
rlabel metal2 s 111430 119200 111486 120000 6 m02_r_data[25]
port 719 nsew signal input
rlabel metal2 s 61198 0 61254 800 6 m02_r_data[26]
port 720 nsew signal input
rlabel metal2 s 58622 119200 58678 120000 6 m02_r_data[27]
port 721 nsew signal input
rlabel metal2 s 428922 0 428978 800 6 m02_r_data[28]
port 722 nsew signal input
rlabel metal2 s 338762 119200 338818 120000 6 m02_r_data[29]
port 723 nsew signal input
rlabel metal2 s 220266 119200 220322 120000 6 m02_r_data[2]
port 724 nsew signal input
rlabel metal2 s 244738 119200 244794 120000 6 m02_r_data[30]
port 725 nsew signal input
rlabel metal2 s 116582 0 116638 800 6 m02_r_data[31]
port 726 nsew signal input
rlabel metal2 s 370962 0 371018 800 6 m02_r_data[3]
port 727 nsew signal input
rlabel metal3 s 0 103368 800 103488 6 m02_r_data[4]
port 728 nsew signal input
rlabel metal2 s 181626 0 181682 800 6 m02_r_data[5]
port 729 nsew signal input
rlabel metal2 s 333610 0 333666 800 6 m02_r_data[6]
port 730 nsew signal input
rlabel metal2 s 162306 0 162362 800 6 m02_r_data[7]
port 731 nsew signal input
rlabel metal2 s 50894 0 50950 800 6 m02_r_data[8]
port 732 nsew signal input
rlabel metal2 s 249246 0 249302 800 6 m02_r_data[9]
port 733 nsew signal input
rlabel metal2 s 46386 0 46442 800 6 m02_r_id[0]
port 734 nsew signal input
rlabel metal2 s 352930 0 352986 800 6 m02_r_id[10]
port 735 nsew signal input
rlabel metal2 s 275006 0 275062 800 6 m02_r_id[11]
port 736 nsew signal input
rlabel metal2 s 320730 0 320786 800 6 m02_r_id[1]
port 737 nsew signal input
rlabel metal2 s 270498 0 270554 800 6 m02_r_id[2]
port 738 nsew signal input
rlabel metal3 s 0 46248 800 46368 6 m02_r_id[3]
port 739 nsew signal input
rlabel metal2 s 379978 0 380034 800 6 m02_r_id[4]
port 740 nsew signal input
rlabel metal3 s 479200 57128 480000 57248 6 m02_r_id[5]
port 741 nsew signal input
rlabel metal2 s 238942 119200 238998 120000 6 m02_r_id[6]
port 742 nsew signal input
rlabel metal2 s 179694 0 179750 800 6 m02_r_id[7]
port 743 nsew signal input
rlabel metal2 s 108854 119200 108910 120000 6 m02_r_id[8]
port 744 nsew signal input
rlabel metal2 s 51538 0 51594 800 6 m02_r_id[9]
port 745 nsew signal input
rlabel metal2 s 85026 119200 85082 120000 6 m02_r_last
port 746 nsew signal input
rlabel metal3 s 479200 35368 480000 35488 6 m02_r_ready
port 747 nsew signal output
rlabel metal3 s 0 84328 800 84448 6 m02_r_resp[0]
port 748 nsew signal input
rlabel metal2 s 5814 0 5870 800 6 m02_r_resp[1]
port 749 nsew signal input
rlabel metal2 s 30286 0 30342 800 6 m02_r_user[-1]
port 750 nsew signal input
rlabel metal2 s 221554 0 221610 800 6 m02_r_user[0]
port 751 nsew signal input
rlabel metal3 s 0 27208 800 27328 6 m02_r_valid
port 752 nsew signal input
rlabel metal2 s 251822 119200 251878 120000 6 m02_w_data[0]
port 753 nsew signal output
rlabel metal3 s 0 65288 800 65408 6 m02_w_data[10]
port 754 nsew signal output
rlabel metal2 s 182914 0 182970 800 6 m02_w_data[11]
port 755 nsew signal output
rlabel metal2 s 223486 0 223542 800 6 m02_w_data[12]
port 756 nsew signal output
rlabel metal2 s 313002 119200 313058 120000 6 m02_w_data[13]
port 757 nsew signal output
rlabel metal2 s 285954 0 286010 800 6 m02_w_data[14]
port 758 nsew signal output
rlabel metal2 s 291106 0 291162 800 6 m02_w_data[15]
port 759 nsew signal output
rlabel metal2 s 308494 0 308550 800 6 m02_w_data[16]
port 760 nsew signal output
rlabel metal2 s 57334 119200 57390 120000 6 m02_w_data[17]
port 761 nsew signal output
rlabel metal2 s 217690 0 217746 800 6 m02_w_data[18]
port 762 nsew signal output
rlabel metal2 s 59266 0 59322 800 6 m02_w_data[19]
port 763 nsew signal output
rlabel metal2 s 117870 119200 117926 120000 6 m02_w_data[1]
port 764 nsew signal output
rlabel metal2 s 316222 119200 316278 120000 6 m02_w_data[20]
port 765 nsew signal output
rlabel metal2 s 430210 0 430266 800 6 m02_w_data[21]
port 766 nsew signal output
rlabel metal2 s 27066 119200 27122 120000 6 m02_w_data[22]
port 767 nsew signal output
rlabel metal2 s 441158 119200 441214 120000 6 m02_w_data[23]
port 768 nsew signal output
rlabel metal2 s 249890 0 249946 800 6 m02_w_data[24]
port 769 nsew signal output
rlabel metal2 s 139122 0 139178 800 6 m02_w_data[25]
port 770 nsew signal output
rlabel metal3 s 479200 23128 480000 23248 6 m02_w_data[26]
port 771 nsew signal output
rlabel metal2 s 14186 119200 14242 120000 6 m02_w_data[27]
port 772 nsew signal output
rlabel metal2 s 94042 119200 94098 120000 6 m02_w_data[28]
port 773 nsew signal output
rlabel metal3 s 479200 31288 480000 31408 6 m02_w_data[29]
port 774 nsew signal output
rlabel metal2 s 200302 0 200358 800 6 m02_w_data[2]
port 775 nsew signal output
rlabel metal2 s 341982 0 342038 800 6 m02_w_data[30]
port 776 nsew signal output
rlabel metal2 s 458546 0 458602 800 6 m02_w_data[31]
port 777 nsew signal output
rlabel metal2 s 147494 0 147550 800 6 m02_w_data[3]
port 778 nsew signal output
rlabel metal2 s 219622 0 219678 800 6 m02_w_data[4]
port 779 nsew signal output
rlabel metal2 s 74722 0 74778 800 6 m02_w_data[5]
port 780 nsew signal output
rlabel metal2 s 101126 119200 101182 120000 6 m02_w_data[6]
port 781 nsew signal output
rlabel metal2 s 434718 0 434774 800 6 m02_w_data[7]
port 782 nsew signal output
rlabel metal3 s 0 43528 800 43648 6 m02_w_data[8]
port 783 nsew signal output
rlabel metal2 s 342626 0 342682 800 6 m02_w_data[9]
port 784 nsew signal output
rlabel metal3 s 479200 688 480000 808 6 m02_w_last
port 785 nsew signal output
rlabel metal2 s 338762 0 338818 800 6 m02_w_ready
port 786 nsew signal input
rlabel metal2 s 448242 0 448298 800 6 m02_w_strb[0]
port 787 nsew signal output
rlabel metal2 s 68926 119200 68982 120000 6 m02_w_strb[1]
port 788 nsew signal output
rlabel metal2 s 423770 119200 423826 120000 6 m02_w_strb[2]
port 789 nsew signal output
rlabel metal2 s 328458 0 328514 800 6 m02_w_strb[3]
port 790 nsew signal output
rlabel metal2 s 169390 0 169446 800 6 m02_w_user[-1]
port 791 nsew signal output
rlabel metal3 s 479200 107448 480000 107568 6 m02_w_user[0]
port 792 nsew signal output
rlabel metal2 s 222842 119200 222898 120000 6 m02_w_valid
port 793 nsew signal output
rlabel metal2 s 251178 0 251234 800 6 rst_n
port 794 nsew signal input
rlabel metal2 s 5814 119200 5870 120000 6 s00_ar_addr[0]
port 795 nsew signal input
rlabel metal2 s 451462 119200 451518 120000 6 s00_ar_addr[10]
port 796 nsew signal input
rlabel metal2 s 282734 119200 282790 120000 6 s00_ar_addr[11]
port 797 nsew signal input
rlabel metal2 s 250534 119200 250590 120000 6 s00_ar_addr[12]
port 798 nsew signal input
rlabel metal2 s 381266 0 381322 800 6 s00_ar_addr[13]
port 799 nsew signal input
rlabel metal2 s 211250 0 211306 800 6 s00_ar_addr[14]
port 800 nsew signal input
rlabel metal2 s 454038 119200 454094 120000 6 s00_ar_addr[15]
port 801 nsew signal input
rlabel metal3 s 0 37408 800 37528 6 s00_ar_addr[16]
port 802 nsew signal input
rlabel metal2 s 71502 0 71558 800 6 s00_ar_addr[17]
port 803 nsew signal input
rlabel metal2 s 256330 119200 256386 120000 6 s00_ar_addr[18]
port 804 nsew signal input
rlabel metal2 s 446954 119200 447010 120000 6 s00_ar_addr[19]
port 805 nsew signal input
rlabel metal2 s 159730 0 159786 800 6 s00_ar_addr[1]
port 806 nsew signal input
rlabel metal3 s 479200 19728 480000 19848 6 s00_ar_addr[20]
port 807 nsew signal input
rlabel metal2 s 149426 119200 149482 120000 6 s00_ar_addr[21]
port 808 nsew signal input
rlabel metal2 s 13542 0 13598 800 6 s00_ar_addr[22]
port 809 nsew signal input
rlabel metal2 s 419262 0 419318 800 6 s00_ar_addr[23]
port 810 nsew signal input
rlabel metal3 s 479200 42848 480000 42968 6 s00_ar_addr[24]
port 811 nsew signal input
rlabel metal2 s 266634 119200 266690 120000 6 s00_ar_addr[25]
port 812 nsew signal input
rlabel metal2 s 196438 0 196494 800 6 s00_ar_addr[26]
port 813 nsew signal input
rlabel metal2 s 405094 0 405150 800 6 s00_ar_addr[27]
port 814 nsew signal input
rlabel metal2 s 43810 0 43866 800 6 s00_ar_addr[28]
port 815 nsew signal input
rlabel metal2 s 208030 0 208086 800 6 s00_ar_addr[29]
port 816 nsew signal input
rlabel metal2 s 424414 0 424470 800 6 s00_ar_addr[2]
port 817 nsew signal input
rlabel metal2 s 103058 119200 103114 120000 6 s00_ar_addr[30]
port 818 nsew signal input
rlabel metal2 s 57978 0 58034 800 6 s00_ar_addr[31]
port 819 nsew signal input
rlabel metal3 s 0 16328 800 16448 6 s00_ar_addr[3]
port 820 nsew signal input
rlabel metal2 s 10322 0 10378 800 6 s00_ar_addr[4]
port 821 nsew signal input
rlabel metal2 s 235722 0 235778 800 6 s00_ar_addr[5]
port 822 nsew signal input
rlabel metal2 s 393502 119200 393558 120000 6 s00_ar_addr[6]
port 823 nsew signal input
rlabel metal2 s 133326 0 133382 800 6 s00_ar_addr[7]
port 824 nsew signal input
rlabel metal2 s 43166 0 43222 800 6 s00_ar_addr[8]
port 825 nsew signal input
rlabel metal2 s 132038 119200 132094 120000 6 s00_ar_addr[9]
port 826 nsew signal input
rlabel metal2 s 69570 119200 69626 120000 6 s00_ar_burst[0]
port 827 nsew signal input
rlabel metal2 s 129462 0 129518 800 6 s00_ar_burst[1]
port 828 nsew signal input
rlabel metal3 s 479200 94528 480000 94648 6 s00_ar_cache[0]
port 829 nsew signal input
rlabel metal2 s 240874 119200 240930 120000 6 s00_ar_cache[1]
port 830 nsew signal input
rlabel metal2 s 467562 119200 467618 120000 6 s00_ar_cache[2]
port 831 nsew signal input
rlabel metal2 s 86314 119200 86370 120000 6 s00_ar_cache[3]
port 832 nsew signal input
rlabel metal2 s 362590 119200 362646 120000 6 s00_ar_id[0]
port 833 nsew signal input
rlabel metal2 s 396722 0 396778 800 6 s00_ar_id[1]
port 834 nsew signal input
rlabel metal2 s 476578 119200 476634 120000 6 s00_ar_id[2]
port 835 nsew signal input
rlabel metal3 s 479200 43528 480000 43648 6 s00_ar_id[3]
port 836 nsew signal input
rlabel metal2 s 346490 0 346546 800 6 s00_ar_id[4]
port 837 nsew signal input
rlabel metal3 s 479200 37408 480000 37528 6 s00_ar_id[5]
port 838 nsew signal input
rlabel metal2 s 103702 119200 103758 120000 6 s00_ar_id[6]
port 839 nsew signal input
rlabel metal2 s 81162 0 81218 800 6 s00_ar_id[7]
port 840 nsew signal input
rlabel metal2 s 417330 119200 417386 120000 6 s00_ar_id[8]
port 841 nsew signal input
rlabel metal2 s 366454 0 366510 800 6 s00_ar_id[9]
port 842 nsew signal input
rlabel metal2 s 182270 119200 182326 120000 6 s00_ar_len[0]
port 843 nsew signal input
rlabel metal2 s 434074 0 434130 800 6 s00_ar_len[1]
port 844 nsew signal input
rlabel metal2 s 369030 0 369086 800 6 s00_ar_len[2]
port 845 nsew signal input
rlabel metal2 s 30930 119200 30986 120000 6 s00_ar_len[3]
port 846 nsew signal input
rlabel metal2 s 468850 119200 468906 120000 6 s00_ar_len[4]
port 847 nsew signal input
rlabel metal2 s 232502 119200 232558 120000 6 s00_ar_len[5]
port 848 nsew signal input
rlabel metal2 s 377402 0 377458 800 6 s00_ar_len[6]
port 849 nsew signal input
rlabel metal2 s 420550 119200 420606 120000 6 s00_ar_len[7]
port 850 nsew signal input
rlabel metal3 s 0 110168 800 110288 6 s00_ar_lock
port 851 nsew signal input
rlabel metal2 s 336186 119200 336242 120000 6 s00_ar_prot[0]
port 852 nsew signal input
rlabel metal2 s 416042 0 416098 800 6 s00_ar_prot[1]
port 853 nsew signal input
rlabel metal2 s 417974 119200 418030 120000 6 s00_ar_prot[2]
port 854 nsew signal input
rlabel metal2 s 45098 0 45154 800 6 s00_ar_qos[0]
port 855 nsew signal input
rlabel metal2 s 400586 0 400642 800 6 s00_ar_qos[1]
port 856 nsew signal input
rlabel metal2 s 105634 0 105690 800 6 s00_ar_qos[2]
port 857 nsew signal input
rlabel metal2 s 142986 119200 143042 120000 6 s00_ar_qos[3]
port 858 nsew signal input
rlabel metal2 s 429566 0 429622 800 6 s00_ar_ready
port 859 nsew signal output
rlabel metal2 s 351642 0 351698 800 6 s00_ar_region[0]
port 860 nsew signal input
rlabel metal3 s 479200 84328 480000 84448 6 s00_ar_region[1]
port 861 nsew signal input
rlabel metal2 s 327814 0 327870 800 6 s00_ar_region[2]
port 862 nsew signal input
rlabel metal2 s 403806 119200 403862 120000 6 s00_ar_region[3]
port 863 nsew signal input
rlabel metal2 s 461766 119200 461822 120000 6 s00_ar_size[0]
port 864 nsew signal input
rlabel metal2 s 410890 0 410946 800 6 s00_ar_size[1]
port 865 nsew signal input
rlabel metal2 s 9678 0 9734 800 6 s00_ar_size[2]
port 866 nsew signal input
rlabel metal2 s 178406 119200 178462 120000 6 s00_ar_user[-1]
port 867 nsew signal input
rlabel metal2 s 171322 0 171378 800 6 s00_ar_user[0]
port 868 nsew signal input
rlabel metal2 s 29642 0 29698 800 6 s00_ar_valid
port 869 nsew signal input
rlabel metal3 s 479200 111528 480000 111648 6 s00_aw_addr[0]
port 870 nsew signal input
rlabel metal2 s 237654 119200 237710 120000 6 s00_aw_addr[10]
port 871 nsew signal input
rlabel metal2 s 148782 119200 148838 120000 6 s00_aw_addr[11]
port 872 nsew signal input
rlabel metal2 s 286598 119200 286654 120000 6 s00_aw_addr[12]
port 873 nsew signal input
rlabel metal2 s 38658 119200 38714 120000 6 s00_aw_addr[13]
port 874 nsew signal input
rlabel metal2 s 264702 0 264758 800 6 s00_aw_addr[14]
port 875 nsew signal input
rlabel metal2 s 432786 0 432842 800 6 s00_aw_addr[15]
port 876 nsew signal input
rlabel metal2 s 56690 119200 56746 120000 6 s00_aw_addr[16]
port 877 nsew signal input
rlabel metal2 s 309138 0 309194 800 6 s00_aw_addr[17]
port 878 nsew signal input
rlabel metal2 s 115294 0 115350 800 6 s00_aw_addr[18]
port 879 nsew signal input
rlabel metal2 s 231214 0 231270 800 6 s00_aw_addr[19]
port 880 nsew signal input
rlabel metal2 s 92110 119200 92166 120000 6 s00_aw_addr[1]
port 881 nsew signal input
rlabel metal3 s 0 10888 800 11008 6 s00_aw_addr[20]
port 882 nsew signal input
rlabel metal2 s 329746 0 329802 800 6 s00_aw_addr[21]
port 883 nsew signal input
rlabel metal3 s 479200 34008 480000 34128 6 s00_aw_addr[22]
port 884 nsew signal input
rlabel metal2 s 374182 119200 374238 120000 6 s00_aw_addr[23]
port 885 nsew signal input
rlabel metal2 s 10966 0 11022 800 6 s00_aw_addr[24]
port 886 nsew signal input
rlabel metal2 s 319442 0 319498 800 6 s00_aw_addr[25]
port 887 nsew signal input
rlabel metal2 s 86958 119200 87014 120000 6 s00_aw_addr[26]
port 888 nsew signal input
rlabel metal2 s 156510 119200 156566 120000 6 s00_aw_addr[27]
port 889 nsew signal input
rlabel metal2 s 412178 119200 412234 120000 6 s00_aw_addr[28]
port 890 nsew signal input
rlabel metal2 s 201590 119200 201646 120000 6 s00_aw_addr[29]
port 891 nsew signal input
rlabel metal2 s 210606 0 210662 800 6 s00_aw_addr[2]
port 892 nsew signal input
rlabel metal2 s 329102 119200 329158 120000 6 s00_aw_addr[30]
port 893 nsew signal input
rlabel metal2 s 63774 0 63830 800 6 s00_aw_addr[31]
port 894 nsew signal input
rlabel metal2 s 112074 119200 112130 120000 6 s00_aw_addr[3]
port 895 nsew signal input
rlabel metal2 s 341338 119200 341394 120000 6 s00_aw_addr[4]
port 896 nsew signal input
rlabel metal2 s 224130 119200 224186 120000 6 s00_aw_addr[5]
port 897 nsew signal input
rlabel metal2 s 233146 0 233202 800 6 s00_aw_addr[6]
port 898 nsew signal input
rlabel metal2 s 9034 0 9090 800 6 s00_aw_addr[7]
port 899 nsew signal input
rlabel metal2 s 81806 0 81862 800 6 s00_aw_addr[8]
port 900 nsew signal input
rlabel metal3 s 479200 40128 480000 40248 6 s00_aw_addr[9]
port 901 nsew signal input
rlabel metal2 s 108210 0 108266 800 6 s00_aw_burst[0]
port 902 nsew signal input
rlabel metal2 s 244094 0 244150 800 6 s00_aw_burst[1]
port 903 nsew signal input
rlabel metal2 s 153290 119200 153346 120000 6 s00_aw_cache[0]
port 904 nsew signal input
rlabel metal2 s 170034 0 170090 800 6 s00_aw_cache[1]
port 905 nsew signal input
rlabel metal2 s 32218 0 32274 800 6 s00_aw_cache[2]
port 906 nsew signal input
rlabel metal2 s 367098 119200 367154 120000 6 s00_aw_cache[3]
port 907 nsew signal input
rlabel metal2 s 120446 119200 120502 120000 6 s00_aw_id[0]
port 908 nsew signal input
rlabel metal2 s 422482 0 422538 800 6 s00_aw_id[1]
port 909 nsew signal input
rlabel metal2 s 300766 0 300822 800 6 s00_aw_id[2]
port 910 nsew signal input
rlabel metal2 s 383842 0 383898 800 6 s00_aw_id[3]
port 911 nsew signal input
rlabel metal2 s 455326 0 455382 800 6 s00_aw_id[4]
port 912 nsew signal input
rlabel metal3 s 479200 32648 480000 32768 6 s00_aw_id[5]
port 913 nsew signal input
rlabel metal2 s 358726 0 358782 800 6 s00_aw_id[6]
port 914 nsew signal input
rlabel metal2 s 9678 119200 9734 120000 6 s00_aw_id[7]
port 915 nsew signal input
rlabel metal2 s 130750 119200 130806 120000 6 s00_aw_id[8]
port 916 nsew signal input
rlabel metal3 s 0 68688 800 68808 6 s00_aw_id[9]
port 917 nsew signal input
rlabel metal2 s 117226 119200 117282 120000 6 s00_aw_len[0]
port 918 nsew signal input
rlabel metal2 s 460478 0 460534 800 6 s00_aw_len[1]
port 919 nsew signal input
rlabel metal2 s 127530 0 127586 800 6 s00_aw_len[2]
port 920 nsew signal input
rlabel metal2 s 70214 119200 70270 120000 6 s00_aw_len[3]
port 921 nsew signal input
rlabel metal3 s 0 17008 800 17128 6 s00_aw_len[4]
port 922 nsew signal input
rlabel metal2 s 384486 0 384542 800 6 s00_aw_len[5]
port 923 nsew signal input
rlabel metal2 s 180982 119200 181038 120000 6 s00_aw_len[6]
port 924 nsew signal input
rlabel metal2 s 175186 0 175242 800 6 s00_aw_len[7]
port 925 nsew signal input
rlabel metal2 s 43810 119200 43866 120000 6 s00_aw_lock
port 926 nsew signal input
rlabel metal2 s 285310 119200 285366 120000 6 s00_aw_prot[0]
port 927 nsew signal input
rlabel metal2 s 428922 119200 428978 120000 6 s00_aw_prot[1]
port 928 nsew signal input
rlabel metal2 s 121090 0 121146 800 6 s00_aw_prot[2]
port 929 nsew signal input
rlabel metal2 s 40590 0 40646 800 6 s00_aw_qos[0]
port 930 nsew signal input
rlabel metal2 s 288530 0 288586 800 6 s00_aw_qos[1]
port 931 nsew signal input
rlabel metal2 s 282090 119200 282146 120000 6 s00_aw_qos[2]
port 932 nsew signal input
rlabel metal3 s 479200 13608 480000 13728 6 s00_aw_qos[3]
port 933 nsew signal input
rlabel metal2 s 303986 0 304042 800 6 s00_aw_ready
port 934 nsew signal output
rlabel metal3 s 479200 119688 480000 119808 6 s00_aw_region[0]
port 935 nsew signal input
rlabel metal2 s 56690 0 56746 800 6 s00_aw_region[1]
port 936 nsew signal input
rlabel metal2 s 388350 119200 388406 120000 6 s00_aw_region[2]
port 937 nsew signal input
rlabel metal2 s 130750 0 130806 800 6 s00_aw_region[3]
port 938 nsew signal input
rlabel metal3 s 0 59168 800 59288 6 s00_aw_size[0]
port 939 nsew signal input
rlabel metal2 s 178406 0 178462 800 6 s00_aw_size[1]
port 940 nsew signal input
rlabel metal2 s 264702 119200 264758 120000 6 s00_aw_size[2]
port 941 nsew signal input
rlabel metal2 s 197082 119200 197138 120000 6 s00_aw_user[-1]
port 942 nsew signal input
rlabel metal2 s 217046 119200 217102 120000 6 s00_aw_user[0]
port 943 nsew signal input
rlabel metal2 s 182914 119200 182970 120000 6 s00_aw_valid
port 944 nsew signal input
rlabel metal3 s 0 50328 800 50448 6 s00_b_id[0]
port 945 nsew signal output
rlabel metal2 s 286598 0 286654 800 6 s00_b_id[1]
port 946 nsew signal output
rlabel metal3 s 479200 97248 480000 97368 6 s00_b_id[2]
port 947 nsew signal output
rlabel metal2 s 329746 119200 329802 120000 6 s00_b_id[3]
port 948 nsew signal output
rlabel metal2 s 245382 119200 245438 120000 6 s00_b_id[4]
port 949 nsew signal output
rlabel metal3 s 479200 36728 480000 36848 6 s00_b_id[5]
port 950 nsew signal output
rlabel metal2 s 372894 0 372950 800 6 s00_b_id[6]
port 951 nsew signal output
rlabel metal2 s 373538 119200 373594 120000 6 s00_b_id[7]
port 952 nsew signal output
rlabel metal3 s 0 13608 800 13728 6 s00_b_id[8]
port 953 nsew signal output
rlabel metal2 s 95330 0 95386 800 6 s00_b_id[9]
port 954 nsew signal output
rlabel metal2 s 121734 119200 121790 120000 6 s00_b_ready
port 955 nsew signal input
rlabel metal2 s 99838 0 99894 800 6 s00_b_resp[0]
port 956 nsew signal output
rlabel metal2 s 463698 0 463754 800 6 s00_b_resp[1]
port 957 nsew signal output
rlabel metal2 s 197726 119200 197782 120000 6 s00_b_user[-1]
port 958 nsew signal output
rlabel metal2 s 393502 0 393558 800 6 s00_b_user[0]
port 959 nsew signal output
rlabel metal3 s 0 102688 800 102808 6 s00_b_valid
port 960 nsew signal output
rlabel metal2 s 387706 0 387762 800 6 s00_r_data[0]
port 961 nsew signal output
rlabel metal2 s 141054 0 141110 800 6 s00_r_data[10]
port 962 nsew signal output
rlabel metal2 s 36726 0 36782 800 6 s00_r_data[11]
port 963 nsew signal output
rlabel metal2 s 457902 119200 457958 120000 6 s00_r_data[12]
port 964 nsew signal output
rlabel metal2 s 302698 119200 302754 120000 6 s00_r_data[13]
port 965 nsew signal output
rlabel metal2 s 334898 0 334954 800 6 s00_r_data[14]
port 966 nsew signal output
rlabel metal3 s 0 112208 800 112328 6 s00_r_data[15]
port 967 nsew signal output
rlabel metal3 s 0 41488 800 41608 6 s00_r_data[16]
port 968 nsew signal output
rlabel metal2 s 158442 0 158498 800 6 s00_r_data[17]
port 969 nsew signal output
rlabel metal2 s 285954 119200 286010 120000 6 s00_r_data[18]
port 970 nsew signal output
rlabel metal3 s 479200 92488 480000 92608 6 s00_r_data[19]
port 971 nsew signal output
rlabel metal2 s 256974 119200 257030 120000 6 s00_r_data[1]
port 972 nsew signal output
rlabel metal2 s 304630 119200 304686 120000 6 s00_r_data[20]
port 973 nsew signal output
rlabel metal2 s 241518 0 241574 800 6 s00_r_data[21]
port 974 nsew signal output
rlabel metal2 s 93398 0 93454 800 6 s00_r_data[22]
port 975 nsew signal output
rlabel metal2 s 398010 0 398066 800 6 s00_r_data[23]
port 976 nsew signal output
rlabel metal2 s 30286 119200 30342 120000 6 s00_r_data[24]
port 977 nsew signal output
rlabel metal2 s 126886 119200 126942 120000 6 s00_r_data[25]
port 978 nsew signal output
rlabel metal2 s 462410 119200 462466 120000 6 s00_r_data[26]
port 979 nsew signal output
rlabel metal2 s 28354 0 28410 800 6 s00_r_data[27]
port 980 nsew signal output
rlabel metal2 s 27066 0 27122 800 6 s00_r_data[28]
port 981 nsew signal output
rlabel metal2 s 186134 0 186190 800 6 s00_r_data[29]
port 982 nsew signal output
rlabel metal2 s 21914 0 21970 800 6 s00_r_data[2]
port 983 nsew signal output
rlabel metal2 s 430854 119200 430910 120000 6 s00_r_data[30]
port 984 nsew signal output
rlabel metal2 s 441802 0 441858 800 6 s00_r_data[31]
port 985 nsew signal output
rlabel metal2 s 298834 119200 298890 120000 6 s00_r_data[3]
port 986 nsew signal output
rlabel metal2 s 92754 119200 92810 120000 6 s00_r_data[4]
port 987 nsew signal output
rlabel metal2 s 336830 119200 336886 120000 6 s00_r_data[5]
port 988 nsew signal output
rlabel metal2 s 407670 0 407726 800 6 s00_r_data[6]
port 989 nsew signal output
rlabel metal2 s 115938 0 115994 800 6 s00_r_data[7]
port 990 nsew signal output
rlabel metal2 s 126242 119200 126298 120000 6 s00_r_data[8]
port 991 nsew signal output
rlabel metal2 s 203522 119200 203578 120000 6 s00_r_data[9]
port 992 nsew signal output
rlabel metal3 s 0 29928 800 30048 6 s00_r_id[0]
port 993 nsew signal output
rlabel metal2 s 118514 119200 118570 120000 6 s00_r_id[1]
port 994 nsew signal output
rlabel metal3 s 0 57808 800 57928 6 s00_r_id[2]
port 995 nsew signal output
rlabel metal2 s 114006 119200 114062 120000 6 s00_r_id[3]
port 996 nsew signal output
rlabel metal2 s 70214 0 70270 800 6 s00_r_id[4]
port 997 nsew signal output
rlabel metal3 s 0 70048 800 70168 6 s00_r_id[5]
port 998 nsew signal output
rlabel metal2 s 284666 0 284722 800 6 s00_r_id[6]
port 999 nsew signal output
rlabel metal2 s 19982 0 20038 800 6 s00_r_id[7]
port 1000 nsew signal output
rlabel metal2 s 256974 0 257030 800 6 s00_r_id[8]
port 1001 nsew signal output
rlabel metal2 s 399298 119200 399354 120000 6 s00_r_id[9]
port 1002 nsew signal output
rlabel metal3 s 0 45568 800 45688 6 s00_r_last
port 1003 nsew signal output
rlabel metal2 s 142342 119200 142398 120000 6 s00_r_ready
port 1004 nsew signal input
rlabel metal3 s 0 31968 800 32088 6 s00_r_resp[0]
port 1005 nsew signal output
rlabel metal2 s 303342 0 303398 800 6 s00_r_resp[1]
port 1006 nsew signal output
rlabel metal3 s 479200 59168 480000 59288 6 s00_r_user[-1]
port 1007 nsew signal output
rlabel metal2 s 53470 0 53526 800 6 s00_r_user[0]
port 1008 nsew signal output
rlabel metal3 s 0 73448 800 73568 6 s00_r_valid
port 1009 nsew signal output
rlabel metal2 s 148782 0 148838 800 6 s00_w_data[0]
port 1010 nsew signal input
rlabel metal2 s 460478 119200 460534 120000 6 s00_w_data[10]
port 1011 nsew signal input
rlabel metal2 s 102414 119200 102470 120000 6 s00_w_data[11]
port 1012 nsew signal input
rlabel metal2 s 230570 119200 230626 120000 6 s00_w_data[12]
port 1013 nsew signal input
rlabel metal3 s 0 108128 800 108248 6 s00_w_data[13]
port 1014 nsew signal input
rlabel metal2 s 394146 0 394202 800 6 s00_w_data[14]
port 1015 nsew signal input
rlabel metal2 s 61842 0 61898 800 6 s00_w_data[15]
port 1016 nsew signal input
rlabel metal3 s 0 6128 800 6248 6 s00_w_data[16]
port 1017 nsew signal input
rlabel metal2 s 472714 0 472770 800 6 s00_w_data[17]
port 1018 nsew signal input
rlabel metal2 s 161018 119200 161074 120000 6 s00_w_data[18]
port 1019 nsew signal input
rlabel metal2 s 198370 0 198426 800 6 s00_w_data[19]
port 1020 nsew signal input
rlabel metal2 s 296902 119200 296958 120000 6 s00_w_data[1]
port 1021 nsew signal input
rlabel metal2 s 68282 119200 68338 120000 6 s00_w_data[20]
port 1022 nsew signal input
rlabel metal3 s 0 91128 800 91248 6 s00_w_data[21]
port 1023 nsew signal input
rlabel metal2 s 122378 119200 122434 120000 6 s00_w_data[22]
port 1024 nsew signal input
rlabel metal2 s 227994 0 228050 800 6 s00_w_data[23]
port 1025 nsew signal input
rlabel metal2 s 430854 0 430910 800 6 s00_w_data[24]
port 1026 nsew signal input
rlabel metal2 s 280158 0 280214 800 6 s00_w_data[25]
port 1027 nsew signal input
rlabel metal3 s 0 86368 800 86488 6 s00_w_data[26]
port 1028 nsew signal input
rlabel metal3 s 479200 72088 480000 72208 6 s00_w_data[27]
port 1029 nsew signal input
rlabel metal2 s 60554 119200 60610 120000 6 s00_w_data[28]
port 1030 nsew signal input
rlabel metal3 s 479200 69368 480000 69488 6 s00_w_data[29]
port 1031 nsew signal input
rlabel metal2 s 408958 119200 409014 120000 6 s00_w_data[2]
port 1032 nsew signal input
rlabel metal3 s 479200 106768 480000 106888 6 s00_w_data[30]
port 1033 nsew signal input
rlabel metal2 s 253110 0 253166 800 6 s00_w_data[31]
port 1034 nsew signal input
rlabel metal2 s 265346 119200 265402 120000 6 s00_w_data[3]
port 1035 nsew signal input
rlabel metal3 s 0 76848 800 76968 6 s00_w_data[4]
port 1036 nsew signal input
rlabel metal2 s 408314 0 408370 800 6 s00_w_data[5]
port 1037 nsew signal input
rlabel metal2 s 199658 0 199714 800 6 s00_w_data[6]
port 1038 nsew signal input
rlabel metal3 s 0 59848 800 59968 6 s00_w_data[7]
port 1039 nsew signal input
rlabel metal2 s 282734 0 282790 800 6 s00_w_data[8]
port 1040 nsew signal input
rlabel metal2 s 662 119200 718 120000 6 s00_w_data[9]
port 1041 nsew signal input
rlabel metal3 s 479200 53728 480000 53848 6 s00_w_last
port 1042 nsew signal input
rlabel metal3 s 479200 7488 480000 7608 6 s00_w_ready
port 1043 nsew signal output
rlabel metal2 s 165526 0 165582 800 6 s00_w_strb[0]
port 1044 nsew signal input
rlabel metal2 s 124310 119200 124366 120000 6 s00_w_strb[1]
port 1045 nsew signal input
rlabel metal2 s 55402 0 55458 800 6 s00_w_strb[2]
port 1046 nsew signal input
rlabel metal2 s 452750 0 452806 800 6 s00_w_strb[3]
port 1047 nsew signal input
rlabel metal2 s 333610 119200 333666 120000 6 s00_w_user[-1]
port 1048 nsew signal input
rlabel metal3 s 479200 78888 480000 79008 6 s00_w_user[0]
port 1049 nsew signal input
rlabel metal2 s 400586 119200 400642 120000 6 s00_w_valid
port 1050 nsew signal input
rlabel metal2 s 327170 119200 327226 120000 6 s01_ar_addr[0]
port 1051 nsew signal input
rlabel metal2 s 315578 0 315634 800 6 s01_ar_addr[10]
port 1052 nsew signal input
rlabel metal2 s 445666 0 445722 800 6 s01_ar_addr[11]
port 1053 nsew signal input
rlabel metal2 s 297546 0 297602 800 6 s01_ar_addr[12]
port 1054 nsew signal input
rlabel metal2 s 135258 0 135314 800 6 s01_ar_addr[13]
port 1055 nsew signal input
rlabel metal3 s 0 101328 800 101448 6 s01_ar_addr[14]
port 1056 nsew signal input
rlabel metal2 s 253754 0 253810 800 6 s01_ar_addr[15]
port 1057 nsew signal input
rlabel metal2 s 215758 0 215814 800 6 s01_ar_addr[16]
port 1058 nsew signal input
rlabel metal2 s 388994 119200 389050 120000 6 s01_ar_addr[17]
port 1059 nsew signal input
rlabel metal2 s 215758 119200 215814 120000 6 s01_ar_addr[18]
port 1060 nsew signal input
rlabel metal2 s 309782 0 309838 800 6 s01_ar_addr[19]
port 1061 nsew signal input
rlabel metal2 s 28998 119200 29054 120000 6 s01_ar_addr[1]
port 1062 nsew signal input
rlabel metal2 s 237010 0 237066 800 6 s01_ar_addr[20]
port 1063 nsew signal input
rlabel metal2 s 60554 0 60610 800 6 s01_ar_addr[21]
port 1064 nsew signal input
rlabel metal2 s 189354 119200 189410 120000 6 s01_ar_addr[22]
port 1065 nsew signal input
rlabel metal2 s 279514 119200 279570 120000 6 s01_ar_addr[23]
port 1066 nsew signal input
rlabel metal2 s 292394 119200 292450 120000 6 s01_ar_addr[24]
port 1067 nsew signal input
rlabel metal2 s 464342 0 464398 800 6 s01_ar_addr[25]
port 1068 nsew signal input
rlabel metal2 s 189998 119200 190054 120000 6 s01_ar_addr[26]
port 1069 nsew signal input
rlabel metal2 s 449530 0 449586 800 6 s01_ar_addr[27]
port 1070 nsew signal input
rlabel metal3 s 0 74128 800 74248 6 s01_ar_addr[28]
port 1071 nsew signal input
rlabel metal2 s 269210 0 269266 800 6 s01_ar_addr[29]
port 1072 nsew signal input
rlabel metal2 s 316866 119200 316922 120000 6 s01_ar_addr[2]
port 1073 nsew signal input
rlabel metal2 s 296258 119200 296314 120000 6 s01_ar_addr[30]
port 1074 nsew signal input
rlabel metal2 s 11610 0 11666 800 6 s01_ar_addr[31]
port 1075 nsew signal input
rlabel metal3 s 0 69368 800 69488 6 s01_ar_addr[3]
port 1076 nsew signal input
rlabel metal2 s 181626 119200 181682 120000 6 s01_ar_addr[4]
port 1077 nsew signal input
rlabel metal2 s 350354 119200 350410 120000 6 s01_ar_addr[5]
port 1078 nsew signal input
rlabel metal2 s 233146 119200 233202 120000 6 s01_ar_addr[6]
port 1079 nsew signal input
rlabel metal2 s 127530 119200 127586 120000 6 s01_ar_addr[7]
port 1080 nsew signal input
rlabel metal2 s 290462 119200 290518 120000 6 s01_ar_addr[8]
port 1081 nsew signal input
rlabel metal2 s 385774 0 385830 800 6 s01_ar_addr[9]
port 1082 nsew signal input
rlabel metal2 s 300122 119200 300178 120000 6 s01_ar_burst[0]
port 1083 nsew signal input
rlabel metal2 s 254398 119200 254454 120000 6 s01_ar_burst[1]
port 1084 nsew signal input
rlabel metal2 s 145562 0 145618 800 6 s01_ar_cache[0]
port 1085 nsew signal input
rlabel metal2 s 35438 0 35494 800 6 s01_ar_cache[1]
port 1086 nsew signal input
rlabel metal3 s 479200 55088 480000 55208 6 s01_ar_cache[2]
port 1087 nsew signal input
rlabel metal2 s 8390 119200 8446 120000 6 s01_ar_cache[3]
port 1088 nsew signal input
rlabel metal2 s 19338 0 19394 800 6 s01_ar_id[0]
port 1089 nsew signal input
rlabel metal2 s 473358 0 473414 800 6 s01_ar_id[1]
port 1090 nsew signal input
rlabel metal2 s 232502 0 232558 800 6 s01_ar_id[2]
port 1091 nsew signal input
rlabel metal2 s 414110 0 414166 800 6 s01_ar_id[3]
port 1092 nsew signal input
rlabel metal2 s 207386 119200 207442 120000 6 s01_ar_id[4]
port 1093 nsew signal input
rlabel metal2 s 190642 0 190698 800 6 s01_ar_id[5]
port 1094 nsew signal input
rlabel metal2 s 161662 0 161718 800 6 s01_ar_id[6]
port 1095 nsew signal input
rlabel metal2 s 354218 119200 354274 120000 6 s01_ar_id[7]
port 1096 nsew signal input
rlabel metal2 s 410246 0 410302 800 6 s01_ar_id[8]
port 1097 nsew signal input
rlabel metal3 s 479200 81608 480000 81728 6 s01_ar_id[9]
port 1098 nsew signal input
rlabel metal3 s 479200 1368 480000 1488 6 s01_ar_len[0]
port 1099 nsew signal input
rlabel metal3 s 479200 61888 480000 62008 6 s01_ar_len[1]
port 1100 nsew signal input
rlabel metal2 s 65062 119200 65118 120000 6 s01_ar_len[2]
port 1101 nsew signal input
rlabel metal2 s 292394 0 292450 800 6 s01_ar_len[3]
port 1102 nsew signal input
rlabel metal2 s 408314 119200 408370 120000 6 s01_ar_len[4]
port 1103 nsew signal input
rlabel metal2 s 363878 0 363934 800 6 s01_ar_len[5]
port 1104 nsew signal input
rlabel metal3 s 479200 52368 480000 52488 6 s01_ar_len[6]
port 1105 nsew signal input
rlabel metal2 s 312358 119200 312414 120000 6 s01_ar_len[7]
port 1106 nsew signal input
rlabel metal2 s 323950 119200 324006 120000 6 s01_ar_lock
port 1107 nsew signal input
rlabel metal2 s 409602 0 409658 800 6 s01_ar_prot[0]
port 1108 nsew signal input
rlabel metal2 s 330390 0 330446 800 6 s01_ar_prot[1]
port 1109 nsew signal input
rlabel metal2 s 248602 119200 248658 120000 6 s01_ar_prot[2]
port 1110 nsew signal input
rlabel metal2 s 200302 119200 200358 120000 6 s01_ar_qos[0]
port 1111 nsew signal input
rlabel metal3 s 479200 18368 480000 18488 6 s01_ar_qos[1]
port 1112 nsew signal input
rlabel metal2 s 206098 0 206154 800 6 s01_ar_qos[2]
port 1113 nsew signal input
rlabel metal3 s 0 23128 800 23248 6 s01_ar_qos[3]
port 1114 nsew signal input
rlabel metal2 s 224130 0 224186 800 6 s01_ar_ready
port 1115 nsew signal output
rlabel metal3 s 479200 62568 480000 62688 6 s01_ar_region[0]
port 1116 nsew signal input
rlabel metal2 s 160374 119200 160430 120000 6 s01_ar_region[1]
port 1117 nsew signal input
rlabel metal2 s 431498 0 431554 800 6 s01_ar_region[2]
port 1118 nsew signal input
rlabel metal2 s 3882 119200 3938 120000 6 s01_ar_region[3]
port 1119 nsew signal input
rlabel metal2 s 461122 0 461178 800 6 s01_ar_size[0]
port 1120 nsew signal input
rlabel metal2 s 110142 119200 110198 120000 6 s01_ar_size[1]
port 1121 nsew signal input
rlabel metal2 s 262126 0 262182 800 6 s01_ar_size[2]
port 1122 nsew signal input
rlabel metal3 s 479200 85008 480000 85128 6 s01_ar_user[-1]
port 1123 nsew signal input
rlabel metal2 s 458546 119200 458602 120000 6 s01_ar_user[0]
port 1124 nsew signal input
rlabel metal2 s 348422 119200 348478 120000 6 s01_ar_valid
port 1125 nsew signal input
rlabel metal2 s 437938 119200 437994 120000 6 s01_aw_addr[0]
port 1126 nsew signal input
rlabel metal3 s 479200 80248 480000 80368 6 s01_aw_addr[10]
port 1127 nsew signal input
rlabel metal2 s 313646 0 313702 800 6 s01_aw_addr[11]
port 1128 nsew signal input
rlabel metal2 s 434074 119200 434130 120000 6 s01_aw_addr[12]
port 1129 nsew signal input
rlabel metal2 s 153290 0 153346 800 6 s01_aw_addr[13]
port 1130 nsew signal input
rlabel metal2 s 279514 0 279570 800 6 s01_aw_addr[14]
port 1131 nsew signal input
rlabel metal2 s 425058 0 425114 800 6 s01_aw_addr[15]
port 1132 nsew signal input
rlabel metal3 s 0 72088 800 72208 6 s01_aw_addr[16]
port 1133 nsew signal input
rlabel metal2 s 39302 119200 39358 120000 6 s01_aw_addr[17]
port 1134 nsew signal input
rlabel metal2 s 459834 119200 459890 120000 6 s01_aw_addr[18]
port 1135 nsew signal input
rlabel metal2 s 151358 0 151414 800 6 s01_aw_addr[19]
port 1136 nsew signal input
rlabel metal2 s 192574 0 192630 800 6 s01_aw_addr[1]
port 1137 nsew signal input
rlabel metal2 s 214470 119200 214526 120000 6 s01_aw_addr[20]
port 1138 nsew signal input
rlabel metal2 s 123022 119200 123078 120000 6 s01_aw_addr[21]
port 1139 nsew signal input
rlabel metal2 s 388350 0 388406 800 6 s01_aw_addr[22]
port 1140 nsew signal input
rlabel metal2 s 474646 119200 474702 120000 6 s01_aw_addr[23]
port 1141 nsew signal input
rlabel metal2 s 47674 119200 47730 120000 6 s01_aw_addr[24]
port 1142 nsew signal input
rlabel metal2 s 476578 0 476634 800 6 s01_aw_addr[25]
port 1143 nsew signal input
rlabel metal2 s 88246 119200 88302 120000 6 s01_aw_addr[26]
port 1144 nsew signal input
rlabel metal2 s 139766 0 139822 800 6 s01_aw_addr[27]
port 1145 nsew signal input
rlabel metal2 s 246670 0 246726 800 6 s01_aw_addr[28]
port 1146 nsew signal input
rlabel metal2 s 3238 0 3294 800 6 s01_aw_addr[29]
port 1147 nsew signal input
rlabel metal2 s 224774 119200 224830 120000 6 s01_aw_addr[2]
port 1148 nsew signal input
rlabel metal3 s 479200 104048 480000 104168 6 s01_aw_addr[30]
port 1149 nsew signal input
rlabel metal2 s 252466 119200 252522 120000 6 s01_aw_addr[31]
port 1150 nsew signal input
rlabel metal2 s 152002 119200 152058 120000 6 s01_aw_addr[3]
port 1151 nsew signal input
rlabel metal2 s 325238 0 325294 800 6 s01_aw_addr[4]
port 1152 nsew signal input
rlabel metal3 s 0 28568 800 28688 6 s01_aw_addr[5]
port 1153 nsew signal input
rlabel metal3 s 479200 30608 480000 30728 6 s01_aw_addr[6]
port 1154 nsew signal input
rlabel metal3 s 479200 54408 480000 54528 6 s01_aw_addr[7]
port 1155 nsew signal input
rlabel metal3 s 479200 112888 480000 113008 6 s01_aw_addr[8]
port 1156 nsew signal input
rlabel metal2 s 179050 119200 179106 120000 6 s01_aw_addr[9]
port 1157 nsew signal input
rlabel metal2 s 383198 119200 383254 120000 6 s01_aw_burst[0]
port 1158 nsew signal input
rlabel metal2 s 141698 0 141754 800 6 s01_aw_burst[1]
port 1159 nsew signal input
rlabel metal2 s 249246 119200 249302 120000 6 s01_aw_cache[0]
port 1160 nsew signal input
rlabel metal3 s 0 51688 800 51808 6 s01_aw_cache[1]
port 1161 nsew signal input
rlabel metal2 s 323306 119200 323362 120000 6 s01_aw_cache[2]
port 1162 nsew signal input
rlabel metal3 s 479200 91808 480000 91928 6 s01_aw_cache[3]
port 1163 nsew signal input
rlabel metal2 s 288530 119200 288586 120000 6 s01_aw_id[0]
port 1164 nsew signal input
rlabel metal2 s 383842 119200 383898 120000 6 s01_aw_id[1]
port 1165 nsew signal input
rlabel metal2 s 358082 0 358138 800 6 s01_aw_id[2]
port 1166 nsew signal input
rlabel metal2 s 287242 119200 287298 120000 6 s01_aw_id[3]
port 1167 nsew signal input
rlabel metal3 s 0 119008 800 119128 6 s01_aw_id[4]
port 1168 nsew signal input
rlabel metal2 s 277582 119200 277638 120000 6 s01_aw_id[5]
port 1169 nsew signal input
rlabel metal2 s 321374 119200 321430 120000 6 s01_aw_id[6]
port 1170 nsew signal input
rlabel metal2 s 428278 119200 428334 120000 6 s01_aw_id[7]
port 1171 nsew signal input
rlabel metal2 s 450818 119200 450874 120000 6 s01_aw_id[8]
port 1172 nsew signal input
rlabel metal2 s 311070 0 311126 800 6 s01_aw_id[9]
port 1173 nsew signal input
rlabel metal2 s 248602 0 248658 800 6 s01_aw_len[0]
port 1174 nsew signal input
rlabel metal2 s 144274 119200 144330 120000 6 s01_aw_len[1]
port 1175 nsew signal input
rlabel metal2 s 168102 0 168158 800 6 s01_aw_len[2]
port 1176 nsew signal input
rlabel metal3 s 479200 90448 480000 90568 6 s01_aw_len[3]
port 1177 nsew signal input
rlabel metal2 s 284022 119200 284078 120000 6 s01_aw_len[4]
port 1178 nsew signal input
rlabel metal2 s 267278 119200 267334 120000 6 s01_aw_len[5]
port 1179 nsew signal input
rlabel metal3 s 479200 21088 480000 21208 6 s01_aw_len[6]
port 1180 nsew signal input
rlabel metal2 s 269210 119200 269266 120000 6 s01_aw_len[7]
port 1181 nsew signal input
rlabel metal3 s 0 3408 800 3528 6 s01_aw_lock
port 1182 nsew signal input
rlabel metal2 s 83094 0 83150 800 6 s01_aw_prot[0]
port 1183 nsew signal input
rlabel metal3 s 0 89088 800 89208 6 s01_aw_prot[1]
port 1184 nsew signal input
rlabel metal3 s 0 2728 800 2848 6 s01_aw_prot[2]
port 1185 nsew signal input
rlabel metal2 s 234434 0 234490 800 6 s01_aw_qos[0]
port 1186 nsew signal input
rlabel metal2 s 477222 0 477278 800 6 s01_aw_qos[1]
port 1187 nsew signal input
rlabel metal2 s 465630 0 465686 800 6 s01_aw_qos[2]
port 1188 nsew signal input
rlabel metal3 s 479200 22448 480000 22568 6 s01_aw_qos[3]
port 1189 nsew signal input
rlabel metal2 s 186134 119200 186190 120000 6 s01_aw_ready
port 1190 nsew signal output
rlabel metal2 s 33506 119200 33562 120000 6 s01_aw_region[0]
port 1191 nsew signal input
rlabel metal2 s 157798 0 157854 800 6 s01_aw_region[1]
port 1192 nsew signal input
rlabel metal2 s 475934 119200 475990 120000 6 s01_aw_region[2]
port 1193 nsew signal input
rlabel metal2 s 206742 0 206798 800 6 s01_aw_region[3]
port 1194 nsew signal input
rlabel metal2 s 50894 119200 50950 120000 6 s01_aw_size[0]
port 1195 nsew signal input
rlabel metal3 s 0 78208 800 78328 6 s01_aw_size[1]
port 1196 nsew signal input
rlabel metal2 s 275650 119200 275706 120000 6 s01_aw_size[2]
port 1197 nsew signal input
rlabel metal3 s 479200 12928 480000 13048 6 s01_aw_user[-1]
port 1198 nsew signal input
rlabel metal2 s 231858 119200 231914 120000 6 s01_aw_user[0]
port 1199 nsew signal input
rlabel metal2 s 189998 0 190054 800 6 s01_aw_valid
port 1200 nsew signal input
rlabel metal2 s 103058 0 103114 800 6 s01_b_id[0]
port 1201 nsew signal output
rlabel metal2 s 403162 119200 403218 120000 6 s01_b_id[1]
port 1202 nsew signal output
rlabel metal2 s 311714 0 311770 800 6 s01_b_id[2]
port 1203 nsew signal output
rlabel metal2 s 455970 119200 456026 120000 6 s01_b_id[3]
port 1204 nsew signal output
rlabel metal2 s 23202 119200 23258 120000 6 s01_b_id[4]
port 1205 nsew signal output
rlabel metal2 s 306562 119200 306618 120000 6 s01_b_id[5]
port 1206 nsew signal output
rlabel metal2 s 215114 119200 215170 120000 6 s01_b_id[6]
port 1207 nsew signal output
rlabel metal2 s 44454 119200 44510 120000 6 s01_b_id[7]
port 1208 nsew signal output
rlabel metal2 s 96618 119200 96674 120000 6 s01_b_id[8]
port 1209 nsew signal output
rlabel metal2 s 365810 0 365866 800 6 s01_b_id[9]
port 1210 nsew signal output
rlabel metal2 s 438582 119200 438638 120000 6 s01_b_ready
port 1211 nsew signal input
rlabel metal2 s 208030 119200 208086 120000 6 s01_b_resp[0]
port 1212 nsew signal output
rlabel metal2 s 160374 0 160430 800 6 s01_b_resp[1]
port 1213 nsew signal output
rlabel metal2 s 88246 0 88302 800 6 s01_b_user[-1]
port 1214 nsew signal output
rlabel metal2 s 479154 119200 479210 120000 6 s01_b_user[0]
port 1215 nsew signal output
rlabel metal3 s 0 107448 800 107568 6 s01_b_valid
port 1216 nsew signal output
rlabel metal2 s 38014 119200 38070 120000 6 s01_r_data[0]
port 1217 nsew signal output
rlabel metal3 s 0 67328 800 67448 6 s01_r_data[10]
port 1218 nsew signal output
rlabel metal3 s 0 75488 800 75608 6 s01_r_data[11]
port 1219 nsew signal output
rlabel metal2 s 415398 119200 415454 120000 6 s01_r_data[12]
port 1220 nsew signal output
rlabel metal2 s 14830 0 14886 800 6 s01_r_data[13]
port 1221 nsew signal output
rlabel metal2 s 204166 0 204222 800 6 s01_r_data[14]
port 1222 nsew signal output
rlabel metal2 s 445022 119200 445078 120000 6 s01_r_data[15]
port 1223 nsew signal output
rlabel metal2 s 80518 119200 80574 120000 6 s01_r_data[16]
port 1224 nsew signal output
rlabel metal3 s 479200 72768 480000 72888 6 s01_r_data[17]
port 1225 nsew signal output
rlabel metal2 s 274362 119200 274418 120000 6 s01_r_data[18]
port 1226 nsew signal output
rlabel metal3 s 0 36728 800 36848 6 s01_r_data[19]
port 1227 nsew signal output
rlabel metal3 s 0 54408 800 54528 6 s01_r_data[1]
port 1228 nsew signal output
rlabel metal2 s 173898 0 173954 800 6 s01_r_data[20]
port 1229 nsew signal output
rlabel metal2 s 475290 0 475346 800 6 s01_r_data[21]
port 1230 nsew signal output
rlabel metal2 s 59266 119200 59322 120000 6 s01_r_data[22]
port 1231 nsew signal output
rlabel metal2 s 140410 0 140466 800 6 s01_r_data[23]
port 1232 nsew signal output
rlabel metal2 s 291750 119200 291806 120000 6 s01_r_data[24]
port 1233 nsew signal output
rlabel metal2 s 325238 119200 325294 120000 6 s01_r_data[25]
port 1234 nsew signal output
rlabel metal2 s 84382 0 84438 800 6 s01_r_data[26]
port 1235 nsew signal output
rlabel metal2 s 307206 119200 307262 120000 6 s01_r_data[27]
port 1236 nsew signal output
rlabel metal3 s 479200 23808 480000 23928 6 s01_r_data[28]
port 1237 nsew signal output
rlabel metal2 s 374826 0 374882 800 6 s01_r_data[29]
port 1238 nsew signal output
rlabel metal2 s 51538 119200 51594 120000 6 s01_r_data[2]
port 1239 nsew signal output
rlabel metal3 s 0 18368 800 18488 6 s01_r_data[30]
port 1240 nsew signal output
rlabel metal2 s 478510 119200 478566 120000 6 s01_r_data[31]
port 1241 nsew signal output
rlabel metal2 s 443734 0 443790 800 6 s01_r_data[3]
port 1242 nsew signal output
rlabel metal2 s 347134 0 347190 800 6 s01_r_data[4]
port 1243 nsew signal output
rlabel metal2 s 314934 119200 314990 120000 6 s01_r_data[5]
port 1244 nsew signal output
rlabel metal2 s 94686 119200 94742 120000 6 s01_r_data[6]
port 1245 nsew signal output
rlabel metal3 s 0 42168 800 42288 6 s01_r_data[7]
port 1246 nsew signal output
rlabel metal2 s 224774 0 224830 800 6 s01_r_data[8]
port 1247 nsew signal output
rlabel metal2 s 78586 119200 78642 120000 6 s01_r_data[9]
port 1248 nsew signal output
rlabel metal2 s 350998 119200 351054 120000 6 s01_r_id[0]
port 1249 nsew signal output
rlabel metal2 s 76654 0 76710 800 6 s01_r_id[1]
port 1250 nsew signal output
rlabel metal2 s 435362 119200 435418 120000 6 s01_r_id[2]
port 1251 nsew signal output
rlabel metal3 s 479200 88408 480000 88528 6 s01_r_id[3]
port 1252 nsew signal output
rlabel metal2 s 229926 0 229982 800 6 s01_r_id[4]
port 1253 nsew signal output
rlabel metal3 s 479200 48968 480000 49088 6 s01_r_id[5]
port 1254 nsew signal output
rlabel metal2 s 134614 119200 134670 120000 6 s01_r_id[6]
port 1255 nsew signal output
rlabel metal2 s 426990 0 427046 800 6 s01_r_id[7]
port 1256 nsew signal output
rlabel metal2 s 467562 0 467618 800 6 s01_r_id[8]
port 1257 nsew signal output
rlabel metal3 s 479200 27888 480000 28008 6 s01_r_id[9]
port 1258 nsew signal output
rlabel metal2 s 137834 0 137890 800 6 s01_r_last
port 1259 nsew signal output
rlabel metal2 s 422482 119200 422538 120000 6 s01_r_ready
port 1260 nsew signal input
rlabel metal2 s 229282 0 229338 800 6 s01_r_resp[0]
port 1261 nsew signal output
rlabel metal2 s 466274 119200 466330 120000 6 s01_r_resp[1]
port 1262 nsew signal output
rlabel metal2 s 202234 119200 202290 120000 6 s01_r_user[-1]
port 1263 nsew signal output
rlabel metal2 s 331034 0 331090 800 6 s01_r_user[0]
port 1264 nsew signal output
rlabel metal3 s 0 38088 800 38208 6 s01_r_valid
port 1265 nsew signal output
rlabel metal2 s 30930 0 30986 800 6 s01_w_data[0]
port 1266 nsew signal input
rlabel metal3 s 0 93848 800 93968 6 s01_w_data[10]
port 1267 nsew signal input
rlabel metal2 s 396078 0 396134 800 6 s01_w_data[11]
port 1268 nsew signal input
rlabel metal3 s 479200 4088 480000 4208 6 s01_w_data[12]
port 1269 nsew signal input
rlabel metal2 s 131394 119200 131450 120000 6 s01_w_data[13]
port 1270 nsew signal input
rlabel metal3 s 479200 114248 480000 114368 6 s01_w_data[14]
port 1271 nsew signal input
rlabel metal2 s 257618 0 257674 800 6 s01_w_data[15]
port 1272 nsew signal input
rlabel metal2 s 34794 0 34850 800 6 s01_w_data[16]
port 1273 nsew signal input
rlabel metal2 s 107566 119200 107622 120000 6 s01_w_data[17]
port 1274 nsew signal input
rlabel metal2 s 275650 0 275706 800 6 s01_w_data[18]
port 1275 nsew signal input
rlabel metal2 s 45742 119200 45798 120000 6 s01_w_data[19]
port 1276 nsew signal input
rlabel metal2 s 291750 0 291806 800 6 s01_w_data[1]
port 1277 nsew signal input
rlabel metal2 s 382554 119200 382610 120000 6 s01_w_data[20]
port 1278 nsew signal input
rlabel metal3 s 479200 2048 480000 2168 6 s01_w_data[21]
port 1279 nsew signal input
rlabel metal2 s 396722 119200 396778 120000 6 s01_w_data[22]
port 1280 nsew signal input
rlabel metal2 s 244738 0 244794 800 6 s01_w_data[23]
port 1281 nsew signal input
rlabel metal2 s 89534 119200 89590 120000 6 s01_w_data[24]
port 1282 nsew signal input
rlabel metal2 s 135902 119200 135958 120000 6 s01_w_data[25]
port 1283 nsew signal input
rlabel metal3 s 0 21088 800 21208 6 s01_w_data[26]
port 1284 nsew signal input
rlabel metal2 s 125598 119200 125654 120000 6 s01_w_data[27]
port 1285 nsew signal input
rlabel metal2 s 63130 0 63186 800 6 s01_w_data[28]
port 1286 nsew signal input
rlabel metal2 s 354862 0 354918 800 6 s01_w_data[29]
port 1287 nsew signal input
rlabel metal2 s 395434 0 395490 800 6 s01_w_data[2]
port 1288 nsew signal input
rlabel metal2 s 385130 119200 385186 120000 6 s01_w_data[30]
port 1289 nsew signal input
rlabel metal3 s 479200 70048 480000 70168 6 s01_w_data[31]
port 1290 nsew signal input
rlabel metal3 s 479200 29928 480000 30048 6 s01_w_data[3]
port 1291 nsew signal input
rlabel metal3 s 0 53728 800 53848 6 s01_w_data[4]
port 1292 nsew signal input
rlabel metal2 s 316866 0 316922 800 6 s01_w_data[5]
port 1293 nsew signal input
rlabel metal2 s 164882 0 164938 800 6 s01_w_data[6]
port 1294 nsew signal input
rlabel metal2 s 145562 119200 145618 120000 6 s01_w_data[7]
port 1295 nsew signal input
rlabel metal2 s 240230 0 240286 800 6 s01_w_data[8]
port 1296 nsew signal input
rlabel metal2 s 332322 0 332378 800 6 s01_w_data[9]
port 1297 nsew signal input
rlabel metal2 s 265346 0 265402 800 6 s01_w_last
port 1298 nsew signal input
rlabel metal3 s 0 9528 800 9648 6 s01_w_ready
port 1299 nsew signal output
rlabel metal2 s 390282 119200 390338 120000 6 s01_w_strb[0]
port 1300 nsew signal input
rlabel metal2 s 218978 0 219034 800 6 s01_w_strb[1]
port 1301 nsew signal input
rlabel metal2 s 479798 0 479854 800 6 s01_w_strb[2]
port 1302 nsew signal input
rlabel metal2 s 412822 0 412878 800 6 s01_w_strb[3]
port 1303 nsew signal input
rlabel metal3 s 479200 51688 480000 51808 6 s01_w_user[-1]
port 1304 nsew signal input
rlabel metal3 s 479200 27208 480000 27328 6 s01_w_user[0]
port 1305 nsew signal input
rlabel metal2 s 162950 0 163006 800 6 s01_w_valid
port 1306 nsew signal input
rlabel metal2 s 6458 0 6514 800 6 s02_ar_addr[0]
port 1307 nsew signal input
rlabel metal2 s 302698 0 302754 800 6 s02_ar_addr[10]
port 1308 nsew signal input
rlabel metal2 s 218334 119200 218390 120000 6 s02_ar_addr[11]
port 1309 nsew signal input
rlabel metal2 s 350354 0 350410 800 6 s02_ar_addr[12]
port 1310 nsew signal input
rlabel metal2 s 258906 119200 258962 120000 6 s02_ar_addr[13]
port 1311 nsew signal input
rlabel metal2 s 18 0 74 800 6 s02_ar_addr[14]
port 1312 nsew signal input
rlabel metal3 s 0 96568 800 96688 6 s02_ar_addr[15]
port 1313 nsew signal input
rlabel metal2 s 426990 119200 427046 120000 6 s02_ar_addr[16]
port 1314 nsew signal input
rlabel metal2 s 227350 0 227406 800 6 s02_ar_addr[17]
port 1315 nsew signal input
rlabel metal3 s 0 62568 800 62688 6 s02_ar_addr[18]
port 1316 nsew signal input
rlabel metal2 s 109498 0 109554 800 6 s02_ar_addr[19]
port 1317 nsew signal input
rlabel metal2 s 165526 119200 165582 120000 6 s02_ar_addr[1]
port 1318 nsew signal input
rlabel metal2 s 318154 0 318210 800 6 s02_ar_addr[20]
port 1319 nsew signal input
rlabel metal3 s 0 95208 800 95328 6 s02_ar_addr[21]
port 1320 nsew signal input
rlabel metal2 s 174542 119200 174598 120000 6 s02_ar_addr[22]
port 1321 nsew signal input
rlabel metal2 s 122378 0 122434 800 6 s02_ar_addr[23]
port 1322 nsew signal input
rlabel metal2 s 262126 119200 262182 120000 6 s02_ar_addr[24]
port 1323 nsew signal input
rlabel metal2 s 325882 0 325938 800 6 s02_ar_addr[25]
port 1324 nsew signal input
rlabel metal3 s 479200 65968 480000 66088 6 s02_ar_addr[26]
port 1325 nsew signal input
rlabel metal2 s 25778 119200 25834 120000 6 s02_ar_addr[27]
port 1326 nsew signal input
rlabel metal2 s 173898 119200 173954 120000 6 s02_ar_addr[28]
port 1327 nsew signal input
rlabel metal2 s 420550 0 420606 800 6 s02_ar_addr[29]
port 1328 nsew signal input
rlabel metal2 s 187422 0 187478 800 6 s02_ar_addr[2]
port 1329 nsew signal input
rlabel metal2 s 220266 0 220322 800 6 s02_ar_addr[30]
port 1330 nsew signal input
rlabel metal2 s 261482 119200 261538 120000 6 s02_ar_addr[31]
port 1331 nsew signal input
rlabel metal3 s 0 33328 800 33448 6 s02_ar_addr[3]
port 1332 nsew signal input
rlabel metal2 s 191286 119200 191342 120000 6 s02_ar_addr[4]
port 1333 nsew signal input
rlabel metal2 s 106278 0 106334 800 6 s02_ar_addr[5]
port 1334 nsew signal input
rlabel metal2 s 432142 119200 432198 120000 6 s02_ar_addr[6]
port 1335 nsew signal input
rlabel metal2 s 299478 0 299534 800 6 s02_ar_addr[7]
port 1336 nsew signal input
rlabel metal2 s 253110 119200 253166 120000 6 s02_ar_addr[8]
port 1337 nsew signal input
rlabel metal2 s 439226 119200 439282 120000 6 s02_ar_addr[9]
port 1338 nsew signal input
rlabel metal3 s 0 1368 800 1488 6 s02_ar_burst[0]
port 1339 nsew signal input
rlabel metal2 s 177762 119200 177818 120000 6 s02_ar_burst[1]
port 1340 nsew signal input
rlabel metal2 s 164238 0 164294 800 6 s02_ar_cache[0]
port 1341 nsew signal input
rlabel metal2 s 14830 119200 14886 120000 6 s02_ar_cache[1]
port 1342 nsew signal input
rlabel metal2 s 295614 0 295670 800 6 s02_ar_cache[2]
port 1343 nsew signal input
rlabel metal2 s 463054 119200 463110 120000 6 s02_ar_cache[3]
port 1344 nsew signal input
rlabel metal2 s 77942 0 77998 800 6 s02_ar_id[0]
port 1345 nsew signal input
rlabel metal2 s 109498 119200 109554 120000 6 s02_ar_id[1]
port 1346 nsew signal input
rlabel metal2 s 233790 0 233846 800 6 s02_ar_id[2]
port 1347 nsew signal input
rlabel metal2 s 207386 0 207442 800 6 s02_ar_id[3]
port 1348 nsew signal input
rlabel metal2 s 299478 119200 299534 120000 6 s02_ar_id[4]
port 1349 nsew signal input
rlabel metal3 s 479200 76848 480000 76968 6 s02_ar_id[5]
port 1350 nsew signal input
rlabel metal2 s 421194 0 421250 800 6 s02_ar_id[6]
port 1351 nsew signal input
rlabel metal2 s 453394 119200 453450 120000 6 s02_ar_id[7]
port 1352 nsew signal input
rlabel metal2 s 256330 0 256386 800 6 s02_ar_id[8]
port 1353 nsew signal input
rlabel metal2 s 142986 0 143042 800 6 s02_ar_id[9]
port 1354 nsew signal input
rlabel metal2 s 139766 119200 139822 120000 6 s02_ar_len[0]
port 1355 nsew signal input
rlabel metal2 s 357438 119200 357494 120000 6 s02_ar_len[1]
port 1356 nsew signal input
rlabel metal3 s 0 38768 800 38888 6 s02_ar_len[2]
port 1357 nsew signal input
rlabel metal3 s 479200 106088 480000 106208 6 s02_ar_len[3]
port 1358 nsew signal input
rlabel metal2 s 324594 0 324650 800 6 s02_ar_len[4]
port 1359 nsew signal input
rlabel metal3 s 479200 10888 480000 11008 6 s02_ar_len[5]
port 1360 nsew signal input
rlabel metal2 s 416042 119200 416098 120000 6 s02_ar_len[6]
port 1361 nsew signal input
rlabel metal2 s 146850 119200 146906 120000 6 s02_ar_len[7]
port 1362 nsew signal input
rlabel metal2 s 31574 0 31630 800 6 s02_ar_lock
port 1363 nsew signal input
rlabel metal2 s 208674 0 208730 800 6 s02_ar_prot[0]
port 1364 nsew signal input
rlabel metal2 s 111430 0 111486 800 6 s02_ar_prot[1]
port 1365 nsew signal input
rlabel metal2 s 455970 0 456026 800 6 s02_ar_prot[2]
port 1366 nsew signal input
rlabel metal2 s 25778 0 25834 800 6 s02_ar_qos[0]
port 1367 nsew signal input
rlabel metal2 s 114650 0 114706 800 6 s02_ar_qos[1]
port 1368 nsew signal input
rlabel metal3 s 0 688 800 808 6 s02_ar_qos[2]
port 1369 nsew signal input
rlabel metal2 s 334254 119200 334310 120000 6 s02_ar_qos[3]
port 1370 nsew signal input
rlabel metal3 s 479200 67328 480000 67448 6 s02_ar_ready
port 1371 nsew signal output
rlabel metal2 s 41234 0 41290 800 6 s02_ar_region[0]
port 1372 nsew signal input
rlabel metal3 s 479200 36048 480000 36168 6 s02_ar_region[1]
port 1373 nsew signal input
rlabel metal2 s 266634 0 266690 800 6 s02_ar_region[2]
port 1374 nsew signal input
rlabel metal2 s 268566 119200 268622 120000 6 s02_ar_region[3]
port 1375 nsew signal input
rlabel metal2 s 246026 0 246082 800 6 s02_ar_size[0]
port 1376 nsew signal input
rlabel metal3 s 479200 112208 480000 112328 6 s02_ar_size[1]
port 1377 nsew signal input
rlabel metal2 s 318798 119200 318854 120000 6 s02_ar_size[2]
port 1378 nsew signal input
rlabel metal2 s 276938 119200 276994 120000 6 s02_ar_user[-1]
port 1379 nsew signal input
rlabel metal2 s 183558 119200 183614 120000 6 s02_ar_user[0]
port 1380 nsew signal input
rlabel metal2 s 325882 119200 325938 120000 6 s02_ar_valid
port 1381 nsew signal input
rlabel metal2 s 54114 119200 54170 120000 6 s02_aw_addr[0]
port 1382 nsew signal input
rlabel metal2 s 124954 0 125010 800 6 s02_aw_addr[10]
port 1383 nsew signal input
rlabel metal2 s 401874 0 401930 800 6 s02_aw_addr[11]
port 1384 nsew signal input
rlabel metal3 s 479200 17688 480000 17808 6 s02_aw_addr[12]
port 1385 nsew signal input
rlabel metal3 s 0 104728 800 104848 6 s02_aw_addr[13]
port 1386 nsew signal input
rlabel metal2 s 139122 119200 139178 120000 6 s02_aw_addr[14]
port 1387 nsew signal input
rlabel metal3 s 0 71408 800 71528 6 s02_aw_addr[15]
port 1388 nsew signal input
rlabel metal2 s 401230 119200 401286 120000 6 s02_aw_addr[16]
port 1389 nsew signal input
rlabel metal2 s 450174 119200 450230 120000 6 s02_aw_addr[17]
port 1390 nsew signal input
rlabel metal2 s 303342 119200 303398 120000 6 s02_aw_addr[18]
port 1391 nsew signal input
rlabel metal2 s 370318 119200 370374 120000 6 s02_aw_addr[19]
port 1392 nsew signal input
rlabel metal2 s 343270 0 343326 800 6 s02_aw_addr[1]
port 1393 nsew signal input
rlabel metal3 s 0 5448 800 5568 6 s02_aw_addr[20]
port 1394 nsew signal input
rlabel metal2 s 329102 0 329158 800 6 s02_aw_addr[21]
port 1395 nsew signal input
rlabel metal2 s 392858 0 392914 800 6 s02_aw_addr[22]
port 1396 nsew signal input
rlabel metal2 s 66350 0 66406 800 6 s02_aw_addr[23]
port 1397 nsew signal input
rlabel metal2 s 101126 0 101182 800 6 s02_aw_addr[24]
port 1398 nsew signal input
rlabel metal2 s 350998 0 351054 800 6 s02_aw_addr[25]
port 1399 nsew signal input
rlabel metal2 s 477866 0 477922 800 6 s02_aw_addr[26]
port 1400 nsew signal input
rlabel metal2 s 410246 119200 410302 120000 6 s02_aw_addr[27]
port 1401 nsew signal input
rlabel metal2 s 168746 119200 168802 120000 6 s02_aw_addr[28]
port 1402 nsew signal input
rlabel metal2 s 153934 119200 153990 120000 6 s02_aw_addr[29]
port 1403 nsew signal input
rlabel metal2 s 97906 119200 97962 120000 6 s02_aw_addr[2]
port 1404 nsew signal input
rlabel metal2 s 123022 0 123078 800 6 s02_aw_addr[30]
port 1405 nsew signal input
rlabel metal2 s 378690 119200 378746 120000 6 s02_aw_addr[31]
port 1406 nsew signal input
rlabel metal2 s 383198 0 383254 800 6 s02_aw_addr[3]
port 1407 nsew signal input
rlabel metal2 s 82450 119200 82506 120000 6 s02_aw_addr[4]
port 1408 nsew signal input
rlabel metal2 s 78586 0 78642 800 6 s02_aw_addr[5]
port 1409 nsew signal input
rlabel metal2 s 425058 119200 425114 120000 6 s02_aw_addr[6]
port 1410 nsew signal input
rlabel metal2 s 247314 119200 247370 120000 6 s02_aw_addr[7]
port 1411 nsew signal input
rlabel metal2 s 226706 119200 226762 120000 6 s02_aw_addr[8]
port 1412 nsew signal input
rlabel metal2 s 291106 119200 291162 120000 6 s02_aw_addr[9]
port 1413 nsew signal input
rlabel metal2 s 310426 119200 310482 120000 6 s02_aw_burst[0]
port 1414 nsew signal input
rlabel metal2 s 313646 119200 313702 120000 6 s02_aw_burst[1]
port 1415 nsew signal input
rlabel metal3 s 0 24488 800 24608 6 s02_aw_cache[0]
port 1416 nsew signal input
rlabel metal2 s 195794 119200 195850 120000 6 s02_aw_cache[1]
port 1417 nsew signal input
rlabel metal3 s 0 52368 800 52488 6 s02_aw_cache[2]
port 1418 nsew signal input
rlabel metal2 s 5170 0 5226 800 6 s02_aw_cache[3]
port 1419 nsew signal input
rlabel metal2 s 316222 0 316278 800 6 s02_aw_id[0]
port 1420 nsew signal input
rlabel metal2 s 214470 0 214526 800 6 s02_aw_id[1]
port 1421 nsew signal input
rlabel metal2 s 426346 0 426402 800 6 s02_aw_id[2]
port 1422 nsew signal input
rlabel metal2 s 239586 119200 239642 120000 6 s02_aw_id[3]
port 1423 nsew signal input
rlabel metal2 s 457258 0 457314 800 6 s02_aw_id[4]
port 1424 nsew signal input
rlabel metal2 s 5170 119200 5226 120000 6 s02_aw_id[5]
port 1425 nsew signal input
rlabel metal2 s 16118 0 16174 800 6 s02_aw_id[6]
port 1426 nsew signal input
rlabel metal2 s 80518 0 80574 800 6 s02_aw_id[7]
port 1427 nsew signal input
rlabel metal2 s 179050 0 179106 800 6 s02_aw_id[8]
port 1428 nsew signal input
rlabel metal2 s 202878 119200 202934 120000 6 s02_aw_id[9]
port 1429 nsew signal input
rlabel metal2 s 321374 0 321430 800 6 s02_aw_len[0]
port 1430 nsew signal input
rlabel metal2 s 152646 0 152702 800 6 s02_aw_len[1]
port 1431 nsew signal input
rlabel metal2 s 300122 0 300178 800 6 s02_aw_len[2]
port 1432 nsew signal input
rlabel metal3 s 0 99288 800 99408 6 s02_aw_len[3]
port 1433 nsew signal input
rlabel metal2 s 412822 119200 412878 120000 6 s02_aw_len[4]
port 1434 nsew signal input
rlabel metal2 s 305918 0 305974 800 6 s02_aw_len[5]
port 1435 nsew signal input
rlabel metal2 s 20626 119200 20682 120000 6 s02_aw_len[6]
port 1436 nsew signal input
rlabel metal2 s 388994 0 389050 800 6 s02_aw_len[7]
port 1437 nsew signal input
rlabel metal2 s 433430 119200 433486 120000 6 s02_aw_lock
port 1438 nsew signal input
rlabel metal2 s 168102 119200 168158 120000 6 s02_aw_prot[0]
port 1439 nsew signal input
rlabel metal3 s 479200 116288 480000 116408 6 s02_aw_prot[1]
port 1440 nsew signal input
rlabel metal2 s 296902 0 296958 800 6 s02_aw_prot[2]
port 1441 nsew signal input
rlabel metal2 s 255042 119200 255098 120000 6 s02_aw_qos[0]
port 1442 nsew signal input
rlabel metal2 s 425702 0 425758 800 6 s02_aw_qos[1]
port 1443 nsew signal input
rlabel metal2 s 147494 119200 147550 120000 6 s02_aw_qos[2]
port 1444 nsew signal input
rlabel metal2 s 357438 0 357494 800 6 s02_aw_qos[3]
port 1445 nsew signal input
rlabel metal2 s 18050 119200 18106 120000 6 s02_aw_ready
port 1446 nsew signal output
rlabel metal2 s 48962 0 49018 800 6 s02_aw_region[0]
port 1447 nsew signal input
rlabel metal3 s 479200 97928 480000 98048 6 s02_aw_region[1]
port 1448 nsew signal input
rlabel metal2 s 215114 0 215170 800 6 s02_aw_region[2]
port 1449 nsew signal input
rlabel metal2 s 445666 119200 445722 120000 6 s02_aw_region[3]
port 1450 nsew signal input
rlabel metal2 s 97262 0 97318 800 6 s02_aw_size[0]
port 1451 nsew signal input
rlabel metal2 s 360014 0 360070 800 6 s02_aw_size[1]
port 1452 nsew signal input
rlabel metal2 s 56046 119200 56102 120000 6 s02_aw_size[2]
port 1453 nsew signal input
rlabel metal2 s 270498 119200 270554 120000 6 s02_aw_user[-1]
port 1454 nsew signal input
rlabel metal2 s 413466 119200 413522 120000 6 s02_aw_user[0]
port 1455 nsew signal input
rlabel metal2 s 48318 119200 48374 120000 6 s02_aw_valid
port 1456 nsew signal input
rlabel metal2 s 83738 119200 83794 120000 6 s02_b_id[0]
port 1457 nsew signal output
rlabel metal2 s 437938 0 437994 800 6 s02_b_id[1]
port 1458 nsew signal output
rlabel metal2 s 32218 119200 32274 120000 6 s02_b_id[2]
port 1459 nsew signal output
rlabel metal3 s 479200 19048 480000 19168 6 s02_b_id[3]
port 1460 nsew signal output
rlabel metal2 s 213826 119200 213882 120000 6 s02_b_id[4]
port 1461 nsew signal output
rlabel metal2 s 138478 119200 138534 120000 6 s02_b_id[5]
port 1462 nsew signal output
rlabel metal3 s 0 116288 800 116408 6 s02_b_id[6]
port 1463 nsew signal output
rlabel metal2 s 34150 0 34206 800 6 s02_b_id[7]
port 1464 nsew signal output
rlabel metal2 s 204810 0 204866 800 6 s02_b_id[8]
port 1465 nsew signal output
rlabel metal2 s 441802 119200 441858 120000 6 s02_b_id[9]
port 1466 nsew signal output
rlabel metal3 s 0 27888 800 28008 6 s02_b_ready
port 1467 nsew signal input
rlabel metal2 s 231858 0 231914 800 6 s02_b_resp[0]
port 1468 nsew signal output
rlabel metal3 s 479200 105408 480000 105528 6 s02_b_resp[1]
port 1469 nsew signal output
rlabel metal2 s 474002 0 474058 800 6 s02_b_user[-1]
port 1470 nsew signal output
rlabel metal2 s 347778 0 347834 800 6 s02_b_user[0]
port 1471 nsew signal output
rlabel metal3 s 0 19048 800 19168 6 s02_b_valid
port 1472 nsew signal output
rlabel metal2 s 332966 119200 333022 120000 6 s02_r_data[0]
port 1473 nsew signal output
rlabel metal2 s 203522 0 203578 800 6 s02_r_data[10]
port 1474 nsew signal output
rlabel metal2 s 289174 0 289230 800 6 s02_r_data[11]
port 1475 nsew signal output
rlabel metal3 s 0 42848 800 42968 6 s02_r_data[12]
port 1476 nsew signal output
rlabel metal2 s 52826 119200 52882 120000 6 s02_r_data[13]
port 1477 nsew signal output
rlabel metal2 s 194506 0 194562 800 6 s02_r_data[14]
port 1478 nsew signal output
rlabel metal2 s 38014 0 38070 800 6 s02_r_data[15]
port 1479 nsew signal output
rlabel metal2 s 136546 119200 136602 120000 6 s02_r_data[16]
port 1480 nsew signal output
rlabel metal3 s 479200 80928 480000 81048 6 s02_r_data[17]
port 1481 nsew signal output
rlabel metal2 s 387062 119200 387118 120000 6 s02_r_data[18]
port 1482 nsew signal output
rlabel metal2 s 136546 0 136602 800 6 s02_r_data[19]
port 1483 nsew signal output
rlabel metal2 s 303986 119200 304042 120000 6 s02_r_data[1]
port 1484 nsew signal output
rlabel metal3 s 479200 17008 480000 17128 6 s02_r_data[20]
port 1485 nsew signal output
rlabel metal2 s 271786 0 271842 800 6 s02_r_data[21]
port 1486 nsew signal output
rlabel metal2 s 300766 119200 300822 120000 6 s02_r_data[22]
port 1487 nsew signal output
rlabel metal2 s 260838 0 260894 800 6 s02_r_data[23]
port 1488 nsew signal output
rlabel metal2 s 110142 0 110198 800 6 s02_r_data[24]
port 1489 nsew signal output
rlabel metal2 s 17406 0 17462 800 6 s02_r_data[25]
port 1490 nsew signal output
rlabel metal2 s 345202 0 345258 800 6 s02_r_data[26]
port 1491 nsew signal output
rlabel metal2 s 437294 0 437350 800 6 s02_r_data[27]
port 1492 nsew signal output
rlabel metal2 s 157154 119200 157210 120000 6 s02_r_data[28]
port 1493 nsew signal output
rlabel metal2 s 434718 119200 434774 120000 6 s02_r_data[29]
port 1494 nsew signal output
rlabel metal3 s 0 20408 800 20528 6 s02_r_data[2]
port 1495 nsew signal output
rlabel metal2 s 2594 119200 2650 120000 6 s02_r_data[30]
port 1496 nsew signal output
rlabel metal3 s 0 114248 800 114368 6 s02_r_data[31]
port 1497 nsew signal output
rlabel metal2 s 14186 0 14242 800 6 s02_r_data[3]
port 1498 nsew signal output
rlabel metal2 s 73434 0 73490 800 6 s02_r_data[4]
port 1499 nsew signal output
rlabel metal3 s 479200 34688 480000 34808 6 s02_r_data[5]
port 1500 nsew signal output
rlabel metal2 s 193862 0 193918 800 6 s02_r_data[6]
port 1501 nsew signal output
rlabel metal2 s 298190 119200 298246 120000 6 s02_r_data[7]
port 1502 nsew signal output
rlabel metal2 s 379978 119200 380034 120000 6 s02_r_data[8]
port 1503 nsew signal output
rlabel metal2 s 90822 119200 90878 120000 6 s02_r_data[9]
port 1504 nsew signal output
rlabel metal2 s 52182 0 52238 800 6 s02_r_id[0]
port 1505 nsew signal output
rlabel metal3 s 479200 56448 480000 56568 6 s02_r_id[1]
port 1506 nsew signal output
rlabel metal2 s 396078 119200 396134 120000 6 s02_r_id[2]
port 1507 nsew signal output
rlabel metal3 s 0 64608 800 64728 6 s02_r_id[3]
port 1508 nsew signal output
rlabel metal3 s 479200 114928 480000 115048 6 s02_r_id[4]
port 1509 nsew signal output
rlabel metal2 s 438582 0 438638 800 6 s02_r_id[5]
port 1510 nsew signal output
rlabel metal2 s 228638 0 228694 800 6 s02_r_id[6]
port 1511 nsew signal output
rlabel metal2 s 363878 119200 363934 120000 6 s02_r_id[7]
port 1512 nsew signal output
rlabel metal2 s 171966 119200 172022 120000 6 s02_r_id[8]
port 1513 nsew signal output
rlabel metal2 s 103702 0 103758 800 6 s02_r_id[9]
port 1514 nsew signal output
rlabel metal3 s 479200 46248 480000 46368 6 s02_r_last
port 1515 nsew signal output
rlabel metal2 s 267278 0 267334 800 6 s02_r_ready
port 1516 nsew signal input
rlabel metal2 s 421838 0 421894 800 6 s02_r_resp[0]
port 1517 nsew signal output
rlabel metal3 s 0 68008 800 68128 6 s02_r_resp[1]
port 1518 nsew signal output
rlabel metal2 s 336830 0 336886 800 6 s02_r_user[-1]
port 1519 nsew signal output
rlabel metal2 s 52826 0 52882 800 6 s02_r_user[0]
port 1520 nsew signal output
rlabel metal2 s 161018 0 161074 800 6 s02_r_valid
port 1521 nsew signal output
rlabel metal2 s 462410 0 462466 800 6 s02_w_data[0]
port 1522 nsew signal input
rlabel metal2 s 366454 119200 366510 120000 6 s02_w_data[10]
port 1523 nsew signal input
rlabel metal2 s 466918 119200 466974 120000 6 s02_w_data[11]
port 1524 nsew signal input
rlabel metal2 s 337474 0 337530 800 6 s02_w_data[12]
port 1525 nsew signal input
rlabel metal2 s 26422 0 26478 800 6 s02_w_data[13]
port 1526 nsew signal input
rlabel metal3 s 479200 21768 480000 21888 6 s02_w_data[14]
port 1527 nsew signal input
rlabel metal2 s 7102 0 7158 800 6 s02_w_data[15]
port 1528 nsew signal input
rlabel metal2 s 464342 119200 464398 120000 6 s02_w_data[16]
port 1529 nsew signal input
rlabel metal2 s 363234 119200 363290 120000 6 s02_w_data[17]
port 1530 nsew signal input
rlabel metal2 s 353574 0 353630 800 6 s02_w_data[18]
port 1531 nsew signal input
rlabel metal2 s 355506 119200 355562 120000 6 s02_w_data[19]
port 1532 nsew signal input
rlabel metal2 s 213182 0 213238 800 6 s02_w_data[1]
port 1533 nsew signal input
rlabel metal3 s 0 32648 800 32768 6 s02_w_data[20]
port 1534 nsew signal input
rlabel metal2 s 211894 0 211950 800 6 s02_w_data[21]
port 1535 nsew signal input
rlabel metal2 s 662 0 718 800 6 s02_w_data[22]
port 1536 nsew signal input
rlabel metal2 s 247958 0 248014 800 6 s02_w_data[23]
port 1537 nsew signal input
rlabel metal3 s 0 95888 800 96008 6 s02_w_data[24]
port 1538 nsew signal input
rlabel metal2 s 100482 119200 100538 120000 6 s02_w_data[25]
port 1539 nsew signal input
rlabel metal2 s 229282 119200 229338 120000 6 s02_w_data[26]
port 1540 nsew signal input
rlabel metal3 s 0 55088 800 55208 6 s02_w_data[27]
port 1541 nsew signal input
rlabel metal2 s 65062 0 65118 800 6 s02_w_data[28]
port 1542 nsew signal input
rlabel metal2 s 23202 0 23258 800 6 s02_w_data[29]
port 1543 nsew signal input
rlabel metal2 s 311070 119200 311126 120000 6 s02_w_data[2]
port 1544 nsew signal input
rlabel metal2 s 243450 119200 243506 120000 6 s02_w_data[30]
port 1545 nsew signal input
rlabel metal2 s 166814 0 166870 800 6 s02_w_data[31]
port 1546 nsew signal input
rlabel metal2 s 367742 119200 367798 120000 6 s02_w_data[3]
port 1547 nsew signal input
rlabel metal2 s 392214 0 392270 800 6 s02_w_data[4]
port 1548 nsew signal input
rlabel metal2 s 54758 119200 54814 120000 6 s02_w_data[5]
port 1549 nsew signal input
rlabel metal3 s 479200 63248 480000 63368 6 s02_w_data[6]
port 1550 nsew signal input
rlabel metal2 s 68282 0 68338 800 6 s02_w_data[7]
port 1551 nsew signal input
rlabel metal2 s 117870 0 117926 800 6 s02_w_data[8]
port 1552 nsew signal input
rlabel metal3 s 0 6808 800 6928 6 s02_w_data[9]
port 1553 nsew signal input
rlabel metal3 s 479200 48288 480000 48408 6 s02_w_last
port 1554 nsew signal input
rlabel metal2 s 183558 0 183614 800 6 s02_w_ready
port 1555 nsew signal output
rlabel metal2 s 368386 119200 368442 120000 6 s02_w_strb[0]
port 1556 nsew signal input
rlabel metal2 s 365810 119200 365866 120000 6 s02_w_strb[1]
port 1557 nsew signal input
rlabel metal2 s 151358 119200 151414 120000 6 s02_w_strb[2]
port 1558 nsew signal input
rlabel metal2 s 206742 119200 206798 120000 6 s02_w_strb[3]
port 1559 nsew signal input
rlabel metal2 s 217046 0 217102 800 6 s02_w_user[-1]
port 1560 nsew signal input
rlabel metal3 s 0 63248 800 63368 6 s02_w_user[0]
port 1561 nsew signal input
rlabel metal2 s 128174 119200 128230 120000 6 s02_w_valid
port 1562 nsew signal input
rlabel metal2 s 444378 0 444434 800 6 test_en_i
port 1563 nsew signal input
rlabel metal4 s 4208 2128 4528 117552 6 vccd1
port 1564 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 117552 6 vccd1
port 1564 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 117552 6 vccd1
port 1564 nsew power bidirectional
rlabel metal4 s 96368 2128 96688 117552 6 vccd1
port 1564 nsew power bidirectional
rlabel metal4 s 127088 2128 127408 117552 6 vccd1
port 1564 nsew power bidirectional
rlabel metal4 s 157808 2128 158128 117552 6 vccd1
port 1564 nsew power bidirectional
rlabel metal4 s 188528 2128 188848 117552 6 vccd1
port 1564 nsew power bidirectional
rlabel metal4 s 219248 2128 219568 117552 6 vccd1
port 1564 nsew power bidirectional
rlabel metal4 s 249968 2128 250288 117552 6 vccd1
port 1564 nsew power bidirectional
rlabel metal4 s 280688 2128 281008 117552 6 vccd1
port 1564 nsew power bidirectional
rlabel metal4 s 311408 2128 311728 117552 6 vccd1
port 1564 nsew power bidirectional
rlabel metal4 s 342128 2128 342448 117552 6 vccd1
port 1564 nsew power bidirectional
rlabel metal4 s 372848 2128 373168 117552 6 vccd1
port 1564 nsew power bidirectional
rlabel metal4 s 403568 2128 403888 117552 6 vccd1
port 1564 nsew power bidirectional
rlabel metal4 s 434288 2128 434608 117552 6 vccd1
port 1564 nsew power bidirectional
rlabel metal4 s 465008 2128 465328 117552 6 vccd1
port 1564 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 117552 6 vssd1
port 1565 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 117552 6 vssd1
port 1565 nsew ground bidirectional
rlabel metal4 s 81008 2128 81328 117552 6 vssd1
port 1565 nsew ground bidirectional
rlabel metal4 s 111728 2128 112048 117552 6 vssd1
port 1565 nsew ground bidirectional
rlabel metal4 s 142448 2128 142768 117552 6 vssd1
port 1565 nsew ground bidirectional
rlabel metal4 s 173168 2128 173488 117552 6 vssd1
port 1565 nsew ground bidirectional
rlabel metal4 s 203888 2128 204208 117552 6 vssd1
port 1565 nsew ground bidirectional
rlabel metal4 s 234608 2128 234928 117552 6 vssd1
port 1565 nsew ground bidirectional
rlabel metal4 s 265328 2128 265648 117552 6 vssd1
port 1565 nsew ground bidirectional
rlabel metal4 s 296048 2128 296368 117552 6 vssd1
port 1565 nsew ground bidirectional
rlabel metal4 s 326768 2128 327088 117552 6 vssd1
port 1565 nsew ground bidirectional
rlabel metal4 s 357488 2128 357808 117552 6 vssd1
port 1565 nsew ground bidirectional
rlabel metal4 s 388208 2128 388528 117552 6 vssd1
port 1565 nsew ground bidirectional
rlabel metal4 s 418928 2128 419248 117552 6 vssd1
port 1565 nsew ground bidirectional
rlabel metal4 s 449648 2128 449968 117552 6 vssd1
port 1565 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 480000 120000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 38342260
string GDS_FILE /home/mbaykenar/Desktop/workspace/mpw7_yonga_soc/openlane/axi_node_intf_wrap/runs/22_09_05_10_40/results/signoff/axi_node_intf_wrap.magic.gds
string GDS_START 1629276
<< end >>

