magic
tech sky130B
magscale 1 2
timestamp 1649977179
use sky130_fd_pr__dfl1sd2__example_55959141808679  sky130_fd_pr__dfl1sd2__example_55959141808679_0
timestamp 1649977179
transform 1 0 100 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfl1sd2__example_55959141808679  sky130_fd_pr__dfl1sd2__example_55959141808679_1
timestamp 1649977179
transform 1 0 256 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfl1sd2__example_55959141808679  sky130_fd_pr__dfl1sd2__example_55959141808679_2
timestamp 1649977179
transform 1 0 412 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfl1sd2__example_55959141808679  sky130_fd_pr__dfl1sd2__example_55959141808679_3
timestamp 1649977179
transform 1 0 568 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfl1sd2__example_55959141808679  sky130_fd_pr__dfl1sd2__example_55959141808679_4
timestamp 1649977179
transform 1 0 724 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfl1sd2__example_55959141808679  sky130_fd_pr__dfl1sd2__example_55959141808679_5
timestamp 1649977179
transform 1 0 880 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfl1sd2__example_55959141808679  sky130_fd_pr__dfl1sd2__example_55959141808679_6
timestamp 1649977179
transform 1 0 1036 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfl1sd2__example_55959141808679  sky130_fd_pr__dfl1sd2__example_55959141808679_7
timestamp 1649977179
transform 1 0 1192 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfl1sd2__example_55959141808679  sky130_fd_pr__dfl1sd2__example_55959141808679_8
timestamp 1649977179
transform 1 0 1348 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfl1sd2__example_55959141808679  sky130_fd_pr__dfl1sd2__example_55959141808679_9
timestamp 1649977179
transform 1 0 1504 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfl1sd2__example_55959141808679  sky130_fd_pr__dfl1sd2__example_55959141808679_10
timestamp 1649977179
transform 1 0 1660 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfl1sd2__example_55959141808679  sky130_fd_pr__dfl1sd2__example_55959141808679_11
timestamp 1649977179
transform 1 0 1816 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfl1sd2__example_55959141808679  sky130_fd_pr__dfl1sd2__example_55959141808679_12
timestamp 1649977179
transform 1 0 1972 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfl1sd2__example_55959141808679  sky130_fd_pr__dfl1sd2__example_55959141808679_13
timestamp 1649977179
transform 1 0 2128 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfl1sd__example_55959141808678  sky130_fd_pr__dfl1sd__example_55959141808678_0
timestamp 1649977179
transform -1 0 0 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfl1sd__example_55959141808678  sky130_fd_pr__dfl1sd__example_55959141808678_1
timestamp 1649977179
transform 1 0 2284 0 1 0
box 0 0 1 1
<< labels >>
flabel comment s 2312 675 2312 675 0 FreeSans 300 0 0 0 D
flabel comment s 2156 675 2156 675 0 FreeSans 300 0 0 0 S
flabel comment s 2000 675 2000 675 0 FreeSans 300 0 0 0 D
flabel comment s 1844 675 1844 675 0 FreeSans 300 0 0 0 S
flabel comment s 1688 675 1688 675 0 FreeSans 300 0 0 0 D
flabel comment s 1532 675 1532 675 0 FreeSans 300 0 0 0 S
flabel comment s 1376 675 1376 675 0 FreeSans 300 0 0 0 D
flabel comment s 1220 675 1220 675 0 FreeSans 300 0 0 0 S
flabel comment s 1064 675 1064 675 0 FreeSans 300 0 0 0 D
flabel comment s 908 675 908 675 0 FreeSans 300 0 0 0 S
flabel comment s 752 675 752 675 0 FreeSans 300 0 0 0 D
flabel comment s 596 675 596 675 0 FreeSans 300 0 0 0 S
flabel comment s 440 675 440 675 0 FreeSans 300 0 0 0 D
flabel comment s 284 675 284 675 0 FreeSans 300 0 0 0 S
flabel comment s 128 675 128 675 0 FreeSans 300 0 0 0 D
flabel comment s -28 675 -28 675 0 FreeSans 300 0 0 0 S
<< properties >>
string GDS_END 11328814
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 11320668
<< end >>
