magic
tech sky130B
magscale 1 2
timestamp 1649977179
<< nwell >>
rect 0 0 466 408
<< pmos >>
rect 89 36 119 372
rect 175 36 205 372
rect 261 36 291 372
rect 347 36 377 372
<< pdiff >>
rect 36 329 89 372
rect 36 295 44 329
rect 78 295 89 329
rect 36 257 89 295
rect 36 223 44 257
rect 78 223 89 257
rect 36 185 89 223
rect 36 151 44 185
rect 78 151 89 185
rect 36 113 89 151
rect 36 79 44 113
rect 78 79 89 113
rect 36 36 89 79
rect 119 329 175 372
rect 119 295 130 329
rect 164 295 175 329
rect 119 257 175 295
rect 119 223 130 257
rect 164 223 175 257
rect 119 185 175 223
rect 119 151 130 185
rect 164 151 175 185
rect 119 113 175 151
rect 119 79 130 113
rect 164 79 175 113
rect 119 36 175 79
rect 205 329 261 372
rect 205 295 216 329
rect 250 295 261 329
rect 205 257 261 295
rect 205 223 216 257
rect 250 223 261 257
rect 205 185 261 223
rect 205 151 216 185
rect 250 151 261 185
rect 205 113 261 151
rect 205 79 216 113
rect 250 79 261 113
rect 205 36 261 79
rect 291 329 347 372
rect 291 295 302 329
rect 336 295 347 329
rect 291 257 347 295
rect 291 223 302 257
rect 336 223 347 257
rect 291 185 347 223
rect 291 151 302 185
rect 336 151 347 185
rect 291 113 347 151
rect 291 79 302 113
rect 336 79 347 113
rect 291 36 347 79
rect 377 329 430 372
rect 377 295 388 329
rect 422 295 430 329
rect 377 257 430 295
rect 377 223 388 257
rect 422 223 430 257
rect 377 185 430 223
rect 377 151 388 185
rect 422 151 430 185
rect 377 113 430 151
rect 377 79 388 113
rect 422 79 430 113
rect 377 36 430 79
<< pdiffc >>
rect 44 295 78 329
rect 44 223 78 257
rect 44 151 78 185
rect 44 79 78 113
rect 130 295 164 329
rect 130 223 164 257
rect 130 151 164 185
rect 130 79 164 113
rect 216 295 250 329
rect 216 223 250 257
rect 216 151 250 185
rect 216 79 250 113
rect 302 295 336 329
rect 302 223 336 257
rect 302 151 336 185
rect 302 79 336 113
rect 388 295 422 329
rect 388 223 422 257
rect 388 151 422 185
rect 388 79 422 113
<< poly >>
rect 89 455 377 471
rect 89 421 114 455
rect 148 421 182 455
rect 216 421 250 455
rect 284 421 318 455
rect 352 421 377 455
rect 89 398 377 421
rect 89 372 119 398
rect 175 372 205 398
rect 261 372 291 398
rect 347 372 377 398
rect 89 10 119 36
rect 175 10 205 36
rect 261 10 291 36
rect 347 10 377 36
<< polycont >>
rect 114 421 148 455
rect 182 421 216 455
rect 250 421 284 455
rect 318 421 352 455
<< locali >>
rect 98 455 368 471
rect 98 421 108 455
rect 148 421 180 455
rect 216 421 250 455
rect 286 421 318 455
rect 358 421 368 455
rect 98 403 368 421
rect 44 329 78 357
rect 44 257 78 295
rect 44 185 78 223
rect 44 113 78 151
rect 44 51 78 79
rect 130 329 164 357
rect 130 257 164 295
rect 130 185 164 223
rect 130 113 164 151
rect 130 51 164 79
rect 216 329 250 357
rect 216 257 250 295
rect 216 185 250 223
rect 216 113 250 151
rect 216 51 250 79
rect 302 329 336 357
rect 302 257 336 295
rect 302 185 336 223
rect 302 113 336 151
rect 302 51 336 79
rect 388 329 422 357
rect 388 257 422 295
rect 388 185 422 223
rect 388 113 422 151
rect 388 51 422 79
<< viali >>
rect 108 421 114 455
rect 114 421 142 455
rect 180 421 182 455
rect 182 421 214 455
rect 252 421 284 455
rect 284 421 286 455
rect 324 421 352 455
rect 352 421 358 455
rect 44 295 78 329
rect 44 223 78 257
rect 44 151 78 185
rect 44 79 78 113
rect 130 295 164 329
rect 130 223 164 257
rect 130 151 164 185
rect 130 79 164 113
rect 216 295 250 329
rect 216 223 250 257
rect 216 151 250 185
rect 216 79 250 113
rect 302 295 336 329
rect 302 223 336 257
rect 302 151 336 185
rect 302 79 336 113
rect 388 295 422 329
rect 388 223 422 257
rect 388 151 422 185
rect 388 79 422 113
<< metal1 >>
rect 96 455 370 467
rect 96 421 108 455
rect 142 421 180 455
rect 214 421 252 455
rect 286 421 324 455
rect 358 421 370 455
rect 96 409 370 421
rect 38 329 84 357
rect 38 295 44 329
rect 78 295 84 329
rect 38 257 84 295
rect 38 223 44 257
rect 78 223 84 257
rect 38 185 84 223
rect 38 151 44 185
rect 78 151 84 185
rect 38 113 84 151
rect 38 79 44 113
rect 78 79 84 113
rect 38 -29 84 79
rect 121 346 173 357
rect 121 282 173 294
rect 121 223 130 230
rect 164 223 173 230
rect 121 185 173 223
rect 121 151 130 185
rect 164 151 173 185
rect 121 113 173 151
rect 121 79 130 113
rect 164 79 173 113
rect 121 51 173 79
rect 210 329 256 357
rect 210 295 216 329
rect 250 295 256 329
rect 210 257 256 295
rect 210 223 216 257
rect 250 223 256 257
rect 210 185 256 223
rect 210 151 216 185
rect 250 151 256 185
rect 210 113 256 151
rect 210 79 216 113
rect 250 79 256 113
rect 210 -29 256 79
rect 293 346 345 357
rect 293 282 345 294
rect 293 223 302 230
rect 336 223 345 230
rect 293 185 345 223
rect 293 151 302 185
rect 336 151 345 185
rect 293 113 345 151
rect 293 79 302 113
rect 336 79 345 113
rect 293 51 345 79
rect 382 329 428 357
rect 382 295 388 329
rect 422 295 428 329
rect 382 257 428 295
rect 382 223 388 257
rect 422 223 428 257
rect 382 185 428 223
rect 382 151 388 185
rect 422 151 428 185
rect 382 113 428 151
rect 382 79 388 113
rect 422 79 428 113
rect 382 -29 428 79
rect 38 -89 428 -29
<< via1 >>
rect 121 329 173 346
rect 121 295 130 329
rect 130 295 164 329
rect 164 295 173 329
rect 121 294 173 295
rect 121 257 173 282
rect 121 230 130 257
rect 130 230 164 257
rect 164 230 173 257
rect 293 329 345 346
rect 293 295 302 329
rect 302 295 336 329
rect 336 295 345 329
rect 293 294 345 295
rect 293 257 345 282
rect 293 230 302 257
rect 302 230 336 257
rect 336 230 345 257
<< metal2 >>
rect 114 356 180 365
rect 114 300 119 356
rect 175 300 180 356
rect 114 294 121 300
rect 173 294 180 300
rect 114 282 180 294
rect 114 276 121 282
rect 173 276 180 282
rect 114 220 119 276
rect 175 220 180 276
rect 114 211 180 220
rect 286 356 352 365
rect 286 300 291 356
rect 347 300 352 356
rect 286 294 293 300
rect 345 294 352 300
rect 286 282 352 294
rect 286 276 293 282
rect 345 276 352 282
rect 286 220 291 276
rect 347 220 352 276
rect 286 211 352 220
<< via2 >>
rect 119 346 175 356
rect 119 300 121 346
rect 121 300 173 346
rect 173 300 175 346
rect 119 230 121 276
rect 121 230 173 276
rect 173 230 175 276
rect 119 220 175 230
rect 291 346 347 356
rect 291 300 293 346
rect 293 300 345 346
rect 345 300 347 346
rect 291 230 293 276
rect 293 230 345 276
rect 345 230 347 276
rect 291 220 347 230
<< metal3 >>
rect 114 356 352 365
rect 114 300 119 356
rect 175 300 291 356
rect 347 300 352 356
rect 114 299 352 300
rect 114 276 180 299
rect 114 220 119 276
rect 175 220 180 276
rect 114 211 180 220
rect 286 276 352 299
rect 286 220 291 276
rect 347 220 352 276
rect 286 211 352 220
<< labels >>
flabel metal3 s 114 299 352 365 0 FreeSans 400 0 0 0 DRAIN
port 2 nsew
flabel metal1 s 96 409 370 467 0 FreeSans 400 0 0 0 GATE
port 3 nsew
flabel metal1 s 38 -89 428 -29 0 FreeSans 400 0 0 0 SOURCE
port 4 nsew
flabel nwell s 80 399 86 406 0 FreeSans 400 0 0 0 BULK
port 1 nsew
<< properties >>
string GDS_END 9297180
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_pr/gds/sky130_fd_pr.gds
string GDS_START 9288876
string path 7.975 8.925 7.975 1.275 
<< end >>
