magic
tech sky130B
magscale 1 2
timestamp 1649977179
<< pwell >>
rect 15 163 1035 817
<< mvnmos >>
rect 241 189 341 791
rect 397 189 497 791
rect 553 189 653 791
rect 709 189 809 791
<< mvndiff >>
rect 181 779 241 791
rect 181 745 196 779
rect 230 745 241 779
rect 181 711 241 745
rect 181 677 196 711
rect 230 677 241 711
rect 181 643 241 677
rect 181 609 196 643
rect 230 609 241 643
rect 181 575 241 609
rect 181 541 196 575
rect 230 541 241 575
rect 181 507 241 541
rect 181 473 196 507
rect 230 473 241 507
rect 181 439 241 473
rect 181 405 196 439
rect 230 405 241 439
rect 181 371 241 405
rect 181 337 196 371
rect 230 337 241 371
rect 181 303 241 337
rect 181 269 196 303
rect 230 269 241 303
rect 181 235 241 269
rect 181 201 196 235
rect 230 201 241 235
rect 181 189 241 201
rect 341 779 397 791
rect 341 745 352 779
rect 386 745 397 779
rect 341 711 397 745
rect 341 677 352 711
rect 386 677 397 711
rect 341 643 397 677
rect 341 609 352 643
rect 386 609 397 643
rect 341 575 397 609
rect 341 541 352 575
rect 386 541 397 575
rect 341 507 397 541
rect 341 473 352 507
rect 386 473 397 507
rect 341 439 397 473
rect 341 405 352 439
rect 386 405 397 439
rect 341 371 397 405
rect 341 337 352 371
rect 386 337 397 371
rect 341 303 397 337
rect 341 269 352 303
rect 386 269 397 303
rect 341 235 397 269
rect 341 201 352 235
rect 386 201 397 235
rect 341 189 397 201
rect 497 779 553 791
rect 497 745 508 779
rect 542 745 553 779
rect 497 711 553 745
rect 497 677 508 711
rect 542 677 553 711
rect 497 643 553 677
rect 497 609 508 643
rect 542 609 553 643
rect 497 575 553 609
rect 497 541 508 575
rect 542 541 553 575
rect 497 507 553 541
rect 497 473 508 507
rect 542 473 553 507
rect 497 439 553 473
rect 497 405 508 439
rect 542 405 553 439
rect 497 371 553 405
rect 497 337 508 371
rect 542 337 553 371
rect 497 303 553 337
rect 497 269 508 303
rect 542 269 553 303
rect 497 235 553 269
rect 497 201 508 235
rect 542 201 553 235
rect 497 189 553 201
rect 653 779 709 791
rect 653 745 664 779
rect 698 745 709 779
rect 653 711 709 745
rect 653 677 664 711
rect 698 677 709 711
rect 653 643 709 677
rect 653 609 664 643
rect 698 609 709 643
rect 653 575 709 609
rect 653 541 664 575
rect 698 541 709 575
rect 653 507 709 541
rect 653 473 664 507
rect 698 473 709 507
rect 653 439 709 473
rect 653 405 664 439
rect 698 405 709 439
rect 653 371 709 405
rect 653 337 664 371
rect 698 337 709 371
rect 653 303 709 337
rect 653 269 664 303
rect 698 269 709 303
rect 653 235 709 269
rect 653 201 664 235
rect 698 201 709 235
rect 653 189 709 201
rect 809 779 869 791
rect 809 745 820 779
rect 854 745 869 779
rect 809 711 869 745
rect 809 677 820 711
rect 854 677 869 711
rect 809 643 869 677
rect 809 609 820 643
rect 854 609 869 643
rect 809 575 869 609
rect 809 541 820 575
rect 854 541 869 575
rect 809 507 869 541
rect 809 473 820 507
rect 854 473 869 507
rect 809 439 869 473
rect 809 405 820 439
rect 854 405 869 439
rect 809 371 869 405
rect 809 337 820 371
rect 854 337 869 371
rect 809 303 869 337
rect 809 269 820 303
rect 854 269 869 303
rect 809 235 869 269
rect 809 201 820 235
rect 854 201 869 235
rect 809 189 869 201
<< mvndiffc >>
rect 196 745 230 779
rect 196 677 230 711
rect 196 609 230 643
rect 196 541 230 575
rect 196 473 230 507
rect 196 405 230 439
rect 196 337 230 371
rect 196 269 230 303
rect 196 201 230 235
rect 352 745 386 779
rect 352 677 386 711
rect 352 609 386 643
rect 352 541 386 575
rect 352 473 386 507
rect 352 405 386 439
rect 352 337 386 371
rect 352 269 386 303
rect 352 201 386 235
rect 508 745 542 779
rect 508 677 542 711
rect 508 609 542 643
rect 508 541 542 575
rect 508 473 542 507
rect 508 405 542 439
rect 508 337 542 371
rect 508 269 542 303
rect 508 201 542 235
rect 664 745 698 779
rect 664 677 698 711
rect 664 609 698 643
rect 664 541 698 575
rect 664 473 698 507
rect 664 405 698 439
rect 664 337 698 371
rect 664 269 698 303
rect 664 201 698 235
rect 820 745 854 779
rect 820 677 854 711
rect 820 609 854 643
rect 820 541 854 575
rect 820 473 854 507
rect 820 405 854 439
rect 820 337 854 371
rect 820 269 854 303
rect 820 201 854 235
<< mvpsubdiff >>
rect 41 779 181 791
rect 41 201 60 779
rect 162 201 181 779
rect 41 189 181 201
rect 869 779 1009 791
rect 869 201 888 779
rect 990 201 1009 779
rect 869 189 1009 201
<< mvpsubdiffcont >>
rect 60 201 162 779
rect 888 201 990 779
<< poly >>
rect 383 959 667 980
rect 190 867 341 883
rect 190 833 206 867
rect 240 833 341 867
rect 383 857 406 959
rect 644 857 667 959
rect 383 841 667 857
rect 709 867 860 883
rect 190 817 341 833
rect 241 791 341 817
rect 397 791 497 841
rect 553 791 653 841
rect 709 833 810 867
rect 844 833 860 867
rect 709 817 860 833
rect 709 791 809 817
rect 241 163 341 189
rect 190 147 341 163
rect 190 113 206 147
rect 240 113 341 147
rect 397 139 497 189
rect 553 139 653 189
rect 709 163 809 189
rect 709 147 860 163
rect 190 97 341 113
rect 383 123 667 139
rect 383 21 406 123
rect 644 21 667 123
rect 709 113 810 147
rect 844 113 860 147
rect 709 97 860 113
rect 383 0 667 21
<< polycont >>
rect 206 833 240 867
rect 406 857 644 959
rect 810 833 844 867
rect 206 113 240 147
rect 406 21 644 123
rect 810 113 844 147
<< locali >>
rect 383 961 667 980
rect 190 867 256 883
rect 190 833 206 867
rect 240 833 256 867
rect 383 855 400 961
rect 650 855 667 961
rect 383 843 667 855
rect 794 867 860 883
rect 190 817 256 833
rect 794 833 810 867
rect 844 833 860 867
rect 794 817 860 833
rect 190 795 230 817
rect 820 795 860 817
rect 41 779 230 795
rect 41 201 60 779
rect 162 745 196 779
rect 162 711 230 745
rect 162 677 196 711
rect 162 643 230 677
rect 162 609 196 643
rect 162 575 230 609
rect 162 541 196 575
rect 162 507 230 541
rect 162 473 196 507
rect 162 439 230 473
rect 162 405 196 439
rect 162 371 230 405
rect 162 337 196 371
rect 162 303 230 337
rect 162 269 196 303
rect 162 235 230 269
rect 162 201 196 235
rect 41 185 230 201
rect 352 779 386 795
rect 352 711 386 725
rect 352 643 386 653
rect 352 575 386 581
rect 352 507 386 509
rect 352 471 386 473
rect 352 399 386 405
rect 352 327 386 337
rect 352 255 386 269
rect 352 185 386 201
rect 508 779 542 795
rect 508 711 542 725
rect 508 643 542 653
rect 508 575 542 581
rect 508 507 542 509
rect 508 471 542 473
rect 508 399 542 405
rect 508 327 542 337
rect 508 255 542 269
rect 508 185 542 201
rect 664 779 698 795
rect 664 711 698 725
rect 664 643 698 653
rect 664 575 698 581
rect 664 507 698 509
rect 664 471 698 473
rect 664 399 698 405
rect 664 327 698 337
rect 664 255 698 269
rect 664 185 698 201
rect 820 779 1009 795
rect 854 745 888 779
rect 820 711 888 745
rect 854 677 888 711
rect 820 643 888 677
rect 854 609 888 643
rect 820 575 888 609
rect 854 541 888 575
rect 820 507 888 541
rect 854 473 888 507
rect 820 439 888 473
rect 854 405 888 439
rect 820 371 888 405
rect 854 337 888 371
rect 820 303 888 337
rect 854 269 888 303
rect 820 235 888 269
rect 854 201 888 235
rect 990 201 1009 779
rect 820 185 1009 201
rect 190 163 230 185
rect 820 163 860 185
rect 190 147 256 163
rect 190 113 206 147
rect 240 113 256 147
rect 794 147 860 163
rect 190 97 256 113
rect 383 125 667 137
rect 383 19 400 125
rect 650 19 667 125
rect 794 113 810 147
rect 844 113 860 147
rect 794 97 860 113
rect 383 0 667 19
<< viali >>
rect 400 959 650 961
rect 400 857 406 959
rect 406 857 644 959
rect 644 857 650 959
rect 400 855 650 857
rect 60 725 94 759
rect 60 653 94 687
rect 60 581 94 615
rect 60 509 94 543
rect 60 437 94 471
rect 60 365 94 399
rect 60 293 94 327
rect 60 221 94 255
rect 352 745 386 759
rect 352 725 386 745
rect 352 677 386 687
rect 352 653 386 677
rect 352 609 386 615
rect 352 581 386 609
rect 352 541 386 543
rect 352 509 386 541
rect 352 439 386 471
rect 352 437 386 439
rect 352 371 386 399
rect 352 365 386 371
rect 352 303 386 327
rect 352 293 386 303
rect 352 235 386 255
rect 352 221 386 235
rect 508 745 542 759
rect 508 725 542 745
rect 508 677 542 687
rect 508 653 542 677
rect 508 609 542 615
rect 508 581 542 609
rect 508 541 542 543
rect 508 509 542 541
rect 508 439 542 471
rect 508 437 542 439
rect 508 371 542 399
rect 508 365 542 371
rect 508 303 542 327
rect 508 293 542 303
rect 508 235 542 255
rect 508 221 542 235
rect 664 745 698 759
rect 664 725 698 745
rect 664 677 698 687
rect 664 653 698 677
rect 664 609 698 615
rect 664 581 698 609
rect 664 541 698 543
rect 664 509 698 541
rect 664 439 698 471
rect 664 437 698 439
rect 664 371 698 399
rect 664 365 698 371
rect 664 303 698 327
rect 664 293 698 303
rect 664 235 698 255
rect 664 221 698 235
rect 956 725 990 759
rect 956 653 990 687
rect 956 581 990 615
rect 956 509 990 543
rect 956 437 990 471
rect 956 365 990 399
rect 956 293 990 327
rect 956 221 990 255
rect 400 123 650 125
rect 400 21 406 123
rect 406 21 644 123
rect 644 21 650 123
rect 400 19 650 21
<< metal1 >>
rect 380 961 670 980
rect 380 855 400 961
rect 650 855 670 961
rect 380 843 670 855
rect 41 759 100 771
rect 41 725 60 759
rect 94 725 100 759
rect 41 687 100 725
rect 41 653 60 687
rect 94 653 100 687
rect 41 615 100 653
rect 41 581 60 615
rect 94 581 100 615
rect 41 543 100 581
rect 41 509 60 543
rect 94 509 100 543
rect 41 471 100 509
rect 41 437 60 471
rect 94 437 100 471
rect 41 399 100 437
rect 41 365 60 399
rect 94 365 100 399
rect 41 327 100 365
rect 41 293 60 327
rect 94 293 100 327
rect 41 255 100 293
rect 41 221 60 255
rect 94 221 100 255
rect 41 209 100 221
rect 343 759 395 771
rect 343 725 352 759
rect 386 725 395 759
rect 343 687 395 725
rect 343 653 352 687
rect 386 653 395 687
rect 343 615 395 653
rect 343 581 352 615
rect 386 581 395 615
rect 343 543 395 581
rect 343 509 352 543
rect 386 509 395 543
rect 343 471 395 509
rect 343 459 352 471
rect 386 459 395 471
rect 343 399 395 407
rect 343 395 352 399
rect 386 395 395 399
rect 343 331 395 343
rect 343 267 395 279
rect 343 209 395 215
rect 499 765 551 771
rect 499 701 551 713
rect 499 637 551 649
rect 499 581 508 585
rect 542 581 551 585
rect 499 573 551 581
rect 499 509 508 521
rect 542 509 551 521
rect 499 471 551 509
rect 499 437 508 471
rect 542 437 551 471
rect 499 399 551 437
rect 499 365 508 399
rect 542 365 551 399
rect 499 327 551 365
rect 499 293 508 327
rect 542 293 551 327
rect 499 255 551 293
rect 499 221 508 255
rect 542 221 551 255
rect 499 209 551 221
rect 655 759 707 771
rect 655 725 664 759
rect 698 725 707 759
rect 655 687 707 725
rect 655 653 664 687
rect 698 653 707 687
rect 655 615 707 653
rect 655 581 664 615
rect 698 581 707 615
rect 655 543 707 581
rect 655 509 664 543
rect 698 509 707 543
rect 655 471 707 509
rect 655 459 664 471
rect 698 459 707 471
rect 655 399 707 407
rect 655 395 664 399
rect 698 395 707 399
rect 655 331 707 343
rect 655 267 707 279
rect 655 209 707 215
rect 950 759 1009 771
rect 950 725 956 759
rect 990 725 1009 759
rect 950 687 1009 725
rect 950 653 956 687
rect 990 653 1009 687
rect 950 615 1009 653
rect 950 581 956 615
rect 990 581 1009 615
rect 950 543 1009 581
rect 950 509 956 543
rect 990 509 1009 543
rect 950 471 1009 509
rect 950 437 956 471
rect 990 437 1009 471
rect 950 399 1009 437
rect 950 365 956 399
rect 990 365 1009 399
rect 950 327 1009 365
rect 950 293 956 327
rect 990 293 1009 327
rect 950 255 1009 293
rect 950 221 956 255
rect 990 221 1009 255
rect 950 209 1009 221
rect 380 125 670 137
rect 380 19 400 125
rect 650 19 670 125
rect 380 0 670 19
<< via1 >>
rect 343 437 352 459
rect 352 437 386 459
rect 386 437 395 459
rect 343 407 395 437
rect 343 365 352 395
rect 352 365 386 395
rect 386 365 395 395
rect 343 343 395 365
rect 343 327 395 331
rect 343 293 352 327
rect 352 293 386 327
rect 386 293 395 327
rect 343 279 395 293
rect 343 255 395 267
rect 343 221 352 255
rect 352 221 386 255
rect 386 221 395 255
rect 343 215 395 221
rect 499 759 551 765
rect 499 725 508 759
rect 508 725 542 759
rect 542 725 551 759
rect 499 713 551 725
rect 499 687 551 701
rect 499 653 508 687
rect 508 653 542 687
rect 542 653 551 687
rect 499 649 551 653
rect 499 615 551 637
rect 499 585 508 615
rect 508 585 542 615
rect 542 585 551 615
rect 499 543 551 573
rect 499 521 508 543
rect 508 521 542 543
rect 542 521 551 543
rect 655 437 664 459
rect 664 437 698 459
rect 698 437 707 459
rect 655 407 707 437
rect 655 365 664 395
rect 664 365 698 395
rect 698 365 707 395
rect 655 343 707 365
rect 655 327 707 331
rect 655 293 664 327
rect 664 293 698 327
rect 698 293 707 327
rect 655 279 707 293
rect 655 255 707 267
rect 655 221 664 255
rect 664 221 698 255
rect 698 221 707 255
rect 655 215 707 221
<< metal2 >>
rect 14 765 1036 771
rect 14 713 499 765
rect 551 713 1036 765
rect 14 701 1036 713
rect 14 649 499 701
rect 551 649 1036 701
rect 14 637 1036 649
rect 14 585 499 637
rect 551 585 1036 637
rect 14 573 1036 585
rect 14 521 499 573
rect 551 521 1036 573
rect 14 515 1036 521
rect 14 459 1036 465
rect 14 407 343 459
rect 395 407 655 459
rect 707 407 1036 459
rect 14 395 1036 407
rect 14 343 343 395
rect 395 343 655 395
rect 707 343 1036 395
rect 14 331 1036 343
rect 14 279 343 331
rect 395 279 655 331
rect 707 279 1036 331
rect 14 267 1036 279
rect 14 215 343 267
rect 395 215 655 267
rect 707 215 1036 267
rect 14 209 1036 215
<< labels >>
flabel metal2 s 36 313 66 417 0 FreeSans 400 90 0 0 SOURCE
port 3 nsew
flabel metal2 s 35 602 70 699 0 FreeSans 400 270 0 0 DRAIN
port 1 nsew
flabel metal1 s 470 85 568 119 0 FreeSans 200 0 0 0 GATE
port 2 nsew
flabel metal1 s 470 855 568 889 0 FreeSans 400 0 0 0 GATE
port 2 nsew
flabel metal1 s 41 466 100 496 0 FreeSans 200 90 0 0 SUBSTRATE
port 4 nsew
flabel metal1 s 950 469 1009 499 0 FreeSans 200 90 0 0 SUBSTRATE
port 4 nsew
flabel comment s 369 490 369 490 0 FreeSans 300 0 0 0 S
flabel comment s 525 490 525 490 0 FreeSans 300 0 0 0 S
flabel comment s 681 490 681 490 0 FreeSans 300 0 0 0 S
flabel comment s 369 490 369 490 0 FreeSans 300 0 0 0 S
flabel comment s 525 490 525 490 0 FreeSans 300 0 0 0 D
flabel comment s 681 490 681 490 0 FreeSans 300 0 0 0 S
flabel comment s 757 462 757 462 0 FreeSans 400 90 0 0 dummy_poly
flabel comment s 287 473 287 473 0 FreeSans 400 90 0 0 dummy_poly
<< properties >>
string GDS_END 8481320
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_pr/gds/sky130_fd_pr.gds
string GDS_START 8464596
<< end >>
