magic
tech sky130A
magscale 1 2
timestamp 1649977179
<< nwell >>
rect -66 377 1122 897
<< pwell >>
rect 4 43 914 283
rect -26 -43 1082 43
<< mvnmos >>
rect 87 107 187 257
rect 254 107 354 257
rect 410 107 510 257
rect 575 107 675 257
rect 731 107 831 257
<< mvpmos >>
rect 87 443 187 743
rect 433 443 533 743
rect 575 443 675 743
rect 731 443 831 743
rect 873 443 973 743
<< mvndiff >>
rect 30 249 87 257
rect 30 215 42 249
rect 76 215 87 249
rect 30 149 87 215
rect 30 115 42 149
rect 76 115 87 149
rect 30 107 87 115
rect 187 249 254 257
rect 187 215 198 249
rect 232 215 254 249
rect 187 149 254 215
rect 187 115 198 149
rect 232 115 254 149
rect 187 107 254 115
rect 354 161 410 257
rect 354 127 365 161
rect 399 127 410 161
rect 354 107 410 127
rect 510 183 575 257
rect 510 149 521 183
rect 555 149 575 183
rect 510 107 575 149
rect 675 177 731 257
rect 675 143 686 177
rect 720 143 731 177
rect 675 107 731 143
rect 831 179 888 257
rect 831 145 842 179
rect 876 145 888 179
rect 831 107 888 145
<< mvpdiff >>
rect 30 735 87 743
rect 30 701 42 735
rect 76 701 87 735
rect 30 652 87 701
rect 30 618 42 652
rect 76 618 87 652
rect 30 568 87 618
rect 30 534 42 568
rect 76 534 87 568
rect 30 485 87 534
rect 30 451 42 485
rect 76 451 87 485
rect 30 443 87 451
rect 187 735 433 743
rect 187 701 198 735
rect 232 701 433 735
rect 187 649 433 701
rect 187 615 198 649
rect 232 615 433 649
rect 187 564 433 615
rect 187 530 198 564
rect 232 530 433 564
rect 187 443 433 530
rect 533 443 575 743
rect 675 735 731 743
rect 675 701 686 735
rect 720 701 731 735
rect 675 652 731 701
rect 675 618 686 652
rect 720 618 731 652
rect 675 568 731 618
rect 675 534 686 568
rect 720 534 731 568
rect 675 485 731 534
rect 675 451 686 485
rect 720 451 731 485
rect 675 443 731 451
rect 831 443 873 743
rect 973 731 1026 743
rect 973 697 984 731
rect 1018 697 1026 731
rect 973 651 1026 697
rect 973 617 984 651
rect 1018 617 1026 651
rect 973 569 1026 617
rect 973 535 984 569
rect 1018 535 1026 569
rect 973 489 1026 535
rect 973 455 984 489
rect 1018 455 1026 489
rect 973 443 1026 455
<< mvndiffc >>
rect 42 215 76 249
rect 42 115 76 149
rect 198 215 232 249
rect 198 115 232 149
rect 365 127 399 161
rect 521 149 555 183
rect 686 143 720 177
rect 842 145 876 179
<< mvpdiffc >>
rect 42 701 76 735
rect 42 618 76 652
rect 42 534 76 568
rect 42 451 76 485
rect 198 701 232 735
rect 198 615 232 649
rect 198 530 232 564
rect 686 701 720 735
rect 686 618 720 652
rect 686 534 720 568
rect 686 451 720 485
rect 984 697 1018 731
rect 984 617 1018 651
rect 984 535 1018 569
rect 984 455 1018 489
<< mvpsubdiff >>
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1056 17
<< mvnsubdiff >>
rect 0 797 31 831
rect 65 797 127 831
rect 161 797 223 831
rect 257 797 319 831
rect 353 797 415 831
rect 449 797 511 831
rect 545 797 607 831
rect 641 797 703 831
rect 737 797 799 831
rect 833 797 895 831
rect 929 797 991 831
rect 1025 797 1056 831
<< mvpsubdiffcont >>
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
<< mvnsubdiffcont >>
rect 31 797 65 831
rect 127 797 161 831
rect 223 797 257 831
rect 319 797 353 831
rect 415 797 449 831
rect 511 797 545 831
rect 607 797 641 831
rect 703 797 737 831
rect 799 797 833 831
rect 895 797 929 831
rect 991 797 1025 831
<< poly >>
rect 87 743 187 769
rect 433 743 533 769
rect 575 743 675 769
rect 731 743 831 769
rect 873 743 973 769
rect 87 335 187 443
rect 433 417 533 443
rect 87 301 133 335
rect 167 301 187 335
rect 87 257 187 301
rect 254 395 354 415
rect 254 361 300 395
rect 334 361 354 395
rect 254 257 354 361
rect 410 395 533 417
rect 410 361 482 395
rect 516 361 533 395
rect 410 283 533 361
rect 575 366 675 443
rect 575 332 603 366
rect 637 332 675 366
rect 410 257 510 283
rect 575 257 675 332
rect 731 366 831 443
rect 731 332 751 366
rect 785 332 831 366
rect 731 257 831 332
rect 873 417 973 443
rect 873 394 980 417
rect 873 360 926 394
rect 960 360 980 394
rect 873 326 980 360
rect 873 292 926 326
rect 960 292 980 326
rect 873 272 980 292
rect 87 81 187 107
rect 254 81 354 107
rect 410 81 510 107
rect 575 81 675 107
rect 731 81 831 107
<< polycont >>
rect 133 301 167 335
rect 300 361 334 395
rect 482 361 516 395
rect 603 332 637 366
rect 751 332 785 366
rect 926 360 960 394
rect 926 292 960 326
<< locali >>
rect 0 797 31 831
rect 65 797 127 831
rect 161 797 223 831
rect 257 797 319 831
rect 353 797 415 831
rect 449 797 511 831
rect 545 797 607 831
rect 641 797 703 831
rect 737 797 799 831
rect 833 797 895 831
rect 929 797 991 831
rect 1025 797 1056 831
rect 25 735 76 751
rect 25 701 42 735
rect 25 652 76 701
rect 25 618 42 652
rect 25 568 76 618
rect 25 534 42 568
rect 25 485 76 534
rect 112 735 650 751
rect 146 701 184 735
rect 232 701 256 735
rect 290 701 328 735
rect 362 701 400 735
rect 434 701 472 735
rect 506 701 544 735
rect 578 701 616 735
rect 112 649 650 701
rect 112 615 198 649
rect 232 615 650 649
rect 112 564 650 615
rect 112 530 198 564
rect 232 530 650 564
rect 686 735 736 751
rect 720 701 736 735
rect 686 652 736 701
rect 720 618 736 652
rect 686 568 736 618
rect 720 534 736 568
rect 686 494 736 534
rect 25 451 42 485
rect 25 249 76 451
rect 117 485 736 494
rect 117 460 686 485
rect 117 335 183 460
rect 720 451 736 485
rect 686 435 736 451
rect 772 735 1034 747
rect 772 701 778 735
rect 812 701 850 735
rect 884 701 922 735
rect 956 731 994 735
rect 956 701 984 731
rect 1028 701 1034 735
rect 772 697 984 701
rect 1018 697 1034 701
rect 772 651 1034 697
rect 772 617 984 651
rect 1018 617 1034 651
rect 772 569 1034 617
rect 772 535 984 569
rect 1018 535 1034 569
rect 772 489 1034 535
rect 772 455 984 489
rect 1018 455 1034 489
rect 772 439 1034 455
rect 284 395 430 411
rect 284 361 300 395
rect 334 361 430 395
rect 284 355 430 361
rect 117 301 133 335
rect 167 319 183 335
rect 167 301 360 319
rect 117 285 360 301
rect 25 215 42 249
rect 25 149 76 215
rect 25 115 42 149
rect 25 99 76 115
rect 112 215 198 249
rect 232 215 290 249
rect 112 149 290 215
rect 326 244 360 285
rect 396 314 430 355
rect 466 395 551 424
rect 466 361 482 395
rect 516 361 551 395
rect 466 350 551 361
rect 591 366 650 424
rect 910 394 976 403
rect 591 332 603 366
rect 637 332 650 366
rect 591 316 650 332
rect 697 366 839 382
rect 697 332 751 366
rect 785 332 839 366
rect 697 316 839 332
rect 910 360 926 394
rect 960 360 976 394
rect 910 326 976 360
rect 396 280 555 314
rect 910 292 926 326
rect 960 292 976 326
rect 910 280 976 292
rect 521 246 976 280
rect 326 210 485 244
rect 607 242 742 246
rect 451 183 571 210
rect 451 176 521 183
rect 112 115 198 149
rect 232 115 290 149
rect 112 113 290 115
rect 146 79 184 113
rect 218 79 256 113
rect 112 73 290 79
rect 349 161 415 174
rect 349 127 365 161
rect 399 127 415 161
rect 349 87 415 127
rect 505 149 521 176
rect 555 149 571 183
rect 505 123 571 149
rect 670 177 736 206
rect 670 143 686 177
rect 720 143 736 177
rect 670 87 736 143
rect 349 53 736 87
rect 778 179 1038 210
rect 778 145 842 179
rect 876 145 1038 179
rect 778 113 1038 145
rect 778 79 783 113
rect 817 79 855 113
rect 889 79 927 113
rect 961 79 999 113
rect 1033 79 1038 113
rect 778 73 1038 79
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1056 17
<< viali >>
rect 31 797 65 831
rect 127 797 161 831
rect 223 797 257 831
rect 319 797 353 831
rect 415 797 449 831
rect 511 797 545 831
rect 607 797 641 831
rect 703 797 737 831
rect 799 797 833 831
rect 895 797 929 831
rect 991 797 1025 831
rect 112 701 146 735
rect 184 701 198 735
rect 198 701 218 735
rect 256 701 290 735
rect 328 701 362 735
rect 400 701 434 735
rect 472 701 506 735
rect 544 701 578 735
rect 616 701 650 735
rect 778 701 812 735
rect 850 701 884 735
rect 922 701 956 735
rect 994 731 1028 735
rect 994 701 1018 731
rect 1018 701 1028 731
rect 112 79 146 113
rect 184 79 218 113
rect 256 79 290 113
rect 783 79 817 113
rect 855 79 889 113
rect 927 79 961 113
rect 999 79 1033 113
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
<< metal1 >>
rect 0 831 1056 837
rect 0 797 31 831
rect 65 797 127 831
rect 161 797 223 831
rect 257 797 319 831
rect 353 797 415 831
rect 449 797 511 831
rect 545 797 607 831
rect 641 797 703 831
rect 737 797 799 831
rect 833 797 895 831
rect 929 797 991 831
rect 1025 797 1056 831
rect 0 791 1056 797
rect 0 735 1056 763
rect 0 701 112 735
rect 146 701 184 735
rect 218 701 256 735
rect 290 701 328 735
rect 362 701 400 735
rect 434 701 472 735
rect 506 701 544 735
rect 578 701 616 735
rect 650 701 778 735
rect 812 701 850 735
rect 884 701 922 735
rect 956 701 994 735
rect 1028 701 1056 735
rect 0 689 1056 701
rect 0 113 1056 125
rect 0 79 112 113
rect 146 79 184 113
rect 218 79 256 113
rect 290 79 783 113
rect 817 79 855 113
rect 889 79 927 113
rect 961 79 999 113
rect 1033 79 1056 113
rect 0 51 1056 79
rect 0 17 1056 23
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1056 17
rect 0 -23 1056 -17
<< labels >>
rlabel comment s 0 0 0 0 4 o22a_1
flabel metal1 s 0 51 1056 125 0 FreeSans 340 0 0 0 VGND
port 5 nsew ground bidirectional
flabel metal1 s 0 0 1056 23 0 FreeSans 340 0 0 0 VNB
port 6 nsew ground bidirectional
flabel metal1 s 0 689 1056 763 0 FreeSans 340 0 0 0 VPWR
port 8 nsew power bidirectional
flabel metal1 s 0 791 1056 814 0 FreeSans 340 0 0 0 VPB
port 7 nsew power bidirectional
flabel locali s 607 242 641 276 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 703 242 737 276 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 703 316 737 350 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 799 316 833 350 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 511 390 545 424 0 FreeSans 340 0 0 0 B1
port 3 nsew signal input
flabel locali s 607 316 641 350 0 FreeSans 340 0 0 0 B2
port 4 nsew signal input
flabel locali s 607 390 641 424 0 FreeSans 340 0 0 0 B2
port 4 nsew signal input
flabel locali s 31 168 65 202 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
flabel locali s 31 242 65 276 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
flabel locali s 31 316 65 350 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
flabel locali s 31 390 65 424 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
flabel locali s 31 464 65 498 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
flabel locali s 31 538 65 572 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
flabel locali s 31 612 65 646 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 1056 814
string GDS_END 398928
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hvl/gds/sky130_fd_sc_hvl.gds
string GDS_START 386192
string LEFclass CORE
string LEFsite unithv
string LEFsymmetry X Y
<< end >>
