magic
tech sky130B
magscale 12 1
timestamp 1598774805
<< metal5 >>
rect 0 0 60 15
<< properties >>
string FIXED_BBOX 0 -30 75 105
<< end >>
