magic
tech sky130A
magscale 1 2
timestamp 1649977179
<< nwell >>
rect -66 377 3042 897
<< pwell >>
rect 2714 283 2972 303
rect 1784 217 2050 283
rect 2448 217 2972 283
rect 7 43 2972 217
rect -26 -43 3002 43
<< mvnmos >>
rect 86 107 186 191
rect 242 107 342 191
rect 384 107 484 191
rect 540 107 640 191
rect 682 107 782 191
rect 838 107 938 191
rect 1104 107 1204 191
rect 1390 107 1490 191
rect 1546 107 1646 191
rect 1688 107 1788 191
rect 1867 107 1967 257
rect 2046 107 2146 191
rect 2210 107 2310 191
rect 2352 107 2452 191
rect 2527 107 2627 257
rect 2793 127 2893 277
<< mvpmos >>
rect 87 593 187 677
rect 243 593 343 677
rect 385 593 485 677
rect 541 593 641 677
rect 683 593 783 677
rect 858 593 958 743
rect 1124 593 1224 743
rect 1390 543 1490 627
rect 1546 543 1646 627
rect 1688 543 1788 627
rect 1867 543 1967 743
rect 2023 543 2123 743
rect 2202 543 2302 627
rect 2352 543 2452 627
rect 2527 543 2627 743
rect 2793 443 2893 743
<< mvndiff >>
rect 1810 191 1867 257
rect 33 166 86 191
rect 33 132 41 166
rect 75 132 86 166
rect 33 107 86 132
rect 186 166 242 191
rect 186 132 197 166
rect 231 132 242 166
rect 186 107 242 132
rect 342 107 384 191
rect 484 166 540 191
rect 484 132 495 166
rect 529 132 540 166
rect 484 107 540 132
rect 640 107 682 191
rect 782 166 838 191
rect 782 132 793 166
rect 827 132 838 166
rect 782 107 838 132
rect 938 166 991 191
rect 938 132 949 166
rect 983 132 991 166
rect 938 107 991 132
rect 1051 166 1104 191
rect 1051 132 1059 166
rect 1093 132 1104 166
rect 1051 107 1104 132
rect 1204 166 1257 191
rect 1204 132 1215 166
rect 1249 132 1257 166
rect 1204 107 1257 132
rect 1317 170 1390 191
rect 1317 136 1329 170
rect 1363 136 1390 170
rect 1317 107 1390 136
rect 1490 170 1546 191
rect 1490 136 1501 170
rect 1535 136 1546 170
rect 1490 107 1546 136
rect 1646 107 1688 191
rect 1788 182 1867 191
rect 1788 148 1822 182
rect 1856 148 1867 182
rect 1788 107 1867 148
rect 1967 191 2024 257
rect 2740 265 2793 277
rect 2474 245 2527 257
rect 2474 211 2482 245
rect 2516 211 2527 245
rect 2474 191 2527 211
rect 1967 182 2046 191
rect 1967 148 1978 182
rect 2012 148 2046 182
rect 1967 107 2046 148
rect 2146 166 2210 191
rect 2146 132 2165 166
rect 2199 132 2210 166
rect 2146 107 2210 132
rect 2310 107 2352 191
rect 2452 153 2527 191
rect 2452 119 2482 153
rect 2516 119 2527 153
rect 2452 107 2527 119
rect 2627 245 2680 257
rect 2627 211 2638 245
rect 2672 211 2680 245
rect 2627 153 2680 211
rect 2627 119 2638 153
rect 2672 119 2680 153
rect 2740 231 2748 265
rect 2782 231 2793 265
rect 2740 173 2793 231
rect 2740 139 2748 173
rect 2782 139 2793 173
rect 2740 127 2793 139
rect 2893 265 2946 277
rect 2893 231 2904 265
rect 2938 231 2946 265
rect 2893 173 2946 231
rect 2893 139 2904 173
rect 2938 139 2946 173
rect 2893 127 2946 139
rect 2627 107 2680 119
<< mvpdiff >>
rect 805 731 858 743
rect 805 697 813 731
rect 847 697 858 731
rect 805 677 858 697
rect 30 652 87 677
rect 30 618 42 652
rect 76 618 87 652
rect 30 593 87 618
rect 187 652 243 677
rect 187 618 198 652
rect 232 618 243 652
rect 187 593 243 618
rect 343 593 385 677
rect 485 652 541 677
rect 485 618 496 652
rect 530 618 541 652
rect 485 593 541 618
rect 641 593 683 677
rect 783 639 858 677
rect 783 605 813 639
rect 847 605 858 639
rect 783 593 858 605
rect 958 731 1011 743
rect 958 697 969 731
rect 1003 697 1011 731
rect 958 639 1011 697
rect 958 605 969 639
rect 1003 605 1011 639
rect 958 593 1011 605
rect 1071 731 1124 743
rect 1071 697 1079 731
rect 1113 697 1124 731
rect 1071 639 1124 697
rect 1071 605 1079 639
rect 1113 605 1124 639
rect 1071 593 1124 605
rect 1224 731 1277 743
rect 1224 697 1235 731
rect 1269 697 1277 731
rect 1224 639 1277 697
rect 1810 735 1867 743
rect 1810 701 1822 735
rect 1856 701 1867 735
rect 1224 605 1235 639
rect 1269 605 1277 639
rect 1810 627 1867 701
rect 1224 593 1277 605
rect 1337 602 1390 627
rect 1337 568 1345 602
rect 1379 568 1390 602
rect 1337 543 1390 568
rect 1490 602 1546 627
rect 1490 568 1501 602
rect 1535 568 1546 602
rect 1490 543 1546 568
rect 1646 543 1688 627
rect 1788 543 1867 627
rect 1967 590 2023 743
rect 1967 556 1978 590
rect 2012 556 2023 590
rect 1967 543 2023 556
rect 2123 627 2180 743
rect 2474 731 2527 743
rect 2474 697 2482 731
rect 2516 697 2527 731
rect 2474 660 2527 697
rect 2474 627 2482 660
rect 2123 599 2202 627
rect 2123 565 2134 599
rect 2168 565 2202 599
rect 2123 543 2202 565
rect 2302 543 2352 627
rect 2452 626 2482 627
rect 2516 626 2527 660
rect 2452 589 2527 626
rect 2452 555 2482 589
rect 2516 555 2527 589
rect 2452 543 2527 555
rect 2627 731 2680 743
rect 2627 697 2638 731
rect 2672 697 2680 731
rect 2627 660 2680 697
rect 2627 626 2638 660
rect 2672 626 2680 660
rect 2627 589 2680 626
rect 2627 555 2638 589
rect 2672 555 2680 589
rect 2627 543 2680 555
rect 2740 731 2793 743
rect 2740 697 2748 731
rect 2782 697 2793 731
rect 2740 651 2793 697
rect 2740 617 2748 651
rect 2782 617 2793 651
rect 2740 569 2793 617
rect 2740 535 2748 569
rect 2782 535 2793 569
rect 2740 489 2793 535
rect 2740 455 2748 489
rect 2782 455 2793 489
rect 2740 443 2793 455
rect 2893 731 2946 743
rect 2893 697 2904 731
rect 2938 697 2946 731
rect 2893 651 2946 697
rect 2893 617 2904 651
rect 2938 617 2946 651
rect 2893 569 2946 617
rect 2893 535 2904 569
rect 2938 535 2946 569
rect 2893 489 2946 535
rect 2893 455 2904 489
rect 2938 455 2946 489
rect 2893 443 2946 455
<< mvndiffc >>
rect 41 132 75 166
rect 197 132 231 166
rect 495 132 529 166
rect 793 132 827 166
rect 949 132 983 166
rect 1059 132 1093 166
rect 1215 132 1249 166
rect 1329 136 1363 170
rect 1501 136 1535 170
rect 1822 148 1856 182
rect 2482 211 2516 245
rect 1978 148 2012 182
rect 2165 132 2199 166
rect 2482 119 2516 153
rect 2638 211 2672 245
rect 2638 119 2672 153
rect 2748 231 2782 265
rect 2748 139 2782 173
rect 2904 231 2938 265
rect 2904 139 2938 173
<< mvpdiffc >>
rect 813 697 847 731
rect 42 618 76 652
rect 198 618 232 652
rect 496 618 530 652
rect 813 605 847 639
rect 969 697 1003 731
rect 969 605 1003 639
rect 1079 697 1113 731
rect 1079 605 1113 639
rect 1235 697 1269 731
rect 1822 701 1856 735
rect 1235 605 1269 639
rect 1345 568 1379 602
rect 1501 568 1535 602
rect 1978 556 2012 590
rect 2482 697 2516 731
rect 2134 565 2168 599
rect 2482 626 2516 660
rect 2482 555 2516 589
rect 2638 697 2672 731
rect 2638 626 2672 660
rect 2638 555 2672 589
rect 2748 697 2782 731
rect 2748 617 2782 651
rect 2748 535 2782 569
rect 2748 455 2782 489
rect 2904 697 2938 731
rect 2904 617 2938 651
rect 2904 535 2938 569
rect 2904 455 2938 489
<< mvpsubdiff >>
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2719 17
rect 2753 -17 2815 17
rect 2849 -17 2911 17
rect 2945 -17 2976 17
<< mvnsubdiff >>
rect 0 797 31 831
rect 65 797 127 831
rect 161 797 223 831
rect 257 797 319 831
rect 353 797 415 831
rect 449 797 511 831
rect 545 797 607 831
rect 641 797 703 831
rect 737 797 799 831
rect 833 797 895 831
rect 929 797 991 831
rect 1025 797 1087 831
rect 1121 797 1183 831
rect 1217 797 1279 831
rect 1313 797 1375 831
rect 1409 797 1471 831
rect 1505 797 1567 831
rect 1601 797 1663 831
rect 1697 797 1759 831
rect 1793 797 1855 831
rect 1889 797 1951 831
rect 1985 797 2047 831
rect 2081 797 2143 831
rect 2177 797 2239 831
rect 2273 797 2335 831
rect 2369 797 2431 831
rect 2465 797 2527 831
rect 2561 797 2623 831
rect 2657 797 2719 831
rect 2753 797 2815 831
rect 2849 797 2911 831
rect 2945 797 2976 831
<< mvpsubdiffcont >>
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
rect 2047 -17 2081 17
rect 2143 -17 2177 17
rect 2239 -17 2273 17
rect 2335 -17 2369 17
rect 2431 -17 2465 17
rect 2527 -17 2561 17
rect 2623 -17 2657 17
rect 2719 -17 2753 17
rect 2815 -17 2849 17
rect 2911 -17 2945 17
<< mvnsubdiffcont >>
rect 31 797 65 831
rect 127 797 161 831
rect 223 797 257 831
rect 319 797 353 831
rect 415 797 449 831
rect 511 797 545 831
rect 607 797 641 831
rect 703 797 737 831
rect 799 797 833 831
rect 895 797 929 831
rect 991 797 1025 831
rect 1087 797 1121 831
rect 1183 797 1217 831
rect 1279 797 1313 831
rect 1375 797 1409 831
rect 1471 797 1505 831
rect 1567 797 1601 831
rect 1663 797 1697 831
rect 1759 797 1793 831
rect 1855 797 1889 831
rect 1951 797 1985 831
rect 2047 797 2081 831
rect 2143 797 2177 831
rect 2239 797 2273 831
rect 2335 797 2369 831
rect 2431 797 2465 831
rect 2527 797 2561 831
rect 2623 797 2657 831
rect 2719 797 2753 831
rect 2815 797 2849 831
rect 2911 797 2945 831
<< poly >>
rect 87 677 187 786
rect 243 677 343 786
rect 858 743 958 769
rect 1124 743 1224 769
rect 1867 743 1967 769
rect 2023 743 2123 769
rect 2527 743 2627 769
rect 2793 743 2893 769
rect 385 677 485 703
rect 541 677 641 703
rect 683 677 783 703
rect 1390 627 1490 653
rect 1546 627 1646 653
rect 1688 627 1788 653
rect 87 571 187 593
rect 243 571 343 593
rect 87 537 343 571
rect 87 471 229 537
rect 385 495 485 593
rect 271 475 421 495
rect 87 418 191 471
rect 86 398 191 418
rect 86 364 137 398
rect 171 364 191 398
rect 86 330 191 364
rect 86 296 137 330
rect 171 296 191 330
rect 271 441 310 475
rect 344 441 421 475
rect 541 453 641 593
rect 271 439 421 441
rect 271 397 364 439
rect 463 397 641 453
rect 683 567 783 593
rect 683 545 790 567
rect 683 511 736 545
rect 770 511 790 545
rect 683 477 790 511
rect 683 443 736 477
rect 770 443 790 477
rect 683 423 790 443
rect 271 317 342 397
rect 406 355 498 397
rect 86 276 191 296
rect 86 191 186 276
rect 242 191 342 317
rect 384 335 498 355
rect 384 301 411 335
rect 445 301 498 335
rect 384 267 498 301
rect 384 233 411 267
rect 445 233 498 267
rect 384 213 498 233
rect 540 335 640 355
rect 540 301 560 335
rect 594 301 640 335
rect 690 317 790 423
rect 858 357 958 593
rect 1124 567 1224 593
rect 1051 545 1224 567
rect 1051 511 1071 545
rect 1105 511 1224 545
rect 2202 627 2302 653
rect 2352 627 2452 653
rect 1390 521 1490 543
rect 1051 477 1224 511
rect 1051 443 1071 477
rect 1105 443 1224 477
rect 1051 423 1224 443
rect 1362 495 1490 521
rect 1362 461 1408 495
rect 1442 461 1490 495
rect 1362 446 1490 461
rect 1546 495 1646 543
rect 1546 461 1592 495
rect 1626 461 1646 495
rect 1362 441 1462 446
rect 1546 435 1646 461
rect 540 267 640 301
rect 540 233 560 267
rect 594 233 640 267
rect 384 191 484 213
rect 540 191 640 233
rect 682 217 790 317
rect 838 337 958 357
rect 1124 399 1224 423
rect 1538 427 1646 435
rect 1538 404 1592 427
rect 1504 399 1592 404
rect 1124 393 1592 399
rect 1626 393 1646 427
rect 1124 355 1646 393
rect 1688 517 1788 543
rect 1688 495 1794 517
rect 1688 461 1740 495
rect 1774 461 1794 495
rect 1688 427 1794 461
rect 1688 393 1740 427
rect 1774 393 1794 427
rect 1688 373 1794 393
rect 838 303 885 337
rect 919 303 958 337
rect 838 269 958 303
rect 838 235 885 269
rect 919 235 958 269
rect 682 191 782 217
rect 838 215 958 235
rect 1104 335 1646 355
rect 1104 301 1124 335
rect 1158 329 1638 335
rect 1158 301 1504 329
rect 1694 313 1794 373
rect 1104 267 1504 301
rect 1104 233 1124 267
rect 1158 255 1504 267
rect 1546 267 1646 287
rect 1158 233 1204 255
rect 838 191 938 215
rect 1104 191 1204 233
rect 1390 191 1490 255
rect 1546 233 1592 267
rect 1626 233 1646 267
rect 1546 191 1646 233
rect 1688 213 1794 313
rect 1867 355 1967 543
rect 2023 495 2123 543
rect 2023 461 2048 495
rect 2082 461 2123 495
rect 2023 441 2123 461
rect 2202 399 2302 543
rect 1867 321 1887 355
rect 1921 321 1967 355
rect 1867 257 1967 321
rect 2009 339 2302 399
rect 2009 305 2025 339
rect 2059 329 2302 339
rect 2352 435 2452 543
rect 2527 517 2627 543
rect 2516 487 2627 517
rect 2516 453 2536 487
rect 2570 453 2627 487
rect 2352 415 2466 435
rect 2352 381 2412 415
rect 2446 381 2466 415
rect 2352 347 2466 381
rect 2516 419 2627 453
rect 2516 385 2536 419
rect 2570 385 2627 419
rect 2793 417 2893 443
rect 2516 365 2627 385
rect 2059 305 2146 329
rect 2009 285 2146 305
rect 2352 313 2412 347
rect 2446 313 2466 347
rect 2352 293 2466 313
rect 1688 191 1788 213
rect 2046 191 2146 285
rect 2210 267 2310 287
rect 2210 233 2254 267
rect 2288 233 2310 267
rect 2210 191 2310 233
rect 2352 191 2452 293
rect 2527 257 2627 365
rect 2669 387 2893 417
rect 2669 353 2689 387
rect 2723 353 2893 387
rect 2669 303 2893 353
rect 2793 277 2893 303
rect 86 81 186 107
rect 242 81 342 107
rect 384 81 484 107
rect 540 81 640 107
rect 682 81 782 107
rect 838 81 938 107
rect 1104 81 1204 107
rect 1390 81 1490 107
rect 1546 81 1646 107
rect 1688 81 1788 107
rect 1867 81 1967 107
rect 2046 81 2146 107
rect 2210 81 2310 107
rect 2352 81 2452 107
rect 2527 81 2627 107
rect 2793 101 2893 127
<< polycont >>
rect 137 364 171 398
rect 137 296 171 330
rect 310 441 344 475
rect 736 511 770 545
rect 736 443 770 477
rect 411 301 445 335
rect 411 233 445 267
rect 560 301 594 335
rect 1071 511 1105 545
rect 1071 443 1105 477
rect 1408 461 1442 495
rect 1592 461 1626 495
rect 560 233 594 267
rect 1592 393 1626 427
rect 1740 461 1774 495
rect 1740 393 1774 427
rect 885 303 919 337
rect 885 235 919 269
rect 1124 301 1158 335
rect 1124 233 1158 267
rect 1592 233 1626 267
rect 2048 461 2082 495
rect 1887 321 1921 355
rect 2025 305 2059 339
rect 2536 453 2570 487
rect 2412 381 2446 415
rect 2536 385 2570 419
rect 2412 313 2446 347
rect 2254 233 2288 267
rect 2689 353 2723 387
<< locali >>
rect 0 797 31 831
rect 65 797 127 831
rect 161 797 223 831
rect 257 797 319 831
rect 353 797 415 831
rect 449 797 511 831
rect 545 797 607 831
rect 641 797 703 831
rect 737 797 799 831
rect 833 797 895 831
rect 929 797 991 831
rect 1025 797 1087 831
rect 1121 797 1183 831
rect 1217 797 1279 831
rect 1313 797 1375 831
rect 1409 797 1471 831
rect 1505 797 1567 831
rect 1601 797 1663 831
rect 1697 797 1759 831
rect 1793 797 1855 831
rect 1889 797 1951 831
rect 1985 797 2047 831
rect 2081 797 2143 831
rect 2177 797 2239 831
rect 2273 797 2335 831
rect 2369 797 2431 831
rect 2465 797 2527 831
rect 2561 797 2623 831
rect 2657 797 2719 831
rect 2753 797 2815 831
rect 2849 797 2911 831
rect 2945 797 2976 831
rect 182 735 372 741
rect 182 701 188 735
rect 222 701 260 735
rect 294 701 332 735
rect 366 701 372 735
rect 25 652 76 685
rect 25 618 42 652
rect 25 253 76 618
rect 182 652 372 701
rect 727 735 917 747
rect 727 701 733 735
rect 767 701 805 735
rect 839 731 877 735
rect 847 701 877 731
rect 911 701 917 735
rect 727 697 813 701
rect 847 697 917 701
rect 182 618 198 652
rect 232 618 372 652
rect 182 585 372 618
rect 480 652 546 685
rect 480 618 496 652
rect 530 619 546 652
rect 727 639 917 697
rect 530 618 680 619
rect 480 585 680 618
rect 727 605 813 639
rect 847 605 917 639
rect 727 589 917 605
rect 953 731 1019 747
rect 953 697 969 731
rect 1003 697 1019 731
rect 953 639 1019 697
rect 953 605 969 639
rect 1003 605 1019 639
rect 121 475 551 504
rect 121 441 310 475
rect 344 441 551 475
rect 646 407 680 585
rect 953 553 1019 605
rect 1063 735 1181 747
rect 1063 701 1069 735
rect 1103 731 1141 735
rect 1113 701 1141 731
rect 1175 701 1181 735
rect 1063 697 1079 701
rect 1113 697 1181 701
rect 1063 639 1181 697
rect 1063 605 1079 639
rect 1113 605 1181 639
rect 1063 589 1181 605
rect 1219 731 1285 747
rect 1219 697 1235 731
rect 1269 701 1285 731
rect 1806 741 1996 751
rect 1806 707 1812 741
rect 1846 735 1884 741
rect 1856 707 1884 735
rect 1918 707 1956 741
rect 1990 707 1996 741
rect 1806 701 1822 707
rect 1856 701 1996 707
rect 2396 735 2586 747
rect 2396 701 2402 735
rect 2436 701 2474 735
rect 2508 731 2546 735
rect 2516 701 2546 731
rect 2580 701 2586 735
rect 1269 697 1465 701
rect 1219 667 1465 697
rect 1219 639 1285 667
rect 1219 605 1235 639
rect 1269 605 1285 639
rect 1219 589 1285 605
rect 1322 602 1395 631
rect 1322 568 1345 602
rect 1379 568 1395 602
rect 720 545 839 553
rect 720 511 736 545
rect 770 511 839 545
rect 953 545 1121 553
rect 953 519 1071 545
rect 720 477 839 511
rect 720 443 736 477
rect 770 443 839 477
rect 1055 511 1071 519
rect 1105 511 1121 545
rect 1055 477 1121 511
rect 1055 443 1071 477
rect 1105 443 1121 477
rect 1322 539 1395 568
rect 1322 407 1356 539
rect 1431 503 1465 667
rect 2064 665 2290 699
rect 1392 495 1465 503
rect 1392 461 1408 495
rect 1442 461 1465 495
rect 1392 445 1465 461
rect 1501 602 1551 635
rect 1535 568 1551 602
rect 1501 535 1551 568
rect 1608 631 2098 665
rect 121 398 610 405
rect 121 364 137 398
rect 171 371 610 398
rect 171 364 359 371
rect 121 330 359 364
rect 544 335 610 371
rect 121 296 137 330
rect 171 296 359 330
rect 121 289 359 296
rect 395 301 411 335
rect 445 301 461 335
rect 395 267 461 301
rect 395 253 411 267
rect 25 233 411 253
rect 445 233 461 267
rect 25 219 461 233
rect 544 301 560 335
rect 594 301 610 335
rect 544 267 610 301
rect 544 233 560 267
rect 594 233 610 267
rect 544 219 610 233
rect 646 373 1356 407
rect 25 166 91 219
rect 646 183 680 373
rect 869 303 885 337
rect 919 303 935 337
rect 869 269 935 303
rect 869 235 885 269
rect 919 235 935 269
rect 1108 335 1174 337
rect 1108 301 1124 335
rect 1158 301 1174 335
rect 1108 267 1174 301
rect 1108 265 1124 267
rect 971 233 1124 265
rect 1158 233 1174 267
rect 971 231 1174 233
rect 25 132 41 166
rect 75 132 91 166
rect 25 103 91 132
rect 181 166 371 183
rect 181 132 197 166
rect 231 132 371 166
rect 181 113 371 132
rect 181 79 187 113
rect 221 79 259 113
rect 293 79 331 113
rect 365 79 371 113
rect 479 166 680 183
rect 479 132 495 166
rect 529 149 680 166
rect 716 166 897 199
rect 971 195 1005 231
rect 1313 199 1356 373
rect 529 132 545 149
rect 479 99 545 132
rect 716 132 793 166
rect 827 132 897 166
rect 716 113 897 132
rect 181 73 371 79
rect 716 79 718 113
rect 752 79 790 113
rect 824 79 862 113
rect 896 79 897 113
rect 933 166 1005 195
rect 933 132 949 166
rect 983 132 1005 166
rect 933 103 1005 132
rect 1043 166 1161 195
rect 1043 132 1059 166
rect 1093 132 1161 166
rect 1043 113 1161 132
rect 716 73 897 79
rect 1043 79 1049 113
rect 1083 79 1121 113
rect 1155 79 1161 113
rect 1043 73 1161 79
rect 1199 166 1265 195
rect 1199 132 1215 166
rect 1249 132 1265 166
rect 1199 87 1265 132
rect 1313 170 1379 199
rect 1313 136 1329 170
rect 1363 136 1379 170
rect 1313 123 1379 136
rect 1415 87 1449 445
rect 1501 355 1535 535
rect 1608 499 1642 631
rect 1962 590 2028 595
rect 1962 556 1978 590
rect 2012 556 2028 590
rect 1962 535 2028 556
rect 1576 495 1642 499
rect 1576 461 1592 495
rect 1626 461 1642 495
rect 1576 427 1642 461
rect 1576 393 1592 427
rect 1626 393 1642 427
rect 1576 391 1642 393
rect 1724 495 1790 511
rect 1724 461 1740 495
rect 1774 461 1790 495
rect 1724 427 1790 461
rect 1724 393 1740 427
rect 1774 425 1790 427
rect 1962 425 1996 535
rect 2064 499 2098 631
rect 2134 599 2215 629
rect 2168 565 2215 599
rect 2134 535 2215 565
rect 2032 495 2098 499
rect 2032 461 2048 495
rect 2082 461 2098 495
rect 1774 393 2129 425
rect 1724 391 2129 393
rect 1501 321 1887 355
rect 1921 321 1937 355
rect 2009 339 2059 355
rect 1501 199 1551 321
rect 2009 305 2025 339
rect 2009 285 2059 305
rect 1485 170 1551 199
rect 1485 136 1501 170
rect 1535 136 1551 170
rect 1485 123 1551 136
rect 1587 267 2059 285
rect 1587 233 1592 267
rect 1626 251 2059 267
rect 1626 233 1642 251
rect 1587 87 1642 233
rect 2095 215 2129 391
rect 1199 53 1642 87
rect 1736 182 1926 215
rect 1736 148 1822 182
rect 1856 148 1926 182
rect 1736 113 1926 148
rect 1736 79 1742 113
rect 1776 79 1814 113
rect 1848 79 1886 113
rect 1920 79 1926 113
rect 1962 182 2129 215
rect 1962 148 1978 182
rect 2012 181 2129 182
rect 2012 148 2028 181
rect 1962 99 2028 148
rect 2165 166 2215 535
rect 2251 267 2290 665
rect 2396 697 2482 701
rect 2516 697 2586 701
rect 2396 660 2586 697
rect 2396 626 2482 660
rect 2516 626 2586 660
rect 2396 589 2586 626
rect 2396 555 2482 589
rect 2516 555 2586 589
rect 2396 539 2586 555
rect 2622 731 2688 747
rect 2622 697 2638 731
rect 2672 697 2688 731
rect 2622 660 2688 697
rect 2622 626 2638 660
rect 2672 626 2688 660
rect 2622 589 2688 626
rect 2622 555 2638 589
rect 2672 555 2688 589
rect 2251 233 2254 267
rect 2288 233 2290 267
rect 2251 217 2290 233
rect 2326 487 2586 503
rect 2326 469 2536 487
rect 2199 133 2215 166
rect 2326 133 2360 469
rect 2520 453 2536 469
rect 2570 453 2586 487
rect 2396 415 2462 431
rect 2396 381 2412 415
rect 2446 381 2462 415
rect 2396 347 2462 381
rect 2520 419 2586 453
rect 2520 385 2536 419
rect 2570 385 2586 419
rect 2520 369 2586 385
rect 2622 403 2688 555
rect 2732 731 2804 747
rect 2732 697 2748 731
rect 2782 697 2804 731
rect 2732 651 2804 697
rect 2732 617 2748 651
rect 2782 617 2804 651
rect 2732 569 2804 617
rect 2732 535 2748 569
rect 2782 535 2804 569
rect 2732 489 2804 535
rect 2732 455 2748 489
rect 2782 455 2804 489
rect 2732 439 2804 455
rect 2840 735 2958 747
rect 2840 701 2846 735
rect 2880 731 2918 735
rect 2880 701 2904 731
rect 2952 701 2958 735
rect 2840 697 2904 701
rect 2938 697 2958 701
rect 2840 651 2958 697
rect 2840 617 2904 651
rect 2938 617 2958 651
rect 2840 569 2958 617
rect 2840 535 2904 569
rect 2938 535 2958 569
rect 2840 489 2958 535
rect 2840 455 2904 489
rect 2938 455 2958 489
rect 2840 439 2958 455
rect 2622 387 2734 403
rect 2396 313 2412 347
rect 2446 331 2462 347
rect 2622 353 2689 387
rect 2723 353 2734 387
rect 2622 337 2734 353
rect 2770 356 2804 439
rect 2622 331 2688 337
rect 2446 313 2688 331
rect 2396 297 2688 313
rect 2770 301 2951 356
rect 2199 132 2360 133
rect 2165 99 2360 132
rect 2396 245 2586 261
rect 2396 211 2482 245
rect 2516 211 2586 245
rect 2396 153 2586 211
rect 2396 119 2482 153
rect 2516 119 2586 153
rect 2396 113 2586 119
rect 1736 73 1926 79
rect 2396 79 2402 113
rect 2436 79 2474 113
rect 2508 79 2546 113
rect 2580 79 2586 113
rect 2622 245 2688 297
rect 2622 211 2638 245
rect 2672 211 2688 245
rect 2622 153 2688 211
rect 2622 119 2638 153
rect 2672 119 2688 153
rect 2732 265 2804 301
rect 2732 231 2748 265
rect 2782 231 2804 265
rect 2732 173 2804 231
rect 2732 139 2748 173
rect 2782 139 2804 173
rect 2732 123 2804 139
rect 2840 231 2904 265
rect 2938 231 2958 265
rect 2840 173 2958 231
rect 2840 139 2904 173
rect 2938 139 2958 173
rect 2622 103 2688 119
rect 2840 113 2958 139
rect 2396 73 2586 79
rect 2840 79 2846 113
rect 2880 79 2918 113
rect 2952 79 2958 113
rect 2840 73 2958 79
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2719 17
rect 2753 -17 2815 17
rect 2849 -17 2911 17
rect 2945 -17 2976 17
<< viali >>
rect 31 797 65 831
rect 127 797 161 831
rect 223 797 257 831
rect 319 797 353 831
rect 415 797 449 831
rect 511 797 545 831
rect 607 797 641 831
rect 703 797 737 831
rect 799 797 833 831
rect 895 797 929 831
rect 991 797 1025 831
rect 1087 797 1121 831
rect 1183 797 1217 831
rect 1279 797 1313 831
rect 1375 797 1409 831
rect 1471 797 1505 831
rect 1567 797 1601 831
rect 1663 797 1697 831
rect 1759 797 1793 831
rect 1855 797 1889 831
rect 1951 797 1985 831
rect 2047 797 2081 831
rect 2143 797 2177 831
rect 2239 797 2273 831
rect 2335 797 2369 831
rect 2431 797 2465 831
rect 2527 797 2561 831
rect 2623 797 2657 831
rect 2719 797 2753 831
rect 2815 797 2849 831
rect 2911 797 2945 831
rect 188 701 222 735
rect 260 701 294 735
rect 332 701 366 735
rect 733 701 767 735
rect 805 731 839 735
rect 805 701 813 731
rect 813 701 839 731
rect 877 701 911 735
rect 1069 731 1103 735
rect 1069 701 1079 731
rect 1079 701 1103 731
rect 1141 701 1175 735
rect 1812 735 1846 741
rect 1812 707 1822 735
rect 1822 707 1846 735
rect 1884 707 1918 741
rect 1956 707 1990 741
rect 2402 701 2436 735
rect 2474 731 2508 735
rect 2474 701 2482 731
rect 2482 701 2508 731
rect 2546 701 2580 735
rect 187 79 221 113
rect 259 79 293 113
rect 331 79 365 113
rect 718 79 752 113
rect 790 79 824 113
rect 862 79 896 113
rect 1049 79 1083 113
rect 1121 79 1155 113
rect 1742 79 1776 113
rect 1814 79 1848 113
rect 1886 79 1920 113
rect 2846 701 2880 735
rect 2918 731 2952 735
rect 2918 701 2938 731
rect 2938 701 2952 731
rect 2402 79 2436 113
rect 2474 79 2508 113
rect 2546 79 2580 113
rect 2846 79 2880 113
rect 2918 79 2952 113
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
rect 2047 -17 2081 17
rect 2143 -17 2177 17
rect 2239 -17 2273 17
rect 2335 -17 2369 17
rect 2431 -17 2465 17
rect 2527 -17 2561 17
rect 2623 -17 2657 17
rect 2719 -17 2753 17
rect 2815 -17 2849 17
rect 2911 -17 2945 17
<< metal1 >>
rect 0 831 2976 837
rect 0 797 31 831
rect 65 797 127 831
rect 161 797 223 831
rect 257 797 319 831
rect 353 797 415 831
rect 449 797 511 831
rect 545 797 607 831
rect 641 797 703 831
rect 737 797 799 831
rect 833 797 895 831
rect 929 797 991 831
rect 1025 797 1087 831
rect 1121 797 1183 831
rect 1217 797 1279 831
rect 1313 797 1375 831
rect 1409 797 1471 831
rect 1505 797 1567 831
rect 1601 797 1663 831
rect 1697 797 1759 831
rect 1793 797 1855 831
rect 1889 797 1951 831
rect 1985 797 2047 831
rect 2081 797 2143 831
rect 2177 797 2239 831
rect 2273 797 2335 831
rect 2369 797 2431 831
rect 2465 797 2527 831
rect 2561 797 2623 831
rect 2657 797 2719 831
rect 2753 797 2815 831
rect 2849 797 2911 831
rect 2945 797 2976 831
rect 0 791 2976 797
rect 0 741 2976 763
rect 0 735 1812 741
rect 0 701 188 735
rect 222 701 260 735
rect 294 701 332 735
rect 366 701 733 735
rect 767 701 805 735
rect 839 701 877 735
rect 911 701 1069 735
rect 1103 701 1141 735
rect 1175 707 1812 735
rect 1846 707 1884 741
rect 1918 707 1956 741
rect 1990 735 2976 741
rect 1990 707 2402 735
rect 1175 701 2402 707
rect 2436 701 2474 735
rect 2508 701 2546 735
rect 2580 701 2846 735
rect 2880 701 2918 735
rect 2952 701 2976 735
rect 0 689 2976 701
rect 0 113 2976 125
rect 0 79 187 113
rect 221 79 259 113
rect 293 79 331 113
rect 365 79 718 113
rect 752 79 790 113
rect 824 79 862 113
rect 896 79 1049 113
rect 1083 79 1121 113
rect 1155 79 1742 113
rect 1776 79 1814 113
rect 1848 79 1886 113
rect 1920 79 2402 113
rect 2436 79 2474 113
rect 2508 79 2546 113
rect 2580 79 2846 113
rect 2880 79 2918 113
rect 2952 79 2976 113
rect 0 51 2976 79
rect 0 17 2976 23
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2719 17
rect 2753 -17 2815 17
rect 2849 -17 2911 17
rect 2945 -17 2976 17
rect 0 -23 2976 -17
<< labels >>
flabel comment s 1340 344 1340 344 0 FreeSans 200 0 0 0 no_jumper_check
rlabel comment s 0 0 0 0 4 sdfxtp_1
flabel metal1 s 0 51 2976 125 0 FreeSans 340 0 0 0 VGND
port 5 nsew ground bidirectional
flabel metal1 s 0 0 2976 23 0 FreeSans 340 0 0 0 VNB
port 6 nsew ground bidirectional
flabel metal1 s 0 689 2976 763 0 FreeSans 340 0 0 0 VPWR
port 8 nsew power bidirectional
flabel metal1 s 0 791 2976 814 0 FreeSans 340 0 0 0 VPB
port 7 nsew power bidirectional
flabel locali s 511 464 545 498 0 FreeSans 340 180 0 0 D
port 2 nsew signal input
flabel locali s 415 464 449 498 0 FreeSans 340 180 0 0 D
port 2 nsew signal input
flabel locali s 319 464 353 498 0 FreeSans 340 180 0 0 D
port 2 nsew signal input
flabel locali s 223 464 257 498 0 FreeSans 340 180 0 0 D
port 2 nsew signal input
flabel locali s 127 464 161 498 0 FreeSans 340 180 0 0 D
port 2 nsew signal input
flabel locali s 799 464 833 498 0 FreeSans 340 180 0 0 SCD
port 3 nsew signal input
flabel locali s 319 316 353 350 0 FreeSans 340 180 0 0 SCE
port 4 nsew signal input
flabel locali s 223 316 257 350 0 FreeSans 340 180 0 0 SCE
port 4 nsew signal input
flabel locali s 127 316 161 350 0 FreeSans 340 180 0 0 SCE
port 4 nsew signal input
flabel locali s 895 242 929 276 0 FreeSans 340 180 0 0 CLK
port 1 nsew clock input
flabel locali s 2911 316 2945 350 0 FreeSans 340 180 0 0 Q
port 9 nsew signal output
flabel locali s 2815 316 2849 350 0 FreeSans 340 180 0 0 Q
port 9 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 2976 814
string GDS_END 672124
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hvl/gds/sky130_fd_sc_hvl.gds
string GDS_START 643136
string LEFclass CORE
string LEFsite unithv
string LEFsymmetry X Y
<< end >>
