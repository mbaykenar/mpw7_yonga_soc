* SKY130 Spice File.
.option scale = 1.0u
.include "invariant.spice"
* Derivative Parameters:
.param
+ c0m4m3_vpp = '9.09375e-03*ic_cap*ic_cap+8.53750e-02*ic_cap+1.00000e+00'
+ c0m5m3_vpp = '5.28125e-03*ic_cap*ic_cap+7.03750e-02*ic_cap+1.00000e+00'
+ c0m5m4_vpp = '9.09375e-03*ic_cap*ic_cap+8.53750e-02*ic_cap+1.00000e+00'
+ c0m5m4_vpp0p4shield = '5.14350e-02*ic_cap*ic_cap+3.04590e-01*ic_cap+1.00000e+00'
+ c1m4m3_vpp = '5.78125e-03*ic_cap*ic_cap+8.16250e-02*ic_cap+1.00000e+00'
+ c1m5m3_vpp = '8.43750e-03*ic_cap*ic_cap+9.02500e-02*ic_cap+1.00000e+00'
+ c1m5m4_vpp = '5.78125e-03*ic_cap*ic_cap+8.16250e-02*ic_cap+1.00000e+00'
+ c1m5m4_vpp0p4shield = '8.44188e-03*ic_cap*ic_cap+9.22675e-02*ic_cap+1.00000e+00'
+ camimc = '2.81250e-19*mim*mim+5.66250e-17*mim+2.00000e-15'
+ cl1d = '-5.50000e-07*ic_cap*ic_cap+-3.00000e-07*ic_cap+5.53000e-05'
+ cl1dsw = '-7.96875e-13*ic_cap*ic_cap+-5.12500e-13*ic_cap+8.23000e-11'
+ cl1f = '-4.15625e-07*ic_cap*ic_cap+-2.37500e-07*ic_cap+3.69000e-05'
+ cl1fsw = '-8.03125e-13*ic_cap*ic_cap+-5.37500e-13*ic_cap+8.30000e-11'
+ cl1p1 = '-1.65000e-06*ic_cap*ic_cap+-8.00000e-07*ic_cap+9.41000e-05'
+ cl1p1f = '-3.03125e-06*ic_cap*ic_cap+-1.62500e-06*ic_cap+2.00000e-04'
+ cl1p1fsw = '-5.90625e-13*ic_cap*ic_cap+-3.12500e-13*ic_cap+8.32000e-11'
+ cl1p1sw = '-7.68750e-13*ic_cap*ic_cap+-5.00000e-13*ic_cap+8.13000e-11'
+ cli2s_vpp = '4.40625e-03*ic_cap*ic_cap+6.91250e-02*ic_cap+1.00000e+00'
+ cm1d = '-3.71875e-07*ic_cap*ic_cap+-2.37500e-07*ic_cap+3.36000e-05'
+ cm1dsw = '-9.06250e-13*ic_cap*ic_cap+-4.75000e-13*ic_cap+1.06000e-10'
+ cm1f = '-3.03125e-07*ic_cap*ic_cap+-1.87500e-07*ic_cap+2.58000e-05'
+ cm1fsw = '-9.59375e-13*ic_cap*ic_cap+-4.87500e-13*ic_cap+1.07000e-10'
+ cm1l1 = '-1.98438e-06*ic_cap*ic_cap+-1.26250e-06*ic_cap+1.14000e-04'
+ cm1l1d = '-2.50000e-06*ic_cap*ic_cap+-1.50000e-06*ic_cap+1.69000e-04'
+ cm1l1dsw = '-6.93750e-13*ic_cap*ic_cap+-4.50000e-13*ic_cap+7.81000e-11'
+ cm1l1f = '-2.37500e-06*ic_cap*ic_cap+-1.50000e-06*ic_cap+1.51000e-04'
+ cm1l1fsw = '-7.09375e-13*ic_cap*ic_cap+-4.62500e-13*ic_cap+7.90000e-11'
+ cm1l1p1 = '-3.59375e-06*ic_cap*ic_cap+-2.12500e-06*ic_cap+2.08000e-04'
+ cm1l1p1sw = '-6.68750e-13*ic_cap*ic_cap+-4.25000e-13*ic_cap+7.71000e-11'
+ cm1l1sw = '-8.09375e-13*ic_cap*ic_cap+-4.87500e-13*ic_cap+1.03000e-10'
+ cm1p1 = '-6.81250e-07*ic_cap*ic_cap+-4.00000e-07*ic_cap+4.48000e-05'
+ cm1p1f = '-2.09375e-06*ic_cap*ic_cap+-1.12500e-06*ic_cap+1.51000e-04'
+ cm1p1fsw = '-6.12500e-13*ic_cap*ic_cap+-3.50000e-13*ic_cap+8.45000e-11'
+ cm1p1sw = '-9.28125e-13*ic_cap*ic_cap+-4.87500e-13*ic_cap+1.06000e-10'
+ cm2d = '-2.15625e-07*ic_cap*ic_cap+-1.37500e-07*ic_cap+2.08000e-05'
+ cm2dsw = '-9.50000e-13*ic_cap*ic_cap+-5.00000e-13*ic_cap+1.07000e-10'
+ cm2f = '-1.90625e-07*ic_cap*ic_cap+-1.12500e-07*ic_cap+1.75000e-05'
+ cm2fsw = '-1.00938e-12*ic_cap*ic_cap+-5.12500e-13*ic_cap+1.08000e-10'
+ cm2l1 = '-4.50000e-07*ic_cap*ic_cap+-3.00000e-07*ic_cap+3.70000e-05'
+ cm2l1d = '-1.00000e-06*ic_cap*ic_cap+-6.00000e-07*ic_cap+9.23000e-05'
+ cm2l1dsw = '-7.43750e-13*ic_cap*ic_cap+-4.75000e-13*ic_cap+8.04000e-11'
+ cm2l1f = '-8.68750e-07*ic_cap*ic_cap+-5.25000e-07*ic_cap+7.40000e-05'
+ cm2l1fsw = '-7.65625e-13*ic_cap*ic_cap+-5.12500e-13*ic_cap+8.14000e-11'
+ cm2l1p1 = '-2.08750e-06*ic_cap*ic_cap+-1.10000e-06*ic_cap+1.31000e-04'
+ cm2l1p1sw = '-7.18750e-13*ic_cap*ic_cap+-4.50000e-13*ic_cap+7.94000e-11'
+ cm2l1sw = '-9.15625e-13*ic_cap*ic_cap+-5.37500e-13*ic_cap+1.06000e-10'
+ cm2m1 = '-2.66250e-06*ic_cap*ic_cap+-1.25000e-06*ic_cap+1.28000e-04'
+ cm2m1d = '-3.06250e-06*ic_cap*ic_cap+-1.50000e-06*ic_cap+1.62000e-04'
+ cm2m1dsw = '-7.96875e-13*ic_cap*ic_cap+-4.37500e-13*ic_cap+1.02000e-10'
+ cm2m1f = '-2.96875e-06*ic_cap*ic_cap+-1.37500e-06*ic_cap+1.54000e-04'
+ cm2m1fsw = '-7.93750e-13*ic_cap*ic_cap+-4.00000e-13*ic_cap+1.02000e-10'
+ cm2m1l1 = '-4.62500e-06*ic_cap*ic_cap+-2.50000e-06*ic_cap+2.42000e-04'
+ cm2m1l1sw = '-7.18750e-13*ic_cap*ic_cap+-4.00000e-13*ic_cap+9.89000e-11'
+ cm2m1p1 = '-3.34375e-06*ic_cap*ic_cap+-1.62500e-06*ic_cap+1.73000e-04'
+ cm2m1p1sw = '-7.50000e-13*ic_cap*ic_cap+-4.25000e-13*ic_cap+1.01000e-10'
+ cm2m1sw = '-8.18750e-13*ic_cap*ic_cap+-5.25000e-13*ic_cap+1.03000e-10'
+ cm2p1 = '-3.15625e-07*ic_cap*ic_cap+-1.87500e-07*ic_cap+2.47000e-05'
+ cm2p1f = '-1.73750e-06*ic_cap*ic_cap+-9.50000e-07*ic_cap+1.31000e-04'
+ cm2p1fsw = '-6.28125e-13*ic_cap*ic_cap+-3.62500e-13*ic_cap+8.53000e-11'
+ cm2p1sw = '-9.62500e-13*ic_cap*ic_cap+-5.25000e-13*ic_cap+1.07000e-10'
+ cm3d = '-1.37500e-07*ic_cap*ic_cap+-7.50000e-08*ic_cap+1.42000e-05'
+ cm3dsw = '-8.53125e-13*ic_cap*ic_cap+-4.62500e-13*ic_cap+1.09000e-10'
+ cm3f = '-1.31250e-07*ic_cap*ic_cap+-7.50000e-08*ic_cap+1.26000e-05'
+ cm3fsw = '-7.78125e-13*ic_cap*ic_cap+-4.62500e-13*ic_cap+1.08000e-10'
+ cm3l1 = '-2.09375e-07*ic_cap*ic_cap+-1.37500e-07*ic_cap+2.02000e-05'
+ cm3l1d = '-7.53125e-07*ic_cap*ic_cap+-4.37500e-07*ic_cap+7.54000e-05'
+ cm3l1dsw = '-7.65625e-13*ic_cap*ic_cap+-4.87500e-13*ic_cap+8.13000e-11'
+ cm3l1f = '-6.21875e-07*ic_cap*ic_cap+-3.62500e-07*ic_cap+5.71000e-05'
+ cm3l1fsw = '-7.75000e-13*ic_cap*ic_cap+-5.25000e-13*ic_cap+8.21000e-11'
+ cm3l1p1 = '-1.83750e-06*ic_cap*ic_cap+-9.25000e-07*ic_cap+1.14000e-04'
+ cm3l1p1sw = '-7.40625e-13*ic_cap*ic_cap+-4.87500e-13*ic_cap+8.04000e-11'
+ cm3l1sw = '-8.15625e-13*ic_cap*ic_cap+-4.62500e-13*ic_cap+1.08000e-10'
+ cm3m1 = '-3.90625e-07*ic_cap*ic_cap+-2.12500e-07*ic_cap+3.29000e-05'
+ cm3m1d = '-7.59375e-07*ic_cap*ic_cap+-4.62500e-07*ic_cap+6.65000e-05'
+ cm3m1dsw = '-8.56250e-13*ic_cap*ic_cap+-5.50000e-13*ic_cap+1.04000e-10'
+ cm3m1f = '-6.90625e-07*ic_cap*ic_cap+-4.12500e-07*ic_cap+5.87000e-05'
+ cm3m1fsw = '-8.93750e-13*ic_cap*ic_cap+-5.00000e-13*ic_cap+1.05000e-10'
+ cm3m1l1 = '-2.37500e-06*ic_cap*ic_cap+-1.50000e-06*ic_cap+1.47000e-04'
+ cm3m1l1sw = '-8.28125e-13*ic_cap*ic_cap+-3.62500e-13*ic_cap+1.02000e-10'
+ cm3m1p1 = '-1.07500e-06*ic_cap*ic_cap+-6.25000e-07*ic_cap+7.78000e-05'
+ cm3m1p1sw = '-8.65625e-13*ic_cap*ic_cap+-5.37500e-13*ic_cap+1.04000e-10'
+ cm3m1sw = '-7.96875e-13*ic_cap*ic_cap+-4.37500e-13*ic_cap+1.07000e-10'
+ cm3m2 = '-1.25000e-06*ic_cap*ic_cap+-6.75000e-07*ic_cap+8.22000e-05'
+ cm3m2_vpp = '2.06250e-03*ic_cap*ic_cap+1.46750e-01*ic_cap+1.00000e+00'
+ cm3m2d = '-1.46563e-06*ic_cap*ic_cap+-8.12500e-07*ic_cap+1.03000e-04'
+ cm3m2dsw = '-8.09375e-13*ic_cap*ic_cap+-4.37500e-13*ic_cap+1.03000e-10'
+ cm3m2f = '-1.45000e-06*ic_cap*ic_cap+-8.00000e-07*ic_cap+9.98000e-05'
+ cm3m2fsw = '-8.18750e-13*ic_cap*ic_cap+-4.00000e-13*ic_cap+1.03000e-10'
+ cm3m2l1 = '-1.69063e-06*ic_cap*ic_cap+-9.62500e-07*ic_cap+1.19000e-04'
+ cm3m2l1sw = '-7.65625e-13*ic_cap*ic_cap+-4.62500e-13*ic_cap+1.02000e-10'
+ cm3m2m1 = '-3.90625e-06*ic_cap*ic_cap+-1.87500e-06*ic_cap+2.10000e-04'
+ cm3m2m1sw = '-7.53125e-13*ic_cap*ic_cap+-4.37500e-13*ic_cap+9.97000e-11'
+ cm3m2p1 = '-1.57188e-06*ic_cap*ic_cap+-8.62500e-07*ic_cap+1.07000e-04'
+ cm3m2p1sw = '-8.90625e-13*ic_cap*ic_cap+-3.87500e-13*ic_cap+1.04000e-10'
+ cm3m2sw = '-7.59375e-13*ic_cap*ic_cap+-4.12500e-13*ic_cap+1.05000e-10'
+ cm3p1 = '-1.71875e-07*ic_cap*ic_cap+-1.12500e-07*ic_cap+1.58000e-05'
+ cm3p1f = '-1.59062e-06*ic_cap*ic_cap+-8.62500e-07*ic_cap+1.22000e-04'
+ cm3p1fsw = '-6.43750e-13*ic_cap*ic_cap+-3.75000e-13*ic_cap+8.58000e-11'
+ cm3p1sw = '-7.90625e-13*ic_cap*ic_cap+-4.62500e-13*ic_cap+1.08000e-10'
+ cm4d = '-7.71875e-08*ic_cap*ic_cap+-4.87500e-08*ic_cap+9.41000e-06'
+ cm4dsw = '-8.12500e-13*ic_cap*ic_cap+-5.00000e-13*ic_cap+1.09000e-10'
+ cm4f = '-7.50000e-08*ic_cap*ic_cap+-4.75000e-08*ic_cap+8.67000e-06'
+ cm4fsw = '-8.09375e-13*ic_cap*ic_cap+-4.87500e-13*ic_cap+1.09000e-10'
+ cm4l1 = '-9.62500e-08*ic_cap*ic_cap+-6.00000e-08*ic_cap+1.17000e-05'
+ cm4l1d = '-6.46875e-07*ic_cap*ic_cap+-3.62500e-07*ic_cap+6.70000e-05'
+ cm4l1dsw = '-7.81250e-13*ic_cap*ic_cap+-5.00000e-13*ic_cap+8.18000e-11'
+ cm4l1f = '-5.09375e-07*ic_cap*ic_cap+-2.87500e-07*ic_cap+4.86000e-05'
+ cm4l1fsw = '-7.87500e-13*ic_cap*ic_cap+-5.25000e-13*ic_cap+8.26000e-11'
+ cm4l1p1 = '-1.75938e-06*ic_cap*ic_cap+-8.62500e-07*ic_cap+1.06000e-04'
+ cm4l1p1sw = '-7.53125e-13*ic_cap*ic_cap+-4.87500e-13*ic_cap+8.08000e-11'
+ cm4l1sw = '-8.28125e-13*ic_cap*ic_cap+-4.87500e-13*ic_cap+1.09000e-10'
+ cm4m1 = '-1.25000e-07*ic_cap*ic_cap+-7.50000e-08*ic_cap+1.51000e-05'
+ cm4m1d = '-5.00000e-07*ic_cap*ic_cap+-3.25000e-07*ic_cap+4.87000e-05'
+ cm4m1dsw = '-9.25000e-13*ic_cap*ic_cap+-5.25000e-13*ic_cap+1.06000e-10'
+ cm4m1f = '-4.28125e-07*ic_cap*ic_cap+-2.62500e-07*ic_cap+4.09000e-05'
+ cm4m1fsw = '-9.75000e-13*ic_cap*ic_cap+-5.25000e-13*ic_cap+1.07000e-10'
+ cm4m1l1 = '-2.09375e-06*ic_cap*ic_cap+-1.37500e-06*ic_cap+1.29000e-04'
+ cm4m1l1sw = '-8.37500e-13*ic_cap*ic_cap+-4.25000e-13*ic_cap+1.03000e-10'
+ cm4m1p1 = '-8.09375e-07*ic_cap*ic_cap+-4.87500e-07*ic_cap+6.00000e-05'
+ cm4m1p1sw = '-9.31250e-13*ic_cap*ic_cap+-5.00000e-13*ic_cap+1.06000e-10'
+ cm4m1sw = '-7.81250e-13*ic_cap*ic_cap+-4.75000e-13*ic_cap+1.08000e-10'
+ cm4m2 = '-1.68750e-07*ic_cap*ic_cap+-1.00000e-07*ic_cap+2.09000e-05'
+ cm4m2d = '-3.84375e-07*ic_cap*ic_cap+-2.37500e-07*ic_cap+4.17000e-05'
+ cm4m2dsw = '-9.25000e-13*ic_cap*ic_cap+-5.25000e-13*ic_cap+1.06000e-10'
+ cm4m2f = '-3.62500e-07*ic_cap*ic_cap+-2.25000e-07*ic_cap+3.84000e-05'
+ cm4m2fsw = '-9.65625e-13*ic_cap*ic_cap+-4.87500e-13*ic_cap+1.07000e-10'
+ cm4m2l1 = '-6.21875e-07*ic_cap*ic_cap+-3.87500e-07*ic_cap+5.79000e-05'
+ cm4m2l1sw = '-8.87500e-13*ic_cap*ic_cap+-5.25000e-13*ic_cap+1.05000e-10'
+ cm4m2m1 = '-2.84062e-06*ic_cap*ic_cap+-1.36250e-06*ic_cap+1.49000e-04'
+ cm4m2m1sw = '-8.65625e-13*ic_cap*ic_cap+-3.62500e-13*ic_cap+1.03000e-10'
+ cm4m2p1 = '-4.84375e-07*ic_cap*ic_cap+-2.87500e-07*ic_cap+4.56000e-05'
+ cm4m2p1sw = '-9.21875e-13*ic_cap*ic_cap+-4.87500e-13*ic_cap+1.06000e-10'
+ cm4m2sw = '-8.09375e-13*ic_cap*ic_cap+-4.62500e-13*ic_cap+1.08000e-10'
+ cm4m3 = '-1.72187e-06*ic_cap*ic_cap+-8.37500e-07*ic_cap+8.85000e-05'
+ cm4m3d = '-1.87812e-06*ic_cap*ic_cap+-9.37500e-07*ic_cap+1.03000e-04'
+ cm4m3dsw = '-6.75000e-13*ic_cap*ic_cap+-4.00000e-13*ic_cap+1.03000e-10'
+ cm4m3f = '-1.84375e-06*ic_cap*ic_cap+-9.25000e-07*ic_cap+1.01000e-04'
+ cm4m3fsw = '-6.62500e-13*ic_cap*ic_cap+-4.00000e-13*ic_cap+1.03000e-10'
+ cm4m3l1 = '-1.95000e-06*ic_cap*ic_cap+-9.75000e-07*ic_cap+1.09000e-04'
+ cm4m3l1sw = '-7.09375e-13*ic_cap*ic_cap+-3.37500e-13*ic_cap+1.03000e-10'
+ cm4m3m1 = '-2.08750e-06*ic_cap*ic_cap+-1.07500e-06*ic_cap+1.21000e-04'
+ cm4m3m1sw = '-6.81250e-13*ic_cap*ic_cap+-3.75000e-13*ic_cap+1.02000e-10'
+ cm4m3m2 = '-3.00000e-06*ic_cap*ic_cap+-1.50000e-06*ic_cap+1.71000e-04'
+ cm4m3m2sw = '-6.34375e-13*ic_cap*ic_cap+-3.62500e-13*ic_cap+9.99000e-11'
+ cm4m3p1 = '-1.87500e-06*ic_cap*ic_cap+-9.50000e-07*ic_cap+1.04000e-04'
+ cm4m3p1sw = '-6.87500e-13*ic_cap*ic_cap+-4.25000e-13*ic_cap+1.03000e-10'
+ cm4m3sw = '-7.37500e-13*ic_cap*ic_cap+-4.50000e-13*ic_cap+1.05000e-10'
+ cm4p1 = '-9.06250e-08*ic_cap*ic_cap+-5.75000e-08*ic_cap+1.01000e-05'
+ cm4p1f = '-1.48437e-06*ic_cap*ic_cap+-8.37500e-07*ic_cap+1.16000e-04'
+ cm4p1fsw = '-6.50000e-13*ic_cap*ic_cap+-3.75000e-13*ic_cap+8.61000e-11'
+ cm4p1sw = '-8.18750e-13*ic_cap*ic_cap+-4.75000e-13*ic_cap+1.09000e-10'
+ cm5d = '-4.96875e-08*ic_cap*ic_cap+-3.12500e-08*ic_cap+6.88000e-06'
+ cm5dsw = '-4.93750e-13*ic_cap*ic_cap+-3.50000e-13*ic_cap+7.84000e-11'
+ cm5f = '-4.96875e-08*ic_cap*ic_cap+-3.12500e-08*ic_cap+6.48000e-06'
+ cm5fsw = '-4.90625e-13*ic_cap*ic_cap+-3.37500e-13*ic_cap+7.85000e-11'
+ cm5l1 = '-5.75000e-08*ic_cap*ic_cap+-3.75000e-08*ic_cap+8.04000e-06'
+ cm5l1d = '-6.06250e-07*ic_cap*ic_cap+-3.50000e-07*ic_cap+6.33000e-05'
+ cm5l1dsw = '-7.90625e-13*ic_cap*ic_cap+-5.12500e-13*ic_cap+8.20000e-11'
+ cm5l1f = '-4.68750e-07*ic_cap*ic_cap+-2.75000e-07*ic_cap+4.49000e-05'
+ cm5l1fsw = '-7.93750e-13*ic_cap*ic_cap+-5.25000e-13*ic_cap+8.28000e-11'
+ cm5l1p1 = '-1.70000e-06*ic_cap*ic_cap+-8.25000e-07*ic_cap+1.02000e-04'
+ cm5l1p1sw = '-7.53125e-13*ic_cap*ic_cap+-4.87500e-13*ic_cap+8.09000e-11'
+ cm5l1sw = '-4.84375e-13*ic_cap*ic_cap+-3.12500e-13*ic_cap+7.80000e-11'
+ cm5m1 = '-6.71875e-08*ic_cap*ic_cap+-4.12500e-08*ic_cap+9.50000e-06'
+ cm5m1d = '-4.40625e-07*ic_cap*ic_cap+-2.87500e-07*ic_cap+4.31000e-05'
+ cm5m1dsw = '-9.15625e-13*ic_cap*ic_cap+-5.37500e-13*ic_cap+1.06000e-10'
+ cm5m1f = '-3.68750e-07*ic_cap*ic_cap+-2.25000e-07*ic_cap+3.53000e-05'
+ cm5m1fsw = '-9.62500e-13*ic_cap*ic_cap+-5.50000e-13*ic_cap+1.07000e-10'
+ cm5m1l1 = '-2.01875e-06*ic_cap*ic_cap+-1.30000e-06*ic_cap+1.23000e-04'
+ cm5m1l1sw = '-8.84375e-13*ic_cap*ic_cap+-4.37500e-13*ic_cap+1.04000e-10'
+ cm5m1p1 = '-7.50000e-07*ic_cap*ic_cap+-4.50000e-07*ic_cap+5.44000e-05'
+ cm5m1p1sw = '-9.28125e-13*ic_cap*ic_cap+-5.12500e-13*ic_cap+1.06000e-10'
+ cm5m1sw = '-4.87500e-13*ic_cap*ic_cap+-3.25000e-13*ic_cap+7.77000e-11'
+ cm5m2 = '-7.50000e-08*ic_cap*ic_cap+-5.00000e-08*ic_cap+1.15000e-05'
+ cm5m2d = '-2.90625e-07*ic_cap*ic_cap+-1.87500e-07*ic_cap+3.23000e-05'
+ cm5m2dsw = '-9.43750e-13*ic_cap*ic_cap+-4.75000e-13*ic_cap+1.07000e-10'
+ cm5m2f = '-2.71875e-07*ic_cap*ic_cap+-1.62500e-07*ic_cap+2.91000e-05'
+ cm5m2fsw = '-9.37500e-13*ic_cap*ic_cap+-4.75000e-13*ic_cap+1.07000e-10'
+ cm5m2l1 = '-5.28125e-07*ic_cap*ic_cap+-3.37500e-07*ic_cap+4.85000e-05'
+ cm5m2l1sw = '-8.65625e-13*ic_cap*ic_cap+-5.37500e-13*ic_cap+1.05000e-10'
+ cm5m2m1 = '-2.70312e-06*ic_cap*ic_cap+-1.31250e-06*ic_cap+1.39000e-04'
+ cm5m2m1sw = '-8.40625e-13*ic_cap*ic_cap+-3.87500e-13*ic_cap+1.03000e-10'
+ cm5m2p1 = '-3.90625e-07*ic_cap*ic_cap+-2.37500e-07*ic_cap+3.62000e-05'
+ cm5m2p1sw = '-9.46875e-13*ic_cap*ic_cap+-4.62500e-13*ic_cap+1.07000e-10'
+ cm5m2sw = '-4.84375e-13*ic_cap*ic_cap+-3.12500e-13*ic_cap+7.74000e-11'
+ cm5m3 = '-1.75000e-07*ic_cap*ic_cap+-1.00000e-07*ic_cap+1.99000e-05'
+ cm5m3d = '-3.09375e-07*ic_cap*ic_cap+-1.87500e-07*ic_cap+3.40000e-05'
+ cm5m3dsw = '-7.59375e-13*ic_cap*ic_cap+-4.37500e-13*ic_cap+1.06000e-10'
+ cm5m3f = '-3.00000e-07*ic_cap*ic_cap+-1.75000e-07*ic_cap+3.24000e-05'
+ cm5m3fsw = '-7.50000e-13*ic_cap*ic_cap+-4.25000e-13*ic_cap+1.06000e-10'
+ cm5m3l1 = '-3.81250e-07*ic_cap*ic_cap+-2.25000e-07*ic_cap+4.00000e-05'
+ cm5m3l1sw = '-7.21875e-13*ic_cap*ic_cap+-4.37500e-13*ic_cap+1.05000e-10'
+ cm5m3m1 = '-5.62500e-07*ic_cap*ic_cap+-3.25000e-07*ic_cap+5.27000e-05'
+ cm5m3m1sw = '-7.65625e-13*ic_cap*ic_cap+-4.12500e-13*ic_cap+1.05000e-10'
+ cm5m3m2 = '-1.42500e-06*ic_cap*ic_cap+-7.75000e-07*ic_cap+1.02000e-04'
+ cm5m3m2sw = '-7.12500e-13*ic_cap*ic_cap+-3.75000e-13*ic_cap+1.03000e-10'
+ cm5m3p1 = '-3.46875e-07*ic_cap*ic_cap+-2.12500e-07*ic_cap+3.57000e-05'
+ cm5m3p1sw = '-7.62500e-13*ic_cap*ic_cap+-4.25000e-13*ic_cap+1.06000e-10'
+ cm5m3sw = '-5.03125e-13*ic_cap*ic_cap+-3.37500e-13*ic_cap+7.76000e-11'
+ cm5m4 = '-1.09687e-06*ic_cap*ic_cap+-5.37500e-07*ic_cap+6.84000e-05'
+ cm5m4d = '-1.17812e-06*ic_cap*ic_cap+-5.87500e-07*ic_cap+7.78000e-05'
+ cm5m4dsw = '-7.09375e-13*ic_cap*ic_cap+-3.87500e-13*ic_cap+1.04000e-10'
+ cm5m4f = '-1.17188e-06*ic_cap*ic_cap+-5.87500e-07*ic_cap+7.70000e-05'
+ cm5m4fsw = '-7.06250e-13*ic_cap*ic_cap+-3.75000e-13*ic_cap+1.04000e-10'
+ cm5m4l1 = '-1.19375e-06*ic_cap*ic_cap+-6.00000e-07*ic_cap+8.01000e-05'
+ cm5m4l1sw = '-7.28125e-13*ic_cap*ic_cap+-4.12500e-13*ic_cap+1.04000e-10'
+ cm5m4m1 = '-1.22500e-06*ic_cap*ic_cap+-6.25000e-07*ic_cap+8.35000e-05'
+ cm5m4m1sw = '-6.75000e-13*ic_cap*ic_cap+-3.75000e-13*ic_cap+1.03000e-10'
+ cm5m4m2 = '-1.26563e-06*ic_cap*ic_cap+-6.37500e-07*ic_cap+8.92000e-05'
+ cm5m4m2sw = '-7.03125e-13*ic_cap*ic_cap+-3.87500e-13*ic_cap+1.03000e-10'
+ cm5m4m3 = '-2.84375e-06*ic_cap*ic_cap+-1.37500e-06*ic_cap+1.57000e-04'
+ cm5m4m3sw = '-6.25000e-13*ic_cap*ic_cap+-3.50000e-13*ic_cap+1.00000e-10'
+ cm5m4p1 = '-1.18750e-06*ic_cap*ic_cap+-6.00000e-07*ic_cap+7.85000e-05'
+ cm5m4p1sw = '-7.18750e-13*ic_cap*ic_cap+-4.00000e-13*ic_cap+1.04000e-10'
+ cm5m4sw = '-7.28125e-13*ic_cap*ic_cap+-4.37500e-13*ic_cap+8.87000e-11'
+ cm5p1 = '-5.71875e-08*ic_cap*ic_cap+-3.62500e-08*ic_cap+7.26000e-06'
+ cm5p1f = '-1.44375e-06*ic_cap*ic_cap+-8.25000e-07*ic_cap+1.13000e-04'
+ cm5p1fsw = '-6.50000e-13*ic_cap*ic_cap+-3.75000e-13*ic_cap+8.61000e-11'
+ cm5p1sw = '-4.81250e-13*ic_cap*ic_cap+-3.25000e-13*ic_cap+7.82000e-11'
+ cnwvc2_cdepmult = '-1.25000e-02*cnwvc+1.00000e+00'
+ cnwvc2_cintmult = '-1.25000e-02*cnwvc+1.00000e+00'
+ cnwvc2_dlc = '-2.50000e-03*cnwvc'
+ cnwvc2_dld = '-1.50000e-04*cnwvc'
+ cnwvc2_dwc = '-5.00000e-03*cnwvc'
+ cnwvc2_tox = '1.32732e-02*cnwvc*cnwvc+5.84020e-01*cnwvc+4.24742e+01'
+ cnwvc2_vt1 = '1.85000e-02*cnwvc+2.00000e-01'
+ cnwvc2_vt2 = '1.85000e-02*cnwvc+3.30000e-01'
+ cnwvc2_vtr = '1.85000e-02*cnwvc+1.40000e-01'
+ cnwvc_cdepmult = '-2.50000e-02*cnwvc+1.00000e+00'
+ cnwvc_cintmult = '-1.25000e-02*cnwvc+1.00000e+00'
+ cnwvc_dlc = '-2.50000e-03*poly_cd'
+ cnwvc_dld = '-2.00000e-04*cnwvc'
+ cnwvc_dwc = '-5.00000e-03*cnwvc'
+ cnwvc_tox = '1.59937e-02*cnwvc*cnwvc+5.75774e-01*cnwvc+4.26499e+01'
+ cnwvc_vt1 = '2.80000e-02*lvp_threshold+3.33300e-01'
+ cnwvc_vt2 = '2.80000e-02*lvp_threshold+2.38095e-01'
+ cnwvc_vtr = '2.80000e-02*lvp_threshold+1.60000e-01'
+ cp1f = '-1.40313e-06*ic_cap*ic_cap+-7.87500e-07*ic_cap+1.06000e-04'
+ cp1fsw = '-6.62500e-13*ic_cap*ic_cap+-3.75000e-13*ic_cap+8.64000e-11'
+ cpl2s_vpp = '6.87500e-03*ic_cap*ic_cap+8.75000e-02*ic_cap+1.00000e+00'
+ cpl2s_vpp0p4shield = '8.62813e-03*ic_cap*ic_cap+9.67375e-02*ic_cap+1.00000e+00'
+ cpmimc = '4.00000e-17*mim+1.90000e-16'
+ crdld = '-2.28125e-08*ic_cap*ic_cap+-1.37500e-08*ic_cap+2.63000e-06'
+ crdldsw = '-5.65625e-13*ic_cap*ic_cap+-3.37500e-13*ic_cap+5.75000e-11'
+ crdlf = '-2.28125e-08*ic_cap*ic_cap+-1.37500e-08*ic_cap+2.57000e-06'
+ crdlfsw = '-5.62500e-13*ic_cap*ic_cap+-3.50000e-13*ic_cap+5.75000e-11'
+ crdll1 = '-2.43750e-08*ic_cap*ic_cap+-1.50000e-08*ic_cap+2.78000e-06'
+ crdll1d = '-5.68750e-07*ic_cap*ic_cap+-3.25000e-07*ic_cap+5.80000e-05'
+ crdll1dsw = '-7.93750e-13*ic_cap*ic_cap+-5.25000e-13*ic_cap+8.22000e-11'
+ crdll1f = '-4.40625e-07*ic_cap*ic_cap+-2.37500e-07*ic_cap+3.97000e-05'
+ crdll1fsw = '-8.06250e-13*ic_cap*ic_cap+-5.25000e-13*ic_cap+8.30000e-11'
+ crdll1p1 = '-1.67813e-06*ic_cap*ic_cap+-8.12500e-07*ic_cap+9.69000e-05'
+ crdll1p1sw = '-7.62500e-13*ic_cap*ic_cap+-5.00000e-13*ic_cap+8.12000e-11'
+ crdll1sw = '-5.62500e-13*ic_cap*ic_cap+-3.50000e-13*ic_cap+5.73000e-11'
+ crdlm1 = '-2.56250e-08*ic_cap*ic_cap+-1.50000e-08*ic_cap+2.93000e-06'
+ crdlm1d = '-3.96875e-07*ic_cap*ic_cap+-2.62500e-07*ic_cap+3.65000e-05'
+ crdlm1dsw = '-9.59375e-13*ic_cap*ic_cap+-5.12500e-13*ic_cap+1.07000e-10'
+ crdlm1f = '-3.25000e-07*ic_cap*ic_cap+-2.00000e-07*ic_cap+2.87000e-05'
+ crdlm1fsw = '-9.43750e-13*ic_cap*ic_cap+-5.25000e-13*ic_cap+1.07000e-10'
+ crdlm1l1 = '-2.01250e-06*ic_cap*ic_cap+-1.27500e-06*ic_cap+1.17000e-04'
+ crdlm1l1sw = '-8.09375e-13*ic_cap*ic_cap+-4.62500e-13*ic_cap+1.03000e-10'
+ crdlm1p1 = '-7.09375e-07*ic_cap*ic_cap+-4.12500e-07*ic_cap+4.78000e-05'
+ crdlm1p1sw = '-9.15625e-13*ic_cap*ic_cap+-5.12500e-13*ic_cap+1.06000e-10'
+ crdlm1sw = '-5.59375e-13*ic_cap*ic_cap+-3.37500e-13*ic_cap+5.71000e-11'
+ crdlm2 = '-2.71875e-08*ic_cap*ic_cap+-1.62500e-08*ic_cap+3.10000e-06'
+ crdlm2d = '-2.40625e-07*ic_cap*ic_cap+-1.62500e-07*ic_cap+2.39000e-05'
+ crdlm2dsw = '-9.40625e-13*ic_cap*ic_cap+-5.37500e-13*ic_cap+1.07000e-10'
+ crdlm2f = '-2.15625e-07*ic_cap*ic_cap+-1.37500e-07*ic_cap+2.06000e-05'
+ crdlm2fsw = '-9.34375e-13*ic_cap*ic_cap+-5.37500e-13*ic_cap+1.07000e-10'
+ crdlm2l1 = '-4.78125e-07*ic_cap*ic_cap+-3.12500e-07*ic_cap+4.01000e-05'
+ crdlm2l1sw = '-9.09375e-13*ic_cap*ic_cap+-5.37500e-13*ic_cap+1.06000e-10'
+ crdlm2m1 = '-2.68125e-06*ic_cap*ic_cap+-1.27500e-06*ic_cap+1.31000e-04'
+ crdlm2m1sw = '-8.12500e-13*ic_cap*ic_cap+-4.25000e-13*ic_cap+1.03000e-10'
+ crdlm2p1 = '-3.40625e-07*ic_cap*ic_cap+-2.12500e-07*ic_cap+2.78000e-05'
+ crdlm2p1sw = '-9.53125e-13*ic_cap*ic_cap+-5.37500e-13*ic_cap+1.07000e-10'
+ crdlm2sw = '-5.59375e-13*ic_cap*ic_cap+-3.37500e-13*ic_cap+5.70000e-11'
+ crdlm3 = '-3.25000e-08*ic_cap*ic_cap+-2.00000e-08*ic_cap+3.50000e-06'
+ crdlm3d = '-1.71875e-07*ic_cap*ic_cap+-1.12500e-07*ic_cap+1.77000e-05'
+ crdlm3dsw = '-7.84375e-13*ic_cap*ic_cap+-4.37500e-13*ic_cap+1.08000e-10'
+ crdlm3f = '-1.62500e-07*ic_cap*ic_cap+-1.00000e-07*ic_cap+1.61000e-05'
+ crdlm3fsw = '-7.84375e-13*ic_cap*ic_cap+-4.37500e-13*ic_cap+1.08000e-10'
+ crdlm3l1 = '-2.43750e-07*ic_cap*ic_cap+-1.50000e-07*ic_cap+2.37000e-05'
+ crdlm3l1sw = '-7.53125e-13*ic_cap*ic_cap+-4.37500e-13*ic_cap+1.07000e-10'
+ crdlm3m1 = '-4.21875e-07*ic_cap*ic_cap+-2.37500e-07*ic_cap+3.64000e-05'
+ crdlm3m1sw = '-7.37500e-13*ic_cap*ic_cap+-4.50000e-13*ic_cap+1.06000e-10'
+ crdlm3m2 = '-1.28750e-06*ic_cap*ic_cap+-7.00000e-07*ic_cap+8.57000e-05'
+ crdlm3m2sw = '-7.43750e-13*ic_cap*ic_cap+-4.25000e-13*ic_cap+1.05000e-10'
+ crdlm3p1 = '-2.12500e-07*ic_cap*ic_cap+-1.25000e-07*ic_cap+1.94000e-05'
+ crdlm3p1sw = '-7.28125e-13*ic_cap*ic_cap+-4.37500e-13*ic_cap+1.07000e-10'
+ crdlm3sw = '-5.59375e-13*ic_cap*ic_cap+-3.37500e-13*ic_cap+5.68000e-11'
+ crdlm4 = '-3.90625e-08*ic_cap*ic_cap+-2.37500e-08*ic_cap+4.00000e-06'
+ crdlm4d = '-1.18750e-07*ic_cap*ic_cap+-7.50000e-08*ic_cap+1.34000e-05'
+ crdlm4dsw = '-8.18750e-13*ic_cap*ic_cap+-4.25000e-13*ic_cap+1.09000e-10'
+ crdlm4f = '-1.15625e-07*ic_cap*ic_cap+-6.25000e-08*ic_cap+1.27000e-05'
+ crdlm4fsw = '-8.15625e-13*ic_cap*ic_cap+-4.37500e-13*ic_cap+1.09000e-10'
+ crdlm4l1 = '-1.34375e-07*ic_cap*ic_cap+-8.75000e-08*ic_cap+1.57000e-05'
+ crdlm4l1sw = '-8.28125e-13*ic_cap*ic_cap+-4.37500e-13*ic_cap+1.09000e-10'
+ crdlm4m1 = '-1.68750e-07*ic_cap*ic_cap+-1.00000e-07*ic_cap+1.91000e-05'
+ crdlm4m1sw = '-7.87500e-13*ic_cap*ic_cap+-4.50000e-13*ic_cap+1.08000e-10'
+ crdlm4m2 = '-2.12500e-07*ic_cap*ic_cap+-1.25000e-07*ic_cap+2.49000e-05'
+ crdlm4m2sw = '-8.18750e-13*ic_cap*ic_cap+-4.75000e-13*ic_cap+1.08000e-10'
+ crdlm4m3 = '-1.75938e-06*ic_cap*ic_cap+-8.62500e-07*ic_cap+9.25000e-05'
+ crdlm4m3sw = '-7.40625e-13*ic_cap*ic_cap+-4.37500e-13*ic_cap+1.05000e-10'
+ crdlm4p1 = '-1.31250e-07*ic_cap*ic_cap+-7.50000e-08*ic_cap+1.41000e-05'
+ crdlm4p1sw = '-8.21875e-13*ic_cap*ic_cap+-4.37500e-13*ic_cap+1.09000e-10'
+ crdlm4sw = '-5.53125e-13*ic_cap*ic_cap+-3.37500e-13*ic_cap+5.66000e-11'
+ crdlm5 = '-6.31250e-08*ic_cap*ic_cap+-3.75000e-08*ic_cap+5.44000e-06'
+ crdlm5d = '-1.15625e-07*ic_cap*ic_cap+-6.25000e-08*ic_cap+1.24000e-05'
+ crdlm5dsw = '-4.62500e-13*ic_cap*ic_cap+-3.00000e-13*ic_cap+7.59000e-11'
+ crdlm5f = '-1.16875e-07*ic_cap*ic_cap+-6.75000e-08*ic_cap+1.20000e-05'
+ crdlm5fsw = '-4.56250e-13*ic_cap*ic_cap+-3.00000e-13*ic_cap+7.60000e-11'
+ crdlm5l1 = '-1.18750e-07*ic_cap*ic_cap+-7.50000e-08*ic_cap+1.35000e-05'
+ crdlm5l1sw = '-4.53125e-13*ic_cap*ic_cap+-3.12500e-13*ic_cap+7.55000e-11'
+ crdlm5m1 = '-1.31250e-07*ic_cap*ic_cap+-7.50000e-08*ic_cap+1.50000e-05'
+ crdlm5m1sw = '-4.53125e-13*ic_cap*ic_cap+-3.12500e-13*ic_cap+7.52000e-11'
+ crdlm5m2 = '-1.40625e-07*ic_cap*ic_cap+-8.75000e-08*ic_cap+1.70000e-05'
+ crdlm5m2sw = '-4.56250e-13*ic_cap*ic_cap+-3.00000e-13*ic_cap+7.49000e-11'
+ crdlm5m3 = '-2.34375e-07*ic_cap*ic_cap+-1.37500e-07*ic_cap+2.53000e-05'
+ crdlm5m3sw = '-4.68750e-13*ic_cap*ic_cap+-3.00000e-13*ic_cap+7.50000e-11'
+ crdlm5m4 = '-1.16250e-06*ic_cap*ic_cap+-5.75000e-07*ic_cap+7.39000e-05'
+ crdlm5m4sw = '-6.90625e-13*ic_cap*ic_cap+-4.12500e-13*ic_cap+8.61000e-11'
+ crdlm5p1 = '-1.18750e-07*ic_cap*ic_cap+-7.50000e-08*ic_cap+1.27000e-05'
+ crdlm5p1sw = '-4.56250e-13*ic_cap*ic_cap+-3.00000e-13*ic_cap+7.57000e-11'
+ crdlm5sw = '-5.56250e-13*ic_cap*ic_cap+-3.50000e-13*ic_cap+5.68000e-11'
+ crdlp1 = '-2.37500e-08*ic_cap*ic_cap+-1.50000e-08*ic_cap+2.68000e-06'
+ crdlp1f = '-1.44688e-06*ic_cap*ic_cap+-7.87500e-07*ic_cap+1.09000e-04'
+ crdlp1fsw = '-6.56250e-13*ic_cap*ic_cap+-3.75000e-13*ic_cap+8.63000e-11'
+ crdlp1sw = '-5.62500e-13*ic_cap*ic_cap+-3.50000e-13*ic_cap+5.74000e-11'
+ crpf_precision = '6.84375e-07*ic_res*ic_res+9.01250e-06*ic_res+1.06000e-04'
+ crpfsw_precision_16_2 = '9.37500e-14*ic_res*ic_res+1.90000e-12*ic_res+6.97000e-11'
+ crpfsw_precision_1_1 = '8.12500e-14*ic_res*ic_res+1.65000e-12*ic_res+5.04000e-11'
+ crpfsw_precision_2_1 = '8.43750e-14*ic_res*ic_res+1.66250e-12*ic_res+5.39000e-11'
+ crpfsw_precision_4_1 = '8.75000e-14*ic_res*ic_res+1.72500e-12*ic_res+5.83000e-11'
+ crpfsw_precision_8_2 = '9.06250e-14*ic_res*ic_res+1.78750e-12*ic_res+6.36000e-11'
+ cvpp2_nhvnative10x4_cor = '-6.25000e-05*ic_cap*ic_cap+-3.42500e-02*ic_cap+1.00000e+00'
+ cvpp2_nhvnative10x4_sub = '1.10250e-16*ic_cap*ic_cap+-1.42900e-15*ic_cap+4.82000e-15'
+ cvpp2_phv5x4_cor = '-6.25000e-05*ic_cap*ic_cap+-3.42500e-02*ic_cap+1.00000e+00'
+ cvpp2_phv5x4_sub = '1.10250e-16*ic_cap*ic_cap+-1.42900e-15*ic_cap+4.82000e-15'
+ cvpp3_cor = '7.50000e-02*ic_cap+1.00000e+00'
+ cvpp4_cor = '7.50000e-02*ic_cap+1.00000e+00'
+ cvpp5_cor = '7.50000e-02*ic_cap+1.00000e+00'
+ cvpp_cor = '-6.25000e-05*ic_cap*ic_cap+3.42500e-02*ic_cap+1.00000e+00'
+ dkbfnpn1x1 = '1.40312e-04*sky130_fd_pr__npn_05v5_all*sky130_fd_pr__npn_05v5_all+-1.28636e-01*sky130_fd_pr__npn_05v5_all+9.85010e-01'
+ dkbfnpn1x2 = '1.40000e-04*sky130_fd_pr__npn_05v5_all*sky130_fd_pr__npn_05v5_all+-1.26493e-01*sky130_fd_pr__npn_05v5_all+9.67590e-01'
+ dkbfnpnpolyhv = '1.25000e-04*sky130_fd_pr__npn_05v5_all*sky130_fd_pr__npn_05v5_all+-1.30750e-01*sky130_fd_pr__npn_05v5_all+1.00000e+00'
+ dkbfpp = '1.54062e-04*pnp_05v5_W0p68L0p68*pnp_05v5_W0p68L0p68+-1.15849e-01*pnp_05v5_W0p68L0p68+9.51540e-01'
+ dkbfpp5x = '-1.19375e-04*pnp_05v5_W0p68L0p68*pnp_05v5_W0p68L0p68+-1.66327e-01*pnp_05v5_W0p68L0p68+1.12880e+00'
+ dkisnpn1x1 = '4.00625e-03*sky130_fd_pr__npn_05v5_all*sky130_fd_pr__npn_05v5_all+-8.62425e-02*sky130_fd_pr__npn_05v5_all+8.79130e-01'
+ dkisnpn1x2 = '4.10969e-03*sky130_fd_pr__npn_05v5_all*sky130_fd_pr__npn_05v5_all+-8.80613e-02*sky130_fd_pr__npn_05v5_all+9.09500e-01'
+ dkisnpnpolyhv = '8.78125e-03*sky130_fd_pr__npn_05v5_all*sky130_fd_pr__npn_05v5_all+-1.37375e-01*sky130_fd_pr__npn_05v5_all+1.00000e+00'
+ dkispp = '1.20531e-03*pnp_05v5_W0p68L0p68*pnp_05v5_W0p68L0p68+-5.95037e-02*pnp_05v5_W0p68L0p68+9.28400e-01'
+ dkispp5x = '-3.81875e-04*pnp_05v5_W0p68L0p68*pnp_05v5_W0p68L0p68+-5.29775e-02*pnp_05v5_W0p68L0p68+1.00460e+00'
+ sky130_fd_pr__model__parasitic__diode_ps2dn__ajunction_mult = '-4.75000e-04*well_diode*well_diode+6.70500e-02*well_diode+9.85800e-01'
+ sky130_fd_pr__model__parasitic__diode_ps2dn__pjunction_mult = '3.98750e-04*well_diode*well_diode+7.84800e-02*well_diode+1.01160e+00'
+ sky130_fd_pr__model__parasitic__diode_pw2dn__ajunction_mult = '1.87500e-04*well_diode*well_diode+7.37500e-02*well_diode+9.82000e-01'
+ sky130_fd_pr__model__parasitic__diode_pw2dn__pjunction_mult = '-7.79688e-04*well_diode*well_diode+1.78588e-02*well_diode+9.63040e-01'
+ sky130_fd_pr__special_nfet_pass_flash__ajunction_mult = '9.37500e-07*lvn_diode*lvn_diode+3.87638e-02*lvn_diode+9.95430e-01'
+ sky130_fd_pr__special_nfet_pass_flash__dlc_diff = '-3.03188e-09*poly_cd'
+ sky130_fd_pr__special_nfet_pass_flash__dwc_diff = '5.63000e-09*diff_cd'
+ sky130_fd_pr__special_nfet_pass_flash__kt1_diff_1 = '-1.06270e-02*lvn_subvt*lvn_subvt+1.13538e-02*lvn_subvt+3.82270e-02'
+ sky130_fd_pr__special_nfet_pass_flash__lint_diff = '-3.03188e-09*poly_cd'
+ sky130_fd_pr__special_nfet_pass_flash__nfactor_diff_0 = '-7.91375e-03*lvn_subvt*lvn_subvt+3.16550e-02*lvn_subvt'
+ sky130_fd_pr__special_nfet_pass_flash__nfactor_diff_1 = '1.41651e-02*lvn_subvt*lvn_subvt+8.47347e-02*lvn_subvt+1.41380e-01'
+ sky130_fd_pr__special_nfet_pass_flash__overlap_mult = '1.18750e-04*lvtox*lvtox+2.44075e-02*lvtox+8.98050e-01'
+ sky130_fd_pr__special_nfet_pass_flash__pjunction_mult = '-9.37500e-07*lvn_diode*lvn_diode+3.97287e-02*lvn_diode+1.02040e+00'
+ sky130_fd_pr__special_nfet_pass_flash__tox_mult = '9.12500e-03*lvtox+1.00000e+00'
+ sky130_fd_pr__special_nfet_pass_flash__u0_diff_0 = '-1.24384e-05*lvn_mobility*lvn_mobility+8.14504e-04*lvn_mobility+2.75840e-03'
+ sky130_fd_pr__special_nfet_pass_flash__u0_diff_1 = '-1.68563e-04*lvn_mobility*lvn_mobility+1.84207e-03*lvn_mobility+1.29560e-03'
+ sky130_fd_pr__special_nfet_pass_flash__voff_diff_0 = '3.09406e-03*lvn_subvt*lvn_subvt+-1.23763e-02*lvn_subvt'
+ sky130_fd_pr__special_nfet_pass_flash__voff_diff_1 = '3.10416e-03*lvn_subvt*lvn_subvt+1.24166e-02*lvn_subvt'
+ sky130_fd_pr__special_nfet_pass_flash__vsat_diff_0 = '1.10588e+03*lvn_saturation*lvn_saturation+9.76162e+03*lvn_saturation+3.85540e+03'
+ sky130_fd_pr__special_nfet_pass_flash__vsat_diff_1 = '-6.14031e+02*lvn_saturation*lvn_saturation+3.55288e+03*lvn_saturation+1.36790e+04'
+ sky130_fd_pr__special_nfet_pass_flash__vth0_diff_0 = '-2.37156e-04*lvn_threshold*lvn_threshold+5.41889e-02*lvn_threshold+-1.56630e-01'
+ sky130_fd_pr__special_nfet_pass_flash__vth0_diff_1 = '-3.54442e-03*lvn_threshold*lvn_threshold+4.54875e-02*lvn_threshold+-5.70930e-03'
+ sky130_fd_pr__special_nfet_pass_flash__wint_diff = '5.63000e-09*diff_cd'
+ sky130_fd_pr__res_high_po__var_mult = '1.25000e+00*ic_res'
+ sky130_fd_pr__res_high_po__var = '1.25000e+00*ic_res'
+ sky130_fd_pr__res_xhigh_po__var_mult = '1.25000e+00*ic_res'
+ mcl1d_ca_w_0_170_s_0_180 = '-5.50000e-07*ic_cap*ic_cap+-3.00000e-07*ic_cap+5.53000e-05'
+ mcl1d_ca_w_0_170_s_0_225 = '-5.50000e-07*ic_cap*ic_cap+-3.00000e-07*ic_cap+5.53000e-05'
+ mcl1d_ca_w_0_170_s_0_270 = '-5.50000e-07*ic_cap*ic_cap+-3.00000e-07*ic_cap+5.53000e-05'
+ mcl1d_ca_w_0_170_s_0_360 = '-5.50000e-07*ic_cap*ic_cap+-3.00000e-07*ic_cap+5.53000e-05'
+ mcl1d_ca_w_0_170_s_0_450 = '-5.50000e-07*ic_cap*ic_cap+-3.00000e-07*ic_cap+5.53000e-05'
+ mcl1d_ca_w_0_170_s_0_540 = '-5.50000e-07*ic_cap*ic_cap+-3.00000e-07*ic_cap+5.53000e-05'
+ mcl1d_ca_w_0_170_s_0_720 = '-5.50000e-07*ic_cap*ic_cap+-3.00000e-07*ic_cap+5.53000e-05'
+ mcl1d_ca_w_0_170_s_1_080 = '-5.50000e-07*ic_cap*ic_cap+-3.00000e-07*ic_cap+5.53000e-05'
+ mcl1d_ca_w_0_170_s_1_980 = '-5.50000e-07*ic_cap*ic_cap+-3.00000e-07*ic_cap+5.53000e-05'
+ mcl1d_ca_w_0_170_s_4_500 = '-5.50000e-07*ic_cap*ic_cap+-3.00000e-07*ic_cap+5.53000e-05'
+ mcl1d_ca_w_1_360_s_0_180 = '-5.50000e-07*ic_cap*ic_cap+-3.00000e-07*ic_cap+5.53000e-05'
+ mcl1d_ca_w_1_360_s_0_225 = '-5.50000e-07*ic_cap*ic_cap+-3.00000e-07*ic_cap+5.53000e-05'
+ mcl1d_ca_w_1_360_s_0_270 = '-5.50000e-07*ic_cap*ic_cap+-3.00000e-07*ic_cap+5.53000e-05'
+ mcl1d_ca_w_1_360_s_0_360 = '-5.50000e-07*ic_cap*ic_cap+-3.00000e-07*ic_cap+5.53000e-05'
+ mcl1d_ca_w_1_360_s_0_450 = '-5.50000e-07*ic_cap*ic_cap+-3.00000e-07*ic_cap+5.53000e-05'
+ mcl1d_ca_w_1_360_s_0_540 = '-5.50000e-07*ic_cap*ic_cap+-3.00000e-07*ic_cap+5.53000e-05'
+ mcl1d_ca_w_1_360_s_0_720 = '-5.50000e-07*ic_cap*ic_cap+-3.00000e-07*ic_cap+5.53000e-05'
+ mcl1d_ca_w_1_360_s_1_080 = '-5.50000e-07*ic_cap*ic_cap+-3.00000e-07*ic_cap+5.53000e-05'
+ mcl1d_ca_w_1_360_s_1_980 = '-5.50000e-07*ic_cap*ic_cap+-3.00000e-07*ic_cap+5.53000e-05'
+ mcl1d_ca_w_1_360_s_4_500 = '-5.50000e-07*ic_cap*ic_cap+-3.00000e-07*ic_cap+5.53000e-05'
+ mcl1d_cc_w_0_170_s_0_180 = '-7.84375e-13*ic_cap*ic_cap+-5.12500e-13*ic_cap+7.74000e-11'
+ mcl1d_cc_w_0_170_s_0_225 = '-5.65625e-13*ic_cap*ic_cap+-3.87500e-13*ic_cap+6.56000e-11'
+ mcl1d_cc_w_0_170_s_0_270 = '-4.31250e-13*ic_cap*ic_cap+-3.00000e-13*ic_cap+5.78000e-11'
+ mcl1d_cc_w_0_170_s_0_360 = '-2.90625e-13*ic_cap*ic_cap+-2.12500e-13*ic_cap+4.66000e-11'
+ mcl1d_cc_w_0_170_s_0_450 = '-1.96875e-13*ic_cap*ic_cap+-1.62500e-13*ic_cap+3.96000e-11'
+ mcl1d_cc_w_0_170_s_0_540 = '-1.43750e-13*ic_cap*ic_cap+-1.25000e-13*ic_cap+3.39000e-11'
+ mcl1d_cc_w_0_170_s_0_720 = '-8.12500e-14*ic_cap*ic_cap+-7.50000e-14*ic_cap+2.64000e-11'
+ mcl1d_cc_w_0_170_s_1_080 = '-1.56250e-14*ic_cap*ic_cap+-3.75000e-14*ic_cap+1.75000e-11'
+ mcl1d_cc_w_0_170_s_1_980 = '1.62500e-14*ic_cap*ic_cap+8.42000e-12'
+ mcl1d_cc_w_0_170_s_4_500 = '1.06250e-14*ic_cap*ic_cap+5.00000e-15*ic_cap+2.28000e-12'
+ mcl1d_cc_w_1_360_s_0_180 = '-7.06250e-13*ic_cap*ic_cap+-4.50000e-13*ic_cap+9.72000e-11'
+ mcl1d_cc_w_1_360_s_0_225 = '-4.96875e-13*ic_cap*ic_cap+-3.37500e-13*ic_cap+8.44000e-11'
+ mcl1d_cc_w_1_360_s_0_270 = '-3.65625e-13*ic_cap*ic_cap+-2.62500e-13*ic_cap+7.51000e-11'
+ mcl1d_cc_w_1_360_s_0_360 = '-2.21875e-13*ic_cap*ic_cap+-1.62500e-13*ic_cap+6.24000e-11'
+ mcl1d_cc_w_1_360_s_0_450 = '-1.40625e-13*ic_cap*ic_cap+-1.12500e-13*ic_cap+5.39000e-11'
+ mcl1d_cc_w_1_360_s_0_540 = '-9.37500e-14*ic_cap*ic_cap+-1.00000e-13*ic_cap+4.76000e-11'
+ mcl1d_cc_w_1_360_s_0_720 = '-3.43750e-14*ic_cap*ic_cap+-3.75000e-14*ic_cap+3.87000e-11'
+ mcl1d_cc_w_1_360_s_1_080 = '1.56250e-14*ic_cap*ic_cap+-1.25000e-14*ic_cap+2.80000e-11'
+ mcl1d_cc_w_1_360_s_1_980 = '3.43750e-14*ic_cap*ic_cap+1.25000e-14*ic_cap+1.55000e-11'
+ mcl1d_cc_w_1_360_s_4_500 = '2.34375e-14*ic_cap*ic_cap+6.25000e-15*ic_cap+5.35000e-12'
+ mcl1d_cf_w_0_170_s_0_180 = '-8.12500e-15*ic_cap*ic_cap+-2.50000e-15*ic_cap+4.83000e-12'
+ mcl1d_cf_w_0_170_s_0_225 = '-1.96875e-14*ic_cap*ic_cap+-1.12500e-14*ic_cap+5.98000e-12'
+ mcl1d_cf_w_0_170_s_0_270 = '-3.09375e-14*ic_cap*ic_cap+-1.62500e-14*ic_cap+7.08000e-12'
+ mcl1d_cf_w_0_170_s_0_360 = '-4.62500e-14*ic_cap*ic_cap+-2.75000e-14*ic_cap+9.37000e-12'
+ mcl1d_cf_w_0_170_s_0_450 = '-7.31250e-14*ic_cap*ic_cap+-4.25000e-14*ic_cap+1.13000e-11'
+ mcl1d_cf_w_0_170_s_0_540 = '-9.37500e-14*ic_cap*ic_cap+-5.00000e-14*ic_cap+1.35000e-11'
+ mcl1d_cf_w_0_170_s_0_720 = '-1.21875e-13*ic_cap*ic_cap+-6.25000e-14*ic_cap+1.70000e-11'
+ mcl1d_cf_w_0_170_s_1_080 = '-1.62500e-13*ic_cap*ic_cap+-1.00000e-13*ic_cap+2.25000e-11'
+ mcl1d_cf_w_0_170_s_1_980 = '-2.06250e-13*ic_cap*ic_cap+-1.25000e-13*ic_cap+3.00000e-11'
+ mcl1d_cf_w_0_170_s_4_500 = '-2.03125e-13*ic_cap*ic_cap+-1.37500e-13*ic_cap+3.59000e-11'
+ mcl1d_cf_w_1_360_s_0_180 = '-8.12500e-15*ic_cap*ic_cap+-2.50000e-15*ic_cap+4.83000e-12'
+ mcl1d_cf_w_1_360_s_0_225 = '-1.96875e-14*ic_cap*ic_cap+-8.75000e-15*ic_cap+5.98000e-12'
+ mcl1d_cf_w_1_360_s_0_270 = '-3.06250e-14*ic_cap*ic_cap+-1.50000e-14*ic_cap+7.11000e-12'
+ mcl1d_cf_w_1_360_s_0_360 = '-5.18750e-14*ic_cap*ic_cap+-2.75000e-14*ic_cap+9.29000e-12'
+ mcl1d_cf_w_1_360_s_0_450 = '-7.18750e-14*ic_cap*ic_cap+-3.75000e-14*ic_cap+1.14000e-11'
+ mcl1d_cf_w_1_360_s_0_540 = '-8.75000e-14*ic_cap*ic_cap+-5.00000e-14*ic_cap+1.33000e-11'
+ mcl1d_cf_w_1_360_s_0_720 = '-1.21875e-13*ic_cap*ic_cap+-6.25000e-14*ic_cap+1.70000e-11'
+ mcl1d_cf_w_1_360_s_1_080 = '-1.62500e-13*ic_cap*ic_cap+-1.00000e-13*ic_cap+2.29000e-11'
+ mcl1d_cf_w_1_360_s_1_980 = '-2.03125e-13*ic_cap*ic_cap+-1.12500e-13*ic_cap+3.25000e-11'
+ mcl1d_cf_w_1_360_s_4_500 = '-2.00000e-13*ic_cap*ic_cap+-1.25000e-13*ic_cap+4.19000e-11'
+ mcl1f_ca_w_0_170_s_0_180 = '-4.15625e-07*ic_cap*ic_cap+-2.37500e-07*ic_cap+3.69000e-05'
+ mcl1f_ca_w_0_170_s_0_225 = '-4.15625e-07*ic_cap*ic_cap+-2.37500e-07*ic_cap+3.69000e-05'
+ mcl1f_ca_w_0_170_s_0_270 = '-4.15625e-07*ic_cap*ic_cap+-2.37500e-07*ic_cap+3.69000e-05'
+ mcl1f_ca_w_0_170_s_0_360 = '-4.15625e-07*ic_cap*ic_cap+-2.37500e-07*ic_cap+3.69000e-05'
+ mcl1f_ca_w_0_170_s_0_450 = '-4.15625e-07*ic_cap*ic_cap+-2.37500e-07*ic_cap+3.69000e-05'
+ mcl1f_ca_w_0_170_s_0_540 = '-4.15625e-07*ic_cap*ic_cap+-2.37500e-07*ic_cap+3.69000e-05'
+ mcl1f_ca_w_0_170_s_0_720 = '-4.15625e-07*ic_cap*ic_cap+-2.37500e-07*ic_cap+3.69000e-05'
+ mcl1f_ca_w_0_170_s_1_080 = '-4.15625e-07*ic_cap*ic_cap+-2.37500e-07*ic_cap+3.69000e-05'
+ mcl1f_ca_w_0_170_s_1_980 = '-4.15625e-07*ic_cap*ic_cap+-2.37500e-07*ic_cap+3.69000e-05'
+ mcl1f_ca_w_0_170_s_4_500 = '-4.15625e-07*ic_cap*ic_cap+-2.37500e-07*ic_cap+3.69000e-05'
+ mcl1f_ca_w_1_360_s_0_180 = '-4.15625e-07*ic_cap*ic_cap+-2.37500e-07*ic_cap+3.69000e-05'
+ mcl1f_ca_w_1_360_s_0_225 = '-4.15625e-07*ic_cap*ic_cap+-2.37500e-07*ic_cap+3.69000e-05'
+ mcl1f_ca_w_1_360_s_0_270 = '-4.15625e-07*ic_cap*ic_cap+-2.37500e-07*ic_cap+3.69000e-05'
+ mcl1f_ca_w_1_360_s_0_360 = '-4.15625e-07*ic_cap*ic_cap+-2.37500e-07*ic_cap+3.69000e-05'
+ mcl1f_ca_w_1_360_s_0_450 = '-4.15625e-07*ic_cap*ic_cap+-2.37500e-07*ic_cap+3.69000e-05'
+ mcl1f_ca_w_1_360_s_0_540 = '-4.15625e-07*ic_cap*ic_cap+-2.37500e-07*ic_cap+3.69000e-05'
+ mcl1f_ca_w_1_360_s_0_720 = '-4.15625e-07*ic_cap*ic_cap+-2.37500e-07*ic_cap+3.69000e-05'
+ mcl1f_ca_w_1_360_s_1_080 = '-4.15625e-07*ic_cap*ic_cap+-2.37500e-07*ic_cap+3.69000e-05'
+ mcl1f_ca_w_1_360_s_1_980 = '-4.15625e-07*ic_cap*ic_cap+-2.37500e-07*ic_cap+3.69000e-05'
+ mcl1f_ca_w_1_360_s_4_500 = '-4.15625e-07*ic_cap*ic_cap+-2.37500e-07*ic_cap+3.69000e-05'
+ mcl1f_cc_w_0_170_s_0_180 = '-7.93750e-13*ic_cap*ic_cap+-5.25000e-13*ic_cap+7.98000e-11'
+ mcl1f_cc_w_0_170_s_0_225 = '-5.87500e-13*ic_cap*ic_cap+-4.00000e-13*ic_cap+6.83000e-11'
+ mcl1f_cc_w_0_170_s_0_270 = '-4.50000e-13*ic_cap*ic_cap+-3.25000e-13*ic_cap+6.07000e-11'
+ mcl1f_cc_w_0_170_s_0_360 = '-3.06250e-13*ic_cap*ic_cap+-2.25000e-13*ic_cap+4.97000e-11'
+ mcl1f_cc_w_0_170_s_0_450 = '-2.09375e-13*ic_cap*ic_cap+-1.62500e-13*ic_cap+4.29000e-11'
+ mcl1f_cc_w_0_170_s_0_540 = '-1.50000e-13*ic_cap*ic_cap+-1.25000e-13*ic_cap+3.73000e-11'
+ mcl1f_cc_w_0_170_s_0_720 = '-8.75000e-14*ic_cap*ic_cap+-7.50000e-14*ic_cap+3.01000e-11'
+ mcl1f_cc_w_0_170_s_1_080 = '-1.87500e-14*ic_cap*ic_cap+-2.50000e-14*ic_cap+2.13000e-11'
+ mcl1f_cc_w_0_170_s_1_980 = '3.12500e-14*ic_cap*ic_cap+1.14000e-11'
+ mcl1f_cc_w_0_170_s_4_500 = '2.59375e-14*ic_cap*ic_cap+1.37500e-14*ic_cap+3.41000e-12'
+ mcl1f_cc_w_1_360_s_0_180 = '-7.18750e-13*ic_cap*ic_cap+-4.25000e-13*ic_cap+1.02000e-10'
+ mcl1f_cc_w_1_360_s_0_225 = '-4.84375e-13*ic_cap*ic_cap+-3.37500e-13*ic_cap+8.88000e-11'
+ mcl1f_cc_w_1_360_s_0_270 = '-3.50000e-13*ic_cap*ic_cap+-2.50000e-13*ic_cap+7.95000e-11'
+ mcl1f_cc_w_1_360_s_0_360 = '-2.06250e-13*ic_cap*ic_cap+-1.50000e-13*ic_cap+6.68000e-11'
+ mcl1f_cc_w_1_360_s_0_450 = '-1.25000e-13*ic_cap*ic_cap+-1.00000e-13*ic_cap+5.83000e-11'
+ mcl1f_cc_w_1_360_s_0_540 = '-7.81250e-14*ic_cap*ic_cap+-6.25000e-14*ic_cap+5.20000e-11'
+ mcl1f_cc_w_1_360_s_0_720 = '-2.18750e-14*ic_cap*ic_cap+-3.75000e-14*ic_cap+4.31000e-11'
+ mcl1f_cc_w_1_360_s_1_080 = '3.12500e-14*ic_cap*ic_cap+3.23000e-11'
+ mcl1f_cc_w_1_360_s_1_980 = '6.56250e-14*ic_cap*ic_cap+3.75000e-14*ic_cap+1.90000e-11'
+ mcl1f_cc_w_1_360_s_4_500 = '4.68750e-14*ic_cap*ic_cap+2.50000e-14*ic_cap+7.05000e-12'
+ mcl1f_cf_w_0_170_s_0_180 = '-1.06250e-14*ic_cap*ic_cap+-5.00000e-15*ic_cap+3.26000e-12'
+ mcl1f_cf_w_0_170_s_0_225 = '-1.87500e-14*ic_cap*ic_cap+-1.00000e-14*ic_cap+4.04000e-12'
+ mcl1f_cf_w_0_170_s_0_270 = '-2.75000e-14*ic_cap*ic_cap+-1.50000e-14*ic_cap+4.81000e-12'
+ mcl1f_cf_w_0_170_s_0_360 = '-4.03125e-14*ic_cap*ic_cap+-2.62500e-14*ic_cap+6.42000e-12'
+ mcl1f_cf_w_0_170_s_0_450 = '-6.15625e-14*ic_cap*ic_cap+-3.37500e-14*ic_cap+7.78000e-12'
+ mcl1f_cf_w_0_170_s_0_540 = '-7.68750e-14*ic_cap*ic_cap+-4.25000e-14*ic_cap+9.40000e-12'
+ mcl1f_cf_w_0_170_s_0_720 = '-1.03125e-13*ic_cap*ic_cap+-6.25000e-14*ic_cap+1.20000e-11'
+ mcl1f_cf_w_0_170_s_1_080 = '-1.50000e-13*ic_cap*ic_cap+-7.50000e-14*ic_cap+1.66000e-11'
+ mcl1f_cf_w_0_170_s_1_980 = '-1.96875e-13*ic_cap*ic_cap+-1.12500e-13*ic_cap+2.36000e-11'
+ mcl1f_cf_w_0_170_s_4_500 = '-2.03125e-13*ic_cap*ic_cap+-1.37500e-13*ic_cap+3.09000e-11'
+ mcl1f_cf_w_1_360_s_0_180 = '-1.06250e-14*ic_cap*ic_cap+-5.00000e-15*ic_cap+3.26000e-12'
+ mcl1f_cf_w_1_360_s_0_225 = '-1.87500e-14*ic_cap*ic_cap+-1.00000e-14*ic_cap+4.04000e-12'
+ mcl1f_cf_w_1_360_s_0_270 = '-2.75000e-14*ic_cap*ic_cap+-1.50000e-14*ic_cap+4.82000e-12'
+ mcl1f_cf_w_1_360_s_0_360 = '-4.43750e-14*ic_cap*ic_cap+-2.50000e-14*ic_cap+6.35000e-12'
+ mcl1f_cf_w_1_360_s_0_450 = '-6.03125e-14*ic_cap*ic_cap+-3.37500e-14*ic_cap+7.83000e-12'
+ mcl1f_cf_w_1_360_s_0_540 = '-7.53125e-14*ic_cap*ic_cap+-4.12500e-14*ic_cap+9.25000e-12'
+ mcl1f_cf_w_1_360_s_0_720 = '-1.00000e-13*ic_cap*ic_cap+-5.00000e-14*ic_cap+1.19000e-11'
+ mcl1f_cf_w_1_360_s_1_080 = '-1.46875e-13*ic_cap*ic_cap+-8.75000e-14*ic_cap+1.67000e-11'
+ mcl1f_cf_w_1_360_s_1_980 = '-1.96875e-13*ic_cap*ic_cap+-1.12500e-13*ic_cap+2.53000e-11'
+ mcl1f_cf_w_1_360_s_4_500 = '-2.03125e-13*ic_cap*ic_cap+-1.37500e-13*ic_cap+3.57000e-11'
+ mcl1p1_ca_w_0_170_s_0_180 = '-1.65000e-06*ic_cap*ic_cap+-8.00000e-07*ic_cap+9.41000e-05'
+ mcl1p1_ca_w_0_170_s_0_225 = '-1.65000e-06*ic_cap*ic_cap+-8.00000e-07*ic_cap+9.41000e-05'
+ mcl1p1_ca_w_0_170_s_0_270 = '-1.65000e-06*ic_cap*ic_cap+-8.00000e-07*ic_cap+9.41000e-05'
+ mcl1p1_ca_w_0_170_s_0_360 = '-1.65000e-06*ic_cap*ic_cap+-8.00000e-07*ic_cap+9.41000e-05'
+ mcl1p1_ca_w_0_170_s_0_450 = '-1.65000e-06*ic_cap*ic_cap+-8.00000e-07*ic_cap+9.41000e-05'
+ mcl1p1_ca_w_0_170_s_0_540 = '-1.65000e-06*ic_cap*ic_cap+-8.00000e-07*ic_cap+9.41000e-05'
+ mcl1p1_ca_w_0_170_s_0_720 = '-1.65000e-06*ic_cap*ic_cap+-8.00000e-07*ic_cap+9.41000e-05'
+ mcl1p1_ca_w_0_170_s_1_080 = '-1.65000e-06*ic_cap*ic_cap+-8.00000e-07*ic_cap+9.41000e-05'
+ mcl1p1_ca_w_0_170_s_1_980 = '-1.65000e-06*ic_cap*ic_cap+-8.00000e-07*ic_cap+9.41000e-05'
+ mcl1p1_ca_w_0_170_s_4_500 = '-1.65000e-06*ic_cap*ic_cap+-8.00000e-07*ic_cap+9.41000e-05'
+ mcl1p1_ca_w_1_360_s_0_180 = '-1.65000e-06*ic_cap*ic_cap+-8.00000e-07*ic_cap+9.41000e-05'
+ mcl1p1_ca_w_1_360_s_0_225 = '-1.65000e-06*ic_cap*ic_cap+-8.00000e-07*ic_cap+9.41000e-05'
+ mcl1p1_ca_w_1_360_s_0_270 = '-1.65000e-06*ic_cap*ic_cap+-8.00000e-07*ic_cap+9.41000e-05'
+ mcl1p1_ca_w_1_360_s_0_360 = '-1.65000e-06*ic_cap*ic_cap+-8.00000e-07*ic_cap+9.41000e-05'
+ mcl1p1_ca_w_1_360_s_0_450 = '-1.65000e-06*ic_cap*ic_cap+-8.00000e-07*ic_cap+9.41000e-05'
+ mcl1p1_ca_w_1_360_s_0_540 = '-1.65000e-06*ic_cap*ic_cap+-8.00000e-07*ic_cap+9.41000e-05'
+ mcl1p1_ca_w_1_360_s_0_720 = '-1.65000e-06*ic_cap*ic_cap+-8.00000e-07*ic_cap+9.41000e-05'
+ mcl1p1_ca_w_1_360_s_1_080 = '-1.65000e-06*ic_cap*ic_cap+-8.00000e-07*ic_cap+9.41000e-05'
+ mcl1p1_ca_w_1_360_s_1_980 = '-1.65000e-06*ic_cap*ic_cap+-8.00000e-07*ic_cap+9.41000e-05'
+ mcl1p1_ca_w_1_360_s_4_500 = '-1.65000e-06*ic_cap*ic_cap+-8.00000e-07*ic_cap+9.41000e-05'
+ mcl1p1_cc_w_0_170_s_0_180 = '-6.81250e-13*ic_cap*ic_cap+-4.50000e-13*ic_cap+7.32000e-11'
+ mcl1p1_cc_w_0_170_s_0_225 = '-4.65625e-13*ic_cap*ic_cap+-3.37500e-13*ic_cap+6.12000e-11'
+ mcl1p1_cc_w_0_170_s_0_270 = '-3.25000e-13*ic_cap*ic_cap+-2.50000e-13*ic_cap+5.32000e-11'
+ mcl1p1_cc_w_0_170_s_0_360 = '-1.75000e-13*ic_cap*ic_cap+-1.50000e-13*ic_cap+4.16000e-11'
+ mcl1p1_cc_w_0_170_s_0_450 = '-8.12500e-14*ic_cap*ic_cap+-1.00000e-13*ic_cap+3.45000e-11'
+ mcl1p1_cc_w_0_170_s_0_540 = '-2.81250e-14*ic_cap*ic_cap+-6.25000e-14*ic_cap+2.86000e-11'
+ mcl1p1_cc_w_0_170_s_0_720 = '3.12500e-14*ic_cap*ic_cap+-2.50000e-14*ic_cap+2.11000e-11'
+ mcl1p1_cc_w_0_170_s_1_080 = '6.87500e-14*ic_cap*ic_cap+2.50000e-14*ic_cap+1.28000e-11'
+ mcl1p1_cc_w_0_170_s_1_980 = '5.62500e-14*ic_cap*ic_cap+2.50000e-14*ic_cap+5.43000e-12'
+ mcl1p1_cc_w_0_170_s_4_500 = '1.90625e-14*ic_cap*ic_cap+1.12500e-14*ic_cap+1.35000e-12'
+ mcl1p1_cc_w_1_360_s_0_180 = '-6.03125e-13*ic_cap*ic_cap+-3.87500e-13*ic_cap+9.13000e-11'
+ mcl1p1_cc_w_1_360_s_0_225 = '-3.87500e-13*ic_cap*ic_cap+-2.75000e-13*ic_cap+7.85000e-11'
+ mcl1p1_cc_w_1_360_s_0_270 = '-2.62500e-13*ic_cap*ic_cap+-2.00000e-13*ic_cap+6.93000e-11'
+ mcl1p1_cc_w_1_360_s_0_360 = '-1.21875e-13*ic_cap*ic_cap+-1.12500e-13*ic_cap+5.66000e-11'
+ mcl1p1_cc_w_1_360_s_0_450 = '-4.06250e-14*ic_cap*ic_cap+-6.25000e-14*ic_cap+4.82000e-11'
+ mcl1p1_cc_w_1_360_s_0_540 = '9.37500e-15*ic_cap*ic_cap+-3.75000e-14*ic_cap+4.19000e-11'
+ mcl1p1_cc_w_1_360_s_0_720 = '5.93750e-14*ic_cap*ic_cap+1.25000e-14*ic_cap+3.32000e-11'
+ mcl1p1_cc_w_1_360_s_1_080 = '9.06250e-14*ic_cap*ic_cap+3.75000e-14*ic_cap+2.31000e-11'
+ mcl1p1_cc_w_1_360_s_1_980 = '8.12500e-14*ic_cap*ic_cap+5.00000e-14*ic_cap+1.19000e-11'
+ mcl1p1_cc_w_1_360_s_4_500 = '3.59375e-14*ic_cap*ic_cap+1.87500e-14*ic_cap+3.90000e-12'
+ mcl1p1_cf_w_0_170_s_0_180 = '-8.25000e-14*ic_cap*ic_cap+-3.75000e-14*ic_cap+8.06000e-12'
+ mcl1p1_cf_w_0_170_s_0_225 = '-1.12812e-13*ic_cap*ic_cap+-5.37500e-14*ic_cap+9.91000e-12'
+ mcl1p1_cf_w_0_170_s_0_270 = '-1.45000e-13*ic_cap*ic_cap+-6.75000e-14*ic_cap+1.17000e-11'
+ mcl1p1_cf_w_0_170_s_0_360 = '-1.90625e-13*ic_cap*ic_cap+-8.75000e-14*ic_cap+1.52000e-11'
+ mcl1p1_cf_w_0_170_s_0_450 = '-2.40625e-13*ic_cap*ic_cap+-1.12500e-13*ic_cap+1.80000e-11'
+ mcl1p1_cf_w_0_170_s_0_540 = '-2.87500e-13*ic_cap*ic_cap+-1.50000e-13*ic_cap+2.12000e-11'
+ mcl1p1_cf_w_0_170_s_0_720 = '-3.37500e-13*ic_cap*ic_cap+-1.75000e-13*ic_cap+2.58000e-11'
+ mcl1p1_cf_w_0_170_s_1_080 = '-3.90625e-13*ic_cap*ic_cap+-2.12500e-13*ic_cap+3.22000e-11'
+ mcl1p1_cf_w_0_170_s_1_980 = '-3.96875e-13*ic_cap*ic_cap+-2.37500e-13*ic_cap+3.89000e-11'
+ mcl1p1_cf_w_0_170_s_4_500 = '-3.62500e-13*ic_cap*ic_cap+-2.25000e-13*ic_cap+4.29000e-11'
+ mcl1p1_cf_w_1_360_s_0_180 = '-8.37500e-14*ic_cap*ic_cap+-3.75000e-14*ic_cap+8.11000e-12'
+ mcl1p1_cf_w_1_360_s_0_225 = '-1.14688e-13*ic_cap*ic_cap+-5.37500e-14*ic_cap+9.97000e-12'
+ mcl1p1_cf_w_1_360_s_0_270 = '-1.46563e-13*ic_cap*ic_cap+-6.87500e-14*ic_cap+1.18000e-11'
+ mcl1p1_cf_w_1_360_s_0_360 = '-1.93750e-13*ic_cap*ic_cap+-1.00000e-13*ic_cap+1.51000e-11'
+ mcl1p1_cf_w_1_360_s_0_450 = '-2.40625e-13*ic_cap*ic_cap+-1.12500e-13*ic_cap+1.82000e-11'
+ mcl1p1_cf_w_1_360_s_0_540 = '-2.84375e-13*ic_cap*ic_cap+-1.37500e-13*ic_cap+2.11000e-11'
+ mcl1p1_cf_w_1_360_s_0_720 = '-3.37500e-13*ic_cap*ic_cap+-1.75000e-13*ic_cap+2.59000e-11'
+ mcl1p1_cf_w_1_360_s_1_080 = '-3.96875e-13*ic_cap*ic_cap+-2.12500e-13*ic_cap+3.31000e-11'
+ mcl1p1_cf_w_1_360_s_1_980 = '-4.21875e-13*ic_cap*ic_cap+-2.37500e-13*ic_cap+4.28000e-11'
+ mcl1p1_cf_w_1_360_s_4_500 = '-3.87500e-13*ic_cap*ic_cap+-2.25000e-13*ic_cap+5.06000e-11'
+ mcl1p1f_ca_w_0_150_s_0_210 = '-3.03125e-06*ic_cap*ic_cap+-1.62500e-06*ic_cap+2.00000e-04'
+ mcl1p1f_ca_w_0_150_s_0_263 = '-3.03125e-06*ic_cap*ic_cap+-1.62500e-06*ic_cap+2.00000e-04'
+ mcl1p1f_ca_w_0_150_s_0_315 = '-3.03125e-06*ic_cap*ic_cap+-1.62500e-06*ic_cap+2.00000e-04'
+ mcl1p1f_ca_w_0_150_s_0_420 = '-3.03125e-06*ic_cap*ic_cap+-1.62500e-06*ic_cap+2.00000e-04'
+ mcl1p1f_ca_w_0_150_s_0_525 = '-3.03125e-06*ic_cap*ic_cap+-1.62500e-06*ic_cap+2.00000e-04'
+ mcl1p1f_ca_w_0_150_s_0_630 = '-3.03125e-06*ic_cap*ic_cap+-1.62500e-06*ic_cap+2.00000e-04'
+ mcl1p1f_ca_w_0_150_s_0_840 = '-3.03125e-06*ic_cap*ic_cap+-1.62500e-06*ic_cap+2.00000e-04'
+ mcl1p1f_ca_w_0_150_s_1_260 = '-3.03125e-06*ic_cap*ic_cap+-1.62500e-06*ic_cap+2.00000e-04'
+ mcl1p1f_ca_w_0_150_s_2_310 = '-3.03125e-06*ic_cap*ic_cap+-1.62500e-06*ic_cap+2.00000e-04'
+ mcl1p1f_ca_w_0_150_s_5_250 = '-3.03125e-06*ic_cap*ic_cap+-1.62500e-06*ic_cap+2.00000e-04'
+ mcl1p1f_ca_w_1_200_s_0_210 = '-3.03125e-06*ic_cap*ic_cap+-1.62500e-06*ic_cap+2.00000e-04'
+ mcl1p1f_ca_w_1_200_s_0_263 = '-3.03125e-06*ic_cap*ic_cap+-1.62500e-06*ic_cap+2.00000e-04'
+ mcl1p1f_ca_w_1_200_s_0_315 = '-3.03125e-06*ic_cap*ic_cap+-1.62500e-06*ic_cap+2.00000e-04'
+ mcl1p1f_ca_w_1_200_s_0_420 = '-3.03125e-06*ic_cap*ic_cap+-1.62500e-06*ic_cap+2.00000e-04'
+ mcl1p1f_ca_w_1_200_s_0_525 = '-3.03125e-06*ic_cap*ic_cap+-1.62500e-06*ic_cap+2.00000e-04'
+ mcl1p1f_ca_w_1_200_s_0_630 = '-3.03125e-06*ic_cap*ic_cap+-1.62500e-06*ic_cap+2.00000e-04'
+ mcl1p1f_ca_w_1_200_s_0_840 = '-3.03125e-06*ic_cap*ic_cap+-1.62500e-06*ic_cap+2.00000e-04'
+ mcl1p1f_ca_w_1_200_s_1_260 = '-3.03125e-06*ic_cap*ic_cap+-1.62500e-06*ic_cap+2.00000e-04'
+ mcl1p1f_ca_w_1_200_s_2_310 = '-3.03125e-06*ic_cap*ic_cap+-1.62500e-06*ic_cap+2.00000e-04'
+ mcl1p1f_ca_w_1_200_s_5_250 = '-3.03125e-06*ic_cap*ic_cap+-1.62500e-06*ic_cap+2.00000e-04'
+ mcl1p1f_cc_w_0_150_s_0_210 = '-3.93750e-13*ic_cap*ic_cap+-2.25000e-13*ic_cap+6.42000e-11'
+ mcl1p1f_cc_w_0_150_s_0_263 = '-1.78125e-13*ic_cap*ic_cap+-1.12500e-13*ic_cap+4.90000e-11'
+ mcl1p1f_cc_w_0_150_s_0_315 = '-6.87500e-14*ic_cap*ic_cap+-5.00000e-14*ic_cap+3.87000e-11'
+ mcl1p1f_cc_w_0_150_s_0_420 = '5.31250e-14*ic_cap*ic_cap+1.25000e-14*ic_cap+2.56000e-11'
+ mcl1p1f_cc_w_0_150_s_0_525 = '1.03125e-13*ic_cap*ic_cap+3.75000e-14*ic_cap+1.74000e-11'
+ mcl1p1f_cc_w_0_150_s_0_630 = '1.15625e-13*ic_cap*ic_cap+6.25000e-14*ic_cap+1.21000e-11'
+ mcl1p1f_cc_w_0_150_s_0_840 = '1.12500e-13*ic_cap*ic_cap+6.75000e-14*ic_cap+5.89000e-12'
+ mcl1p1f_cc_w_0_150_s_1_260 = '5.65625e-14*ic_cap*ic_cap+4.12500e-14*ic_cap+1.52000e-12'
+ mcl1p1f_cc_w_0_150_s_2_310 = '4.84375e-15*ic_cap*ic_cap+1.87500e-15*ic_cap+1.10000e-13'
+ mcl1p1f_cc_w_0_150_s_5_250 = '-3.12500e-16*ic_cap*ic_cap+4.03897e-28*ic_cap+5.00000e-15'
+ mcl1p1f_cc_w_1_200_s_0_210 = '-2.93750e-13*ic_cap*ic_cap+-1.50000e-13*ic_cap+6.64000e-11'
+ mcl1p1f_cc_w_1_200_s_0_263 = '-1.00000e-13*ic_cap*ic_cap+-7.50000e-14*ic_cap+5.07000e-11'
+ mcl1p1f_cc_w_1_200_s_0_315 = '6.25000e-15*ic_cap*ic_cap+-2.50000e-14*ic_cap+4.02000e-11'
+ mcl1p1f_cc_w_1_200_s_0_420 = '1.06250e-13*ic_cap*ic_cap+5.00000e-14*ic_cap+2.66000e-11'
+ mcl1p1f_cc_w_1_200_s_0_525 = '1.50000e-13*ic_cap*ic_cap+1.00000e-13*ic_cap+1.81000e-11'
+ mcl1p1f_cc_w_1_200_s_0_630 = '1.56250e-13*ic_cap*ic_cap+7.50000e-14*ic_cap+1.26000e-11'
+ mcl1p1f_cc_w_1_200_s_0_840 = '1.37500e-13*ic_cap*ic_cap+8.75000e-14*ic_cap+6.20000e-12'
+ mcl1p1f_cc_w_1_200_s_1_260 = '6.87500e-14*ic_cap*ic_cap+5.00000e-14*ic_cap+1.60000e-12'
+ mcl1p1f_cc_w_1_200_s_2_310 = '3.12500e-15*ic_cap*ic_cap+-3.15544e-30*ic_cap+1.50000e-13'
+ mcl1p1f_cf_w_0_150_s_0_210 = '-2.06250e-13*ic_cap*ic_cap+-1.00000e-13*ic_cap+1.91000e-11'
+ mcl1p1f_cf_w_0_150_s_0_263 = '-2.62500e-13*ic_cap*ic_cap+-1.25000e-13*ic_cap+2.32000e-11'
+ mcl1p1f_cf_w_0_150_s_0_315 = '-3.03125e-13*ic_cap*ic_cap+-1.62500e-13*ic_cap+2.68000e-11'
+ mcl1p1f_cf_w_0_150_s_0_420 = '-3.81250e-13*ic_cap*ic_cap+-2.00000e-13*ic_cap+3.33000e-11'
+ mcl1p1f_cf_w_0_150_s_0_525 = '-4.34375e-13*ic_cap*ic_cap+-2.37500e-13*ic_cap+3.84000e-11'
+ mcl1p1f_cf_w_0_150_s_0_630 = '-4.62500e-13*ic_cap*ic_cap+-2.50000e-13*ic_cap+4.23000e-11'
+ mcl1p1f_cf_w_0_150_s_0_840 = '-4.68750e-13*ic_cap*ic_cap+-2.75000e-13*ic_cap+4.74000e-11'
+ mcl1p1f_cf_w_0_150_s_1_260 = '-4.25000e-13*ic_cap*ic_cap+-2.50000e-13*ic_cap+5.15000e-11'
+ mcl1p1f_cf_w_0_150_s_2_310 = '-3.84375e-13*ic_cap*ic_cap+-2.12500e-13*ic_cap+5.29000e-11'
+ mcl1p1f_cf_w_0_150_s_5_250 = '-3.75000e-13*ic_cap*ic_cap+-2.00000e-13*ic_cap+5.30000e-11'
+ mcl1p1f_cf_w_1_200_s_0_210 = '-2.00000e-13*ic_cap*ic_cap+-1.00000e-13*ic_cap+1.90000e-11'
+ mcl1p1f_cf_w_1_200_s_0_263 = '-2.56250e-13*ic_cap*ic_cap+-1.25000e-13*ic_cap+2.31000e-11'
+ mcl1p1f_cf_w_1_200_s_0_315 = '-3.09375e-13*ic_cap*ic_cap+-1.62500e-13*ic_cap+2.69000e-11'
+ mcl1p1f_cf_w_1_200_s_0_420 = '-3.81250e-13*ic_cap*ic_cap+-2.00000e-13*ic_cap+3.34000e-11'
+ mcl1p1f_cf_w_1_200_s_0_525 = '-4.25000e-13*ic_cap*ic_cap+-2.25000e-13*ic_cap+3.86000e-11'
+ mcl1p1f_cf_w_1_200_s_0_630 = '-4.46875e-13*ic_cap*ic_cap+-2.37500e-13*ic_cap+4.26000e-11'
+ mcl1p1f_cf_w_1_200_s_0_840 = '-4.56250e-13*ic_cap*ic_cap+-2.50000e-13*ic_cap+4.80000e-11'
+ mcl1p1f_cf_w_1_200_s_1_260 = '-4.06250e-13*ic_cap*ic_cap+-2.25000e-13*ic_cap+5.23000e-11'
+ mcl1p1f_cf_w_1_200_s_2_310 = '-3.46875e-13*ic_cap*ic_cap+-1.87500e-13*ic_cap+5.37000e-11'
+ mcl1p1f_cf_w_1_200_s_5_250 = '-3.40625e-13*ic_cap*ic_cap+-1.87500e-13*ic_cap+5.38000e-11'
+ mcm1d_ca_w_0_140_s_0_140 = '-3.71875e-07*ic_cap*ic_cap+-2.37500e-07*ic_cap+3.36000e-05'
+ mcm1d_ca_w_0_140_s_0_175 = '-3.71875e-07*ic_cap*ic_cap+-2.37500e-07*ic_cap+3.36000e-05'
+ mcm1d_ca_w_0_140_s_0_210 = '-3.71875e-07*ic_cap*ic_cap+-2.37500e-07*ic_cap+3.36000e-05'
+ mcm1d_ca_w_0_140_s_0_280 = '-3.71875e-07*ic_cap*ic_cap+-2.37500e-07*ic_cap+3.36000e-05'
+ mcm1d_ca_w_0_140_s_0_350 = '-3.71875e-07*ic_cap*ic_cap+-2.37500e-07*ic_cap+3.36000e-05'
+ mcm1d_ca_w_0_140_s_0_420 = '-3.71875e-07*ic_cap*ic_cap+-2.37500e-07*ic_cap+3.36000e-05'
+ mcm1d_ca_w_0_140_s_0_560 = '-3.71875e-07*ic_cap*ic_cap+-2.37500e-07*ic_cap+3.36000e-05'
+ mcm1d_ca_w_0_140_s_0_840 = '-3.71875e-07*ic_cap*ic_cap+-2.37500e-07*ic_cap+3.36000e-05'
+ mcm1d_ca_w_0_140_s_1_540 = '-3.71875e-07*ic_cap*ic_cap+-2.37500e-07*ic_cap+3.36000e-05'
+ mcm1d_ca_w_0_140_s_3_500 = '-3.71875e-07*ic_cap*ic_cap+-2.37500e-07*ic_cap+3.36000e-05'
+ mcm1d_ca_w_1_120_s_0_140 = '-3.71875e-07*ic_cap*ic_cap+-2.37500e-07*ic_cap+3.36000e-05'
+ mcm1d_ca_w_1_120_s_0_175 = '-3.71875e-07*ic_cap*ic_cap+-2.37500e-07*ic_cap+3.36000e-05'
+ mcm1d_ca_w_1_120_s_0_210 = '-3.71875e-07*ic_cap*ic_cap+-2.37500e-07*ic_cap+3.36000e-05'
+ mcm1d_ca_w_1_120_s_0_280 = '-3.71875e-07*ic_cap*ic_cap+-2.37500e-07*ic_cap+3.36000e-05'
+ mcm1d_ca_w_1_120_s_0_350 = '-3.71875e-07*ic_cap*ic_cap+-2.37500e-07*ic_cap+3.36000e-05'
+ mcm1d_ca_w_1_120_s_0_420 = '-3.71875e-07*ic_cap*ic_cap+-2.37500e-07*ic_cap+3.36000e-05'
+ mcm1d_ca_w_1_120_s_0_560 = '-3.71875e-07*ic_cap*ic_cap+-2.37500e-07*ic_cap+3.36000e-05'
+ mcm1d_ca_w_1_120_s_0_840 = '-3.71875e-07*ic_cap*ic_cap+-2.37500e-07*ic_cap+3.36000e-05'
+ mcm1d_ca_w_1_120_s_1_540 = '-3.71875e-07*ic_cap*ic_cap+-2.37500e-07*ic_cap+3.36000e-05'
+ mcm1d_ca_w_1_120_s_3_500 = '-3.71875e-07*ic_cap*ic_cap+-2.37500e-07*ic_cap+3.36000e-05'
+ mcm1d_cc_w_0_140_s_0_140 = '-9.21875e-13*ic_cap*ic_cap+-4.62500e-13*ic_cap+1.04000e-10'
+ mcm1d_cc_w_0_140_s_0_175 = '-8.53125e-13*ic_cap*ic_cap+-5.87500e-13*ic_cap+1.02000e-10'
+ mcm1d_cc_w_0_140_s_0_210 = '-7.34375e-13*ic_cap*ic_cap+-4.62500e-13*ic_cap+9.66000e-11'
+ mcm1d_cc_w_0_140_s_0_280 = '-5.93750e-13*ic_cap*ic_cap+-3.75000e-13*ic_cap+8.60000e-11'
+ mcm1d_cc_w_0_140_s_0_350 = '-4.40625e-13*ic_cap*ic_cap+-3.12500e-13*ic_cap+7.46000e-11'
+ mcm1d_cc_w_0_140_s_0_420 = '-3.43750e-13*ic_cap*ic_cap+-2.75000e-13*ic_cap+6.53000e-11'
+ mcm1d_cc_w_0_140_s_0_560 = '-2.06250e-13*ic_cap*ic_cap+-1.25000e-13*ic_cap+5.27000e-11'
+ mcm1d_cc_w_0_140_s_0_840 = '-8.43750e-14*ic_cap*ic_cap+-6.25000e-14*ic_cap+3.84000e-11'
+ mcm1d_cc_w_0_140_s_1_540 = '9.37500e-15*ic_cap*ic_cap+1.25000e-14*ic_cap+2.23000e-11'
+ mcm1d_cc_w_0_140_s_3_500 = '3.93750e-14*ic_cap*ic_cap+2.75000e-14*ic_cap+8.26000e-12'
+ mcm1d_cc_w_1_120_s_0_140 = '-8.43750e-13*ic_cap*ic_cap+-3.75000e-13*ic_cap+1.28000e-10'
+ mcm1d_cc_w_1_120_s_0_175 = '-7.50000e-13*ic_cap*ic_cap+-2.50000e-13*ic_cap+1.24000e-10'
+ mcm1d_cc_w_1_120_s_0_210 = '-6.56250e-13*ic_cap*ic_cap+-3.75000e-13*ic_cap+1.18000e-10'
+ mcm1d_cc_w_1_120_s_0_280 = '-4.84375e-13*ic_cap*ic_cap+-2.87500e-13*ic_cap+1.04000e-10'
+ mcm1d_cc_w_1_120_s_0_350 = '-3.84375e-13*ic_cap*ic_cap+-2.62500e-13*ic_cap+9.17000e-11'
+ mcm1d_cc_w_1_120_s_0_420 = '-2.84375e-13*ic_cap*ic_cap+-2.12500e-13*ic_cap+8.11000e-11'
+ mcm1d_cc_w_1_120_s_0_560 = '-1.37500e-13*ic_cap*ic_cap+-1.00000e-13*ic_cap+6.60000e-11'
+ mcm1d_cc_w_1_120_s_0_840 = '-4.37500e-14*ic_cap*ic_cap+-2.50000e-14*ic_cap+4.91000e-11'
+ mcm1d_cc_w_1_120_s_1_540 = '3.75000e-14*ic_cap*ic_cap+2.50000e-14*ic_cap+3.01000e-11'
+ mcm1d_cc_w_1_120_s_3_500 = '5.93750e-14*ic_cap*ic_cap+3.75000e-14*ic_cap+1.26000e-11'
+ mcm1d_cf_w_0_140_s_0_140 = '-4.06250e-15*ic_cap*ic_cap+-3.75000e-15*ic_cap+2.32000e-12'
+ mcm1d_cf_w_0_140_s_0_175 = '-1.00000e-14*ic_cap*ic_cap+-7.50000e-15*ic_cap+2.90000e-12'
+ mcm1d_cf_w_0_140_s_0_210 = '-1.68750e-14*ic_cap*ic_cap+-1.25000e-14*ic_cap+3.49000e-12'
+ mcm1d_cf_w_0_140_s_0_280 = '-2.90625e-14*ic_cap*ic_cap+-2.12500e-14*ic_cap+4.62000e-12'
+ mcm1d_cf_w_0_140_s_0_350 = '-4.21875e-14*ic_cap*ic_cap+-2.87500e-14*ic_cap+5.73000e-12'
+ mcm1d_cf_w_0_140_s_0_420 = '-5.34375e-14*ic_cap*ic_cap+-3.62500e-14*ic_cap+6.87000e-12'
+ mcm1d_cf_w_0_140_s_0_560 = '-7.50000e-14*ic_cap*ic_cap+-4.75000e-14*ic_cap+8.91000e-12'
+ mcm1d_cf_w_0_140_s_0_840 = '-1.18750e-13*ic_cap*ic_cap+-7.50000e-14*ic_cap+1.28000e-11'
+ mcm1d_cf_w_0_140_s_1_540 = '-1.81250e-13*ic_cap*ic_cap+-1.25000e-13*ic_cap+2.05000e-11'
+ mcm1d_cf_w_0_140_s_3_500 = '-2.31250e-13*ic_cap*ic_cap+-1.50000e-13*ic_cap+3.15000e-11'
+ mcm1d_cf_w_1_120_s_0_140 = '-5.62500e-15*ic_cap*ic_cap+-5.00000e-15*ic_cap+2.39000e-12'
+ mcm1d_cf_w_1_120_s_0_175 = '-1.09375e-14*ic_cap*ic_cap+-8.75000e-15*ic_cap+2.96000e-12'
+ mcm1d_cf_w_1_120_s_0_210 = '-1.75000e-14*ic_cap*ic_cap+-1.25000e-14*ic_cap+3.54000e-12'
+ mcm1d_cf_w_1_120_s_0_280 = '-3.00000e-14*ic_cap*ic_cap+-2.25000e-14*ic_cap+4.68000e-12'
+ mcm1d_cf_w_1_120_s_0_350 = '-4.18750e-14*ic_cap*ic_cap+-3.00000e-14*ic_cap+5.80000e-12'
+ mcm1d_cf_w_1_120_s_0_420 = '-5.37500e-14*ic_cap*ic_cap+-3.75000e-14*ic_cap+6.89000e-12'
+ mcm1d_cf_w_1_120_s_0_560 = '-7.59375e-14*ic_cap*ic_cap+-5.12500e-14*ic_cap+8.99000e-12'
+ mcm1d_cf_w_1_120_s_0_840 = '-1.12500e-13*ic_cap*ic_cap+-7.50000e-14*ic_cap+1.29000e-11'
+ mcm1d_cf_w_1_120_s_1_540 = '-1.81250e-13*ic_cap*ic_cap+-1.25000e-13*ic_cap+2.09000e-11'
+ mcm1d_cf_w_1_120_s_3_500 = '-2.28125e-13*ic_cap*ic_cap+-1.62500e-13*ic_cap+3.36000e-11'
+ mcm1f_ca_w_0_140_s_0_140 = '-3.03125e-07*ic_cap*ic_cap+-1.87500e-07*ic_cap+2.58000e-05'
+ mcm1f_ca_w_0_140_s_0_175 = '-3.03125e-07*ic_cap*ic_cap+-1.87500e-07*ic_cap+2.58000e-05'
+ mcm1f_ca_w_0_140_s_0_210 = '-3.03125e-07*ic_cap*ic_cap+-1.87500e-07*ic_cap+2.58000e-05'
+ mcm1f_ca_w_0_140_s_0_280 = '-3.03125e-07*ic_cap*ic_cap+-1.87500e-07*ic_cap+2.58000e-05'
+ mcm1f_ca_w_0_140_s_0_350 = '-3.03125e-07*ic_cap*ic_cap+-1.87500e-07*ic_cap+2.58000e-05'
+ mcm1f_ca_w_0_140_s_0_420 = '-3.03125e-07*ic_cap*ic_cap+-1.87500e-07*ic_cap+2.58000e-05'
+ mcm1f_ca_w_0_140_s_0_560 = '-3.03125e-07*ic_cap*ic_cap+-1.87500e-07*ic_cap+2.58000e-05'
+ mcm1f_ca_w_0_140_s_0_840 = '-3.03125e-07*ic_cap*ic_cap+-1.87500e-07*ic_cap+2.58000e-05'
+ mcm1f_ca_w_0_140_s_1_540 = '-3.03125e-07*ic_cap*ic_cap+-1.87500e-07*ic_cap+2.58000e-05'
+ mcm1f_ca_w_0_140_s_3_500 = '-3.03125e-07*ic_cap*ic_cap+-1.87500e-07*ic_cap+2.58000e-05'
+ mcm1f_ca_w_1_120_s_0_140 = '-3.03125e-07*ic_cap*ic_cap+-1.87500e-07*ic_cap+2.58000e-05'
+ mcm1f_ca_w_1_120_s_0_175 = '-3.03125e-07*ic_cap*ic_cap+-1.87500e-07*ic_cap+2.58000e-05'
+ mcm1f_ca_w_1_120_s_0_210 = '-3.03125e-07*ic_cap*ic_cap+-1.87500e-07*ic_cap+2.58000e-05'
+ mcm1f_ca_w_1_120_s_0_280 = '-3.03125e-07*ic_cap*ic_cap+-1.87500e-07*ic_cap+2.58000e-05'
+ mcm1f_ca_w_1_120_s_0_350 = '-3.03125e-07*ic_cap*ic_cap+-1.87500e-07*ic_cap+2.58000e-05'
+ mcm1f_ca_w_1_120_s_0_420 = '-3.03125e-07*ic_cap*ic_cap+-1.87500e-07*ic_cap+2.58000e-05'
+ mcm1f_ca_w_1_120_s_0_560 = '-3.03125e-07*ic_cap*ic_cap+-1.87500e-07*ic_cap+2.58000e-05'
+ mcm1f_ca_w_1_120_s_0_840 = '-3.03125e-07*ic_cap*ic_cap+-1.87500e-07*ic_cap+2.58000e-05'
+ mcm1f_ca_w_1_120_s_1_540 = '-3.03125e-07*ic_cap*ic_cap+-1.87500e-07*ic_cap+2.58000e-05'
+ mcm1f_ca_w_1_120_s_3_500 = '-3.03125e-07*ic_cap*ic_cap+-1.87500e-07*ic_cap+2.58000e-05'
+ mcm1f_cc_w_0_140_s_0_140 = '-9.40625e-13*ic_cap*ic_cap+-4.87500e-13*ic_cap+1.05000e-10'
+ mcm1f_cc_w_0_140_s_0_175 = '-8.62500e-13*ic_cap*ic_cap+-5.75000e-13*ic_cap+1.03000e-10'
+ mcm1f_cc_w_0_140_s_0_210 = '-7.65625e-13*ic_cap*ic_cap+-4.37500e-13*ic_cap+9.77000e-11'
+ mcm1f_cc_w_0_140_s_0_280 = '-6.18750e-13*ic_cap*ic_cap+-4.25000e-13*ic_cap+8.76000e-11'
+ mcm1f_cc_w_0_140_s_0_350 = '-4.68750e-13*ic_cap*ic_cap+-3.00000e-13*ic_cap+7.63000e-11'
+ mcm1f_cc_w_0_140_s_0_420 = '-3.71875e-13*ic_cap*ic_cap+-2.62500e-13*ic_cap+6.70000e-11'
+ mcm1f_cc_w_0_140_s_0_560 = '-2.12500e-13*ic_cap*ic_cap+-1.50000e-13*ic_cap+5.45000e-11'
+ mcm1f_cc_w_0_140_s_0_840 = '-9.06250e-14*ic_cap*ic_cap+-6.25000e-14*ic_cap+4.05000e-11'
+ mcm1f_cc_w_0_140_s_1_540 = '6.25000e-15*ic_cap*ic_cap+2.47000e-11'
+ mcm1f_cc_w_0_140_s_3_500 = '5.00000e-14*ic_cap*ic_cap+2.50000e-14*ic_cap+1.00000e-11'
+ mcm1f_cc_w_1_120_s_0_140 = '-8.75000e-13*ic_cap*ic_cap+-5.00000e-13*ic_cap+1.31000e-10'
+ mcm1f_cc_w_1_120_s_0_175 = '-7.81250e-13*ic_cap*ic_cap+-3.75000e-13*ic_cap+1.27000e-10'
+ mcm1f_cc_w_1_120_s_0_210 = '-7.18750e-13*ic_cap*ic_cap+-3.75000e-13*ic_cap+1.21000e-10'
+ mcm1f_cc_w_1_120_s_0_280 = '-5.09375e-13*ic_cap*ic_cap+-2.87500e-13*ic_cap+1.07000e-10'
+ mcm1f_cc_w_1_120_s_0_350 = '-3.90625e-13*ic_cap*ic_cap+-2.62500e-13*ic_cap+9.46000e-11'
+ mcm1f_cc_w_1_120_s_0_420 = '-2.81250e-13*ic_cap*ic_cap+-2.25000e-13*ic_cap+8.38000e-11'
+ mcm1f_cc_w_1_120_s_0_560 = '-1.43750e-13*ic_cap*ic_cap+-1.00000e-13*ic_cap+6.88000e-11'
+ mcm1f_cc_w_1_120_s_0_840 = '-4.06250e-14*ic_cap*ic_cap+-3.75000e-14*ic_cap+5.20000e-11'
+ mcm1f_cc_w_1_120_s_1_540 = '4.37500e-14*ic_cap*ic_cap+2.50000e-14*ic_cap+3.29000e-11'
+ mcm1f_cc_w_1_120_s_3_500 = '7.50000e-14*ic_cap*ic_cap+5.00000e-14*ic_cap+1.47000e-11'
+ mcm1f_cf_w_0_140_s_0_140 = '-4.68750e-15*ic_cap*ic_cap+-3.75000e-15*ic_cap+1.79000e-12'
+ mcm1f_cf_w_0_140_s_0_175 = '-9.06250e-15*ic_cap*ic_cap+-6.25000e-15*ic_cap+2.23000e-12'
+ mcm1f_cf_w_0_140_s_0_210 = '-1.43750e-14*ic_cap*ic_cap+-1.00000e-14*ic_cap+2.68000e-12'
+ mcm1f_cf_w_0_140_s_0_280 = '-2.46875e-14*ic_cap*ic_cap+-1.62500e-14*ic_cap+3.56000e-12'
+ mcm1f_cf_w_0_140_s_0_350 = '-3.50000e-14*ic_cap*ic_cap+-2.25000e-14*ic_cap+4.42000e-12'
+ mcm1f_cf_w_0_140_s_0_420 = '-4.40625e-14*ic_cap*ic_cap+-2.87500e-14*ic_cap+5.31000e-12'
+ mcm1f_cf_w_0_140_s_0_560 = '-6.37500e-14*ic_cap*ic_cap+-4.00000e-14*ic_cap+6.93000e-12'
+ mcm1f_cf_w_0_140_s_0_840 = '-9.65625e-14*ic_cap*ic_cap+-6.12500e-14*ic_cap+1.00000e-11'
+ mcm1f_cf_w_0_140_s_1_540 = '-1.56250e-13*ic_cap*ic_cap+-1.00000e-13*ic_cap+1.65000e-11'
+ mcm1f_cf_w_0_140_s_3_500 = '-2.18750e-13*ic_cap*ic_cap+-1.50000e-13*ic_cap+2.70000e-11'
+ mcm1f_cf_w_1_120_s_0_140 = '-4.68750e-15*ic_cap*ic_cap+-3.75000e-15*ic_cap+1.82000e-12'
+ mcm1f_cf_w_1_120_s_0_175 = '-1.06250e-14*ic_cap*ic_cap+-7.50000e-15*ic_cap+2.28000e-12'
+ mcm1f_cf_w_1_120_s_0_210 = '-1.56250e-14*ic_cap*ic_cap+-1.00000e-14*ic_cap+2.72000e-12'
+ mcm1f_cf_w_1_120_s_0_280 = '-2.62500e-14*ic_cap*ic_cap+-1.75000e-14*ic_cap+3.61000e-12'
+ mcm1f_cf_w_1_120_s_0_350 = '-3.53125e-14*ic_cap*ic_cap+-2.37500e-14*ic_cap+4.47000e-12'
+ mcm1f_cf_w_1_120_s_0_420 = '-4.56250e-14*ic_cap*ic_cap+-3.00000e-14*ic_cap+5.33000e-12'
+ mcm1f_cf_w_1_120_s_0_560 = '-6.40625e-14*ic_cap*ic_cap+-4.12500e-14*ic_cap+6.98000e-12'
+ mcm1f_cf_w_1_120_s_0_840 = '-9.75000e-14*ic_cap*ic_cap+-6.25000e-14*ic_cap+1.01000e-11'
+ mcm1f_cf_w_1_120_s_1_540 = '-1.62500e-13*ic_cap*ic_cap+-1.00000e-13*ic_cap+1.69000e-11'
+ mcm1f_cf_w_1_120_s_3_500 = '-2.31250e-13*ic_cap*ic_cap+-1.50000e-13*ic_cap+2.88000e-11'
+ mcm1l1_ca_w_0_140_s_0_140 = '-1.98438e-06*ic_cap*ic_cap+-1.26250e-06*ic_cap+1.14000e-04'
+ mcm1l1_ca_w_0_140_s_0_175 = '-1.98438e-06*ic_cap*ic_cap+-1.26250e-06*ic_cap+1.14000e-04'
+ mcm1l1_ca_w_0_140_s_0_210 = '-1.98438e-06*ic_cap*ic_cap+-1.26250e-06*ic_cap+1.14000e-04'
+ mcm1l1_ca_w_0_140_s_0_280 = '-1.98438e-06*ic_cap*ic_cap+-1.26250e-06*ic_cap+1.14000e-04'
+ mcm1l1_ca_w_0_140_s_0_350 = '-1.98438e-06*ic_cap*ic_cap+-1.26250e-06*ic_cap+1.14000e-04'
+ mcm1l1_ca_w_0_140_s_0_420 = '-1.98438e-06*ic_cap*ic_cap+-1.26250e-06*ic_cap+1.14000e-04'
+ mcm1l1_ca_w_0_140_s_0_560 = '-1.98438e-06*ic_cap*ic_cap+-1.26250e-06*ic_cap+1.14000e-04'
+ mcm1l1_ca_w_0_140_s_0_840 = '-1.98438e-06*ic_cap*ic_cap+-1.26250e-06*ic_cap+1.14000e-04'
+ mcm1l1_ca_w_0_140_s_1_540 = '-1.98438e-06*ic_cap*ic_cap+-1.26250e-06*ic_cap+1.14000e-04'
+ mcm1l1_ca_w_0_140_s_3_500 = '-1.98438e-06*ic_cap*ic_cap+-1.26250e-06*ic_cap+1.14000e-04'
+ mcm1l1_ca_w_1_120_s_0_140 = '-1.98438e-06*ic_cap*ic_cap+-1.26250e-06*ic_cap+1.14000e-04'
+ mcm1l1_ca_w_1_120_s_0_175 = '-1.98438e-06*ic_cap*ic_cap+-1.26250e-06*ic_cap+1.14000e-04'
+ mcm1l1_ca_w_1_120_s_0_210 = '-1.98438e-06*ic_cap*ic_cap+-1.26250e-06*ic_cap+1.14000e-04'
+ mcm1l1_ca_w_1_120_s_0_280 = '-1.98438e-06*ic_cap*ic_cap+-1.26250e-06*ic_cap+1.14000e-04'
+ mcm1l1_ca_w_1_120_s_0_350 = '-1.98438e-06*ic_cap*ic_cap+-1.26250e-06*ic_cap+1.14000e-04'
+ mcm1l1_ca_w_1_120_s_0_420 = '-1.98438e-06*ic_cap*ic_cap+-1.26250e-06*ic_cap+1.14000e-04'
+ mcm1l1_ca_w_1_120_s_0_560 = '-1.98438e-06*ic_cap*ic_cap+-1.26250e-06*ic_cap+1.14000e-04'
+ mcm1l1_ca_w_1_120_s_0_840 = '-1.98438e-06*ic_cap*ic_cap+-1.26250e-06*ic_cap+1.14000e-04'
+ mcm1l1_ca_w_1_120_s_1_540 = '-1.98438e-06*ic_cap*ic_cap+-1.26250e-06*ic_cap+1.14000e-04'
+ mcm1l1_ca_w_1_120_s_3_500 = '-1.98438e-06*ic_cap*ic_cap+-1.26250e-06*ic_cap+1.14000e-04'
+ mcm1l1_cc_w_0_140_s_0_140 = '-7.59375e-13*ic_cap*ic_cap+-4.37500e-13*ic_cap+9.58000e-11'
+ mcm1l1_cc_w_0_140_s_0_175 = '-7.21875e-13*ic_cap*ic_cap+-4.62500e-13*ic_cap+9.38000e-11'
+ mcm1l1_cc_w_0_140_s_0_210 = '-6.00000e-13*ic_cap*ic_cap+-3.25000e-13*ic_cap+8.80000e-11'
+ mcm1l1_cc_w_0_140_s_0_280 = '-4.28125e-13*ic_cap*ic_cap+-2.37500e-13*ic_cap+7.59000e-11'
+ mcm1l1_cc_w_0_140_s_0_350 = '-3.06250e-13*ic_cap*ic_cap+-2.25000e-13*ic_cap+6.44000e-11'
+ mcm1l1_cc_w_0_140_s_0_420 = '-1.96875e-13*ic_cap*ic_cap+-1.37500e-13*ic_cap+5.44000e-11'
+ mcm1l1_cc_w_0_140_s_0_560 = '-8.12500e-14*ic_cap*ic_cap+-2.50000e-14*ic_cap+4.13000e-11'
+ mcm1l1_cc_w_0_140_s_0_840 = '9.37500e-15*ic_cap*ic_cap+1.25000e-14*ic_cap+2.70000e-11'
+ mcm1l1_cc_w_0_140_s_1_540 = '4.68750e-14*ic_cap*ic_cap+6.25000e-14*ic_cap+1.25000e-11'
+ mcm1l1_cc_w_0_140_s_3_500 = '1.93750e-14*ic_cap*ic_cap+2.75000e-14*ic_cap+3.55000e-12'
+ mcm1l1_cc_w_1_120_s_0_140 = '-7.81250e-13*ic_cap*ic_cap+-3.75000e-13*ic_cap+1.15000e-10'
+ mcm1l1_cc_w_1_120_s_0_175 = '-6.06250e-13*ic_cap*ic_cap+-4.25000e-13*ic_cap+1.10000e-10'
+ mcm1l1_cc_w_1_120_s_0_210 = '-5.56250e-13*ic_cap*ic_cap+-3.00000e-13*ic_cap+1.04000e-10'
+ mcm1l1_cc_w_1_120_s_0_280 = '-4.06250e-13*ic_cap*ic_cap+-2.25000e-13*ic_cap+9.04000e-11'
+ mcm1l1_cc_w_1_120_s_0_350 = '-2.28125e-13*ic_cap*ic_cap+-1.12500e-13*ic_cap+7.72000e-11'
+ mcm1l1_cc_w_1_120_s_0_420 = '-1.75000e-13*ic_cap*ic_cap+-1.25000e-13*ic_cap+6.73000e-11'
+ mcm1l1_cc_w_1_120_s_0_560 = '-5.93750e-14*ic_cap*ic_cap+-1.25000e-14*ic_cap+5.26000e-11'
+ mcm1l1_cc_w_1_120_s_0_840 = '3.43750e-14*ic_cap*ic_cap+3.75000e-14*ic_cap+3.64000e-11'
+ mcm1l1_cc_w_1_120_s_1_540 = '5.62500e-14*ic_cap*ic_cap+5.00000e-14*ic_cap+1.97000e-11'
+ mcm1l1_cc_w_1_120_s_3_500 = '3.12500e-14*ic_cap*ic_cap+2.50000e-14*ic_cap+7.00000e-12'
+ mcm1l1_cf_w_0_140_s_0_140 = '-6.31250e-14*ic_cap*ic_cap+-5.25000e-14*ic_cap+7.43000e-12'
+ mcm1l1_cf_w_0_140_s_0_175 = '-9.62500e-14*ic_cap*ic_cap+-7.25000e-14*ic_cap+9.39000e-12'
+ mcm1l1_cf_w_0_140_s_0_210 = '-1.30625e-13*ic_cap*ic_cap+-9.25000e-14*ic_cap+1.13000e-11'
+ mcm1l1_cf_w_0_140_s_0_280 = '-1.84375e-13*ic_cap*ic_cap+-1.37500e-13*ic_cap+1.48000e-11'
+ mcm1l1_cf_w_0_140_s_0_350 = '-2.37500e-13*ic_cap*ic_cap+-1.75000e-13*ic_cap+1.81000e-11'
+ mcm1l1_cf_w_0_140_s_0_420 = '-2.81250e-13*ic_cap*ic_cap+-2.00000e-13*ic_cap+2.12000e-11'
+ mcm1l1_cf_w_0_140_s_0_560 = '-3.53125e-13*ic_cap*ic_cap+-2.37500e-13*ic_cap+2.65000e-11'
+ mcm1l1_cf_w_0_140_s_0_840 = '-4.40625e-13*ic_cap*ic_cap+-3.12500e-13*ic_cap+3.47000e-11'
+ mcm1l1_cf_w_0_140_s_1_540 = '-5.00000e-13*ic_cap*ic_cap+-3.50000e-13*ic_cap+4.62000e-11'
+ mcm1l1_cf_w_0_140_s_3_500 = '-4.96875e-13*ic_cap*ic_cap+-3.37500e-13*ic_cap+5.51000e-11'
+ mcm1l1_cf_w_1_120_s_0_140 = '-6.62500e-14*ic_cap*ic_cap+-5.25000e-14*ic_cap+7.56000e-12'
+ mcm1l1_cf_w_1_120_s_0_175 = '-9.84375e-14*ic_cap*ic_cap+-7.62500e-14*ic_cap+9.50000e-12'
+ mcm1l1_cf_w_1_120_s_0_210 = '-1.31563e-13*ic_cap*ic_cap+-9.37500e-14*ic_cap+1.14000e-11'
+ mcm1l1_cf_w_1_120_s_0_280 = '-1.87500e-13*ic_cap*ic_cap+-1.25000e-13*ic_cap+1.49000e-11'
+ mcm1l1_cf_w_1_120_s_0_350 = '-2.40625e-13*ic_cap*ic_cap+-1.62500e-13*ic_cap+1.82000e-11'
+ mcm1l1_cf_w_1_120_s_0_420 = '-2.87500e-13*ic_cap*ic_cap+-2.00000e-13*ic_cap+2.13000e-11'
+ mcm1l1_cf_w_1_120_s_0_560 = '-3.56250e-13*ic_cap*ic_cap+-2.50000e-13*ic_cap+2.66000e-11'
+ mcm1l1_cf_w_1_120_s_0_840 = '-4.43750e-13*ic_cap*ic_cap+-3.00000e-13*ic_cap+3.50000e-11'
+ mcm1l1_cf_w_1_120_s_1_540 = '-5.12500e-13*ic_cap*ic_cap+-3.75000e-13*ic_cap+4.74000e-11'
+ mcm1l1_cf_w_1_120_s_3_500 = '-5.18750e-13*ic_cap*ic_cap+-3.50000e-13*ic_cap+5.94000e-11'
+ mcm1l1d_ca_w_0_170_s_0_180 = '-2.50000e-06*ic_cap*ic_cap+-1.50000e-06*ic_cap+1.69000e-04'
+ mcm1l1d_ca_w_0_170_s_0_225 = '-2.50000e-06*ic_cap*ic_cap+-1.50000e-06*ic_cap+1.69000e-04'
+ mcm1l1d_ca_w_0_170_s_0_270 = '-2.50000e-06*ic_cap*ic_cap+-1.50000e-06*ic_cap+1.69000e-04'
+ mcm1l1d_ca_w_0_170_s_0_360 = '-2.50000e-06*ic_cap*ic_cap+-1.50000e-06*ic_cap+1.69000e-04'
+ mcm1l1d_ca_w_0_170_s_0_450 = '-2.50000e-06*ic_cap*ic_cap+-1.50000e-06*ic_cap+1.69000e-04'
+ mcm1l1d_ca_w_0_170_s_0_540 = '-2.50000e-06*ic_cap*ic_cap+-1.50000e-06*ic_cap+1.69000e-04'
+ mcm1l1d_ca_w_0_170_s_0_720 = '-2.50000e-06*ic_cap*ic_cap+-1.50000e-06*ic_cap+1.69000e-04'
+ mcm1l1d_ca_w_0_170_s_1_080 = '-2.50000e-06*ic_cap*ic_cap+-1.50000e-06*ic_cap+1.69000e-04'
+ mcm1l1d_ca_w_0_170_s_1_980 = '-2.50000e-06*ic_cap*ic_cap+-1.50000e-06*ic_cap+1.69000e-04'
+ mcm1l1d_ca_w_0_170_s_4_500 = '-2.50000e-06*ic_cap*ic_cap+-1.50000e-06*ic_cap+1.69000e-04'
+ mcm1l1d_ca_w_1_360_s_0_180 = '-2.50000e-06*ic_cap*ic_cap+-1.50000e-06*ic_cap+1.69000e-04'
+ mcm1l1d_ca_w_1_360_s_0_225 = '-2.50000e-06*ic_cap*ic_cap+-1.50000e-06*ic_cap+1.69000e-04'
+ mcm1l1d_ca_w_1_360_s_0_270 = '-2.50000e-06*ic_cap*ic_cap+-1.50000e-06*ic_cap+1.69000e-04'
+ mcm1l1d_ca_w_1_360_s_0_360 = '-2.50000e-06*ic_cap*ic_cap+-1.50000e-06*ic_cap+1.69000e-04'
+ mcm1l1d_ca_w_1_360_s_0_450 = '-2.50000e-06*ic_cap*ic_cap+-1.50000e-06*ic_cap+1.69000e-04'
+ mcm1l1d_ca_w_1_360_s_0_540 = '-2.50000e-06*ic_cap*ic_cap+-1.50000e-06*ic_cap+1.69000e-04'
+ mcm1l1d_ca_w_1_360_s_0_720 = '-2.50000e-06*ic_cap*ic_cap+-1.50000e-06*ic_cap+1.69000e-04'
+ mcm1l1d_ca_w_1_360_s_1_080 = '-2.50000e-06*ic_cap*ic_cap+-1.50000e-06*ic_cap+1.69000e-04'
+ mcm1l1d_ca_w_1_360_s_1_980 = '-2.50000e-06*ic_cap*ic_cap+-1.50000e-06*ic_cap+1.69000e-04'
+ mcm1l1d_ca_w_1_360_s_4_500 = '-2.50000e-06*ic_cap*ic_cap+-1.50000e-06*ic_cap+1.69000e-04'
+ mcm1l1d_cc_w_0_170_s_0_180 = '-5.90625e-13*ic_cap*ic_cap+-3.87500e-13*ic_cap+6.40000e-11'
+ mcm1l1d_cc_w_0_170_s_0_225 = '-3.68750e-13*ic_cap*ic_cap+-2.50000e-13*ic_cap+5.15000e-11'
+ mcm1l1d_cc_w_0_170_s_0_270 = '-2.34375e-13*ic_cap*ic_cap+-1.62500e-13*ic_cap+4.25000e-11'
+ mcm1l1d_cc_w_0_170_s_0_360 = '-7.81250e-14*ic_cap*ic_cap+-6.25000e-14*ic_cap+3.03000e-11'
+ mcm1l1d_cc_w_0_170_s_0_450 = '-3.12500e-15*ic_cap*ic_cap+-1.25000e-14*ic_cap+2.25000e-11'
+ mcm1l1d_cc_w_0_170_s_0_540 = '4.37500e-14*ic_cap*ic_cap+2.50000e-14*ic_cap+1.69000e-11'
+ mcm1l1d_cc_w_0_170_s_0_720 = '7.62500e-14*ic_cap*ic_cap+5.00000e-14*ic_cap+9.88000e-12'
+ mcm1l1d_cc_w_0_170_s_1_080 = '6.78125e-14*ic_cap*ic_cap+5.12500e-14*ic_cap+3.53000e-12'
+ mcm1l1d_cc_w_0_170_s_1_980 = '1.43750e-14*ic_cap*ic_cap+1.75000e-14*ic_cap+3.45000e-13'
+ mcm1l1d_cc_w_0_170_s_4_500 = '1.56250e-16*ic_cap*ic_cap+-3.12500e-15*ic_cap+3.00000e-14'
+ mcm1l1d_cc_w_1_360_s_0_180 = '-4.78125e-13*ic_cap*ic_cap+-2.62500e-13*ic_cap+6.78000e-11'
+ mcm1l1d_cc_w_1_360_s_0_225 = '-2.56250e-13*ic_cap*ic_cap+-1.75000e-13*ic_cap+5.46000e-11'
+ mcm1l1d_cc_w_1_360_s_0_270 = '-1.46875e-13*ic_cap*ic_cap+-8.75000e-14*ic_cap+4.53000e-11'
+ mcm1l1d_cc_w_1_360_s_0_450 = '7.18750e-14*ic_cap*ic_cap+3.75000e-14*ic_cap+2.40000e-11'
+ mcm1l1d_cc_w_1_360_s_0_540 = '9.37500e-14*ic_cap*ic_cap+5.00000e-14*ic_cap+1.83000e-11'
+ mcm1l1d_cc_w_1_360_s_0_720 = '1.21875e-13*ic_cap*ic_cap+8.75000e-14*ic_cap+1.07000e-11'
+ mcm1l1d_cc_w_1_360_s_1_080 = '8.75000e-14*ic_cap*ic_cap+7.50000e-14*ic_cap+3.90000e-12'
+ mcm1l1d_cc_w_1_360_s_1_980 = '2.21875e-14*ic_cap*ic_cap+2.00000e-14*ic_cap+3.50000e-13'
+ mcm1l1d_cc_w_1_360_s_4_500 = '1.56250e-15*ic_cap*ic_cap+6.25000e-15*ic_cap+1.29000e-26'
+ mcm1l1d_cf_w_0_170_s_0_180 = '-1.00000e-13*ic_cap*ic_cap+-7.50000e-14*ic_cap+1.41000e-11'
+ mcm1l1d_cf_w_0_170_s_0_225 = '-1.43750e-13*ic_cap*ic_cap+-1.00000e-13*ic_cap+1.72000e-11'
+ mcm1l1d_cf_w_0_170_s_0_270 = '-1.87500e-13*ic_cap*ic_cap+-1.25000e-13*ic_cap+2.01000e-11'
+ mcm1l1d_cf_w_0_170_s_0_360 = '-2.53125e-13*ic_cap*ic_cap+-1.62500e-13*ic_cap+2.53000e-11'
+ mcm1l1d_cf_w_0_170_s_0_450 = '-3.03125e-13*ic_cap*ic_cap+-2.12500e-13*ic_cap+2.96000e-11'
+ mcm1l1d_cf_w_0_170_s_0_540 = '-3.37500e-13*ic_cap*ic_cap+-2.25000e-13*ic_cap+3.32000e-11'
+ mcm1l1d_cf_w_0_170_s_0_720 = '-3.78125e-13*ic_cap*ic_cap+-2.62500e-13*ic_cap+3.85000e-11'
+ mcm1l1d_cf_w_0_170_s_1_080 = '-3.87500e-13*ic_cap*ic_cap+-2.75000e-13*ic_cap+4.41000e-11'
+ mcm1l1d_cf_w_0_170_s_1_980 = '-3.43750e-13*ic_cap*ic_cap+-2.50000e-13*ic_cap+4.72000e-11'
+ mcm1l1d_cf_w_0_170_s_4_500 = '-3.28125e-13*ic_cap*ic_cap+-2.37500e-13*ic_cap+4.75000e-11'
+ mcm1l1d_cf_w_1_360_s_0_180 = '-1.00000e-13*ic_cap*ic_cap+-7.50000e-14*ic_cap+1.40000e-11'
+ mcm1l1d_cf_w_1_360_s_0_225 = '-1.43750e-13*ic_cap*ic_cap+-1.00000e-13*ic_cap+1.71000e-11'
+ mcm1l1d_cf_w_1_360_s_0_270 = '-1.81250e-13*ic_cap*ic_cap+-1.25000e-13*ic_cap+2.00000e-11'
+ mcm1l1d_cf_w_1_360_s_0_360 = '-2.43750e-13*ic_cap*ic_cap+-1.75000e-13*ic_cap+2.52000e-11'
+ mcm1l1d_cf_w_1_360_s_0_450 = '-2.93750e-13*ic_cap*ic_cap+-2.00000e-13*ic_cap+2.97000e-11'
+ mcm1l1d_cf_w_1_360_s_0_540 = '-3.25000e-13*ic_cap*ic_cap+-2.25000e-13*ic_cap+3.34000e-11'
+ mcm1l1d_cf_w_1_360_s_0_720 = '-3.62500e-13*ic_cap*ic_cap+-2.50000e-13*ic_cap+3.90000e-11'
+ mcm1l1d_cf_w_1_360_s_1_080 = '-3.53125e-13*ic_cap*ic_cap+-2.62500e-13*ic_cap+4.49000e-11'
+ mcm1l1d_cf_w_1_360_s_1_980 = '-2.96875e-13*ic_cap*ic_cap+-2.12500e-13*ic_cap+4.83000e-11'
+ mcm1l1d_cf_w_1_360_s_4_500 = '-2.71875e-13*ic_cap*ic_cap+-1.87500e-13*ic_cap+4.86000e-11'
+ mcm1l1f_ca_w_0_170_s_0_180 = '-2.37500e-06*ic_cap*ic_cap+-1.50000e-06*ic_cap+1.51000e-04'
+ mcm1l1f_ca_w_0_170_s_0_225 = '-2.37500e-06*ic_cap*ic_cap+-1.50000e-06*ic_cap+1.51000e-04'
+ mcm1l1f_ca_w_0_170_s_0_270 = '-2.37500e-06*ic_cap*ic_cap+-1.50000e-06*ic_cap+1.51000e-04'
+ mcm1l1f_ca_w_0_170_s_0_360 = '-2.37500e-06*ic_cap*ic_cap+-1.50000e-06*ic_cap+1.51000e-04'
+ mcm1l1f_ca_w_0_170_s_0_450 = '-2.37500e-06*ic_cap*ic_cap+-1.50000e-06*ic_cap+1.51000e-04'
+ mcm1l1f_ca_w_0_170_s_0_540 = '-2.37500e-06*ic_cap*ic_cap+-1.50000e-06*ic_cap+1.51000e-04'
+ mcm1l1f_ca_w_0_170_s_0_720 = '-2.37500e-06*ic_cap*ic_cap+-1.50000e-06*ic_cap+1.51000e-04'
+ mcm1l1f_ca_w_0_170_s_1_080 = '-2.37500e-06*ic_cap*ic_cap+-1.50000e-06*ic_cap+1.51000e-04'
+ mcm1l1f_ca_w_0_170_s_1_980 = '-2.37500e-06*ic_cap*ic_cap+-1.50000e-06*ic_cap+1.51000e-04'
+ mcm1l1f_ca_w_0_170_s_4_500 = '-2.37500e-06*ic_cap*ic_cap+-1.50000e-06*ic_cap+1.51000e-04'
+ mcm1l1f_ca_w_1_360_s_0_180 = '-2.37500e-06*ic_cap*ic_cap+-1.50000e-06*ic_cap+1.51000e-04'
+ mcm1l1f_ca_w_1_360_s_0_225 = '-2.37500e-06*ic_cap*ic_cap+-1.50000e-06*ic_cap+1.51000e-04'
+ mcm1l1f_ca_w_1_360_s_0_270 = '-2.37500e-06*ic_cap*ic_cap+-1.50000e-06*ic_cap+1.51000e-04'
+ mcm1l1f_ca_w_1_360_s_0_360 = '-2.37500e-06*ic_cap*ic_cap+-1.50000e-06*ic_cap+1.51000e-04'
+ mcm1l1f_ca_w_1_360_s_0_450 = '-2.37500e-06*ic_cap*ic_cap+-1.50000e-06*ic_cap+1.51000e-04'
+ mcm1l1f_ca_w_1_360_s_0_540 = '-2.37500e-06*ic_cap*ic_cap+-1.50000e-06*ic_cap+1.51000e-04'
+ mcm1l1f_ca_w_1_360_s_0_720 = '-2.37500e-06*ic_cap*ic_cap+-1.50000e-06*ic_cap+1.51000e-04'
+ mcm1l1f_ca_w_1_360_s_1_080 = '-2.37500e-06*ic_cap*ic_cap+-1.50000e-06*ic_cap+1.51000e-04'
+ mcm1l1f_ca_w_1_360_s_1_980 = '-2.37500e-06*ic_cap*ic_cap+-1.50000e-06*ic_cap+1.51000e-04'
+ mcm1l1f_ca_w_1_360_s_4_500 = '-2.37500e-06*ic_cap*ic_cap+-1.50000e-06*ic_cap+1.51000e-04'
+ mcm1l1f_cc_w_0_170_s_0_180 = '-6.06250e-13*ic_cap*ic_cap+-3.75000e-13*ic_cap+6.64000e-11'
+ mcm1l1f_cc_w_0_170_s_0_225 = '-3.78125e-13*ic_cap*ic_cap+-2.62500e-13*ic_cap+5.39000e-11'
+ mcm1l1f_cc_w_0_170_s_0_270 = '-2.43750e-13*ic_cap*ic_cap+-1.75000e-13*ic_cap+4.51000e-11'
+ mcm1l1f_cc_w_0_170_s_0_360 = '-9.37500e-14*ic_cap*ic_cap+-7.50000e-14*ic_cap+3.31000e-11'
+ mcm1l1f_cc_w_0_170_s_0_450 = '-3.12500e-15*ic_cap*ic_cap+-1.25000e-14*ic_cap+2.52000e-11'
+ mcm1l1f_cc_w_0_170_s_0_540 = '4.06250e-14*ic_cap*ic_cap+1.25000e-14*ic_cap+1.96000e-11'
+ mcm1l1f_cc_w_0_170_s_0_720 = '8.43750e-14*ic_cap*ic_cap+3.75000e-14*ic_cap+1.22000e-11'
+ mcm1l1f_cc_w_0_170_s_1_080 = '8.18750e-14*ic_cap*ic_cap+5.50000e-14*ic_cap+5.14000e-12'
+ mcm1l1f_cc_w_0_170_s_1_980 = '2.87500e-14*ic_cap*ic_cap+2.75000e-14*ic_cap+7.00000e-13'
+ mcm1l1f_cc_w_0_170_s_4_500 = '2.81250e-15*ic_cap*ic_cap+-1.25000e-15*ic_cap'
+ mcm1l1f_cc_w_1_360_s_0_180 = '-4.68750e-13*ic_cap*ic_cap+-2.50000e-13*ic_cap+7.19000e-11'
+ mcm1l1f_cc_w_1_360_s_0_225 = '-2.53125e-13*ic_cap*ic_cap+-1.37500e-13*ic_cap+5.86000e-11'
+ mcm1l1f_cc_w_1_360_s_0_270 = '-1.25000e-13*ic_cap*ic_cap+-7.50000e-14*ic_cap+4.93000e-11'
+ mcm1l1f_cc_w_1_360_s_0_360 = '9.37500e-15*ic_cap*ic_cap+1.25000e-14*ic_cap+3.65000e-11'
+ mcm1l1f_cc_w_1_360_s_0_450 = '8.12500e-14*ic_cap*ic_cap+5.00000e-14*ic_cap+2.80000e-11'
+ mcm1l1f_cc_w_1_360_s_0_540 = '1.21875e-13*ic_cap*ic_cap+8.75000e-14*ic_cap+2.19000e-11'
+ mcm1l1f_cc_w_1_360_s_0_720 = '1.46875e-13*ic_cap*ic_cap+8.75000e-14*ic_cap+1.39000e-11'
+ mcm1l1f_cc_w_1_360_s_1_080 = '1.26563e-13*ic_cap*ic_cap+9.12500e-14*ic_cap+5.95000e-12'
+ mcm1l1f_cc_w_1_360_s_1_980 = '4.43750e-14*ic_cap*ic_cap+3.12500e-14*ic_cap+8.15000e-13'
+ mcm1l1f_cc_w_1_360_s_4_500 = '2.81250e-15*ic_cap*ic_cap+7.50000e-15*ic_cap'
+ mcm1l1f_cf_w_0_170_s_0_180 = '-1.06250e-13*ic_cap*ic_cap+-7.50000e-14*ic_cap+1.26000e-11'
+ mcm1l1f_cf_w_0_170_s_0_225 = '-1.40625e-13*ic_cap*ic_cap+-1.12500e-13*ic_cap+1.53000e-11'
+ mcm1l1f_cf_w_0_170_s_0_270 = '-1.81250e-13*ic_cap*ic_cap+-1.25000e-13*ic_cap+1.79000e-11'
+ mcm1l1f_cf_w_0_170_s_0_360 = '-2.40625e-13*ic_cap*ic_cap+-1.62500e-13*ic_cap+2.27000e-11'
+ mcm1l1f_cf_w_0_170_s_0_450 = '-2.93750e-13*ic_cap*ic_cap+-2.00000e-13*ic_cap+2.67000e-11'
+ mcm1l1f_cf_w_0_170_s_0_540 = '-3.31250e-13*ic_cap*ic_cap+-2.25000e-13*ic_cap+3.02000e-11'
+ mcm1l1f_cf_w_0_170_s_0_720 = '-3.78125e-13*ic_cap*ic_cap+-2.62500e-13*ic_cap+3.55000e-11'
+ mcm1l1f_cf_w_0_170_s_1_080 = '-3.96875e-13*ic_cap*ic_cap+-2.87500e-13*ic_cap+4.15000e-11'
+ mcm1l1f_cf_w_0_170_s_1_980 = '-3.59375e-13*ic_cap*ic_cap+-2.62500e-13*ic_cap+4.57000e-11'
+ mcm1l1f_cf_w_0_170_s_4_500 = '-3.28125e-13*ic_cap*ic_cap+-2.37500e-13*ic_cap+4.63000e-11'
+ mcm1l1f_cf_w_1_360_s_0_180 = '-1.00000e-13*ic_cap*ic_cap+-7.50000e-14*ic_cap+1.25000e-11'
+ mcm1l1f_cf_w_1_360_s_0_225 = '-1.43750e-13*ic_cap*ic_cap+-1.00000e-13*ic_cap+1.53000e-11'
+ mcm1l1f_cf_w_1_360_s_0_270 = '-1.75000e-13*ic_cap*ic_cap+-1.25000e-13*ic_cap+1.79000e-11'
+ mcm1l1f_cf_w_1_360_s_0_360 = '-2.40625e-13*ic_cap*ic_cap+-1.62500e-13*ic_cap+2.27000e-11'
+ mcm1l1f_cf_w_1_360_s_0_450 = '-2.93750e-13*ic_cap*ic_cap+-2.00000e-13*ic_cap+2.69000e-11'
+ mcm1l1f_cf_w_1_360_s_0_540 = '-3.31250e-13*ic_cap*ic_cap+-2.25000e-13*ic_cap+3.05000e-11'
+ mcm1l1f_cf_w_1_360_s_0_720 = '-3.65625e-13*ic_cap*ic_cap+-2.62500e-13*ic_cap+3.60000e-11'
+ mcm1l1f_cf_w_1_360_s_1_080 = '-3.71875e-13*ic_cap*ic_cap+-2.62500e-13*ic_cap+4.26000e-11'
+ mcm1l1f_cf_w_1_360_s_1_980 = '-3.12500e-13*ic_cap*ic_cap+-2.25000e-13*ic_cap+4.75000e-11'
+ mcm1l1f_cf_w_1_360_s_4_500 = '-2.71875e-13*ic_cap*ic_cap+-1.87500e-13*ic_cap+4.83000e-11'
+ mcm1l1p1_ca_w_0_170_s_0_180 = '-3.59375e-06*ic_cap*ic_cap+-2.12500e-06*ic_cap+2.08000e-04'
+ mcm1l1p1_ca_w_0_170_s_0_225 = '-3.59375e-06*ic_cap*ic_cap+-2.12500e-06*ic_cap+2.08000e-04'
+ mcm1l1p1_ca_w_0_170_s_0_270 = '-3.59375e-06*ic_cap*ic_cap+-2.12500e-06*ic_cap+2.08000e-04'
+ mcm1l1p1_ca_w_0_170_s_0_360 = '-3.59375e-06*ic_cap*ic_cap+-2.12500e-06*ic_cap+2.08000e-04'
+ mcm1l1p1_ca_w_0_170_s_0_450 = '-3.59375e-06*ic_cap*ic_cap+-2.12500e-06*ic_cap+2.08000e-04'
+ mcm1l1p1_ca_w_0_170_s_0_540 = '-3.59375e-06*ic_cap*ic_cap+-2.12500e-06*ic_cap+2.08000e-04'
+ mcm1l1p1_ca_w_0_170_s_0_720 = '-3.59375e-06*ic_cap*ic_cap+-2.12500e-06*ic_cap+2.08000e-04'
+ mcm1l1p1_ca_w_0_170_s_1_080 = '-3.59375e-06*ic_cap*ic_cap+-2.12500e-06*ic_cap+2.08000e-04'
+ mcm1l1p1_ca_w_0_170_s_1_980 = '-3.59375e-06*ic_cap*ic_cap+-2.12500e-06*ic_cap+2.08000e-04'
+ mcm1l1p1_ca_w_0_170_s_4_500 = '-3.59375e-06*ic_cap*ic_cap+-2.12500e-06*ic_cap+2.08000e-04'
+ mcm1l1p1_ca_w_1_360_s_0_180 = '-3.59375e-06*ic_cap*ic_cap+-2.12500e-06*ic_cap+2.08000e-04'
+ mcm1l1p1_ca_w_1_360_s_0_225 = '-3.59375e-06*ic_cap*ic_cap+-2.12500e-06*ic_cap+2.08000e-04'
+ mcm1l1p1_ca_w_1_360_s_0_270 = '-3.59375e-06*ic_cap*ic_cap+-2.12500e-06*ic_cap+2.08000e-04'
+ mcm1l1p1_ca_w_1_360_s_0_360 = '-3.59375e-06*ic_cap*ic_cap+-2.12500e-06*ic_cap+2.08000e-04'
+ mcm1l1p1_ca_w_1_360_s_0_450 = '-3.59375e-06*ic_cap*ic_cap+-2.12500e-06*ic_cap+2.08000e-04'
+ mcm1l1p1_ca_w_1_360_s_0_540 = '-3.59375e-06*ic_cap*ic_cap+-2.12500e-06*ic_cap+2.08000e-04'
+ mcm1l1p1_ca_w_1_360_s_0_720 = '-3.59375e-06*ic_cap*ic_cap+-2.12500e-06*ic_cap+2.08000e-04'
+ mcm1l1p1_ca_w_1_360_s_1_080 = '-3.59375e-06*ic_cap*ic_cap+-2.12500e-06*ic_cap+2.08000e-04'
+ mcm1l1p1_ca_w_1_360_s_1_980 = '-3.59375e-06*ic_cap*ic_cap+-2.12500e-06*ic_cap+2.08000e-04'
+ mcm1l1p1_ca_w_1_360_s_4_500 = '-3.59375e-06*ic_cap*ic_cap+-2.12500e-06*ic_cap+2.08000e-04'
+ mcm1l1p1_cc_w_0_170_s_0_180 = '-4.87500e-13*ic_cap*ic_cap+-3.25000e-13*ic_cap+5.98000e-11'
+ mcm1l1p1_cc_w_0_170_s_0_225 = '-2.68750e-13*ic_cap*ic_cap+-2.00000e-13*ic_cap+4.72000e-11'
+ mcm1l1p1_cc_w_0_170_s_0_270 = '-1.28125e-13*ic_cap*ic_cap+-1.12500e-13*ic_cap+3.81000e-11'
+ mcm1l1p1_cc_w_0_170_s_0_360 = '1.87500e-14*ic_cap*ic_cap+-2.50000e-14*ic_cap+2.60000e-11'
+ mcm1l1p1_cc_w_0_170_s_0_450 = '9.37500e-14*ic_cap*ic_cap+5.00000e-14*ic_cap+1.82000e-11'
+ mcm1l1p1_cc_w_0_170_s_0_540 = '1.25000e-13*ic_cap*ic_cap+5.00000e-14*ic_cap+1.30000e-11'
+ mcm1l1p1_cc_w_0_170_s_0_720 = '1.30313e-13*ic_cap*ic_cap+7.62500e-14*ic_cap+6.77000e-12'
+ mcm1l1p1_cc_w_0_170_s_1_080 = '8.21875e-14*ic_cap*ic_cap+5.87500e-14*ic_cap+1.87000e-12'
+ mcm1l1p1_cc_w_0_170_s_1_980 = '1.23438e-14*ic_cap*ic_cap+1.31250e-14*ic_cap+9.50000e-14'
+ mcm1l1p1_cc_w_0_170_s_4_500 = '9.37500e-16*ic_cap*ic_cap+2.50000e-15*ic_cap'
+ mcm1l1p1_cc_w_1_360_s_0_180 = '-3.62500e-13*ic_cap*ic_cap+-2.25000e-13*ic_cap+6.16000e-11'
+ mcm1l1p1_cc_w_1_360_s_0_225 = '-1.50000e-13*ic_cap*ic_cap+-1.25000e-13*ic_cap+4.86000e-11'
+ mcm1l1p1_cc_w_1_360_s_0_270 = '-2.81250e-14*ic_cap*ic_cap+-3.75000e-14*ic_cap+3.93000e-11'
+ mcm1l1p1_cc_w_1_360_s_0_360 = '9.06250e-14*ic_cap*ic_cap+3.75000e-14*ic_cap+2.69000e-11'
+ mcm1l1p1_cc_w_1_360_s_0_450 = '1.59375e-13*ic_cap*ic_cap+8.75000e-14*ic_cap+1.88000e-11'
+ mcm1l1p1_cc_w_1_360_s_0_540 = '1.75000e-13*ic_cap*ic_cap+1.00000e-13*ic_cap+1.35000e-11'
+ mcm1l1p1_cc_w_1_360_s_0_720 = '1.67187e-13*ic_cap*ic_cap+1.06250e-13*ic_cap+7.00000e-12'
+ mcm1l1p1_cc_w_1_360_s_1_080 = '1.00000e-13*ic_cap*ic_cap+7.50000e-14*ic_cap+1.95000e-12'
+ mcm1l1p1_cc_w_1_360_s_1_980 = '1.09375e-14*ic_cap*ic_cap+6.25000e-15*ic_cap+1.50000e-13'
+ mcm1l1p1_cc_w_1_360_s_4_500 = '1.56250e-15*ic_cap*ic_cap+6.25000e-15*ic_cap'
+ mcm1l1p1_cf_w_0_170_s_0_180 = '-1.78125e-13*ic_cap*ic_cap+-1.12500e-13*ic_cap+1.73000e-11'
+ mcm1l1p1_cf_w_0_170_s_0_225 = '-2.31250e-13*ic_cap*ic_cap+-1.50000e-13*ic_cap+2.09000e-11'
+ mcm1l1p1_cf_w_0_170_s_0_270 = '-2.87500e-13*ic_cap*ic_cap+-1.75000e-13*ic_cap+2.43000e-11'
+ mcm1l1p1_cf_w_0_170_s_0_360 = '-3.75000e-13*ic_cap*ic_cap+-2.25000e-13*ic_cap+3.03000e-11'
+ mcm1l1p1_cf_w_0_170_s_0_450 = '-4.40625e-13*ic_cap*ic_cap+-2.62500e-13*ic_cap+3.51000e-11'
+ mcm1l1p1_cf_w_0_170_s_0_540 = '-4.75000e-13*ic_cap*ic_cap+-3.00000e-13*ic_cap+3.89000e-11'
+ mcm1l1p1_cf_w_0_170_s_0_720 = '-5.00000e-13*ic_cap*ic_cap+-3.25000e-13*ic_cap+4.40000e-11'
+ mcm1l1p1_cf_w_0_170_s_1_080 = '-4.71875e-13*ic_cap*ic_cap+-3.12500e-13*ic_cap+4.85000e-11'
+ mcm1l1p1_cf_w_0_170_s_1_980 = '-4.12500e-13*ic_cap*ic_cap+-2.75000e-13*ic_cap+5.03000e-11'
+ mcm1l1p1_cf_w_0_170_s_4_500 = '-4.03125e-13*ic_cap*ic_cap+-2.62500e-13*ic_cap+5.04000e-11'
+ mcm1l1p1_cf_w_1_360_s_0_180 = '-1.71875e-13*ic_cap*ic_cap+-1.12500e-13*ic_cap+1.71000e-11'
+ mcm1l1p1_cf_w_1_360_s_0_225 = '-2.31250e-13*ic_cap*ic_cap+-1.50000e-13*ic_cap+2.08000e-11'
+ mcm1l1p1_cf_w_1_360_s_0_270 = '-2.87500e-13*ic_cap*ic_cap+-1.75000e-13*ic_cap+2.43000e-11'
+ mcm1l1p1_cf_w_1_360_s_0_360 = '-3.65625e-13*ic_cap*ic_cap+-2.12500e-13*ic_cap+3.02000e-11'
+ mcm1l1p1_cf_w_1_360_s_0_450 = '-4.28125e-13*ic_cap*ic_cap+-2.62500e-13*ic_cap+3.52000e-11'
+ mcm1l1p1_cf_w_1_360_s_0_540 = '-4.59375e-13*ic_cap*ic_cap+-2.87500e-13*ic_cap+3.90000e-11'
+ mcm1l1p1_cf_w_1_360_s_0_720 = '-4.78125e-13*ic_cap*ic_cap+-3.12500e-13*ic_cap+4.43000e-11'
+ mcm1l1p1_cf_w_1_360_s_1_080 = '-4.40625e-13*ic_cap*ic_cap+-2.87500e-13*ic_cap+4.90000e-11'
+ mcm1l1p1_cf_w_1_360_s_1_980 = '-3.59375e-13*ic_cap*ic_cap+-2.37500e-13*ic_cap+5.08000e-11'
+ mcm1l1p1_cf_w_1_360_s_4_500 = '-3.43750e-13*ic_cap*ic_cap+-2.25000e-13*ic_cap+5.08000e-11'
+ mcm1p1_ca_w_0_140_s_0_140 = '-6.81250e-07*ic_cap*ic_cap+-4.00000e-07*ic_cap+4.48000e-05'
+ mcm1p1_ca_w_0_140_s_0_175 = '-6.81250e-07*ic_cap*ic_cap+-4.00000e-07*ic_cap+4.48000e-05'
+ mcm1p1_ca_w_0_140_s_0_210 = '-6.81250e-07*ic_cap*ic_cap+-4.00000e-07*ic_cap+4.48000e-05'
+ mcm1p1_ca_w_0_140_s_0_280 = '-6.81250e-07*ic_cap*ic_cap+-4.00000e-07*ic_cap+4.48000e-05'
+ mcm1p1_ca_w_0_140_s_0_350 = '-6.81250e-07*ic_cap*ic_cap+-4.00000e-07*ic_cap+4.48000e-05'
+ mcm1p1_ca_w_0_140_s_0_420 = '-6.81250e-07*ic_cap*ic_cap+-4.00000e-07*ic_cap+4.48000e-05'
+ mcm1p1_ca_w_0_140_s_0_560 = '-6.81250e-07*ic_cap*ic_cap+-4.00000e-07*ic_cap+4.48000e-05'
+ mcm1p1_ca_w_0_140_s_0_840 = '-6.81250e-07*ic_cap*ic_cap+-4.00000e-07*ic_cap+4.48000e-05'
+ mcm1p1_ca_w_0_140_s_1_540 = '-6.81250e-07*ic_cap*ic_cap+-4.00000e-07*ic_cap+4.48000e-05'
+ mcm1p1_ca_w_0_140_s_3_500 = '-6.81250e-07*ic_cap*ic_cap+-4.00000e-07*ic_cap+4.48000e-05'
+ mcm1p1_ca_w_1_120_s_0_140 = '-6.81250e-07*ic_cap*ic_cap+-4.00000e-07*ic_cap+4.48000e-05'
+ mcm1p1_ca_w_1_120_s_0_175 = '-6.81250e-07*ic_cap*ic_cap+-4.00000e-07*ic_cap+4.48000e-05'
+ mcm1p1_ca_w_1_120_s_0_210 = '-6.81250e-07*ic_cap*ic_cap+-4.00000e-07*ic_cap+4.48000e-05'
+ mcm1p1_ca_w_1_120_s_0_280 = '-6.81250e-07*ic_cap*ic_cap+-4.00000e-07*ic_cap+4.48000e-05'
+ mcm1p1_ca_w_1_120_s_0_350 = '-6.81250e-07*ic_cap*ic_cap+-4.00000e-07*ic_cap+4.48000e-05'
+ mcm1p1_ca_w_1_120_s_0_420 = '-6.81250e-07*ic_cap*ic_cap+-4.00000e-07*ic_cap+4.48000e-05'
+ mcm1p1_ca_w_1_120_s_0_560 = '-6.81250e-07*ic_cap*ic_cap+-4.00000e-07*ic_cap+4.48000e-05'
+ mcm1p1_ca_w_1_120_s_0_840 = '-6.81250e-07*ic_cap*ic_cap+-4.00000e-07*ic_cap+4.48000e-05'
+ mcm1p1_ca_w_1_120_s_1_540 = '-6.81250e-07*ic_cap*ic_cap+-4.00000e-07*ic_cap+4.48000e-05'
+ mcm1p1_ca_w_1_120_s_3_500 = '-6.81250e-07*ic_cap*ic_cap+-4.00000e-07*ic_cap+4.48000e-05'
+ mcm1p1_cc_w_0_140_s_0_140 = '-9.12500e-13*ic_cap*ic_cap+-4.75000e-13*ic_cap+1.03000e-10'
+ mcm1p1_cc_w_0_140_s_0_175 = '-8.56250e-13*ic_cap*ic_cap+-5.00000e-13*ic_cap+1.01000e-10'
+ mcm1p1_cc_w_0_140_s_0_210 = '-6.81250e-13*ic_cap*ic_cap+-4.75000e-13*ic_cap+9.50000e-11'
+ mcm1p1_cc_w_0_140_s_0_280 = '-5.62500e-13*ic_cap*ic_cap+-3.00000e-13*ic_cap+8.43000e-11'
+ mcm1p1_cc_w_0_140_s_0_350 = '-4.00000e-13*ic_cap*ic_cap+-2.75000e-13*ic_cap+7.26000e-11'
+ mcm1p1_cc_w_0_140_s_0_420 = '-2.75000e-13*ic_cap*ic_cap+-2.25000e-13*ic_cap+6.31000e-11'
+ mcm1p1_cc_w_0_140_s_0_560 = '-1.50000e-13*ic_cap*ic_cap+-1.00000e-13*ic_cap+5.03000e-11'
+ mcm1p1_cc_w_0_140_s_0_840 = '-2.50000e-14*ic_cap*ic_cap+-2.50000e-14*ic_cap+3.57000e-11'
+ mcm1p1_cc_w_0_140_s_1_540 = '5.93750e-14*ic_cap*ic_cap+3.75000e-14*ic_cap+1.96000e-11'
+ mcm1p1_cc_w_0_140_s_3_500 = '6.09375e-14*ic_cap*ic_cap+4.37500e-14*ic_cap+6.59000e-12'
+ mcm1p1_cc_w_1_120_s_0_140 = '-7.81250e-13*ic_cap*ic_cap+-3.75000e-13*ic_cap+1.25000e-10'
+ mcm1p1_cc_w_1_120_s_0_175 = '-7.18750e-13*ic_cap*ic_cap+-3.75000e-13*ic_cap+1.21000e-10'
+ mcm1p1_cc_w_1_120_s_0_210 = '-5.62500e-13*ic_cap*ic_cap+-2.50000e-13*ic_cap+1.14000e-10'
+ mcm1p1_cc_w_1_120_s_0_280 = '-4.37500e-13*ic_cap*ic_cap+-2.50000e-13*ic_cap+1.01000e-10'
+ mcm1p1_cc_w_1_120_s_0_350 = '-2.96875e-13*ic_cap*ic_cap+-1.87500e-13*ic_cap+8.83000e-11'
+ mcm1p1_cc_w_1_120_s_0_420 = '-1.96875e-13*ic_cap*ic_cap+-1.62500e-13*ic_cap+7.77000e-11'
+ mcm1p1_cc_w_1_120_s_0_560 = '-7.81250e-14*ic_cap*ic_cap+-6.25000e-14*ic_cap+6.27000e-11'
+ mcm1p1_cc_w_1_120_s_0_840 = '1.87500e-14*ic_cap*ic_cap+4.59000e-11'
+ mcm1p1_cc_w_1_120_s_1_540 = '8.75000e-14*ic_cap*ic_cap+5.00000e-14*ic_cap+2.71000e-11'
+ mcm1p1_cc_w_1_120_s_3_500 = '8.12500e-14*ic_cap*ic_cap+5.00000e-14*ic_cap+1.07000e-11'
+ mcm1p1_cf_w_0_140_s_0_140 = '-2.03125e-14*ic_cap*ic_cap+-1.37500e-14*ic_cap+3.09000e-12'
+ mcm1p1_cf_w_0_140_s_0_175 = '-3.18750e-14*ic_cap*ic_cap+-2.00000e-14*ic_cap+3.87000e-12'
+ mcm1p1_cf_w_0_140_s_0_210 = '-4.37500e-14*ic_cap*ic_cap+-2.75000e-14*ic_cap+4.64000e-12'
+ mcm1p1_cf_w_0_140_s_0_280 = '-6.56250e-14*ic_cap*ic_cap+-4.00000e-14*ic_cap+6.14000e-12'
+ mcm1p1_cf_w_0_140_s_0_350 = '-8.78125e-14*ic_cap*ic_cap+-5.37500e-14*ic_cap+7.60000e-12'
+ mcm1p1_cf_w_0_140_s_0_420 = '-1.07813e-13*ic_cap*ic_cap+-6.87500e-14*ic_cap+9.06000e-12'
+ mcm1p1_cf_w_0_140_s_0_560 = '-1.45313e-13*ic_cap*ic_cap+-8.87500e-14*ic_cap+1.17000e-11'
+ mcm1p1_cf_w_0_140_s_0_840 = '-2.06250e-13*ic_cap*ic_cap+-1.25000e-13*ic_cap+1.65000e-11'
+ mcm1p1_cf_w_0_140_s_1_540 = '-2.96875e-13*ic_cap*ic_cap+-1.87500e-13*ic_cap+2.55000e-11'
+ mcm1p1_cf_w_0_140_s_3_500 = '-3.31250e-13*ic_cap*ic_cap+-2.25000e-13*ic_cap+3.65000e-11'
+ mcm1p1_cf_w_1_120_s_0_140 = '-2.28125e-14*ic_cap*ic_cap+-1.37500e-14*ic_cap+3.22000e-12'
+ mcm1p1_cf_w_1_120_s_0_175 = '-3.46875e-14*ic_cap*ic_cap+-2.12500e-14*ic_cap+4.00000e-12'
+ mcm1p1_cf_w_1_120_s_0_210 = '-4.71875e-14*ic_cap*ic_cap+-2.87500e-14*ic_cap+4.77000e-12'
+ mcm1p1_cf_w_1_120_s_0_280 = '-6.78125e-14*ic_cap*ic_cap+-4.12500e-14*ic_cap+6.26000e-12'
+ mcm1p1_cf_w_1_120_s_0_350 = '-8.87500e-14*ic_cap*ic_cap+-5.50000e-14*ic_cap+7.72000e-12'
+ mcm1p1_cf_w_1_120_s_0_420 = '-1.10625e-13*ic_cap*ic_cap+-6.75000e-14*ic_cap+9.16000e-12'
+ mcm1p1_cf_w_1_120_s_0_560 = '-1.45000e-13*ic_cap*ic_cap+-9.00000e-14*ic_cap+1.18000e-11'
+ mcm1p1_cf_w_1_120_s_0_840 = '-2.15625e-13*ic_cap*ic_cap+-1.37500e-13*ic_cap+1.68000e-11'
+ mcm1p1_cf_w_1_120_s_1_540 = '-2.96875e-13*ic_cap*ic_cap+-1.87500e-13*ic_cap+2.61000e-11'
+ mcm1p1_cf_w_1_120_s_3_500 = '-3.43750e-13*ic_cap*ic_cap+-2.25000e-13*ic_cap+3.92000e-11'
+ mcm1p1f_ca_w_0_150_s_0_210 = '-2.09375e-06*ic_cap*ic_cap+-1.12500e-06*ic_cap+1.51000e-04'
+ mcm1p1f_ca_w_0_150_s_0_263 = '-2.09375e-06*ic_cap*ic_cap+-1.12500e-06*ic_cap+1.51000e-04'
+ mcm1p1f_ca_w_0_150_s_0_315 = '-2.09375e-06*ic_cap*ic_cap+-1.12500e-06*ic_cap+1.51000e-04'
+ mcm1p1f_ca_w_0_150_s_0_420 = '-2.09375e-06*ic_cap*ic_cap+-1.12500e-06*ic_cap+1.51000e-04'
+ mcm1p1f_ca_w_0_150_s_0_525 = '-2.09375e-06*ic_cap*ic_cap+-1.12500e-06*ic_cap+1.51000e-04'
+ mcm1p1f_ca_w_0_150_s_0_630 = '-2.09375e-06*ic_cap*ic_cap+-1.12500e-06*ic_cap+1.51000e-04'
+ mcm1p1f_ca_w_0_150_s_0_840 = '-2.09375e-06*ic_cap*ic_cap+-1.12500e-06*ic_cap+1.51000e-04'
+ mcm1p1f_ca_w_0_150_s_1_260 = '-2.09375e-06*ic_cap*ic_cap+-1.12500e-06*ic_cap+1.51000e-04'
+ mcm1p1f_ca_w_0_150_s_2_310 = '-2.09375e-06*ic_cap*ic_cap+-1.12500e-06*ic_cap+1.51000e-04'
+ mcm1p1f_ca_w_0_150_s_5_250 = '-2.09375e-06*ic_cap*ic_cap+-1.12500e-06*ic_cap+1.51000e-04'
+ mcm1p1f_ca_w_1_200_s_0_210 = '-2.09375e-06*ic_cap*ic_cap+-1.12500e-06*ic_cap+1.51000e-04'
+ mcm1p1f_ca_w_1_200_s_0_263 = '-2.09375e-06*ic_cap*ic_cap+-1.12500e-06*ic_cap+1.51000e-04'
+ mcm1p1f_ca_w_1_200_s_0_315 = '-2.09375e-06*ic_cap*ic_cap+-1.12500e-06*ic_cap+1.51000e-04'
+ mcm1p1f_ca_w_1_200_s_0_420 = '-2.09375e-06*ic_cap*ic_cap+-1.12500e-06*ic_cap+1.51000e-04'
+ mcm1p1f_ca_w_1_200_s_0_525 = '-2.09375e-06*ic_cap*ic_cap+-1.12500e-06*ic_cap+1.51000e-04'
+ mcm1p1f_ca_w_1_200_s_0_630 = '-2.09375e-06*ic_cap*ic_cap+-1.12500e-06*ic_cap+1.51000e-04'
+ mcm1p1f_ca_w_1_200_s_0_840 = '-2.09375e-06*ic_cap*ic_cap+-1.12500e-06*ic_cap+1.51000e-04'
+ mcm1p1f_ca_w_1_200_s_1_260 = '-2.09375e-06*ic_cap*ic_cap+-1.12500e-06*ic_cap+1.51000e-04'
+ mcm1p1f_ca_w_1_200_s_2_310 = '-2.09375e-06*ic_cap*ic_cap+-1.12500e-06*ic_cap+1.51000e-04'
+ mcm1p1f_ca_w_1_200_s_5_250 = '-2.09375e-06*ic_cap*ic_cap+-1.12500e-06*ic_cap+1.51000e-04'
+ mcm1p1f_cc_w_0_150_s_0_210 = '-4.78125e-13*ic_cap*ic_cap+-2.62500e-13*ic_cap+6.98000e-11'
+ mcm1p1f_cc_w_0_150_s_0_263 = '-2.75000e-13*ic_cap*ic_cap+-1.50000e-13*ic_cap+5.50000e-11'
+ mcm1p1f_cc_w_0_150_s_0_315 = '-1.53125e-13*ic_cap*ic_cap+-8.75000e-14*ic_cap+4.48000e-11'
+ mcm1p1f_cc_w_0_150_s_0_420 = '-2.18750e-14*ic_cap*ic_cap+-1.25000e-14*ic_cap+3.17000e-11'
+ mcm1p1f_cc_w_0_150_s_0_525 = '4.37500e-14*ic_cap*ic_cap+2.50000e-14*ic_cap+2.33000e-11'
+ mcm1p1f_cc_w_0_150_s_0_630 = '7.50000e-14*ic_cap*ic_cap+5.00000e-14*ic_cap+1.75000e-11'
+ mcm1p1f_cc_w_0_150_s_0_840 = '9.37500e-14*ic_cap*ic_cap+7.50000e-14*ic_cap+1.03000e-11'
+ mcm1p1f_cc_w_0_150_s_1_260 = '7.78125e-14*ic_cap*ic_cap+5.37500e-14*ic_cap+3.78000e-12'
+ mcm1p1f_cc_w_0_150_s_2_310 = '2.12500e-14*ic_cap*ic_cap+1.87500e-14*ic_cap+3.70000e-13'
+ mcm1p1f_cc_w_0_150_s_5_250 = '-1.09375e-15*ic_cap*ic_cap+-6.25000e-16*ic_cap+4.00000e-14'
+ mcm1p1f_cc_w_1_200_s_0_210 = '-3.65625e-13*ic_cap*ic_cap+-1.87500e-13*ic_cap+7.52000e-11'
+ mcm1p1f_cc_w_1_200_s_0_263 = '-1.62500e-13*ic_cap*ic_cap+-7.50000e-14*ic_cap+5.93000e-11'
+ mcm1p1f_cc_w_1_200_s_0_315 = '-5.93750e-14*ic_cap*ic_cap+-1.25000e-14*ic_cap+4.87000e-11'
+ mcm1p1f_cc_w_1_200_s_0_420 = '6.25000e-14*ic_cap*ic_cap+5.00000e-14*ic_cap+3.46000e-11'
+ mcm1p1f_cc_w_1_200_s_0_525 = '1.12500e-13*ic_cap*ic_cap+7.50000e-14*ic_cap+2.57000e-11'
+ mcm1p1f_cc_w_1_200_s_0_630 = '1.34375e-13*ic_cap*ic_cap+8.75000e-14*ic_cap+1.95000e-11'
+ mcm1p1f_cc_w_1_200_s_0_840 = '1.43750e-13*ic_cap*ic_cap+1.00000e-13*ic_cap+1.16000e-11'
+ mcm1p1f_cc_w_1_200_s_1_260 = '1.08438e-13*ic_cap*ic_cap+7.62500e-14*ic_cap+4.37000e-12'
+ mcm1p1f_cc_w_1_200_s_2_310 = '2.96875e-14*ic_cap*ic_cap+2.37500e-14*ic_cap+4.60000e-13'
+ mcm1p1f_cc_w_1_200_s_5_250 = '2.18750e-15*ic_cap*ic_cap+3.75000e-15*ic_cap'
+ mcm1p1f_cf_w_0_150_s_0_210 = '-1.40625e-13*ic_cap*ic_cap+-8.75000e-14*ic_cap+1.48000e-11'
+ mcm1p1f_cf_w_0_150_s_0_263 = '-1.84375e-13*ic_cap*ic_cap+-1.12500e-13*ic_cap+1.80000e-11'
+ mcm1p1f_cf_w_0_150_s_0_315 = '-2.18750e-13*ic_cap*ic_cap+-1.25000e-13*ic_cap+2.09000e-11'
+ mcm1p1f_cf_w_0_150_s_0_420 = '-2.84375e-13*ic_cap*ic_cap+-1.62500e-13*ic_cap+2.64000e-11'
+ mcm1p1f_cf_w_0_150_s_0_525 = '-3.28125e-13*ic_cap*ic_cap+-1.87500e-13*ic_cap+3.09000e-11'
+ mcm1p1f_cf_w_0_150_s_0_630 = '-3.53125e-13*ic_cap*ic_cap+-2.12500e-13*ic_cap+3.45000e-11'
+ mcm1p1f_cf_w_0_150_s_0_840 = '-3.90625e-13*ic_cap*ic_cap+-2.37500e-13*ic_cap+4.00000e-11'
+ mcm1p1f_cf_w_0_150_s_1_260 = '-3.90625e-13*ic_cap*ic_cap+-2.37500e-13*ic_cap+4.57000e-11'
+ mcm1p1f_cf_w_0_150_s_2_310 = '-3.37500e-13*ic_cap*ic_cap+-2.00000e-13*ic_cap+4.88000e-11'
+ mcm1p1f_cf_w_0_150_s_5_250 = '-3.15625e-13*ic_cap*ic_cap+-1.87500e-13*ic_cap+4.92000e-11'
+ mcm1p1f_cf_w_1_200_s_0_210 = '-1.40625e-13*ic_cap*ic_cap+-8.75000e-14*ic_cap+1.47000e-11'
+ mcm1p1f_cf_w_1_200_s_0_263 = '-1.75000e-13*ic_cap*ic_cap+-1.00000e-13*ic_cap+1.79000e-11'
+ mcm1p1f_cf_w_1_200_s_0_315 = '-2.12500e-13*ic_cap*ic_cap+-1.25000e-13*ic_cap+2.09000e-11'
+ mcm1p1f_cf_w_1_200_s_0_420 = '-2.78125e-13*ic_cap*ic_cap+-1.62500e-13*ic_cap+2.64000e-11'
+ mcm1p1f_cf_w_1_200_s_0_525 = '-3.21875e-13*ic_cap*ic_cap+-1.87500e-13*ic_cap+3.11000e-11'
+ mcm1p1f_cf_w_1_200_s_0_630 = '-3.50000e-13*ic_cap*ic_cap+-2.00000e-13*ic_cap+3.49000e-11'
+ mcm1p1f_cf_w_1_200_s_0_840 = '-3.81250e-13*ic_cap*ic_cap+-2.25000e-13*ic_cap+4.07000e-11'
+ mcm1p1f_cf_w_1_200_s_1_260 = '-3.75000e-13*ic_cap*ic_cap+-2.25000e-13*ic_cap+4.70000e-11'
+ mcm1p1f_cf_w_1_200_s_2_310 = '-3.00000e-13*ic_cap*ic_cap+-1.75000e-13*ic_cap+5.07000e-11'
+ mcm1p1f_cf_w_1_200_s_5_250 = '-2.68750e-13*ic_cap*ic_cap+-1.50000e-13*ic_cap+5.11000e-11'
+ mcm2d_ca_w_0_140_s_0_140 = '-2.15625e-07*ic_cap*ic_cap+-1.37500e-07*ic_cap+2.08000e-05'
+ mcm2d_ca_w_0_140_s_0_175 = '-2.15625e-07*ic_cap*ic_cap+-1.37500e-07*ic_cap+2.08000e-05'
+ mcm2d_ca_w_0_140_s_0_210 = '-2.15625e-07*ic_cap*ic_cap+-1.37500e-07*ic_cap+2.08000e-05'
+ mcm2d_ca_w_0_140_s_0_280 = '-2.15625e-07*ic_cap*ic_cap+-1.37500e-07*ic_cap+2.08000e-05'
+ mcm2d_ca_w_0_140_s_0_350 = '-2.15625e-07*ic_cap*ic_cap+-1.37500e-07*ic_cap+2.08000e-05'
+ mcm2d_ca_w_0_140_s_0_420 = '-2.15625e-07*ic_cap*ic_cap+-1.37500e-07*ic_cap+2.08000e-05'
+ mcm2d_ca_w_0_140_s_0_560 = '-2.15625e-07*ic_cap*ic_cap+-1.37500e-07*ic_cap+2.08000e-05'
+ mcm2d_ca_w_0_140_s_0_840 = '-2.15625e-07*ic_cap*ic_cap+-1.37500e-07*ic_cap+2.08000e-05'
+ mcm2d_ca_w_0_140_s_1_540 = '-2.15625e-07*ic_cap*ic_cap+-1.37500e-07*ic_cap+2.08000e-05'
+ mcm2d_ca_w_0_140_s_3_500 = '-2.15625e-07*ic_cap*ic_cap+-1.37500e-07*ic_cap+2.08000e-05'
+ mcm2d_ca_w_1_120_s_0_140 = '-2.15625e-07*ic_cap*ic_cap+-1.37500e-07*ic_cap+2.08000e-05'
+ mcm2d_ca_w_1_120_s_0_175 = '-2.15625e-07*ic_cap*ic_cap+-1.37500e-07*ic_cap+2.08000e-05'
+ mcm2d_ca_w_1_120_s_0_210 = '-2.15625e-07*ic_cap*ic_cap+-1.37500e-07*ic_cap+2.08000e-05'
+ mcm2d_ca_w_1_120_s_0_280 = '-2.15625e-07*ic_cap*ic_cap+-1.37500e-07*ic_cap+2.08000e-05'
+ mcm2d_ca_w_1_120_s_0_350 = '-2.15625e-07*ic_cap*ic_cap+-1.37500e-07*ic_cap+2.08000e-05'
+ mcm2d_ca_w_1_120_s_0_420 = '-2.15625e-07*ic_cap*ic_cap+-1.37500e-07*ic_cap+2.08000e-05'
+ mcm2d_ca_w_1_120_s_0_560 = '-2.15625e-07*ic_cap*ic_cap+-1.37500e-07*ic_cap+2.08000e-05'
+ mcm2d_ca_w_1_120_s_0_840 = '-2.15625e-07*ic_cap*ic_cap+-1.37500e-07*ic_cap+2.08000e-05'
+ mcm2d_ca_w_1_120_s_1_540 = '-2.15625e-07*ic_cap*ic_cap+-1.37500e-07*ic_cap+2.08000e-05'
+ mcm2d_ca_w_1_120_s_3_500 = '-2.15625e-07*ic_cap*ic_cap+-1.37500e-07*ic_cap+2.08000e-05'
+ mcm2d_cc_w_0_140_s_0_140 = '-9.12500e-13*ic_cap*ic_cap+-5.00000e-13*ic_cap+1.05000e-10'
+ mcm2d_cc_w_0_140_s_0_175 = '-8.59375e-13*ic_cap*ic_cap+-5.62500e-13*ic_cap+1.03000e-10'
+ mcm2d_cc_w_0_140_s_0_210 = '-7.68750e-13*ic_cap*ic_cap+-4.25000e-13*ic_cap+9.82000e-11'
+ mcm2d_cc_w_0_140_s_0_280 = '-6.34375e-13*ic_cap*ic_cap+-3.87500e-13*ic_cap+8.83000e-11'
+ mcm2d_cc_w_0_140_s_0_350 = '-4.84375e-13*ic_cap*ic_cap+-3.37500e-13*ic_cap+7.70000e-11'
+ mcm2d_cc_w_0_140_s_0_420 = '-3.62500e-13*ic_cap*ic_cap+-2.50000e-13*ic_cap+6.74000e-11'
+ mcm2d_cc_w_0_140_s_0_560 = '-2.21875e-13*ic_cap*ic_cap+-1.62500e-13*ic_cap+5.52000e-11'
+ mcm2d_cc_w_0_140_s_0_840 = '-1.06250e-13*ic_cap*ic_cap+-7.50000e-14*ic_cap+4.16000e-11'
+ mcm2d_cc_w_0_140_s_3_500 = '4.37500e-14*ic_cap*ic_cap+2.50000e-14*ic_cap+1.14000e-11'
+ mcm2d_cc_w_1_120_s_0_140 = '-8.75000e-13*ic_cap*ic_cap+-5.00000e-13*ic_cap+1.32000e-10'
+ mcm2d_cc_w_1_120_s_0_175 = '-7.81250e-13*ic_cap*ic_cap+-3.75000e-13*ic_cap+1.28000e-10'
+ mcm2d_cc_w_1_120_s_0_210 = '-6.87500e-13*ic_cap*ic_cap+-2.50000e-13*ic_cap+1.22000e-10'
+ mcm2d_cc_w_1_120_s_0_280 = '-5.21875e-13*ic_cap*ic_cap+-3.37500e-13*ic_cap+1.08000e-10'
+ mcm2d_cc_w_1_120_s_0_350 = '-3.78125e-13*ic_cap*ic_cap+-2.37500e-13*ic_cap+9.54000e-11'
+ mcm2d_cc_w_1_120_s_0_420 = '-2.90625e-13*ic_cap*ic_cap+-2.37500e-13*ic_cap+8.50000e-11'
+ mcm2d_cc_w_1_120_s_0_560 = '-1.50000e-13*ic_cap*ic_cap+-1.00000e-13*ic_cap+7.00000e-11'
+ mcm2d_cc_w_1_120_s_0_840 = '-4.68750e-14*ic_cap*ic_cap+-3.75000e-14*ic_cap+5.33000e-11'
+ mcm2d_cc_w_1_120_s_1_540 = '3.12500e-14*ic_cap*ic_cap+2.50000e-14*ic_cap+3.45000e-11'
+ mcm2d_cc_w_1_120_s_3_500 = '6.25000e-14*ic_cap*ic_cap+5.00000e-14*ic_cap+1.63000e-11'
+ mcm2d_cf_w_0_140_s_0_140 = '-1.25000e-15*ic_cap*ic_cap+-2.50000e-15*ic_cap+1.45000e-12'
+ mcm2d_cf_w_0_140_s_0_175 = '-5.00000e-15*ic_cap*ic_cap+-5.00000e-15*ic_cap+1.81000e-12'
+ mcm2d_cf_w_0_140_s_0_210 = '-9.06250e-15*ic_cap*ic_cap+-6.25000e-15*ic_cap+2.18000e-12'
+ mcm2d_cf_w_0_140_s_0_280 = '-1.62500e-14*ic_cap*ic_cap+-1.00000e-14*ic_cap+2.89000e-12'
+ mcm2d_cf_w_0_140_s_0_350 = '-2.37500e-14*ic_cap*ic_cap+-1.50000e-14*ic_cap+3.59000e-12'
+ mcm2d_cf_w_0_140_s_0_420 = '-3.09375e-14*ic_cap*ic_cap+-2.12500e-14*ic_cap+4.32000e-12'
+ mcm2d_cf_w_0_140_s_0_560 = '-4.34375e-14*ic_cap*ic_cap+-3.12500e-14*ic_cap+5.62000e-12'
+ mcm2d_cf_w_0_140_s_0_840 = '-7.00000e-14*ic_cap*ic_cap+-4.50000e-14*ic_cap+8.21000e-12'
+ mcm2d_cf_w_0_140_s_1_540 = '-1.12500e-13*ic_cap*ic_cap+-7.50000e-14*ic_cap+1.37000e-11'
+ mcm2d_cf_w_0_140_s_3_500 = '-1.71875e-13*ic_cap*ic_cap+-1.12500e-13*ic_cap+2.35000e-11'
+ mcm2d_cf_w_1_120_s_0_140 = '-2.18750e-15*ic_cap*ic_cap+-1.25000e-15*ic_cap+1.49000e-12'
+ mcm2d_cf_w_1_120_s_0_175 = '-5.62500e-15*ic_cap*ic_cap+-5.00000e-15*ic_cap+1.85000e-12'
+ mcm2d_cf_w_1_120_s_0_210 = '-9.37500e-15*ic_cap*ic_cap+-7.50000e-15*ic_cap+2.21000e-12'
+ mcm2d_cf_w_1_120_s_0_280 = '-1.65625e-14*ic_cap*ic_cap+-1.12500e-14*ic_cap+2.92000e-12'
+ mcm2d_cf_w_1_120_s_0_350 = '-2.40625e-14*ic_cap*ic_cap+-1.62500e-14*ic_cap+3.63000e-12'
+ mcm2d_cf_w_1_120_s_0_420 = '-3.06250e-14*ic_cap*ic_cap+-2.00000e-14*ic_cap+4.32000e-12'
+ mcm2d_cf_w_1_120_s_0_560 = '-4.43750e-14*ic_cap*ic_cap+-3.00000e-14*ic_cap+5.68000e-12'
+ mcm2d_cf_w_1_120_s_0_840 = '-6.93750e-14*ic_cap*ic_cap+-4.50000e-14*ic_cap+8.27000e-12'
+ mcm2d_cf_w_1_120_s_1_540 = '-1.18750e-13*ic_cap*ic_cap+-7.50000e-14*ic_cap+1.40000e-11'
+ mcm2d_cf_w_1_120_s_3_500 = '-1.84375e-13*ic_cap*ic_cap+-1.12500e-13*ic_cap+2.50000e-11'
+ mcm2f_ca_w_0_140_s_0_140 = '-1.90625e-07*ic_cap*ic_cap+-1.12500e-07*ic_cap+1.75000e-05'
+ mcm2f_ca_w_0_140_s_0_175 = '-1.90625e-07*ic_cap*ic_cap+-1.12500e-07*ic_cap+1.75000e-05'
+ mcm2f_ca_w_0_140_s_0_210 = '-1.90625e-07*ic_cap*ic_cap+-1.12500e-07*ic_cap+1.75000e-05'
+ mcm2f_ca_w_0_140_s_0_280 = '-1.90625e-07*ic_cap*ic_cap+-1.12500e-07*ic_cap+1.75000e-05'
+ mcm2f_ca_w_0_140_s_0_350 = '-1.90625e-07*ic_cap*ic_cap+-1.12500e-07*ic_cap+1.75000e-05'
+ mcm2f_ca_w_0_140_s_0_420 = '-1.90625e-07*ic_cap*ic_cap+-1.12500e-07*ic_cap+1.75000e-05'
+ mcm2f_ca_w_0_140_s_0_560 = '-1.90625e-07*ic_cap*ic_cap+-1.12500e-07*ic_cap+1.75000e-05'
+ mcm2f_ca_w_0_140_s_0_840 = '-1.90625e-07*ic_cap*ic_cap+-1.12500e-07*ic_cap+1.75000e-05'
+ mcm2f_ca_w_0_140_s_1_540 = '-1.90625e-07*ic_cap*ic_cap+-1.12500e-07*ic_cap+1.75000e-05'
+ mcm2f_ca_w_0_140_s_3_500 = '-1.90625e-07*ic_cap*ic_cap+-1.12500e-07*ic_cap+1.75000e-05'
+ mcm2f_ca_w_1_120_s_0_140 = '-1.90625e-07*ic_cap*ic_cap+-1.12500e-07*ic_cap+1.75000e-05'
+ mcm2f_ca_w_1_120_s_0_175 = '-1.90625e-07*ic_cap*ic_cap+-1.12500e-07*ic_cap+1.75000e-05'
+ mcm2f_ca_w_1_120_s_0_210 = '-1.90625e-07*ic_cap*ic_cap+-1.12500e-07*ic_cap+1.75000e-05'
+ mcm2f_ca_w_1_120_s_0_280 = '-1.90625e-07*ic_cap*ic_cap+-1.12500e-07*ic_cap+1.75000e-05'
+ mcm2f_ca_w_1_120_s_0_350 = '-1.90625e-07*ic_cap*ic_cap+-1.12500e-07*ic_cap+1.75000e-05'
+ mcm2f_ca_w_1_120_s_0_420 = '-1.90625e-07*ic_cap*ic_cap+-1.12500e-07*ic_cap+1.75000e-05'
+ mcm2f_ca_w_1_120_s_0_560 = '-1.90625e-07*ic_cap*ic_cap+-1.12500e-07*ic_cap+1.75000e-05'
+ mcm2f_ca_w_1_120_s_0_840 = '-1.90625e-07*ic_cap*ic_cap+-1.12500e-07*ic_cap+1.75000e-05'
+ mcm2f_ca_w_1_120_s_1_540 = '-1.90625e-07*ic_cap*ic_cap+-1.12500e-07*ic_cap+1.75000e-05'
+ mcm2f_ca_w_1_120_s_3_500 = '-1.90625e-07*ic_cap*ic_cap+-1.12500e-07*ic_cap+1.75000e-05'
+ mcm2f_cc_w_0_140_s_0_140 = '-1.02188e-12*ic_cap*ic_cap+-5.12500e-13*ic_cap+1.07000e-10'
+ mcm2f_cc_w_0_140_s_0_175 = '-9.03125e-13*ic_cap*ic_cap+-5.37500e-13*ic_cap+1.04000e-10'
+ mcm2f_cc_w_0_140_s_0_210 = '-7.68750e-13*ic_cap*ic_cap+-4.50000e-13*ic_cap+9.87000e-11'
+ mcm2f_cc_w_0_140_s_0_280 = '-6.21875e-13*ic_cap*ic_cap+-4.37500e-13*ic_cap+8.88000e-11'
+ mcm2f_cc_w_0_140_s_0_350 = '-4.81250e-13*ic_cap*ic_cap+-3.25000e-13*ic_cap+7.76000e-11'
+ mcm2f_cc_w_0_140_s_0_420 = '-3.84375e-13*ic_cap*ic_cap+-2.62500e-13*ic_cap+6.85000e-11'
+ mcm2f_cc_w_0_140_s_0_560 = '-2.37500e-13*ic_cap*ic_cap+-1.50000e-13*ic_cap+5.62000e-11'
+ mcm2f_cc_w_0_140_s_0_840 = '-1.03125e-13*ic_cap*ic_cap+-8.75000e-14*ic_cap+4.26000e-11'
+ mcm2f_cc_w_0_140_s_1_540 = '-6.25000e-15*ic_cap*ic_cap+2.74000e-11'
+ mcm2f_cc_w_0_140_s_3_500 = '4.68750e-14*ic_cap*ic_cap+3.75000e-14*ic_cap+1.27000e-11'
+ mcm2f_cc_w_1_120_s_0_140 = '-8.43750e-13*ic_cap*ic_cap+-3.75000e-13*ic_cap+1.33000e-10'
+ mcm2f_cc_w_1_120_s_0_175 = '-7.81250e-13*ic_cap*ic_cap+-3.75000e-13*ic_cap+1.29000e-10'
+ mcm2f_cc_w_1_120_s_0_210 = '-6.56250e-13*ic_cap*ic_cap+-3.75000e-13*ic_cap+1.23000e-10'
+ mcm2f_cc_w_1_120_s_0_280 = '-5.40625e-13*ic_cap*ic_cap+-4.12500e-13*ic_cap+1.10000e-10'
+ mcm2f_cc_w_1_120_s_0_350 = '-3.87500e-13*ic_cap*ic_cap+-2.50000e-13*ic_cap+9.70000e-11'
+ mcm2f_cc_w_1_120_s_0_420 = '-2.87500e-13*ic_cap*ic_cap+-2.50000e-13*ic_cap+8.65000e-11'
+ mcm2f_cc_w_1_120_s_0_560 = '-1.56250e-13*ic_cap*ic_cap+-1.00000e-13*ic_cap+7.16000e-11'
+ mcm2f_cc_w_1_120_s_0_840 = '-4.68750e-14*ic_cap*ic_cap+-3.75000e-14*ic_cap+5.50000e-11'
+ mcm2f_cc_w_1_120_s_1_540 = '3.12500e-14*ic_cap*ic_cap+2.50000e-14*ic_cap+3.62000e-11'
+ mcm2f_cc_w_1_120_s_3_500 = '7.50000e-14*ic_cap*ic_cap+5.00000e-14*ic_cap+1.79000e-11'
+ mcm2f_cf_w_0_140_s_0_140 = '-1.56250e-15*ic_cap*ic_cap+-1.25000e-15*ic_cap+1.22000e-12'
+ mcm2f_cf_w_0_140_s_0_175 = '-5.31250e-15*ic_cap*ic_cap+-3.75000e-15*ic_cap+1.53000e-12'
+ mcm2f_cf_w_0_140_s_0_210 = '-8.75000e-15*ic_cap*ic_cap+-5.00000e-15*ic_cap+1.84000e-12'
+ mcm2f_cf_w_0_140_s_0_280 = '-1.50000e-14*ic_cap*ic_cap+-1.00000e-14*ic_cap+2.44000e-12'
+ mcm2f_cf_w_0_140_s_0_350 = '-2.15625e-14*ic_cap*ic_cap+-1.37500e-14*ic_cap+3.03000e-12'
+ mcm2f_cf_w_0_140_s_0_420 = '-2.78125e-14*ic_cap*ic_cap+-1.87500e-14*ic_cap+3.65000e-12'
+ mcm2f_cf_w_0_140_s_0_560 = '-4.03125e-14*ic_cap*ic_cap+-2.62500e-14*ic_cap+4.77000e-12'
+ mcm2f_cf_w_0_140_s_0_840 = '-6.37500e-14*ic_cap*ic_cap+-4.00000e-14*ic_cap+6.98000e-12'
+ mcm2f_cf_w_0_140_s_1_540 = '-1.11563e-13*ic_cap*ic_cap+-7.12500e-14*ic_cap+1.19000e-11'
+ mcm2f_cf_w_0_140_s_3_500 = '-1.71875e-13*ic_cap*ic_cap+-1.12500e-13*ic_cap+2.10000e-11'
+ mcm2f_cf_w_1_120_s_0_140 = '-2.50000e-15*ic_cap*ic_cap+-2.50000e-15*ic_cap+1.25000e-12'
+ mcm2f_cf_w_1_120_s_0_175 = '-5.31250e-15*ic_cap*ic_cap+-3.75000e-15*ic_cap+1.55000e-12'
+ mcm2f_cf_w_1_120_s_0_210 = '-9.06250e-15*ic_cap*ic_cap+-6.25000e-15*ic_cap+1.86000e-12'
+ mcm2f_cf_w_1_120_s_0_280 = '-1.59375e-14*ic_cap*ic_cap+-1.12500e-14*ic_cap+2.47000e-12'
+ mcm2f_cf_w_1_120_s_0_350 = '-2.18750e-14*ic_cap*ic_cap+-1.50000e-14*ic_cap+3.06000e-12'
+ mcm2f_cf_w_1_120_s_0_420 = '-2.90625e-14*ic_cap*ic_cap+-1.87500e-14*ic_cap+3.66000e-12'
+ mcm2f_cf_w_1_120_s_0_560 = '-4.06250e-14*ic_cap*ic_cap+-2.75000e-14*ic_cap+4.81000e-12'
+ mcm2f_cf_w_1_120_s_0_840 = '-6.50000e-14*ic_cap*ic_cap+-4.00000e-14*ic_cap+7.06000e-12'
+ mcm2f_cf_w_1_120_s_1_540 = '-1.12813e-13*ic_cap*ic_cap+-7.62500e-14*ic_cap+1.21000e-11'
+ mcm2f_cf_w_1_120_s_3_500 = '-1.78125e-13*ic_cap*ic_cap+-1.12500e-13*ic_cap+2.22000e-11'
+ mcm2l1_ca_w_0_140_s_0_140 = '-4.50000e-07*ic_cap*ic_cap+-3.00000e-07*ic_cap+3.70000e-05'
+ mcm2l1_ca_w_0_140_s_0_175 = '-4.50000e-07*ic_cap*ic_cap+-3.00000e-07*ic_cap+3.70000e-05'
+ mcm2l1_ca_w_0_140_s_0_210 = '-4.50000e-07*ic_cap*ic_cap+-3.00000e-07*ic_cap+3.70000e-05'
+ mcm2l1_ca_w_0_140_s_0_280 = '-4.50000e-07*ic_cap*ic_cap+-3.00000e-07*ic_cap+3.70000e-05'
+ mcm2l1_ca_w_0_140_s_0_350 = '-4.50000e-07*ic_cap*ic_cap+-3.00000e-07*ic_cap+3.70000e-05'
+ mcm2l1_ca_w_0_140_s_0_420 = '-4.50000e-07*ic_cap*ic_cap+-3.00000e-07*ic_cap+3.70000e-05'
+ mcm2l1_ca_w_0_140_s_0_560 = '-4.50000e-07*ic_cap*ic_cap+-3.00000e-07*ic_cap+3.70000e-05'
+ mcm2l1_ca_w_0_140_s_0_840 = '-4.50000e-07*ic_cap*ic_cap+-3.00000e-07*ic_cap+3.70000e-05'
+ mcm2l1_ca_w_0_140_s_1_540 = '-4.50000e-07*ic_cap*ic_cap+-3.00000e-07*ic_cap+3.70000e-05'
+ mcm2l1_ca_w_0_140_s_3_500 = '-4.50000e-07*ic_cap*ic_cap+-3.00000e-07*ic_cap+3.70000e-05'
+ mcm2l1_ca_w_1_120_s_0_140 = '-4.50000e-07*ic_cap*ic_cap+-3.00000e-07*ic_cap+3.70000e-05'
+ mcm2l1_ca_w_1_120_s_0_175 = '-4.50000e-07*ic_cap*ic_cap+-3.00000e-07*ic_cap+3.70000e-05'
+ mcm2l1_ca_w_1_120_s_0_210 = '-4.50000e-07*ic_cap*ic_cap+-3.00000e-07*ic_cap+3.70000e-05'
+ mcm2l1_ca_w_1_120_s_0_280 = '-4.50000e-07*ic_cap*ic_cap+-3.00000e-07*ic_cap+3.70000e-05'
+ mcm2l1_ca_w_1_120_s_0_350 = '-4.50000e-07*ic_cap*ic_cap+-3.00000e-07*ic_cap+3.70000e-05'
+ mcm2l1_ca_w_1_120_s_0_420 = '-4.50000e-07*ic_cap*ic_cap+-3.00000e-07*ic_cap+3.70000e-05'
+ mcm2l1_ca_w_1_120_s_0_560 = '-4.50000e-07*ic_cap*ic_cap+-3.00000e-07*ic_cap+3.70000e-05'
+ mcm2l1_ca_w_1_120_s_0_840 = '-4.50000e-07*ic_cap*ic_cap+-3.00000e-07*ic_cap+3.70000e-05'
+ mcm2l1_ca_w_1_120_s_1_540 = '-4.50000e-07*ic_cap*ic_cap+-3.00000e-07*ic_cap+3.70000e-05'
+ mcm2l1_ca_w_1_120_s_3_500 = '-4.50000e-07*ic_cap*ic_cap+-3.00000e-07*ic_cap+3.70000e-05'
+ mcm2l1_cc_w_0_140_s_0_140 = '-8.81250e-13*ic_cap*ic_cap+-5.25000e-13*ic_cap+1.03000e-10'
+ mcm2l1_cc_w_0_140_s_0_175 = '-8.87500e-13*ic_cap*ic_cap+-5.25000e-13*ic_cap+1.02000e-10'
+ mcm2l1_cc_w_0_140_s_0_210 = '-7.31250e-13*ic_cap*ic_cap+-4.50000e-13*ic_cap+9.62000e-11'
+ mcm2l1_cc_w_0_140_s_0_280 = '-5.71875e-13*ic_cap*ic_cap+-3.37500e-13*ic_cap+8.51000e-11'
+ mcm2l1_cc_w_0_140_s_0_350 = '-4.28125e-13*ic_cap*ic_cap+-3.12500e-13*ic_cap+7.38000e-11'
+ mcm2l1_cc_w_0_140_s_0_420 = '-3.18750e-13*ic_cap*ic_cap+-2.00000e-13*ic_cap+6.44000e-11'
+ mcm2l1_cc_w_0_140_s_0_560 = '-1.78125e-13*ic_cap*ic_cap+-1.12500e-13*ic_cap+5.15000e-11'
+ mcm2l1_cc_w_0_140_s_0_840 = '-5.62500e-14*ic_cap*ic_cap+-5.00000e-14*ic_cap+3.71000e-11'
+ mcm2l1_cc_w_0_140_s_1_540 = '2.50000e-14*ic_cap*ic_cap+2.50000e-14*ic_cap+2.11000e-11'
+ mcm2l1_cc_w_0_140_s_3_500 = '4.50000e-14*ic_cap*ic_cap+3.75000e-14*ic_cap+7.54000e-12'
+ mcm2l1_cc_w_1_120_s_0_140 = '-8.43750e-13*ic_cap*ic_cap+-3.75000e-13*ic_cap+1.27000e-10'
+ mcm2l1_cc_w_1_120_s_0_175 = '-6.87500e-13*ic_cap*ic_cap+-5.00000e-13*ic_cap+1.22000e-10'
+ mcm2l1_cc_w_1_120_s_0_210 = '-6.25000e-13*ic_cap*ic_cap+-2.50000e-13*ic_cap+1.16000e-10'
+ mcm2l1_cc_w_1_120_s_0_280 = '-4.37500e-13*ic_cap*ic_cap+-2.50000e-13*ic_cap+1.02000e-10'
+ mcm2l1_cc_w_1_120_s_0_350 = '-3.25000e-13*ic_cap*ic_cap+-2.25000e-13*ic_cap+8.96000e-11'
+ mcm2l1_cc_w_1_120_s_0_420 = '-2.40625e-13*ic_cap*ic_cap+-1.37500e-13*ic_cap+7.92000e-11'
+ mcm2l1_cc_w_1_120_s_0_560 = '-1.09375e-13*ic_cap*ic_cap+-6.25000e-14*ic_cap+6.41000e-11'
+ mcm2l1_cc_w_1_120_s_0_840 = '-6.25000e-15*ic_cap*ic_cap+4.73000e-11'
+ mcm2l1_cc_w_1_120_s_1_540 = '5.31250e-14*ic_cap*ic_cap+3.75000e-14*ic_cap+2.86000e-11'
+ mcm2l1_cc_w_1_120_s_3_500 = '6.25000e-14*ic_cap*ic_cap+5.00000e-14*ic_cap+1.18000e-11'
+ mcm2l1_cf_w_0_140_s_0_140 = '-7.18750e-15*ic_cap*ic_cap+-6.25000e-15*ic_cap+2.54000e-12'
+ mcm2l1_cf_w_0_140_s_0_175 = '-1.50000e-14*ic_cap*ic_cap+-1.00000e-14*ic_cap+3.18000e-12'
+ mcm2l1_cf_w_0_140_s_0_210 = '-2.31250e-14*ic_cap*ic_cap+-1.75000e-14*ic_cap+3.83000e-12'
+ mcm2l1_cf_w_0_140_s_0_280 = '-3.78125e-14*ic_cap*ic_cap+-2.62500e-14*ic_cap+5.07000e-12'
+ mcm2l1_cf_w_0_140_s_0_350 = '-5.21875e-14*ic_cap*ic_cap+-3.87500e-14*ic_cap+6.28000e-12'
+ mcm2l1_cf_w_0_140_s_0_420 = '-6.71875e-14*ic_cap*ic_cap+-4.62500e-14*ic_cap+7.51000e-12'
+ mcm2l1_cf_w_0_140_s_0_560 = '-9.25000e-14*ic_cap*ic_cap+-6.50000e-14*ic_cap+9.75000e-12'
+ mcm2l1_cf_w_0_140_s_0_840 = '-1.34375e-13*ic_cap*ic_cap+-8.75000e-14*ic_cap+1.38000e-11'
+ mcm2l1_cf_w_0_140_s_1_540 = '-2.09375e-13*ic_cap*ic_cap+-1.37500e-13*ic_cap+2.20000e-11'
+ mcm2l1_cf_w_0_140_s_3_500 = '-2.50000e-13*ic_cap*ic_cap+-1.75000e-13*ic_cap+3.29000e-11'
+ mcm2l1_cf_w_1_120_s_0_140 = '-7.50000e-15*ic_cap*ic_cap+-7.50000e-15*ic_cap+2.57000e-12'
+ mcm2l1_cf_w_1_120_s_0_175 = '-1.50000e-14*ic_cap*ic_cap+-1.25000e-14*ic_cap+3.21000e-12'
+ mcm2l1_cf_w_1_120_s_0_210 = '-2.31250e-14*ic_cap*ic_cap+-1.75000e-14*ic_cap+3.85000e-12'
+ mcm2l1_cf_w_1_120_s_0_280 = '-3.81250e-14*ic_cap*ic_cap+-2.75000e-14*ic_cap+5.10000e-12'
+ mcm2l1_cf_w_1_120_s_0_350 = '-5.21875e-14*ic_cap*ic_cap+-3.62500e-14*ic_cap+6.32000e-12'
+ mcm2l1_cf_w_1_120_s_0_420 = '-6.71875e-14*ic_cap*ic_cap+-4.62500e-14*ic_cap+7.52000e-12'
+ mcm2l1_cf_w_1_120_s_0_560 = '-9.21875e-14*ic_cap*ic_cap+-6.12500e-14*ic_cap+9.79000e-12'
+ mcm2l1_cf_w_1_120_s_0_840 = '-1.37500e-13*ic_cap*ic_cap+-1.00000e-13*ic_cap+1.40000e-11'
+ mcm2l1_cf_w_1_120_s_1_540 = '-2.12500e-13*ic_cap*ic_cap+-1.50000e-13*ic_cap+2.25000e-11'
+ mcm2l1_cf_w_1_120_s_3_500 = '-2.62500e-13*ic_cap*ic_cap+-1.75000e-13*ic_cap+3.52000e-11'
+ mcm2l1d_ca_w_0_170_s_0_180 = '-1.00000e-06*ic_cap*ic_cap+-6.00000e-07*ic_cap+9.23000e-05'
+ mcm2l1d_ca_w_0_170_s_0_225 = '-1.00000e-06*ic_cap*ic_cap+-6.00000e-07*ic_cap+9.23000e-05'
+ mcm2l1d_ca_w_0_170_s_0_270 = '-1.00000e-06*ic_cap*ic_cap+-6.00000e-07*ic_cap+9.23000e-05'
+ mcm2l1d_ca_w_0_170_s_0_360 = '-1.00000e-06*ic_cap*ic_cap+-6.00000e-07*ic_cap+9.23000e-05'
+ mcm2l1d_ca_w_0_170_s_0_450 = '-1.00000e-06*ic_cap*ic_cap+-6.00000e-07*ic_cap+9.23000e-05'
+ mcm2l1d_ca_w_0_170_s_0_540 = '-1.00000e-06*ic_cap*ic_cap+-6.00000e-07*ic_cap+9.23000e-05'
+ mcm2l1d_ca_w_0_170_s_0_720 = '-1.00000e-06*ic_cap*ic_cap+-6.00000e-07*ic_cap+9.23000e-05'
+ mcm2l1d_ca_w_0_170_s_1_080 = '-1.00000e-06*ic_cap*ic_cap+-6.00000e-07*ic_cap+9.23000e-05'
+ mcm2l1d_ca_w_0_170_s_1_980 = '-1.00000e-06*ic_cap*ic_cap+-6.00000e-07*ic_cap+9.23000e-05'
+ mcm2l1d_ca_w_0_170_s_4_500 = '-1.00000e-06*ic_cap*ic_cap+-6.00000e-07*ic_cap+9.23000e-05'
+ mcm2l1d_ca_w_1_360_s_0_180 = '-1.00000e-06*ic_cap*ic_cap+-6.00000e-07*ic_cap+9.23000e-05'
+ mcm2l1d_ca_w_1_360_s_0_225 = '-1.00000e-06*ic_cap*ic_cap+-6.00000e-07*ic_cap+9.23000e-05'
+ mcm2l1d_ca_w_1_360_s_0_270 = '-1.00000e-06*ic_cap*ic_cap+-6.00000e-07*ic_cap+9.23000e-05'
+ mcm2l1d_ca_w_1_360_s_0_360 = '-1.00000e-06*ic_cap*ic_cap+-6.00000e-07*ic_cap+9.23000e-05'
+ mcm2l1d_ca_w_1_360_s_0_450 = '-1.00000e-06*ic_cap*ic_cap+-6.00000e-07*ic_cap+9.23000e-05'
+ mcm2l1d_ca_w_1_360_s_0_540 = '-1.00000e-06*ic_cap*ic_cap+-6.00000e-07*ic_cap+9.23000e-05'
+ mcm2l1d_ca_w_1_360_s_0_720 = '-1.00000e-06*ic_cap*ic_cap+-6.00000e-07*ic_cap+9.23000e-05'
+ mcm2l1d_ca_w_1_360_s_1_080 = '-1.00000e-06*ic_cap*ic_cap+-6.00000e-07*ic_cap+9.23000e-05'
+ mcm2l1d_ca_w_1_360_s_1_980 = '-1.00000e-06*ic_cap*ic_cap+-6.00000e-07*ic_cap+9.23000e-05'
+ mcm2l1d_ca_w_1_360_s_4_500 = '-1.00000e-06*ic_cap*ic_cap+-6.00000e-07*ic_cap+9.23000e-05'
+ mcm2l1d_cc_w_0_170_s_0_180 = '-7.21875e-13*ic_cap*ic_cap+-4.62500e-13*ic_cap+7.24000e-11'
+ mcm2l1d_cc_w_0_170_s_0_225 = '-5.03125e-13*ic_cap*ic_cap+-3.37500e-13*ic_cap+6.02000e-11'
+ mcm2l1d_cc_w_0_170_s_0_270 = '-3.53125e-13*ic_cap*ic_cap+-2.62500e-13*ic_cap+5.14000e-11'
+ mcm2l1d_cc_w_0_170_s_0_360 = '-1.96875e-13*ic_cap*ic_cap+-1.62500e-13*ic_cap+3.94000e-11'
+ mcm2l1d_cc_w_0_170_s_0_450 = '-1.03125e-13*ic_cap*ic_cap+-8.75000e-14*ic_cap+3.15000e-11'
+ mcm2l1d_cc_w_0_170_s_0_540 = '-5.00000e-14*ic_cap*ic_cap+-5.00000e-14*ic_cap+2.56000e-11'
+ mcm2l1d_cc_w_0_170_s_0_720 = '1.25000e-14*ic_cap*ic_cap+1.76000e-11'
+ mcm2l1d_cc_w_0_170_s_1_080 = '5.93750e-14*ic_cap*ic_cap+2.75000e-14*ic_cap+8.77000e-12'
+ mcm2l1d_cc_w_0_170_s_1_980 = '4.12500e-14*ic_cap*ic_cap+2.50000e-14*ic_cap+1.71000e-12'
+ mcm2l1d_cc_w_0_170_s_4_500 = '2.50000e-15*ic_cap*ic_cap+2.50000e-15*ic_cap+4.50000e-14'
+ mcm2l1d_cc_w_1_360_s_0_180 = '-5.59375e-13*ic_cap*ic_cap+-3.37500e-13*ic_cap+7.96000e-11'
+ mcm2l1d_cc_w_1_360_s_0_225 = '-3.46875e-13*ic_cap*ic_cap+-2.37500e-13*ic_cap+6.65000e-11'
+ mcm2l1d_cc_w_1_360_s_0_270 = '-2.21875e-13*ic_cap*ic_cap+-1.62500e-13*ic_cap+5.70000e-11'
+ mcm2l1d_cc_w_1_360_s_0_360 = '-7.18750e-14*ic_cap*ic_cap+-6.25000e-14*ic_cap+4.39000e-11'
+ mcm2l1d_cc_w_1_360_s_0_450 = '6.25000e-15*ic_cap*ic_cap+3.51000e-11'
+ mcm2l1d_cc_w_1_360_s_0_540 = '5.00000e-14*ic_cap*ic_cap+2.50000e-14*ic_cap+2.87000e-11'
+ mcm2l1d_cc_w_1_360_s_0_720 = '9.68750e-14*ic_cap*ic_cap+6.25000e-14*ic_cap+1.98000e-11'
+ mcm2l1d_cc_w_1_360_s_1_080 = '1.06250e-13*ic_cap*ic_cap+7.50000e-14*ic_cap+1.01000e-11'
+ mcm2l1d_cc_w_1_360_s_1_980 = '6.31250e-14*ic_cap*ic_cap+4.50000e-14*ic_cap+1.97000e-12'
+ mcm2l1d_cc_w_1_360_s_4_500 = '1.87500e-15*ic_cap*ic_cap+6.25000e-15*ic_cap+9.50000e-14'
+ mcm2l1d_cf_w_0_170_s_0_180 = '-2.28125e-14*ic_cap*ic_cap+-1.37500e-14*ic_cap+8.03000e-12'
+ mcm2l1d_cf_w_0_170_s_0_225 = '-4.28125e-14*ic_cap*ic_cap+-2.87500e-14*ic_cap+9.90000e-12'
+ mcm2l1d_cf_w_0_170_s_0_270 = '-6.56250e-14*ic_cap*ic_cap+-3.75000e-14*ic_cap+1.17000e-11'
+ mcm2l1d_cf_w_0_170_s_0_360 = '-9.68750e-14*ic_cap*ic_cap+-6.25000e-14*ic_cap+1.52000e-11'
+ mcm2l1d_cf_w_0_170_s_0_450 = '-1.37500e-13*ic_cap*ic_cap+-7.50000e-14*ic_cap+1.83000e-11'
+ mcm2l1d_cf_w_0_170_s_0_540 = '-1.62500e-13*ic_cap*ic_cap+-1.00000e-13*ic_cap+2.11000e-11'
+ mcm2l1d_cf_w_0_170_s_0_720 = '-2.06250e-13*ic_cap*ic_cap+-1.25000e-13*ic_cap+2.58000e-11'
+ mcm2l1d_cf_w_0_170_s_1_080 = '-2.53125e-13*ic_cap*ic_cap+-1.62500e-13*ic_cap+3.23000e-11'
+ mcm2l1d_cf_w_0_170_s_1_980 = '-2.46875e-13*ic_cap*ic_cap+-1.62500e-13*ic_cap+3.85000e-11'
+ mcm2l1d_cf_w_0_170_s_4_500 = '-2.06250e-13*ic_cap*ic_cap+-1.50000e-13*ic_cap+4.01000e-11'
+ mcm2l1d_cf_w_1_360_s_0_180 = '-2.15625e-14*ic_cap*ic_cap+-1.37500e-14*ic_cap+7.99000e-12'
+ mcm2l1d_cf_w_1_360_s_0_225 = '-4.25000e-14*ic_cap*ic_cap+-2.75000e-14*ic_cap+9.88000e-12'
+ mcm2l1d_cf_w_1_360_s_0_270 = '-5.93750e-14*ic_cap*ic_cap+-3.75000e-14*ic_cap+1.17000e-11'
+ mcm2l1d_cf_w_1_360_s_0_360 = '-1.03125e-13*ic_cap*ic_cap+-6.25000e-14*ic_cap+1.52000e-11'
+ mcm2l1d_cf_w_1_360_s_0_450 = '-1.31250e-13*ic_cap*ic_cap+-7.50000e-14*ic_cap+1.84000e-11'
+ mcm2l1d_cf_w_1_360_s_0_540 = '-1.62500e-13*ic_cap*ic_cap+-1.00000e-13*ic_cap+2.13000e-11'
+ mcm2l1d_cf_w_1_360_s_0_720 = '-2.00000e-13*ic_cap*ic_cap+-1.25000e-13*ic_cap+2.63000e-11'
+ mcm2l1d_cf_w_1_360_s_1_080 = '-2.37500e-13*ic_cap*ic_cap+-1.50000e-13*ic_cap+3.33000e-11'
+ mcm2l1d_cf_w_1_360_s_1_980 = '-2.09375e-13*ic_cap*ic_cap+-1.37500e-13*ic_cap+4.04000e-11'
+ mcm2l1d_cf_w_1_360_s_4_500 = '-1.56250e-13*ic_cap*ic_cap+-1.00000e-13*ic_cap+4.23000e-11'
+ mcm2l1f_ca_w_0_170_s_0_180 = '-8.68750e-07*ic_cap*ic_cap+-5.25000e-07*ic_cap+7.40000e-05'
+ mcm2l1f_ca_w_0_170_s_0_225 = '-8.68750e-07*ic_cap*ic_cap+-5.25000e-07*ic_cap+7.40000e-05'
+ mcm2l1f_ca_w_0_170_s_0_270 = '-8.68750e-07*ic_cap*ic_cap+-5.25000e-07*ic_cap+7.40000e-05'
+ mcm2l1f_ca_w_0_170_s_0_360 = '-8.68750e-07*ic_cap*ic_cap+-5.25000e-07*ic_cap+7.40000e-05'
+ mcm2l1f_ca_w_0_170_s_0_450 = '-8.68750e-07*ic_cap*ic_cap+-5.25000e-07*ic_cap+7.40000e-05'
+ mcm2l1f_ca_w_0_170_s_0_540 = '-8.68750e-07*ic_cap*ic_cap+-5.25000e-07*ic_cap+7.40000e-05'
+ mcm2l1f_ca_w_0_170_s_0_720 = '-8.68750e-07*ic_cap*ic_cap+-5.25000e-07*ic_cap+7.40000e-05'
+ mcm2l1f_ca_w_0_170_s_1_080 = '-8.68750e-07*ic_cap*ic_cap+-5.25000e-07*ic_cap+7.40000e-05'
+ mcm2l1f_ca_w_0_170_s_1_980 = '-8.68750e-07*ic_cap*ic_cap+-5.25000e-07*ic_cap+7.40000e-05'
+ mcm2l1f_ca_w_0_170_s_4_500 = '-8.68750e-07*ic_cap*ic_cap+-5.25000e-07*ic_cap+7.40000e-05'
+ mcm2l1f_ca_w_1_360_s_0_180 = '-8.68750e-07*ic_cap*ic_cap+-5.25000e-07*ic_cap+7.40000e-05'
+ mcm2l1f_ca_w_1_360_s_0_225 = '-8.68750e-07*ic_cap*ic_cap+-5.25000e-07*ic_cap+7.40000e-05'
+ mcm2l1f_ca_w_1_360_s_0_270 = '-8.68750e-07*ic_cap*ic_cap+-5.25000e-07*ic_cap+7.40000e-05'
+ mcm2l1f_ca_w_1_360_s_0_360 = '-8.68750e-07*ic_cap*ic_cap+-5.25000e-07*ic_cap+7.40000e-05'
+ mcm2l1f_ca_w_1_360_s_0_450 = '-8.68750e-07*ic_cap*ic_cap+-5.25000e-07*ic_cap+7.40000e-05'
+ mcm2l1f_ca_w_1_360_s_0_540 = '-8.68750e-07*ic_cap*ic_cap+-5.25000e-07*ic_cap+7.40000e-05'
+ mcm2l1f_ca_w_1_360_s_0_720 = '-8.68750e-07*ic_cap*ic_cap+-5.25000e-07*ic_cap+7.40000e-05'
+ mcm2l1f_ca_w_1_360_s_1_080 = '-8.68750e-07*ic_cap*ic_cap+-5.25000e-07*ic_cap+7.40000e-05'
+ mcm2l1f_ca_w_1_360_s_1_980 = '-8.68750e-07*ic_cap*ic_cap+-5.25000e-07*ic_cap+7.40000e-05'
+ mcm2l1f_ca_w_1_360_s_4_500 = '-8.68750e-07*ic_cap*ic_cap+-5.25000e-07*ic_cap+7.40000e-05'
+ mcm2l1f_cc_w_0_170_s_0_180 = '-7.40625e-13*ic_cap*ic_cap+-4.87500e-13*ic_cap+7.49000e-11'
+ mcm2l1f_cc_w_0_170_s_0_225 = '-5.15625e-13*ic_cap*ic_cap+-3.62500e-13*ic_cap+6.27000e-11'
+ mcm2l1f_cc_w_0_170_s_0_270 = '-3.65625e-13*ic_cap*ic_cap+-2.62500e-13*ic_cap+5.41000e-11'
+ mcm2l1f_cc_w_0_170_s_0_360 = '-2.12500e-13*ic_cap*ic_cap+-1.50000e-13*ic_cap+4.24000e-11'
+ mcm2l1f_cc_w_0_170_s_0_450 = '-1.06250e-13*ic_cap*ic_cap+-1.00000e-13*ic_cap+3.45000e-11'
+ mcm2l1f_cc_w_0_170_s_0_540 = '-5.93750e-14*ic_cap*ic_cap+-6.25000e-14*ic_cap+2.87000e-11'
+ mcm2l1f_cc_w_0_170_s_0_720 = '1.56250e-14*ic_cap*ic_cap+-1.25000e-14*ic_cap+2.06000e-11'
+ mcm2l1f_cc_w_0_170_s_1_080 = '6.87500e-14*ic_cap*ic_cap+2.50000e-14*ic_cap+1.13000e-11'
+ mcm2l1f_cc_w_0_170_s_1_980 = '6.06250e-14*ic_cap*ic_cap+4.00000e-14*ic_cap+2.81000e-12'
+ mcm2l1f_cc_w_0_170_s_4_500 = '5.93750e-15*ic_cap*ic_cap+5.00000e-15*ic_cap+9.50000e-14'
+ mcm2l1f_cc_w_1_360_s_0_180 = '-5.53125e-13*ic_cap*ic_cap+-3.37500e-13*ic_cap+8.41000e-11'
+ mcm2l1f_cc_w_1_360_s_0_225 = '-3.37500e-13*ic_cap*ic_cap+-2.25000e-13*ic_cap+7.09000e-11'
+ mcm2l1f_cc_w_1_360_s_0_270 = '-2.06250e-13*ic_cap*ic_cap+-1.50000e-13*ic_cap+6.14000e-11'
+ mcm2l1f_cc_w_1_360_s_0_360 = '-6.25000e-14*ic_cap*ic_cap+-5.00000e-14*ic_cap+4.83000e-11'
+ mcm2l1f_cc_w_1_360_s_0_450 = '1.87500e-14*ic_cap*ic_cap+3.94000e-11'
+ mcm2l1f_cc_w_1_360_s_0_540 = '6.25000e-14*ic_cap*ic_cap+2.50000e-14*ic_cap+3.29000e-11'
+ mcm2l1f_cc_w_1_360_s_0_720 = '1.15625e-13*ic_cap*ic_cap+6.25000e-14*ic_cap+2.37000e-11'
+ mcm2l1f_cc_w_1_360_s_1_080 = '1.34375e-13*ic_cap*ic_cap+8.75000e-14*ic_cap+1.32000e-11'
+ mcm2l1f_cc_w_1_360_s_1_980 = '9.40625e-14*ic_cap*ic_cap+6.37500e-14*ic_cap+3.32000e-12'
+ mcm2l1f_cc_w_1_360_s_4_500 = '6.87500e-15*ic_cap*ic_cap+1.00000e-14*ic_cap+1.30000e-13'
+ mcm2l1f_cf_w_0_170_s_0_180 = '-2.40625e-14*ic_cap*ic_cap+-1.62500e-14*ic_cap+6.47000e-12'
+ mcm2l1f_cf_w_0_170_s_0_225 = '-4.34375e-14*ic_cap*ic_cap+-2.87500e-14*ic_cap+8.02000e-12'
+ mcm2l1f_cf_w_0_170_s_0_270 = '-6.09375e-14*ic_cap*ic_cap+-3.87500e-14*ic_cap+9.48000e-12'
+ mcm2l1f_cf_w_0_170_s_0_360 = '-9.06250e-14*ic_cap*ic_cap+-6.25000e-14*ic_cap+1.24000e-11'
+ mcm2l1f_cf_w_0_170_s_0_450 = '-1.25000e-13*ic_cap*ic_cap+-7.50000e-14*ic_cap+1.50000e-11'
+ mcm2l1f_cf_w_0_170_s_0_540 = '-1.53125e-13*ic_cap*ic_cap+-8.75000e-14*ic_cap+1.75000e-11'
+ mcm2l1f_cf_w_0_170_s_0_720 = '-1.93750e-13*ic_cap*ic_cap+-1.25000e-13*ic_cap+2.17000e-11'
+ mcm2l1f_cf_w_0_170_s_1_080 = '-2.43750e-13*ic_cap*ic_cap+-1.50000e-13*ic_cap+2.79000e-11'
+ mcm2l1f_cf_w_0_170_s_1_980 = '-2.50000e-13*ic_cap*ic_cap+-1.75000e-13*ic_cap+3.50000e-11'
+ mcm2l1f_cf_w_0_170_s_4_500 = '-2.03125e-13*ic_cap*ic_cap+-1.37500e-13*ic_cap+3.76000e-11'
+ mcm2l1f_cf_w_1_360_s_0_180 = '-2.34375e-14*ic_cap*ic_cap+-1.62500e-14*ic_cap+6.43000e-12'
+ mcm2l1f_cf_w_1_360_s_0_225 = '-4.15625e-14*ic_cap*ic_cap+-2.62500e-14*ic_cap+7.97000e-12'
+ mcm2l1f_cf_w_1_360_s_0_270 = '-5.93750e-14*ic_cap*ic_cap+-3.75000e-14*ic_cap+9.48000e-12'
+ mcm2l1f_cf_w_1_360_s_0_360 = '-9.37500e-14*ic_cap*ic_cap+-5.00000e-14*ic_cap+1.24000e-11'
+ mcm2l1f_cf_w_1_360_s_0_450 = '-1.25000e-13*ic_cap*ic_cap+-7.50000e-14*ic_cap+1.51000e-11'
+ mcm2l1f_cf_w_1_360_s_0_540 = '-1.46875e-13*ic_cap*ic_cap+-8.75000e-14*ic_cap+1.76000e-11'
+ mcm2l1f_cf_w_1_360_s_0_720 = '-1.93750e-13*ic_cap*ic_cap+-1.25000e-13*ic_cap+2.21000e-11'
+ mcm2l1f_cf_w_1_360_s_1_080 = '-2.34375e-13*ic_cap*ic_cap+-1.62500e-13*ic_cap+2.88000e-11'
+ mcm2l1f_cf_w_1_360_s_1_980 = '-2.25000e-13*ic_cap*ic_cap+-1.50000e-13*ic_cap+3.70000e-11'
+ mcm2l1f_cf_w_1_360_s_4_500 = '-1.50000e-13*ic_cap*ic_cap+-1.00000e-13*ic_cap+4.01000e-11'
+ mcm2l1p1_ca_w_0_170_s_0_180 = '-2.08750e-06*ic_cap*ic_cap+-1.10000e-06*ic_cap+1.31000e-04'
+ mcm2l1p1_ca_w_0_170_s_0_225 = '-2.08750e-06*ic_cap*ic_cap+-1.10000e-06*ic_cap+1.31000e-04'
+ mcm2l1p1_ca_w_0_170_s_0_270 = '-2.08750e-06*ic_cap*ic_cap+-1.10000e-06*ic_cap+1.31000e-04'
+ mcm2l1p1_ca_w_0_170_s_0_360 = '-2.08750e-06*ic_cap*ic_cap+-1.10000e-06*ic_cap+1.31000e-04'
+ mcm2l1p1_ca_w_0_170_s_0_450 = '-2.08750e-06*ic_cap*ic_cap+-1.10000e-06*ic_cap+1.31000e-04'
+ mcm2l1p1_ca_w_0_170_s_0_540 = '-2.08750e-06*ic_cap*ic_cap+-1.10000e-06*ic_cap+1.31000e-04'
+ mcm2l1p1_ca_w_0_170_s_0_720 = '-2.08750e-06*ic_cap*ic_cap+-1.10000e-06*ic_cap+1.31000e-04'
+ mcm2l1p1_ca_w_0_170_s_1_080 = '-2.08750e-06*ic_cap*ic_cap+-1.10000e-06*ic_cap+1.31000e-04'
+ mcm2l1p1_ca_w_0_170_s_1_980 = '-2.08750e-06*ic_cap*ic_cap+-1.10000e-06*ic_cap+1.31000e-04'
+ mcm2l1p1_ca_w_0_170_s_4_500 = '-2.08750e-06*ic_cap*ic_cap+-1.10000e-06*ic_cap+1.31000e-04'
+ mcm2l1p1_ca_w_1_360_s_0_180 = '-2.08750e-06*ic_cap*ic_cap+-1.10000e-06*ic_cap+1.31000e-04'
+ mcm2l1p1_ca_w_1_360_s_0_225 = '-2.08750e-06*ic_cap*ic_cap+-1.10000e-06*ic_cap+1.31000e-04'
+ mcm2l1p1_ca_w_1_360_s_0_270 = '-2.08750e-06*ic_cap*ic_cap+-1.10000e-06*ic_cap+1.31000e-04'
+ mcm2l1p1_ca_w_1_360_s_0_360 = '-2.08750e-06*ic_cap*ic_cap+-1.10000e-06*ic_cap+1.31000e-04'
+ mcm2l1p1_ca_w_1_360_s_0_450 = '-2.08750e-06*ic_cap*ic_cap+-1.10000e-06*ic_cap+1.31000e-04'
+ mcm2l1p1_ca_w_1_360_s_0_540 = '-2.08750e-06*ic_cap*ic_cap+-1.10000e-06*ic_cap+1.31000e-04'
+ mcm2l1p1_ca_w_1_360_s_0_720 = '-2.08750e-06*ic_cap*ic_cap+-1.10000e-06*ic_cap+1.31000e-04'
+ mcm2l1p1_ca_w_1_360_s_1_080 = '-2.08750e-06*ic_cap*ic_cap+-1.10000e-06*ic_cap+1.31000e-04'
+ mcm2l1p1_ca_w_1_360_s_1_980 = '-2.08750e-06*ic_cap*ic_cap+-1.10000e-06*ic_cap+1.31000e-04'
+ mcm2l1p1_ca_w_1_360_s_4_500 = '-2.08750e-06*ic_cap*ic_cap+-1.10000e-06*ic_cap+1.31000e-04'
+ mcm2l1p1_cc_w_0_170_s_0_180 = '-6.25000e-13*ic_cap*ic_cap+-4.00000e-13*ic_cap+6.82000e-11'
+ mcm2l1p1_cc_w_0_170_s_0_225 = '-3.84375e-13*ic_cap*ic_cap+-2.87500e-13*ic_cap+5.56000e-11'
+ mcm2l1p1_cc_w_0_170_s_0_270 = '-2.46875e-13*ic_cap*ic_cap+-2.12500e-13*ic_cap+4.68000e-11'
+ mcm2l1p1_cc_w_0_170_s_0_360 = '-8.75000e-14*ic_cap*ic_cap+-1.00000e-13*ic_cap+3.47000e-11'
+ mcm2l1p1_cc_w_0_170_s_0_450 = '-5.00000e-14*ic_cap+2.68000e-11'
+ mcm2l1p1_cc_w_0_170_s_0_540 = '5.00000e-14*ic_cap*ic_cap+2.10000e-11'
+ mcm2l1p1_cc_w_0_170_s_0_720 = '9.68750e-14*ic_cap*ic_cap+3.75000e-14*ic_cap+1.34000e-11'
+ mcm2l1p1_cc_w_0_170_s_1_080 = '1.03125e-13*ic_cap*ic_cap+5.50000e-14*ic_cap+5.79000e-12'
+ mcm2l1p1_cc_w_0_170_s_1_980 = '4.31250e-14*ic_cap*ic_cap+3.00000e-14*ic_cap+8.00000e-13'
+ mcm2l1p1_cc_w_0_170_s_4_500 = '2.50000e-15*ic_cap*ic_cap+1.25000e-15*ic_cap+5.00000e-15'
+ mcm2l1p1_cc_w_1_360_s_0_180 = '-4.56250e-13*ic_cap*ic_cap+-3.00000e-13*ic_cap+7.38000e-11'
+ mcm2l1p1_cc_w_1_360_s_0_225 = '-2.46875e-13*ic_cap*ic_cap+-1.87500e-13*ic_cap+6.07000e-11'
+ mcm2l1p1_cc_w_1_360_s_0_270 = '-1.18750e-13*ic_cap*ic_cap+-1.00000e-13*ic_cap+5.13000e-11'
+ mcm2l1p1_cc_w_1_360_s_0_360 = '2.81250e-14*ic_cap*ic_cap+-1.25000e-14*ic_cap+3.83000e-11'
+ mcm2l1p1_cc_w_1_360_s_0_450 = '9.68750e-14*ic_cap*ic_cap+3.75000e-14*ic_cap+2.97000e-11'
+ mcm2l1p1_cc_w_1_360_s_0_540 = '1.37500e-13*ic_cap*ic_cap+7.50000e-14*ic_cap+2.35000e-11'
+ mcm2l1p1_cc_w_1_360_s_0_720 = '1.65625e-13*ic_cap*ic_cap+8.75000e-14*ic_cap+1.52000e-11'
+ mcm2l1p1_cc_w_1_360_s_1_080 = '1.53125e-13*ic_cap*ic_cap+9.00000e-14*ic_cap+6.72000e-12'
+ mcm2l1p1_cc_w_1_360_s_1_980 = '5.59375e-14*ic_cap*ic_cap+4.25000e-14*ic_cap+9.95000e-13'
+ mcm2l1p1_cc_w_1_360_s_4_500 = '-1.40625e-15*ic_cap*ic_cap+-3.12500e-15*ic_cap+6.00000e-14'
+ mcm2l1p1_cf_w_0_170_s_0_180 = '-9.43750e-14*ic_cap*ic_cap+-4.75000e-14*ic_cap+1.12000e-11'
+ mcm2l1p1_cf_w_0_170_s_0_225 = '-1.37500e-13*ic_cap*ic_cap+-7.50000e-14*ic_cap+1.38000e-11'
+ mcm2l1p1_cf_w_0_170_s_0_270 = '-1.75000e-13*ic_cap*ic_cap+-1.00000e-13*ic_cap+1.62000e-11'
+ mcm2l1p1_cf_w_0_170_s_0_360 = '-2.40625e-13*ic_cap*ic_cap+-1.37500e-13*ic_cap+2.08000e-11'
+ mcm2l1p1_cf_w_0_170_s_0_450 = '-2.96875e-13*ic_cap*ic_cap+-1.62500e-13*ic_cap+2.46000e-11'
+ mcm2l1p1_cf_w_0_170_s_0_540 = '-3.37500e-13*ic_cap*ic_cap+-1.75000e-13*ic_cap+2.80000e-11'
+ mcm2l1p1_cf_w_0_170_s_0_720 = '-3.90625e-13*ic_cap*ic_cap+-2.12500e-13*ic_cap+3.33000e-11'
+ mcm2l1p1_cf_w_0_170_s_1_080 = '-4.15625e-13*ic_cap*ic_cap+-2.37500e-13*ic_cap+3.95000e-11'
+ mcm2l1p1_cf_w_0_170_s_1_980 = '-3.68750e-13*ic_cap*ic_cap+-2.25000e-13*ic_cap+4.41000e-11'
+ mcm2l1p1_cf_w_0_170_s_4_500 = '-3.31250e-13*ic_cap*ic_cap+-2.00000e-13*ic_cap+4.49000e-11'
+ mcm2l1p1_cf_w_1_360_s_0_180 = '-9.62500e-14*ic_cap*ic_cap+-4.75000e-14*ic_cap+1.12000e-11'
+ mcm2l1p1_cf_w_1_360_s_0_225 = '-1.31250e-13*ic_cap*ic_cap+-7.50000e-14*ic_cap+1.37000e-11'
+ mcm2l1p1_cf_w_1_360_s_0_270 = '-1.71875e-13*ic_cap*ic_cap+-8.75000e-14*ic_cap+1.62000e-11'
+ mcm2l1p1_cf_w_1_360_s_0_360 = '-2.37500e-13*ic_cap*ic_cap+-1.25000e-13*ic_cap+2.07000e-11'
+ mcm2l1p1_cf_w_1_360_s_0_450 = '-2.87500e-13*ic_cap*ic_cap+-1.50000e-13*ic_cap+2.47000e-11'
+ mcm2l1p1_cf_w_1_360_s_0_540 = '-3.28125e-13*ic_cap*ic_cap+-1.87500e-13*ic_cap+2.82000e-11'
+ mcm2l1p1_cf_w_1_360_s_0_720 = '-3.71875e-13*ic_cap*ic_cap+-2.12500e-13*ic_cap+3.37000e-11'
+ mcm2l1p1_cf_w_1_360_s_1_080 = '-3.96875e-13*ic_cap*ic_cap+-2.37500e-13*ic_cap+4.06000e-11'
+ mcm2l1p1_cf_w_1_360_s_1_980 = '-3.18750e-13*ic_cap*ic_cap+-2.00000e-13*ic_cap+4.59000e-11'
+ mcm2l1p1_cf_w_1_360_s_4_500 = '-2.68750e-13*ic_cap*ic_cap+-1.50000e-13*ic_cap+4.69000e-11'
+ mcm2m1_ca_w_0_140_s_0_140 = '-2.66250e-06*ic_cap*ic_cap+-1.25000e-06*ic_cap+1.28000e-04'
+ mcm2m1_ca_w_0_140_s_0_175 = '-2.66250e-06*ic_cap*ic_cap+-1.25000e-06*ic_cap+1.28000e-04'
+ mcm2m1_ca_w_0_140_s_0_210 = '-2.66250e-06*ic_cap*ic_cap+-1.25000e-06*ic_cap+1.28000e-04'
+ mcm2m1_ca_w_0_140_s_0_280 = '-2.66250e-06*ic_cap*ic_cap+-1.25000e-06*ic_cap+1.28000e-04'
+ mcm2m1_ca_w_0_140_s_0_350 = '-2.66250e-06*ic_cap*ic_cap+-1.25000e-06*ic_cap+1.28000e-04'
+ mcm2m1_ca_w_0_140_s_0_420 = '-2.66250e-06*ic_cap*ic_cap+-1.25000e-06*ic_cap+1.28000e-04'
+ mcm2m1_ca_w_0_140_s_0_560 = '-2.66250e-06*ic_cap*ic_cap+-1.25000e-06*ic_cap+1.28000e-04'
+ mcm2m1_ca_w_0_140_s_0_840 = '-2.66250e-06*ic_cap*ic_cap+-1.25000e-06*ic_cap+1.28000e-04'
+ mcm2m1_ca_w_0_140_s_1_540 = '-2.66250e-06*ic_cap*ic_cap+-1.25000e-06*ic_cap+1.28000e-04'
+ mcm2m1_ca_w_0_140_s_3_500 = '-2.66250e-06*ic_cap*ic_cap+-1.25000e-06*ic_cap+1.28000e-04'
+ mcm2m1_ca_w_1_120_s_0_140 = '-2.66250e-06*ic_cap*ic_cap+-1.25000e-06*ic_cap+1.28000e-04'
+ mcm2m1_ca_w_1_120_s_0_175 = '-2.66250e-06*ic_cap*ic_cap+-1.25000e-06*ic_cap+1.28000e-04'
+ mcm2m1_ca_w_1_120_s_0_210 = '-2.66250e-06*ic_cap*ic_cap+-1.25000e-06*ic_cap+1.28000e-04'
+ mcm2m1_ca_w_1_120_s_0_280 = '-2.66250e-06*ic_cap*ic_cap+-1.25000e-06*ic_cap+1.28000e-04'
+ mcm2m1_ca_w_1_120_s_0_350 = '-2.66250e-06*ic_cap*ic_cap+-1.25000e-06*ic_cap+1.28000e-04'
+ mcm2m1_ca_w_1_120_s_0_420 = '-2.66250e-06*ic_cap*ic_cap+-1.25000e-06*ic_cap+1.28000e-04'
+ mcm2m1_ca_w_1_120_s_0_560 = '-2.66250e-06*ic_cap*ic_cap+-1.25000e-06*ic_cap+1.28000e-04'
+ mcm2m1_ca_w_1_120_s_0_840 = '-2.66250e-06*ic_cap*ic_cap+-1.25000e-06*ic_cap+1.28000e-04'
+ mcm2m1_ca_w_1_120_s_1_540 = '-2.66250e-06*ic_cap*ic_cap+-1.25000e-06*ic_cap+1.28000e-04'
+ mcm2m1_ca_w_1_120_s_3_500 = '-2.66250e-06*ic_cap*ic_cap+-1.25000e-06*ic_cap+1.28000e-04'
+ mcm2m1_cc_w_0_140_s_0_140 = '-7.06250e-13*ic_cap*ic_cap+-4.75000e-13*ic_cap+9.46000e-11'
+ mcm2m1_cc_w_0_140_s_0_175 = '-6.71875e-13*ic_cap*ic_cap+-4.62500e-13*ic_cap+9.27000e-11'
+ mcm2m1_cc_w_0_140_s_0_210 = '-5.50000e-13*ic_cap*ic_cap+-3.25000e-13*ic_cap+8.69000e-11'
+ mcm2m1_cc_w_0_140_s_0_280 = '-3.78125e-13*ic_cap*ic_cap+-2.37500e-13*ic_cap+7.48000e-11'
+ mcm2m1_cc_w_0_140_s_0_350 = '-2.50000e-13*ic_cap*ic_cap+-2.25000e-13*ic_cap+6.32000e-11'
+ mcm2m1_cc_w_0_140_s_0_420 = '-1.40625e-13*ic_cap*ic_cap+-1.37500e-13*ic_cap+5.31000e-11'
+ mcm2m1_cc_w_0_140_s_0_560 = '-2.18750e-14*ic_cap*ic_cap+-6.25000e-14*ic_cap+4.01000e-11'
+ mcm2m1_cc_w_0_140_s_0_840 = '5.31250e-14*ic_cap*ic_cap+1.25000e-14*ic_cap+2.60000e-11'
+ mcm2m1_cc_w_0_140_s_1_540 = '6.87500e-14*ic_cap*ic_cap+5.00000e-14*ic_cap+1.19000e-11'
+ mcm2m1_cc_w_0_140_s_3_500 = '2.65625e-14*ic_cap*ic_cap+1.87500e-14*ic_cap+3.35000e-12'
+ mcm2m1_cc_w_1_120_s_0_140 = '-6.56250e-13*ic_cap*ic_cap+-3.75000e-13*ic_cap+1.13000e-10'
+ mcm2m1_cc_w_1_120_s_0_175 = '-5.90625e-13*ic_cap*ic_cap+-3.62500e-13*ic_cap+1.09000e-10'
+ mcm2m1_cc_w_1_120_s_0_210 = '-4.50000e-13*ic_cap*ic_cap+-3.25000e-13*ic_cap+1.02000e-10'
+ mcm2m1_cc_w_1_120_s_0_280 = '-3.46875e-13*ic_cap*ic_cap+-2.12500e-13*ic_cap+8.91000e-11'
+ mcm2m1_cc_w_1_120_s_0_350 = '-2.00000e-13*ic_cap*ic_cap+-1.75000e-13*ic_cap+7.62000e-11'
+ mcm2m1_cc_w_1_120_s_0_420 = '-1.18750e-13*ic_cap*ic_cap+-1.25000e-13*ic_cap+6.60000e-11'
+ mcm2m1_cc_w_1_120_s_0_560 = '-6.25000e-15*ic_cap*ic_cap+-2.50000e-14*ic_cap+5.15000e-11'
+ mcm2m1_cc_w_1_120_s_0_840 = '7.18750e-14*ic_cap*ic_cap+3.75000e-14*ic_cap+3.55000e-11'
+ mcm2m1_cc_w_1_120_s_1_540 = '8.12500e-14*ic_cap*ic_cap+5.00000e-14*ic_cap+1.90000e-11'
+ mcm2m1_cc_w_1_120_s_3_500 = '3.90625e-14*ic_cap*ic_cap+3.12500e-14*ic_cap+6.75000e-12'
+ mcm2m1_cf_w_0_140_s_0_140 = '-1.00938e-13*ic_cap*ic_cap+-5.12500e-14*ic_cap+8.24000e-12'
+ mcm2m1_cf_w_0_140_s_0_175 = '-1.43750e-13*ic_cap*ic_cap+-7.00000e-14*ic_cap+1.04000e-11'
+ mcm2m1_cf_w_0_140_s_0_210 = '-1.86250e-13*ic_cap*ic_cap+-9.00000e-14*ic_cap+1.25000e-11'
+ mcm2m1_cf_w_0_140_s_0_280 = '-2.68750e-13*ic_cap*ic_cap+-1.25000e-13*ic_cap+1.65000e-11'
+ mcm2m1_cf_w_0_140_s_0_350 = '-3.34375e-13*ic_cap*ic_cap+-1.62500e-13*ic_cap+2.01000e-11'
+ mcm2m1_cf_w_0_140_s_0_420 = '-3.87500e-13*ic_cap*ic_cap+-2.00000e-13*ic_cap+2.34000e-11'
+ mcm2m1_cf_w_0_140_s_0_560 = '-4.75000e-13*ic_cap*ic_cap+-2.50000e-13*ic_cap+2.91000e-11'
+ mcm2m1_cf_w_0_140_s_0_840 = '-5.81250e-13*ic_cap*ic_cap+-3.00000e-13*ic_cap+3.77000e-11'
+ mcm2m1_cf_w_0_140_s_1_540 = '-6.46875e-13*ic_cap*ic_cap+-3.37500e-13*ic_cap+4.94000e-11'
+ mcm2m1_cf_w_0_140_s_3_500 = '-6.31250e-13*ic_cap*ic_cap+-3.25000e-13*ic_cap+5.79000e-11'
+ mcm2m1_cf_w_1_120_s_0_140 = '-1.00625e-13*ic_cap*ic_cap+-4.75000e-14*ic_cap+8.25000e-12'
+ mcm2m1_cf_w_1_120_s_0_175 = '-1.48750e-13*ic_cap*ic_cap+-7.00000e-14*ic_cap+1.05000e-11'
+ mcm2m1_cf_w_1_120_s_0_210 = '-1.85000e-13*ic_cap*ic_cap+-9.00000e-14*ic_cap+1.25000e-11'
+ mcm2m1_cf_w_1_120_s_0_280 = '-2.68750e-13*ic_cap*ic_cap+-1.25000e-13*ic_cap+1.65000e-11'
+ mcm2m1_cf_w_1_120_s_0_350 = '-3.34375e-13*ic_cap*ic_cap+-1.62500e-13*ic_cap+2.01000e-11'
+ mcm2m1_cf_w_1_120_s_0_420 = '-3.90625e-13*ic_cap*ic_cap+-1.87500e-13*ic_cap+2.34000e-11'
+ mcm2m1_cf_w_1_120_s_0_560 = '-4.71875e-13*ic_cap*ic_cap+-2.37500e-13*ic_cap+2.91000e-11'
+ mcm2m1_cf_w_1_120_s_0_840 = '-5.75000e-13*ic_cap*ic_cap+-3.00000e-13*ic_cap+3.78000e-11'
+ mcm2m1_cf_w_1_120_s_1_540 = '-6.56250e-13*ic_cap*ic_cap+-3.50000e-13*ic_cap+5.05000e-11'
+ mcm2m1_cf_w_1_120_s_3_500 = '-6.56250e-13*ic_cap*ic_cap+-3.50000e-13*ic_cap+6.23000e-11'
+ mcm2m1d_ca_w_0_140_s_0_140 = '-3.06250e-06*ic_cap*ic_cap+-1.50000e-06*ic_cap+1.62000e-04'
+ mcm2m1d_ca_w_0_140_s_0_175 = '-3.06250e-06*ic_cap*ic_cap+-1.50000e-06*ic_cap+1.62000e-04'
+ mcm2m1d_ca_w_0_140_s_0_210 = '-3.06250e-06*ic_cap*ic_cap+-1.50000e-06*ic_cap+1.62000e-04'
+ mcm2m1d_ca_w_0_140_s_0_280 = '-3.06250e-06*ic_cap*ic_cap+-1.50000e-06*ic_cap+1.62000e-04'
+ mcm2m1d_ca_w_0_140_s_0_350 = '-3.06250e-06*ic_cap*ic_cap+-1.50000e-06*ic_cap+1.62000e-04'
+ mcm2m1d_ca_w_0_140_s_0_420 = '-3.06250e-06*ic_cap*ic_cap+-1.50000e-06*ic_cap+1.62000e-04'
+ mcm2m1d_ca_w_0_140_s_0_560 = '-3.06250e-06*ic_cap*ic_cap+-1.50000e-06*ic_cap+1.62000e-04'
+ mcm2m1d_ca_w_0_140_s_0_840 = '-3.06250e-06*ic_cap*ic_cap+-1.50000e-06*ic_cap+1.62000e-04'
+ mcm2m1d_ca_w_0_140_s_1_540 = '-3.06250e-06*ic_cap*ic_cap+-1.50000e-06*ic_cap+1.62000e-04'
+ mcm2m1d_ca_w_0_140_s_3_500 = '-3.06250e-06*ic_cap*ic_cap+-1.50000e-06*ic_cap+1.62000e-04'
+ mcm2m1d_ca_w_1_120_s_0_140 = '-3.06250e-06*ic_cap*ic_cap+-1.50000e-06*ic_cap+1.62000e-04'
+ mcm2m1d_ca_w_1_120_s_0_175 = '-3.06250e-06*ic_cap*ic_cap+-1.50000e-06*ic_cap+1.62000e-04'
+ mcm2m1d_ca_w_1_120_s_0_210 = '-3.06250e-06*ic_cap*ic_cap+-1.50000e-06*ic_cap+1.62000e-04'
+ mcm2m1d_ca_w_1_120_s_0_280 = '-3.06250e-06*ic_cap*ic_cap+-1.50000e-06*ic_cap+1.62000e-04'
+ mcm2m1d_ca_w_1_120_s_0_350 = '-3.06250e-06*ic_cap*ic_cap+-1.50000e-06*ic_cap+1.62000e-04'
+ mcm2m1d_ca_w_1_120_s_0_420 = '-3.06250e-06*ic_cap*ic_cap+-1.50000e-06*ic_cap+1.62000e-04'
+ mcm2m1d_ca_w_1_120_s_0_560 = '-3.06250e-06*ic_cap*ic_cap+-1.50000e-06*ic_cap+1.62000e-04'
+ mcm2m1d_ca_w_1_120_s_0_840 = '-3.06250e-06*ic_cap*ic_cap+-1.50000e-06*ic_cap+1.62000e-04'
+ mcm2m1d_ca_w_1_120_s_1_540 = '-3.06250e-06*ic_cap*ic_cap+-1.50000e-06*ic_cap+1.62000e-04'
+ mcm2m1d_ca_w_1_120_s_3_500 = '-3.06250e-06*ic_cap*ic_cap+-1.50000e-06*ic_cap+1.62000e-04'
+ mcm2m1d_cc_w_0_140_s_0_140 = '-6.71875e-13*ic_cap*ic_cap+-3.87500e-13*ic_cap+9.13000e-11'
+ mcm2m1d_cc_w_0_140_s_0_175 = '-6.62500e-13*ic_cap*ic_cap+-3.25000e-13*ic_cap+8.90000e-11'
+ mcm2m1d_cc_w_0_140_s_0_210 = '-5.37500e-13*ic_cap*ic_cap+-3.50000e-13*ic_cap+8.32000e-11'
+ mcm2m1d_cc_w_0_140_s_0_280 = '-3.12500e-13*ic_cap*ic_cap+-2.75000e-13*ic_cap+6.98000e-11'
+ mcm2m1d_cc_w_0_140_s_0_350 = '-2.09375e-13*ic_cap*ic_cap+-1.62500e-13*ic_cap+5.79000e-11'
+ mcm2m1d_cc_w_0_140_s_0_420 = '-1.12500e-13*ic_cap*ic_cap+-7.50000e-14*ic_cap+4.76000e-11'
+ mcm2m1d_cc_w_0_140_s_0_560 = '1.87500e-14*ic_cap*ic_cap+3.33000e-11'
+ mcm2m1d_cc_w_0_140_s_0_840 = '1.09375e-13*ic_cap*ic_cap+6.25000e-14*ic_cap+1.78000e-11'
+ mcm2m1d_cc_w_0_140_s_1_540 = '9.03125e-14*ic_cap*ic_cap+5.87500e-14*ic_cap+4.57000e-12'
+ mcm2m1d_cc_w_0_140_s_3_500 = '1.10937e-14*ic_cap*ic_cap+8.12500e-15*ic_cap+1.75000e-13'
+ mcm2m1d_cc_w_1_120_s_0_140 = '-5.09375e-13*ic_cap*ic_cap+-3.12500e-13*ic_cap+9.89000e-11'
+ mcm2m1d_cc_w_1_120_s_0_175 = '-5.00000e-13*ic_cap*ic_cap+-2.50000e-13*ic_cap+9.56000e-11'
+ mcm2m1d_cc_w_1_120_s_0_210 = '-3.78125e-13*ic_cap*ic_cap+-2.62500e-13*ic_cap+8.86000e-11'
+ mcm2m1d_cc_w_1_120_s_0_280 = '-2.31250e-13*ic_cap*ic_cap+-1.50000e-13*ic_cap+7.49000e-11'
+ mcm2m1d_cc_w_1_120_s_0_350 = '-1.09375e-13*ic_cap*ic_cap+-8.75000e-14*ic_cap+6.19000e-11'
+ mcm2m1d_cc_w_1_120_s_0_420 = '-1.56250e-14*ic_cap*ic_cap+-3.75000e-14*ic_cap+5.10000e-11'
+ mcm2m1d_cc_w_1_120_s_0_560 = '8.75000e-14*ic_cap*ic_cap+2.50000e-14*ic_cap+3.58000e-11'
+ mcm2m1d_cc_w_1_120_s_0_840 = '1.50000e-13*ic_cap*ic_cap+1.00000e-13*ic_cap+1.95000e-11'
+ mcm2m1d_cc_w_1_120_s_1_540 = '1.12500e-13*ic_cap*ic_cap+7.25000e-14*ic_cap+5.09000e-12'
+ mcm2m1d_cc_w_1_120_s_3_500 = '1.37500e-14*ic_cap*ic_cap+7.50000e-15*ic_cap+1.70000e-13'
+ mcm2m1d_cf_w_0_140_s_0_140 = '-1.01562e-13*ic_cap*ic_cap+-4.87500e-14*ic_cap+1.03000e-11'
+ mcm2m1d_cf_w_0_140_s_0_175 = '-1.43750e-13*ic_cap*ic_cap+-7.50000e-14*ic_cap+1.27000e-11'
+ mcm2m1d_cf_w_0_140_s_0_210 = '-1.78125e-13*ic_cap*ic_cap+-8.75000e-14*ic_cap+1.50000e-11'
+ mcm2m1d_cf_w_0_140_s_0_280 = '-2.53125e-13*ic_cap*ic_cap+-1.37500e-13*ic_cap+1.95000e-11'
+ mcm2m1d_cf_w_0_140_s_0_350 = '-3.09375e-13*ic_cap*ic_cap+-1.62500e-13*ic_cap+2.36000e-11'
+ mcm2m1d_cf_w_0_140_s_0_420 = '-3.68750e-13*ic_cap*ic_cap+-2.00000e-13*ic_cap+2.76000e-11'
+ mcm2m1d_cf_w_0_140_s_0_560 = '-4.46875e-13*ic_cap*ic_cap+-2.37500e-13*ic_cap+3.41000e-11'
+ mcm2m1d_cf_w_0_140_s_0_840 = '-5.40625e-13*ic_cap*ic_cap+-3.12500e-13*ic_cap+4.39000e-11'
+ mcm2m1d_cf_w_0_140_s_1_540 = '-5.68750e-13*ic_cap*ic_cap+-3.25000e-13*ic_cap+5.53000e-11'
+ mcm2m1d_cf_w_0_140_s_3_500 = '-5.06250e-13*ic_cap*ic_cap+-3.00000e-13*ic_cap+5.99000e-11'
+ mcm2m1d_cf_w_1_120_s_0_140 = '-1.03437e-13*ic_cap*ic_cap+-5.12500e-14*ic_cap+1.04000e-11'
+ mcm2m1d_cf_w_1_120_s_0_175 = '-1.43750e-13*ic_cap*ic_cap+-7.50000e-14*ic_cap+1.28000e-11'
+ mcm2m1d_cf_w_1_120_s_0_210 = '-1.78125e-13*ic_cap*ic_cap+-8.75000e-14*ic_cap+1.51000e-11'
+ mcm2m1d_cf_w_1_120_s_0_280 = '-2.43750e-13*ic_cap*ic_cap+-1.25000e-13*ic_cap+1.95000e-11'
+ mcm2m1d_cf_w_1_120_s_0_350 = '-3.09375e-13*ic_cap*ic_cap+-1.62500e-13*ic_cap+2.37000e-11'
+ mcm2m1d_cf_w_1_120_s_0_420 = '-3.59375e-13*ic_cap*ic_cap+-1.87500e-13*ic_cap+2.76000e-11'
+ mcm2m1d_cf_w_1_120_s_0_560 = '-4.46875e-13*ic_cap*ic_cap+-2.37500e-13*ic_cap+3.44000e-11'
+ mcm2m1d_cf_w_1_120_s_0_840 = '-5.34375e-13*ic_cap*ic_cap+-3.12500e-13*ic_cap+4.44000e-11'
+ mcm2m1d_cf_w_1_120_s_1_540 = '-5.59375e-13*ic_cap*ic_cap+-3.12500e-13*ic_cap+5.64000e-11'
+ mcm2m1d_cf_w_1_120_s_3_500 = '-4.71875e-13*ic_cap*ic_cap+-2.87500e-13*ic_cap+6.15000e-11'
+ mcm2m1f_ca_w_0_140_s_0_140 = '-2.96875e-06*ic_cap*ic_cap+-1.37500e-06*ic_cap+1.54000e-04'
+ mcm2m1f_ca_w_0_140_s_0_175 = '-2.96875e-06*ic_cap*ic_cap+-1.37500e-06*ic_cap+1.54000e-04'
+ mcm2m1f_ca_w_0_140_s_0_210 = '-2.96875e-06*ic_cap*ic_cap+-1.37500e-06*ic_cap+1.54000e-04'
+ mcm2m1f_ca_w_0_140_s_0_280 = '-2.96875e-06*ic_cap*ic_cap+-1.37500e-06*ic_cap+1.54000e-04'
+ mcm2m1f_ca_w_0_140_s_0_350 = '-2.96875e-06*ic_cap*ic_cap+-1.37500e-06*ic_cap+1.54000e-04'
+ mcm2m1f_ca_w_0_140_s_0_420 = '-2.96875e-06*ic_cap*ic_cap+-1.37500e-06*ic_cap+1.54000e-04'
+ mcm2m1f_ca_w_0_140_s_0_560 = '-2.96875e-06*ic_cap*ic_cap+-1.37500e-06*ic_cap+1.54000e-04'
+ mcm2m1f_ca_w_0_140_s_0_840 = '-2.96875e-06*ic_cap*ic_cap+-1.37500e-06*ic_cap+1.54000e-04'
+ mcm2m1f_ca_w_0_140_s_1_540 = '-2.96875e-06*ic_cap*ic_cap+-1.37500e-06*ic_cap+1.54000e-04'
+ mcm2m1f_ca_w_0_140_s_3_500 = '-2.96875e-06*ic_cap*ic_cap+-1.37500e-06*ic_cap+1.54000e-04'
+ mcm2m1f_ca_w_1_120_s_0_140 = '-2.96875e-06*ic_cap*ic_cap+-1.37500e-06*ic_cap+1.54000e-04'
+ mcm2m1f_ca_w_1_120_s_0_175 = '-2.96875e-06*ic_cap*ic_cap+-1.37500e-06*ic_cap+1.54000e-04'
+ mcm2m1f_ca_w_1_120_s_0_210 = '-2.96875e-06*ic_cap*ic_cap+-1.37500e-06*ic_cap+1.54000e-04'
+ mcm2m1f_ca_w_1_120_s_0_280 = '-2.96875e-06*ic_cap*ic_cap+-1.37500e-06*ic_cap+1.54000e-04'
+ mcm2m1f_ca_w_1_120_s_0_350 = '-2.96875e-06*ic_cap*ic_cap+-1.37500e-06*ic_cap+1.54000e-04'
+ mcm2m1f_ca_w_1_120_s_0_420 = '-2.96875e-06*ic_cap*ic_cap+-1.37500e-06*ic_cap+1.54000e-04'
+ mcm2m1f_ca_w_1_120_s_0_560 = '-2.96875e-06*ic_cap*ic_cap+-1.37500e-06*ic_cap+1.54000e-04'
+ mcm2m1f_ca_w_1_120_s_0_840 = '-2.96875e-06*ic_cap*ic_cap+-1.37500e-06*ic_cap+1.54000e-04'
+ mcm2m1f_ca_w_1_120_s_1_540 = '-2.96875e-06*ic_cap*ic_cap+-1.37500e-06*ic_cap+1.54000e-04'
+ mcm2m1f_ca_w_1_120_s_3_500 = '-2.96875e-06*ic_cap*ic_cap+-1.37500e-06*ic_cap+1.54000e-04'
+ mcm2m1f_cc_w_0_140_s_0_140 = '-6.84375e-13*ic_cap*ic_cap+-3.62500e-13*ic_cap+9.21000e-11'
+ mcm2m1f_cc_w_0_140_s_0_175 = '-6.62500e-13*ic_cap*ic_cap+-3.00000e-13*ic_cap+9.00000e-11'
+ mcm2m1f_cc_w_0_140_s_0_210 = '-5.56250e-13*ic_cap*ic_cap+-3.50000e-13*ic_cap+8.45000e-11'
+ mcm2m1f_cc_w_0_140_s_0_280 = '-3.25000e-13*ic_cap*ic_cap+-3.00000e-13*ic_cap+7.12000e-11'
+ mcm2m1f_cc_w_0_140_s_0_350 = '-2.18750e-13*ic_cap*ic_cap+-1.75000e-13*ic_cap+5.93000e-11'
+ mcm2m1f_cc_w_0_140_s_0_420 = '-1.15625e-13*ic_cap*ic_cap+-1.12500e-13*ic_cap+4.91000e-11'
+ mcm2m1f_cc_w_0_140_s_0_560 = '1.25000e-14*ic_cap*ic_cap+-2.50000e-14*ic_cap+3.50000e-11'
+ mcm2m1f_cc_w_0_140_s_0_840 = '1.00000e-13*ic_cap*ic_cap+5.00000e-14*ic_cap+1.97000e-11'
+ mcm2m1f_cc_w_0_140_s_1_540 = '9.59375e-14*ic_cap*ic_cap+6.12500e-14*ic_cap+5.79000e-12'
+ mcm2m1f_cc_w_0_140_s_3_500 = '1.81250e-14*ic_cap*ic_cap+1.50000e-14*ic_cap+3.20000e-13'
+ mcm2m1f_cc_w_1_120_s_0_140 = '-4.93750e-13*ic_cap*ic_cap+-2.50000e-13*ic_cap+1.01000e-10'
+ mcm2m1f_cc_w_1_120_s_0_175 = '-5.12500e-13*ic_cap*ic_cap+-2.75000e-13*ic_cap+9.83000e-11'
+ mcm2m1f_cc_w_1_120_s_0_210 = '-3.84375e-13*ic_cap*ic_cap+-2.62500e-13*ic_cap+9.13000e-11'
+ mcm2m1f_cc_w_1_120_s_0_280 = '-2.28125e-13*ic_cap*ic_cap+-1.62500e-13*ic_cap+7.75000e-11'
+ mcm2m1f_cc_w_1_120_s_0_350 = '-1.28125e-13*ic_cap*ic_cap+-1.12500e-13*ic_cap+6.48000e-11'
+ mcm2m1f_cc_w_1_120_s_0_420 = '-3.12500e-14*ic_cap*ic_cap+-5.00000e-14*ic_cap+5.39000e-11'
+ mcm2m1f_cc_w_1_120_s_0_560 = '8.75000e-14*ic_cap*ic_cap+5.00000e-14*ic_cap+3.86000e-11'
+ mcm2m1f_cc_w_1_120_s_0_840 = '1.53125e-13*ic_cap*ic_cap+8.75000e-14*ic_cap+2.21000e-11'
+ mcm2m1f_cc_w_1_120_s_1_540 = '1.28437e-13*ic_cap*ic_cap+8.12500e-14*ic_cap+6.77000e-12'
+ mcm2m1f_cc_w_1_120_s_3_500 = '2.35938e-14*ic_cap*ic_cap+1.43750e-14*ic_cap+3.65000e-13'
+ mcm2m1f_cf_w_0_140_s_0_140 = '-1.03125e-13*ic_cap*ic_cap+-5.00000e-14*ic_cap+9.79000e-12'
+ mcm2m1f_cf_w_0_140_s_0_175 = '-1.40938e-13*ic_cap*ic_cap+-6.37500e-14*ic_cap+1.20000e-11'
+ mcm2m1f_cf_w_0_140_s_0_210 = '-1.71875e-13*ic_cap*ic_cap+-8.75000e-14*ic_cap+1.42000e-11'
+ mcm2m1f_cf_w_0_140_s_0_280 = '-2.43750e-13*ic_cap*ic_cap+-1.25000e-13*ic_cap+1.84000e-11'
+ mcm2m1f_cf_w_0_140_s_0_350 = '-3.03125e-13*ic_cap*ic_cap+-1.62500e-13*ic_cap+2.23000e-11'
+ mcm2m1f_cf_w_0_140_s_0_420 = '-3.59375e-13*ic_cap*ic_cap+-1.87500e-13*ic_cap+2.61000e-11'
+ mcm2m1f_cf_w_0_140_s_0_560 = '-4.37500e-13*ic_cap*ic_cap+-2.25000e-13*ic_cap+3.22000e-11'
+ mcm2m1f_cf_w_0_140_s_0_840 = '-5.34375e-13*ic_cap*ic_cap+-2.87500e-13*ic_cap+4.17000e-11'
+ mcm2m1f_cf_w_0_140_s_1_540 = '-5.68750e-13*ic_cap*ic_cap+-3.25000e-13*ic_cap+5.32000e-11'
+ mcm2m1f_cf_w_0_140_s_3_500 = '-5.00000e-13*ic_cap*ic_cap+-3.00000e-13*ic_cap+5.86000e-11'
+ mcm2m1f_cf_w_1_120_s_0_140 = '-1.01562e-13*ic_cap*ic_cap+-4.87500e-14*ic_cap+9.82000e-12'
+ mcm2m1f_cf_w_1_120_s_0_175 = '-1.41562e-13*ic_cap*ic_cap+-6.62500e-14*ic_cap+1.21000e-11'
+ mcm2m1f_cf_w_1_120_s_0_210 = '-1.78125e-13*ic_cap*ic_cap+-8.75000e-14*ic_cap+1.43000e-11'
+ mcm2m1f_cf_w_1_120_s_0_280 = '-2.37500e-13*ic_cap*ic_cap+-1.25000e-13*ic_cap+1.84000e-11'
+ mcm2m1f_cf_w_1_120_s_0_350 = '-3.00000e-13*ic_cap*ic_cap+-1.50000e-13*ic_cap+2.24000e-11'
+ mcm2m1f_cf_w_1_120_s_0_420 = '-3.53125e-13*ic_cap*ic_cap+-1.87500e-13*ic_cap+2.61000e-11'
+ mcm2m1f_cf_w_1_120_s_0_560 = '-4.34375e-13*ic_cap*ic_cap+-2.37500e-13*ic_cap+3.25000e-11'
+ mcm2m1f_cf_w_1_120_s_0_840 = '-5.21875e-13*ic_cap*ic_cap+-2.87500e-13*ic_cap+4.21000e-11'
+ mcm2m1f_cf_w_1_120_s_1_540 = '-5.50000e-13*ic_cap*ic_cap+-3.25000e-13*ic_cap+5.43000e-11'
+ mcm2m1f_cf_w_1_120_s_3_500 = '-4.75000e-13*ic_cap*ic_cap+-2.75000e-13*ic_cap+6.08000e-11'
+ mcm2m1l1_ca_w_0_140_s_0_140 = '-4.62500e-06*ic_cap*ic_cap+-2.50000e-06*ic_cap+2.42000e-04'
+ mcm2m1l1_ca_w_0_140_s_0_175 = '-4.62500e-06*ic_cap*ic_cap+-2.50000e-06*ic_cap+2.42000e-04'
+ mcm2m1l1_ca_w_0_140_s_0_210 = '-4.62500e-06*ic_cap*ic_cap+-2.50000e-06*ic_cap+2.42000e-04'
+ mcm2m1l1_ca_w_0_140_s_0_280 = '-4.62500e-06*ic_cap*ic_cap+-2.50000e-06*ic_cap+2.42000e-04'
+ mcm2m1l1_ca_w_0_140_s_0_350 = '-4.62500e-06*ic_cap*ic_cap+-2.50000e-06*ic_cap+2.42000e-04'
+ mcm2m1l1_ca_w_0_140_s_0_420 = '-4.62500e-06*ic_cap*ic_cap+-2.50000e-06*ic_cap+2.42000e-04'
+ mcm2m1l1_ca_w_0_140_s_0_560 = '-4.62500e-06*ic_cap*ic_cap+-2.50000e-06*ic_cap+2.42000e-04'
+ mcm2m1l1_ca_w_0_140_s_0_840 = '-4.62500e-06*ic_cap*ic_cap+-2.50000e-06*ic_cap+2.42000e-04'
+ mcm2m1l1_ca_w_0_140_s_1_540 = '-4.62500e-06*ic_cap*ic_cap+-2.50000e-06*ic_cap+2.42000e-04'
+ mcm2m1l1_ca_w_0_140_s_3_500 = '-4.62500e-06*ic_cap*ic_cap+-2.50000e-06*ic_cap+2.42000e-04'
+ mcm2m1l1_ca_w_1_120_s_0_140 = '-4.62500e-06*ic_cap*ic_cap+-2.50000e-06*ic_cap+2.42000e-04'
+ mcm2m1l1_ca_w_1_120_s_0_175 = '-4.62500e-06*ic_cap*ic_cap+-2.50000e-06*ic_cap+2.42000e-04'
+ mcm2m1l1_ca_w_1_120_s_0_210 = '-4.62500e-06*ic_cap*ic_cap+-2.50000e-06*ic_cap+2.42000e-04'
+ mcm2m1l1_ca_w_1_120_s_0_280 = '-4.62500e-06*ic_cap*ic_cap+-2.50000e-06*ic_cap+2.42000e-04'
+ mcm2m1l1_ca_w_1_120_s_0_350 = '-4.62500e-06*ic_cap*ic_cap+-2.50000e-06*ic_cap+2.42000e-04'
+ mcm2m1l1_ca_w_1_120_s_0_420 = '-4.62500e-06*ic_cap*ic_cap+-2.50000e-06*ic_cap+2.42000e-04'
+ mcm2m1l1_ca_w_1_120_s_0_560 = '-4.62500e-06*ic_cap*ic_cap+-2.50000e-06*ic_cap+2.42000e-04'
+ mcm2m1l1_ca_w_1_120_s_0_840 = '-4.62500e-06*ic_cap*ic_cap+-2.50000e-06*ic_cap+2.42000e-04'
+ mcm2m1l1_ca_w_1_120_s_1_540 = '-4.62500e-06*ic_cap*ic_cap+-2.50000e-06*ic_cap+2.42000e-04'
+ mcm2m1l1_ca_w_1_120_s_3_500 = '-4.62500e-06*ic_cap*ic_cap+-2.50000e-06*ic_cap+2.42000e-04'
+ mcm2m1l1_cc_w_0_140_s_0_140 = '-5.56250e-13*ic_cap*ic_cap+-3.00000e-13*ic_cap+8.35000e-11'
+ mcm2m1l1_cc_w_0_140_s_0_175 = '-5.06250e-13*ic_cap*ic_cap+-2.25000e-13*ic_cap+8.06000e-11'
+ mcm2m1l1_cc_w_0_140_s_0_210 = '-3.56250e-13*ic_cap*ic_cap+-3.00000e-13*ic_cap+7.38000e-11'
+ mcm2m1l1_cc_w_0_140_s_0_280 = '-1.90625e-13*ic_cap*ic_cap+-1.37500e-13*ic_cap+6.02000e-11'
+ mcm2m1l1_cc_w_0_140_s_0_350 = '-6.25000e-14*ic_cap*ic_cap+-5.00000e-14*ic_cap+4.74000e-11'
+ mcm2m1l1_cc_w_0_140_s_0_420 = '4.06250e-14*ic_cap*ic_cap+3.75000e-14*ic_cap+3.68000e-11'
+ mcm2m1l1_cc_w_0_140_s_0_560 = '1.43750e-13*ic_cap*ic_cap+1.00000e-13*ic_cap+2.26000e-11'
+ mcm2m1l1_cc_w_0_140_s_0_840 = '1.68125e-13*ic_cap*ic_cap+1.25000e-13*ic_cap+8.81000e-12'
+ mcm2m1l1_cc_w_0_140_s_1_540 = '5.46875e-14*ic_cap*ic_cap+4.50000e-14*ic_cap+9.45000e-13'
+ mcm2m1l1_cc_w_0_140_s_3_500 = '1.71875e-15*ic_cap*ic_cap+-4.37500e-15*ic_cap+2.50000e-14'
+ mcm2m1l1_cc_w_1_120_s_0_140 = '-3.93750e-13*ic_cap*ic_cap+-1.50000e-13*ic_cap+8.49000e-11'
+ mcm2m1l1_cc_w_1_120_s_0_175 = '-3.81250e-13*ic_cap*ic_cap+-1.50000e-13*ic_cap+8.16000e-11'
+ mcm2m1l1_cc_w_1_120_s_0_210 = '-2.87500e-13*ic_cap*ic_cap+-1.50000e-13*ic_cap+7.54000e-11'
+ mcm2m1l1_cc_w_1_120_s_0_280 = '-1.03125e-13*ic_cap*ic_cap+-6.25000e-14*ic_cap+6.07000e-11'
+ mcm2m1l1_cc_w_1_120_s_0_350 = '3.12500e-15*ic_cap*ic_cap+1.25000e-14*ic_cap+4.79000e-11'
+ mcm2m1l1_cc_w_1_120_s_0_420 = '9.37500e-14*ic_cap*ic_cap+1.25000e-13*ic_cap+3.72000e-11'
+ mcm2m1l1_cc_w_1_120_s_0_560 = '1.78125e-13*ic_cap*ic_cap+1.37500e-13*ic_cap+2.28000e-11'
+ mcm2m1l1_cc_w_1_120_s_0_840 = '1.81250e-13*ic_cap*ic_cap+1.25000e-13*ic_cap+9.00000e-12'
+ mcm2m1l1_cc_w_1_120_s_1_540 = '5.78125e-14*ic_cap*ic_cap+5.62500e-14*ic_cap+9.50000e-13'
+ mcm2m1l1_cf_w_0_140_s_0_140 = '-1.62500e-13*ic_cap*ic_cap+-1.00000e-13*ic_cap+1.54000e-11'
+ mcm2m1l1_cf_w_0_140_s_0_175 = '-2.28125e-13*ic_cap*ic_cap+-1.37500e-13*ic_cap+1.92000e-11'
+ mcm2m1l1_cf_w_0_140_s_0_210 = '-2.90625e-13*ic_cap*ic_cap+-1.62500e-13*ic_cap+2.28000e-11'
+ mcm2m1l1_cf_w_0_140_s_0_280 = '-4.03125e-13*ic_cap*ic_cap+-2.37500e-13*ic_cap+2.96000e-11'
+ mcm2m1l1_cf_w_0_140_s_0_350 = '-5.12500e-13*ic_cap*ic_cap+-3.00000e-13*ic_cap+3.60000e-11'
+ mcm2m1l1_cf_w_0_140_s_0_420 = '-5.90625e-13*ic_cap*ic_cap+-3.62500e-13*ic_cap+4.16000e-11'
+ mcm2m1l1_cf_w_0_140_s_0_560 = '-7.15625e-13*ic_cap*ic_cap+-4.37500e-13*ic_cap+5.08000e-11'
+ mcm2m1l1_cf_w_0_140_s_0_840 = '-8.03125e-13*ic_cap*ic_cap+-4.87500e-13*ic_cap+6.23000e-11'
+ mcm2m1l1_cf_w_0_140_s_1_540 = '-7.40625e-13*ic_cap*ic_cap+-4.62500e-13*ic_cap+7.06000e-11'
+ mcm2m1l1_cf_w_0_140_s_3_500 = '-6.87500e-13*ic_cap*ic_cap+-4.25000e-13*ic_cap+7.20000e-11'
+ mcm2m1l1_cf_w_1_120_s_0_140 = '-1.62500e-13*ic_cap*ic_cap+-1.00000e-13*ic_cap+1.55000e-11'
+ mcm2m1l1_cf_w_1_120_s_0_175 = '-2.28125e-13*ic_cap*ic_cap+-1.37500e-13*ic_cap+1.93000e-11'
+ mcm2m1l1_cf_w_1_120_s_0_210 = '-2.93750e-13*ic_cap*ic_cap+-1.75000e-13*ic_cap+2.29000e-11'
+ mcm2m1l1_cf_w_1_120_s_0_280 = '-4.03125e-13*ic_cap*ic_cap+-2.37500e-13*ic_cap+2.97000e-11'
+ mcm2m1l1_cf_w_1_120_s_0_350 = '-5.00000e-13*ic_cap*ic_cap+-3.00000e-13*ic_cap+3.60000e-11'
+ mcm2m1l1_cf_w_1_120_s_0_420 = '-5.87500e-13*ic_cap*ic_cap+-3.50000e-13*ic_cap+4.17000e-11'
+ mcm2m1l1_cf_w_1_120_s_0_560 = '-7.06250e-13*ic_cap*ic_cap+-4.25000e-13*ic_cap+5.10000e-11'
+ mcm2m1l1_cf_w_1_120_s_0_840 = '-7.87500e-13*ic_cap*ic_cap+-4.75000e-13*ic_cap+6.26000e-11'
+ mcm2m1l1_cf_w_1_120_s_1_540 = '-7.09375e-13*ic_cap*ic_cap+-4.37500e-13*ic_cap+7.09000e-11'
+ mcm2m1l1_cf_w_1_120_s_3_500 = '-6.62500e-13*ic_cap*ic_cap+-4.00000e-13*ic_cap+7.24000e-11'
+ mcm2m1p1_ca_w_0_140_s_0_140 = '-3.34375e-06*ic_cap*ic_cap+-1.62500e-06*ic_cap+1.73000e-04'
+ mcm2m1p1_ca_w_0_140_s_0_175 = '-3.34375e-06*ic_cap*ic_cap+-1.62500e-06*ic_cap+1.73000e-04'
+ mcm2m1p1_ca_w_0_140_s_0_210 = '-3.34375e-06*ic_cap*ic_cap+-1.62500e-06*ic_cap+1.73000e-04'
+ mcm2m1p1_ca_w_0_140_s_0_280 = '-3.34375e-06*ic_cap*ic_cap+-1.62500e-06*ic_cap+1.73000e-04'
+ mcm2m1p1_ca_w_0_140_s_0_350 = '-3.34375e-06*ic_cap*ic_cap+-1.62500e-06*ic_cap+1.73000e-04'
+ mcm2m1p1_ca_w_0_140_s_0_420 = '-3.34375e-06*ic_cap*ic_cap+-1.62500e-06*ic_cap+1.73000e-04'
+ mcm2m1p1_ca_w_0_140_s_0_560 = '-3.34375e-06*ic_cap*ic_cap+-1.62500e-06*ic_cap+1.73000e-04'
+ mcm2m1p1_ca_w_0_140_s_0_840 = '-3.34375e-06*ic_cap*ic_cap+-1.62500e-06*ic_cap+1.73000e-04'
+ mcm2m1p1_ca_w_0_140_s_1_540 = '-3.34375e-06*ic_cap*ic_cap+-1.62500e-06*ic_cap+1.73000e-04'
+ mcm2m1p1_ca_w_0_140_s_3_500 = '-3.34375e-06*ic_cap*ic_cap+-1.62500e-06*ic_cap+1.73000e-04'
+ mcm2m1p1_ca_w_1_120_s_0_140 = '-3.34375e-06*ic_cap*ic_cap+-1.62500e-06*ic_cap+1.73000e-04'
+ mcm2m1p1_ca_w_1_120_s_0_175 = '-3.34375e-06*ic_cap*ic_cap+-1.62500e-06*ic_cap+1.73000e-04'
+ mcm2m1p1_ca_w_1_120_s_0_210 = '-3.34375e-06*ic_cap*ic_cap+-1.62500e-06*ic_cap+1.73000e-04'
+ mcm2m1p1_ca_w_1_120_s_0_280 = '-3.34375e-06*ic_cap*ic_cap+-1.62500e-06*ic_cap+1.73000e-04'
+ mcm2m1p1_ca_w_1_120_s_0_350 = '-3.34375e-06*ic_cap*ic_cap+-1.62500e-06*ic_cap+1.73000e-04'
+ mcm2m1p1_ca_w_1_120_s_0_420 = '-3.34375e-06*ic_cap*ic_cap+-1.62500e-06*ic_cap+1.73000e-04'
+ mcm2m1p1_ca_w_1_120_s_0_560 = '-3.34375e-06*ic_cap*ic_cap+-1.62500e-06*ic_cap+1.73000e-04'
+ mcm2m1p1_ca_w_1_120_s_0_840 = '-3.34375e-06*ic_cap*ic_cap+-1.62500e-06*ic_cap+1.73000e-04'
+ mcm2m1p1_ca_w_1_120_s_1_540 = '-3.34375e-06*ic_cap*ic_cap+-1.62500e-06*ic_cap+1.73000e-04'
+ mcm2m1p1_ca_w_1_120_s_3_500 = '-3.34375e-06*ic_cap*ic_cap+-1.62500e-06*ic_cap+1.73000e-04'
+ mcm2m1p1_cc_w_0_140_s_0_140 = '-6.53125e-13*ic_cap*ic_cap+-3.62500e-13*ic_cap+9.03000e-11'
+ mcm2m1p1_cc_w_0_140_s_0_175 = '-6.31250e-13*ic_cap*ic_cap+-3.00000e-13*ic_cap+8.77000e-11'
+ mcm2m1p1_cc_w_0_140_s_0_210 = '-4.75000e-13*ic_cap*ic_cap+-3.25000e-13*ic_cap+8.13000e-11'
+ mcm2m1p1_cc_w_0_140_s_0_280 = '-2.65625e-13*ic_cap*ic_cap+-2.62500e-13*ic_cap+6.80000e-11'
+ mcm2m1p1_cc_w_0_140_s_0_350 = '-1.59375e-13*ic_cap*ic_cap+-1.37500e-13*ic_cap+5.59000e-11'
+ mcm2m1p1_cc_w_0_140_s_0_420 = '-5.93750e-14*ic_cap*ic_cap+-3.75000e-14*ic_cap+4.55000e-11'
+ mcm2m1p1_cc_w_0_140_s_0_560 = '8.12500e-14*ic_cap*ic_cap+2.50000e-14*ic_cap+3.09000e-11'
+ mcm2m1p1_cc_w_0_140_s_0_840 = '1.56250e-13*ic_cap*ic_cap+7.50000e-14*ic_cap+1.56000e-11'
+ mcm2m1p1_cc_w_0_140_s_1_540 = '1.05000e-13*ic_cap*ic_cap+7.00000e-14*ic_cap+3.31000e-12'
+ mcm2m1p1_cc_w_0_140_s_3_500 = '6.40625e-15*ic_cap*ic_cap+5.62500e-15*ic_cap+1.25000e-13'
+ mcm2m1p1_cc_w_1_120_s_0_140 = '-4.31250e-13*ic_cap*ic_cap+-2.50000e-13*ic_cap+9.55000e-11'
+ mcm2m1p1_cc_w_1_120_s_0_175 = '-4.34375e-13*ic_cap*ic_cap+-1.87500e-13*ic_cap+9.24000e-11'
+ mcm2m1p1_cc_w_1_120_s_0_210 = '-3.68750e-13*ic_cap*ic_cap+-2.00000e-13*ic_cap+8.64000e-11'
+ mcm2m1p1_cc_w_1_120_s_0_280 = '-1.65625e-13*ic_cap*ic_cap+-1.12500e-13*ic_cap+7.16000e-11'
+ mcm2m1p1_cc_w_1_120_s_0_350 = '-5.93750e-14*ic_cap*ic_cap+-1.25000e-14*ic_cap+5.87000e-11'
+ mcm2m1p1_cc_w_1_120_s_0_420 = '3.12500e-14*ic_cap*ic_cap+4.79000e-11'
+ mcm2m1p1_cc_w_1_120_s_0_560 = '1.59375e-13*ic_cap*ic_cap+8.75000e-14*ic_cap+3.25000e-11'
+ mcm2m1p1_cc_w_1_120_s_0_840 = '2.03125e-13*ic_cap*ic_cap+1.12500e-13*ic_cap+1.66000e-11'
+ mcm2m1p1_cc_w_1_120_s_1_540 = '1.26250e-13*ic_cap*ic_cap+9.00000e-14*ic_cap+3.54000e-12'
+ mcm2m1p1_cc_w_1_120_s_3_500 = '9.06250e-15*ic_cap*ic_cap+7.50000e-15*ic_cap+1.20000e-13'
+ mcm2m1p1_cf_w_0_140_s_0_140 = '-1.19688e-13*ic_cap*ic_cap+-5.87500e-14*ic_cap+1.11000e-11'
+ mcm2m1p1_cf_w_0_140_s_0_175 = '-1.65625e-13*ic_cap*ic_cap+-8.75000e-14*ic_cap+1.37000e-11'
+ mcm2m1p1_cf_w_0_140_s_0_210 = '-2.06250e-13*ic_cap*ic_cap+-1.00000e-13*ic_cap+1.62000e-11'
+ mcm2m1p1_cf_w_0_140_s_0_280 = '-2.87500e-13*ic_cap*ic_cap+-1.50000e-13*ic_cap+2.10000e-11'
+ mcm2m1p1_cf_w_0_140_s_0_350 = '-3.46875e-13*ic_cap*ic_cap+-1.87500e-13*ic_cap+2.54000e-11'
+ mcm2m1p1_cf_w_0_140_s_0_420 = '-4.15625e-13*ic_cap*ic_cap+-2.37500e-13*ic_cap+2.97000e-11'
+ mcm2m1p1_cf_w_0_140_s_0_560 = '-5.12500e-13*ic_cap*ic_cap+-2.75000e-13*ic_cap+3.67000e-11'
+ mcm2m1p1_cf_w_0_140_s_0_840 = '-6.12500e-13*ic_cap*ic_cap+-3.50000e-13*ic_cap+4.70000e-11'
+ mcm2m1p1_cf_w_0_140_s_1_540 = '-6.15625e-13*ic_cap*ic_cap+-3.87500e-13*ic_cap+5.80000e-11'
+ mcm2m1p1_cf_w_0_140_s_3_500 = '-5.43750e-13*ic_cap*ic_cap+-3.00000e-13*ic_cap+6.16000e-11'
+ mcm2m1p1_cf_w_1_120_s_0_140 = '-1.19063e-13*ic_cap*ic_cap+-5.87500e-14*ic_cap+1.12000e-11'
+ mcm2m1p1_cf_w_1_120_s_0_175 = '-1.65625e-13*ic_cap*ic_cap+-8.75000e-14*ic_cap+1.38000e-11'
+ mcm2m1p1_cf_w_1_120_s_0_210 = '-2.09375e-13*ic_cap*ic_cap+-1.12500e-13*ic_cap+1.63000e-11'
+ mcm2m1p1_cf_w_1_120_s_0_280 = '-2.84375e-13*ic_cap*ic_cap+-1.37500e-13*ic_cap+2.11000e-11'
+ mcm2m1p1_cf_w_1_120_s_0_350 = '-3.53125e-13*ic_cap*ic_cap+-1.87500e-13*ic_cap+2.56000e-11'
+ mcm2m1p1_cf_w_1_120_s_0_420 = '-4.12500e-13*ic_cap*ic_cap+-2.25000e-13*ic_cap+2.98000e-11'
+ mcm2m1p1_cf_w_1_120_s_0_560 = '-5.09375e-13*ic_cap*ic_cap+-2.87500e-13*ic_cap+3.70000e-11'
+ mcm2m1p1_cf_w_1_120_s_0_840 = '-6.06250e-13*ic_cap*ic_cap+-3.50000e-13*ic_cap+4.75000e-11'
+ mcm2m1p1_cf_w_1_120_s_1_540 = '-5.93750e-13*ic_cap*ic_cap+-3.75000e-13*ic_cap+5.88000e-11'
+ mcm2m1p1_cf_w_1_120_s_3_500 = '-5.06250e-13*ic_cap*ic_cap+-2.75000e-13*ic_cap+6.28000e-11'
+ mcm2p1_ca_w_0_140_s_0_140 = '-3.15625e-07*ic_cap*ic_cap+-1.87500e-07*ic_cap+2.47000e-05'
+ mcm2p1_ca_w_0_140_s_0_175 = '-3.15625e-07*ic_cap*ic_cap+-1.87500e-07*ic_cap+2.47000e-05'
+ mcm2p1_ca_w_0_140_s_0_210 = '-3.15625e-07*ic_cap*ic_cap+-1.87500e-07*ic_cap+2.47000e-05'
+ mcm2p1_ca_w_0_140_s_0_280 = '-3.15625e-07*ic_cap*ic_cap+-1.87500e-07*ic_cap+2.47000e-05'
+ mcm2p1_ca_w_0_140_s_0_350 = '-3.15625e-07*ic_cap*ic_cap+-1.87500e-07*ic_cap+2.47000e-05'
+ mcm2p1_ca_w_0_140_s_0_420 = '-3.15625e-07*ic_cap*ic_cap+-1.87500e-07*ic_cap+2.47000e-05'
+ mcm2p1_ca_w_0_140_s_0_560 = '-3.15625e-07*ic_cap*ic_cap+-1.87500e-07*ic_cap+2.47000e-05'
+ mcm2p1_ca_w_0_140_s_0_840 = '-3.15625e-07*ic_cap*ic_cap+-1.87500e-07*ic_cap+2.47000e-05'
+ mcm2p1_ca_w_0_140_s_1_540 = '-3.15625e-07*ic_cap*ic_cap+-1.87500e-07*ic_cap+2.47000e-05'
+ mcm2p1_ca_w_0_140_s_3_500 = '-3.15625e-07*ic_cap*ic_cap+-1.87500e-07*ic_cap+2.47000e-05'
+ mcm2p1_ca_w_1_120_s_0_140 = '-3.15625e-07*ic_cap*ic_cap+-1.87500e-07*ic_cap+2.47000e-05'
+ mcm2p1_ca_w_1_120_s_0_175 = '-3.15625e-07*ic_cap*ic_cap+-1.87500e-07*ic_cap+2.47000e-05'
+ mcm2p1_ca_w_1_120_s_0_210 = '-3.15625e-07*ic_cap*ic_cap+-1.87500e-07*ic_cap+2.47000e-05'
+ mcm2p1_ca_w_1_120_s_0_280 = '-3.15625e-07*ic_cap*ic_cap+-1.87500e-07*ic_cap+2.47000e-05'
+ mcm2p1_ca_w_1_120_s_0_350 = '-3.15625e-07*ic_cap*ic_cap+-1.87500e-07*ic_cap+2.47000e-05'
+ mcm2p1_ca_w_1_120_s_0_420 = '-3.15625e-07*ic_cap*ic_cap+-1.87500e-07*ic_cap+2.47000e-05'
+ mcm2p1_ca_w_1_120_s_0_560 = '-3.15625e-07*ic_cap*ic_cap+-1.87500e-07*ic_cap+2.47000e-05'
+ mcm2p1_ca_w_1_120_s_0_840 = '-3.15625e-07*ic_cap*ic_cap+-1.87500e-07*ic_cap+2.47000e-05'
+ mcm2p1_ca_w_1_120_s_1_540 = '-3.15625e-07*ic_cap*ic_cap+-1.87500e-07*ic_cap+2.47000e-05'
+ mcm2p1_ca_w_1_120_s_3_500 = '-3.15625e-07*ic_cap*ic_cap+-1.87500e-07*ic_cap+2.47000e-05'
+ mcm2p1_cc_w_0_140_s_0_140 = '-9.37500e-13*ic_cap*ic_cap+-5.25000e-13*ic_cap+1.05000e-10'
+ mcm2p1_cc_w_0_140_s_0_175 = '-8.78125e-13*ic_cap*ic_cap+-5.62500e-13*ic_cap+1.03000e-10'
+ mcm2p1_cc_w_0_140_s_0_210 = '-7.56250e-13*ic_cap*ic_cap+-4.25000e-13*ic_cap+9.77000e-11'
+ mcm2p1_cc_w_0_140_s_0_280 = '-6.21875e-13*ic_cap*ic_cap+-3.87500e-13*ic_cap+8.77000e-11'
+ mcm2p1_cc_w_0_140_s_0_350 = '-4.53125e-13*ic_cap*ic_cap+-3.12500e-13*ic_cap+7.60000e-11'
+ mcm2p1_cc_w_0_140_s_0_420 = '-3.25000e-13*ic_cap*ic_cap+-2.25000e-13*ic_cap+6.66000e-11'
+ mcm2p1_cc_w_0_140_s_0_560 = '-2.12500e-13*ic_cap*ic_cap+-1.25000e-13*ic_cap+5.44000e-11'
+ mcm2p1_cc_w_0_140_s_0_840 = '-7.81250e-14*ic_cap*ic_cap+-6.25000e-14*ic_cap+4.04000e-11'
+ mcm2p1_cc_w_0_140_s_1_540 = '2.81250e-14*ic_cap*ic_cap+1.25000e-14*ic_cap+2.46000e-11'
+ mcm2p1_cc_w_0_140_s_3_500 = '6.56250e-14*ic_cap*ic_cap+3.75000e-14*ic_cap+1.01000e-11'
+ mcm2p1_cc_w_1_120_s_0_140 = '-7.81250e-13*ic_cap*ic_cap+-3.75000e-13*ic_cap+1.30000e-10'
+ mcm2p1_cc_w_1_120_s_0_175 = '-7.18750e-13*ic_cap*ic_cap+-3.75000e-13*ic_cap+1.26000e-10'
+ mcm2p1_cc_w_1_120_s_0_210 = '-6.25000e-13*ic_cap*ic_cap+-2.50000e-13*ic_cap+1.20000e-10'
+ mcm2p1_cc_w_1_120_s_0_280 = '-5.21875e-13*ic_cap*ic_cap+-3.37500e-13*ic_cap+1.07000e-10'
+ mcm2p1_cc_w_1_120_s_0_350 = '-3.46875e-13*ic_cap*ic_cap+-2.12500e-13*ic_cap+9.38000e-11'
+ mcm2p1_cc_w_1_120_s_0_420 = '-2.46875e-13*ic_cap*ic_cap+-1.37500e-13*ic_cap+8.32000e-11'
+ mcm2p1_cc_w_1_120_s_0_560 = '-1.25000e-13*ic_cap*ic_cap+-7.50000e-14*ic_cap+6.85000e-11'
+ mcm2p1_cc_w_1_120_s_0_840 = '-1.56250e-14*ic_cap*ic_cap+-1.25000e-14*ic_cap+5.16000e-11'
+ mcm2p1_cc_w_1_120_s_1_540 = '6.25000e-14*ic_cap*ic_cap+5.00000e-14*ic_cap+3.27000e-11'
+ mcm2p1_cc_w_1_120_s_3_500 = '8.43750e-14*ic_cap*ic_cap+6.25000e-14*ic_cap+1.48000e-11'
+ mcm2p1_cf_w_0_140_s_0_140 = '-6.25000e-15*ic_cap*ic_cap+-5.00000e-15*ic_cap+1.72000e-12'
+ mcm2p1_cf_w_0_140_s_0_175 = '-1.09375e-14*ic_cap*ic_cap+-8.75000e-15*ic_cap+2.14000e-12'
+ mcm2p1_cf_w_0_140_s_0_210 = '-1.71875e-14*ic_cap*ic_cap+-1.12500e-14*ic_cap+2.58000e-12'
+ mcm2p1_cf_w_0_140_s_0_280 = '-2.75000e-14*ic_cap*ic_cap+-1.75000e-14*ic_cap+3.42000e-12'
+ mcm2p1_cf_w_0_140_s_0_350 = '-3.78125e-14*ic_cap*ic_cap+-2.37500e-14*ic_cap+4.24000e-12'
+ mcm2p1_cf_w_0_140_s_0_420 = '-4.84375e-14*ic_cap*ic_cap+-3.12500e-14*ic_cap+5.10000e-12'
+ mcm2p1_cf_w_0_140_s_0_560 = '-6.81250e-14*ic_cap*ic_cap+-4.25000e-14*ic_cap+6.65000e-12'
+ mcm2p1_cf_w_0_140_s_0_840 = '-1.02500e-13*ic_cap*ic_cap+-6.25000e-14*ic_cap+9.62000e-12'
+ mcm2p1_cf_w_0_140_s_1_540 = '-1.65625e-13*ic_cap*ic_cap+-1.12500e-13*ic_cap+1.59000e-11'
+ mcm2p1_cf_w_0_140_s_3_500 = '-2.31250e-13*ic_cap*ic_cap+-1.50000e-13*ic_cap+2.62000e-11'
+ mcm2p1_cf_w_1_120_s_0_140 = '-7.18750e-15*ic_cap*ic_cap+-6.25000e-15*ic_cap+1.78000e-12'
+ mcm2p1_cf_w_1_120_s_0_175 = '-1.28125e-14*ic_cap*ic_cap+-8.75000e-15*ic_cap+2.21000e-12'
+ mcm2p1_cf_w_1_120_s_0_210 = '-1.84375e-14*ic_cap*ic_cap+-1.12500e-14*ic_cap+2.64000e-12'
+ mcm2p1_cf_w_1_120_s_0_280 = '-2.87500e-14*ic_cap*ic_cap+-1.75000e-14*ic_cap+3.48000e-12'
+ mcm2p1_cf_w_1_120_s_0_350 = '-3.90625e-14*ic_cap*ic_cap+-2.37500e-14*ic_cap+4.31000e-12'
+ mcm2p1_cf_w_1_120_s_0_420 = '-4.96875e-14*ic_cap*ic_cap+-2.87500e-14*ic_cap+5.14000e-12'
+ mcm2p1_cf_w_1_120_s_0_560 = '-6.84375e-14*ic_cap*ic_cap+-4.37500e-14*ic_cap+6.72000e-12'
+ mcm2p1_cf_w_1_120_s_0_840 = '-1.03750e-13*ic_cap*ic_cap+-6.25000e-14*ic_cap+9.73000e-12'
+ mcm2p1_cf_w_1_120_s_1_540 = '-1.68750e-13*ic_cap*ic_cap+-1.00000e-13*ic_cap+1.62000e-11'
+ mcm2p1_cf_w_1_120_s_3_500 = '-2.40625e-13*ic_cap*ic_cap+-1.62500e-13*ic_cap+2.79000e-11'
+ mcm2p1f_ca_w_0_150_s_0_210 = '-1.73750e-06*ic_cap*ic_cap+-9.50000e-07*ic_cap+1.31000e-04'
+ mcm2p1f_ca_w_0_150_s_0_263 = '-1.73750e-06*ic_cap*ic_cap+-9.50000e-07*ic_cap+1.31000e-04'
+ mcm2p1f_ca_w_0_150_s_0_315 = '-1.73750e-06*ic_cap*ic_cap+-9.50000e-07*ic_cap+1.31000e-04'
+ mcm2p1f_ca_w_0_150_s_0_420 = '-1.73750e-06*ic_cap*ic_cap+-9.50000e-07*ic_cap+1.31000e-04'
+ mcm2p1f_ca_w_0_150_s_0_525 = '-1.73750e-06*ic_cap*ic_cap+-9.50000e-07*ic_cap+1.31000e-04'
+ mcm2p1f_ca_w_0_150_s_0_630 = '-1.73750e-06*ic_cap*ic_cap+-9.50000e-07*ic_cap+1.31000e-04'
+ mcm2p1f_ca_w_0_150_s_0_840 = '-1.73750e-06*ic_cap*ic_cap+-9.50000e-07*ic_cap+1.31000e-04'
+ mcm2p1f_ca_w_0_150_s_1_260 = '-1.73750e-06*ic_cap*ic_cap+-9.50000e-07*ic_cap+1.31000e-04'
+ mcm2p1f_ca_w_0_150_s_2_310 = '-1.73750e-06*ic_cap*ic_cap+-9.50000e-07*ic_cap+1.31000e-04'
+ mcm2p1f_ca_w_0_150_s_5_250 = '-1.73750e-06*ic_cap*ic_cap+-9.50000e-07*ic_cap+1.31000e-04'
+ mcm2p1f_ca_w_1_200_s_0_210 = '-1.73750e-06*ic_cap*ic_cap+-9.50000e-07*ic_cap+1.31000e-04'
+ mcm2p1f_ca_w_1_200_s_0_263 = '-1.73750e-06*ic_cap*ic_cap+-9.50000e-07*ic_cap+1.31000e-04'
+ mcm2p1f_ca_w_1_200_s_0_315 = '-1.73750e-06*ic_cap*ic_cap+-9.50000e-07*ic_cap+1.31000e-04'
+ mcm2p1f_ca_w_1_200_s_0_420 = '-1.73750e-06*ic_cap*ic_cap+-9.50000e-07*ic_cap+1.31000e-04'
+ mcm2p1f_ca_w_1_200_s_0_525 = '-1.73750e-06*ic_cap*ic_cap+-9.50000e-07*ic_cap+1.31000e-04'
+ mcm2p1f_ca_w_1_200_s_0_630 = '-1.73750e-06*ic_cap*ic_cap+-9.50000e-07*ic_cap+1.31000e-04'
+ mcm2p1f_ca_w_1_200_s_0_840 = '-1.73750e-06*ic_cap*ic_cap+-9.50000e-07*ic_cap+1.31000e-04'
+ mcm2p1f_ca_w_1_200_s_1_260 = '-1.73750e-06*ic_cap*ic_cap+-9.50000e-07*ic_cap+1.31000e-04'
+ mcm2p1f_ca_w_1_200_s_2_310 = '-1.73750e-06*ic_cap*ic_cap+-9.50000e-07*ic_cap+1.31000e-04'
+ mcm2p1f_ca_w_1_200_s_5_250 = '-1.73750e-06*ic_cap*ic_cap+-9.50000e-07*ic_cap+1.31000e-04'
+ mcm2p1f_cc_w_0_150_s_0_210 = '-5.18750e-13*ic_cap*ic_cap+-3.00000e-13*ic_cap+7.25000e-11'
+ mcm2p1f_cc_w_0_150_s_0_263 = '-3.28125e-13*ic_cap*ic_cap+-1.87500e-13*ic_cap+5.80000e-11'
+ mcm2p1f_cc_w_0_150_s_0_315 = '-2.00000e-13*ic_cap*ic_cap+-1.25000e-13*ic_cap+4.81000e-11'
+ mcm2p1f_cc_w_0_150_s_0_420 = '-8.12500e-14*ic_cap*ic_cap+-5.00000e-14*ic_cap+3.53000e-11'
+ mcm2p1f_cc_w_0_150_s_0_525 = '-1.56250e-14*ic_cap*ic_cap+-1.25000e-14*ic_cap+2.71000e-11'
+ mcm2p1f_cc_w_0_150_s_0_630 = '2.50000e-14*ic_cap*ic_cap+2.50000e-14*ic_cap+2.13000e-11'
+ mcm2p1f_cc_w_0_150_s_0_840 = '5.93750e-14*ic_cap*ic_cap+3.75000e-14*ic_cap+1.37000e-11'
+ mcm2p1f_cc_w_0_150_s_1_260 = '5.96875e-14*ic_cap*ic_cap+4.12500e-14*ic_cap+6.29000e-12'
+ mcm2p1f_cc_w_0_150_s_2_310 = '3.21875e-14*ic_cap*ic_cap+1.87500e-14*ic_cap+1.12000e-12'
+ mcm2p1f_cc_w_0_150_s_5_250 = '7.81250e-16*ic_cap*ic_cap+4.37500e-15*ic_cap+5.00000e-14'
+ mcm2p1f_cc_w_1_200_s_0_210 = '-4.31250e-13*ic_cap*ic_cap+-2.25000e-13*ic_cap+8.17000e-11'
+ mcm2p1f_cc_w_1_200_s_0_263 = '-2.37500e-13*ic_cap*ic_cap+-1.25000e-13*ic_cap+6.59000e-11'
+ mcm2p1f_cc_w_1_200_s_0_315 = '-1.21875e-13*ic_cap*ic_cap+-6.25000e-14*ic_cap+5.52000e-11'
+ mcm2p1f_cc_w_1_200_s_0_525 = '5.62500e-14*ic_cap*ic_cap+2.50000e-14*ic_cap+3.20000e-11'
+ mcm2p1f_cc_w_1_200_s_0_630 = '8.43750e-14*ic_cap*ic_cap+6.25000e-14*ic_cap+2.56000e-11'
+ mcm2p1f_cc_w_1_200_s_0_840 = '1.15625e-13*ic_cap*ic_cap+6.25000e-14*ic_cap+1.70000e-11'
+ mcm2p1f_cc_w_1_200_s_1_260 = '1.08437e-13*ic_cap*ic_cap+6.37500e-14*ic_cap+8.21000e-12'
+ mcm2p1f_cc_w_1_200_s_2_310 = '5.25000e-14*ic_cap*ic_cap+4.00000e-14*ic_cap+1.59000e-12'
+ mcm2p1f_cc_w_1_200_s_5_250 = '4.21875e-15*ic_cap*ic_cap+3.12500e-15*ic_cap+3.50000e-14'
+ mcm2p1f_cf_w_0_150_s_0_210 = '-1.09375e-13*ic_cap*ic_cap+-6.25000e-14*ic_cap+1.28000e-11'
+ mcm2p1f_cf_w_0_150_s_0_263 = '-1.46875e-13*ic_cap*ic_cap+-8.75000e-14*ic_cap+1.56000e-11'
+ mcm2p1f_cf_w_0_150_s_0_315 = '-1.75000e-13*ic_cap*ic_cap+-1.00000e-13*ic_cap+1.82000e-11'
+ mcm2p1f_cf_w_0_150_s_0_420 = '-2.28125e-13*ic_cap*ic_cap+-1.37500e-13*ic_cap+2.30000e-11'
+ mcm2p1f_cf_w_0_150_s_0_525 = '-2.71875e-13*ic_cap*ic_cap+-1.62500e-13*ic_cap+2.71000e-11'
+ mcm2p1f_cf_w_0_150_s_0_630 = '-3.00000e-13*ic_cap*ic_cap+-1.75000e-13*ic_cap+3.05000e-11'
+ mcm2p1f_cf_w_0_150_s_0_840 = '-3.31250e-13*ic_cap*ic_cap+-2.00000e-13*ic_cap+3.58000e-11'
+ mcm2p1f_cf_w_0_150_s_1_260 = '-3.46875e-13*ic_cap*ic_cap+-2.12500e-13*ic_cap+4.20000e-11'
+ mcm2p1f_cf_w_0_150_s_2_310 = '-3.21875e-13*ic_cap*ic_cap+-1.87500e-13*ic_cap+4.67000e-11'
+ mcm2p1f_cf_w_0_150_s_5_250 = '-2.93750e-13*ic_cap*ic_cap+-1.75000e-13*ic_cap+4.78000e-11'
+ mcm2p1f_cf_w_1_200_s_0_210 = '-1.09375e-13*ic_cap*ic_cap+-6.25000e-14*ic_cap+1.27000e-11'
+ mcm2p1f_cf_w_1_200_s_0_263 = '-1.43750e-13*ic_cap*ic_cap+-7.50000e-14*ic_cap+1.56000e-11'
+ mcm2p1f_cf_w_1_200_s_0_315 = '-1.75000e-13*ic_cap*ic_cap+-1.00000e-13*ic_cap+1.82000e-11'
+ mcm2p1f_cf_w_1_200_s_0_420 = '-2.25000e-13*ic_cap*ic_cap+-1.25000e-13*ic_cap+2.30000e-11'
+ mcm2p1f_cf_w_1_200_s_0_525 = '-2.62500e-13*ic_cap*ic_cap+-1.50000e-13*ic_cap+2.72000e-11'
+ mcm2p1f_cf_w_1_200_s_0_630 = '-2.93750e-13*ic_cap*ic_cap+-1.75000e-13*ic_cap+3.08000e-11'
+ mcm2p1f_cf_w_1_200_s_0_840 = '-3.28125e-13*ic_cap*ic_cap+-1.87500e-13*ic_cap+3.65000e-11'
+ mcm2p1f_cf_w_1_200_s_1_260 = '-3.43750e-13*ic_cap*ic_cap+-2.00000e-13*ic_cap+4.36000e-11'
+ mcm2p1f_cf_w_1_200_s_2_310 = '-3.03125e-13*ic_cap*ic_cap+-1.87500e-13*ic_cap+4.97000e-11'
+ mcm2p1f_cf_w_1_200_s_5_250 = '-2.56250e-13*ic_cap*ic_cap+-1.50000e-13*ic_cap+5.12000e-11'
+ mcm3d_ca_w_0_300_s_0_300 = '-1.37500e-07*ic_cap*ic_cap+-7.50000e-08*ic_cap+1.42000e-05'
+ mcm3d_ca_w_0_300_s_0_360 = '-1.37500e-07*ic_cap*ic_cap+-7.50000e-08*ic_cap+1.42000e-05'
+ mcm3d_ca_w_0_300_s_0_450 = '-1.37500e-07*ic_cap*ic_cap+-7.50000e-08*ic_cap+1.42000e-05'
+ mcm3d_ca_w_0_300_s_0_600 = '-1.37500e-07*ic_cap*ic_cap+-7.50000e-08*ic_cap+1.42000e-05'
+ mcm3d_ca_w_0_300_s_0_800 = '-1.37500e-07*ic_cap*ic_cap+-7.50000e-08*ic_cap+1.42000e-05'
+ mcm3d_ca_w_0_300_s_1_000 = '-1.37500e-07*ic_cap*ic_cap+-7.50000e-08*ic_cap+1.42000e-05'
+ mcm3d_ca_w_0_300_s_1_200 = '-1.37500e-07*ic_cap*ic_cap+-7.50000e-08*ic_cap+1.42000e-05'
+ mcm3d_ca_w_0_300_s_2_100 = '-1.37500e-07*ic_cap*ic_cap+-7.50000e-08*ic_cap+1.42000e-05'
+ mcm3d_ca_w_0_300_s_3_300 = '-1.37500e-07*ic_cap*ic_cap+-7.50000e-08*ic_cap+1.42000e-05'
+ mcm3d_ca_w_0_300_s_9_000 = '-1.37500e-07*ic_cap*ic_cap+-7.50000e-08*ic_cap+1.42000e-05'
+ mcm3d_ca_w_2_400_s_0_300 = '-1.37500e-07*ic_cap*ic_cap+-7.50000e-08*ic_cap+1.42000e-05'
+ mcm3d_ca_w_2_400_s_0_360 = '-1.37500e-07*ic_cap*ic_cap+-7.50000e-08*ic_cap+1.42000e-05'
+ mcm3d_ca_w_2_400_s_0_450 = '-1.37500e-07*ic_cap*ic_cap+-7.50000e-08*ic_cap+1.42000e-05'
+ mcm3d_ca_w_2_400_s_0_600 = '-1.37500e-07*ic_cap*ic_cap+-7.50000e-08*ic_cap+1.42000e-05'
+ mcm3d_ca_w_2_400_s_0_800 = '-1.37500e-07*ic_cap*ic_cap+-7.50000e-08*ic_cap+1.42000e-05'
+ mcm3d_ca_w_2_400_s_1_000 = '-1.37500e-07*ic_cap*ic_cap+-7.50000e-08*ic_cap+1.42000e-05'
+ mcm3d_ca_w_2_400_s_1_200 = '-1.37500e-07*ic_cap*ic_cap+-7.50000e-08*ic_cap+1.42000e-05'
+ mcm3d_ca_w_2_400_s_2_100 = '-1.37500e-07*ic_cap*ic_cap+-7.50000e-08*ic_cap+1.42000e-05'
+ mcm3d_ca_w_2_400_s_3_300 = '-1.37500e-07*ic_cap*ic_cap+-7.50000e-08*ic_cap+1.42000e-05'
+ mcm3d_ca_w_2_400_s_9_000 = '-1.37500e-07*ic_cap*ic_cap+-7.50000e-08*ic_cap+1.42000e-05'
+ mcm3d_cc_w_0_300_s_0_300 = '-7.90625e-13*ic_cap*ic_cap+-4.62500e-13*ic_cap+1.06000e-10'
+ mcm3d_cc_w_0_300_s_0_360 = '-6.93750e-13*ic_cap*ic_cap+-4.00000e-13*ic_cap+9.90000e-11'
+ mcm3d_cc_w_0_300_s_0_450 = '-5.75000e-13*ic_cap*ic_cap+-3.50000e-13*ic_cap+8.93000e-11'
+ mcm3d_cc_w_0_300_s_0_600 = '-4.43750e-13*ic_cap*ic_cap+-2.75000e-13*ic_cap+7.68000e-11'
+ mcm3d_cc_w_0_300_s_0_800 = '-3.06250e-13*ic_cap*ic_cap+-2.25000e-13*ic_cap+6.46000e-11'
+ mcm3d_cc_w_0_300_s_1_000 = '-2.21875e-13*ic_cap*ic_cap+-1.62500e-13*ic_cap+5.55000e-11'
+ mcm3d_cc_w_0_300_s_1_200 = '-1.65625e-13*ic_cap*ic_cap+-1.12500e-13*ic_cap+4.86000e-11'
+ mcm3d_cc_w_0_300_s_2_100 = '-5.31250e-14*ic_cap*ic_cap+-3.75000e-14*ic_cap+3.16000e-11'
+ mcm3d_cc_w_0_300_s_3_300 = '-6.25000e-15*ic_cap*ic_cap+2.16000e-11'
+ mcm3d_cc_w_0_300_s_9_000 = '2.59375e-14*ic_cap*ic_cap+1.87500e-14*ic_cap+6.17000e-12'
+ mcm3d_cc_w_2_400_s_0_300 = '-7.18750e-13*ic_cap*ic_cap+-3.75000e-13*ic_cap+1.30000e-10'
+ mcm3d_cc_w_2_400_s_0_360 = '-6.25000e-13*ic_cap*ic_cap+-2.50000e-13*ic_cap+1.22000e-10'
+ mcm3d_cc_w_2_400_s_0_450 = '-5.00000e-13*ic_cap*ic_cap+-2.50000e-13*ic_cap+1.11000e-10'
+ mcm3d_cc_w_2_400_s_0_600 = '-3.68750e-13*ic_cap*ic_cap+-2.00000e-13*ic_cap+9.60000e-11'
+ mcm3d_cc_w_2_400_s_0_800 = '-2.43750e-13*ic_cap*ic_cap+-1.50000e-13*ic_cap+8.14000e-11'
+ mcm3d_cc_w_2_400_s_1_000 = '-1.65625e-13*ic_cap*ic_cap+-1.12500e-13*ic_cap+7.06000e-11'
+ mcm3d_cc_w_2_400_s_1_200 = '-1.12500e-13*ic_cap*ic_cap+-7.50000e-14*ic_cap+6.25000e-11'
+ mcm3d_cc_w_2_400_s_2_100 = '-1.56250e-14*ic_cap*ic_cap+-1.25000e-14*ic_cap+4.22000e-11'
+ mcm3d_cc_w_2_400_s_3_300 = '2.18750e-14*ic_cap*ic_cap+1.25000e-14*ic_cap+2.95000e-11'
+ mcm3d_cc_w_2_400_s_9_000 = '3.56250e-14*ic_cap*ic_cap+2.50000e-14*ic_cap+9.73000e-12'
+ mcm3d_cf_w_0_300_s_0_300 = '-5.31250e-15*ic_cap*ic_cap+-3.75000e-15*ic_cap+2.09000e-12'
+ mcm3d_cf_w_0_300_s_0_360 = '-9.06250e-15*ic_cap*ic_cap+-6.25000e-15*ic_cap+2.50000e-12'
+ mcm3d_cf_w_0_300_s_0_450 = '-1.46875e-14*ic_cap*ic_cap+-8.75000e-15*ic_cap+3.13000e-12'
+ mcm3d_cf_w_0_300_s_0_600 = '-2.34375e-14*ic_cap*ic_cap+-1.62500e-14*ic_cap+4.15000e-12'
+ mcm3d_cf_w_0_300_s_0_800 = '-3.65625e-14*ic_cap*ic_cap+-2.37500e-14*ic_cap+5.39000e-12'
+ mcm3d_cf_w_0_300_s_1_000 = '-4.78125e-14*ic_cap*ic_cap+-3.12500e-14*ic_cap+6.64000e-12'
+ mcm3d_cf_w_0_300_s_1_200 = '-5.81250e-14*ic_cap*ic_cap+-3.75000e-14*ic_cap+7.84000e-12'
+ mcm3d_cf_w_0_300_s_2_100 = '-1.03125e-13*ic_cap*ic_cap+-6.25000e-14*ic_cap+1.31000e-11'
+ mcm3d_cf_w_0_300_s_3_300 = '-1.34375e-13*ic_cap*ic_cap+-8.75000e-14*ic_cap+1.80000e-11'
+ mcm3d_cf_w_0_300_s_9_000 = '-1.78125e-13*ic_cap*ic_cap+-1.12500e-13*ic_cap+2.99000e-11'
+ mcm3d_cf_w_2_400_s_0_300 = '-6.25000e-15*ic_cap*ic_cap+-5.00000e-15*ic_cap+2.14000e-12'
+ mcm3d_cf_w_2_400_s_0_360 = '-1.00000e-14*ic_cap*ic_cap+-7.50000e-15*ic_cap+2.55000e-12'
+ mcm3d_cf_w_2_400_s_0_450 = '-1.59375e-14*ic_cap*ic_cap+-1.12500e-14*ic_cap+3.16000e-12'
+ mcm3d_cf_w_2_400_s_0_600 = '-2.46875e-14*ic_cap*ic_cap+-1.62500e-14*ic_cap+4.15000e-12'
+ mcm3d_cf_w_2_400_s_0_800 = '-3.68750e-14*ic_cap*ic_cap+-2.50000e-14*ic_cap+5.45000e-12'
+ mcm3d_cf_w_2_400_s_1_000 = '-4.84375e-14*ic_cap*ic_cap+-3.12500e-14*ic_cap+6.72000e-12'
+ mcm3d_cf_w_2_400_s_1_200 = '-5.84375e-14*ic_cap*ic_cap+-3.87500e-14*ic_cap+7.94000e-12'
+ mcm3d_cf_w_2_400_s_2_100 = '-1.00000e-13*ic_cap*ic_cap+-7.50000e-14*ic_cap+1.30000e-11'
+ mcm3d_cf_w_2_400_s_3_300 = '-1.40625e-13*ic_cap*ic_cap+-8.75000e-14*ic_cap+1.86000e-11'
+ mcm3d_cf_w_2_400_s_9_000 = '-1.81250e-13*ic_cap*ic_cap+-1.25000e-13*ic_cap+3.28000e-11'
+ mcm3f_ca_w_0_300_s_0_300 = '-1.31250e-07*ic_cap*ic_cap+-7.50000e-08*ic_cap+1.26000e-05'
+ mcm3f_ca_w_0_300_s_0_360 = '-1.31250e-07*ic_cap*ic_cap+-7.50000e-08*ic_cap+1.26000e-05'
+ mcm3f_ca_w_0_300_s_0_450 = '-1.31250e-07*ic_cap*ic_cap+-7.50000e-08*ic_cap+1.26000e-05'
+ mcm3f_ca_w_0_300_s_0_600 = '-1.31250e-07*ic_cap*ic_cap+-7.50000e-08*ic_cap+1.26000e-05'
+ mcm3f_ca_w_0_300_s_0_800 = '-1.31250e-07*ic_cap*ic_cap+-7.50000e-08*ic_cap+1.26000e-05'
+ mcm3f_ca_w_0_300_s_1_000 = '-1.31250e-07*ic_cap*ic_cap+-7.50000e-08*ic_cap+1.26000e-05'
+ mcm3f_ca_w_0_300_s_1_200 = '-1.31250e-07*ic_cap*ic_cap+-7.50000e-08*ic_cap+1.26000e-05'
+ mcm3f_ca_w_0_300_s_2_100 = '-1.31250e-07*ic_cap*ic_cap+-7.50000e-08*ic_cap+1.26000e-05'
+ mcm3f_ca_w_0_300_s_3_300 = '-1.31250e-07*ic_cap*ic_cap+-7.50000e-08*ic_cap+1.26000e-05'
+ mcm3f_ca_w_0_300_s_9_000 = '-1.31250e-07*ic_cap*ic_cap+-7.50000e-08*ic_cap+1.26000e-05'
+ mcm3f_ca_w_2_400_s_0_300 = '-1.31250e-07*ic_cap*ic_cap+-7.50000e-08*ic_cap+1.26000e-05'
+ mcm3f_ca_w_2_400_s_0_360 = '-1.31250e-07*ic_cap*ic_cap+-7.50000e-08*ic_cap+1.26000e-05'
+ mcm3f_ca_w_2_400_s_0_450 = '-1.31250e-07*ic_cap*ic_cap+-7.50000e-08*ic_cap+1.26000e-05'
+ mcm3f_ca_w_2_400_s_0_600 = '-1.31250e-07*ic_cap*ic_cap+-7.50000e-08*ic_cap+1.26000e-05'
+ mcm3f_ca_w_2_400_s_0_800 = '-1.31250e-07*ic_cap*ic_cap+-7.50000e-08*ic_cap+1.26000e-05'
+ mcm3f_ca_w_2_400_s_1_000 = '-1.31250e-07*ic_cap*ic_cap+-7.50000e-08*ic_cap+1.26000e-05'
+ mcm3f_ca_w_2_400_s_1_200 = '-1.31250e-07*ic_cap*ic_cap+-7.50000e-08*ic_cap+1.26000e-05'
+ mcm3f_ca_w_2_400_s_2_100 = '-1.31250e-07*ic_cap*ic_cap+-7.50000e-08*ic_cap+1.26000e-05'
+ mcm3f_ca_w_2_400_s_3_300 = '-1.31250e-07*ic_cap*ic_cap+-7.50000e-08*ic_cap+1.26000e-05'
+ mcm3f_ca_w_2_400_s_9_000 = '-1.31250e-07*ic_cap*ic_cap+-7.50000e-08*ic_cap+1.26000e-05'
+ mcm3f_cc_w_0_300_s_0_300 = '-7.62500e-13*ic_cap*ic_cap+-4.50000e-13*ic_cap+1.06000e-10'
+ mcm3f_cc_w_0_300_s_0_360 = '-7.00000e-13*ic_cap*ic_cap+-4.00000e-13*ic_cap+9.95000e-11'
+ mcm3f_cc_w_0_300_s_0_450 = '-5.81250e-13*ic_cap*ic_cap+-3.50000e-13*ic_cap+8.98000e-11'
+ mcm3f_cc_w_0_300_s_0_600 = '-4.40625e-13*ic_cap*ic_cap+-2.87500e-13*ic_cap+7.73000e-11'
+ mcm3f_cc_w_0_300_s_0_800 = '-3.12500e-13*ic_cap*ic_cap+-2.25000e-13*ic_cap+6.53000e-11'
+ mcm3f_cc_w_0_300_s_1_000 = '-2.25000e-13*ic_cap*ic_cap+-1.50000e-13*ic_cap+5.62000e-11'
+ mcm3f_cc_w_0_300_s_1_200 = '-1.68750e-13*ic_cap*ic_cap+-1.25000e-13*ic_cap+4.95000e-11'
+ mcm3f_cc_w_0_300_s_2_100 = '-5.93750e-14*ic_cap*ic_cap+-3.75000e-14*ic_cap+3.26000e-11'
+ mcm3f_cc_w_0_300_s_3_300 = '-3.12500e-15*ic_cap*ic_cap+-1.25000e-14*ic_cap+2.26000e-11'
+ mcm3f_cc_w_0_300_s_9_000 = '3.06250e-14*ic_cap*ic_cap+2.25000e-14*ic_cap+6.81000e-12'
+ mcm3f_cc_w_2_400_s_0_300 = '-7.50000e-13*ic_cap*ic_cap+-5.00000e-13*ic_cap+1.32000e-10'
+ mcm3f_cc_w_2_400_s_0_360 = '-6.25000e-13*ic_cap*ic_cap+-2.50000e-13*ic_cap+1.23000e-10'
+ mcm3f_cc_w_2_400_s_0_450 = '-5.00000e-13*ic_cap*ic_cap+-2.50000e-13*ic_cap+1.12000e-10'
+ mcm3f_cc_w_2_400_s_0_600 = '-3.65625e-13*ic_cap*ic_cap+-2.12500e-13*ic_cap+9.72000e-11'
+ mcm3f_cc_w_2_400_s_0_800 = '-2.43750e-13*ic_cap*ic_cap+-1.50000e-13*ic_cap+8.27000e-11'
+ mcm3f_cc_w_2_400_s_1_000 = '-1.68750e-13*ic_cap*ic_cap+-1.25000e-13*ic_cap+7.19000e-11'
+ mcm3f_cc_w_2_400_s_1_200 = '-1.15625e-13*ic_cap*ic_cap+-8.75000e-14*ic_cap+6.38000e-11'
+ mcm3f_cc_w_2_400_s_2_100 = '-1.56250e-14*ic_cap*ic_cap+-1.25000e-14*ic_cap+4.35000e-11'
+ mcm3f_cc_w_2_400_s_3_300 = '3.12500e-14*ic_cap*ic_cap+2.50000e-14*ic_cap+3.06000e-11'
+ mcm3f_cc_w_2_400_s_9_000 = '4.68750e-14*ic_cap*ic_cap+3.75000e-14*ic_cap+1.05000e-11'
+ mcm3f_cf_w_0_300_s_0_300 = '-5.93750e-15*ic_cap*ic_cap+-3.75000e-15*ic_cap+1.86000e-12'
+ mcm3f_cf_w_0_300_s_0_360 = '-9.06250e-15*ic_cap*ic_cap+-6.25000e-15*ic_cap+2.22000e-12'
+ mcm3f_cf_w_0_300_s_0_450 = '-1.46875e-14*ic_cap*ic_cap+-8.75000e-15*ic_cap+2.79000e-12'
+ mcm3f_cf_w_0_300_s_0_600 = '-2.31250e-14*ic_cap*ic_cap+-1.50000e-14*ic_cap+3.70000e-12'
+ mcm3f_cf_w_0_300_s_0_800 = '-3.50000e-14*ic_cap*ic_cap+-2.25000e-14*ic_cap+4.80000e-12'
+ mcm3f_cf_w_0_300_s_1_000 = '-4.59375e-14*ic_cap*ic_cap+-2.87500e-14*ic_cap+5.93000e-12'
+ mcm3f_cf_w_0_300_s_1_200 = '-5.56250e-14*ic_cap*ic_cap+-3.50000e-14*ic_cap+7.00000e-12'
+ mcm3f_cf_w_0_300_s_2_100 = '-9.68750e-14*ic_cap*ic_cap+-6.25000e-14*ic_cap+1.18000e-11'
+ mcm3f_cf_w_0_300_s_3_300 = '-1.34375e-13*ic_cap*ic_cap+-8.75000e-14*ic_cap+1.64000e-11'
+ mcm3f_cf_w_0_300_s_9_000 = '-1.81250e-13*ic_cap*ic_cap+-1.25000e-13*ic_cap+2.82000e-11'
+ mcm3f_cf_w_2_400_s_0_300 = '-5.93750e-15*ic_cap*ic_cap+-3.75000e-15*ic_cap+1.89000e-12'
+ mcm3f_cf_w_2_400_s_0_360 = '-1.00000e-14*ic_cap*ic_cap+-7.50000e-15*ic_cap+2.26000e-12'
+ mcm3f_cf_w_2_400_s_0_450 = '-1.50000e-14*ic_cap*ic_cap+-1.00000e-14*ic_cap+2.80000e-12'
+ mcm3f_cf_w_2_400_s_0_600 = '-2.37500e-14*ic_cap*ic_cap+-1.50000e-14*ic_cap+3.69000e-12'
+ mcm3f_cf_w_2_400_s_0_800 = '-3.56250e-14*ic_cap*ic_cap+-2.25000e-14*ic_cap+4.86000e-12'
+ mcm3f_cf_w_2_400_s_1_000 = '-4.65625e-14*ic_cap*ic_cap+-2.87500e-14*ic_cap+6.00000e-12'
+ mcm3f_cf_w_2_400_s_1_200 = '-5.71875e-14*ic_cap*ic_cap+-3.62500e-14*ic_cap+7.11000e-12'
+ mcm3f_cf_w_2_400_s_2_100 = '-9.65625e-14*ic_cap*ic_cap+-6.12500e-14*ic_cap+1.17000e-11'
+ mcm3f_cf_w_2_400_s_3_300 = '-1.34375e-13*ic_cap*ic_cap+-8.75000e-14*ic_cap+1.69000e-11'
+ mcm3f_cf_w_2_400_s_9_000 = '-1.87500e-13*ic_cap*ic_cap+-1.25000e-13*ic_cap+3.09000e-11'
+ mcm3l1_ca_w_0_300_s_0_300 = '-2.09375e-07*ic_cap*ic_cap+-1.37500e-07*ic_cap+2.02000e-05'
+ mcm3l1_ca_w_0_300_s_0_360 = '-2.09375e-07*ic_cap*ic_cap+-1.37500e-07*ic_cap+2.02000e-05'
+ mcm3l1_ca_w_0_300_s_0_450 = '-2.09375e-07*ic_cap*ic_cap+-1.37500e-07*ic_cap+2.02000e-05'
+ mcm3l1_ca_w_0_300_s_0_600 = '-2.09375e-07*ic_cap*ic_cap+-1.37500e-07*ic_cap+2.02000e-05'
+ mcm3l1_ca_w_0_300_s_0_800 = '-2.09375e-07*ic_cap*ic_cap+-1.37500e-07*ic_cap+2.02000e-05'
+ mcm3l1_ca_w_0_300_s_1_000 = '-2.09375e-07*ic_cap*ic_cap+-1.37500e-07*ic_cap+2.02000e-05'
+ mcm3l1_ca_w_0_300_s_1_200 = '-2.09375e-07*ic_cap*ic_cap+-1.37500e-07*ic_cap+2.02000e-05'
+ mcm3l1_ca_w_0_300_s_2_100 = '-2.09375e-07*ic_cap*ic_cap+-1.37500e-07*ic_cap+2.02000e-05'
+ mcm3l1_ca_w_0_300_s_3_300 = '-2.09375e-07*ic_cap*ic_cap+-1.37500e-07*ic_cap+2.02000e-05'
+ mcm3l1_ca_w_0_300_s_9_000 = '-2.09375e-07*ic_cap*ic_cap+-1.37500e-07*ic_cap+2.02000e-05'
+ mcm3l1_ca_w_2_400_s_0_300 = '-2.09375e-07*ic_cap*ic_cap+-1.37500e-07*ic_cap+2.02000e-05'
+ mcm3l1_ca_w_2_400_s_0_360 = '-2.09375e-07*ic_cap*ic_cap+-1.37500e-07*ic_cap+2.02000e-05'
+ mcm3l1_ca_w_2_400_s_0_450 = '-2.09375e-07*ic_cap*ic_cap+-1.37500e-07*ic_cap+2.02000e-05'
+ mcm3l1_ca_w_2_400_s_0_600 = '-2.09375e-07*ic_cap*ic_cap+-1.37500e-07*ic_cap+2.02000e-05'
+ mcm3l1_ca_w_2_400_s_0_800 = '-2.09375e-07*ic_cap*ic_cap+-1.37500e-07*ic_cap+2.02000e-05'
+ mcm3l1_ca_w_2_400_s_1_000 = '-2.09375e-07*ic_cap*ic_cap+-1.37500e-07*ic_cap+2.02000e-05'
+ mcm3l1_ca_w_2_400_s_1_200 = '-2.09375e-07*ic_cap*ic_cap+-1.37500e-07*ic_cap+2.02000e-05'
+ mcm3l1_ca_w_2_400_s_2_100 = '-2.09375e-07*ic_cap*ic_cap+-1.37500e-07*ic_cap+2.02000e-05'
+ mcm3l1_ca_w_2_400_s_3_300 = '-2.09375e-07*ic_cap*ic_cap+-1.37500e-07*ic_cap+2.02000e-05'
+ mcm3l1_ca_w_2_400_s_9_000 = '-2.09375e-07*ic_cap*ic_cap+-1.37500e-07*ic_cap+2.02000e-05'
+ mcm3l1_cc_w_0_300_s_0_300 = '-8.03125e-13*ic_cap*ic_cap+-4.62500e-13*ic_cap+1.05000e-10'
+ mcm3l1_cc_w_0_300_s_0_360 = '-6.71875e-13*ic_cap*ic_cap+-4.12500e-13*ic_cap+9.73000e-11'
+ mcm3l1_cc_w_0_300_s_0_450 = '-5.53125e-13*ic_cap*ic_cap+-3.37500e-13*ic_cap+8.75000e-11'
+ mcm3l1_cc_w_0_300_s_0_600 = '-4.25000e-13*ic_cap*ic_cap+-2.75000e-13*ic_cap+7.49000e-11'
+ mcm3l1_cc_w_0_300_s_0_800 = '-2.87500e-13*ic_cap*ic_cap+-2.00000e-13*ic_cap+6.24000e-11'
+ mcm3l1_cc_w_0_300_s_1_000 = '-2.09375e-13*ic_cap*ic_cap+-1.37500e-13*ic_cap+5.32000e-11'
+ mcm3l1_cc_w_0_300_s_1_200 = '-1.53125e-13*ic_cap*ic_cap+-1.12500e-13*ic_cap+4.62000e-11'
+ mcm3l1_cc_w_0_300_s_2_100 = '-4.06250e-14*ic_cap*ic_cap+-1.25000e-14*ic_cap+2.86000e-11'
+ mcm3l1_cc_w_0_300_s_3_300 = '6.25000e-15*ic_cap*ic_cap+1.86000e-11'
+ mcm3l1_cc_w_0_300_s_9_000 = '1.96875e-14*ic_cap*ic_cap+1.62500e-14*ic_cap+4.69000e-12'
+ mcm3l1_cc_w_2_400_s_0_300 = '-7.18750e-13*ic_cap*ic_cap+-3.75000e-13*ic_cap+1.27000e-10'
+ mcm3l1_cc_w_2_400_s_0_360 = '-5.93750e-13*ic_cap*ic_cap+-3.75000e-13*ic_cap+1.18000e-10'
+ mcm3l1_cc_w_2_400_s_0_450 = '-4.90625e-13*ic_cap*ic_cap+-2.12500e-13*ic_cap+1.07000e-10'
+ mcm3l1_cc_w_2_400_s_0_600 = '-3.62500e-13*ic_cap*ic_cap+-2.00000e-13*ic_cap+9.24000e-11'
+ mcm3l1_cc_w_2_400_s_0_800 = '-2.28125e-13*ic_cap*ic_cap+-1.37500e-13*ic_cap+7.77000e-11'
+ mcm3l1_cc_w_2_400_s_1_000 = '-1.50000e-13*ic_cap*ic_cap+-1.00000e-13*ic_cap+6.68000e-11'
+ mcm3l1_cc_w_2_400_s_1_200 = '-9.68750e-14*ic_cap*ic_cap+-6.25000e-14*ic_cap+5.87000e-11'
+ mcm3l1_cc_w_2_400_s_2_100 = '-1.25000e-14*ic_cap*ic_cap+3.86000e-11'
+ mcm3l1_cc_w_2_400_s_3_300 = '3.12500e-14*ic_cap*ic_cap+2.50000e-14*ic_cap+2.60000e-11'
+ mcm3l1_cc_w_2_400_s_9_000 = '2.96875e-14*ic_cap*ic_cap+1.87500e-14*ic_cap+7.85000e-12'
+ mcm3l1_cf_w_0_300_s_0_300 = '-9.37500e-15*ic_cap*ic_cap+-7.50000e-15*ic_cap+2.95000e-12'
+ mcm3l1_cf_w_0_300_s_0_360 = '-1.53125e-14*ic_cap*ic_cap+-1.12500e-14*ic_cap+3.52000e-12'
+ mcm3l1_cf_w_0_300_s_0_450 = '-2.28125e-14*ic_cap*ic_cap+-1.62500e-14*ic_cap+4.38000e-12'
+ mcm3l1_cf_w_0_300_s_0_600 = '-3.62500e-14*ic_cap*ic_cap+-2.50000e-14*ic_cap+5.78000e-12'
+ mcm3l1_cf_w_0_300_s_0_800 = '-5.37500e-14*ic_cap*ic_cap+-3.50000e-14*ic_cap+7.48000e-12'
+ mcm3l1_cf_w_0_300_s_1_000 = '-6.90625e-14*ic_cap*ic_cap+-4.62500e-14*ic_cap+9.16000e-12'
+ mcm3l1_cf_w_0_300_s_1_200 = '-8.56250e-14*ic_cap*ic_cap+-5.50000e-14*ic_cap+1.08000e-11'
+ mcm3l1_cf_w_0_300_s_2_100 = '-1.34375e-13*ic_cap*ic_cap+-8.75000e-14*ic_cap+1.74000e-11'
+ mcm3l1_cf_w_0_300_s_3_300 = '-1.71875e-13*ic_cap*ic_cap+-1.12500e-13*ic_cap+2.32000e-11'
+ mcm3l1_cf_w_0_300_s_9_000 = '-1.96875e-13*ic_cap*ic_cap+-1.37500e-13*ic_cap+3.48000e-11'
+ mcm3l1_cf_w_2_400_s_0_300 = '-1.00000e-14*ic_cap*ic_cap+-7.50000e-15*ic_cap+2.99000e-12'
+ mcm3l1_cf_w_2_400_s_0_360 = '-1.59375e-14*ic_cap*ic_cap+-1.12500e-14*ic_cap+3.56000e-12'
+ mcm3l1_cf_w_2_400_s_0_450 = '-2.43750e-14*ic_cap*ic_cap+-1.75000e-14*ic_cap+4.41000e-12'
+ mcm3l1_cf_w_2_400_s_0_600 = '-3.75000e-14*ic_cap*ic_cap+-2.50000e-14*ic_cap+5.78000e-12'
+ mcm3l1_cf_w_2_400_s_0_800 = '-5.40625e-14*ic_cap*ic_cap+-3.62500e-14*ic_cap+7.55000e-12'
+ mcm3l1_cf_w_2_400_s_1_000 = '-6.93750e-14*ic_cap*ic_cap+-4.75000e-14*ic_cap+9.25000e-12'
+ mcm3l1_cf_w_2_400_s_1_200 = '-8.53125e-14*ic_cap*ic_cap+-5.62500e-14*ic_cap+1.09000e-11'
+ mcm3l1_cf_w_2_400_s_2_100 = '-1.31250e-13*ic_cap*ic_cap+-1.00000e-13*ic_cap+1.73000e-11'
+ mcm3l1_cf_w_2_400_s_3_300 = '-1.71875e-13*ic_cap*ic_cap+-1.12500e-13*ic_cap+2.40000e-11'
+ mcm3l1_cf_w_2_400_s_9_000 = '-2.00000e-13*ic_cap*ic_cap+-1.50000e-13*ic_cap+3.84000e-11'
+ mcm3l1d_ca_w_0_170_s_0_180 = '-7.53125e-07*ic_cap*ic_cap+-4.37500e-07*ic_cap+7.54000e-05'
+ mcm3l1d_ca_w_0_170_s_0_225 = '-7.53125e-07*ic_cap*ic_cap+-4.37500e-07*ic_cap+7.54000e-05'
+ mcm3l1d_ca_w_0_170_s_0_270 = '-7.53125e-07*ic_cap*ic_cap+-4.37500e-07*ic_cap+7.54000e-05'
+ mcm3l1d_ca_w_0_170_s_0_360 = '-7.53125e-07*ic_cap*ic_cap+-4.37500e-07*ic_cap+7.54000e-05'
+ mcm3l1d_ca_w_0_170_s_0_450 = '-7.53125e-07*ic_cap*ic_cap+-4.37500e-07*ic_cap+7.54000e-05'
+ mcm3l1d_ca_w_0_170_s_0_540 = '-7.53125e-07*ic_cap*ic_cap+-4.37500e-07*ic_cap+7.54000e-05'
+ mcm3l1d_ca_w_0_170_s_0_720 = '-7.53125e-07*ic_cap*ic_cap+-4.37500e-07*ic_cap+7.54000e-05'
+ mcm3l1d_ca_w_0_170_s_1_080 = '-7.53125e-07*ic_cap*ic_cap+-4.37500e-07*ic_cap+7.54000e-05'
+ mcm3l1d_ca_w_0_170_s_1_980 = '-7.53125e-07*ic_cap*ic_cap+-4.37500e-07*ic_cap+7.54000e-05'
+ mcm3l1d_ca_w_0_170_s_4_500 = '-7.53125e-07*ic_cap*ic_cap+-4.37500e-07*ic_cap+7.54000e-05'
+ mcm3l1d_ca_w_1_360_s_0_180 = '-7.53125e-07*ic_cap*ic_cap+-4.37500e-07*ic_cap+7.54000e-05'
+ mcm3l1d_ca_w_1_360_s_0_225 = '-7.53125e-07*ic_cap*ic_cap+-4.37500e-07*ic_cap+7.54000e-05'
+ mcm3l1d_ca_w_1_360_s_0_270 = '-7.53125e-07*ic_cap*ic_cap+-4.37500e-07*ic_cap+7.54000e-05'
+ mcm3l1d_ca_w_1_360_s_0_360 = '-7.53125e-07*ic_cap*ic_cap+-4.37500e-07*ic_cap+7.54000e-05'
+ mcm3l1d_ca_w_1_360_s_0_450 = '-7.53125e-07*ic_cap*ic_cap+-4.37500e-07*ic_cap+7.54000e-05'
+ mcm3l1d_ca_w_1_360_s_0_540 = '-7.53125e-07*ic_cap*ic_cap+-4.37500e-07*ic_cap+7.54000e-05'
+ mcm3l1d_ca_w_1_360_s_0_720 = '-7.53125e-07*ic_cap*ic_cap+-4.37500e-07*ic_cap+7.54000e-05'
+ mcm3l1d_ca_w_1_360_s_1_080 = '-7.53125e-07*ic_cap*ic_cap+-4.37500e-07*ic_cap+7.54000e-05'
+ mcm3l1d_ca_w_1_360_s_1_980 = '-7.53125e-07*ic_cap*ic_cap+-4.37500e-07*ic_cap+7.54000e-05'
+ mcm3l1d_ca_w_1_360_s_4_500 = '-7.53125e-07*ic_cap*ic_cap+-4.37500e-07*ic_cap+7.54000e-05'
+ mcm3l1d_cc_w_0_170_s_0_180 = '-7.53125e-13*ic_cap*ic_cap+-4.87500e-13*ic_cap+7.47000e-11'
+ mcm3l1d_cc_w_0_170_s_0_225 = '-5.31250e-13*ic_cap*ic_cap+-3.75000e-13*ic_cap+6.26000e-11'
+ mcm3l1d_cc_w_0_170_s_0_270 = '-3.93750e-13*ic_cap*ic_cap+-2.75000e-13*ic_cap+5.43000e-11'
+ mcm3l1d_cc_w_0_170_s_0_360 = '-2.40625e-13*ic_cap*ic_cap+-1.87500e-13*ic_cap+4.25000e-11'
+ mcm3l1d_cc_w_0_170_s_0_450 = '-1.46875e-13*ic_cap*ic_cap+-1.12500e-13*ic_cap+3.49000e-11'
+ mcm3l1d_cc_w_0_170_s_0_540 = '-9.06250e-14*ic_cap*ic_cap+-8.75000e-14*ic_cap+2.90000e-11'
+ mcm3l1d_cc_w_0_170_s_0_720 = '-2.18750e-14*ic_cap*ic_cap+-3.75000e-14*ic_cap+2.10000e-11'
+ mcm3l1d_cc_w_0_170_s_1_080 = '3.12500e-14*ic_cap*ic_cap+1.19000e-11'
+ mcm3l1d_cc_w_0_170_s_1_980 = '4.37500e-14*ic_cap*ic_cap+2.50000e-14*ic_cap+3.34000e-12'
+ mcm3l1d_cc_w_0_170_s_4_500 = '7.18750e-15*ic_cap*ic_cap+5.00000e-15*ic_cap+1.60000e-13'
+ mcm3l1d_cc_w_1_360_s_0_180 = '-6.12500e-13*ic_cap*ic_cap+-4.00000e-13*ic_cap+8.58000e-11'
+ mcm3l1d_cc_w_1_360_s_0_225 = '-3.87500e-13*ic_cap*ic_cap+-2.75000e-13*ic_cap+7.25000e-11'
+ mcm3l1d_cc_w_1_360_s_0_270 = '-2.65625e-13*ic_cap*ic_cap+-1.87500e-13*ic_cap+6.31000e-11'
+ mcm3l1d_cc_w_1_360_s_0_360 = '-1.21875e-13*ic_cap*ic_cap+-1.12500e-13*ic_cap+5.01000e-11'
+ mcm3l1d_cc_w_1_360_s_0_450 = '-3.75000e-14*ic_cap*ic_cap+-5.00000e-14*ic_cap+4.12000e-11'
+ mcm3l1d_cc_w_1_360_s_0_540 = '1.56250e-14*ic_cap*ic_cap+-1.25000e-14*ic_cap+3.46000e-11'
+ mcm3l1d_cc_w_1_360_s_0_720 = '6.25000e-14*ic_cap*ic_cap+2.50000e-14*ic_cap+2.55000e-11'
+ mcm3l1d_cc_w_1_360_s_1_080 = '1.06250e-13*ic_cap*ic_cap+5.00000e-14*ic_cap+1.48000e-11'
+ mcm3l1d_cc_w_1_360_s_1_980 = '8.00000e-14*ic_cap*ic_cap+5.25000e-14*ic_cap+4.42000e-12'
+ mcm3l1d_cc_w_1_360_s_4_500 = '1.29687e-14*ic_cap*ic_cap+1.31250e-14*ic_cap+1.80000e-13'
+ mcm3l1d_cf_w_0_170_s_0_180 = '-1.21875e-14*ic_cap*ic_cap+-6.25000e-15*ic_cap+6.60000e-12'
+ mcm3l1d_cf_w_0_170_s_0_225 = '-2.81250e-14*ic_cap*ic_cap+-1.75000e-14*ic_cap+8.16000e-12'
+ mcm3l1d_cf_w_0_170_s_0_270 = '-4.46875e-14*ic_cap*ic_cap+-2.62500e-14*ic_cap+9.66000e-12'
+ mcm3l1d_cf_w_0_170_s_0_360 = '-7.18750e-14*ic_cap*ic_cap+-3.75000e-14*ic_cap+1.27000e-11'
+ mcm3l1d_cf_w_0_170_s_0_450 = '-1.00000e-13*ic_cap*ic_cap+-5.00000e-14*ic_cap+1.52000e-11'
+ mcm3l1d_cf_w_0_170_s_0_540 = '-1.25000e-13*ic_cap*ic_cap+-7.50000e-14*ic_cap+1.78000e-11'
+ mcm3l1d_cf_w_0_170_s_0_720 = '-1.59375e-13*ic_cap*ic_cap+-8.75000e-14*ic_cap+2.20000e-11'
+ mcm3l1d_cf_w_0_170_s_1_080 = '-2.06250e-13*ic_cap*ic_cap+-1.25000e-13*ic_cap+2.82000e-11'
+ mcm3l1d_cf_w_0_170_s_1_980 = '-2.25000e-13*ic_cap*ic_cap+-1.50000e-13*ic_cap+3.54000e-11'
+ mcm3l1d_cf_w_0_170_s_4_500 = '-1.96875e-13*ic_cap*ic_cap+-1.37500e-13*ic_cap+3.85000e-11'
+ mcm3l1d_cf_w_1_360_s_0_180 = '-1.15625e-14*ic_cap*ic_cap+-6.25000e-15*ic_cap+6.57000e-12'
+ mcm3l1d_cf_w_1_360_s_0_225 = '-2.78125e-14*ic_cap*ic_cap+-1.62500e-14*ic_cap+8.14000e-12'
+ mcm3l1d_cf_w_1_360_s_0_270 = '-4.31250e-14*ic_cap*ic_cap+-2.50000e-14*ic_cap+9.67000e-12'
+ mcm3l1d_cf_w_1_360_s_0_360 = '-7.18750e-14*ic_cap*ic_cap+-3.75000e-14*ic_cap+1.26000e-11'
+ mcm3l1d_cf_w_1_360_s_0_450 = '-9.68750e-14*ic_cap*ic_cap+-6.25000e-14*ic_cap+1.53000e-11'
+ mcm3l1d_cf_w_1_360_s_0_540 = '-1.25000e-13*ic_cap*ic_cap+-7.50000e-14*ic_cap+1.79000e-11'
+ mcm3l1d_cf_w_1_360_s_0_720 = '-1.62500e-13*ic_cap*ic_cap+-1.00000e-13*ic_cap+2.24000e-11'
+ mcm3l1d_cf_w_1_360_s_1_080 = '-2.00000e-13*ic_cap*ic_cap+-1.25000e-13*ic_cap+2.92000e-11'
+ mcm3l1d_cf_w_1_360_s_1_980 = '-2.03125e-13*ic_cap*ic_cap+-1.37500e-13*ic_cap+3.78000e-11'
+ mcm3l1d_cf_w_1_360_s_4_500 = '-1.46875e-13*ic_cap*ic_cap+-8.75000e-14*ic_cap+4.19000e-11'
+ mcm3l1f_ca_w_0_170_s_0_180 = '-6.21875e-07*ic_cap*ic_cap+-3.62500e-07*ic_cap+5.71000e-05'
+ mcm3l1f_ca_w_0_170_s_0_225 = '-6.21875e-07*ic_cap*ic_cap+-3.62500e-07*ic_cap+5.71000e-05'
+ mcm3l1f_ca_w_0_170_s_0_270 = '-6.21875e-07*ic_cap*ic_cap+-3.62500e-07*ic_cap+5.71000e-05'
+ mcm3l1f_ca_w_0_170_s_0_360 = '-6.21875e-07*ic_cap*ic_cap+-3.62500e-07*ic_cap+5.71000e-05'
+ mcm3l1f_ca_w_0_170_s_0_450 = '-6.21875e-07*ic_cap*ic_cap+-3.62500e-07*ic_cap+5.71000e-05'
+ mcm3l1f_ca_w_0_170_s_0_540 = '-6.21875e-07*ic_cap*ic_cap+-3.62500e-07*ic_cap+5.71000e-05'
+ mcm3l1f_ca_w_0_170_s_0_720 = '-6.21875e-07*ic_cap*ic_cap+-3.62500e-07*ic_cap+5.71000e-05'
+ mcm3l1f_ca_w_0_170_s_1_080 = '-6.21875e-07*ic_cap*ic_cap+-3.62500e-07*ic_cap+5.71000e-05'
+ mcm3l1f_ca_w_0_170_s_1_980 = '-6.21875e-07*ic_cap*ic_cap+-3.62500e-07*ic_cap+5.71000e-05'
+ mcm3l1f_ca_w_0_170_s_4_500 = '-6.21875e-07*ic_cap*ic_cap+-3.62500e-07*ic_cap+5.71000e-05'
+ mcm3l1f_ca_w_1_360_s_0_180 = '-6.21875e-07*ic_cap*ic_cap+-3.62500e-07*ic_cap+5.71000e-05'
+ mcm3l1f_ca_w_1_360_s_0_225 = '-6.21875e-07*ic_cap*ic_cap+-3.62500e-07*ic_cap+5.71000e-05'
+ mcm3l1f_ca_w_1_360_s_0_270 = '-6.21875e-07*ic_cap*ic_cap+-3.62500e-07*ic_cap+5.71000e-05'
+ mcm3l1f_ca_w_1_360_s_0_360 = '-6.21875e-07*ic_cap*ic_cap+-3.62500e-07*ic_cap+5.71000e-05'
+ mcm3l1f_ca_w_1_360_s_0_450 = '-6.21875e-07*ic_cap*ic_cap+-3.62500e-07*ic_cap+5.71000e-05'
+ mcm3l1f_ca_w_1_360_s_0_540 = '-6.21875e-07*ic_cap*ic_cap+-3.62500e-07*ic_cap+5.71000e-05'
+ mcm3l1f_ca_w_1_360_s_0_720 = '-6.21875e-07*ic_cap*ic_cap+-3.62500e-07*ic_cap+5.71000e-05'
+ mcm3l1f_ca_w_1_360_s_1_080 = '-6.21875e-07*ic_cap*ic_cap+-3.62500e-07*ic_cap+5.71000e-05'
+ mcm3l1f_ca_w_1_360_s_1_980 = '-6.21875e-07*ic_cap*ic_cap+-3.62500e-07*ic_cap+5.71000e-05'
+ mcm3l1f_ca_w_1_360_s_4_500 = '-6.21875e-07*ic_cap*ic_cap+-3.62500e-07*ic_cap+5.71000e-05'
+ mcm3l1f_cc_w_0_170_s_0_180 = '-7.62500e-13*ic_cap*ic_cap+-5.00000e-13*ic_cap+7.71000e-11'
+ mcm3l1f_cc_w_0_170_s_0_225 = '-5.53125e-13*ic_cap*ic_cap+-3.62500e-13*ic_cap+6.52000e-11'
+ mcm3l1f_cc_w_0_170_s_0_270 = '-4.03125e-13*ic_cap*ic_cap+-2.87500e-13*ic_cap+5.70000e-11'
+ mcm3l1f_cc_w_0_170_s_0_360 = '-2.56250e-13*ic_cap*ic_cap+-1.75000e-13*ic_cap+4.55000e-11'
+ mcm3l1f_cc_w_0_170_s_0_450 = '-1.59375e-13*ic_cap*ic_cap+-1.37500e-13*ic_cap+3.81000e-11'
+ mcm3l1f_cc_w_0_170_s_0_540 = '-9.68750e-14*ic_cap*ic_cap+-8.75000e-14*ic_cap+3.22000e-11'
+ mcm3l1f_cc_w_0_170_s_0_720 = '-2.50000e-14*ic_cap*ic_cap+-5.00000e-14*ic_cap+2.43000e-11'
+ mcm3l1f_cc_w_0_170_s_1_080 = '4.06250e-14*ic_cap*ic_cap+1.25000e-14*ic_cap+1.48000e-11'
+ mcm3l1f_cc_w_0_170_s_1_980 = '6.21875e-14*ic_cap*ic_cap+3.37500e-14*ic_cap+4.96000e-12'
+ mcm3l1f_cc_w_0_170_s_4_500 = '1.50000e-14*ic_cap*ic_cap+1.12500e-14*ic_cap+3.10000e-13'
+ mcm3l1f_cc_w_1_360_s_0_180 = '-5.96875e-13*ic_cap*ic_cap+-3.87500e-13*ic_cap+9.02000e-11'
+ mcm3l1f_cc_w_1_360_s_0_225 = '-3.78125e-13*ic_cap*ic_cap+-2.62500e-13*ic_cap+7.69000e-11'
+ mcm3l1f_cc_w_1_360_s_0_270 = '-2.53125e-13*ic_cap*ic_cap+-1.87500e-13*ic_cap+6.75000e-11'
+ mcm3l1f_cc_w_1_360_s_0_360 = '-1.03125e-13*ic_cap*ic_cap+-8.75000e-14*ic_cap+5.44000e-11'
+ mcm3l1f_cc_w_1_360_s_0_450 = '-2.18750e-14*ic_cap*ic_cap+-3.75000e-14*ic_cap+4.55000e-11'
+ mcm3l1f_cc_w_1_360_s_0_540 = '2.50000e-14*ic_cap*ic_cap+3.89000e-11'
+ mcm3l1f_cc_w_1_360_s_0_720 = '8.43750e-14*ic_cap*ic_cap+3.75000e-14*ic_cap+2.95000e-11'
+ mcm3l1f_cc_w_1_360_s_1_080 = '1.25000e-13*ic_cap*ic_cap+7.50000e-14*ic_cap+1.83000e-11'
+ mcm3l1f_cc_w_1_360_s_1_980 = '1.11563e-13*ic_cap*ic_cap+6.62500e-14*ic_cap+6.38000e-12'
+ mcm3l1f_cc_w_1_360_s_4_500 = '2.43750e-14*ic_cap*ic_cap+1.87500e-14*ic_cap+3.95000e-13'
+ mcm3l1f_cf_w_0_170_s_0_180 = '-1.37500e-14*ic_cap*ic_cap+-7.50000e-15*ic_cap+5.03000e-12'
+ mcm3l1f_cf_w_0_170_s_0_225 = '-2.84375e-14*ic_cap*ic_cap+-1.62500e-14*ic_cap+6.25000e-12'
+ mcm3l1f_cf_w_0_170_s_0_270 = '-4.09375e-14*ic_cap*ic_cap+-2.62500e-14*ic_cap+7.41000e-12'
+ mcm3l1f_cf_w_0_170_s_0_360 = '-6.53125e-14*ic_cap*ic_cap+-3.62500e-14*ic_cap+9.84000e-12'
+ mcm3l1f_cf_w_0_170_s_0_450 = '-8.75000e-14*ic_cap*ic_cap+-5.00000e-14*ic_cap+1.18000e-11'
+ mcm3l1f_cf_w_0_170_s_0_540 = '-1.09375e-13*ic_cap*ic_cap+-6.25000e-14*ic_cap+1.40000e-11'
+ mcm3l1f_cf_w_0_170_s_0_720 = '-1.46875e-13*ic_cap*ic_cap+-8.75000e-14*ic_cap+1.76000e-11'
+ mcm3l1f_cf_w_0_170_s_1_080 = '-1.93750e-13*ic_cap*ic_cap+-1.25000e-13*ic_cap+2.32000e-11'
+ mcm3l1f_cf_w_0_170_s_1_980 = '-2.31250e-13*ic_cap*ic_cap+-1.50000e-13*ic_cap+3.10000e-11'
+ mcm3l1f_cf_w_0_170_s_4_500 = '-1.90625e-13*ic_cap*ic_cap+-1.37500e-13*ic_cap+3.53000e-11'
+ mcm3l1f_cf_w_1_360_s_0_180 = '-1.40625e-14*ic_cap*ic_cap+-8.75000e-15*ic_cap+5.01000e-12'
+ mcm3l1f_cf_w_1_360_s_0_225 = '-2.71875e-14*ic_cap*ic_cap+-1.62500e-14*ic_cap+6.22000e-12'
+ mcm3l1f_cf_w_1_360_s_0_270 = '-4.03125e-14*ic_cap*ic_cap+-2.37500e-14*ic_cap+7.41000e-12'
+ mcm3l1f_cf_w_1_360_s_0_360 = '-6.53125e-14*ic_cap*ic_cap+-3.87500e-14*ic_cap+9.72000e-12'
+ mcm3l1f_cf_w_1_360_s_0_450 = '-8.75000e-14*ic_cap*ic_cap+-5.00000e-14*ic_cap+1.19000e-11'
+ mcm3l1f_cf_w_1_360_s_0_540 = '-1.09375e-13*ic_cap*ic_cap+-6.25000e-14*ic_cap+1.40000e-11'
+ mcm3l1f_cf_w_1_360_s_0_720 = '-1.46875e-13*ic_cap*ic_cap+-8.75000e-14*ic_cap+1.78000e-11'
+ mcm3l1f_cf_w_1_360_s_1_080 = '-1.90625e-13*ic_cap*ic_cap+-1.12500e-13*ic_cap+2.40000e-11'
+ mcm3l1f_cf_w_1_360_s_1_980 = '-2.15625e-13*ic_cap*ic_cap+-1.37500e-13*ic_cap+3.31000e-11'
+ mcm3l1f_cf_w_1_360_s_4_500 = '-1.40625e-13*ic_cap*ic_cap+-8.75000e-14*ic_cap+3.86000e-11'
+ mcm3l1p1_ca_w_0_170_s_0_180 = '-1.83750e-06*ic_cap*ic_cap+-9.25000e-07*ic_cap+1.14000e-04'
+ mcm3l1p1_ca_w_0_170_s_0_225 = '-1.83750e-06*ic_cap*ic_cap+-9.25000e-07*ic_cap+1.14000e-04'
+ mcm3l1p1_ca_w_0_170_s_0_270 = '-1.83750e-06*ic_cap*ic_cap+-9.25000e-07*ic_cap+1.14000e-04'
+ mcm3l1p1_ca_w_0_170_s_0_360 = '-1.83750e-06*ic_cap*ic_cap+-9.25000e-07*ic_cap+1.14000e-04'
+ mcm3l1p1_ca_w_0_170_s_0_450 = '-1.83750e-06*ic_cap*ic_cap+-9.25000e-07*ic_cap+1.14000e-04'
+ mcm3l1p1_ca_w_0_170_s_0_540 = '-1.83750e-06*ic_cap*ic_cap+-9.25000e-07*ic_cap+1.14000e-04'
+ mcm3l1p1_ca_w_0_170_s_0_720 = '-1.83750e-06*ic_cap*ic_cap+-9.25000e-07*ic_cap+1.14000e-04'
+ mcm3l1p1_ca_w_0_170_s_1_080 = '-1.83750e-06*ic_cap*ic_cap+-9.25000e-07*ic_cap+1.14000e-04'
+ mcm3l1p1_ca_w_0_170_s_1_980 = '-1.83750e-06*ic_cap*ic_cap+-9.25000e-07*ic_cap+1.14000e-04'
+ mcm3l1p1_ca_w_0_170_s_4_500 = '-1.83750e-06*ic_cap*ic_cap+-9.25000e-07*ic_cap+1.14000e-04'
+ mcm3l1p1_ca_w_1_360_s_0_180 = '-1.83750e-06*ic_cap*ic_cap+-9.25000e-07*ic_cap+1.14000e-04'
+ mcm3l1p1_ca_w_1_360_s_0_225 = '-1.83750e-06*ic_cap*ic_cap+-9.25000e-07*ic_cap+1.14000e-04'
+ mcm3l1p1_ca_w_1_360_s_0_270 = '-1.83750e-06*ic_cap*ic_cap+-9.25000e-07*ic_cap+1.14000e-04'
+ mcm3l1p1_ca_w_1_360_s_0_360 = '-1.83750e-06*ic_cap*ic_cap+-9.25000e-07*ic_cap+1.14000e-04'
+ mcm3l1p1_ca_w_1_360_s_0_450 = '-1.83750e-06*ic_cap*ic_cap+-9.25000e-07*ic_cap+1.14000e-04'
+ mcm3l1p1_ca_w_1_360_s_0_540 = '-1.83750e-06*ic_cap*ic_cap+-9.25000e-07*ic_cap+1.14000e-04'
+ mcm3l1p1_ca_w_1_360_s_0_720 = '-1.83750e-06*ic_cap*ic_cap+-9.25000e-07*ic_cap+1.14000e-04'
+ mcm3l1p1_ca_w_1_360_s_1_080 = '-1.83750e-06*ic_cap*ic_cap+-9.25000e-07*ic_cap+1.14000e-04'
+ mcm3l1p1_ca_w_1_360_s_1_980 = '-1.83750e-06*ic_cap*ic_cap+-9.25000e-07*ic_cap+1.14000e-04'
+ mcm3l1p1_ca_w_1_360_s_4_500 = '-1.83750e-06*ic_cap*ic_cap+-9.25000e-07*ic_cap+1.14000e-04'
+ mcm3l1p1_cc_w_0_170_s_0_180 = '-6.50000e-13*ic_cap*ic_cap+-4.50000e-13*ic_cap+7.05000e-11'
+ mcm3l1p1_cc_w_0_170_s_0_225 = '-4.31250e-13*ic_cap*ic_cap+-3.25000e-13*ic_cap+5.82000e-11'
+ mcm3l1p1_cc_w_0_170_s_0_270 = '-2.81250e-13*ic_cap*ic_cap+-2.25000e-13*ic_cap+4.96000e-11'
+ mcm3l1p1_cc_w_0_170_s_0_360 = '-1.25000e-13*ic_cap*ic_cap+-1.25000e-13*ic_cap+3.76000e-11'
+ mcm3l1p1_cc_w_0_170_s_0_450 = '-3.75000e-14*ic_cap*ic_cap+-7.50000e-14*ic_cap+3.00000e-11'
+ mcm3l1p1_cc_w_0_170_s_0_540 = '6.25000e-15*ic_cap*ic_cap+-2.50000e-14*ic_cap+2.42000e-11'
+ mcm3l1p1_cc_w_0_170_s_0_720 = '7.18750e-14*ic_cap*ic_cap+1.25000e-14*ic_cap+1.64000e-11'
+ mcm3l1p1_cc_w_0_170_s_1_080 = '9.00000e-14*ic_cap*ic_cap+4.00000e-14*ic_cap+8.31000e-12'
+ mcm3l1p1_cc_w_0_170_s_1_980 = '5.37500e-14*ic_cap*ic_cap+3.00000e-14*ic_cap+1.89000e-12'
+ mcm3l1p1_cc_w_0_170_s_4_500 = '5.78125e-15*ic_cap*ic_cap+4.37500e-15*ic_cap+7.00000e-14'
+ mcm3l1p1_cc_w_1_360_s_0_180 = '-4.96875e-13*ic_cap*ic_cap+-3.37500e-13*ic_cap+7.98000e-11'
+ mcm3l1p1_cc_w_1_360_s_0_225 = '-2.87500e-13*ic_cap*ic_cap+-2.25000e-13*ic_cap+6.68000e-11'
+ mcm3l1p1_cc_w_1_360_s_0_270 = '-1.53125e-13*ic_cap*ic_cap+-1.37500e-13*ic_cap+5.72000e-11'
+ mcm3l1p1_cc_w_1_360_s_0_360 = '-1.25000e-14*ic_cap*ic_cap+-2.50000e-14*ic_cap+4.43000e-11'
+ mcm3l1p1_cc_w_1_360_s_0_450 = '6.25000e-14*ic_cap*ic_cap+3.56000e-11'
+ mcm3l1p1_cc_w_1_360_s_0_540 = '1.09375e-13*ic_cap*ic_cap+3.75000e-14*ic_cap+2.92000e-11'
+ mcm3l1p1_cc_w_1_360_s_0_720 = '1.50000e-13*ic_cap*ic_cap+7.50000e-14*ic_cap+2.05000e-11'
+ mcm3l1p1_cc_w_1_360_s_1_080 = '1.59375e-13*ic_cap*ic_cap+8.75000e-14*ic_cap+1.09000e-11'
+ mcm3l1p1_cc_w_1_360_s_1_980 = '8.84375e-14*ic_cap*ic_cap+6.87500e-14*ic_cap+2.72000e-12'
+ mcm3l1p1_cc_w_1_360_s_4_500 = '9.21875e-15*ic_cap*ic_cap+-6.25000e-16*ic_cap+1.05000e-13'
+ mcm3l1p1_cf_w_0_170_s_0_180 = '-8.68750e-14*ic_cap*ic_cap+-4.25000e-14*ic_cap+9.84000e-12'
+ mcm3l1p1_cf_w_0_170_s_0_225 = '-1.22500e-13*ic_cap*ic_cap+-6.50000e-14*ic_cap+1.21000e-11'
+ mcm3l1p1_cf_w_0_170_s_0_270 = '-1.56250e-13*ic_cap*ic_cap+-7.50000e-14*ic_cap+1.42000e-11'
+ mcm3l1p1_cf_w_0_170_s_0_360 = '-2.15625e-13*ic_cap*ic_cap+-1.12500e-13*ic_cap+1.84000e-11'
+ mcm3l1p1_cf_w_0_170_s_0_450 = '-2.65625e-13*ic_cap*ic_cap+-1.37500e-13*ic_cap+2.18000e-11'
+ mcm3l1p1_cf_w_0_170_s_0_540 = '-3.09375e-13*ic_cap*ic_cap+-1.62500e-13*ic_cap+2.51000e-11'
+ mcm3l1p1_cf_w_0_170_s_0_720 = '-3.62500e-13*ic_cap*ic_cap+-2.00000e-13*ic_cap+3.01000e-11'
+ mcm3l1p1_cf_w_0_170_s_1_080 = '-4.03125e-13*ic_cap*ic_cap+-2.37500e-13*ic_cap+3.65000e-11'
+ mcm3l1p1_cf_w_0_170_s_1_980 = '-3.75000e-13*ic_cap*ic_cap+-2.25000e-13*ic_cap+4.22000e-11'
+ mcm3l1p1_cf_w_0_170_s_4_500 = '-3.31250e-13*ic_cap*ic_cap+-2.00000e-13*ic_cap+4.40000e-11'
+ mcm3l1p1_cf_w_1_360_s_0_180 = '-8.59375e-14*ic_cap*ic_cap+-4.12500e-14*ic_cap+9.83000e-12'
+ mcm3l1p1_cf_w_1_360_s_0_225 = '-1.21250e-13*ic_cap*ic_cap+-6.00000e-14*ic_cap+1.21000e-11'
+ mcm3l1p1_cf_w_1_360_s_0_270 = '-1.50000e-13*ic_cap*ic_cap+-7.50000e-14*ic_cap+1.42000e-11'
+ mcm3l1p1_cf_w_1_360_s_0_360 = '-2.15625e-13*ic_cap*ic_cap+-1.12500e-13*ic_cap+1.83000e-11'
+ mcm3l1p1_cf_w_1_360_s_0_450 = '-2.59375e-13*ic_cap*ic_cap+-1.37500e-13*ic_cap+2.19000e-11'
+ mcm3l1p1_cf_w_1_360_s_0_540 = '-3.03125e-13*ic_cap*ic_cap+-1.62500e-13*ic_cap+2.52000e-11'
+ mcm3l1p1_cf_w_1_360_s_0_720 = '-3.53125e-13*ic_cap*ic_cap+-1.87500e-13*ic_cap+3.05000e-11'
+ mcm3l1p1_cf_w_1_360_s_1_080 = '-3.93750e-13*ic_cap*ic_cap+-2.25000e-13*ic_cap+3.78000e-11'
+ mcm3l1p1_cf_w_1_360_s_1_980 = '-3.53125e-13*ic_cap*ic_cap+-2.12500e-13*ic_cap+4.51000e-11'
+ mcm3l1p1_cf_w_1_360_s_4_500 = '-2.84375e-13*ic_cap*ic_cap+-1.62500e-13*ic_cap+4.77000e-11'
+ mcm3m1_ca_w_0_300_s_0_300 = '-3.90625e-07*ic_cap*ic_cap+-2.12500e-07*ic_cap+3.29000e-05'
+ mcm3m1_ca_w_0_300_s_0_360 = '-3.90625e-07*ic_cap*ic_cap+-2.12500e-07*ic_cap+3.29000e-05'
+ mcm3m1_ca_w_0_300_s_0_450 = '-3.90625e-07*ic_cap*ic_cap+-2.12500e-07*ic_cap+3.29000e-05'
+ mcm3m1_ca_w_0_300_s_0_600 = '-3.90625e-07*ic_cap*ic_cap+-2.12500e-07*ic_cap+3.29000e-05'
+ mcm3m1_ca_w_0_300_s_0_800 = '-3.90625e-07*ic_cap*ic_cap+-2.12500e-07*ic_cap+3.29000e-05'
+ mcm3m1_ca_w_0_300_s_1_000 = '-3.90625e-07*ic_cap*ic_cap+-2.12500e-07*ic_cap+3.29000e-05'
+ mcm3m1_ca_w_0_300_s_1_200 = '-3.90625e-07*ic_cap*ic_cap+-2.12500e-07*ic_cap+3.29000e-05'
+ mcm3m1_ca_w_0_300_s_2_100 = '-3.90625e-07*ic_cap*ic_cap+-2.12500e-07*ic_cap+3.29000e-05'
+ mcm3m1_ca_w_0_300_s_3_300 = '-3.90625e-07*ic_cap*ic_cap+-2.12500e-07*ic_cap+3.29000e-05'
+ mcm3m1_ca_w_0_300_s_9_000 = '-3.90625e-07*ic_cap*ic_cap+-2.12500e-07*ic_cap+3.29000e-05'
+ mcm3m1_ca_w_2_400_s_0_300 = '-3.90625e-07*ic_cap*ic_cap+-2.12500e-07*ic_cap+3.29000e-05'
+ mcm3m1_ca_w_2_400_s_0_360 = '-3.90625e-07*ic_cap*ic_cap+-2.12500e-07*ic_cap+3.29000e-05'
+ mcm3m1_ca_w_2_400_s_0_450 = '-3.90625e-07*ic_cap*ic_cap+-2.12500e-07*ic_cap+3.29000e-05'
+ mcm3m1_ca_w_2_400_s_0_600 = '-3.90625e-07*ic_cap*ic_cap+-2.12500e-07*ic_cap+3.29000e-05'
+ mcm3m1_ca_w_2_400_s_0_800 = '-3.90625e-07*ic_cap*ic_cap+-2.12500e-07*ic_cap+3.29000e-05'
+ mcm3m1_ca_w_2_400_s_1_000 = '-3.90625e-07*ic_cap*ic_cap+-2.12500e-07*ic_cap+3.29000e-05'
+ mcm3m1_ca_w_2_400_s_1_200 = '-3.90625e-07*ic_cap*ic_cap+-2.12500e-07*ic_cap+3.29000e-05'
+ mcm3m1_ca_w_2_400_s_2_100 = '-3.90625e-07*ic_cap*ic_cap+-2.12500e-07*ic_cap+3.29000e-05'
+ mcm3m1_ca_w_2_400_s_3_300 = '-3.90625e-07*ic_cap*ic_cap+-2.12500e-07*ic_cap+3.29000e-05'
+ mcm3m1_ca_w_2_400_s_9_000 = '-3.90625e-07*ic_cap*ic_cap+-2.12500e-07*ic_cap+3.29000e-05'
+ mcm3m1_cc_w_0_300_s_0_300 = '-7.56250e-13*ic_cap*ic_cap+-4.25000e-13*ic_cap+1.02000e-10'
+ mcm3m1_cc_w_0_300_s_0_360 = '-6.40625e-13*ic_cap*ic_cap+-3.62500e-13*ic_cap+9.42000e-11'
+ mcm3m1_cc_w_0_300_s_0_450 = '-5.18750e-13*ic_cap*ic_cap+-3.25000e-13*ic_cap+8.43000e-11'
+ mcm3m1_cc_w_0_300_s_0_600 = '-3.81250e-13*ic_cap*ic_cap+-2.50000e-13*ic_cap+7.13000e-11'
+ mcm3m1_cc_w_0_300_s_0_800 = '-2.59375e-13*ic_cap*ic_cap+-1.62500e-13*ic_cap+5.87000e-11'
+ mcm3m1_cc_w_0_300_s_1_000 = '-1.68750e-13*ic_cap*ic_cap+-1.25000e-13*ic_cap+4.91000e-11'
+ mcm3m1_cc_w_0_300_s_1_200 = '-1.12500e-13*ic_cap*ic_cap+-7.50000e-14*ic_cap+4.20000e-11'
+ mcm3m1_cc_w_0_300_s_2_100 = '-1.56250e-14*ic_cap*ic_cap+-1.25000e-14*ic_cap+2.43000e-11'
+ mcm3m1_cc_w_0_300_s_3_300 = '1.87500e-14*ic_cap*ic_cap+1.48000e-11'
+ mcm3m1_cc_w_0_300_s_9_000 = '1.09375e-14*ic_cap*ic_cap+3.75000e-15*ic_cap+3.27000e-12'
+ mcm3m1_cc_w_2_400_s_0_300 = '-6.56250e-13*ic_cap*ic_cap+-3.75000e-13*ic_cap+1.21000e-10'
+ mcm3m1_cc_w_2_400_s_0_360 = '-5.93750e-13*ic_cap*ic_cap+-3.75000e-13*ic_cap+1.13000e-10'
+ mcm3m1_cc_w_2_400_s_0_450 = '-4.71875e-13*ic_cap*ic_cap+-2.37500e-13*ic_cap+1.02000e-10'
+ mcm3m1_cc_w_2_400_s_0_600 = '-3.31250e-13*ic_cap*ic_cap+-2.00000e-13*ic_cap+8.70000e-11'
+ mcm3m1_cc_w_2_400_s_0_800 = '-2.06250e-13*ic_cap*ic_cap+-1.50000e-13*ic_cap+7.25000e-11'
+ mcm3m1_cc_w_2_400_s_1_000 = '-1.31250e-13*ic_cap*ic_cap+-1.00000e-13*ic_cap+6.18000e-11'
+ mcm3m1_cc_w_2_400_s_1_200 = '-8.43750e-14*ic_cap*ic_cap+-6.25000e-14*ic_cap+5.38000e-11'
+ mcm3m1_cc_w_2_400_s_2_100 = '3.12500e-15*ic_cap*ic_cap+-1.25000e-14*ic_cap+3.39000e-11'
+ mcm3m1_cc_w_2_400_s_3_300 = '2.18750e-14*ic_cap*ic_cap+1.25000e-14*ic_cap+2.20000e-11'
+ mcm3m1_cc_w_2_400_s_9_000 = '2.18750e-14*ic_cap*ic_cap+1.25000e-14*ic_cap+6.00000e-12'
+ mcm3m1_cf_w_0_300_s_0_300 = '-2.28125e-14*ic_cap*ic_cap+-1.37500e-14*ic_cap+4.72000e-12'
+ mcm3m1_cf_w_0_300_s_0_360 = '-3.34375e-14*ic_cap*ic_cap+-1.87500e-14*ic_cap+5.62000e-12'
+ mcm3m1_cf_w_0_300_s_0_450 = '-4.68750e-14*ic_cap*ic_cap+-2.75000e-14*ic_cap+6.94000e-12'
+ mcm3m1_cf_w_0_300_s_0_600 = '-6.96875e-14*ic_cap*ic_cap+-3.87500e-14*ic_cap+9.07000e-12'
+ mcm3m1_cf_w_0_300_s_0_800 = '-9.56250e-14*ic_cap*ic_cap+-5.75000e-14*ic_cap+1.16000e-11'
+ mcm3m1_cf_w_0_300_s_1_000 = '-1.25000e-13*ic_cap*ic_cap+-7.50000e-14*ic_cap+1.41000e-11'
+ mcm3m1_cf_w_0_300_s_1_200 = '-1.46875e-13*ic_cap*ic_cap+-8.75000e-14*ic_cap+1.64000e-11'
+ mcm3m1_cf_w_0_300_s_2_100 = '-2.06250e-13*ic_cap*ic_cap+-1.25000e-13*ic_cap+2.51000e-11'
+ mcm3m1_cf_w_0_300_s_3_300 = '-2.43750e-13*ic_cap*ic_cap+-1.50000e-13*ic_cap+3.17000e-11'
+ mcm3m1_cf_w_0_300_s_9_000 = '-2.50000e-13*ic_cap*ic_cap+-1.50000e-13*ic_cap+4.21000e-11'
+ mcm3m1_cf_w_2_400_s_0_300 = '-2.25000e-14*ic_cap*ic_cap+-1.25000e-14*ic_cap+4.73000e-12'
+ mcm3m1_cf_w_2_400_s_0_360 = '-3.34375e-14*ic_cap*ic_cap+-1.87500e-14*ic_cap+5.64000e-12'
+ mcm3m1_cf_w_2_400_s_0_450 = '-4.78125e-14*ic_cap*ic_cap+-2.87500e-14*ic_cap+6.95000e-12'
+ mcm3m1_cf_w_2_400_s_0_600 = '-7.03125e-14*ic_cap*ic_cap+-4.12500e-14*ic_cap+9.05000e-12'
+ mcm3m1_cf_w_2_400_s_0_800 = '-9.65625e-14*ic_cap*ic_cap+-6.12500e-14*ic_cap+1.17000e-11'
+ mcm3m1_cf_w_2_400_s_1_000 = '-1.21875e-13*ic_cap*ic_cap+-6.25000e-14*ic_cap+1.42000e-11'
+ mcm3m1_cf_w_2_400_s_1_200 = '-1.43750e-13*ic_cap*ic_cap+-7.50000e-14*ic_cap+1.65000e-11'
+ mcm3m1_cf_w_2_400_s_2_100 = '-2.00000e-13*ic_cap*ic_cap+-1.25000e-13*ic_cap+2.49000e-11'
+ mcm3m1_cf_w_2_400_s_3_300 = '-2.37500e-13*ic_cap*ic_cap+-1.50000e-13*ic_cap+3.27000e-11'
+ mcm3m1_cf_w_2_400_s_9_000 = '-2.46875e-13*ic_cap*ic_cap+-1.62500e-13*ic_cap+4.65000e-11'
+ mcm3m1d_ca_w_0_140_s_0_140 = '-7.59375e-07*ic_cap*ic_cap+-4.62500e-07*ic_cap+6.65000e-05'
+ mcm3m1d_ca_w_0_140_s_0_175 = '-7.59375e-07*ic_cap*ic_cap+-4.62500e-07*ic_cap+6.65000e-05'
+ mcm3m1d_ca_w_0_140_s_0_210 = '-7.59375e-07*ic_cap*ic_cap+-4.62500e-07*ic_cap+6.65000e-05'
+ mcm3m1d_ca_w_0_140_s_0_280 = '-7.59375e-07*ic_cap*ic_cap+-4.62500e-07*ic_cap+6.65000e-05'
+ mcm3m1d_ca_w_0_140_s_0_350 = '-7.59375e-07*ic_cap*ic_cap+-4.62500e-07*ic_cap+6.65000e-05'
+ mcm3m1d_ca_w_0_140_s_0_420 = '-7.59375e-07*ic_cap*ic_cap+-4.62500e-07*ic_cap+6.65000e-05'
+ mcm3m1d_ca_w_0_140_s_0_560 = '-7.59375e-07*ic_cap*ic_cap+-4.62500e-07*ic_cap+6.65000e-05'
+ mcm3m1d_ca_w_0_140_s_0_840 = '-7.59375e-07*ic_cap*ic_cap+-4.62500e-07*ic_cap+6.65000e-05'
+ mcm3m1d_ca_w_0_140_s_1_540 = '-7.59375e-07*ic_cap*ic_cap+-4.62500e-07*ic_cap+6.65000e-05'
+ mcm3m1d_ca_w_0_140_s_3_500 = '-7.59375e-07*ic_cap*ic_cap+-4.62500e-07*ic_cap+6.65000e-05'
+ mcm3m1d_ca_w_1_120_s_0_140 = '-7.59375e-07*ic_cap*ic_cap+-4.62500e-07*ic_cap+6.65000e-05'
+ mcm3m1d_ca_w_1_120_s_0_175 = '-7.59375e-07*ic_cap*ic_cap+-4.62500e-07*ic_cap+6.65000e-05'
+ mcm3m1d_ca_w_1_120_s_0_210 = '-7.59375e-07*ic_cap*ic_cap+-4.62500e-07*ic_cap+6.65000e-05'
+ mcm3m1d_ca_w_1_120_s_0_280 = '-7.59375e-07*ic_cap*ic_cap+-4.62500e-07*ic_cap+6.65000e-05'
+ mcm3m1d_ca_w_1_120_s_0_350 = '-7.59375e-07*ic_cap*ic_cap+-4.62500e-07*ic_cap+6.65000e-05'
+ mcm3m1d_ca_w_1_120_s_0_420 = '-7.59375e-07*ic_cap*ic_cap+-4.62500e-07*ic_cap+6.65000e-05'
+ mcm3m1d_ca_w_1_120_s_0_560 = '-7.59375e-07*ic_cap*ic_cap+-4.62500e-07*ic_cap+6.65000e-05'
+ mcm3m1d_ca_w_1_120_s_0_840 = '-7.59375e-07*ic_cap*ic_cap+-4.62500e-07*ic_cap+6.65000e-05'
+ mcm3m1d_ca_w_1_120_s_1_540 = '-7.59375e-07*ic_cap*ic_cap+-4.62500e-07*ic_cap+6.65000e-05'
+ mcm3m1d_ca_w_1_120_s_3_500 = '-7.59375e-07*ic_cap*ic_cap+-4.62500e-07*ic_cap+6.65000e-05'
+ mcm3m1d_cc_w_0_140_s_0_140 = '-8.68750e-13*ic_cap*ic_cap+-5.25000e-13*ic_cap+9.98000e-11'
+ mcm3m1d_cc_w_0_140_s_0_175 = '-8.46875e-13*ic_cap*ic_cap+-3.37500e-13*ic_cap+9.81000e-11'
+ mcm3m1d_cc_w_0_140_s_0_210 = '-7.03125e-13*ic_cap*ic_cap+-4.37500e-13*ic_cap+9.26000e-11'
+ mcm3m1d_cc_w_0_140_s_0_280 = '-5.06250e-13*ic_cap*ic_cap+-3.75000e-13*ic_cap+8.03000e-11'
+ mcm3m1d_cc_w_0_140_s_0_350 = '-4.09375e-13*ic_cap*ic_cap+-2.37500e-13*ic_cap+6.89000e-11'
+ mcm3m1d_cc_w_0_140_s_0_420 = '-2.53125e-13*ic_cap*ic_cap+-1.87500e-13*ic_cap+5.84000e-11'
+ mcm3m1d_cc_w_0_140_s_0_560 = '-1.00000e-13*ic_cap*ic_cap+-7.50000e-14*ic_cap+4.41000e-11'
+ mcm3m1d_cc_w_0_140_s_0_840 = '1.56250e-14*ic_cap*ic_cap+-1.25000e-14*ic_cap+2.81000e-11'
+ mcm3m1d_cc_w_0_140_s_1_540 = '9.06250e-14*ic_cap*ic_cap+6.25000e-14*ic_cap+1.07000e-11'
+ mcm3m1d_cc_w_0_140_s_3_500 = '3.34375e-14*ic_cap*ic_cap+2.62500e-14*ic_cap+9.30000e-13'
+ mcm3m1d_cc_w_1_120_s_0_140 = '-7.50000e-13*ic_cap*ic_cap+-5.00000e-13*ic_cap+1.15000e-10'
+ mcm3m1d_cc_w_1_120_s_0_175 = '-7.12500e-13*ic_cap*ic_cap+-3.50000e-13*ic_cap+1.11000e-10'
+ mcm3m1d_cc_w_1_120_s_0_210 = '-5.31250e-13*ic_cap*ic_cap+-3.50000e-13*ic_cap+1.03000e-10'
+ mcm3m1d_cc_w_1_120_s_0_280 = '-3.34375e-13*ic_cap*ic_cap+-2.12500e-13*ic_cap+8.87000e-11'
+ mcm3m1d_cc_w_1_120_s_0_350 = '-2.62500e-13*ic_cap*ic_cap+-1.75000e-13*ic_cap+7.63000e-11'
+ mcm3m1d_cc_w_1_120_s_0_420 = '-1.43750e-13*ic_cap*ic_cap+-7.50000e-14*ic_cap+6.51000e-11'
+ mcm3m1d_cc_w_1_120_s_0_560 = '-9.37500e-15*ic_cap*ic_cap+-1.25000e-14*ic_cap+4.92000e-11'
+ mcm3m1d_cc_w_1_120_s_0_840 = '9.37500e-14*ic_cap*ic_cap+5.00000e-14*ic_cap+3.11000e-11'
+ mcm3m1d_cc_w_1_120_s_1_540 = '1.37500e-13*ic_cap*ic_cap+7.50000e-14*ic_cap+1.20000e-11'
+ mcm3m1d_cc_w_1_120_s_3_500 = '4.09375e-14*ic_cap*ic_cap+3.87500e-14*ic_cap+1.08000e-12'
+ mcm3m1d_cf_w_0_140_s_0_140 = '-1.00000e-14*ic_cap*ic_cap+-7.50000e-15*ic_cap+4.57000e-12'
+ mcm3m1d_cf_w_0_140_s_0_175 = '-2.25000e-14*ic_cap*ic_cap+-1.50000e-14*ic_cap+5.69000e-12'
+ mcm3m1d_cf_w_0_140_s_0_210 = '-3.31250e-14*ic_cap*ic_cap+-2.25000e-14*ic_cap+6.82000e-12'
+ mcm3m1d_cf_w_0_140_s_0_280 = '-5.93750e-14*ic_cap*ic_cap+-3.75000e-14*ic_cap+9.01000e-12'
+ mcm3m1d_cf_w_0_140_s_0_350 = '-8.78125e-14*ic_cap*ic_cap+-5.12500e-14*ic_cap+1.12000e-11'
+ mcm3m1d_cf_w_0_140_s_0_420 = '-1.06250e-13*ic_cap*ic_cap+-7.50000e-14*ic_cap+1.33000e-11'
+ mcm3m1d_cf_w_0_140_s_0_560 = '-1.46875e-13*ic_cap*ic_cap+-8.75000e-14*ic_cap+1.72000e-11'
+ mcm3m1d_cf_w_0_140_s_0_840 = '-2.15625e-13*ic_cap*ic_cap+-1.37500e-13*ic_cap+2.40000e-11'
+ mcm3m1d_cf_w_0_140_s_1_540 = '-2.93750e-13*ic_cap*ic_cap+-2.00000e-13*ic_cap+3.53000e-11'
+ mcm3m1d_cf_w_0_140_s_3_500 = '-2.75000e-13*ic_cap*ic_cap+-1.75000e-13*ic_cap+4.43000e-11'
+ mcm3m1d_cf_w_1_120_s_0_140 = '-1.00000e-14*ic_cap*ic_cap+-5.00000e-15*ic_cap+4.62000e-12'
+ mcm3m1d_cf_w_1_120_s_0_175 = '-2.25000e-14*ic_cap*ic_cap+-1.50000e-14*ic_cap+5.75000e-12'
+ mcm3m1d_cf_w_1_120_s_0_210 = '-3.65625e-14*ic_cap*ic_cap+-2.37500e-14*ic_cap+6.88000e-12'
+ mcm3m1d_cf_w_1_120_s_0_280 = '-6.00000e-14*ic_cap*ic_cap+-4.00000e-14*ic_cap+9.07000e-12'
+ mcm3m1d_cf_w_1_120_s_0_350 = '-8.78125e-14*ic_cap*ic_cap+-5.12500e-14*ic_cap+1.13000e-11'
+ mcm3m1d_cf_w_1_120_s_0_420 = '-1.06250e-13*ic_cap*ic_cap+-7.50000e-14*ic_cap+1.33000e-11'
+ mcm3m1d_cf_w_1_120_s_0_560 = '-1.46875e-13*ic_cap*ic_cap+-8.75000e-14*ic_cap+1.73000e-11'
+ mcm3m1d_cf_w_1_120_s_0_840 = '-2.15625e-13*ic_cap*ic_cap+-1.37500e-13*ic_cap+2.43000e-11'
+ mcm3m1d_cf_w_1_120_s_1_540 = '-2.96875e-13*ic_cap*ic_cap+-1.87500e-13*ic_cap+3.64000e-11'
+ mcm3m1d_cf_w_1_120_s_3_500 = '-2.40625e-13*ic_cap*ic_cap+-1.62500e-13*ic_cap+4.62000e-11'
+ mcm3m1f_ca_w_0_140_s_0_140 = '-6.90625e-07*ic_cap*ic_cap+-4.12500e-07*ic_cap+5.87000e-05'
+ mcm3m1f_ca_w_0_140_s_0_175 = '-6.90625e-07*ic_cap*ic_cap+-4.12500e-07*ic_cap+5.87000e-05'
+ mcm3m1f_ca_w_0_140_s_0_210 = '-6.90625e-07*ic_cap*ic_cap+-4.12500e-07*ic_cap+5.87000e-05'
+ mcm3m1f_ca_w_0_140_s_0_280 = '-6.90625e-07*ic_cap*ic_cap+-4.12500e-07*ic_cap+5.87000e-05'
+ mcm3m1f_ca_w_0_140_s_0_350 = '-6.90625e-07*ic_cap*ic_cap+-4.12500e-07*ic_cap+5.87000e-05'
+ mcm3m1f_ca_w_0_140_s_0_420 = '-6.90625e-07*ic_cap*ic_cap+-4.12500e-07*ic_cap+5.87000e-05'
+ mcm3m1f_ca_w_0_140_s_0_560 = '-6.90625e-07*ic_cap*ic_cap+-4.12500e-07*ic_cap+5.87000e-05'
+ mcm3m1f_ca_w_0_140_s_0_840 = '-6.90625e-07*ic_cap*ic_cap+-4.12500e-07*ic_cap+5.87000e-05'
+ mcm3m1f_ca_w_0_140_s_1_540 = '-6.90625e-07*ic_cap*ic_cap+-4.12500e-07*ic_cap+5.87000e-05'
+ mcm3m1f_ca_w_0_140_s_3_500 = '-6.90625e-07*ic_cap*ic_cap+-4.12500e-07*ic_cap+5.87000e-05'
+ mcm3m1f_ca_w_1_120_s_0_140 = '-6.90625e-07*ic_cap*ic_cap+-4.12500e-07*ic_cap+5.87000e-05'
+ mcm3m1f_ca_w_1_120_s_0_175 = '-6.90625e-07*ic_cap*ic_cap+-4.12500e-07*ic_cap+5.87000e-05'
+ mcm3m1f_ca_w_1_120_s_0_210 = '-6.90625e-07*ic_cap*ic_cap+-4.12500e-07*ic_cap+5.87000e-05'
+ mcm3m1f_ca_w_1_120_s_0_280 = '-6.90625e-07*ic_cap*ic_cap+-4.12500e-07*ic_cap+5.87000e-05'
+ mcm3m1f_ca_w_1_120_s_0_350 = '-6.90625e-07*ic_cap*ic_cap+-4.12500e-07*ic_cap+5.87000e-05'
+ mcm3m1f_ca_w_1_120_s_0_420 = '-6.90625e-07*ic_cap*ic_cap+-4.12500e-07*ic_cap+5.87000e-05'
+ mcm3m1f_ca_w_1_120_s_0_560 = '-6.90625e-07*ic_cap*ic_cap+-4.12500e-07*ic_cap+5.87000e-05'
+ mcm3m1f_ca_w_1_120_s_0_840 = '-6.90625e-07*ic_cap*ic_cap+-4.12500e-07*ic_cap+5.87000e-05'
+ mcm3m1f_ca_w_1_120_s_1_540 = '-6.90625e-07*ic_cap*ic_cap+-4.12500e-07*ic_cap+5.87000e-05'
+ mcm3m1f_ca_w_1_120_s_3_500 = '-6.90625e-07*ic_cap*ic_cap+-4.12500e-07*ic_cap+5.87000e-05'
+ mcm3m1f_cc_w_0_140_s_0_140 = '-8.84375e-13*ic_cap*ic_cap+-4.87500e-13*ic_cap+1.01000e-10'
+ mcm3m1f_cc_w_0_140_s_0_175 = '-8.56250e-13*ic_cap*ic_cap+-3.50000e-13*ic_cap+9.91000e-11'
+ mcm3m1f_cc_w_0_140_s_0_210 = '-7.31250e-13*ic_cap*ic_cap+-4.00000e-13*ic_cap+9.37000e-11'
+ mcm3m1f_cc_w_0_140_s_0_280 = '-5.21875e-13*ic_cap*ic_cap+-3.62500e-13*ic_cap+8.17000e-11'
+ mcm3m1f_cc_w_0_140_s_0_350 = '-4.15625e-13*ic_cap*ic_cap+-2.62500e-13*ic_cap+7.03000e-11'
+ mcm3m1f_cc_w_0_140_s_0_420 = '-2.62500e-13*ic_cap*ic_cap+-1.75000e-13*ic_cap+5.99000e-11'
+ mcm3m1f_cc_w_0_140_s_0_560 = '-1.25000e-13*ic_cap*ic_cap+-7.50000e-14*ic_cap+4.61000e-11'
+ mcm3m1f_cc_w_0_140_s_0_840 = '1.56250e-14*ic_cap*ic_cap+-1.25000e-14*ic_cap+3.00000e-11'
+ mcm3m1f_cc_w_0_140_s_1_540 = '8.75000e-14*ic_cap*ic_cap+5.00000e-14*ic_cap+1.25000e-11'
+ mcm3m1f_cc_w_0_140_s_3_500 = '4.53125e-14*ic_cap*ic_cap+3.37500e-14*ic_cap+1.40000e-12'
+ mcm3m1f_cc_w_1_120_s_0_140 = '-6.25000e-13*ic_cap*ic_cap+-5.00000e-13*ic_cap+1.16000e-10'
+ mcm3m1f_cc_w_1_120_s_0_175 = '-6.87500e-13*ic_cap*ic_cap+-2.50000e-13*ic_cap+1.13000e-10'
+ mcm3m1f_cc_w_1_120_s_0_210 = '-5.40625e-13*ic_cap*ic_cap+-3.37500e-13*ic_cap+1.06000e-10'
+ mcm3m1f_cc_w_1_120_s_0_280 = '-3.53125e-13*ic_cap*ic_cap+-2.12500e-13*ic_cap+9.17000e-11'
+ mcm3m1f_cc_w_1_120_s_0_350 = '-2.62500e-13*ic_cap*ic_cap+-2.00000e-13*ic_cap+7.90000e-11'
+ mcm3m1f_cc_w_1_120_s_0_420 = '-1.53125e-13*ic_cap*ic_cap+-1.12500e-13*ic_cap+6.80000e-11'
+ mcm3m1f_cc_w_1_120_s_0_560 = '-1.25000e-14*ic_cap*ic_cap+-2.50000e-14*ic_cap+5.21000e-11'
+ mcm3m1f_cc_w_1_120_s_0_840 = '1.00000e-13*ic_cap*ic_cap+5.00000e-14*ic_cap+3.39000e-11'
+ mcm3m1f_cc_w_1_120_s_1_540 = '1.40625e-13*ic_cap*ic_cap+8.75000e-14*ic_cap+1.43000e-11'
+ mcm3m1f_cc_w_1_120_s_3_500 = '6.15625e-14*ic_cap*ic_cap+4.62500e-14*ic_cap+1.61000e-12'
+ mcm3m1f_cf_w_0_140_s_0_140 = '-1.00000e-14*ic_cap*ic_cap+-7.50000e-15*ic_cap+4.03000e-12'
+ mcm3m1f_cf_w_0_140_s_0_175 = '-2.15625e-14*ic_cap*ic_cap+-1.37500e-14*ic_cap+5.02000e-12'
+ mcm3m1f_cf_w_0_140_s_0_210 = '-3.15625e-14*ic_cap*ic_cap+-1.87500e-14*ic_cap+6.02000e-12'
+ mcm3m1f_cf_w_0_140_s_0_280 = '-5.53125e-14*ic_cap*ic_cap+-3.37500e-14*ic_cap+7.95000e-12'
+ mcm3m1f_cf_w_0_140_s_0_350 = '-7.81250e-14*ic_cap*ic_cap+-5.00000e-14*ic_cap+9.85000e-12'
+ mcm3m1f_cf_w_0_140_s_0_420 = '-1.01875e-13*ic_cap*ic_cap+-5.75000e-14*ic_cap+1.18000e-11'
+ mcm3m1f_cf_w_0_140_s_0_560 = '-1.34375e-13*ic_cap*ic_cap+-8.75000e-14*ic_cap+1.52000e-11'
+ mcm3m1f_cf_w_0_140_s_0_840 = '-2.00000e-13*ic_cap*ic_cap+-1.25000e-13*ic_cap+2.14000e-11'
+ mcm3m1f_cf_w_0_140_s_1_540 = '-2.93750e-13*ic_cap*ic_cap+-1.75000e-13*ic_cap+3.23000e-11'
+ mcm3m1f_cf_w_0_140_s_3_500 = '-2.75000e-13*ic_cap*ic_cap+-1.75000e-13*ic_cap+4.19000e-11'
+ mcm3m1f_cf_w_1_120_s_0_140 = '-9.68750e-15*ic_cap*ic_cap+-6.25000e-15*ic_cap+4.06000e-12'
+ mcm3m1f_cf_w_1_120_s_0_175 = '-2.15625e-14*ic_cap*ic_cap+-1.37500e-14*ic_cap+5.06000e-12'
+ mcm3m1f_cf_w_1_120_s_0_210 = '-3.37500e-14*ic_cap*ic_cap+-1.75000e-14*ic_cap+6.05000e-12'
+ mcm3m1f_cf_w_1_120_s_0_280 = '-5.43750e-14*ic_cap*ic_cap+-3.50000e-14*ic_cap+7.99000e-12'
+ mcm3m1f_cf_w_1_120_s_0_350 = '-7.81250e-14*ic_cap*ic_cap+-4.50000e-14*ic_cap+9.92000e-12'
+ mcm3m1f_cf_w_1_120_s_0_420 = '-9.78125e-14*ic_cap*ic_cap+-6.62500e-14*ic_cap+1.18000e-11'
+ mcm3m1f_cf_w_1_120_s_0_560 = '-1.40625e-13*ic_cap*ic_cap+-8.75000e-14*ic_cap+1.54000e-11'
+ mcm3m1f_cf_w_1_120_s_0_840 = '-2.00000e-13*ic_cap*ic_cap+-1.25000e-13*ic_cap+2.17000e-11'
+ mcm3m1f_cf_w_1_120_s_1_540 = '-2.90625e-13*ic_cap*ic_cap+-1.87500e-13*ic_cap+3.33000e-11'
+ mcm3m1f_cf_w_1_120_s_3_500 = '-2.50000e-13*ic_cap*ic_cap+-1.75000e-13*ic_cap+4.41000e-11'
+ mcm3m1l1_ca_w_0_140_s_0_140 = '-2.37500e-06*ic_cap*ic_cap+-1.50000e-06*ic_cap+1.47000e-04'
+ mcm3m1l1_ca_w_0_140_s_0_175 = '-2.37500e-06*ic_cap*ic_cap+-1.50000e-06*ic_cap+1.47000e-04'
+ mcm3m1l1_ca_w_0_140_s_0_210 = '-2.37500e-06*ic_cap*ic_cap+-1.50000e-06*ic_cap+1.47000e-04'
+ mcm3m1l1_ca_w_0_140_s_0_280 = '-2.37500e-06*ic_cap*ic_cap+-1.50000e-06*ic_cap+1.47000e-04'
+ mcm3m1l1_ca_w_0_140_s_0_350 = '-2.37500e-06*ic_cap*ic_cap+-1.50000e-06*ic_cap+1.47000e-04'
+ mcm3m1l1_ca_w_0_140_s_0_420 = '-2.37500e-06*ic_cap*ic_cap+-1.50000e-06*ic_cap+1.47000e-04'
+ mcm3m1l1_ca_w_0_140_s_0_560 = '-2.37500e-06*ic_cap*ic_cap+-1.50000e-06*ic_cap+1.47000e-04'
+ mcm3m1l1_ca_w_0_140_s_0_840 = '-2.37500e-06*ic_cap*ic_cap+-1.50000e-06*ic_cap+1.47000e-04'
+ mcm3m1l1_ca_w_0_140_s_1_540 = '-2.37500e-06*ic_cap*ic_cap+-1.50000e-06*ic_cap+1.47000e-04'
+ mcm3m1l1_ca_w_0_140_s_3_500 = '-2.37500e-06*ic_cap*ic_cap+-1.50000e-06*ic_cap+1.47000e-04'
+ mcm3m1l1_ca_w_1_120_s_0_140 = '-2.37500e-06*ic_cap*ic_cap+-1.50000e-06*ic_cap+1.47000e-04'
+ mcm3m1l1_ca_w_1_120_s_0_175 = '-2.37500e-06*ic_cap*ic_cap+-1.50000e-06*ic_cap+1.47000e-04'
+ mcm3m1l1_ca_w_1_120_s_0_210 = '-2.37500e-06*ic_cap*ic_cap+-1.50000e-06*ic_cap+1.47000e-04'
+ mcm3m1l1_ca_w_1_120_s_0_280 = '-2.37500e-06*ic_cap*ic_cap+-1.50000e-06*ic_cap+1.47000e-04'
+ mcm3m1l1_ca_w_1_120_s_0_350 = '-2.37500e-06*ic_cap*ic_cap+-1.50000e-06*ic_cap+1.47000e-04'
+ mcm3m1l1_ca_w_1_120_s_0_420 = '-2.37500e-06*ic_cap*ic_cap+-1.50000e-06*ic_cap+1.47000e-04'
+ mcm3m1l1_ca_w_1_120_s_0_560 = '-2.37500e-06*ic_cap*ic_cap+-1.50000e-06*ic_cap+1.47000e-04'
+ mcm3m1l1_ca_w_1_120_s_0_840 = '-2.37500e-06*ic_cap*ic_cap+-1.50000e-06*ic_cap+1.47000e-04'
+ mcm3m1l1_ca_w_1_120_s_1_540 = '-2.37500e-06*ic_cap*ic_cap+-1.50000e-06*ic_cap+1.47000e-04'
+ mcm3m1l1_ca_w_1_120_s_3_500 = '-2.37500e-06*ic_cap*ic_cap+-1.50000e-06*ic_cap+1.47000e-04'
+ mcm3m1l1_cc_w_0_140_s_0_140 = '-7.56250e-13*ic_cap*ic_cap+-3.00000e-13*ic_cap+9.23000e-11'
+ mcm3m1l1_cc_w_0_140_s_0_175 = '-7.12500e-13*ic_cap*ic_cap+-3.00000e-13*ic_cap+8.99000e-11'
+ mcm3m1l1_cc_w_0_140_s_0_210 = '-5.53125e-13*ic_cap*ic_cap+-3.37500e-13*ic_cap+8.35000e-11'
+ mcm3m1l1_cc_w_0_140_s_0_280 = '-3.59375e-13*ic_cap*ic_cap+-2.37500e-13*ic_cap+7.03000e-11'
+ mcm3m1l1_cc_w_0_140_s_0_350 = '-2.40625e-13*ic_cap*ic_cap+-1.12500e-13*ic_cap+5.81000e-11'
+ mcm3m1l1_cc_w_0_140_s_0_420 = '-1.28125e-13*ic_cap*ic_cap+-3.75000e-14*ic_cap+4.76000e-11'
+ mcm3m1l1_cc_w_0_140_s_0_560 = '9.37500e-15*ic_cap*ic_cap+1.25000e-14*ic_cap+3.32000e-11'
+ mcm3m1l1_cc_w_0_140_s_0_840 = '1.06250e-13*ic_cap*ic_cap+7.50000e-14*ic_cap+1.76000e-11'
+ mcm3m1l1_cc_w_0_140_s_1_540 = '8.43750e-14*ic_cap*ic_cap+6.75000e-14*ic_cap+4.42000e-12'
+ mcm3m1l1_cc_w_0_140_s_3_500 = '5.46875e-15*ic_cap*ic_cap+9.37500e-15*ic_cap+2.10000e-13'
+ mcm3m1l1_cc_w_1_120_s_0_140 = '-5.28125e-13*ic_cap*ic_cap+-4.12500e-13*ic_cap+9.93000e-11'
+ mcm3m1l1_cc_w_1_120_s_0_175 = '-5.84375e-13*ic_cap*ic_cap+-1.62500e-13*ic_cap+9.67000e-11'
+ mcm3m1l1_cc_w_1_120_s_0_210 = '-4.25000e-13*ic_cap*ic_cap+-2.00000e-13*ic_cap+8.96000e-11'
+ mcm3m1l1_cc_w_1_120_s_0_280 = '-2.43750e-13*ic_cap*ic_cap+-1.00000e-13*ic_cap+7.50000e-11'
+ mcm3m1l1_cc_w_1_120_s_0_350 = '-1.37500e-13*ic_cap*ic_cap+-7.50000e-14*ic_cap+6.21000e-11'
+ mcm3m1l1_cc_w_1_120_s_0_420 = '-4.37500e-14*ic_cap*ic_cap+5.11000e-11'
+ mcm3m1l1_cc_w_1_120_s_0_560 = '8.12500e-14*ic_cap*ic_cap+7.50000e-14*ic_cap+3.58000e-11'
+ mcm3m1l1_cc_w_1_120_s_0_840 = '1.53125e-13*ic_cap*ic_cap+1.12500e-13*ic_cap+1.93000e-11'
+ mcm3m1l1_cc_w_1_120_s_1_540 = '1.13750e-13*ic_cap*ic_cap+9.50000e-14*ic_cap+4.97000e-12'
+ mcm3m1l1_cc_w_1_120_s_3_500 = '7.18750e-15*ic_cap*ic_cap+1.12500e-14*ic_cap+2.35000e-13'
+ mcm3m1l1_cf_w_0_140_s_0_140 = '-6.90625e-14*ic_cap*ic_cap+-5.37500e-14*ic_cap+9.69000e-12'
+ mcm3m1l1_cf_w_0_140_s_0_175 = '-1.09375e-13*ic_cap*ic_cap+-8.75000e-14*ic_cap+1.22000e-11'
+ mcm3m1l1_cf_w_0_140_s_0_210 = '-1.43750e-13*ic_cap*ic_cap+-1.00000e-13*ic_cap+1.46000e-11'
+ mcm3m1l1_cf_w_0_140_s_0_280 = '-2.15625e-13*ic_cap*ic_cap+-1.62500e-13*ic_cap+1.92000e-11'
+ mcm3m1l1_cf_w_0_140_s_0_350 = '-2.87500e-13*ic_cap*ic_cap+-2.00000e-13*ic_cap+2.36000e-11'
+ mcm3m1l1_cf_w_0_140_s_0_420 = '-3.43750e-13*ic_cap*ic_cap+-2.25000e-13*ic_cap+2.76000e-11'
+ mcm3m1l1_cf_w_0_140_s_0_560 = '-4.21875e-13*ic_cap*ic_cap+-2.87500e-13*ic_cap+3.45000e-11'
+ mcm3m1l1_cf_w_0_140_s_0_840 = '-5.25000e-13*ic_cap*ic_cap+-3.50000e-13*ic_cap+4.47000e-11'
+ mcm3m1l1_cf_w_0_140_s_1_540 = '-5.62500e-13*ic_cap*ic_cap+-3.75000e-13*ic_cap+5.63000e-11'
+ mcm3m1l1_cf_w_0_140_s_3_500 = '-5.03125e-13*ic_cap*ic_cap+-3.37500e-13*ic_cap+6.09000e-11'
+ mcm3m1l1_cf_w_1_120_s_0_140 = '-6.87500e-14*ic_cap*ic_cap+-5.50000e-14*ic_cap+9.78000e-12'
+ mcm3m1l1_cf_w_1_120_s_0_175 = '-1.09375e-13*ic_cap*ic_cap+-8.75000e-14*ic_cap+1.23000e-11'
+ mcm3m1l1_cf_w_1_120_s_0_210 = '-1.50000e-13*ic_cap*ic_cap+-1.00000e-13*ic_cap+1.47000e-11'
+ mcm3m1l1_cf_w_1_120_s_0_280 = '-2.15625e-13*ic_cap*ic_cap+-1.62500e-13*ic_cap+1.93000e-11'
+ mcm3m1l1_cf_w_1_120_s_0_350 = '-2.78125e-13*ic_cap*ic_cap+-1.87500e-13*ic_cap+2.36000e-11'
+ mcm3m1l1_cf_w_1_120_s_0_420 = '-3.34375e-13*ic_cap*ic_cap+-2.37500e-13*ic_cap+2.76000e-11'
+ mcm3m1l1_cf_w_1_120_s_0_560 = '-4.25000e-13*ic_cap*ic_cap+-2.75000e-13*ic_cap+3.47000e-11'
+ mcm3m1l1_cf_w_1_120_s_0_840 = '-5.25000e-13*ic_cap*ic_cap+-3.50000e-13*ic_cap+4.52000e-11'
+ mcm3m1l1_cf_w_1_120_s_1_540 = '-5.50000e-13*ic_cap*ic_cap+-3.75000e-13*ic_cap+5.75000e-11'
+ mcm3m1l1_cf_w_1_120_s_3_500 = '-4.71875e-13*ic_cap*ic_cap+-3.12500e-13*ic_cap+6.25000e-11'
+ mcm3m1p1_ca_w_0_140_s_0_140 = '-1.07500e-06*ic_cap*ic_cap+-6.25000e-07*ic_cap+7.78000e-05'
+ mcm3m1p1_ca_w_0_140_s_0_175 = '-1.07500e-06*ic_cap*ic_cap+-6.25000e-07*ic_cap+7.78000e-05'
+ mcm3m1p1_ca_w_0_140_s_0_210 = '-1.07500e-06*ic_cap*ic_cap+-6.25000e-07*ic_cap+7.78000e-05'
+ mcm3m1p1_ca_w_0_140_s_0_280 = '-1.07500e-06*ic_cap*ic_cap+-6.25000e-07*ic_cap+7.78000e-05'
+ mcm3m1p1_ca_w_0_140_s_0_350 = '-1.07500e-06*ic_cap*ic_cap+-6.25000e-07*ic_cap+7.78000e-05'
+ mcm3m1p1_ca_w_0_140_s_0_420 = '-1.07500e-06*ic_cap*ic_cap+-6.25000e-07*ic_cap+7.78000e-05'
+ mcm3m1p1_ca_w_0_140_s_0_560 = '-1.07500e-06*ic_cap*ic_cap+-6.25000e-07*ic_cap+7.78000e-05'
+ mcm3m1p1_ca_w_0_140_s_0_840 = '-1.07500e-06*ic_cap*ic_cap+-6.25000e-07*ic_cap+7.78000e-05'
+ mcm3m1p1_ca_w_0_140_s_1_540 = '-1.07500e-06*ic_cap*ic_cap+-6.25000e-07*ic_cap+7.78000e-05'
+ mcm3m1p1_ca_w_0_140_s_3_500 = '-1.07500e-06*ic_cap*ic_cap+-6.25000e-07*ic_cap+7.78000e-05'
+ mcm3m1p1_ca_w_1_120_s_0_140 = '-1.07500e-06*ic_cap*ic_cap+-6.25000e-07*ic_cap+7.78000e-05'
+ mcm3m1p1_ca_w_1_120_s_0_175 = '-1.07500e-06*ic_cap*ic_cap+-6.25000e-07*ic_cap+7.78000e-05'
+ mcm3m1p1_ca_w_1_120_s_0_210 = '-1.07500e-06*ic_cap*ic_cap+-6.25000e-07*ic_cap+7.78000e-05'
+ mcm3m1p1_ca_w_1_120_s_0_280 = '-1.07500e-06*ic_cap*ic_cap+-6.25000e-07*ic_cap+7.78000e-05'
+ mcm3m1p1_ca_w_1_120_s_0_350 = '-1.07500e-06*ic_cap*ic_cap+-6.25000e-07*ic_cap+7.78000e-05'
+ mcm3m1p1_ca_w_1_120_s_0_420 = '-1.07500e-06*ic_cap*ic_cap+-6.25000e-07*ic_cap+7.78000e-05'
+ mcm3m1p1_ca_w_1_120_s_0_560 = '-1.07500e-06*ic_cap*ic_cap+-6.25000e-07*ic_cap+7.78000e-05'
+ mcm3m1p1_ca_w_1_120_s_0_840 = '-1.07500e-06*ic_cap*ic_cap+-6.25000e-07*ic_cap+7.78000e-05'
+ mcm3m1p1_ca_w_1_120_s_1_540 = '-1.07500e-06*ic_cap*ic_cap+-6.25000e-07*ic_cap+7.78000e-05'
+ mcm3m1p1_ca_w_1_120_s_3_500 = '-1.07500e-06*ic_cap*ic_cap+-6.25000e-07*ic_cap+7.78000e-05'
+ mcm3m1p1_cc_w_0_140_s_0_140 = '-8.37500e-13*ic_cap*ic_cap+-5.25000e-13*ic_cap+9.86000e-11'
+ mcm3m1p1_cc_w_0_140_s_0_175 = '-7.78125e-13*ic_cap*ic_cap+-5.37500e-13*ic_cap+9.67000e-11'
+ mcm3m1p1_cc_w_0_140_s_0_210 = '-6.34375e-13*ic_cap*ic_cap+-3.87500e-13*ic_cap+9.06000e-11'
+ mcm3m1p1_cc_w_0_140_s_0_280 = '-4.59375e-13*ic_cap*ic_cap+-3.37500e-13*ic_cap+7.85000e-11'
+ mcm3m1p1_cc_w_0_140_s_0_350 = '-3.25000e-13*ic_cap*ic_cap+-2.25000e-13*ic_cap+6.65000e-11'
+ mcm3m1p1_cc_w_0_140_s_0_420 = '-2.09375e-13*ic_cap*ic_cap+-1.87500e-13*ic_cap+5.61000e-11'
+ mcm3m1p1_cc_w_0_140_s_0_560 = '-5.93750e-14*ic_cap*ic_cap+-6.25000e-14*ic_cap+4.20000e-11'
+ mcm3m1p1_cc_w_0_140_s_0_840 = '6.87500e-14*ic_cap*ic_cap+2.50000e-14*ic_cap+2.56000e-11'
+ mcm3m1p1_cc_w_0_140_s_1_540 = '1.19375e-13*ic_cap*ic_cap+7.50000e-14*ic_cap+8.79000e-12'
+ mcm3m1p1_cc_w_0_140_s_3_500 = '3.09375e-14*ic_cap*ic_cap+2.62500e-14*ic_cap+5.90000e-13'
+ mcm3m1p1_cc_w_1_120_s_0_140 = '-5.87500e-13*ic_cap*ic_cap+-3.50000e-13*ic_cap+1.10000e-10'
+ mcm3m1p1_cc_w_1_120_s_0_175 = '-6.03125e-13*ic_cap*ic_cap+-2.87500e-13*ic_cap+1.07000e-10'
+ mcm3m1p1_cc_w_1_120_s_0_210 = '-4.46875e-13*ic_cap*ic_cap+-2.62500e-13*ic_cap+9.98000e-11'
+ mcm3m1p1_cc_w_1_120_s_0_280 = '-2.65625e-13*ic_cap*ic_cap+-1.87500e-13*ic_cap+8.54000e-11'
+ mcm3m1p1_cc_w_1_120_s_0_350 = '-1.68750e-13*ic_cap*ic_cap+-1.00000e-13*ic_cap+7.26000e-11'
+ mcm3m1p1_cc_w_1_120_s_0_420 = '-5.93750e-14*ic_cap*ic_cap+-8.75000e-14*ic_cap+6.14000e-11'
+ mcm3m1p1_cc_w_1_120_s_0_560 = '5.62500e-14*ic_cap*ic_cap+2.50000e-14*ic_cap+4.58000e-11'
+ mcm3m1p1_cc_w_1_120_s_0_840 = '1.46875e-13*ic_cap*ic_cap+8.75000e-14*ic_cap+2.81000e-11'
+ mcm3m1p1_cc_w_1_120_s_1_540 = '1.67500e-13*ic_cap*ic_cap+1.12500e-13*ic_cap+9.77000e-12'
+ mcm3m1p1_cc_w_1_120_s_3_500 = '4.03125e-14*ic_cap*ic_cap+3.00000e-14*ic_cap+6.25000e-13'
+ mcm3m1p1_cf_w_0_140_s_0_140 = '-2.59375e-14*ic_cap*ic_cap+-1.62500e-14*ic_cap+5.34000e-12'
+ mcm3m1p1_cf_w_0_140_s_0_175 = '-4.43750e-14*ic_cap*ic_cap+-2.75000e-14*ic_cap+6.66000e-12'
+ mcm3m1p1_cf_w_0_140_s_0_210 = '-6.03125e-14*ic_cap*ic_cap+-3.87500e-14*ic_cap+7.99000e-12'
+ mcm3m1p1_cf_w_0_140_s_0_280 = '-9.37500e-14*ic_cap*ic_cap+-6.00000e-14*ic_cap+1.05000e-11'
+ mcm3m1p1_cf_w_0_140_s_0_350 = '-1.28125e-13*ic_cap*ic_cap+-8.75000e-14*ic_cap+1.30000e-11'
+ mcm3m1p1_cf_w_0_140_s_0_420 = '-1.59375e-13*ic_cap*ic_cap+-8.75000e-14*ic_cap+1.54000e-11'
+ mcm3m1p1_cf_w_0_140_s_0_560 = '-2.15625e-13*ic_cap*ic_cap+-1.37500e-13*ic_cap+1.99000e-11'
+ mcm3m1p1_cf_w_0_140_s_0_840 = '-3.03125e-13*ic_cap*ic_cap+-1.87500e-13*ic_cap+2.75000e-11'
+ mcm3m1p1_cf_w_0_140_s_1_540 = '-3.84375e-13*ic_cap*ic_cap+-2.37500e-13*ic_cap+3.93000e-11'
+ mcm3m1p1_cf_w_0_140_s_3_500 = '-3.34375e-13*ic_cap*ic_cap+-2.12500e-13*ic_cap+4.72000e-11'
+ mcm3m1p1_cf_w_1_120_s_0_140 = '-2.71875e-14*ic_cap*ic_cap+-1.87500e-14*ic_cap+5.45000e-12'
+ mcm3m1p1_cf_w_1_120_s_0_175 = '-4.46875e-14*ic_cap*ic_cap+-3.12500e-14*ic_cap+6.77000e-12'
+ mcm3m1p1_cf_w_1_120_s_0_210 = '-6.40625e-14*ic_cap*ic_cap+-3.87500e-14*ic_cap+8.09000e-12'
+ mcm3m1p1_cf_w_1_120_s_0_280 = '-9.40625e-14*ic_cap*ic_cap+-6.12500e-14*ic_cap+1.06000e-11'
+ mcm3m1p1_cf_w_1_120_s_0_350 = '-1.34375e-13*ic_cap*ic_cap+-8.75000e-14*ic_cap+1.32000e-11'
+ mcm3m1p1_cf_w_1_120_s_0_420 = '-1.62500e-13*ic_cap*ic_cap+-1.00000e-13*ic_cap+1.56000e-11'
+ mcm3m1p1_cf_w_1_120_s_0_560 = '-2.18750e-13*ic_cap*ic_cap+-1.25000e-13*ic_cap+2.01000e-11'
+ mcm3m1p1_cf_w_1_120_s_0_840 = '-3.03125e-13*ic_cap*ic_cap+-1.87500e-13*ic_cap+2.79000e-11'
+ mcm3m1p1_cf_w_1_120_s_1_540 = '-3.87500e-13*ic_cap*ic_cap+-2.50000e-13*ic_cap+4.05000e-11'
+ mcm3m1p1_cf_w_1_120_s_3_500 = '-3.00000e-13*ic_cap*ic_cap+-2.00000e-13*ic_cap+4.89000e-11'
+ mcm3m2_ca_w_0_300_s_0_300 = '-1.25000e-06*ic_cap*ic_cap+-6.75000e-07*ic_cap+8.22000e-05'
+ mcm3m2_ca_w_0_300_s_0_360 = '-1.25000e-06*ic_cap*ic_cap+-6.75000e-07*ic_cap+8.22000e-05'
+ mcm3m2_ca_w_0_300_s_0_450 = '-1.25000e-06*ic_cap*ic_cap+-6.75000e-07*ic_cap+8.22000e-05'
+ mcm3m2_ca_w_0_300_s_0_600 = '-1.25000e-06*ic_cap*ic_cap+-6.75000e-07*ic_cap+8.22000e-05'
+ mcm3m2_ca_w_0_300_s_0_800 = '-1.25000e-06*ic_cap*ic_cap+-6.75000e-07*ic_cap+8.22000e-05'
+ mcm3m2_ca_w_0_300_s_1_000 = '-1.25000e-06*ic_cap*ic_cap+-6.75000e-07*ic_cap+8.22000e-05'
+ mcm3m2_ca_w_0_300_s_1_200 = '-1.25000e-06*ic_cap*ic_cap+-6.75000e-07*ic_cap+8.22000e-05'
+ mcm3m2_ca_w_0_300_s_2_100 = '-1.25000e-06*ic_cap*ic_cap+-6.75000e-07*ic_cap+8.22000e-05'
+ mcm3m2_ca_w_0_300_s_3_300 = '-1.25000e-06*ic_cap*ic_cap+-6.75000e-07*ic_cap+8.22000e-05'
+ mcm3m2_ca_w_0_300_s_9_000 = '-1.25000e-06*ic_cap*ic_cap+-6.75000e-07*ic_cap+8.22000e-05'
+ mcm3m2_ca_w_2_400_s_0_300 = '-1.25000e-06*ic_cap*ic_cap+-6.75000e-07*ic_cap+8.22000e-05'
+ mcm3m2_ca_w_2_400_s_0_360 = '-1.25000e-06*ic_cap*ic_cap+-6.75000e-07*ic_cap+8.22000e-05'
+ mcm3m2_ca_w_2_400_s_0_450 = '-1.25000e-06*ic_cap*ic_cap+-6.75000e-07*ic_cap+8.22000e-05'
+ mcm3m2_ca_w_2_400_s_0_600 = '-1.25000e-06*ic_cap*ic_cap+-6.75000e-07*ic_cap+8.22000e-05'
+ mcm3m2_ca_w_2_400_s_0_800 = '-1.25000e-06*ic_cap*ic_cap+-6.75000e-07*ic_cap+8.22000e-05'
+ mcm3m2_ca_w_2_400_s_1_000 = '-1.25000e-06*ic_cap*ic_cap+-6.75000e-07*ic_cap+8.22000e-05'
+ mcm3m2_ca_w_2_400_s_1_200 = '-1.25000e-06*ic_cap*ic_cap+-6.75000e-07*ic_cap+8.22000e-05'
+ mcm3m2_ca_w_2_400_s_2_100 = '-1.25000e-06*ic_cap*ic_cap+-6.75000e-07*ic_cap+8.22000e-05'
+ mcm3m2_ca_w_2_400_s_3_300 = '-1.25000e-06*ic_cap*ic_cap+-6.75000e-07*ic_cap+8.22000e-05'
+ mcm3m2_ca_w_2_400_s_9_000 = '-1.25000e-06*ic_cap*ic_cap+-6.75000e-07*ic_cap+8.22000e-05'
+ mcm3m2_cc_w_0_300_s_0_300 = '-6.65625e-13*ic_cap*ic_cap+-3.62500e-13*ic_cap+9.39000e-11'
+ mcm3m2_cc_w_0_300_s_0_360 = '-5.59375e-13*ic_cap*ic_cap+-3.12500e-13*ic_cap+8.63000e-11'
+ mcm3m2_cc_w_0_300_s_0_450 = '-4.50000e-13*ic_cap*ic_cap+-2.75000e-13*ic_cap+7.63000e-11'
+ mcm3m2_cc_w_0_300_s_0_600 = '-3.15625e-13*ic_cap*ic_cap+-1.87500e-13*ic_cap+6.30000e-11'
+ mcm3m2_cc_w_0_300_s_0_800 = '-1.93750e-13*ic_cap*ic_cap+-1.50000e-13*ic_cap+5.03000e-11'
+ mcm3m2_cc_w_0_300_s_1_000 = '-1.25000e-13*ic_cap*ic_cap+-1.00000e-13*ic_cap+4.10000e-11'
+ mcm3m2_cc_w_0_300_s_1_200 = '-8.75000e-14*ic_cap*ic_cap+-7.50000e-14*ic_cap+3.42000e-11'
+ mcm3m2_cc_w_0_300_s_2_100 = '-1.56250e-14*ic_cap*ic_cap+-1.25000e-14*ic_cap+1.76000e-11'
+ mcm3m2_cc_w_0_300_s_9_000 = '3.12500e-15*ic_cap*ic_cap+1.95000e-12'
+ mcm3m2_cc_w_2_400_s_0_300 = '-6.40625e-13*ic_cap*ic_cap+-3.12500e-13*ic_cap+1.11000e-10'
+ mcm3m2_cc_w_2_400_s_0_360 = '-5.40625e-13*ic_cap*ic_cap+-2.87500e-13*ic_cap+1.03000e-10'
+ mcm3m2_cc_w_2_400_s_0_450 = '-4.25000e-13*ic_cap*ic_cap+-2.50000e-13*ic_cap+9.20000e-11'
+ mcm3m2_cc_w_2_400_s_0_600 = '-2.96875e-13*ic_cap*ic_cap+-1.62500e-13*ic_cap+7.76000e-11'
+ mcm3m2_cc_w_2_400_s_0_800 = '-1.75000e-13*ic_cap*ic_cap+-1.25000e-13*ic_cap+6.33000e-11'
+ mcm3m2_cc_w_2_400_s_1_000 = '-1.18750e-13*ic_cap*ic_cap+-1.00000e-13*ic_cap+5.31000e-11'
+ mcm3m2_cc_w_2_400_s_1_200 = '-7.81250e-14*ic_cap*ic_cap+-6.25000e-14*ic_cap+4.56000e-11'
+ mcm3m2_cc_w_2_400_s_2_100 = '-9.37500e-15*ic_cap*ic_cap+-1.25000e-14*ic_cap+2.72000e-11'
+ mcm3m2_cc_w_2_400_s_3_300 = '6.25000e-15*ic_cap*ic_cap+1.68000e-11'
+ mcm3m2_cc_w_2_400_s_9_000 = '4.68750e-15*ic_cap*ic_cap+6.25000e-15*ic_cap+4.25000e-12'
+ mcm3m2_cf_w_0_300_s_0_300 = '-9.21875e-14*ic_cap*ic_cap+-4.87500e-14*ic_cap+1.11000e-11'
+ mcm3m2_cf_w_0_300_s_0_360 = '-1.15625e-13*ic_cap*ic_cap+-6.25000e-14*ic_cap+1.30000e-11'
+ mcm3m2_cf_w_0_300_s_0_450 = '-1.50000e-13*ic_cap*ic_cap+-7.50000e-14*ic_cap+1.57000e-11'
+ mcm3m2_cf_w_0_300_s_0_600 = '-1.96875e-13*ic_cap*ic_cap+-1.12500e-13*ic_cap+1.99000e-11'
+ mcm3m2_cf_w_0_300_s_0_800 = '-2.46875e-13*ic_cap*ic_cap+-1.37500e-13*ic_cap+2.45000e-11'
+ mcm3m2_cf_w_0_300_s_1_000 = '-2.78125e-13*ic_cap*ic_cap+-1.62500e-13*ic_cap+2.85000e-11'
+ mcm3m2_cf_w_0_300_s_1_200 = '-3.03125e-13*ic_cap*ic_cap+-1.87500e-13*ic_cap+3.19000e-11'
+ mcm3m2_cf_w_0_300_s_2_100 = '-3.62500e-13*ic_cap*ic_cap+-2.25000e-13*ic_cap+4.31000e-11'
+ mcm3m2_cf_w_0_300_s_3_300 = '-3.75000e-13*ic_cap*ic_cap+-2.25000e-13*ic_cap+4.95000e-11'
+ mcm3m2_cf_w_0_300_s_9_000 = '-3.84375e-13*ic_cap*ic_cap+-2.37500e-13*ic_cap+5.72000e-11'
+ mcm3m2_cf_w_2_400_s_0_300 = '-9.09375e-14*ic_cap*ic_cap+-4.87500e-14*ic_cap+1.11000e-11'
+ mcm3m2_cf_w_2_400_s_0_360 = '-1.15625e-13*ic_cap*ic_cap+-6.25000e-14*ic_cap+1.30000e-11'
+ mcm3m2_cf_w_2_400_s_0_450 = '-1.46875e-13*ic_cap*ic_cap+-8.75000e-14*ic_cap+1.57000e-11'
+ mcm3m2_cf_w_2_400_s_0_600 = '-1.96875e-13*ic_cap*ic_cap+-1.12500e-13*ic_cap+1.98000e-11'
+ mcm3m2_cf_w_2_400_s_0_800 = '-2.40625e-13*ic_cap*ic_cap+-1.37500e-13*ic_cap+2.45000e-11'
+ mcm3m2_cf_w_2_400_s_1_000 = '-2.81250e-13*ic_cap*ic_cap+-1.50000e-13*ic_cap+2.86000e-11'
+ mcm3m2_cf_w_2_400_s_1_200 = '-3.00000e-13*ic_cap*ic_cap+-1.75000e-13*ic_cap+3.20000e-11'
+ mcm3m2_cf_w_2_400_s_2_100 = '-3.46875e-13*ic_cap*ic_cap+-2.12500e-13*ic_cap+4.29000e-11'
+ mcm3m2_cf_w_2_400_s_3_300 = '-3.71875e-13*ic_cap*ic_cap+-2.12500e-13*ic_cap+5.12000e-11'
+ mcm3m2_cf_w_2_400_s_9_000 = '-3.75000e-13*ic_cap*ic_cap+-2.25000e-13*ic_cap+6.29000e-11'
+ mcm3m2d_ca_w_0_140_s_0_140 = '-1.46563e-06*ic_cap*ic_cap+-8.12500e-07*ic_cap+1.03000e-04'
+ mcm3m2d_ca_w_0_140_s_0_175 = '-1.46563e-06*ic_cap*ic_cap+-8.12500e-07*ic_cap+1.03000e-04'
+ mcm3m2d_ca_w_0_140_s_0_210 = '-1.46563e-06*ic_cap*ic_cap+-8.12500e-07*ic_cap+1.03000e-04'
+ mcm3m2d_ca_w_0_140_s_0_280 = '-1.46563e-06*ic_cap*ic_cap+-8.12500e-07*ic_cap+1.03000e-04'
+ mcm3m2d_ca_w_0_140_s_0_350 = '-1.46563e-06*ic_cap*ic_cap+-8.12500e-07*ic_cap+1.03000e-04'
+ mcm3m2d_ca_w_0_140_s_0_420 = '-1.46563e-06*ic_cap*ic_cap+-8.12500e-07*ic_cap+1.03000e-04'
+ mcm3m2d_ca_w_0_140_s_0_560 = '-1.46563e-06*ic_cap*ic_cap+-8.12500e-07*ic_cap+1.03000e-04'
+ mcm3m2d_ca_w_0_140_s_0_840 = '-1.46563e-06*ic_cap*ic_cap+-8.12500e-07*ic_cap+1.03000e-04'
+ mcm3m2d_ca_w_0_140_s_1_540 = '-1.46563e-06*ic_cap*ic_cap+-8.12500e-07*ic_cap+1.03000e-04'
+ mcm3m2d_ca_w_0_140_s_3_500 = '-1.46563e-06*ic_cap*ic_cap+-8.12500e-07*ic_cap+1.03000e-04'
+ mcm3m2d_ca_w_1_120_s_0_140 = '-1.46563e-06*ic_cap*ic_cap+-8.12500e-07*ic_cap+1.03000e-04'
+ mcm3m2d_ca_w_1_120_s_0_175 = '-1.46563e-06*ic_cap*ic_cap+-8.12500e-07*ic_cap+1.03000e-04'
+ mcm3m2d_ca_w_1_120_s_0_210 = '-1.46563e-06*ic_cap*ic_cap+-8.12500e-07*ic_cap+1.03000e-04'
+ mcm3m2d_ca_w_1_120_s_0_280 = '-1.46563e-06*ic_cap*ic_cap+-8.12500e-07*ic_cap+1.03000e-04'
+ mcm3m2d_ca_w_1_120_s_0_350 = '-1.46563e-06*ic_cap*ic_cap+-8.12500e-07*ic_cap+1.03000e-04'
+ mcm3m2d_ca_w_1_120_s_0_420 = '-1.46563e-06*ic_cap*ic_cap+-8.12500e-07*ic_cap+1.03000e-04'
+ mcm3m2d_ca_w_1_120_s_0_560 = '-1.46563e-06*ic_cap*ic_cap+-8.12500e-07*ic_cap+1.03000e-04'
+ mcm3m2d_ca_w_1_120_s_0_840 = '-1.46563e-06*ic_cap*ic_cap+-8.12500e-07*ic_cap+1.03000e-04'
+ mcm3m2d_ca_w_1_120_s_1_540 = '-1.46563e-06*ic_cap*ic_cap+-8.12500e-07*ic_cap+1.03000e-04'
+ mcm3m2d_ca_w_1_120_s_3_500 = '-1.46563e-06*ic_cap*ic_cap+-8.12500e-07*ic_cap+1.03000e-04'
+ mcm3m2d_cc_w_0_140_s_0_140 = '-7.65625e-13*ic_cap*ic_cap+-4.12500e-13*ic_cap+9.60000e-11'
+ mcm3m2d_cc_w_0_140_s_0_175 = '-7.46875e-13*ic_cap*ic_cap+-3.62500e-13*ic_cap+9.41000e-11'
+ mcm3m2d_cc_w_0_140_s_0_210 = '-6.25000e-13*ic_cap*ic_cap+-4.00000e-13*ic_cap+8.84000e-11'
+ mcm3m2d_cc_w_0_140_s_0_280 = '-4.31250e-13*ic_cap*ic_cap+-3.50000e-13*ic_cap+7.58000e-11'
+ mcm3m2d_cc_w_0_140_s_0_350 = '-3.18750e-13*ic_cap*ic_cap+-2.50000e-13*ic_cap+6.40000e-11'
+ mcm3m2d_cc_w_0_140_s_0_420 = '-2.03125e-13*ic_cap*ic_cap+-1.37500e-13*ic_cap+5.36000e-11'
+ mcm3m2d_cc_w_0_140_s_0_560 = '-6.56250e-14*ic_cap*ic_cap+-6.25000e-14*ic_cap+3.96000e-11'
+ mcm3m2d_cc_w_0_140_s_0_840 = '5.31250e-14*ic_cap*ic_cap+1.25000e-14*ic_cap+2.37000e-11'
+ mcm3m2d_cc_w_0_140_s_1_540 = '8.34375e-14*ic_cap*ic_cap+5.12500e-14*ic_cap+8.11000e-12'
+ mcm3m2d_cc_w_0_140_s_3_500 = '2.26563e-14*ic_cap*ic_cap+1.68750e-14*ic_cap+6.60000e-13'
+ mcm3m2d_cc_w_1_120_s_0_140 = '-6.09375e-13*ic_cap*ic_cap+-3.62500e-13*ic_cap+1.07000e-10'
+ mcm3m2d_cc_w_1_120_s_0_175 = '-6.65625e-13*ic_cap*ic_cap+-2.87500e-13*ic_cap+1.05000e-10'
+ mcm3m2d_cc_w_1_120_s_0_210 = '-4.87500e-13*ic_cap*ic_cap+-2.75000e-13*ic_cap+9.73000e-11'
+ mcm3m2d_cc_w_1_120_s_0_280 = '-3.21875e-13*ic_cap*ic_cap+-1.87500e-13*ic_cap+8.32000e-11'
+ mcm3m2d_cc_w_1_120_s_0_350 = '-2.06250e-13*ic_cap*ic_cap+-1.50000e-13*ic_cap+7.03000e-11'
+ mcm3m2d_cc_w_1_120_s_0_420 = '-1.03125e-13*ic_cap*ic_cap+-8.75000e-14*ic_cap+5.93000e-11'
+ mcm3m2d_cc_w_1_120_s_0_560 = '3.12500e-14*ic_cap*ic_cap+4.37000e-11'
+ mcm3m2d_cc_w_1_120_s_0_840 = '1.06250e-13*ic_cap*ic_cap+7.50000e-14*ic_cap+2.66000e-11'
+ mcm3m2d_cc_w_1_120_s_1_540 = '1.25625e-13*ic_cap*ic_cap+7.50000e-14*ic_cap+9.39000e-12'
+ mcm3m2d_cc_w_1_120_s_3_500 = '3.46875e-14*ic_cap*ic_cap+2.87500e-14*ic_cap+7.50000e-13'
+ mcm3m2d_cf_w_0_140_s_0_140 = '-3.62500e-14*ic_cap*ic_cap+-2.00000e-14*ic_cap+6.81000e-12'
+ mcm3m2d_cf_w_0_140_s_0_175 = '-5.78125e-14*ic_cap*ic_cap+-3.12500e-14*ic_cap+8.42000e-12'
+ mcm3m2d_cf_w_0_140_s_0_210 = '-7.59375e-14*ic_cap*ic_cap+-4.12500e-14*ic_cap+1.00000e-11'
+ mcm3m2d_cf_w_0_140_s_0_280 = '-1.15625e-13*ic_cap*ic_cap+-6.25000e-14*ic_cap+1.30000e-11'
+ mcm3m2d_cf_w_0_140_s_0_350 = '-1.53125e-13*ic_cap*ic_cap+-8.75000e-14*ic_cap+1.60000e-11'
+ mcm3m2d_cf_w_0_140_s_0_420 = '-1.90625e-13*ic_cap*ic_cap+-1.12500e-13*ic_cap+1.89000e-11'
+ mcm3m2d_cf_w_0_140_s_0_560 = '-2.46875e-13*ic_cap*ic_cap+-1.37500e-13*ic_cap+2.39000e-11'
+ mcm3m2d_cf_w_0_140_s_0_840 = '-3.25000e-13*ic_cap*ic_cap+-2.00000e-13*ic_cap+3.21000e-11'
+ mcm3m2d_cf_w_0_140_s_1_540 = '-3.90625e-13*ic_cap*ic_cap+-2.37500e-13*ic_cap+4.38000e-11'
+ mcm3m2d_cf_w_0_140_s_3_500 = '-3.40625e-13*ic_cap*ic_cap+-2.12500e-13*ic_cap+5.08000e-11'
+ mcm3m2d_cf_w_1_120_s_0_140 = '-3.59375e-14*ic_cap*ic_cap+-1.87500e-14*ic_cap+6.85000e-12'
+ mcm3m2d_cf_w_1_120_s_0_175 = '-5.78125e-14*ic_cap*ic_cap+-3.37500e-14*ic_cap+8.48000e-12'
+ mcm3m2d_cf_w_1_120_s_0_210 = '-7.50000e-14*ic_cap*ic_cap+-4.25000e-14*ic_cap+1.00000e-11'
+ mcm3m2d_cf_w_1_120_s_0_280 = '-1.15625e-13*ic_cap*ic_cap+-6.25000e-14*ic_cap+1.31000e-11'
+ mcm3m2d_cf_w_1_120_s_0_350 = '-1.53125e-13*ic_cap*ic_cap+-8.75000e-14*ic_cap+1.61000e-11'
+ mcm3m2d_cf_w_1_120_s_0_420 = '-1.81250e-13*ic_cap*ic_cap+-1.00000e-13*ic_cap+1.89000e-11'
+ mcm3m2d_cf_w_1_120_s_0_560 = '-2.43750e-13*ic_cap*ic_cap+-1.50000e-13*ic_cap+2.41000e-11'
+ mcm3m2d_cf_w_1_120_s_0_840 = '-3.21875e-13*ic_cap*ic_cap+-1.87500e-13*ic_cap+3.25000e-11'
+ mcm3m2d_cf_w_1_120_s_1_540 = '-3.75000e-13*ic_cap*ic_cap+-2.25000e-13*ic_cap+4.48000e-11'
+ mcm3m2d_cf_w_1_120_s_3_500 = '-3.12500e-13*ic_cap*ic_cap+-2.00000e-13*ic_cap+5.30000e-11'
+ mcm3m2f_ca_w_0_140_s_0_140 = '-1.45000e-06*ic_cap*ic_cap+-8.00000e-07*ic_cap+9.98000e-05'
+ mcm3m2f_ca_w_0_140_s_0_175 = '-1.45000e-06*ic_cap*ic_cap+-8.00000e-07*ic_cap+9.98000e-05'
+ mcm3m2f_ca_w_0_140_s_0_210 = '-1.45000e-06*ic_cap*ic_cap+-8.00000e-07*ic_cap+9.98000e-05'
+ mcm3m2f_ca_w_0_140_s_0_280 = '-1.45000e-06*ic_cap*ic_cap+-8.00000e-07*ic_cap+9.98000e-05'
+ mcm3m2f_ca_w_0_140_s_0_350 = '-1.45000e-06*ic_cap*ic_cap+-8.00000e-07*ic_cap+9.98000e-05'
+ mcm3m2f_ca_w_0_140_s_0_420 = '-1.45000e-06*ic_cap*ic_cap+-8.00000e-07*ic_cap+9.98000e-05'
+ mcm3m2f_ca_w_0_140_s_0_560 = '-1.45000e-06*ic_cap*ic_cap+-8.00000e-07*ic_cap+9.98000e-05'
+ mcm3m2f_ca_w_0_140_s_0_840 = '-1.45000e-06*ic_cap*ic_cap+-8.00000e-07*ic_cap+9.98000e-05'
+ mcm3m2f_ca_w_0_140_s_1_540 = '-1.45000e-06*ic_cap*ic_cap+-8.00000e-07*ic_cap+9.98000e-05'
+ mcm3m2f_ca_w_0_140_s_3_500 = '-1.45000e-06*ic_cap*ic_cap+-8.00000e-07*ic_cap+9.98000e-05'
+ mcm3m2f_ca_w_1_120_s_0_140 = '-1.45000e-06*ic_cap*ic_cap+-8.00000e-07*ic_cap+9.98000e-05'
+ mcm3m2f_ca_w_1_120_s_0_175 = '-1.45000e-06*ic_cap*ic_cap+-8.00000e-07*ic_cap+9.98000e-05'
+ mcm3m2f_ca_w_1_120_s_0_210 = '-1.45000e-06*ic_cap*ic_cap+-8.00000e-07*ic_cap+9.98000e-05'
+ mcm3m2f_ca_w_1_120_s_0_280 = '-1.45000e-06*ic_cap*ic_cap+-8.00000e-07*ic_cap+9.98000e-05'
+ mcm3m2f_ca_w_1_120_s_0_350 = '-1.45000e-06*ic_cap*ic_cap+-8.00000e-07*ic_cap+9.98000e-05'
+ mcm3m2f_ca_w_1_120_s_0_420 = '-1.45000e-06*ic_cap*ic_cap+-8.00000e-07*ic_cap+9.98000e-05'
+ mcm3m2f_ca_w_1_120_s_0_560 = '-1.45000e-06*ic_cap*ic_cap+-8.00000e-07*ic_cap+9.98000e-05'
+ mcm3m2f_ca_w_1_120_s_0_840 = '-1.45000e-06*ic_cap*ic_cap+-8.00000e-07*ic_cap+9.98000e-05'
+ mcm3m2f_ca_w_1_120_s_1_540 = '-1.45000e-06*ic_cap*ic_cap+-8.00000e-07*ic_cap+9.98000e-05'
+ mcm3m2f_ca_w_1_120_s_3_500 = '-1.45000e-06*ic_cap*ic_cap+-8.00000e-07*ic_cap+9.98000e-05'
+ mcm3m2f_cc_w_0_140_s_0_140 = '-7.75000e-13*ic_cap*ic_cap+-3.75000e-13*ic_cap+9.63000e-11'
+ mcm3m2f_cc_w_0_140_s_0_175 = '-7.34375e-13*ic_cap*ic_cap+-4.12500e-13*ic_cap+9.45000e-11'
+ mcm3m2f_cc_w_0_140_s_0_210 = '-6.25000e-13*ic_cap*ic_cap+-4.25000e-13*ic_cap+8.87000e-11'
+ mcm3m2f_cc_w_0_140_s_0_280 = '-4.37500e-13*ic_cap*ic_cap+-3.50000e-13*ic_cap+7.64000e-11'
+ mcm3m2f_cc_w_0_140_s_0_350 = '-3.18750e-13*ic_cap*ic_cap+-2.75000e-13*ic_cap+6.46000e-11'
+ mcm3m2f_cc_w_0_140_s_0_420 = '-2.09375e-13*ic_cap*ic_cap+-1.12500e-13*ic_cap+5.44000e-11'
+ mcm3m2f_cc_w_0_140_s_0_560 = '-6.87500e-14*ic_cap*ic_cap+-5.00000e-14*ic_cap+4.04000e-11'
+ mcm3m2f_cc_w_0_140_s_0_840 = '4.06250e-14*ic_cap*ic_cap+3.75000e-14*ic_cap+2.47000e-11'
+ mcm3m2f_cc_w_0_140_s_1_540 = '8.25000e-14*ic_cap*ic_cap+5.00000e-14*ic_cap+8.98000e-12'
+ mcm3m2f_cc_w_0_140_s_3_500 = '2.87500e-14*ic_cap*ic_cap+2.12500e-14*ic_cap+8.85000e-13'
+ mcm3m2f_cc_w_1_120_s_0_140 = '-6.00000e-13*ic_cap*ic_cap+-3.75000e-13*ic_cap+1.08000e-10'
+ mcm3m2f_cc_w_1_120_s_0_175 = '-6.46875e-13*ic_cap*ic_cap+-2.87500e-13*ic_cap+1.06000e-10'
+ mcm3m2f_cc_w_1_120_s_0_210 = '-4.93750e-13*ic_cap*ic_cap+-3.25000e-13*ic_cap+9.88000e-11'
+ mcm3m2f_cc_w_1_120_s_0_280 = '-3.15625e-13*ic_cap*ic_cap+-2.12500e-13*ic_cap+8.46000e-11'
+ mcm3m2f_cc_w_1_120_s_0_350 = '-2.15625e-13*ic_cap*ic_cap+-1.37500e-13*ic_cap+7.19000e-11'
+ mcm3m2f_cc_w_1_120_s_0_420 = '-1.03125e-13*ic_cap*ic_cap+-8.75000e-14*ic_cap+6.08000e-11'
+ mcm3m2f_cc_w_1_120_s_0_560 = '2.50000e-14*ic_cap*ic_cap+4.53000e-11'
+ mcm3m2f_cc_w_1_120_s_0_840 = '1.12500e-13*ic_cap*ic_cap+5.00000e-14*ic_cap+2.81000e-11'
+ mcm3m2f_cc_w_1_120_s_1_540 = '1.28125e-13*ic_cap*ic_cap+8.75000e-14*ic_cap+1.07000e-11'
+ mcm3m2f_cc_w_1_120_s_3_500 = '4.15625e-14*ic_cap*ic_cap+3.37500e-14*ic_cap+1.09000e-12'
+ mcm3m2f_cf_w_0_140_s_0_140 = '-3.65625e-14*ic_cap*ic_cap+-1.87500e-14*ic_cap+6.58000e-12'
+ mcm3m2f_cf_w_0_140_s_0_175 = '-5.78125e-14*ic_cap*ic_cap+-3.12500e-14*ic_cap+8.13000e-12'
+ mcm3m2f_cf_w_0_140_s_0_210 = '-7.65625e-14*ic_cap*ic_cap+-4.12500e-14*ic_cap+9.67000e-12'
+ mcm3m2f_cf_w_0_140_s_0_280 = '-1.15625e-13*ic_cap*ic_cap+-6.25000e-14*ic_cap+1.26000e-11'
+ mcm3m2f_cf_w_0_140_s_0_350 = '-1.50000e-13*ic_cap*ic_cap+-7.50000e-14*ic_cap+1.54000e-11'
+ mcm3m2f_cf_w_0_140_s_0_420 = '-1.84375e-13*ic_cap*ic_cap+-1.12500e-13*ic_cap+1.82000e-11'
+ mcm3m2f_cf_w_0_140_s_0_560 = '-2.40625e-13*ic_cap*ic_cap+-1.37500e-13*ic_cap+2.31000e-11'
+ mcm3m2f_cf_w_0_140_s_0_840 = '-3.25000e-13*ic_cap*ic_cap+-1.75000e-13*ic_cap+3.11000e-11'
+ mcm3m2f_cf_w_0_140_s_1_540 = '-3.84375e-13*ic_cap*ic_cap+-2.37500e-13*ic_cap+4.26000e-11'
+ mcm3m2f_cf_w_0_140_s_3_500 = '-3.43750e-13*ic_cap*ic_cap+-2.25000e-13*ic_cap+5.01000e-11'
+ mcm3m2f_cf_w_1_120_s_0_140 = '-3.56250e-14*ic_cap*ic_cap+-2.00000e-14*ic_cap+6.61000e-12'
+ mcm3m2f_cf_w_1_120_s_0_175 = '-5.68750e-14*ic_cap*ic_cap+-3.25000e-14*ic_cap+8.17000e-12'
+ mcm3m2f_cf_w_1_120_s_0_210 = '-7.71875e-14*ic_cap*ic_cap+-4.12500e-14*ic_cap+9.69000e-12'
+ mcm3m2f_cf_w_1_120_s_0_280 = '-1.15625e-13*ic_cap*ic_cap+-6.25000e-14*ic_cap+1.27000e-11'
+ mcm3m2f_cf_w_1_120_s_0_350 = '-1.46875e-13*ic_cap*ic_cap+-8.75000e-14*ic_cap+1.55000e-11'
+ mcm3m2f_cf_w_1_120_s_0_420 = '-1.78125e-13*ic_cap*ic_cap+-1.12500e-13*ic_cap+1.82000e-11'
+ mcm3m2f_cf_w_1_120_s_0_560 = '-2.34375e-13*ic_cap*ic_cap+-1.37500e-13*ic_cap+2.32000e-11'
+ mcm3m2f_cf_w_1_120_s_0_840 = '-3.15625e-13*ic_cap*ic_cap+-1.87500e-13*ic_cap+3.14000e-11'
+ mcm3m2f_cf_w_1_120_s_1_540 = '-3.78125e-13*ic_cap*ic_cap+-2.12500e-13*ic_cap+4.37000e-11'
+ mcm3m2f_cf_w_1_120_s_3_500 = '-3.18750e-13*ic_cap*ic_cap+-2.00000e-13*ic_cap+5.26000e-11'
+ mcm3m2l1_ca_w_0_140_s_0_140 = '-1.69063e-06*ic_cap*ic_cap+-9.62500e-07*ic_cap+1.19000e-04'
+ mcm3m2l1_ca_w_0_140_s_0_175 = '-1.69063e-06*ic_cap*ic_cap+-9.62500e-07*ic_cap+1.19000e-04'
+ mcm3m2l1_ca_w_0_140_s_0_210 = '-1.69063e-06*ic_cap*ic_cap+-9.62500e-07*ic_cap+1.19000e-04'
+ mcm3m2l1_ca_w_0_140_s_0_280 = '-1.69063e-06*ic_cap*ic_cap+-9.62500e-07*ic_cap+1.19000e-04'
+ mcm3m2l1_ca_w_0_140_s_0_350 = '-1.69063e-06*ic_cap*ic_cap+-9.62500e-07*ic_cap+1.19000e-04'
+ mcm3m2l1_ca_w_0_140_s_0_420 = '-1.69063e-06*ic_cap*ic_cap+-9.62500e-07*ic_cap+1.19000e-04'
+ mcm3m2l1_ca_w_0_140_s_0_560 = '-1.69063e-06*ic_cap*ic_cap+-9.62500e-07*ic_cap+1.19000e-04'
+ mcm3m2l1_ca_w_0_140_s_0_840 = '-1.69063e-06*ic_cap*ic_cap+-9.62500e-07*ic_cap+1.19000e-04'
+ mcm3m2l1_ca_w_0_140_s_1_540 = '-1.69063e-06*ic_cap*ic_cap+-9.62500e-07*ic_cap+1.19000e-04'
+ mcm3m2l1_ca_w_0_140_s_3_500 = '-1.69063e-06*ic_cap*ic_cap+-9.62500e-07*ic_cap+1.19000e-04'
+ mcm3m2l1_ca_w_1_120_s_0_140 = '-1.69063e-06*ic_cap*ic_cap+-9.62500e-07*ic_cap+1.19000e-04'
+ mcm3m2l1_ca_w_1_120_s_0_175 = '-1.69063e-06*ic_cap*ic_cap+-9.62500e-07*ic_cap+1.19000e-04'
+ mcm3m2l1_ca_w_1_120_s_0_210 = '-1.69063e-06*ic_cap*ic_cap+-9.62500e-07*ic_cap+1.19000e-04'
+ mcm3m2l1_ca_w_1_120_s_0_280 = '-1.69063e-06*ic_cap*ic_cap+-9.62500e-07*ic_cap+1.19000e-04'
+ mcm3m2l1_ca_w_1_120_s_0_350 = '-1.69063e-06*ic_cap*ic_cap+-9.62500e-07*ic_cap+1.19000e-04'
+ mcm3m2l1_ca_w_1_120_s_0_420 = '-1.69063e-06*ic_cap*ic_cap+-9.62500e-07*ic_cap+1.19000e-04'
+ mcm3m2l1_ca_w_1_120_s_0_560 = '-1.69063e-06*ic_cap*ic_cap+-9.62500e-07*ic_cap+1.19000e-04'
+ mcm3m2l1_ca_w_1_120_s_0_840 = '-1.69063e-06*ic_cap*ic_cap+-9.62500e-07*ic_cap+1.19000e-04'
+ mcm3m2l1_ca_w_1_120_s_1_540 = '-1.69063e-06*ic_cap*ic_cap+-9.62500e-07*ic_cap+1.19000e-04'
+ mcm3m2l1_ca_w_1_120_s_3_500 = '-1.69063e-06*ic_cap*ic_cap+-9.62500e-07*ic_cap+1.19000e-04'
+ mcm3m2l1_cc_w_0_140_s_0_140 = '-7.46875e-13*ic_cap*ic_cap+-4.37500e-13*ic_cap+9.45000e-11'
+ mcm3m2l1_cc_w_0_140_s_0_175 = '-7.28125e-13*ic_cap*ic_cap+-3.87500e-13*ic_cap+9.21000e-11'
+ mcm3m2l1_cc_w_0_140_s_0_210 = '-6.00000e-13*ic_cap*ic_cap+-4.00000e-13*ic_cap+8.62000e-11'
+ mcm3m2l1_cc_w_0_140_s_0_280 = '-4.06250e-13*ic_cap*ic_cap+-3.00000e-13*ic_cap+7.32000e-11'
+ mcm3m2l1_cc_w_0_140_s_0_350 = '-2.62500e-13*ic_cap*ic_cap+-2.00000e-13*ic_cap+6.08000e-11'
+ mcm3m2l1_cc_w_0_140_s_0_420 = '-1.71875e-13*ic_cap*ic_cap+-1.87500e-13*ic_cap+5.06000e-11'
+ mcm3m2l1_cc_w_0_140_s_0_560 = '-1.25000e-14*ic_cap*ic_cap+3.58000e-11'
+ mcm3m2l1_cc_w_0_140_s_0_840 = '8.75000e-14*ic_cap*ic_cap+5.00000e-14*ic_cap+1.98000e-11'
+ mcm3m2l1_cc_w_0_140_s_1_540 = '9.53125e-14*ic_cap*ic_cap+6.87500e-14*ic_cap+5.20000e-12'
+ mcm3m2l1_cc_w_0_140_s_3_500 = '1.07813e-14*ic_cap*ic_cap+8.12500e-15*ic_cap+2.10000e-13'
+ mcm3m2l1_cc_w_1_120_s_0_140 = '-5.78125e-13*ic_cap*ic_cap+-3.37500e-13*ic_cap+1.02000e-10'
+ mcm3m2l1_cc_w_1_120_s_0_175 = '-5.43750e-13*ic_cap*ic_cap+-2.25000e-13*ic_cap+9.84000e-11'
+ mcm3m2l1_cc_w_1_120_s_0_210 = '-4.40625e-13*ic_cap*ic_cap+-2.62500e-13*ic_cap+9.19000e-11'
+ mcm3m2l1_cc_w_1_120_s_0_280 = '-2.56250e-13*ic_cap*ic_cap+-1.75000e-13*ic_cap+7.72000e-11'
+ mcm3m2l1_cc_w_1_120_s_0_350 = '-1.34375e-13*ic_cap*ic_cap+-8.75000e-14*ic_cap+6.42000e-11'
+ mcm3m2l1_cc_w_1_120_s_0_420 = '-3.75000e-14*ic_cap*ic_cap+-5.00000e-14*ic_cap+5.32000e-11'
+ mcm3m2l1_cc_w_1_120_s_0_560 = '6.25000e-14*ic_cap*ic_cap+5.00000e-14*ic_cap+3.79000e-11'
+ mcm3m2l1_cc_w_1_120_s_0_840 = '1.50000e-13*ic_cap*ic_cap+1.00000e-13*ic_cap+2.09000e-11'
+ mcm3m2l1_cc_w_1_120_s_1_540 = '1.21562e-13*ic_cap*ic_cap+9.12500e-14*ic_cap+5.55000e-12'
+ mcm3m2l1_cc_w_1_120_s_3_500 = '1.26562e-14*ic_cap*ic_cap+1.43750e-14*ic_cap+2.35000e-13'
+ mcm3m2l1_cf_w_0_140_s_0_140 = '-4.18750e-14*ic_cap*ic_cap+-2.50000e-14*ic_cap+7.89000e-12'
+ mcm3m2l1_cf_w_0_140_s_0_175 = '-6.78125e-14*ic_cap*ic_cap+-3.87500e-14*ic_cap+9.79000e-12'
+ mcm3m2l1_cf_w_0_140_s_0_210 = '-8.84375e-14*ic_cap*ic_cap+-5.37500e-14*ic_cap+1.16000e-11'
+ mcm3m2l1_cf_w_0_140_s_0_280 = '-1.37500e-13*ic_cap*ic_cap+-7.50000e-14*ic_cap+1.52000e-11'
+ mcm3m2l1_cf_w_0_140_s_0_350 = '-1.84375e-13*ic_cap*ic_cap+-1.12500e-13*ic_cap+1.87000e-11'
+ mcm3m2l1_cf_w_0_140_s_0_420 = '-2.28125e-13*ic_cap*ic_cap+-1.37500e-13*ic_cap+2.21000e-11'
+ mcm3m2l1_cf_w_0_140_s_0_560 = '-2.93750e-13*ic_cap*ic_cap+-1.75000e-13*ic_cap+2.78000e-11'
+ mcm3m2l1_cf_w_0_140_s_0_840 = '-3.87500e-13*ic_cap*ic_cap+-2.25000e-13*ic_cap+3.71000e-11'
+ mcm3m2l1_cf_w_0_140_s_1_540 = '-4.31250e-13*ic_cap*ic_cap+-2.75000e-13*ic_cap+4.89000e-11'
+ mcm3m2l1_cf_w_0_140_s_3_500 = '-3.59375e-13*ic_cap*ic_cap+-2.37500e-13*ic_cap+5.38000e-11'
+ mcm3m2l1_cf_w_1_120_s_0_140 = '-4.12500e-14*ic_cap*ic_cap+-2.50000e-14*ic_cap+7.93000e-12'
+ mcm3m2l1_cf_w_1_120_s_0_175 = '-6.71875e-14*ic_cap*ic_cap+-4.12500e-14*ic_cap+9.84000e-12'
+ mcm3m2l1_cf_w_1_120_s_0_210 = '-9.37500e-14*ic_cap*ic_cap+-5.00000e-14*ic_cap+1.17000e-11'
+ mcm3m2l1_cf_w_1_120_s_0_280 = '-1.40625e-13*ic_cap*ic_cap+-8.75000e-14*ic_cap+1.53000e-11'
+ mcm3m2l1_cf_w_1_120_s_0_350 = '-1.84375e-13*ic_cap*ic_cap+-1.12500e-13*ic_cap+1.88000e-11'
+ mcm3m2l1_cf_w_1_120_s_0_420 = '-2.21875e-13*ic_cap*ic_cap+-1.12500e-13*ic_cap+2.21000e-11'
+ mcm3m2l1_cf_w_1_120_s_0_560 = '-2.93750e-13*ic_cap*ic_cap+-1.75000e-13*ic_cap+2.81000e-11'
+ mcm3m2l1_cf_w_1_120_s_0_840 = '-3.87500e-13*ic_cap*ic_cap+-2.25000e-13*ic_cap+3.76000e-11'
+ mcm3m2l1_cf_w_1_120_s_1_540 = '-4.03125e-13*ic_cap*ic_cap+-2.62500e-13*ic_cap+4.96000e-11'
+ mcm3m2l1_cf_w_1_120_s_3_500 = '-3.18750e-13*ic_cap*ic_cap+-2.00000e-13*ic_cap+5.51000e-11'
+ mcm3m2m1_ca_w_0_140_s_0_140 = '-3.90625e-06*ic_cap*ic_cap+-1.87500e-06*ic_cap+2.10000e-04'
+ mcm3m2m1_ca_w_0_140_s_0_175 = '-3.90625e-06*ic_cap*ic_cap+-1.87500e-06*ic_cap+2.10000e-04'
+ mcm3m2m1_ca_w_0_140_s_0_210 = '-3.90625e-06*ic_cap*ic_cap+-1.87500e-06*ic_cap+2.10000e-04'
+ mcm3m2m1_ca_w_0_140_s_0_280 = '-3.90625e-06*ic_cap*ic_cap+-1.87500e-06*ic_cap+2.10000e-04'
+ mcm3m2m1_ca_w_0_140_s_0_350 = '-3.90625e-06*ic_cap*ic_cap+-1.87500e-06*ic_cap+2.10000e-04'
+ mcm3m2m1_ca_w_0_140_s_0_420 = '-3.90625e-06*ic_cap*ic_cap+-1.87500e-06*ic_cap+2.10000e-04'
+ mcm3m2m1_ca_w_0_140_s_0_560 = '-3.90625e-06*ic_cap*ic_cap+-1.87500e-06*ic_cap+2.10000e-04'
+ mcm3m2m1_ca_w_0_140_s_0_840 = '-3.90625e-06*ic_cap*ic_cap+-1.87500e-06*ic_cap+2.10000e-04'
+ mcm3m2m1_ca_w_0_140_s_1_540 = '-3.90625e-06*ic_cap*ic_cap+-1.87500e-06*ic_cap+2.10000e-04'
+ mcm3m2m1_ca_w_0_140_s_3_500 = '-3.90625e-06*ic_cap*ic_cap+-1.87500e-06*ic_cap+2.10000e-04'
+ mcm3m2m1_ca_w_1_120_s_0_140 = '-3.90625e-06*ic_cap*ic_cap+-1.87500e-06*ic_cap+2.10000e-04'
+ mcm3m2m1_ca_w_1_120_s_0_175 = '-3.90625e-06*ic_cap*ic_cap+-1.87500e-06*ic_cap+2.10000e-04'
+ mcm3m2m1_ca_w_1_120_s_0_210 = '-3.90625e-06*ic_cap*ic_cap+-1.87500e-06*ic_cap+2.10000e-04'
+ mcm3m2m1_ca_w_1_120_s_0_280 = '-3.90625e-06*ic_cap*ic_cap+-1.87500e-06*ic_cap+2.10000e-04'
+ mcm3m2m1_ca_w_1_120_s_0_350 = '-3.90625e-06*ic_cap*ic_cap+-1.87500e-06*ic_cap+2.10000e-04'
+ mcm3m2m1_ca_w_1_120_s_0_420 = '-3.90625e-06*ic_cap*ic_cap+-1.87500e-06*ic_cap+2.10000e-04'
+ mcm3m2m1_ca_w_1_120_s_0_560 = '-3.90625e-06*ic_cap*ic_cap+-1.87500e-06*ic_cap+2.10000e-04'
+ mcm3m2m1_ca_w_1_120_s_0_840 = '-3.90625e-06*ic_cap*ic_cap+-1.87500e-06*ic_cap+2.10000e-04'
+ mcm3m2m1_ca_w_1_120_s_1_540 = '-3.90625e-06*ic_cap*ic_cap+-1.87500e-06*ic_cap+2.10000e-04'
+ mcm3m2m1_ca_w_1_120_s_3_500 = '-3.90625e-06*ic_cap*ic_cap+-1.87500e-06*ic_cap+2.10000e-04'
+ mcm3m2m1_cc_w_0_140_s_0_140 = '-6.18750e-13*ic_cap*ic_cap+-3.75000e-13*ic_cap+8.61000e-11'
+ mcm3m2m1_cc_w_0_140_s_0_175 = '-5.37500e-13*ic_cap*ic_cap+-3.00000e-13*ic_cap+8.31000e-11'
+ mcm3m2m1_cc_w_0_140_s_0_210 = '-4.09375e-13*ic_cap*ic_cap+-3.12500e-13*ic_cap+7.67000e-11'
+ mcm3m2m1_cc_w_0_140_s_0_280 = '-2.12500e-13*ic_cap*ic_cap+-1.75000e-13*ic_cap+6.27000e-11'
+ mcm3m2m1_cc_w_0_140_s_0_350 = '-9.06250e-14*ic_cap*ic_cap+-1.37500e-13*ic_cap+5.02000e-11'
+ mcm3m2m1_cc_w_0_140_s_0_420 = '2.18750e-14*ic_cap*ic_cap+-1.25000e-14*ic_cap+3.93000e-11'
+ mcm3m2m1_cc_w_0_140_s_0_560 = '1.34375e-13*ic_cap*ic_cap+3.75000e-14*ic_cap+2.50000e-11'
+ mcm3m2m1_cc_w_0_140_s_0_840 = '1.62500e-13*ic_cap*ic_cap+1.00000e-13*ic_cap+1.07000e-11'
+ mcm3m2m1_cc_w_0_140_s_1_540 = '6.65625e-14*ic_cap*ic_cap+4.37500e-14*ic_cap+1.40000e-12'
+ mcm3m2m1_cc_w_0_140_s_3_500 = '2.34375e-15*ic_cap*ic_cap+-1.87500e-15*ic_cap+3.00000e-14'
+ mcm3m2m1_cc_w_1_120_s_0_140 = '-4.59375e-13*ic_cap*ic_cap+-3.12500e-13*ic_cap+8.88000e-11'
+ mcm3m2m1_cc_w_1_120_s_0_175 = '-4.37500e-13*ic_cap*ic_cap+-2.50000e-13*ic_cap+8.57000e-11'
+ mcm3m2m1_cc_w_1_120_s_0_210 = '-3.09375e-13*ic_cap*ic_cap+-1.37500e-13*ic_cap+7.85000e-11'
+ mcm3m2m1_cc_w_1_120_s_0_280 = '-1.21875e-13*ic_cap*ic_cap+-1.37500e-13*ic_cap+6.38000e-11'
+ mcm3m2m1_cc_w_1_120_s_0_350 = '-2.50000e-14*ic_cap*ic_cap+5.11000e-11'
+ mcm3m2m1_cc_w_1_120_s_0_420 = '8.12500e-14*ic_cap*ic_cap+2.50000e-14*ic_cap+4.03000e-11'
+ mcm3m2m1_cc_w_1_120_s_0_560 = '1.78125e-13*ic_cap*ic_cap+8.75000e-14*ic_cap+2.57000e-11'
+ mcm3m2m1_cc_w_1_120_s_0_840 = '1.90625e-13*ic_cap*ic_cap+1.12500e-13*ic_cap+1.09000e-11'
+ mcm3m2m1_cc_w_1_120_s_1_540 = '7.50000e-14*ic_cap*ic_cap+6.25000e-14*ic_cap+1.40000e-12'
+ mcm3m2m1_cc_w_1_120_s_3_500 = '1.56250e-15*ic_cap*ic_cap+6.25000e-15*ic_cap+5.00000e-14'
+ mcm3m2m1_cf_w_0_140_s_0_140 = '-1.34375e-13*ic_cap*ic_cap+-6.25000e-14*ic_cap+1.36000e-11'
+ mcm3m2m1_cf_w_0_140_s_0_175 = '-1.93750e-13*ic_cap*ic_cap+-1.00000e-13*ic_cap+1.70000e-11'
+ mcm3m2m1_cf_w_0_140_s_0_210 = '-2.59375e-13*ic_cap*ic_cap+-1.37500e-13*ic_cap+2.04000e-11'
+ mcm3m2m1_cf_w_0_140_s_0_280 = '-3.71875e-13*ic_cap*ic_cap+-1.87500e-13*ic_cap+2.67000e-11'
+ mcm3m2m1_cf_w_0_140_s_0_350 = '-4.56250e-13*ic_cap*ic_cap+-2.25000e-13*ic_cap+3.24000e-11'
+ mcm3m2m1_cf_w_0_140_s_0_420 = '-5.50000e-13*ic_cap*ic_cap+-3.00000e-13*ic_cap+3.78000e-11'
+ mcm3m2m1_cf_w_0_140_s_0_560 = '-6.59375e-13*ic_cap*ic_cap+-3.62500e-13*ic_cap+4.64000e-11'
+ mcm3m2m1_cf_w_0_140_s_0_840 = '-7.68750e-13*ic_cap*ic_cap+-4.25000e-13*ic_cap+5.79000e-11'
+ mcm3m2m1_cf_w_0_140_s_1_540 = '-7.21875e-13*ic_cap*ic_cap+-4.12500e-13*ic_cap+6.72000e-11'
+ mcm3m2m1_cf_w_0_140_s_3_500 = '-6.59375e-13*ic_cap*ic_cap+-3.62500e-13*ic_cap+6.92000e-11'
+ mcm3m2m1_cf_w_1_120_s_0_140 = '-1.34375e-13*ic_cap*ic_cap+-6.25000e-14*ic_cap+1.36000e-11'
+ mcm3m2m1_cf_w_1_120_s_0_175 = '-2.00000e-13*ic_cap*ic_cap+-1.00000e-13*ic_cap+1.71000e-11'
+ mcm3m2m1_cf_w_1_120_s_0_210 = '-2.56250e-13*ic_cap*ic_cap+-1.25000e-13*ic_cap+2.04000e-11'
+ mcm3m2m1_cf_w_1_120_s_0_280 = '-3.65625e-13*ic_cap*ic_cap+-1.87500e-13*ic_cap+2.67000e-11'
+ mcm3m2m1_cf_w_1_120_s_0_350 = '-4.68750e-13*ic_cap*ic_cap+-2.25000e-13*ic_cap+3.26000e-11'
+ mcm3m2m1_cf_w_1_120_s_0_420 = '-5.37500e-13*ic_cap*ic_cap+-2.75000e-13*ic_cap+3.78000e-11'
+ mcm3m2m1_cf_w_1_120_s_0_560 = '-6.62500e-13*ic_cap*ic_cap+-3.50000e-13*ic_cap+4.67000e-11'
+ mcm3m2m1_cf_w_1_120_s_0_840 = '-7.62500e-13*ic_cap*ic_cap+-4.25000e-13*ic_cap+5.84000e-11'
+ mcm3m2m1_cf_w_1_120_s_1_540 = '-6.96875e-13*ic_cap*ic_cap+-3.87500e-13*ic_cap+6.78000e-11'
+ mcm3m2m1_cf_w_1_120_s_3_500 = '-6.40625e-13*ic_cap*ic_cap+-3.37500e-13*ic_cap+6.98000e-11'
+ mcm3m2p1_ca_w_0_140_s_0_140 = '-1.57188e-06*ic_cap*ic_cap+-8.62500e-07*ic_cap+1.07000e-04'
+ mcm3m2p1_ca_w_0_140_s_0_175 = '-1.57188e-06*ic_cap*ic_cap+-8.62500e-07*ic_cap+1.07000e-04'
+ mcm3m2p1_ca_w_0_140_s_0_210 = '-1.57188e-06*ic_cap*ic_cap+-8.62500e-07*ic_cap+1.07000e-04'
+ mcm3m2p1_ca_w_0_140_s_0_280 = '-1.57188e-06*ic_cap*ic_cap+-8.62500e-07*ic_cap+1.07000e-04'
+ mcm3m2p1_ca_w_0_140_s_0_350 = '-1.57188e-06*ic_cap*ic_cap+-8.62500e-07*ic_cap+1.07000e-04'
+ mcm3m2p1_ca_w_0_140_s_0_420 = '-1.57188e-06*ic_cap*ic_cap+-8.62500e-07*ic_cap+1.07000e-04'
+ mcm3m2p1_ca_w_0_140_s_0_560 = '-1.57188e-06*ic_cap*ic_cap+-8.62500e-07*ic_cap+1.07000e-04'
+ mcm3m2p1_ca_w_0_140_s_0_840 = '-1.57188e-06*ic_cap*ic_cap+-8.62500e-07*ic_cap+1.07000e-04'
+ mcm3m2p1_ca_w_0_140_s_1_540 = '-1.57188e-06*ic_cap*ic_cap+-8.62500e-07*ic_cap+1.07000e-04'
+ mcm3m2p1_ca_w_0_140_s_3_500 = '-1.57188e-06*ic_cap*ic_cap+-8.62500e-07*ic_cap+1.07000e-04'
+ mcm3m2p1_ca_w_1_120_s_0_140 = '-1.57188e-06*ic_cap*ic_cap+-8.62500e-07*ic_cap+1.07000e-04'
+ mcm3m2p1_ca_w_1_120_s_0_175 = '-1.57188e-06*ic_cap*ic_cap+-8.62500e-07*ic_cap+1.07000e-04'
+ mcm3m2p1_ca_w_1_120_s_0_210 = '-1.57188e-06*ic_cap*ic_cap+-8.62500e-07*ic_cap+1.07000e-04'
+ mcm3m2p1_ca_w_1_120_s_0_280 = '-1.57188e-06*ic_cap*ic_cap+-8.62500e-07*ic_cap+1.07000e-04'
+ mcm3m2p1_ca_w_1_120_s_0_350 = '-1.57188e-06*ic_cap*ic_cap+-8.62500e-07*ic_cap+1.07000e-04'
+ mcm3m2p1_ca_w_1_120_s_0_420 = '-1.57188e-06*ic_cap*ic_cap+-8.62500e-07*ic_cap+1.07000e-04'
+ mcm3m2p1_ca_w_1_120_s_0_560 = '-1.57188e-06*ic_cap*ic_cap+-8.62500e-07*ic_cap+1.07000e-04'
+ mcm3m2p1_ca_w_1_120_s_0_840 = '-1.57188e-06*ic_cap*ic_cap+-8.62500e-07*ic_cap+1.07000e-04'
+ mcm3m2p1_ca_w_1_120_s_1_540 = '-1.57188e-06*ic_cap*ic_cap+-8.62500e-07*ic_cap+1.07000e-04'
+ mcm3m2p1_ca_w_1_120_s_3_500 = '-1.57188e-06*ic_cap*ic_cap+-8.62500e-07*ic_cap+1.07000e-04'
+ mcm3m2p1_cc_w_0_140_s_0_140 = '-8.53125e-13*ic_cap*ic_cap+-3.62500e-13*ic_cap+9.70000e-11'
+ mcm3m2p1_cc_w_0_140_s_0_175 = '-7.40625e-13*ic_cap*ic_cap+-4.12500e-13*ic_cap+9.36000e-11'
+ mcm3m2p1_cc_w_0_140_s_0_210 = '-5.96875e-13*ic_cap*ic_cap+-4.12500e-13*ic_cap+8.75000e-11'
+ mcm3m2p1_cc_w_0_140_s_0_280 = '-4.28125e-13*ic_cap*ic_cap+-3.12500e-13*ic_cap+7.52000e-11'
+ mcm3m2p1_cc_w_0_140_s_0_350 = '-2.84375e-13*ic_cap*ic_cap+-2.37500e-13*ic_cap+6.30000e-11'
+ mcm3m2p1_cc_w_0_140_s_0_420 = '-1.68750e-13*ic_cap*ic_cap+-1.50000e-13*ic_cap+5.27000e-11'
+ mcm3m2p1_cc_w_0_140_s_0_560 = '-3.12500e-14*ic_cap*ic_cap+-5.00000e-14*ic_cap+3.85000e-11'
+ mcm3m2p1_cc_w_0_140_s_0_840 = '6.87500e-14*ic_cap*ic_cap+2.50000e-14*ic_cap+2.27000e-11'
+ mcm3m2p1_cc_w_0_140_s_1_540 = '1.01250e-13*ic_cap*ic_cap+6.00000e-14*ic_cap+7.25000e-12'
+ mcm3m2p1_cc_w_0_140_s_3_500 = '2.29687e-14*ic_cap*ic_cap+1.81250e-14*ic_cap+4.75000e-13'
+ mcm3m2p1_cc_w_1_120_s_0_140 = '-6.00000e-13*ic_cap*ic_cap+-2.75000e-13*ic_cap+1.06000e-10'
+ mcm3m2p1_cc_w_1_120_s_0_175 = '-6.06250e-13*ic_cap*ic_cap+-2.75000e-13*ic_cap+1.03000e-10'
+ mcm3m2p1_cc_w_1_120_s_0_210 = '-4.50000e-13*ic_cap*ic_cap+-3.00000e-13*ic_cap+9.58000e-11'
+ mcm3m2p1_cc_w_1_120_s_0_280 = '-2.93750e-13*ic_cap*ic_cap+-1.75000e-13*ic_cap+8.16000e-11'
+ mcm3m2p1_cc_w_1_120_s_0_350 = '-1.62500e-13*ic_cap*ic_cap+-1.50000e-13*ic_cap+6.87000e-11'
+ mcm3m2p1_cc_w_1_120_s_0_420 = '-7.50000e-14*ic_cap*ic_cap+-7.50000e-14*ic_cap+5.77000e-11'
+ mcm3m2p1_cc_w_1_120_s_0_560 = '6.25000e-14*ic_cap*ic_cap+2.50000e-14*ic_cap+4.20000e-11'
+ mcm3m2p1_cc_w_1_120_s_0_840 = '1.43750e-13*ic_cap*ic_cap+1.00000e-13*ic_cap+2.49000e-11'
+ mcm3m2p1_cc_w_1_120_s_1_540 = '1.46250e-13*ic_cap*ic_cap+1.00000e-13*ic_cap+8.16000e-12'
+ mcm3m2p1_cc_w_1_120_s_3_500 = '2.95312e-14*ic_cap*ic_cap+2.31250e-14*ic_cap+5.15000e-13'
+ mcm3m2p1_cf_w_0_140_s_0_140 = '-4.09375e-14*ic_cap*ic_cap+-2.37500e-14*ic_cap+7.08000e-12'
+ mcm3m2p1_cf_w_0_140_s_0_175 = '-6.46875e-14*ic_cap*ic_cap+-3.37500e-14*ic_cap+8.76000e-12'
+ mcm3m2p1_cf_w_0_140_s_0_210 = '-8.43750e-14*ic_cap*ic_cap+-5.00000e-14*ic_cap+1.04000e-11'
+ mcm3m2p1_cf_w_0_140_s_0_280 = '-1.31250e-13*ic_cap*ic_cap+-7.50000e-14*ic_cap+1.36000e-11'
+ mcm3m2p1_cf_w_0_140_s_0_350 = '-1.68750e-13*ic_cap*ic_cap+-1.00000e-13*ic_cap+1.67000e-11'
+ mcm3m2p1_cf_w_0_140_s_0_420 = '-2.03125e-13*ic_cap*ic_cap+-1.12500e-13*ic_cap+1.96000e-11'
+ mcm3m2p1_cf_w_0_140_s_0_560 = '-2.65625e-13*ic_cap*ic_cap+-1.62500e-13*ic_cap+2.48000e-11'
+ mcm3m2p1_cf_w_0_140_s_0_840 = '-3.50000e-13*ic_cap*ic_cap+-2.25000e-13*ic_cap+3.33000e-11'
+ mcm3m2p1_cf_w_0_140_s_1_540 = '-4.12500e-13*ic_cap*ic_cap+-2.50000e-13*ic_cap+4.51000e-11'
+ mcm3m2p1_cf_w_0_140_s_3_500 = '-3.56250e-13*ic_cap*ic_cap+-2.25000e-13*ic_cap+5.16000e-11'
+ mcm3m2p1_cf_w_1_120_s_0_140 = '-4.03125e-14*ic_cap*ic_cap+-2.37500e-14*ic_cap+7.13000e-12'
+ mcm3m2p1_cf_w_1_120_s_0_175 = '-6.37500e-14*ic_cap*ic_cap+-3.75000e-14*ic_cap+8.82000e-12'
+ mcm3m2p1_cf_w_1_120_s_0_210 = '-8.78125e-14*ic_cap*ic_cap+-4.87500e-14*ic_cap+1.05000e-11'
+ mcm3m2p1_cf_w_1_120_s_0_280 = '-1.31250e-13*ic_cap*ic_cap+-7.50000e-14*ic_cap+1.37000e-11'
+ mcm3m2p1_cf_w_1_120_s_0_350 = '-1.68750e-13*ic_cap*ic_cap+-1.00000e-13*ic_cap+1.68000e-11'
+ mcm3m2p1_cf_w_1_120_s_0_420 = '-2.00000e-13*ic_cap*ic_cap+-1.25000e-13*ic_cap+1.97000e-11'
+ mcm3m2p1_cf_w_1_120_s_0_560 = '-2.68750e-13*ic_cap*ic_cap+-1.50000e-13*ic_cap+2.51000e-11'
+ mcm3m2p1_cf_w_1_120_s_0_840 = '-3.50000e-13*ic_cap*ic_cap+-2.00000e-13*ic_cap+3.37000e-11'
+ mcm3m2p1_cf_w_1_120_s_1_540 = '-4.03125e-13*ic_cap*ic_cap+-2.37500e-13*ic_cap+4.62000e-11'
+ mcm3m2p1_cf_w_1_120_s_3_500 = '-3.18750e-13*ic_cap*ic_cap+-2.00000e-13*ic_cap+5.35000e-11'
+ mcm3p1_ca_w_0_300_s_0_300 = '-1.71875e-07*ic_cap*ic_cap+-1.12500e-07*ic_cap+1.58000e-05'
+ mcm3p1_ca_w_0_300_s_0_360 = '-1.71875e-07*ic_cap*ic_cap+-1.12500e-07*ic_cap+1.58000e-05'
+ mcm3p1_ca_w_0_300_s_0_450 = '-1.71875e-07*ic_cap*ic_cap+-1.12500e-07*ic_cap+1.58000e-05'
+ mcm3p1_ca_w_0_300_s_0_600 = '-1.71875e-07*ic_cap*ic_cap+-1.12500e-07*ic_cap+1.58000e-05'
+ mcm3p1_ca_w_0_300_s_0_800 = '-1.71875e-07*ic_cap*ic_cap+-1.12500e-07*ic_cap+1.58000e-05'
+ mcm3p1_ca_w_0_300_s_1_000 = '-1.71875e-07*ic_cap*ic_cap+-1.12500e-07*ic_cap+1.58000e-05'
+ mcm3p1_ca_w_0_300_s_1_200 = '-1.71875e-07*ic_cap*ic_cap+-1.12500e-07*ic_cap+1.58000e-05'
+ mcm3p1_ca_w_0_300_s_2_100 = '-1.71875e-07*ic_cap*ic_cap+-1.12500e-07*ic_cap+1.58000e-05'
+ mcm3p1_ca_w_0_300_s_3_300 = '-1.71875e-07*ic_cap*ic_cap+-1.12500e-07*ic_cap+1.58000e-05'
+ mcm3p1_ca_w_0_300_s_9_000 = '-1.71875e-07*ic_cap*ic_cap+-1.12500e-07*ic_cap+1.58000e-05'
+ mcm3p1_ca_w_2_400_s_0_300 = '-1.71875e-07*ic_cap*ic_cap+-1.12500e-07*ic_cap+1.58000e-05'
+ mcm3p1_ca_w_2_400_s_0_360 = '-1.71875e-07*ic_cap*ic_cap+-1.12500e-07*ic_cap+1.58000e-05'
+ mcm3p1_ca_w_2_400_s_0_450 = '-1.71875e-07*ic_cap*ic_cap+-1.12500e-07*ic_cap+1.58000e-05'
+ mcm3p1_ca_w_2_400_s_0_600 = '-1.71875e-07*ic_cap*ic_cap+-1.12500e-07*ic_cap+1.58000e-05'
+ mcm3p1_ca_w_2_400_s_0_800 = '-1.71875e-07*ic_cap*ic_cap+-1.12500e-07*ic_cap+1.58000e-05'
+ mcm3p1_ca_w_2_400_s_1_000 = '-1.71875e-07*ic_cap*ic_cap+-1.12500e-07*ic_cap+1.58000e-05'
+ mcm3p1_ca_w_2_400_s_1_200 = '-1.71875e-07*ic_cap*ic_cap+-1.12500e-07*ic_cap+1.58000e-05'
+ mcm3p1_ca_w_2_400_s_2_100 = '-1.71875e-07*ic_cap*ic_cap+-1.12500e-07*ic_cap+1.58000e-05'
+ mcm3p1_ca_w_2_400_s_3_300 = '-1.71875e-07*ic_cap*ic_cap+-1.12500e-07*ic_cap+1.58000e-05'
+ mcm3p1_ca_w_2_400_s_9_000 = '-1.71875e-07*ic_cap*ic_cap+-1.12500e-07*ic_cap+1.58000e-05'
+ mcm3p1_cc_w_0_300_s_0_300 = '-8.06250e-13*ic_cap*ic_cap+-4.50000e-13*ic_cap+1.06000e-10'
+ mcm3p1_cc_w_0_300_s_0_360 = '-6.75000e-13*ic_cap*ic_cap+-4.00000e-13*ic_cap+9.84000e-11'
+ mcm3p1_cc_w_0_300_s_0_450 = '-5.68750e-13*ic_cap*ic_cap+-3.50000e-13*ic_cap+8.89000e-11'
+ mcm3p1_cc_w_0_300_s_0_600 = '-4.28125e-13*ic_cap*ic_cap+-2.62500e-13*ic_cap+7.62000e-11'
+ mcm3p1_cc_w_0_300_s_0_800 = '-3.00000e-13*ic_cap*ic_cap+-2.25000e-13*ic_cap+6.40000e-11'
+ mcm3p1_cc_w_0_300_s_1_000 = '-2.12500e-13*ic_cap*ic_cap+-1.50000e-13*ic_cap+5.48000e-11'
+ mcm3p1_cc_w_0_300_s_1_200 = '-1.53125e-13*ic_cap*ic_cap+-1.12500e-13*ic_cap+4.79000e-11'
+ mcm3p1_cc_w_0_300_s_2_100 = '-3.75000e-14*ic_cap*ic_cap+-2.50000e-14*ic_cap+3.07000e-11'
+ mcm3p1_cc_w_0_300_s_3_300 = '1.25000e-14*ic_cap*ic_cap+2.06000e-11'
+ mcm3p1_cc_w_0_300_s_9_000 = '2.68750e-14*ic_cap*ic_cap+2.25000e-14*ic_cap+5.69000e-12'
+ mcm3p1_cc_w_2_400_s_0_300 = '-6.87500e-13*ic_cap*ic_cap+-5.00000e-13*ic_cap+1.29000e-10'
+ mcm3p1_cc_w_2_400_s_0_360 = '-6.25000e-13*ic_cap*ic_cap+-2.50000e-13*ic_cap+1.21000e-10'
+ mcm3p1_cc_w_2_400_s_0_450 = '-4.37500e-13*ic_cap*ic_cap+-2.50000e-13*ic_cap+1.09000e-10'
+ mcm3p1_cc_w_2_400_s_0_600 = '-3.59375e-13*ic_cap*ic_cap+-2.12500e-13*ic_cap+9.49000e-11'
+ mcm3p1_cc_w_2_400_s_0_800 = '-2.21875e-13*ic_cap*ic_cap+-1.37500e-13*ic_cap+8.02000e-11'
+ mcm3p1_cc_w_2_400_s_1_000 = '-1.43750e-13*ic_cap*ic_cap+-1.00000e-13*ic_cap+6.94000e-11'
+ mcm3p1_cc_w_2_400_s_1_200 = '-9.06250e-14*ic_cap*ic_cap+-6.25000e-14*ic_cap+6.13000e-11'
+ mcm3p1_cc_w_2_400_s_2_100 = '6.25000e-15*ic_cap*ic_cap+4.10000e-11'
+ mcm3p1_cc_w_2_400_s_3_300 = '4.06250e-14*ic_cap*ic_cap+1.25000e-14*ic_cap+2.83000e-11'
+ mcm3p1_cc_w_2_400_s_9_000 = '4.59375e-14*ic_cap*ic_cap+2.37500e-14*ic_cap+9.05000e-12'
+ mcm3p1_cf_w_0_300_s_0_300 = '-9.68750e-15*ic_cap*ic_cap+-6.25000e-15*ic_cap+2.34000e-12'
+ mcm3p1_cf_w_0_300_s_0_360 = '-1.50000e-14*ic_cap*ic_cap+-1.00000e-14*ic_cap+2.80000e-12'
+ mcm3p1_cf_w_0_300_s_0_450 = '-2.21875e-14*ic_cap*ic_cap+-1.37500e-14*ic_cap+3.50000e-12'
+ mcm3p1_cf_w_0_300_s_0_600 = '-3.34375e-14*ic_cap*ic_cap+-2.12500e-14*ic_cap+4.63000e-12'
+ mcm3p1_cf_w_0_300_s_0_800 = '-4.87500e-14*ic_cap*ic_cap+-3.00000e-14*ic_cap+6.00000e-12'
+ mcm3p1_cf_w_0_300_s_1_000 = '-6.37500e-14*ic_cap*ic_cap+-4.00000e-14*ic_cap+7.39000e-12'
+ mcm3p1_cf_w_0_300_s_1_200 = '-7.59375e-14*ic_cap*ic_cap+-4.87500e-14*ic_cap+8.70000e-12'
+ mcm3p1_cf_w_0_300_s_2_100 = '-1.28125e-13*ic_cap*ic_cap+-8.75000e-14*ic_cap+1.44000e-11'
+ mcm3p1_cf_w_0_300_s_3_300 = '-1.65625e-13*ic_cap*ic_cap+-1.12500e-13*ic_cap+1.96000e-11'
+ mcm3p1_cf_w_0_300_s_9_000 = '-2.03125e-13*ic_cap*ic_cap+-1.37500e-13*ic_cap+3.15000e-11'
+ mcm3p1_cf_w_2_400_s_0_300 = '-1.12500e-14*ic_cap*ic_cap+-7.50000e-15*ic_cap+2.42000e-12'
+ mcm3p1_cf_w_2_400_s_0_360 = '-1.56250e-14*ic_cap*ic_cap+-1.00000e-14*ic_cap+2.87000e-12'
+ mcm3p1_cf_w_2_400_s_0_450 = '-2.31250e-14*ic_cap*ic_cap+-1.50000e-14*ic_cap+3.55000e-12'
+ mcm3p1_cf_w_2_400_s_0_600 = '-3.53125e-14*ic_cap*ic_cap+-2.12500e-14*ic_cap+4.66000e-12'
+ mcm3p1_cf_w_2_400_s_0_800 = '-5.03125e-14*ic_cap*ic_cap+-3.12500e-14*ic_cap+6.10000e-12'
+ mcm3p1_cf_w_2_400_s_1_000 = '-6.43750e-14*ic_cap*ic_cap+-4.00000e-14*ic_cap+7.49000e-12'
+ mcm3p1_cf_w_2_400_s_1_200 = '-7.78125e-14*ic_cap*ic_cap+-4.87500e-14*ic_cap+8.85000e-12'
+ mcm3p1_cf_w_2_400_s_2_100 = '-1.25000e-13*ic_cap*ic_cap+-7.50000e-14*ic_cap+1.43000e-11'
+ mcm3p1_cf_w_2_400_s_3_300 = '-1.71875e-13*ic_cap*ic_cap+-1.12500e-13*ic_cap+2.03000e-11'
+ mcm3p1_cf_w_2_400_s_9_000 = '-2.09375e-13*ic_cap*ic_cap+-1.37500e-13*ic_cap+3.46000e-11'
+ mcm3p1f_ca_w_0_150_s_0_210 = '-1.59062e-06*ic_cap*ic_cap+-8.62500e-07*ic_cap+1.22000e-04'
+ mcm3p1f_ca_w_0_150_s_0_263 = '-1.59062e-06*ic_cap*ic_cap+-8.62500e-07*ic_cap+1.22000e-04'
+ mcm3p1f_ca_w_0_150_s_0_315 = '-1.59062e-06*ic_cap*ic_cap+-8.62500e-07*ic_cap+1.22000e-04'
+ mcm3p1f_ca_w_0_150_s_0_420 = '-1.59062e-06*ic_cap*ic_cap+-8.62500e-07*ic_cap+1.22000e-04'
+ mcm3p1f_ca_w_0_150_s_0_525 = '-1.59062e-06*ic_cap*ic_cap+-8.62500e-07*ic_cap+1.22000e-04'
+ mcm3p1f_ca_w_0_150_s_0_630 = '-1.59062e-06*ic_cap*ic_cap+-8.62500e-07*ic_cap+1.22000e-04'
+ mcm3p1f_ca_w_0_150_s_0_840 = '-1.59062e-06*ic_cap*ic_cap+-8.62500e-07*ic_cap+1.22000e-04'
+ mcm3p1f_ca_w_0_150_s_1_260 = '-1.59062e-06*ic_cap*ic_cap+-8.62500e-07*ic_cap+1.22000e-04'
+ mcm3p1f_ca_w_0_150_s_2_310 = '-1.59062e-06*ic_cap*ic_cap+-8.62500e-07*ic_cap+1.22000e-04'
+ mcm3p1f_ca_w_0_150_s_5_250 = '-1.59062e-06*ic_cap*ic_cap+-8.62500e-07*ic_cap+1.22000e-04'
+ mcm3p1f_ca_w_1_200_s_0_210 = '-1.59062e-06*ic_cap*ic_cap+-8.62500e-07*ic_cap+1.22000e-04'
+ mcm3p1f_ca_w_1_200_s_0_263 = '-1.59062e-06*ic_cap*ic_cap+-8.62500e-07*ic_cap+1.22000e-04'
+ mcm3p1f_ca_w_1_200_s_0_315 = '-1.59062e-06*ic_cap*ic_cap+-8.62500e-07*ic_cap+1.22000e-04'
+ mcm3p1f_ca_w_1_200_s_0_420 = '-1.59062e-06*ic_cap*ic_cap+-8.62500e-07*ic_cap+1.22000e-04'
+ mcm3p1f_ca_w_1_200_s_0_525 = '-1.59062e-06*ic_cap*ic_cap+-8.62500e-07*ic_cap+1.22000e-04'
+ mcm3p1f_ca_w_1_200_s_0_630 = '-1.59062e-06*ic_cap*ic_cap+-8.62500e-07*ic_cap+1.22000e-04'
+ mcm3p1f_ca_w_1_200_s_0_840 = '-1.59062e-06*ic_cap*ic_cap+-8.62500e-07*ic_cap+1.22000e-04'
+ mcm3p1f_ca_w_1_200_s_1_260 = '-1.59062e-06*ic_cap*ic_cap+-8.62500e-07*ic_cap+1.22000e-04'
+ mcm3p1f_ca_w_1_200_s_2_310 = '-1.59062e-06*ic_cap*ic_cap+-8.62500e-07*ic_cap+1.22000e-04'
+ mcm3p1f_ca_w_1_200_s_5_250 = '-1.59062e-06*ic_cap*ic_cap+-8.62500e-07*ic_cap+1.22000e-04'
+ mcm3p1f_cc_w_0_150_s_0_210 = '-5.40625e-13*ic_cap*ic_cap+-3.12500e-13*ic_cap+7.38000e-11'
+ mcm3p1f_cc_w_0_150_s_0_263 = '-3.46875e-13*ic_cap*ic_cap+-2.12500e-13*ic_cap+5.94000e-11'
+ mcm3p1f_cc_w_0_150_s_0_315 = '-2.34375e-13*ic_cap*ic_cap+-1.37500e-13*ic_cap+4.99000e-11'
+ mcm3p1f_cc_w_0_150_s_0_420 = '-1.06250e-13*ic_cap*ic_cap+-7.50000e-14*ic_cap+3.71000e-11'
+ mcm3p1f_cc_w_0_150_s_0_525 = '-4.37500e-14*ic_cap*ic_cap+-2.50000e-14*ic_cap+2.91000e-11'
+ mcm3p1f_cc_w_0_150_s_0_630 = '-6.25000e-15*ic_cap*ic_cap+2.34000e-11'
+ mcm3p1f_cc_w_0_150_s_0_840 = '3.43750e-14*ic_cap*ic_cap+1.25000e-14*ic_cap+1.58000e-11'
+ mcm3p1f_cc_w_0_150_s_1_260 = '4.46875e-14*ic_cap*ic_cap+3.37500e-14*ic_cap+7.92000e-12'
+ mcm3p1f_cc_w_0_150_s_2_310 = '3.06250e-14*ic_cap*ic_cap+2.00000e-14*ic_cap+1.95000e-12'
+ mcm3p1f_cc_w_0_150_s_5_250 = '4.53125e-15*ic_cap*ic_cap+1.87500e-15*ic_cap+1.05000e-13'
+ mcm3p1f_cc_w_1_200_s_0_210 = '-4.81250e-13*ic_cap*ic_cap+-2.75000e-13*ic_cap+8.57000e-11'
+ mcm3p1f_cc_w_1_200_s_0_263 = '-2.75000e-13*ic_cap*ic_cap+-1.50000e-13*ic_cap+6.98000e-11'
+ mcm3p1f_cc_w_1_200_s_0_315 = '-1.68750e-13*ic_cap*ic_cap+-1.00000e-13*ic_cap+5.93000e-11'
+ mcm3p1f_cc_w_1_200_s_0_420 = '-4.06250e-14*ic_cap*ic_cap+-1.25000e-14*ic_cap+4.51000e-11'
+ mcm3p1f_cc_w_1_200_s_0_525 = '2.18750e-14*ic_cap*ic_cap+1.25000e-14*ic_cap+3.60000e-11'
+ mcm3p1f_cc_w_1_200_s_0_630 = '4.37500e-14*ic_cap*ic_cap+2.50000e-14*ic_cap+2.96000e-11'
+ mcm3p1f_cc_w_1_200_s_0_840 = '8.12500e-14*ic_cap*ic_cap+5.00000e-14*ic_cap+2.08000e-11'
+ mcm3p1f_cc_w_1_200_s_1_260 = '9.37500e-14*ic_cap*ic_cap+7.50000e-14*ic_cap+1.13000e-11'
+ mcm3p1f_cc_w_1_200_s_2_310 = '5.65625e-14*ic_cap*ic_cap+3.87500e-14*ic_cap+3.11000e-12'
+ mcm3p1f_cc_w_1_200_s_5_250 = '8.43750e-15*ic_cap*ic_cap+2.50000e-15*ic_cap+1.50000e-13'
+ mcm3p1f_cf_w_0_150_s_0_210 = '-9.68750e-14*ic_cap*ic_cap+-6.25000e-14*ic_cap+1.19000e-11'
+ mcm3p1f_cf_w_0_150_s_0_263 = '-1.31250e-13*ic_cap*ic_cap+-7.50000e-14*ic_cap+1.45000e-11'
+ mcm3p1f_cf_w_0_150_s_0_315 = '-1.59375e-13*ic_cap*ic_cap+-8.75000e-14*ic_cap+1.69000e-11'
+ mcm3p1f_cf_w_0_150_s_0_420 = '-2.03125e-13*ic_cap*ic_cap+-1.12500e-13*ic_cap+2.14000e-11'
+ mcm3p1f_cf_w_0_150_s_0_525 = '-2.46875e-13*ic_cap*ic_cap+-1.37500e-13*ic_cap+2.53000e-11'
+ mcm3p1f_cf_w_0_150_s_0_630 = '-2.71875e-13*ic_cap*ic_cap+-1.62500e-13*ic_cap+2.85000e-11'
+ mcm3p1f_cf_w_0_150_s_0_840 = '-3.06250e-13*ic_cap*ic_cap+-1.75000e-13*ic_cap+3.37000e-11'
+ mcm3p1f_cf_w_0_150_s_1_260 = '-3.25000e-13*ic_cap*ic_cap+-2.00000e-13*ic_cap+4.01000e-11'
+ mcm3p1f_cf_w_0_150_s_2_310 = '-3.15625e-13*ic_cap*ic_cap+-1.87500e-13*ic_cap+4.55000e-11'
+ mcm3p1f_cf_w_0_150_s_5_250 = '-2.87500e-13*ic_cap*ic_cap+-1.75000e-13*ic_cap+4.73000e-11'
+ mcm3p1f_cf_w_1_200_s_0_210 = '-1.03125e-13*ic_cap*ic_cap+-6.25000e-14*ic_cap+1.19000e-11'
+ mcm3p1f_cf_w_1_200_s_0_263 = '-1.31250e-13*ic_cap*ic_cap+-7.50000e-14*ic_cap+1.45000e-11'
+ mcm3p1f_cf_w_1_200_s_0_315 = '-1.53125e-13*ic_cap*ic_cap+-8.75000e-14*ic_cap+1.69000e-11'
+ mcm3p1f_cf_w_1_200_s_0_420 = '-2.03125e-13*ic_cap*ic_cap+-1.12500e-13*ic_cap+2.14000e-11'
+ mcm3p1f_cf_w_1_200_s_0_525 = '-2.40625e-13*ic_cap*ic_cap+-1.37500e-13*ic_cap+2.54000e-11'
+ mcm3p1f_cf_w_1_200_s_0_630 = '-2.65625e-13*ic_cap*ic_cap+-1.62500e-13*ic_cap+2.88000e-11'
+ mcm3p1f_cf_w_1_200_s_0_840 = '-3.03125e-13*ic_cap*ic_cap+-1.87500e-13*ic_cap+3.44000e-11'
+ mcm3p1f_cf_w_1_200_s_1_260 = '-3.25000e-13*ic_cap*ic_cap+-2.00000e-13*ic_cap+4.16000e-11'
+ mcm3p1f_cf_w_1_200_s_2_310 = '-3.09375e-13*ic_cap*ic_cap+-1.87500e-13*ic_cap+4.90000e-11'
+ mcm3p1f_cf_w_1_200_s_5_250 = '-2.59375e-13*ic_cap*ic_cap+-1.62500e-13*ic_cap+5.19000e-11'
+ mcm4d_ca_w_0_300_s_0_300 = '-7.71875e-08*ic_cap*ic_cap+-4.87500e-08*ic_cap+9.41000e-06'
+ mcm4d_ca_w_0_300_s_0_360 = '-7.71875e-08*ic_cap*ic_cap+-4.87500e-08*ic_cap+9.41000e-06'
+ mcm4d_ca_w_0_300_s_0_450 = '-7.71875e-08*ic_cap*ic_cap+-4.87500e-08*ic_cap+9.41000e-06'
+ mcm4d_ca_w_0_300_s_0_600 = '-7.71875e-08*ic_cap*ic_cap+-4.87500e-08*ic_cap+9.41000e-06'
+ mcm4d_ca_w_0_300_s_0_800 = '-7.71875e-08*ic_cap*ic_cap+-4.87500e-08*ic_cap+9.41000e-06'
+ mcm4d_ca_w_0_300_s_1_000 = '-7.71875e-08*ic_cap*ic_cap+-4.87500e-08*ic_cap+9.41000e-06'
+ mcm4d_ca_w_0_300_s_1_200 = '-7.71875e-08*ic_cap*ic_cap+-4.87500e-08*ic_cap+9.41000e-06'
+ mcm4d_ca_w_0_300_s_2_100 = '-7.71875e-08*ic_cap*ic_cap+-4.87500e-08*ic_cap+9.41000e-06'
+ mcm4d_ca_w_0_300_s_3_300 = '-7.71875e-08*ic_cap*ic_cap+-4.87500e-08*ic_cap+9.41000e-06'
+ mcm4d_ca_w_0_300_s_9_000 = '-7.71875e-08*ic_cap*ic_cap+-4.87500e-08*ic_cap+9.41000e-06'
+ mcm4d_ca_w_2_400_s_0_300 = '-7.71875e-08*ic_cap*ic_cap+-4.87500e-08*ic_cap+9.41000e-06'
+ mcm4d_ca_w_2_400_s_0_360 = '-7.71875e-08*ic_cap*ic_cap+-4.87500e-08*ic_cap+9.41000e-06'
+ mcm4d_ca_w_2_400_s_0_450 = '-7.71875e-08*ic_cap*ic_cap+-4.87500e-08*ic_cap+9.41000e-06'
+ mcm4d_ca_w_2_400_s_0_600 = '-7.71875e-08*ic_cap*ic_cap+-4.87500e-08*ic_cap+9.41000e-06'
+ mcm4d_ca_w_2_400_s_0_800 = '-7.71875e-08*ic_cap*ic_cap+-4.87500e-08*ic_cap+9.41000e-06'
+ mcm4d_ca_w_2_400_s_1_000 = '-7.71875e-08*ic_cap*ic_cap+-4.87500e-08*ic_cap+9.41000e-06'
+ mcm4d_ca_w_2_400_s_1_200 = '-7.71875e-08*ic_cap*ic_cap+-4.87500e-08*ic_cap+9.41000e-06'
+ mcm4d_ca_w_2_400_s_2_100 = '-7.71875e-08*ic_cap*ic_cap+-4.87500e-08*ic_cap+9.41000e-06'
+ mcm4d_ca_w_2_400_s_3_300 = '-7.71875e-08*ic_cap*ic_cap+-4.87500e-08*ic_cap+9.41000e-06'
+ mcm4d_ca_w_2_400_s_9_000 = '-7.71875e-08*ic_cap*ic_cap+-4.87500e-08*ic_cap+9.41000e-06'
+ mcm4d_cc_w_0_300_s_0_300 = '-8.34375e-13*ic_cap*ic_cap+-4.87500e-13*ic_cap+1.08000e-10'
+ mcm4d_cc_w_0_300_s_0_360 = '-7.50000e-13*ic_cap*ic_cap+-4.50000e-13*ic_cap+1.01000e-10'
+ mcm4d_cc_w_0_300_s_0_450 = '-6.21875e-13*ic_cap*ic_cap+-3.62500e-13*ic_cap+9.14000e-11'
+ mcm4d_cc_w_0_300_s_0_600 = '-4.93750e-13*ic_cap*ic_cap+-3.00000e-13*ic_cap+7.93000e-11'
+ mcm4d_cc_w_0_300_s_0_800 = '-3.62500e-13*ic_cap*ic_cap+-2.25000e-13*ic_cap+6.75000e-11'
+ mcm4d_cc_w_0_300_s_1_000 = '-2.87500e-13*ic_cap*ic_cap+-1.75000e-13*ic_cap+5.87000e-11'
+ mcm4d_cc_w_0_300_s_1_200 = '-2.28125e-13*ic_cap*ic_cap+-1.37500e-13*ic_cap+5.20000e-11'
+ mcm4d_cc_w_0_300_s_2_100 = '-1.09375e-13*ic_cap*ic_cap+-8.75000e-14*ic_cap+3.54000e-11'
+ mcm4d_cc_w_0_300_s_3_300 = '-4.68750e-14*ic_cap*ic_cap+-3.75000e-14*ic_cap+2.53000e-11'
+ mcm4d_cc_w_0_300_s_9_000 = '1.65625e-14*ic_cap*ic_cap+1.12500e-14*ic_cap+8.44000e-12'
+ mcm4d_cc_w_2_400_s_0_300 = '-8.43750e-13*ic_cap*ic_cap+-3.75000e-13*ic_cap+1.36000e-10'
+ mcm4d_cc_w_2_400_s_0_360 = '-7.18750e-13*ic_cap*ic_cap+-3.75000e-13*ic_cap+1.27000e-10'
+ mcm4d_cc_w_2_400_s_0_450 = '-6.56250e-13*ic_cap*ic_cap+-3.75000e-13*ic_cap+1.17000e-10'
+ mcm4d_cc_w_2_400_s_0_600 = '-4.25000e-13*ic_cap*ic_cap+-2.75000e-13*ic_cap+1.01000e-10'
+ mcm4d_cc_w_2_400_s_0_800 = '-3.25000e-13*ic_cap*ic_cap+-2.00000e-13*ic_cap+8.67000e-11'
+ mcm4d_cc_w_2_400_s_1_000 = '-2.43750e-13*ic_cap*ic_cap+-1.75000e-13*ic_cap+7.59000e-11'
+ mcm4d_cc_w_2_400_s_1_200 = '-1.90625e-13*ic_cap*ic_cap+-1.37500e-13*ic_cap+6.77000e-11'
+ mcm4d_cc_w_2_400_s_2_100 = '-7.50000e-14*ic_cap*ic_cap+-5.00000e-14*ic_cap+4.69000e-11'
+ mcm4d_cc_w_2_400_s_3_300 = '-1.56250e-14*ic_cap*ic_cap+-1.25000e-14*ic_cap+3.36000e-11'
+ mcm4d_cc_w_2_400_s_9_000 = '3.12500e-14*ic_cap*ic_cap+2.50000e-14*ic_cap+1.23000e-11'
+ mcm4d_cf_w_0_300_s_0_300 = '-9.37500e-16*ic_cap*ic_cap+-1.25000e-15*ic_cap+1.39000e-12'
+ mcm4d_cf_w_0_300_s_0_360 = '-3.43750e-15*ic_cap*ic_cap+-3.75000e-15*ic_cap+1.67000e-12'
+ mcm4d_cf_w_0_300_s_0_450 = '-6.87500e-15*ic_cap*ic_cap+-5.00000e-15*ic_cap+2.10000e-12'
+ mcm4d_cf_w_0_300_s_0_600 = '-1.21875e-14*ic_cap*ic_cap+-8.75000e-15*ic_cap+2.80000e-12'
+ mcm4d_cf_w_0_300_s_0_800 = '-1.93750e-14*ic_cap*ic_cap+-1.25000e-14*ic_cap+3.63000e-12'
+ mcm4d_cf_w_0_300_s_1_000 = '-2.68750e-14*ic_cap*ic_cap+-1.75000e-14*ic_cap+4.49000e-12'
+ mcm4d_cf_w_0_300_s_1_200 = '-3.34375e-14*ic_cap*ic_cap+-2.12500e-14*ic_cap+5.34000e-12'
+ mcm4d_cf_w_0_300_s_2_100 = '-5.93750e-14*ic_cap*ic_cap+-3.75000e-14*ic_cap+9.13000e-12'
+ mcm4d_cf_w_0_300_s_3_300 = '-8.43750e-14*ic_cap*ic_cap+-6.25000e-14*ic_cap+1.29000e-11'
+ mcm4d_cf_w_0_300_s_9_000 = '-1.40625e-13*ic_cap*ic_cap+-8.75000e-14*ic_cap+2.42000e-11'
+ mcm4d_cf_w_2_400_s_0_300 = '-1.56250e-15*ic_cap*ic_cap+-1.25000e-15*ic_cap+1.42000e-12'
+ mcm4d_cf_w_2_400_s_0_360 = '-3.75000e-15*ic_cap*ic_cap+-2.50000e-15*ic_cap+1.69000e-12'
+ mcm4d_cf_w_2_400_s_0_450 = '-6.87500e-15*ic_cap*ic_cap+-5.00000e-15*ic_cap+2.10000e-12'
+ mcm4d_cf_w_2_400_s_0_600 = '-1.25000e-14*ic_cap*ic_cap+-7.50000e-15*ic_cap+2.78000e-12'
+ mcm4d_cf_w_2_400_s_0_800 = '-1.96875e-14*ic_cap*ic_cap+-1.37500e-14*ic_cap+3.67000e-12'
+ mcm4d_cf_w_2_400_s_1_000 = '-2.68750e-14*ic_cap*ic_cap+-1.75000e-14*ic_cap+4.54000e-12'
+ mcm4d_cf_w_2_400_s_1_200 = '-3.40625e-14*ic_cap*ic_cap+-2.12500e-14*ic_cap+5.40000e-12'
+ mcm4d_cf_w_2_400_s_2_100 = '-6.03125e-14*ic_cap*ic_cap+-3.87500e-14*ic_cap+9.02000e-12'
+ mcm4d_cf_w_2_400_s_3_300 = '-9.06250e-14*ic_cap*ic_cap+-6.25000e-14*ic_cap+1.33000e-11'
+ mcm4d_cf_w_2_400_s_9_000 = '-1.43750e-13*ic_cap*ic_cap+-1.00000e-13*ic_cap+2.63000e-11'
+ mcm4f_ca_w_0_300_s_0_300 = '-7.50000e-08*ic_cap*ic_cap+-4.75000e-08*ic_cap+8.67000e-06'
+ mcm4f_ca_w_0_300_s_0_360 = '-7.50000e-08*ic_cap*ic_cap+-4.75000e-08*ic_cap+8.67000e-06'
+ mcm4f_ca_w_0_300_s_0_450 = '-7.50000e-08*ic_cap*ic_cap+-4.75000e-08*ic_cap+8.67000e-06'
+ mcm4f_ca_w_0_300_s_0_600 = '-7.50000e-08*ic_cap*ic_cap+-4.75000e-08*ic_cap+8.67000e-06'
+ mcm4f_ca_w_0_300_s_0_800 = '-7.50000e-08*ic_cap*ic_cap+-4.75000e-08*ic_cap+8.67000e-06'
+ mcm4f_ca_w_0_300_s_1_000 = '-7.50000e-08*ic_cap*ic_cap+-4.75000e-08*ic_cap+8.67000e-06'
+ mcm4f_ca_w_0_300_s_1_200 = '-7.50000e-08*ic_cap*ic_cap+-4.75000e-08*ic_cap+8.67000e-06'
+ mcm4f_ca_w_0_300_s_2_100 = '-7.50000e-08*ic_cap*ic_cap+-4.75000e-08*ic_cap+8.67000e-06'
+ mcm4f_ca_w_0_300_s_3_300 = '-7.50000e-08*ic_cap*ic_cap+-4.75000e-08*ic_cap+8.67000e-06'
+ mcm4f_ca_w_0_300_s_9_000 = '-7.50000e-08*ic_cap*ic_cap+-4.75000e-08*ic_cap+8.67000e-06'
+ mcm4f_ca_w_2_400_s_0_300 = '-7.50000e-08*ic_cap*ic_cap+-4.75000e-08*ic_cap+8.67000e-06'
+ mcm4f_ca_w_2_400_s_0_360 = '-7.50000e-08*ic_cap*ic_cap+-4.75000e-08*ic_cap+8.67000e-06'
+ mcm4f_ca_w_2_400_s_0_450 = '-7.50000e-08*ic_cap*ic_cap+-4.75000e-08*ic_cap+8.67000e-06'
+ mcm4f_ca_w_2_400_s_0_600 = '-7.50000e-08*ic_cap*ic_cap+-4.75000e-08*ic_cap+8.67000e-06'
+ mcm4f_ca_w_2_400_s_0_800 = '-7.50000e-08*ic_cap*ic_cap+-4.75000e-08*ic_cap+8.67000e-06'
+ mcm4f_ca_w_2_400_s_1_000 = '-7.50000e-08*ic_cap*ic_cap+-4.75000e-08*ic_cap+8.67000e-06'
+ mcm4f_ca_w_2_400_s_1_200 = '-7.50000e-08*ic_cap*ic_cap+-4.75000e-08*ic_cap+8.67000e-06'
+ mcm4f_ca_w_2_400_s_2_100 = '-7.50000e-08*ic_cap*ic_cap+-4.75000e-08*ic_cap+8.67000e-06'
+ mcm4f_ca_w_2_400_s_3_300 = '-7.50000e-08*ic_cap*ic_cap+-4.75000e-08*ic_cap+8.67000e-06'
+ mcm4f_ca_w_2_400_s_9_000 = '-7.50000e-08*ic_cap*ic_cap+-4.75000e-08*ic_cap+8.67000e-06'
+ mcm4f_cc_w_0_300_s_0_300 = '-8.21875e-13*ic_cap*ic_cap+-4.87500e-13*ic_cap+1.08000e-10'
+ mcm4f_cc_w_0_300_s_0_360 = '-7.37500e-13*ic_cap*ic_cap+-4.50000e-13*ic_cap+1.01000e-10'
+ mcm4f_cc_w_0_300_s_0_450 = '-6.28125e-13*ic_cap*ic_cap+-3.62500e-13*ic_cap+9.17000e-11'
+ mcm4f_cc_w_0_300_s_0_600 = '-4.96875e-13*ic_cap*ic_cap+-3.12500e-13*ic_cap+7.96000e-11'
+ mcm4f_cc_w_0_300_s_0_800 = '-3.65625e-13*ic_cap*ic_cap+-2.37500e-13*ic_cap+6.78000e-11'
+ mcm4f_cc_w_0_300_s_1_000 = '-2.84375e-13*ic_cap*ic_cap+-1.87500e-13*ic_cap+5.90000e-11'
+ mcm4f_cc_w_0_300_s_1_200 = '-2.28125e-13*ic_cap*ic_cap+-1.37500e-13*ic_cap+5.24000e-11'
+ mcm4f_cc_w_0_300_s_2_100 = '-1.12500e-13*ic_cap*ic_cap+-7.50000e-14*ic_cap+3.60000e-11'
+ mcm4f_cc_w_0_300_s_3_300 = '-4.37500e-14*ic_cap*ic_cap+-2.50000e-14*ic_cap+2.59000e-11'
+ mcm4f_cc_w_0_300_s_9_000 = '1.96875e-14*ic_cap*ic_cap+1.37500e-14*ic_cap+8.98000e-12'
+ mcm4f_cc_w_2_400_s_0_300 = '-8.12500e-13*ic_cap*ic_cap+-5.00000e-13*ic_cap+1.36000e-10'
+ mcm4f_cc_w_2_400_s_0_360 = '-7.18750e-13*ic_cap*ic_cap+-3.75000e-13*ic_cap+1.28000e-10'
+ mcm4f_cc_w_2_400_s_0_450 = '-5.93750e-13*ic_cap*ic_cap+-3.75000e-13*ic_cap+1.17000e-10'
+ mcm4f_cc_w_2_400_s_0_600 = '-4.43750e-13*ic_cap*ic_cap+-2.75000e-13*ic_cap+1.02000e-10'
+ mcm4f_cc_w_2_400_s_0_800 = '-3.31250e-13*ic_cap*ic_cap+-2.00000e-13*ic_cap+8.75000e-11'
+ mcm4f_cc_w_2_400_s_1_000 = '-2.43750e-13*ic_cap*ic_cap+-1.75000e-13*ic_cap+7.66000e-11'
+ mcm4f_cc_w_2_400_s_1_200 = '-1.84375e-13*ic_cap*ic_cap+-1.37500e-13*ic_cap+6.84000e-11'
+ mcm4f_cc_w_2_400_s_2_100 = '-7.18750e-14*ic_cap*ic_cap+-3.75000e-14*ic_cap+4.77000e-11'
+ mcm4f_cc_w_2_400_s_3_300 = '-9.37500e-15*ic_cap*ic_cap+-1.25000e-14*ic_cap+3.44000e-11'
+ mcm4f_cc_w_2_400_s_9_000 = '4.06250e-14*ic_cap*ic_cap+1.25000e-14*ic_cap+1.29000e-11'
+ mcm4f_cf_w_0_300_s_0_300 = '-2.18750e-15*ic_cap*ic_cap+-1.25000e-15*ic_cap+1.29000e-12'
+ mcm4f_cf_w_0_300_s_0_360 = '-4.06250e-15*ic_cap*ic_cap+-3.75000e-15*ic_cap+1.54000e-12'
+ mcm4f_cf_w_0_300_s_0_450 = '-7.50000e-15*ic_cap*ic_cap+-5.00000e-15*ic_cap+1.94000e-12'
+ mcm4f_cf_w_0_300_s_0_600 = '-1.25000e-14*ic_cap*ic_cap+-7.50000e-15*ic_cap+2.59000e-12'
+ mcm4f_cf_w_0_300_s_0_800 = '-1.90625e-14*ic_cap*ic_cap+-1.12500e-14*ic_cap+3.35000e-12'
+ mcm4f_cf_w_0_300_s_1_000 = '-2.71875e-14*ic_cap*ic_cap+-1.62500e-14*ic_cap+4.16000e-12'
+ mcm4f_cf_w_0_300_s_1_200 = '-3.34375e-14*ic_cap*ic_cap+-2.12500e-14*ic_cap+4.94000e-12'
+ mcm4f_cf_w_0_300_s_2_100 = '-5.84375e-14*ic_cap*ic_cap+-3.87500e-14*ic_cap+8.49000e-12'
+ mcm4f_cf_w_0_300_s_3_300 = '-8.75000e-14*ic_cap*ic_cap+-5.00000e-14*ic_cap+1.21000e-11'
+ mcm4f_cf_w_0_300_s_9_000 = '-1.43750e-13*ic_cap*ic_cap+-1.00000e-13*ic_cap+2.31000e-11'
+ mcm4f_cf_w_2_400_s_0_300 = '-2.50000e-15*ic_cap*ic_cap+-2.50000e-15*ic_cap+1.31000e-12'
+ mcm4f_cf_w_2_400_s_0_360 = '-4.37500e-15*ic_cap*ic_cap+-2.50000e-15*ic_cap+1.56000e-12'
+ mcm4f_cf_w_2_400_s_0_450 = '-7.50000e-15*ic_cap*ic_cap+-5.00000e-15*ic_cap+1.94000e-12'
+ mcm4f_cf_w_2_400_s_0_600 = '-1.34375e-14*ic_cap*ic_cap+-8.75000e-15*ic_cap+2.57000e-12'
+ mcm4f_cf_w_2_400_s_0_800 = '-2.00000e-14*ic_cap*ic_cap+-1.25000e-14*ic_cap+3.39000e-12'
+ mcm4f_cf_w_2_400_s_1_000 = '-2.65625e-14*ic_cap*ic_cap+-1.62500e-14*ic_cap+4.20000e-12'
+ mcm4f_cf_w_2_400_s_1_200 = '-3.34375e-14*ic_cap*ic_cap+-2.12500e-14*ic_cap+4.99000e-12'
+ mcm4f_cf_w_2_400_s_2_100 = '-6.00000e-14*ic_cap*ic_cap+-3.75000e-14*ic_cap+8.38000e-12'
+ mcm4f_cf_w_2_400_s_3_300 = '-8.75000e-14*ic_cap*ic_cap+-5.00000e-14*ic_cap+1.24000e-11'
+ mcm4f_cf_w_2_400_s_9_000 = '-1.50000e-13*ic_cap*ic_cap+-1.00000e-13*ic_cap+2.51000e-11'
+ mcm4l1_ca_w_0_300_s_0_300 = '-9.62500e-08*ic_cap*ic_cap+-6.00000e-08*ic_cap+1.17000e-05'
+ mcm4l1_ca_w_0_300_s_0_360 = '-9.62500e-08*ic_cap*ic_cap+-6.00000e-08*ic_cap+1.17000e-05'
+ mcm4l1_ca_w_0_300_s_0_450 = '-9.62500e-08*ic_cap*ic_cap+-6.00000e-08*ic_cap+1.17000e-05'
+ mcm4l1_ca_w_0_300_s_0_600 = '-9.62500e-08*ic_cap*ic_cap+-6.00000e-08*ic_cap+1.17000e-05'
+ mcm4l1_ca_w_0_300_s_0_800 = '-9.62500e-08*ic_cap*ic_cap+-6.00000e-08*ic_cap+1.17000e-05'
+ mcm4l1_ca_w_0_300_s_1_000 = '-9.62500e-08*ic_cap*ic_cap+-6.00000e-08*ic_cap+1.17000e-05'
+ mcm4l1_ca_w_0_300_s_1_200 = '-9.62500e-08*ic_cap*ic_cap+-6.00000e-08*ic_cap+1.17000e-05'
+ mcm4l1_ca_w_0_300_s_2_100 = '-9.62500e-08*ic_cap*ic_cap+-6.00000e-08*ic_cap+1.17000e-05'
+ mcm4l1_ca_w_0_300_s_3_300 = '-9.62500e-08*ic_cap*ic_cap+-6.00000e-08*ic_cap+1.17000e-05'
+ mcm4l1_ca_w_0_300_s_9_000 = '-9.62500e-08*ic_cap*ic_cap+-6.00000e-08*ic_cap+1.17000e-05'
+ mcm4l1_ca_w_2_400_s_0_300 = '-9.62500e-08*ic_cap*ic_cap+-6.00000e-08*ic_cap+1.17000e-05'
+ mcm4l1_ca_w_2_400_s_0_360 = '-9.62500e-08*ic_cap*ic_cap+-6.00000e-08*ic_cap+1.17000e-05'
+ mcm4l1_ca_w_2_400_s_0_450 = '-9.62500e-08*ic_cap*ic_cap+-6.00000e-08*ic_cap+1.17000e-05'
+ mcm4l1_ca_w_2_400_s_0_600 = '-9.62500e-08*ic_cap*ic_cap+-6.00000e-08*ic_cap+1.17000e-05'
+ mcm4l1_ca_w_2_400_s_0_800 = '-9.62500e-08*ic_cap*ic_cap+-6.00000e-08*ic_cap+1.17000e-05'
+ mcm4l1_ca_w_2_400_s_1_000 = '-9.62500e-08*ic_cap*ic_cap+-6.00000e-08*ic_cap+1.17000e-05'
+ mcm4l1_ca_w_2_400_s_1_200 = '-9.62500e-08*ic_cap*ic_cap+-6.00000e-08*ic_cap+1.17000e-05'
+ mcm4l1_ca_w_2_400_s_2_100 = '-9.62500e-08*ic_cap*ic_cap+-6.00000e-08*ic_cap+1.17000e-05'
+ mcm4l1_ca_w_2_400_s_3_300 = '-9.62500e-08*ic_cap*ic_cap+-6.00000e-08*ic_cap+1.17000e-05'
+ mcm4l1_ca_w_2_400_s_9_000 = '-9.62500e-08*ic_cap*ic_cap+-6.00000e-08*ic_cap+1.17000e-05'
+ mcm4l1_cc_w_0_300_s_0_300 = '-8.68750e-13*ic_cap*ic_cap+-4.75000e-13*ic_cap+1.08000e-10'
+ mcm4l1_cc_w_0_300_s_0_360 = '-7.18750e-13*ic_cap*ic_cap+-4.25000e-13*ic_cap+1.00000e-10'
+ mcm4l1_cc_w_0_300_s_0_450 = '-6.15625e-13*ic_cap*ic_cap+-3.62500e-13*ic_cap+9.07000e-11'
+ mcm4l1_cc_w_0_300_s_0_600 = '-4.87500e-13*ic_cap*ic_cap+-3.00000e-13*ic_cap+7.85000e-11'
+ mcm4l1_cc_w_0_300_s_0_800 = '-3.53125e-13*ic_cap*ic_cap+-2.37500e-13*ic_cap+6.65000e-11'
+ mcm4l1_cc_w_0_300_s_1_000 = '-2.81250e-13*ic_cap*ic_cap+-1.75000e-13*ic_cap+5.76000e-11'
+ mcm4l1_cc_w_0_300_s_1_200 = '-2.18750e-13*ic_cap*ic_cap+-1.50000e-13*ic_cap+5.08000e-11'
+ mcm4l1_cc_w_0_300_s_2_100 = '-9.68750e-14*ic_cap*ic_cap+-6.25000e-14*ic_cap+3.38000e-11'
+ mcm4l1_cc_w_0_300_s_3_300 = '-3.75000e-14*ic_cap*ic_cap+-2.50000e-14*ic_cap+2.35000e-11'
+ mcm4l1_cc_w_0_300_s_9_000 = '1.43750e-14*ic_cap*ic_cap+1.25000e-14*ic_cap+7.13000e-12'
+ mcm4l1_cc_w_2_400_s_0_300 = '-8.12500e-13*ic_cap*ic_cap+-5.00000e-13*ic_cap+1.34000e-10'
+ mcm4l1_cc_w_2_400_s_0_360 = '-6.56250e-13*ic_cap*ic_cap+-3.75000e-13*ic_cap+1.25000e-10'
+ mcm4l1_cc_w_2_400_s_0_450 = '-5.93750e-13*ic_cap*ic_cap+-3.75000e-13*ic_cap+1.14000e-10'
+ mcm4l1_cc_w_2_400_s_0_600 = '-4.53125e-13*ic_cap*ic_cap+-2.62500e-13*ic_cap+9.95000e-11'
+ mcm4l1_cc_w_2_400_s_0_800 = '-3.18750e-13*ic_cap*ic_cap+-2.00000e-13*ic_cap+8.47000e-11'
+ mcm4l1_cc_w_2_400_s_1_000 = '-2.37500e-13*ic_cap*ic_cap+-1.50000e-13*ic_cap+7.38000e-11'
+ mcm4l1_cc_w_2_400_s_1_200 = '-1.84375e-13*ic_cap*ic_cap+-1.12500e-13*ic_cap+6.56000e-11'
+ mcm4l1_cc_w_2_400_s_2_100 = '-6.56250e-14*ic_cap*ic_cap+-3.75000e-14*ic_cap+4.47000e-11'
+ mcm4l1_cc_w_2_400_s_3_300 = '-1.25000e-14*ic_cap*ic_cap+3.14000e-11'
+ mcm4l1_cc_w_2_400_s_9_000 = '2.50000e-14*ic_cap*ic_cap+2.50000e-14*ic_cap+1.07000e-11'
+ mcm4l1_cf_w_0_300_s_0_300 = '-1.56250e-15*ic_cap*ic_cap+-1.25000e-15*ic_cap+1.73000e-12'
+ mcm4l1_cf_w_0_300_s_0_360 = '-4.37500e-15*ic_cap*ic_cap+-2.50000e-15*ic_cap+2.07000e-12'
+ mcm4l1_cf_w_0_300_s_0_450 = '-8.43750e-15*ic_cap*ic_cap+-6.25000e-15*ic_cap+2.60000e-12'
+ mcm4l1_cf_w_0_300_s_0_600 = '-1.50000e-14*ic_cap*ic_cap+-1.00000e-14*ic_cap+3.46000e-12'
+ mcm4l1_cf_w_0_300_s_0_800 = '-2.40625e-14*ic_cap*ic_cap+-1.62500e-14*ic_cap+4.48000e-12'
+ mcm4l1_cf_w_0_300_s_1_000 = '-3.31250e-14*ic_cap*ic_cap+-2.25000e-14*ic_cap+5.53000e-12'
+ mcm4l1_cf_w_0_300_s_1_200 = '-4.03125e-14*ic_cap*ic_cap+-2.62500e-14*ic_cap+6.55000e-12'
+ mcm4l1_cf_w_0_300_s_2_100 = '-6.81250e-14*ic_cap*ic_cap+-4.75000e-14*ic_cap+1.10000e-11'
+ mcm4l1_cf_w_0_300_s_3_300 = '-1.03125e-13*ic_cap*ic_cap+-6.25000e-14*ic_cap+1.55000e-11'
+ mcm4l1_cf_w_0_300_s_9_000 = '-1.53125e-13*ic_cap*ic_cap+-1.12500e-13*ic_cap+2.73000e-11'
+ mcm4l1_cf_w_2_400_s_0_300 = '-1.87500e-15*ic_cap*ic_cap+-2.50000e-15*ic_cap+1.75000e-12'
+ mcm4l1_cf_w_2_400_s_0_360 = '-4.68750e-15*ic_cap*ic_cap+-3.75000e-15*ic_cap+2.09000e-12'
+ mcm4l1_cf_w_2_400_s_0_450 = '-9.06250e-15*ic_cap*ic_cap+-6.25000e-15*ic_cap+2.60000e-12'
+ mcm4l1_cf_w_2_400_s_0_600 = '-1.56250e-14*ic_cap*ic_cap+-1.00000e-14*ic_cap+3.43000e-12'
+ mcm4l1_cf_w_2_400_s_0_800 = '-2.40625e-14*ic_cap*ic_cap+-1.62500e-14*ic_cap+4.52000e-12'
+ mcm4l1_cf_w_2_400_s_1_000 = '-3.25000e-14*ic_cap*ic_cap+-2.25000e-14*ic_cap+5.58000e-12'
+ mcm4l1_cf_w_2_400_s_1_200 = '-4.06250e-14*ic_cap*ic_cap+-2.75000e-14*ic_cap+6.62000e-12'
+ mcm4l1_cf_w_2_400_s_2_100 = '-7.43750e-14*ic_cap*ic_cap+-4.75000e-14*ic_cap+1.10000e-11'
+ mcm4l1_cf_w_2_400_s_3_300 = '-1.06250e-13*ic_cap*ic_cap+-7.50000e-14*ic_cap+1.60000e-11'
+ mcm4l1_cf_w_2_400_s_9_000 = '-1.53125e-13*ic_cap*ic_cap+-1.12500e-13*ic_cap+2.98000e-11'
+ mcm4l1d_ca_w_0_170_s_0_180 = '-6.46875e-07*ic_cap*ic_cap+-3.62500e-07*ic_cap+6.70000e-05'
+ mcm4l1d_ca_w_0_170_s_0_225 = '-6.46875e-07*ic_cap*ic_cap+-3.62500e-07*ic_cap+6.70000e-05'
+ mcm4l1d_ca_w_0_170_s_0_270 = '-6.46875e-07*ic_cap*ic_cap+-3.62500e-07*ic_cap+6.70000e-05'
+ mcm4l1d_ca_w_0_170_s_0_360 = '-6.46875e-07*ic_cap*ic_cap+-3.62500e-07*ic_cap+6.70000e-05'
+ mcm4l1d_ca_w_0_170_s_0_450 = '-6.46875e-07*ic_cap*ic_cap+-3.62500e-07*ic_cap+6.70000e-05'
+ mcm4l1d_ca_w_0_170_s_0_540 = '-6.46875e-07*ic_cap*ic_cap+-3.62500e-07*ic_cap+6.70000e-05'
+ mcm4l1d_ca_w_0_170_s_0_720 = '-6.46875e-07*ic_cap*ic_cap+-3.62500e-07*ic_cap+6.70000e-05'
+ mcm4l1d_ca_w_0_170_s_1_080 = '-6.46875e-07*ic_cap*ic_cap+-3.62500e-07*ic_cap+6.70000e-05'
+ mcm4l1d_ca_w_0_170_s_1_980 = '-6.46875e-07*ic_cap*ic_cap+-3.62500e-07*ic_cap+6.70000e-05'
+ mcm4l1d_ca_w_0_170_s_4_500 = '-6.46875e-07*ic_cap*ic_cap+-3.62500e-07*ic_cap+6.70000e-05'
+ mcm4l1d_ca_w_1_360_s_0_180 = '-6.46875e-07*ic_cap*ic_cap+-3.62500e-07*ic_cap+6.70000e-05'
+ mcm4l1d_ca_w_1_360_s_0_225 = '-6.46875e-07*ic_cap*ic_cap+-3.62500e-07*ic_cap+6.70000e-05'
+ mcm4l1d_ca_w_1_360_s_0_270 = '-6.46875e-07*ic_cap*ic_cap+-3.62500e-07*ic_cap+6.70000e-05'
+ mcm4l1d_ca_w_1_360_s_0_360 = '-6.46875e-07*ic_cap*ic_cap+-3.62500e-07*ic_cap+6.70000e-05'
+ mcm4l1d_ca_w_1_360_s_0_450 = '-6.46875e-07*ic_cap*ic_cap+-3.62500e-07*ic_cap+6.70000e-05'
+ mcm4l1d_ca_w_1_360_s_0_540 = '-6.46875e-07*ic_cap*ic_cap+-3.62500e-07*ic_cap+6.70000e-05'
+ mcm4l1d_ca_w_1_360_s_0_720 = '-6.46875e-07*ic_cap*ic_cap+-3.62500e-07*ic_cap+6.70000e-05'
+ mcm4l1d_ca_w_1_360_s_1_080 = '-6.46875e-07*ic_cap*ic_cap+-3.62500e-07*ic_cap+6.70000e-05'
+ mcm4l1d_ca_w_1_360_s_1_980 = '-6.46875e-07*ic_cap*ic_cap+-3.62500e-07*ic_cap+6.70000e-05'
+ mcm4l1d_ca_w_1_360_s_4_500 = '-6.46875e-07*ic_cap*ic_cap+-3.62500e-07*ic_cap+6.70000e-05'
+ mcm4l1d_cc_w_0_170_s_0_180 = '-7.68750e-13*ic_cap*ic_cap+-5.00000e-13*ic_cap+7.59000e-11'
+ mcm4l1d_cc_w_0_170_s_0_225 = '-5.50000e-13*ic_cap*ic_cap+-3.75000e-13*ic_cap+6.39000e-11'
+ mcm4l1d_cc_w_0_170_s_0_270 = '-4.12500e-13*ic_cap*ic_cap+-3.00000e-13*ic_cap+5.58000e-11'
+ mcm4l1d_cc_w_0_170_s_0_360 = '-2.62500e-13*ic_cap*ic_cap+-2.00000e-13*ic_cap+4.42000e-11'
+ mcm4l1d_cc_w_0_170_s_0_450 = '-1.71875e-13*ic_cap*ic_cap+-1.37500e-13*ic_cap+3.68000e-11'
+ mcm4l1d_cc_w_0_170_s_0_540 = '-1.12500e-13*ic_cap*ic_cap+-1.00000e-13*ic_cap+3.09000e-11'
+ mcm4l1d_cc_w_0_170_s_0_720 = '-4.68750e-14*ic_cap*ic_cap+-6.25000e-14*ic_cap+2.31000e-11'
+ mcm4l1d_cc_w_0_170_s_1_080 = '9.37500e-15*ic_cap*ic_cap+-1.25000e-14*ic_cap+1.40000e-11'
+ mcm4l1d_cc_w_0_170_s_1_980 = '3.37500e-14*ic_cap*ic_cap+1.50000e-14*ic_cap+4.91000e-12'
+ mcm4l1d_cc_w_0_170_s_4_500 = '1.12500e-14*ic_cap*ic_cap+7.50000e-15*ic_cap+4.70000e-13'
+ mcm4l1d_cc_w_1_360_s_0_180 = '-6.56250e-13*ic_cap*ic_cap+-4.25000e-13*ic_cap+9.01000e-11'
+ mcm4l1d_cc_w_1_360_s_0_225 = '-4.37500e-13*ic_cap*ic_cap+-3.00000e-13*ic_cap+7.69000e-11'
+ mcm4l1d_cc_w_1_360_s_0_270 = '-3.06250e-13*ic_cap*ic_cap+-2.25000e-13*ic_cap+6.75000e-11'
+ mcm4l1d_cc_w_1_360_s_0_360 = '-1.62500e-13*ic_cap*ic_cap+-1.25000e-13*ic_cap+5.45000e-11'
+ mcm4l1d_cc_w_1_360_s_0_450 = '-8.12500e-14*ic_cap*ic_cap+-7.50000e-14*ic_cap+4.57000e-11'
+ mcm4l1d_cc_w_1_360_s_0_540 = '-3.12500e-14*ic_cap*ic_cap+-5.00000e-14*ic_cap+3.92000e-11'
+ mcm4l1d_cc_w_1_360_s_0_720 = '3.12500e-14*ic_cap*ic_cap+2.99000e-11'
+ mcm4l1d_cc_w_1_360_s_1_080 = '7.18750e-14*ic_cap*ic_cap+3.75000e-14*ic_cap+1.90000e-11'
+ mcm4l1d_cc_w_1_360_s_1_980 = '7.31250e-14*ic_cap*ic_cap+4.00000e-14*ic_cap+7.34000e-12'
+ mcm4l1d_cc_w_1_360_s_4_500 = '2.31250e-14*ic_cap*ic_cap+2.00000e-14*ic_cap+7.80000e-13'
+ mcm4l1d_cf_w_0_170_s_0_180 = '-7.81250e-15*ic_cap*ic_cap+-3.75000e-15*ic_cap+5.86000e-12'
+ mcm4l1d_cf_w_0_170_s_0_225 = '-2.18750e-14*ic_cap*ic_cap+-1.25000e-14*ic_cap+7.26000e-12'
+ mcm4l1d_cf_w_0_170_s_0_270 = '-3.59375e-14*ic_cap*ic_cap+-2.12500e-14*ic_cap+8.60000e-12'
+ mcm4l1d_cf_w_0_170_s_0_360 = '-6.25000e-14*ic_cap*ic_cap+-2.50000e-14*ic_cap+1.14000e-11'
+ mcm4l1d_cf_w_0_170_s_0_450 = '-8.12500e-14*ic_cap*ic_cap+-5.00000e-14*ic_cap+1.36000e-11'
+ mcm4l1d_cf_w_0_170_s_0_540 = '-1.09375e-13*ic_cap*ic_cap+-6.25000e-14*ic_cap+1.61000e-11'
+ mcm4l1d_cf_w_0_170_s_0_720 = '-1.40625e-13*ic_cap*ic_cap+-8.75000e-14*ic_cap+2.00000e-11'
+ mcm4l1d_cf_w_0_170_s_1_080 = '-1.84375e-13*ic_cap*ic_cap+-1.12500e-13*ic_cap+2.60000e-11'
+ mcm4l1d_cf_w_0_170_s_1_980 = '-2.15625e-13*ic_cap*ic_cap+-1.37500e-13*ic_cap+3.35000e-11'
+ mcm4l1d_cf_w_0_170_s_4_500 = '-1.93750e-13*ic_cap*ic_cap+-1.25000e-13*ic_cap+3.76000e-11'
+ mcm4l1d_cf_w_1_360_s_0_180 = '-7.81250e-15*ic_cap*ic_cap+-3.75000e-15*ic_cap+5.85000e-12'
+ mcm4l1d_cf_w_1_360_s_0_225 = '-2.18750e-14*ic_cap*ic_cap+-1.00000e-14*ic_cap+7.25000e-12'
+ mcm4l1d_cf_w_1_360_s_0_270 = '-3.53125e-14*ic_cap*ic_cap+-1.87500e-14*ic_cap+8.62000e-12'
+ mcm4l1d_cf_w_1_360_s_0_360 = '-5.93750e-14*ic_cap*ic_cap+-3.75000e-14*ic_cap+1.12000e-11'
+ mcm4l1d_cf_w_1_360_s_0_450 = '-8.12500e-14*ic_cap*ic_cap+-5.00000e-14*ic_cap+1.37000e-11'
+ mcm4l1d_cf_w_1_360_s_0_540 = '-1.06250e-13*ic_cap*ic_cap+-5.00000e-14*ic_cap+1.61000e-11'
+ mcm4l1d_cf_w_1_360_s_0_720 = '-1.37500e-13*ic_cap*ic_cap+-7.50000e-14*ic_cap+2.02000e-11'
+ mcm4l1d_cf_w_1_360_s_1_080 = '-1.78125e-13*ic_cap*ic_cap+-1.12500e-13*ic_cap+2.68000e-11'
+ mcm4l1d_cf_w_1_360_s_1_980 = '-2.00000e-13*ic_cap*ic_cap+-1.25000e-13*ic_cap+3.60000e-11'
+ mcm4l1d_cf_w_1_360_s_4_500 = '-1.62500e-13*ic_cap*ic_cap+-1.00000e-13*ic_cap+4.22000e-11'
+ mcm4l1f_ca_w_0_170_s_0_180 = '-5.09375e-07*ic_cap*ic_cap+-2.87500e-07*ic_cap+4.86000e-05'
+ mcm4l1f_ca_w_0_170_s_0_225 = '-5.09375e-07*ic_cap*ic_cap+-2.87500e-07*ic_cap+4.86000e-05'
+ mcm4l1f_ca_w_0_170_s_0_270 = '-5.09375e-07*ic_cap*ic_cap+-2.87500e-07*ic_cap+4.86000e-05'
+ mcm4l1f_ca_w_0_170_s_0_360 = '-5.09375e-07*ic_cap*ic_cap+-2.87500e-07*ic_cap+4.86000e-05'
+ mcm4l1f_ca_w_0_170_s_0_450 = '-5.09375e-07*ic_cap*ic_cap+-2.87500e-07*ic_cap+4.86000e-05'
+ mcm4l1f_ca_w_0_170_s_0_540 = '-5.09375e-07*ic_cap*ic_cap+-2.87500e-07*ic_cap+4.86000e-05'
+ mcm4l1f_ca_w_0_170_s_0_720 = '-5.09375e-07*ic_cap*ic_cap+-2.87500e-07*ic_cap+4.86000e-05'
+ mcm4l1f_ca_w_0_170_s_1_080 = '-5.09375e-07*ic_cap*ic_cap+-2.87500e-07*ic_cap+4.86000e-05'
+ mcm4l1f_ca_w_0_170_s_1_980 = '-5.09375e-07*ic_cap*ic_cap+-2.87500e-07*ic_cap+4.86000e-05'
+ mcm4l1f_ca_w_0_170_s_4_500 = '-5.09375e-07*ic_cap*ic_cap+-2.87500e-07*ic_cap+4.86000e-05'
+ mcm4l1f_ca_w_1_360_s_0_180 = '-5.09375e-07*ic_cap*ic_cap+-2.87500e-07*ic_cap+4.86000e-05'
+ mcm4l1f_ca_w_1_360_s_0_225 = '-5.09375e-07*ic_cap*ic_cap+-2.87500e-07*ic_cap+4.86000e-05'
+ mcm4l1f_ca_w_1_360_s_0_270 = '-5.09375e-07*ic_cap*ic_cap+-2.87500e-07*ic_cap+4.86000e-05'
+ mcm4l1f_ca_w_1_360_s_0_360 = '-5.09375e-07*ic_cap*ic_cap+-2.87500e-07*ic_cap+4.86000e-05'
+ mcm4l1f_ca_w_1_360_s_0_450 = '-5.09375e-07*ic_cap*ic_cap+-2.87500e-07*ic_cap+4.86000e-05'
+ mcm4l1f_ca_w_1_360_s_0_540 = '-5.09375e-07*ic_cap*ic_cap+-2.87500e-07*ic_cap+4.86000e-05'
+ mcm4l1f_ca_w_1_360_s_0_720 = '-5.09375e-07*ic_cap*ic_cap+-2.87500e-07*ic_cap+4.86000e-05'
+ mcm4l1f_ca_w_1_360_s_1_080 = '-5.09375e-07*ic_cap*ic_cap+-2.87500e-07*ic_cap+4.86000e-05'
+ mcm4l1f_ca_w_1_360_s_1_980 = '-5.09375e-07*ic_cap*ic_cap+-2.87500e-07*ic_cap+4.86000e-05'
+ mcm4l1f_ca_w_1_360_s_4_500 = '-5.09375e-07*ic_cap*ic_cap+-2.87500e-07*ic_cap+4.86000e-05'
+ mcm4l1f_cc_w_0_170_s_0_180 = '-7.78125e-13*ic_cap*ic_cap+-5.12500e-13*ic_cap+7.83000e-11'
+ mcm4l1f_cc_w_0_170_s_0_225 = '-5.75000e-13*ic_cap*ic_cap+-3.75000e-13*ic_cap+6.66000e-11'
+ mcm4l1f_cc_w_0_170_s_0_270 = '-4.25000e-13*ic_cap*ic_cap+-3.00000e-13*ic_cap+5.85000e-11'
+ mcm4l1f_cc_w_0_170_s_0_360 = '-2.75000e-13*ic_cap*ic_cap+-2.00000e-13*ic_cap+4.72000e-11'
+ mcm4l1f_cc_w_0_170_s_0_450 = '-1.81250e-13*ic_cap*ic_cap+-1.50000e-13*ic_cap+4.00000e-11'
+ mcm4l1f_cc_w_0_170_s_0_540 = '-1.28125e-13*ic_cap*ic_cap+-1.12500e-13*ic_cap+3.43000e-11'
+ mcm4l1f_cc_w_0_170_s_0_720 = '-5.62500e-14*ic_cap*ic_cap+-5.00000e-14*ic_cap+2.66000e-11'
+ mcm4l1f_cc_w_0_170_s_1_080 = '9.37500e-15*ic_cap*ic_cap+-1.25000e-14*ic_cap+1.73000e-11'
+ mcm4l1f_cc_w_0_170_s_1_980 = '5.12500e-14*ic_cap*ic_cap+2.25000e-14*ic_cap+6.95000e-12'
+ mcm4l1f_cc_w_0_170_s_4_500 = '2.12500e-14*ic_cap*ic_cap+1.37500e-14*ic_cap+8.15000e-13'
+ mcm4l1f_cc_w_1_360_s_0_180 = '-6.46875e-13*ic_cap*ic_cap+-4.37500e-13*ic_cap+9.45000e-11'
+ mcm4l1f_cc_w_1_360_s_0_225 = '-4.15625e-13*ic_cap*ic_cap+-2.87500e-13*ic_cap+8.12000e-11'
+ mcm4l1f_cc_w_1_360_s_0_270 = '-2.96875e-13*ic_cap*ic_cap+-2.12500e-13*ic_cap+7.19000e-11'
+ mcm4l1f_cc_w_1_360_s_0_360 = '-1.46875e-13*ic_cap*ic_cap+-1.12500e-13*ic_cap+5.89000e-11'
+ mcm4l1f_cc_w_1_360_s_0_450 = '-6.25000e-14*ic_cap*ic_cap+-7.50000e-14*ic_cap+5.00000e-11'
+ mcm4l1f_cc_w_1_360_s_0_540 = '-1.56250e-14*ic_cap*ic_cap+-3.75000e-14*ic_cap+4.35000e-11'
+ mcm4l1f_cc_w_1_360_s_0_720 = '4.68750e-14*ic_cap*ic_cap+1.25000e-14*ic_cap+3.41000e-11'
+ mcm4l1f_cc_w_1_360_s_1_080 = '9.37500e-14*ic_cap*ic_cap+5.00000e-14*ic_cap+2.28000e-11'
+ mcm4l1f_cc_w_1_360_s_1_980 = '9.93750e-14*ic_cap*ic_cap+6.25000e-14*ic_cap+9.76000e-12'
+ mcm4l1f_cc_w_1_360_s_4_500 = '3.81250e-14*ic_cap*ic_cap+2.75000e-14*ic_cap+1.23000e-12'
+ mcm4l1f_cf_w_0_170_s_0_180 = '-1.00000e-14*ic_cap*ic_cap+-5.00000e-15*ic_cap+4.30000e-12'
+ mcm4l1f_cf_w_0_170_s_0_225 = '-2.21875e-14*ic_cap*ic_cap+-1.12500e-14*ic_cap+5.34000e-12'
+ mcm4l1f_cf_w_0_170_s_0_270 = '-3.18750e-14*ic_cap*ic_cap+-2.00000e-14*ic_cap+6.33000e-12'
+ mcm4l1f_cf_w_0_170_s_0_360 = '-5.34375e-14*ic_cap*ic_cap+-2.87500e-14*ic_cap+8.48000e-12'
+ mcm4l1f_cf_w_0_170_s_0_450 = '-7.46875e-14*ic_cap*ic_cap+-4.37500e-14*ic_cap+1.02000e-11'
+ mcm4l1f_cf_w_0_170_s_0_540 = '-8.75000e-14*ic_cap*ic_cap+-5.00000e-14*ic_cap+1.21000e-11'
+ mcm4l1f_cf_w_0_170_s_0_720 = '-1.25000e-13*ic_cap*ic_cap+-7.50000e-14*ic_cap+1.54000e-11'
+ mcm4l1f_cf_w_0_170_s_1_080 = '-1.68750e-13*ic_cap*ic_cap+-1.00000e-13*ic_cap+2.06000e-11'
+ mcm4l1f_cf_w_0_170_s_1_980 = '-2.09375e-13*ic_cap*ic_cap+-1.37500e-13*ic_cap+2.83000e-11'
+ mcm4l1f_cf_w_0_170_s_4_500 = '-1.93750e-13*ic_cap*ic_cap+-1.25000e-13*ic_cap+3.39000e-11'
+ mcm4l1f_cf_w_1_360_s_0_180 = '-1.03125e-14*ic_cap*ic_cap+-6.25000e-15*ic_cap+4.29000e-12'
+ mcm4l1f_cf_w_1_360_s_0_225 = '-2.09375e-14*ic_cap*ic_cap+-1.12500e-14*ic_cap+5.32000e-12'
+ mcm4l1f_cf_w_1_360_s_0_270 = '-3.18750e-14*ic_cap*ic_cap+-1.75000e-14*ic_cap+6.35000e-12'
+ mcm4l1f_cf_w_1_360_s_0_360 = '-5.21875e-14*ic_cap*ic_cap+-3.12500e-14*ic_cap+8.33000e-12'
+ mcm4l1f_cf_w_1_360_s_0_450 = '-6.87500e-14*ic_cap*ic_cap+-4.25000e-14*ic_cap+1.02000e-11'
+ mcm4l1f_cf_w_1_360_s_0_540 = '-9.37500e-14*ic_cap*ic_cap+-5.00000e-14*ic_cap+1.21000e-11'
+ mcm4l1f_cf_w_1_360_s_0_720 = '-1.18750e-13*ic_cap*ic_cap+-7.50000e-14*ic_cap+1.54000e-11'
+ mcm4l1f_cf_w_1_360_s_1_080 = '-1.62500e-13*ic_cap*ic_cap+-1.00000e-13*ic_cap+2.11000e-11'
+ mcm4l1f_cf_w_1_360_s_1_980 = '-2.00000e-13*ic_cap*ic_cap+-1.25000e-13*ic_cap+3.03000e-11'
+ mcm4l1f_cf_w_1_360_s_4_500 = '-1.62500e-13*ic_cap*ic_cap+-1.00000e-13*ic_cap+3.80000e-11'
+ mcm4l1p1_ca_w_0_170_s_0_180 = '-1.75938e-06*ic_cap*ic_cap+-8.62500e-07*ic_cap+1.06000e-04'
+ mcm4l1p1_ca_w_0_170_s_0_225 = '-1.75938e-06*ic_cap*ic_cap+-8.62500e-07*ic_cap+1.06000e-04'
+ mcm4l1p1_ca_w_0_170_s_0_270 = '-1.75938e-06*ic_cap*ic_cap+-8.62500e-07*ic_cap+1.06000e-04'
+ mcm4l1p1_ca_w_0_170_s_0_360 = '-1.75938e-06*ic_cap*ic_cap+-8.62500e-07*ic_cap+1.06000e-04'
+ mcm4l1p1_ca_w_0_170_s_0_450 = '-1.75938e-06*ic_cap*ic_cap+-8.62500e-07*ic_cap+1.06000e-04'
+ mcm4l1p1_ca_w_0_170_s_0_540 = '-1.75938e-06*ic_cap*ic_cap+-8.62500e-07*ic_cap+1.06000e-04'
+ mcm4l1p1_ca_w_0_170_s_0_720 = '-1.75938e-06*ic_cap*ic_cap+-8.62500e-07*ic_cap+1.06000e-04'
+ mcm4l1p1_ca_w_0_170_s_1_080 = '-1.75938e-06*ic_cap*ic_cap+-8.62500e-07*ic_cap+1.06000e-04'
+ mcm4l1p1_ca_w_0_170_s_1_980 = '-1.75938e-06*ic_cap*ic_cap+-8.62500e-07*ic_cap+1.06000e-04'
+ mcm4l1p1_ca_w_0_170_s_4_500 = '-1.75938e-06*ic_cap*ic_cap+-8.62500e-07*ic_cap+1.06000e-04'
+ mcm4l1p1_ca_w_1_360_s_0_180 = '-1.75938e-06*ic_cap*ic_cap+-8.62500e-07*ic_cap+1.06000e-04'
+ mcm4l1p1_ca_w_1_360_s_0_225 = '-1.75938e-06*ic_cap*ic_cap+-8.62500e-07*ic_cap+1.06000e-04'
+ mcm4l1p1_ca_w_1_360_s_0_270 = '-1.75938e-06*ic_cap*ic_cap+-8.62500e-07*ic_cap+1.06000e-04'
+ mcm4l1p1_ca_w_1_360_s_0_360 = '-1.75938e-06*ic_cap*ic_cap+-8.62500e-07*ic_cap+1.06000e-04'
+ mcm4l1p1_ca_w_1_360_s_0_450 = '-1.75938e-06*ic_cap*ic_cap+-8.62500e-07*ic_cap+1.06000e-04'
+ mcm4l1p1_ca_w_1_360_s_0_540 = '-1.75938e-06*ic_cap*ic_cap+-8.62500e-07*ic_cap+1.06000e-04'
+ mcm4l1p1_ca_w_1_360_s_0_720 = '-1.75938e-06*ic_cap*ic_cap+-8.62500e-07*ic_cap+1.06000e-04'
+ mcm4l1p1_ca_w_1_360_s_1_080 = '-1.75938e-06*ic_cap*ic_cap+-8.62500e-07*ic_cap+1.06000e-04'
+ mcm4l1p1_ca_w_1_360_s_1_980 = '-1.75938e-06*ic_cap*ic_cap+-8.62500e-07*ic_cap+1.06000e-04'
+ mcm4l1p1_ca_w_1_360_s_4_500 = '-1.75938e-06*ic_cap*ic_cap+-8.62500e-07*ic_cap+1.06000e-04'
+ mcm4l1p1_cc_w_0_170_s_0_180 = '-6.71875e-13*ic_cap*ic_cap+-4.37500e-13*ic_cap+7.17000e-11'
+ mcm4l1p1_cc_w_0_170_s_0_225 = '-4.46875e-13*ic_cap*ic_cap+-3.12500e-13*ic_cap+5.95000e-11'
+ mcm4l1p1_cc_w_0_170_s_0_270 = '-3.03125e-13*ic_cap*ic_cap+-2.37500e-13*ic_cap+5.11000e-11'
+ mcm4l1p1_cc_w_0_170_s_0_360 = '-1.46875e-13*ic_cap*ic_cap+-1.37500e-13*ic_cap+3.92000e-11'
+ mcm4l1p1_cc_w_0_170_s_0_450 = '-5.62500e-14*ic_cap*ic_cap+-7.50000e-14*ic_cap+3.18000e-11'
+ mcm4l1p1_cc_w_0_170_s_0_540 = '-6.25000e-15*ic_cap*ic_cap+-5.00000e-14*ic_cap+2.59000e-11'
+ mcm4l1p1_cc_w_0_170_s_0_720 = '4.68750e-14*ic_cap*ic_cap+-1.25000e-14*ic_cap+1.83000e-11'
+ mcm4l1p1_cc_w_0_170_s_1_080 = '7.81250e-14*ic_cap*ic_cap+3.75000e-14*ic_cap+1.00000e-11'
+ mcm4l1p1_cc_w_0_170_s_1_980 = '5.53125e-14*ic_cap*ic_cap+2.87500e-14*ic_cap+2.96000e-12'
+ mcm4l1p1_cc_w_0_170_s_4_500 = '8.43750e-15*ic_cap*ic_cap+7.50000e-15*ic_cap+2.65000e-13'
+ mcm4l1p1_cc_w_1_360_s_0_180 = '-5.43750e-13*ic_cap*ic_cap+-3.50000e-13*ic_cap+8.41000e-11'
+ mcm4l1p1_cc_w_1_360_s_0_225 = '-3.31250e-13*ic_cap*ic_cap+-2.50000e-13*ic_cap+7.11000e-11'
+ mcm4l1p1_cc_w_1_360_s_0_270 = '-2.03125e-13*ic_cap*ic_cap+-1.62500e-13*ic_cap+6.17000e-11'
+ mcm4l1p1_cc_w_1_360_s_0_360 = '-5.62500e-14*ic_cap*ic_cap+-7.50000e-14*ic_cap+4.88000e-11'
+ mcm4l1p1_cc_w_1_360_s_0_450 = '2.18750e-14*ic_cap*ic_cap+-1.25000e-14*ic_cap+4.00000e-11'
+ mcm4l1p1_cc_w_1_360_s_0_540 = '6.56250e-14*ic_cap*ic_cap+1.25000e-14*ic_cap+3.37000e-11'
+ mcm4l1p1_cc_w_1_360_s_0_720 = '1.15625e-13*ic_cap*ic_cap+3.75000e-14*ic_cap+2.48000e-11'
+ mcm4l1p1_cc_w_1_360_s_1_080 = '1.31250e-13*ic_cap*ic_cap+7.50000e-14*ic_cap+1.48000e-11'
+ mcm4l1p1_cc_w_1_360_s_1_980 = '9.65625e-14*ic_cap*ic_cap+5.87500e-14*ic_cap+5.02000e-12'
+ mcm4l1p1_cc_w_1_360_s_4_500 = '2.00000e-14*ic_cap*ic_cap+1.25000e-14*ic_cap+4.55000e-13'
+ mcm4l1p1_cf_w_0_170_s_0_180 = '-8.34375e-14*ic_cap*ic_cap+-3.87500e-14*ic_cap+9.12000e-12'
+ mcm4l1p1_cf_w_0_170_s_0_225 = '-1.16563e-13*ic_cap*ic_cap+-5.62500e-14*ic_cap+1.12000e-11'
+ mcm4l1p1_cf_w_0_170_s_0_270 = '-1.50000e-13*ic_cap*ic_cap+-7.50000e-14*ic_cap+1.32000e-11'
+ mcm4l1p1_cf_w_0_170_s_0_360 = '-2.06250e-13*ic_cap*ic_cap+-1.00000e-13*ic_cap+1.72000e-11'
+ mcm4l1p1_cf_w_0_170_s_0_450 = '-2.56250e-13*ic_cap*ic_cap+-1.25000e-13*ic_cap+2.03000e-11'
+ mcm4l1p1_cf_w_0_170_s_0_540 = '-2.93750e-13*ic_cap*ic_cap+-1.50000e-13*ic_cap+2.35000e-11'
+ mcm4l1p1_cf_w_0_170_s_0_720 = '-3.40625e-13*ic_cap*ic_cap+-1.87500e-13*ic_cap+2.83000e-11'
+ mcm4l1p1_cf_w_0_170_s_1_080 = '-3.93750e-13*ic_cap*ic_cap+-2.25000e-13*ic_cap+3.48000e-11'
+ mcm4l1p1_cf_w_0_170_s_1_980 = '-3.75000e-13*ic_cap*ic_cap+-2.25000e-13*ic_cap+4.10000e-11'
+ mcm4l1p1_cf_w_0_170_s_4_500 = '-3.43750e-13*ic_cap*ic_cap+-2.00000e-13*ic_cap+4.37000e-11'
+ mcm4l1p1_cf_w_1_360_s_0_180 = '-8.34375e-14*ic_cap*ic_cap+-3.87500e-14*ic_cap+9.16000e-12'
+ mcm4l1p1_cf_w_1_360_s_0_225 = '-1.19063e-13*ic_cap*ic_cap+-5.62500e-14*ic_cap+1.13000e-11'
+ mcm4l1p1_cf_w_1_360_s_0_270 = '-1.50000e-13*ic_cap*ic_cap+-7.50000e-14*ic_cap+1.33000e-11'
+ mcm4l1p1_cf_w_1_360_s_0_360 = '-2.00000e-13*ic_cap*ic_cap+-1.00000e-13*ic_cap+1.70000e-11'
+ mcm4l1p1_cf_w_1_360_s_0_450 = '-2.50000e-13*ic_cap*ic_cap+-1.25000e-13*ic_cap+2.05000e-11'
+ mcm4l1p1_cf_w_1_360_s_0_540 = '-2.93750e-13*ic_cap*ic_cap+-1.50000e-13*ic_cap+2.36000e-11'
+ mcm4l1p1_cf_w_1_360_s_0_720 = '-3.40625e-13*ic_cap*ic_cap+-1.87500e-13*ic_cap+2.87000e-11'
+ mcm4l1p1_cf_w_1_360_s_1_080 = '-3.96875e-13*ic_cap*ic_cap+-2.12500e-13*ic_cap+3.61000e-11'
+ mcm4l1p1_cf_w_1_360_s_1_980 = '-3.87500e-13*ic_cap*ic_cap+-2.25000e-13*ic_cap+4.46000e-11'
+ mcm4l1p1_cf_w_1_360_s_4_500 = '-3.18750e-13*ic_cap*ic_cap+-1.75000e-13*ic_cap+4.90000e-11'
+ mcm4m1_ca_w_0_300_s_0_300 = '-1.25000e-07*ic_cap*ic_cap+-7.50000e-08*ic_cap+1.51000e-05'
+ mcm4m1_ca_w_0_300_s_0_360 = '-1.25000e-07*ic_cap*ic_cap+-7.50000e-08*ic_cap+1.51000e-05'
+ mcm4m1_ca_w_0_300_s_0_450 = '-1.25000e-07*ic_cap*ic_cap+-7.50000e-08*ic_cap+1.51000e-05'
+ mcm4m1_ca_w_0_300_s_0_600 = '-1.25000e-07*ic_cap*ic_cap+-7.50000e-08*ic_cap+1.51000e-05'
+ mcm4m1_ca_w_0_300_s_0_800 = '-1.25000e-07*ic_cap*ic_cap+-7.50000e-08*ic_cap+1.51000e-05'
+ mcm4m1_ca_w_0_300_s_1_000 = '-1.25000e-07*ic_cap*ic_cap+-7.50000e-08*ic_cap+1.51000e-05'
+ mcm4m1_ca_w_0_300_s_1_200 = '-1.25000e-07*ic_cap*ic_cap+-7.50000e-08*ic_cap+1.51000e-05'
+ mcm4m1_ca_w_0_300_s_2_100 = '-1.25000e-07*ic_cap*ic_cap+-7.50000e-08*ic_cap+1.51000e-05'
+ mcm4m1_ca_w_0_300_s_3_300 = '-1.25000e-07*ic_cap*ic_cap+-7.50000e-08*ic_cap+1.51000e-05'
+ mcm4m1_ca_w_0_300_s_9_000 = '-1.25000e-07*ic_cap*ic_cap+-7.50000e-08*ic_cap+1.51000e-05'
+ mcm4m1_ca_w_2_400_s_0_300 = '-1.25000e-07*ic_cap*ic_cap+-7.50000e-08*ic_cap+1.51000e-05'
+ mcm4m1_ca_w_2_400_s_0_360 = '-1.25000e-07*ic_cap*ic_cap+-7.50000e-08*ic_cap+1.51000e-05'
+ mcm4m1_ca_w_2_400_s_0_450 = '-1.25000e-07*ic_cap*ic_cap+-7.50000e-08*ic_cap+1.51000e-05'
+ mcm4m1_ca_w_2_400_s_0_600 = '-1.25000e-07*ic_cap*ic_cap+-7.50000e-08*ic_cap+1.51000e-05'
+ mcm4m1_ca_w_2_400_s_0_800 = '-1.25000e-07*ic_cap*ic_cap+-7.50000e-08*ic_cap+1.51000e-05'
+ mcm4m1_ca_w_2_400_s_1_000 = '-1.25000e-07*ic_cap*ic_cap+-7.50000e-08*ic_cap+1.51000e-05'
+ mcm4m1_ca_w_2_400_s_1_200 = '-1.25000e-07*ic_cap*ic_cap+-7.50000e-08*ic_cap+1.51000e-05'
+ mcm4m1_ca_w_2_400_s_2_100 = '-1.25000e-07*ic_cap*ic_cap+-7.50000e-08*ic_cap+1.51000e-05'
+ mcm4m1_ca_w_2_400_s_3_300 = '-1.25000e-07*ic_cap*ic_cap+-7.50000e-08*ic_cap+1.51000e-05'
+ mcm4m1_ca_w_2_400_s_9_000 = '-1.25000e-07*ic_cap*ic_cap+-7.50000e-08*ic_cap+1.51000e-05'
+ mcm4m1_cc_w_0_300_s_0_300 = '-7.90625e-13*ic_cap*ic_cap+-4.62500e-13*ic_cap+1.06000e-10'
+ mcm4m1_cc_w_0_300_s_0_360 = '-7.31250e-13*ic_cap*ic_cap+-4.00000e-13*ic_cap+9.94000e-11'
+ mcm4m1_cc_w_0_300_s_0_450 = '-6.12500e-13*ic_cap*ic_cap+-3.50000e-13*ic_cap+8.98000e-11'
+ mcm4m1_cc_w_0_300_s_0_600 = '-4.75000e-13*ic_cap*ic_cap+-3.00000e-13*ic_cap+7.73000e-11'
+ mcm4m1_cc_w_0_300_s_0_800 = '-3.40625e-13*ic_cap*ic_cap+-2.12500e-13*ic_cap+6.51000e-11'
+ mcm4m1_cc_w_0_300_s_1_000 = '-2.65625e-13*ic_cap*ic_cap+-1.62500e-13*ic_cap+5.61000e-11'
+ mcm4m1_cc_w_0_300_s_1_200 = '-2.06250e-13*ic_cap*ic_cap+-1.25000e-13*ic_cap+4.92000e-11'
+ mcm4m1_cc_w_0_300_s_2_100 = '-9.06250e-14*ic_cap*ic_cap+-6.25000e-14*ic_cap+3.18000e-11'
+ mcm4m1_cc_w_0_300_s_3_300 = '-3.12500e-14*ic_cap*ic_cap+-2.50000e-14*ic_cap+2.14000e-11'
+ mcm4m1_cc_w_0_300_s_9_000 = '6.56250e-15*ic_cap*ic_cap+8.75000e-15*ic_cap+5.86000e-12'
+ mcm4m1_cc_w_2_400_s_0_300 = '-8.43750e-13*ic_cap*ic_cap+-3.75000e-13*ic_cap+1.32000e-10'
+ mcm4m1_cc_w_2_400_s_0_360 = '-7.18750e-13*ic_cap*ic_cap+-3.75000e-13*ic_cap+1.23000e-10'
+ mcm4m1_cc_w_2_400_s_0_450 = '-5.93750e-13*ic_cap*ic_cap+-3.75000e-13*ic_cap+1.12000e-10'
+ mcm4m1_cc_w_2_400_s_0_600 = '-4.46875e-13*ic_cap*ic_cap+-2.62500e-13*ic_cap+9.70000e-11'
+ mcm4m1_cc_w_2_400_s_0_800 = '-3.06250e-13*ic_cap*ic_cap+-2.00000e-13*ic_cap+8.21000e-11'
+ mcm4m1_cc_w_2_400_s_1_000 = '-2.25000e-13*ic_cap*ic_cap+-1.50000e-13*ic_cap+7.12000e-11'
+ mcm4m1_cc_w_2_400_s_1_200 = '-1.75000e-13*ic_cap*ic_cap+-1.25000e-13*ic_cap+6.30000e-11'
+ mcm4m1_cc_w_2_400_s_2_100 = '-6.25000e-14*ic_cap*ic_cap+-5.00000e-14*ic_cap+4.21000e-11'
+ mcm4m1_cc_w_2_400_s_3_300 = '-9.37500e-15*ic_cap*ic_cap+-1.25000e-14*ic_cap+2.89000e-11'
+ mcm4m1_cc_w_2_400_s_9_000 = '1.93750e-14*ic_cap*ic_cap+1.75000e-14*ic_cap+9.10000e-12'
+ mcm4m1_cf_w_0_300_s_0_300 = '-2.81250e-15*ic_cap*ic_cap+-1.25000e-15*ic_cap+2.22000e-12'
+ mcm4m1_cf_w_0_300_s_0_360 = '-5.93750e-15*ic_cap*ic_cap+-3.75000e-15*ic_cap+2.65000e-12'
+ mcm4m1_cf_w_0_300_s_0_450 = '-1.12500e-14*ic_cap*ic_cap+-7.50000e-15*ic_cap+3.32000e-12'
+ mcm4m1_cf_w_0_300_s_0_600 = '-1.93750e-14*ic_cap*ic_cap+-1.25000e-14*ic_cap+4.40000e-12'
+ mcm4m1_cf_w_0_300_s_0_800 = '-3.09375e-14*ic_cap*ic_cap+-1.87500e-14*ic_cap+5.70000e-12'
+ mcm4m1_cf_w_0_300_s_1_000 = '-4.25000e-14*ic_cap*ic_cap+-2.50000e-14*ic_cap+7.02000e-12'
+ mcm4m1_cf_w_0_300_s_1_200 = '-5.25000e-14*ic_cap*ic_cap+-3.00000e-14*ic_cap+8.29000e-12'
+ mcm4m1_cf_w_0_300_s_2_100 = '-8.75000e-14*ic_cap*ic_cap+-5.00000e-14*ic_cap+1.37000e-11'
+ mcm4m1_cf_w_0_300_s_3_300 = '-1.25000e-13*ic_cap*ic_cap+-7.50000e-14*ic_cap+1.89000e-11'
+ mcm4m1_cf_w_0_300_s_9_000 = '-1.65625e-13*ic_cap*ic_cap+-1.12500e-13*ic_cap+3.09000e-11'
+ mcm4m1_cf_w_2_400_s_0_300 = '-2.81250e-15*ic_cap*ic_cap+-1.25000e-15*ic_cap+2.23000e-12'
+ mcm4m1_cf_w_2_400_s_0_360 = '-5.93750e-15*ic_cap*ic_cap+-3.75000e-15*ic_cap+2.66000e-12'
+ mcm4m1_cf_w_2_400_s_0_450 = '-1.15625e-14*ic_cap*ic_cap+-8.75000e-15*ic_cap+3.31000e-12'
+ mcm4m1_cf_w_2_400_s_0_600 = '-2.00000e-14*ic_cap*ic_cap+-1.25000e-14*ic_cap+4.36000e-12'
+ mcm4m1_cf_w_2_400_s_0_800 = '-3.12500e-14*ic_cap*ic_cap+-2.00000e-14*ic_cap+5.74000e-12'
+ mcm4m1_cf_w_2_400_s_1_000 = '-4.15625e-14*ic_cap*ic_cap+-2.62500e-14*ic_cap+7.07000e-12'
+ mcm4m1_cf_w_2_400_s_1_200 = '-5.12500e-14*ic_cap*ic_cap+-3.25000e-14*ic_cap+8.35000e-12'
+ mcm4m1_cf_w_2_400_s_2_100 = '-8.75000e-14*ic_cap*ic_cap+-5.00000e-14*ic_cap+1.36000e-11'
+ mcm4m1_cf_w_2_400_s_3_300 = '-1.25000e-13*ic_cap*ic_cap+-7.50000e-14*ic_cap+1.95000e-11'
+ mcm4m1_cf_w_2_400_s_9_000 = '-1.65625e-13*ic_cap*ic_cap+-1.12500e-13*ic_cap+3.39000e-11'
+ mcm4m1d_ca_w_0_140_s_0_140 = '-5.00000e-07*ic_cap*ic_cap+-3.25000e-07*ic_cap+4.87000e-05'
+ mcm4m1d_ca_w_0_140_s_0_175 = '-5.00000e-07*ic_cap*ic_cap+-3.25000e-07*ic_cap+4.87000e-05'
+ mcm4m1d_ca_w_0_140_s_0_210 = '-5.00000e-07*ic_cap*ic_cap+-3.25000e-07*ic_cap+4.87000e-05'
+ mcm4m1d_ca_w_0_140_s_0_280 = '-5.00000e-07*ic_cap*ic_cap+-3.25000e-07*ic_cap+4.87000e-05'
+ mcm4m1d_ca_w_0_140_s_0_350 = '-5.00000e-07*ic_cap*ic_cap+-3.25000e-07*ic_cap+4.87000e-05'
+ mcm4m1d_ca_w_0_140_s_0_420 = '-5.00000e-07*ic_cap*ic_cap+-3.25000e-07*ic_cap+4.87000e-05'
+ mcm4m1d_ca_w_0_140_s_0_560 = '-5.00000e-07*ic_cap*ic_cap+-3.25000e-07*ic_cap+4.87000e-05'
+ mcm4m1d_ca_w_0_140_s_0_840 = '-5.00000e-07*ic_cap*ic_cap+-3.25000e-07*ic_cap+4.87000e-05'
+ mcm4m1d_ca_w_0_140_s_1_540 = '-5.00000e-07*ic_cap*ic_cap+-3.25000e-07*ic_cap+4.87000e-05'
+ mcm4m1d_ca_w_0_140_s_3_500 = '-5.00000e-07*ic_cap*ic_cap+-3.25000e-07*ic_cap+4.87000e-05'
+ mcm4m1d_ca_w_1_120_s_0_140 = '-5.00000e-07*ic_cap*ic_cap+-3.25000e-07*ic_cap+4.87000e-05'
+ mcm4m1d_ca_w_1_120_s_0_175 = '-5.00000e-07*ic_cap*ic_cap+-3.25000e-07*ic_cap+4.87000e-05'
+ mcm4m1d_ca_w_1_120_s_0_210 = '-5.00000e-07*ic_cap*ic_cap+-3.25000e-07*ic_cap+4.87000e-05'
+ mcm4m1d_ca_w_1_120_s_0_280 = '-5.00000e-07*ic_cap*ic_cap+-3.25000e-07*ic_cap+4.87000e-05'
+ mcm4m1d_ca_w_1_120_s_0_350 = '-5.00000e-07*ic_cap*ic_cap+-3.25000e-07*ic_cap+4.87000e-05'
+ mcm4m1d_ca_w_1_120_s_0_420 = '-5.00000e-07*ic_cap*ic_cap+-3.25000e-07*ic_cap+4.87000e-05'
+ mcm4m1d_ca_w_1_120_s_0_560 = '-5.00000e-07*ic_cap*ic_cap+-3.25000e-07*ic_cap+4.87000e-05'
+ mcm4m1d_ca_w_1_120_s_0_840 = '-5.00000e-07*ic_cap*ic_cap+-3.25000e-07*ic_cap+4.87000e-05'
+ mcm4m1d_ca_w_1_120_s_1_540 = '-5.00000e-07*ic_cap*ic_cap+-3.25000e-07*ic_cap+4.87000e-05'
+ mcm4m1d_ca_w_1_120_s_3_500 = '-5.00000e-07*ic_cap*ic_cap+-3.25000e-07*ic_cap+4.87000e-05'
+ mcm4m1d_cc_w_0_140_s_0_140 = '-9.46875e-13*ic_cap*ic_cap+-5.12500e-13*ic_cap+1.03000e-10'
+ mcm4m1d_cc_w_0_140_s_0_175 = '-8.18750e-13*ic_cap*ic_cap+-5.75000e-13*ic_cap+1.00000e-10'
+ mcm4m1d_cc_w_0_140_s_0_210 = '-7.65625e-13*ic_cap*ic_cap+-4.12500e-13*ic_cap+9.52000e-11'
+ mcm4m1d_cc_w_0_140_s_0_280 = '-5.53125e-13*ic_cap*ic_cap+-3.87500e-13*ic_cap+8.35000e-11'
+ mcm4m1d_cc_w_0_140_s_0_350 = '-4.37500e-13*ic_cap*ic_cap+-3.00000e-13*ic_cap+7.19000e-11'
+ mcm4m1d_cc_w_0_140_s_0_420 = '-3.21875e-13*ic_cap*ic_cap+-1.87500e-13*ic_cap+6.21000e-11'
+ mcm4m1d_cc_w_0_140_s_0_560 = '-1.53125e-13*ic_cap*ic_cap+-1.37500e-13*ic_cap+4.83000e-11'
+ mcm4m1d_cc_w_0_140_s_0_840 = '-3.75000e-14*ic_cap*ic_cap+-2.50000e-14*ic_cap+3.29000e-11'
+ mcm4m1d_cc_w_0_140_s_1_540 = '5.31250e-14*ic_cap*ic_cap+3.75000e-14*ic_cap+1.53000e-11'
+ mcm4m1d_cc_w_0_140_s_3_500 = '4.53125e-14*ic_cap*ic_cap+3.37500e-14*ic_cap+2.56000e-12'
+ mcm4m1d_cc_w_1_120_s_0_140 = '-7.50000e-13*ic_cap*ic_cap+-5.00000e-13*ic_cap+1.20000e-10'
+ mcm4m1d_cc_w_1_120_s_0_175 = '-7.50000e-13*ic_cap*ic_cap+-2.50000e-13*ic_cap+1.17000e-10'
+ mcm4m1d_cc_w_1_120_s_0_210 = '-5.90625e-13*ic_cap*ic_cap+-3.62500e-13*ic_cap+1.10000e-10'
+ mcm4m1d_cc_w_1_120_s_0_280 = '-4.15625e-13*ic_cap*ic_cap+-2.62500e-13*ic_cap+9.59000e-11'
+ mcm4m1d_cc_w_1_120_s_0_350 = '-3.18750e-13*ic_cap*ic_cap+-1.75000e-13*ic_cap+8.32000e-11'
+ mcm4m1d_cc_w_1_120_s_0_420 = '-1.87500e-13*ic_cap*ic_cap+-1.50000e-13*ic_cap+7.20000e-11'
+ mcm4m1d_cc_w_1_120_s_0_560 = '-9.06250e-14*ic_cap*ic_cap+-3.75000e-14*ic_cap+5.66000e-11'
+ mcm4m1d_cc_w_1_120_s_0_840 = '3.12500e-14*ic_cap*ic_cap+2.50000e-14*ic_cap+3.84000e-11'
+ mcm4m1d_cc_w_1_120_s_1_540 = '1.03125e-13*ic_cap*ic_cap+6.25000e-14*ic_cap+1.83000e-11'
+ mcm4m1d_cc_w_1_120_s_3_500 = '6.75000e-14*ic_cap*ic_cap+5.00000e-14*ic_cap+3.17000e-12'
+ mcm4m1d_cf_w_0_140_s_0_140 = '-2.18750e-15*ic_cap*ic_cap+-3.75000e-15*ic_cap+3.37000e-12'
+ mcm4m1d_cf_w_0_140_s_0_175 = '-1.09375e-14*ic_cap*ic_cap+-8.75000e-15*ic_cap+4.21000e-12'
+ mcm4m1d_cf_w_0_140_s_0_210 = '-1.87500e-14*ic_cap*ic_cap+-1.25000e-14*ic_cap+5.06000e-12'
+ mcm4m1d_cf_w_0_140_s_0_280 = '-3.62500e-14*ic_cap*ic_cap+-2.50000e-14*ic_cap+6.70000e-12'
+ mcm4m1d_cf_w_0_140_s_0_350 = '-5.34375e-14*ic_cap*ic_cap+-3.62500e-14*ic_cap+8.31000e-12'
+ mcm4m1d_cf_w_0_140_s_0_420 = '-7.00000e-14*ic_cap*ic_cap+-4.50000e-14*ic_cap+9.94000e-12'
+ mcm4m1d_cf_w_0_140_s_0_560 = '-9.68750e-14*ic_cap*ic_cap+-6.25000e-14*ic_cap+1.29000e-11'
+ mcm4m1d_cf_w_0_140_s_0_840 = '-1.50000e-13*ic_cap*ic_cap+-1.00000e-13*ic_cap+1.83000e-11'
+ mcm4m1d_cf_w_0_140_s_1_540 = '-2.25000e-13*ic_cap*ic_cap+-1.50000e-13*ic_cap+2.83000e-11'
+ mcm4m1d_cf_w_0_140_s_3_500 = '-2.40625e-13*ic_cap*ic_cap+-1.62500e-13*ic_cap+3.90000e-11'
+ mcm4m1d_cf_w_1_120_s_0_140 = '-3.43750e-15*ic_cap*ic_cap+-1.25000e-15*ic_cap+3.44000e-12'
+ mcm4m1d_cf_w_1_120_s_0_175 = '-1.18750e-14*ic_cap*ic_cap+-7.50000e-15*ic_cap+4.28000e-12'
+ mcm4m1d_cf_w_1_120_s_0_210 = '-2.12500e-14*ic_cap*ic_cap+-1.50000e-14*ic_cap+5.12000e-12'
+ mcm4m1d_cf_w_1_120_s_0_280 = '-3.78125e-14*ic_cap*ic_cap+-2.62500e-14*ic_cap+6.77000e-12'
+ mcm4m1d_cf_w_1_120_s_0_350 = '-5.40625e-14*ic_cap*ic_cap+-3.62500e-14*ic_cap+8.39000e-12'
+ mcm4m1d_cf_w_1_120_s_0_420 = '-7.03125e-14*ic_cap*ic_cap+-4.62500e-14*ic_cap+9.98000e-12'
+ mcm4m1d_cf_w_1_120_s_0_560 = '-9.68750e-14*ic_cap*ic_cap+-6.25000e-14*ic_cap+1.30000e-11'
+ mcm4m1d_cf_w_1_120_s_0_840 = '-1.53125e-13*ic_cap*ic_cap+-8.75000e-14*ic_cap+1.86000e-11'
+ mcm4m1d_cf_w_1_120_s_1_540 = '-2.28125e-13*ic_cap*ic_cap+-1.37500e-13*ic_cap+2.92000e-11'
+ mcm4m1d_cf_w_1_120_s_3_500 = '-2.28125e-13*ic_cap*ic_cap+-1.62500e-13*ic_cap+4.14000e-11'
+ mcm4m1f_ca_w_0_140_s_0_140 = '-4.28125e-07*ic_cap*ic_cap+-2.62500e-07*ic_cap+4.09000e-05'
+ mcm4m1f_ca_w_0_140_s_0_175 = '-4.28125e-07*ic_cap*ic_cap+-2.62500e-07*ic_cap+4.09000e-05'
+ mcm4m1f_ca_w_0_140_s_0_210 = '-4.28125e-07*ic_cap*ic_cap+-2.62500e-07*ic_cap+4.09000e-05'
+ mcm4m1f_ca_w_0_140_s_0_280 = '-4.28125e-07*ic_cap*ic_cap+-2.62500e-07*ic_cap+4.09000e-05'
+ mcm4m1f_ca_w_0_140_s_0_350 = '-4.28125e-07*ic_cap*ic_cap+-2.62500e-07*ic_cap+4.09000e-05'
+ mcm4m1f_ca_w_0_140_s_0_420 = '-4.28125e-07*ic_cap*ic_cap+-2.62500e-07*ic_cap+4.09000e-05'
+ mcm4m1f_ca_w_0_140_s_0_560 = '-4.28125e-07*ic_cap*ic_cap+-2.62500e-07*ic_cap+4.09000e-05'
+ mcm4m1f_ca_w_0_140_s_0_840 = '-4.28125e-07*ic_cap*ic_cap+-2.62500e-07*ic_cap+4.09000e-05'
+ mcm4m1f_ca_w_0_140_s_1_540 = '-4.28125e-07*ic_cap*ic_cap+-2.62500e-07*ic_cap+4.09000e-05'
+ mcm4m1f_ca_w_0_140_s_3_500 = '-4.28125e-07*ic_cap*ic_cap+-2.62500e-07*ic_cap+4.09000e-05'
+ mcm4m1f_ca_w_1_120_s_0_140 = '-4.28125e-07*ic_cap*ic_cap+-2.62500e-07*ic_cap+4.09000e-05'
+ mcm4m1f_ca_w_1_120_s_0_175 = '-4.28125e-07*ic_cap*ic_cap+-2.62500e-07*ic_cap+4.09000e-05'
+ mcm4m1f_ca_w_1_120_s_0_210 = '-4.28125e-07*ic_cap*ic_cap+-2.62500e-07*ic_cap+4.09000e-05'
+ mcm4m1f_ca_w_1_120_s_0_280 = '-4.28125e-07*ic_cap*ic_cap+-2.62500e-07*ic_cap+4.09000e-05'
+ mcm4m1f_ca_w_1_120_s_0_350 = '-4.28125e-07*ic_cap*ic_cap+-2.62500e-07*ic_cap+4.09000e-05'
+ mcm4m1f_ca_w_1_120_s_0_420 = '-4.28125e-07*ic_cap*ic_cap+-2.62500e-07*ic_cap+4.09000e-05'
+ mcm4m1f_ca_w_1_120_s_0_560 = '-4.28125e-07*ic_cap*ic_cap+-2.62500e-07*ic_cap+4.09000e-05'
+ mcm4m1f_ca_w_1_120_s_0_840 = '-4.28125e-07*ic_cap*ic_cap+-2.62500e-07*ic_cap+4.09000e-05'
+ mcm4m1f_ca_w_1_120_s_1_540 = '-4.28125e-07*ic_cap*ic_cap+-2.62500e-07*ic_cap+4.09000e-05'
+ mcm4m1f_ca_w_1_120_s_3_500 = '-4.28125e-07*ic_cap*ic_cap+-2.62500e-07*ic_cap+4.09000e-05'
+ mcm4m1f_cc_w_0_140_s_0_140 = '-9.62500e-13*ic_cap*ic_cap+-5.25000e-13*ic_cap+1.04000e-10'
+ mcm4m1f_cc_w_0_140_s_0_175 = '-8.93750e-13*ic_cap*ic_cap+-6.00000e-13*ic_cap+1.02000e-10'
+ mcm4m1f_cc_w_0_140_s_0_210 = '-7.78125e-13*ic_cap*ic_cap+-4.12500e-13*ic_cap+9.63000e-11'
+ mcm4m1f_cc_w_0_140_s_0_280 = '-5.62500e-13*ic_cap*ic_cap+-4.00000e-13*ic_cap+8.48000e-11'
+ mcm4m1f_cc_w_0_140_s_0_350 = '-4.40625e-13*ic_cap*ic_cap+-2.62500e-13*ic_cap+7.33000e-11'
+ mcm4m1f_cc_w_0_140_s_0_420 = '-3.34375e-13*ic_cap*ic_cap+-1.87500e-13*ic_cap+6.36000e-11'
+ mcm4m1f_cc_w_0_140_s_0_560 = '-1.78125e-13*ic_cap*ic_cap+-1.12500e-13*ic_cap+5.03000e-11'
+ mcm4m1f_cc_w_0_140_s_0_840 = '-5.00000e-14*ic_cap*ic_cap+-5.00000e-14*ic_cap+3.51000e-11'
+ mcm4m1f_cc_w_0_140_s_1_540 = '5.00000e-14*ic_cap*ic_cap+2.50000e-14*ic_cap+1.74000e-11'
+ mcm4m1f_cc_w_0_140_s_3_500 = '5.71875e-14*ic_cap*ic_cap+3.87500e-14*ic_cap+3.40000e-12'
+ mcm4m1f_cc_w_1_120_s_0_140 = '-7.50000e-13*ic_cap*ic_cap+-5.00000e-13*ic_cap+1.23000e-10'
+ mcm4m1f_cc_w_1_120_s_0_175 = '-7.81250e-13*ic_cap*ic_cap+-3.75000e-13*ic_cap+1.20000e-10'
+ mcm4m1f_cc_w_1_120_s_0_210 = '-5.93750e-13*ic_cap*ic_cap+-3.75000e-13*ic_cap+1.13000e-10'
+ mcm4m1f_cc_w_1_120_s_0_280 = '-4.31250e-13*ic_cap*ic_cap+-2.50000e-13*ic_cap+9.88000e-11'
+ mcm4m1f_cc_w_1_120_s_0_350 = '-3.21875e-13*ic_cap*ic_cap+-1.87500e-13*ic_cap+8.60000e-11'
+ mcm4m1f_cc_w_1_120_s_0_420 = '-2.18750e-13*ic_cap*ic_cap+-1.25000e-13*ic_cap+7.51000e-11'
+ mcm4m1f_cc_w_1_120_s_0_560 = '-7.81250e-14*ic_cap*ic_cap+-6.25000e-14*ic_cap+5.93000e-11'
+ mcm4m1f_cc_w_1_120_s_0_840 = '3.43750e-14*ic_cap*ic_cap+1.25000e-14*ic_cap+4.12000e-11'
+ mcm4m1f_cc_w_1_120_s_1_540 = '1.18750e-13*ic_cap*ic_cap+7.50000e-14*ic_cap+2.07000e-11'
+ mcm4m1f_cc_w_1_120_s_3_500 = '8.37500e-14*ic_cap*ic_cap+5.75000e-14*ic_cap+4.21000e-12'
+ mcm4m1f_cf_w_0_140_s_0_140 = '-2.81250e-15*ic_cap*ic_cap+-3.75000e-15*ic_cap+2.84000e-12'
+ mcm4m1f_cf_w_0_140_s_0_175 = '-1.00000e-14*ic_cap*ic_cap+-7.50000e-15*ic_cap+3.54000e-12'
+ mcm4m1f_cf_w_0_140_s_0_210 = '-1.59375e-14*ic_cap*ic_cap+-1.12500e-14*ic_cap+4.25000e-12'
+ mcm4m1f_cf_w_0_140_s_0_280 = '-3.18750e-14*ic_cap*ic_cap+-2.00000e-14*ic_cap+5.64000e-12'
+ mcm4m1f_cf_w_0_140_s_0_350 = '-4.65625e-14*ic_cap*ic_cap+-2.87500e-14*ic_cap+7.00000e-12'
+ mcm4m1f_cf_w_0_140_s_0_420 = '-6.09375e-14*ic_cap*ic_cap+-3.87500e-14*ic_cap+8.39000e-12'
+ mcm4m1f_cf_w_0_140_s_0_560 = '-8.90625e-14*ic_cap*ic_cap+-5.37500e-14*ic_cap+1.10000e-11'
+ mcm4m1f_cf_w_0_140_s_0_840 = '-1.34375e-13*ic_cap*ic_cap+-8.75000e-14*ic_cap+1.57000e-11'
+ mcm4m1f_cf_w_0_140_s_1_540 = '-2.09375e-13*ic_cap*ic_cap+-1.37500e-13*ic_cap+2.48000e-11'
+ mcm4m1f_cf_w_0_140_s_3_500 = '-2.43750e-13*ic_cap*ic_cap+-1.50000e-13*ic_cap+3.59000e-11'
+ mcm4m1f_cf_w_1_120_s_0_140 = '-3.43750e-15*ic_cap*ic_cap+-3.75000e-15*ic_cap+2.88000e-12'
+ mcm4m1f_cf_w_1_120_s_0_175 = '-1.00000e-14*ic_cap*ic_cap+-7.50000e-15*ic_cap+3.58000e-12'
+ mcm4m1f_cf_w_1_120_s_0_210 = '-1.84375e-14*ic_cap*ic_cap+-1.12500e-14*ic_cap+4.29000e-12'
+ mcm4m1f_cf_w_1_120_s_0_280 = '-3.21875e-14*ic_cap*ic_cap+-2.12500e-14*ic_cap+5.68000e-12'
+ mcm4m1f_cf_w_1_120_s_0_350 = '-4.65625e-14*ic_cap*ic_cap+-2.87500e-14*ic_cap+7.06000e-12'
+ mcm4m1f_cf_w_1_120_s_0_420 = '-5.96875e-14*ic_cap*ic_cap+-4.12500e-14*ic_cap+8.40000e-12'
+ mcm4m1f_cf_w_1_120_s_0_560 = '-8.68750e-14*ic_cap*ic_cap+-5.25000e-14*ic_cap+1.10000e-11'
+ mcm4m1f_cf_w_1_120_s_0_840 = '-1.37500e-13*ic_cap*ic_cap+-7.50000e-14*ic_cap+1.59000e-11'
+ mcm4m1f_cf_w_1_120_s_1_540 = '-2.15625e-13*ic_cap*ic_cap+-1.37500e-13*ic_cap+2.56000e-11'
+ mcm4m1f_cf_w_1_120_s_3_500 = '-2.28125e-13*ic_cap*ic_cap+-1.62500e-13*ic_cap+3.82000e-11'
+ mcm4m1l1_ca_w_0_140_s_0_140 = '-2.09375e-06*ic_cap*ic_cap+-1.37500e-06*ic_cap+1.29000e-04'
+ mcm4m1l1_ca_w_0_140_s_0_175 = '-2.09375e-06*ic_cap*ic_cap+-1.37500e-06*ic_cap+1.29000e-04'
+ mcm4m1l1_ca_w_0_140_s_0_210 = '-2.09375e-06*ic_cap*ic_cap+-1.37500e-06*ic_cap+1.29000e-04'
+ mcm4m1l1_ca_w_0_140_s_0_280 = '-2.09375e-06*ic_cap*ic_cap+-1.37500e-06*ic_cap+1.29000e-04'
+ mcm4m1l1_ca_w_0_140_s_0_350 = '-2.09375e-06*ic_cap*ic_cap+-1.37500e-06*ic_cap+1.29000e-04'
+ mcm4m1l1_ca_w_0_140_s_0_420 = '-2.09375e-06*ic_cap*ic_cap+-1.37500e-06*ic_cap+1.29000e-04'
+ mcm4m1l1_ca_w_0_140_s_0_560 = '-2.09375e-06*ic_cap*ic_cap+-1.37500e-06*ic_cap+1.29000e-04'
+ mcm4m1l1_ca_w_0_140_s_0_840 = '-2.09375e-06*ic_cap*ic_cap+-1.37500e-06*ic_cap+1.29000e-04'
+ mcm4m1l1_ca_w_0_140_s_1_540 = '-2.09375e-06*ic_cap*ic_cap+-1.37500e-06*ic_cap+1.29000e-04'
+ mcm4m1l1_ca_w_0_140_s_3_500 = '-2.09375e-06*ic_cap*ic_cap+-1.37500e-06*ic_cap+1.29000e-04'
+ mcm4m1l1_ca_w_1_120_s_0_140 = '-2.09375e-06*ic_cap*ic_cap+-1.37500e-06*ic_cap+1.29000e-04'
+ mcm4m1l1_ca_w_1_120_s_0_175 = '-2.09375e-06*ic_cap*ic_cap+-1.37500e-06*ic_cap+1.29000e-04'
+ mcm4m1l1_ca_w_1_120_s_0_210 = '-2.09375e-06*ic_cap*ic_cap+-1.37500e-06*ic_cap+1.29000e-04'
+ mcm4m1l1_ca_w_1_120_s_0_280 = '-2.09375e-06*ic_cap*ic_cap+-1.37500e-06*ic_cap+1.29000e-04'
+ mcm4m1l1_ca_w_1_120_s_0_350 = '-2.09375e-06*ic_cap*ic_cap+-1.37500e-06*ic_cap+1.29000e-04'
+ mcm4m1l1_ca_w_1_120_s_0_420 = '-2.09375e-06*ic_cap*ic_cap+-1.37500e-06*ic_cap+1.29000e-04'
+ mcm4m1l1_ca_w_1_120_s_0_560 = '-2.09375e-06*ic_cap*ic_cap+-1.37500e-06*ic_cap+1.29000e-04'
+ mcm4m1l1_ca_w_1_120_s_0_840 = '-2.09375e-06*ic_cap*ic_cap+-1.37500e-06*ic_cap+1.29000e-04'
+ mcm4m1l1_ca_w_1_120_s_1_540 = '-2.09375e-06*ic_cap*ic_cap+-1.37500e-06*ic_cap+1.29000e-04'
+ mcm4m1l1_ca_w_1_120_s_3_500 = '-2.09375e-06*ic_cap*ic_cap+-1.37500e-06*ic_cap+1.29000e-04'
+ mcm4m1l1_cc_w_0_140_s_0_140 = '-7.93750e-13*ic_cap*ic_cap+-3.75000e-13*ic_cap+9.48000e-11'
+ mcm4m1l1_cc_w_0_140_s_0_175 = '-7.56250e-13*ic_cap*ic_cap+-3.25000e-13*ic_cap+9.24000e-11'
+ mcm4m1l1_cc_w_0_140_s_0_210 = '-6.03125e-13*ic_cap*ic_cap+-3.12500e-13*ic_cap+8.59000e-11'
+ mcm4m1l1_cc_w_0_140_s_0_280 = '-4.06250e-13*ic_cap*ic_cap+-2.50000e-13*ic_cap+7.35000e-11'
+ mcm4m1l1_cc_w_0_140_s_0_350 = '-3.00000e-13*ic_cap*ic_cap+-2.25000e-13*ic_cap+6.15000e-11'
+ mcm4m1l1_cc_w_0_140_s_0_420 = '-1.65625e-13*ic_cap*ic_cap+-1.37500e-13*ic_cap+5.10000e-11'
+ mcm4m1l1_cc_w_0_140_s_0_560 = '-4.06250e-14*ic_cap*ic_cap+-1.25000e-14*ic_cap+3.72000e-11'
+ mcm4m1l1_cc_w_0_140_s_0_840 = '5.00000e-14*ic_cap*ic_cap+5.00000e-14*ic_cap+2.20000e-11'
+ mcm4m1l1_cc_w_0_140_s_1_540 = '7.21875e-14*ic_cap*ic_cap+5.87500e-14*ic_cap+7.54000e-12'
+ mcm4m1l1_cc_w_0_140_s_3_500 = '1.92187e-14*ic_cap*ic_cap+1.81250e-14*ic_cap+7.50000e-13'
+ mcm4m1l1_cc_w_1_120_s_0_140 = '-6.18750e-13*ic_cap*ic_cap+-2.75000e-13*ic_cap+1.06000e-10'
+ mcm4m1l1_cc_w_1_120_s_0_175 = '-6.31250e-13*ic_cap*ic_cap+-2.00000e-13*ic_cap+1.03000e-10'
+ mcm4m1l1_cc_w_1_120_s_0_210 = '-4.81250e-13*ic_cap*ic_cap+-2.50000e-13*ic_cap+9.61000e-11'
+ mcm4m1l1_cc_w_1_120_s_0_280 = '-3.03125e-13*ic_cap*ic_cap+-1.37500e-13*ic_cap+8.18000e-11'
+ mcm4m1l1_cc_w_1_120_s_0_350 = '-2.09375e-13*ic_cap*ic_cap+-8.75000e-14*ic_cap+6.92000e-11'
+ mcm4m1l1_cc_w_1_120_s_0_420 = '-9.06250e-14*ic_cap*ic_cap+-6.25000e-14*ic_cap+5.81000e-11'
+ mcm4m1l1_cc_w_1_120_s_0_560 = '1.25000e-14*ic_cap*ic_cap+2.50000e-14*ic_cap+4.30000e-11'
+ mcm4m1l1_cc_w_1_120_s_0_840 = '1.00000e-13*ic_cap*ic_cap+1.00000e-13*ic_cap+2.62000e-11'
+ mcm4m1l1_cc_w_1_120_s_1_540 = '1.02500e-13*ic_cap*ic_cap+8.75000e-14*ic_cap+9.81000e-12'
+ mcm4m1l1_cc_w_1_120_s_3_500 = '3.34375e-14*ic_cap*ic_cap+3.12500e-14*ic_cap+1.05000e-12'
+ mcm4m1l1_cf_w_0_140_s_0_140 = '-6.12500e-14*ic_cap*ic_cap+-5.00000e-14*ic_cap+8.49000e-12'
+ mcm4m1l1_cf_w_0_140_s_0_175 = '-9.62500e-14*ic_cap*ic_cap+-7.00000e-14*ic_cap+1.07000e-11'
+ mcm4m1l1_cf_w_0_140_s_0_210 = '-1.31250e-13*ic_cap*ic_cap+-1.00000e-13*ic_cap+1.29000e-11'
+ mcm4m1l1_cf_w_0_140_s_0_280 = '-1.90625e-13*ic_cap*ic_cap+-1.37500e-13*ic_cap+1.69000e-11'
+ mcm4m1l1_cf_w_0_140_s_0_350 = '-2.50000e-13*ic_cap*ic_cap+-1.75000e-13*ic_cap+2.07000e-11'
+ mcm4m1l1_cf_w_0_140_s_0_420 = '-2.96875e-13*ic_cap*ic_cap+-2.12500e-13*ic_cap+2.42000e-11'
+ mcm4m1l1_cf_w_0_140_s_0_560 = '-3.75000e-13*ic_cap*ic_cap+-2.50000e-13*ic_cap+3.04000e-11'
+ mcm4m1l1_cf_w_0_140_s_0_840 = '-4.68750e-13*ic_cap*ic_cap+-3.25000e-13*ic_cap+3.97000e-11'
+ mcm4m1l1_cf_w_0_140_s_1_540 = '-5.25000e-13*ic_cap*ic_cap+-3.75000e-13*ic_cap+5.16000e-11'
+ mcm4m1l1_cf_w_0_140_s_3_500 = '-4.93750e-13*ic_cap*ic_cap+-3.25000e-13*ic_cap+5.84000e-11'
+ mcm4m1l1_cf_w_1_120_s_0_140 = '-6.40625e-14*ic_cap*ic_cap+-5.12500e-14*ic_cap+8.63000e-12'
+ mcm4m1l1_cf_w_1_120_s_0_175 = '-9.59375e-14*ic_cap*ic_cap+-7.37500e-14*ic_cap+1.08000e-11'
+ mcm4m1l1_cf_w_1_120_s_0_210 = '-1.34375e-13*ic_cap*ic_cap+-8.75000e-14*ic_cap+1.30000e-11'
+ mcm4m1l1_cf_w_1_120_s_0_280 = '-1.90625e-13*ic_cap*ic_cap+-1.37500e-13*ic_cap+1.70000e-11'
+ mcm4m1l1_cf_w_1_120_s_0_350 = '-2.50000e-13*ic_cap*ic_cap+-1.75000e-13*ic_cap+2.08000e-11'
+ mcm4m1l1_cf_w_1_120_s_0_420 = '-2.93750e-13*ic_cap*ic_cap+-2.00000e-13*ic_cap+2.43000e-11'
+ mcm4m1l1_cf_w_1_120_s_0_560 = '-3.78125e-13*ic_cap*ic_cap+-2.62500e-13*ic_cap+3.05000e-11'
+ mcm4m1l1_cf_w_1_120_s_0_840 = '-4.75000e-13*ic_cap*ic_cap+-3.25000e-13*ic_cap+4.01000e-11'
+ mcm4m1l1_cf_w_1_120_s_1_540 = '-5.31250e-13*ic_cap*ic_cap+-3.75000e-13*ic_cap+5.30000e-11'
+ mcm4m1l1_cf_w_1_120_s_3_500 = '-4.71875e-13*ic_cap*ic_cap+-3.37500e-13*ic_cap+6.13000e-11'
+ mcm4m1p1_ca_w_0_140_s_0_140 = '-8.09375e-07*ic_cap*ic_cap+-4.87500e-07*ic_cap+6.00000e-05'
+ mcm4m1p1_ca_w_0_140_s_0_175 = '-8.09375e-07*ic_cap*ic_cap+-4.87500e-07*ic_cap+6.00000e-05'
+ mcm4m1p1_ca_w_0_140_s_0_210 = '-8.09375e-07*ic_cap*ic_cap+-4.87500e-07*ic_cap+6.00000e-05'
+ mcm4m1p1_ca_w_0_140_s_0_280 = '-8.09375e-07*ic_cap*ic_cap+-4.87500e-07*ic_cap+6.00000e-05'
+ mcm4m1p1_ca_w_0_140_s_0_350 = '-8.09375e-07*ic_cap*ic_cap+-4.87500e-07*ic_cap+6.00000e-05'
+ mcm4m1p1_ca_w_0_140_s_0_420 = '-8.09375e-07*ic_cap*ic_cap+-4.87500e-07*ic_cap+6.00000e-05'
+ mcm4m1p1_ca_w_0_140_s_0_560 = '-8.09375e-07*ic_cap*ic_cap+-4.87500e-07*ic_cap+6.00000e-05'
+ mcm4m1p1_ca_w_0_140_s_0_840 = '-8.09375e-07*ic_cap*ic_cap+-4.87500e-07*ic_cap+6.00000e-05'
+ mcm4m1p1_ca_w_0_140_s_1_540 = '-8.09375e-07*ic_cap*ic_cap+-4.87500e-07*ic_cap+6.00000e-05'
+ mcm4m1p1_ca_w_0_140_s_3_500 = '-8.09375e-07*ic_cap*ic_cap+-4.87500e-07*ic_cap+6.00000e-05'
+ mcm4m1p1_ca_w_1_120_s_0_140 = '-8.09375e-07*ic_cap*ic_cap+-4.87500e-07*ic_cap+6.00000e-05'
+ mcm4m1p1_ca_w_1_120_s_0_175 = '-8.09375e-07*ic_cap*ic_cap+-4.87500e-07*ic_cap+6.00000e-05'
+ mcm4m1p1_ca_w_1_120_s_0_210 = '-8.09375e-07*ic_cap*ic_cap+-4.87500e-07*ic_cap+6.00000e-05'
+ mcm4m1p1_ca_w_1_120_s_0_280 = '-8.09375e-07*ic_cap*ic_cap+-4.87500e-07*ic_cap+6.00000e-05'
+ mcm4m1p1_ca_w_1_120_s_0_350 = '-8.09375e-07*ic_cap*ic_cap+-4.87500e-07*ic_cap+6.00000e-05'
+ mcm4m1p1_ca_w_1_120_s_0_420 = '-8.09375e-07*ic_cap*ic_cap+-4.87500e-07*ic_cap+6.00000e-05'
+ mcm4m1p1_ca_w_1_120_s_0_560 = '-8.09375e-07*ic_cap*ic_cap+-4.87500e-07*ic_cap+6.00000e-05'
+ mcm4m1p1_ca_w_1_120_s_0_840 = '-8.09375e-07*ic_cap*ic_cap+-4.87500e-07*ic_cap+6.00000e-05'
+ mcm4m1p1_ca_w_1_120_s_1_540 = '-8.09375e-07*ic_cap*ic_cap+-4.87500e-07*ic_cap+6.00000e-05'
+ mcm4m1p1_ca_w_1_120_s_3_500 = '-8.09375e-07*ic_cap*ic_cap+-4.87500e-07*ic_cap+6.00000e-05'
+ mcm4m1p1_cc_w_0_140_s_0_140 = '-9.21875e-13*ic_cap*ic_cap+-4.87500e-13*ic_cap+1.02000e-10'
+ mcm4m1p1_cc_w_0_140_s_0_175 = '-8.09375e-13*ic_cap*ic_cap+-5.62500e-13*ic_cap+9.91000e-11'
+ mcm4m1p1_cc_w_0_140_s_0_210 = '-6.96875e-13*ic_cap*ic_cap+-3.62500e-13*ic_cap+9.32000e-11'
+ mcm4m1p1_cc_w_0_140_s_0_280 = '-5.12500e-13*ic_cap*ic_cap+-3.25000e-13*ic_cap+8.17000e-11'
+ mcm4m1p1_cc_w_0_140_s_0_350 = '-3.53125e-13*ic_cap*ic_cap+-2.37500e-13*ic_cap+6.97000e-11'
+ mcm4m1p1_cc_w_0_140_s_0_420 = '-2.75000e-13*ic_cap*ic_cap+-1.75000e-13*ic_cap+6.00000e-11'
+ mcm4m1p1_cc_w_0_140_s_0_560 = '-1.15625e-13*ic_cap*ic_cap+-8.75000e-14*ic_cap+4.62000e-11'
+ mcm4m1p1_cc_w_0_140_s_0_840 = '1.87500e-14*ic_cap*ic_cap+3.03000e-11'
+ mcm4m1p1_cc_w_0_140_s_1_540 = '9.68750e-14*ic_cap*ic_cap+6.25000e-14*ic_cap+1.31000e-11'
+ mcm4m1p1_cc_w_0_140_s_3_500 = '4.90625e-14*ic_cap*ic_cap+3.62500e-14*ic_cap+1.84000e-12'
+ mcm4m1p1_cc_w_1_120_s_0_140 = '-7.18750e-13*ic_cap*ic_cap+-3.75000e-13*ic_cap+1.17000e-10'
+ mcm4m1p1_cc_w_1_120_s_0_175 = '-6.25000e-13*ic_cap*ic_cap+-2.50000e-13*ic_cap+1.13000e-10'
+ mcm4m1p1_cc_w_1_120_s_0_210 = '-5.43750e-13*ic_cap*ic_cap+-3.50000e-13*ic_cap+1.07000e-10'
+ mcm4m1p1_cc_w_1_120_s_0_280 = '-3.43750e-13*ic_cap*ic_cap+-2.25000e-13*ic_cap+9.24000e-11'
+ mcm4m1p1_cc_w_1_120_s_0_350 = '-2.37500e-13*ic_cap*ic_cap+-1.50000e-13*ic_cap+7.96000e-11'
+ mcm4m1p1_cc_w_1_120_s_0_420 = '-1.43750e-13*ic_cap*ic_cap+-1.00000e-13*ic_cap+6.88000e-11'
+ mcm4m1p1_cc_w_1_120_s_0_560 = '-3.12500e-15*ic_cap*ic_cap+-1.25000e-14*ic_cap+5.30000e-11'
+ mcm4m1p1_cc_w_1_120_s_0_840 = '9.37500e-14*ic_cap*ic_cap+5.00000e-14*ic_cap+3.52000e-11'
+ mcm4m1p1_cc_w_1_120_s_1_540 = '1.46875e-13*ic_cap*ic_cap+8.75000e-14*ic_cap+1.57000e-11'
+ mcm4m1p1_cc_w_1_120_s_3_500 = '6.93750e-14*ic_cap*ic_cap+4.75000e-14*ic_cap+2.33000e-12'
+ mcm4m1p1_cf_w_0_140_s_0_140 = '-1.90625e-14*ic_cap*ic_cap+-1.37500e-14*ic_cap+4.15000e-12'
+ mcm4m1p1_cf_w_0_140_s_0_175 = '-3.28125e-14*ic_cap*ic_cap+-2.12500e-14*ic_cap+5.18000e-12'
+ mcm4m1p1_cf_w_0_140_s_0_210 = '-4.59375e-14*ic_cap*ic_cap+-2.87500e-14*ic_cap+6.23000e-12'
+ mcm4m1p1_cf_w_0_140_s_0_280 = '-7.34375e-14*ic_cap*ic_cap+-4.37500e-14*ic_cap+8.23000e-12'
+ mcm4m1p1_cf_w_0_140_s_0_350 = '-9.96875e-14*ic_cap*ic_cap+-6.12500e-14*ic_cap+1.02000e-11'
+ mcm4m1p1_cf_w_0_140_s_0_420 = '-1.23750e-13*ic_cap*ic_cap+-7.00000e-14*ic_cap+1.21000e-11'
+ mcm4m1p1_cf_w_0_140_s_0_560 = '-1.68750e-13*ic_cap*ic_cap+-1.00000e-13*ic_cap+1.57000e-11'
+ mcm4m1p1_cf_w_0_140_s_0_840 = '-2.43750e-13*ic_cap*ic_cap+-1.50000e-13*ic_cap+2.20000e-11'
+ mcm4m1p1_cf_w_0_140_s_1_540 = '-3.28125e-13*ic_cap*ic_cap+-2.12500e-13*ic_cap+3.28000e-11'
+ mcm4m1p1_cf_w_0_140_s_3_500 = '-3.21875e-13*ic_cap*ic_cap+-2.12500e-13*ic_cap+4.27000e-11'
+ mcm4m1p1_cf_w_1_120_s_0_140 = '-2.28125e-14*ic_cap*ic_cap+-1.62500e-14*ic_cap+4.31000e-12'
+ mcm4m1p1_cf_w_1_120_s_0_175 = '-3.50000e-14*ic_cap*ic_cap+-2.25000e-14*ic_cap+5.32000e-12'
+ mcm4m1p1_cf_w_1_120_s_0_210 = '-4.90625e-14*ic_cap*ic_cap+-3.12500e-14*ic_cap+6.34000e-12'
+ mcm4m1p1_cf_w_1_120_s_0_280 = '-7.43750e-14*ic_cap*ic_cap+-4.75000e-14*ic_cap+8.35000e-12'
+ mcm4m1p1_cf_w_1_120_s_0_350 = '-9.93750e-14*ic_cap*ic_cap+-6.25000e-14*ic_cap+1.03000e-11'
+ mcm4m1p1_cf_w_1_120_s_0_420 = '-1.24375e-13*ic_cap*ic_cap+-7.25000e-14*ic_cap+1.22000e-11'
+ mcm4m1p1_cf_w_1_120_s_0_560 = '-1.71875e-13*ic_cap*ic_cap+-1.12500e-13*ic_cap+1.59000e-11'
+ mcm4m1p1_cf_w_1_120_s_0_840 = '-2.43750e-13*ic_cap*ic_cap+-1.50000e-13*ic_cap+2.23000e-11'
+ mcm4m1p1_cf_w_1_120_s_1_540 = '-3.34375e-13*ic_cap*ic_cap+-2.12500e-13*ic_cap+3.38000e-11'
+ mcm4m1p1_cf_w_1_120_s_3_500 = '-3.06250e-13*ic_cap*ic_cap+-2.00000e-13*ic_cap+4.52000e-11'
+ mcm4m2_ca_w_0_300_s_0_300 = '-1.68750e-07*ic_cap*ic_cap+-1.00000e-07*ic_cap+2.09000e-05'
+ mcm4m2_ca_w_0_300_s_0_360 = '-1.68750e-07*ic_cap*ic_cap+-1.00000e-07*ic_cap+2.09000e-05'
+ mcm4m2_ca_w_0_300_s_0_450 = '-1.68750e-07*ic_cap*ic_cap+-1.00000e-07*ic_cap+2.09000e-05'
+ mcm4m2_ca_w_0_300_s_0_600 = '-1.68750e-07*ic_cap*ic_cap+-1.00000e-07*ic_cap+2.09000e-05'
+ mcm4m2_ca_w_0_300_s_0_800 = '-1.68750e-07*ic_cap*ic_cap+-1.00000e-07*ic_cap+2.09000e-05'
+ mcm4m2_ca_w_0_300_s_1_000 = '-1.68750e-07*ic_cap*ic_cap+-1.00000e-07*ic_cap+2.09000e-05'
+ mcm4m2_ca_w_0_300_s_1_200 = '-1.68750e-07*ic_cap*ic_cap+-1.00000e-07*ic_cap+2.09000e-05'
+ mcm4m2_ca_w_0_300_s_2_100 = '-1.68750e-07*ic_cap*ic_cap+-1.00000e-07*ic_cap+2.09000e-05'
+ mcm4m2_ca_w_0_300_s_3_300 = '-1.68750e-07*ic_cap*ic_cap+-1.00000e-07*ic_cap+2.09000e-05'
+ mcm4m2_ca_w_0_300_s_9_000 = '-1.68750e-07*ic_cap*ic_cap+-1.00000e-07*ic_cap+2.09000e-05'
+ mcm4m2_ca_w_2_400_s_0_300 = '-1.68750e-07*ic_cap*ic_cap+-1.00000e-07*ic_cap+2.09000e-05'
+ mcm4m2_ca_w_2_400_s_0_360 = '-1.68750e-07*ic_cap*ic_cap+-1.00000e-07*ic_cap+2.09000e-05'
+ mcm4m2_ca_w_2_400_s_0_450 = '-1.68750e-07*ic_cap*ic_cap+-1.00000e-07*ic_cap+2.09000e-05'
+ mcm4m2_ca_w_2_400_s_0_600 = '-1.68750e-07*ic_cap*ic_cap+-1.00000e-07*ic_cap+2.09000e-05'
+ mcm4m2_ca_w_2_400_s_0_800 = '-1.68750e-07*ic_cap*ic_cap+-1.00000e-07*ic_cap+2.09000e-05'
+ mcm4m2_ca_w_2_400_s_1_000 = '-1.68750e-07*ic_cap*ic_cap+-1.00000e-07*ic_cap+2.09000e-05'
+ mcm4m2_ca_w_2_400_s_1_200 = '-1.68750e-07*ic_cap*ic_cap+-1.00000e-07*ic_cap+2.09000e-05'
+ mcm4m2_ca_w_2_400_s_2_100 = '-1.68750e-07*ic_cap*ic_cap+-1.00000e-07*ic_cap+2.09000e-05'
+ mcm4m2_ca_w_2_400_s_3_300 = '-1.68750e-07*ic_cap*ic_cap+-1.00000e-07*ic_cap+2.09000e-05'
+ mcm4m2_ca_w_2_400_s_9_000 = '-1.68750e-07*ic_cap*ic_cap+-1.00000e-07*ic_cap+2.09000e-05'
+ mcm4m2_cc_w_0_300_s_0_300 = '-8.09375e-13*ic_cap*ic_cap+-4.62500e-13*ic_cap+1.05000e-10'
+ mcm4m2_cc_w_0_300_s_0_360 = '-7.06250e-13*ic_cap*ic_cap+-4.00000e-13*ic_cap+9.77000e-11'
+ mcm4m2_cc_w_0_300_s_0_450 = '-5.90625e-13*ic_cap*ic_cap+-3.62500e-13*ic_cap+8.80000e-11'
+ mcm4m2_cc_w_0_300_s_0_600 = '-4.62500e-13*ic_cap*ic_cap+-3.00000e-13*ic_cap+7.54000e-11'
+ mcm4m2_cc_w_0_300_s_0_800 = '-3.34375e-13*ic_cap*ic_cap+-2.12500e-13*ic_cap+6.31000e-11'
+ mcm4m2_cc_w_0_300_s_1_000 = '-2.56250e-13*ic_cap*ic_cap+-1.75000e-13*ic_cap+5.38000e-11'
+ mcm4m2_cc_w_0_300_s_1_200 = '-2.00000e-13*ic_cap*ic_cap+-1.25000e-13*ic_cap+4.68000e-11'
+ mcm4m2_cc_w_0_300_s_2_100 = '-8.12500e-14*ic_cap*ic_cap+-5.00000e-14*ic_cap+2.90000e-11'
+ mcm4m2_cc_w_0_300_s_3_300 = '-3.75000e-14*ic_cap*ic_cap+-2.50000e-14*ic_cap+1.88000e-11'
+ mcm4m2_cc_w_0_300_s_9_000 = '4.68750e-15*ic_cap*ic_cap+3.75000e-15*ic_cap+4.49000e-12'
+ mcm4m2_cc_w_2_400_s_0_300 = '-8.12500e-13*ic_cap*ic_cap+-5.00000e-13*ic_cap+1.28000e-10'
+ mcm4m2_cc_w_2_400_s_0_360 = '-7.18750e-13*ic_cap*ic_cap+-3.75000e-13*ic_cap+1.20000e-10'
+ mcm4m2_cc_w_2_400_s_0_450 = '-5.34375e-13*ic_cap*ic_cap+-3.87500e-13*ic_cap+1.08000e-10'
+ mcm4m2_cc_w_2_400_s_0_600 = '-4.40625e-13*ic_cap*ic_cap+-2.62500e-13*ic_cap+9.36000e-11'
+ mcm4m2_cc_w_2_400_s_0_800 = '-3.09375e-13*ic_cap*ic_cap+-1.87500e-13*ic_cap+7.88000e-11'
+ mcm4m2_cc_w_2_400_s_1_000 = '-2.28125e-13*ic_cap*ic_cap+-1.62500e-13*ic_cap+6.78000e-11'
+ mcm4m2_cc_w_2_400_s_1_200 = '-1.65625e-13*ic_cap*ic_cap+-1.12500e-13*ic_cap+5.95000e-11'
+ mcm4m2_cc_w_2_400_s_2_100 = '-6.87500e-14*ic_cap*ic_cap+-5.00000e-14*ic_cap+3.89000e-11'
+ mcm4m2_cc_w_2_400_s_3_300 = '-1.87500e-14*ic_cap*ic_cap+-2.50000e-14*ic_cap+2.59000e-11'
+ mcm4m2_cc_w_2_400_s_9_000 = '1.25000e-14*ic_cap*ic_cap+1.25000e-14*ic_cap+7.40000e-12'
+ mcm4m2_cf_w_0_300_s_0_300 = '-2.18750e-15*ic_cap*ic_cap+-1.25000e-15*ic_cap+3.04000e-12'
+ mcm4m2_cf_w_0_300_s_0_360 = '-6.87500e-15*ic_cap*ic_cap+-5.00000e-15*ic_cap+3.63000e-12'
+ mcm4m2_cf_w_0_300_s_0_450 = '-1.34375e-14*ic_cap*ic_cap+-8.75000e-15*ic_cap+4.52000e-12'
+ mcm4m2_cf_w_0_300_s_0_600 = '-2.43750e-14*ic_cap*ic_cap+-1.50000e-14*ic_cap+5.97000e-12'
+ mcm4m2_cf_w_0_300_s_0_800 = '-3.93750e-14*ic_cap*ic_cap+-2.50000e-14*ic_cap+7.72000e-12'
+ mcm4m2_cf_w_0_300_s_1_000 = '-5.28125e-14*ic_cap*ic_cap+-3.12500e-14*ic_cap+9.44000e-12'
+ mcm4m2_cf_w_0_300_s_1_200 = '-6.59375e-14*ic_cap*ic_cap+-3.87500e-14*ic_cap+1.11000e-11'
+ mcm4m2_cf_w_0_300_s_2_100 = '-1.03125e-13*ic_cap*ic_cap+-6.25000e-14*ic_cap+1.78000e-11'
+ mcm4m2_cf_w_0_300_s_3_300 = '-1.40625e-13*ic_cap*ic_cap+-8.75000e-14*ic_cap+2.38000e-11'
+ mcm4m2_cf_w_0_300_s_9_000 = '-1.78125e-13*ic_cap*ic_cap+-1.12500e-13*ic_cap+3.56000e-11'
+ mcm4m2_cf_w_2_400_s_0_300 = '-2.18750e-15*ic_cap*ic_cap+-1.25000e-15*ic_cap+3.05000e-12'
+ mcm4m2_cf_w_2_400_s_0_360 = '-6.87500e-15*ic_cap*ic_cap+-5.00000e-15*ic_cap+3.64000e-12'
+ mcm4m2_cf_w_2_400_s_0_450 = '-1.40625e-14*ic_cap*ic_cap+-8.75000e-15*ic_cap+4.52000e-12'
+ mcm4m2_cf_w_2_400_s_0_600 = '-2.46875e-14*ic_cap*ic_cap+-1.62500e-14*ic_cap+5.93000e-12'
+ mcm4m2_cf_w_2_400_s_0_800 = '-3.87500e-14*ic_cap*ic_cap+-2.50000e-14*ic_cap+7.76000e-12'
+ mcm4m2_cf_w_2_400_s_1_000 = '-5.28125e-14*ic_cap*ic_cap+-3.37500e-14*ic_cap+9.53000e-12'
+ mcm4m2_cf_w_2_400_s_1_200 = '-6.56250e-14*ic_cap*ic_cap+-3.75000e-14*ic_cap+1.12000e-11'
+ mcm4m2_cf_w_2_400_s_2_100 = '-1.06250e-13*ic_cap*ic_cap+-7.50000e-14*ic_cap+1.78000e-11'
+ mcm4m2_cf_w_2_400_s_3_300 = '-1.40625e-13*ic_cap*ic_cap+-8.75000e-14*ic_cap+2.46000e-11'
+ mcm4m2_cf_w_2_400_s_9_000 = '-1.71875e-13*ic_cap*ic_cap+-1.12500e-13*ic_cap+3.92000e-11'
+ mcm4m2d_ca_w_0_140_s_0_140 = '-3.84375e-07*ic_cap*ic_cap+-2.37500e-07*ic_cap+4.17000e-05'
+ mcm4m2d_ca_w_0_140_s_0_175 = '-3.84375e-07*ic_cap*ic_cap+-2.37500e-07*ic_cap+4.17000e-05'
+ mcm4m2d_ca_w_0_140_s_0_210 = '-3.84375e-07*ic_cap*ic_cap+-2.37500e-07*ic_cap+4.17000e-05'
+ mcm4m2d_ca_w_0_140_s_0_280 = '-3.84375e-07*ic_cap*ic_cap+-2.37500e-07*ic_cap+4.17000e-05'
+ mcm4m2d_ca_w_0_140_s_0_350 = '-3.84375e-07*ic_cap*ic_cap+-2.37500e-07*ic_cap+4.17000e-05'
+ mcm4m2d_ca_w_0_140_s_0_420 = '-3.84375e-07*ic_cap*ic_cap+-2.37500e-07*ic_cap+4.17000e-05'
+ mcm4m2d_ca_w_0_140_s_0_560 = '-3.84375e-07*ic_cap*ic_cap+-2.37500e-07*ic_cap+4.17000e-05'
+ mcm4m2d_ca_w_0_140_s_0_840 = '-3.84375e-07*ic_cap*ic_cap+-2.37500e-07*ic_cap+4.17000e-05'
+ mcm4m2d_ca_w_0_140_s_1_540 = '-3.84375e-07*ic_cap*ic_cap+-2.37500e-07*ic_cap+4.17000e-05'
+ mcm4m2d_ca_w_0_140_s_3_500 = '-3.84375e-07*ic_cap*ic_cap+-2.37500e-07*ic_cap+4.17000e-05'
+ mcm4m2d_ca_w_1_120_s_0_140 = '-3.84375e-07*ic_cap*ic_cap+-2.37500e-07*ic_cap+4.17000e-05'
+ mcm4m2d_ca_w_1_120_s_0_175 = '-3.84375e-07*ic_cap*ic_cap+-2.37500e-07*ic_cap+4.17000e-05'
+ mcm4m2d_ca_w_1_120_s_0_210 = '-3.84375e-07*ic_cap*ic_cap+-2.37500e-07*ic_cap+4.17000e-05'
+ mcm4m2d_ca_w_1_120_s_0_280 = '-3.84375e-07*ic_cap*ic_cap+-2.37500e-07*ic_cap+4.17000e-05'
+ mcm4m2d_ca_w_1_120_s_0_350 = '-3.84375e-07*ic_cap*ic_cap+-2.37500e-07*ic_cap+4.17000e-05'
+ mcm4m2d_ca_w_1_120_s_0_420 = '-3.84375e-07*ic_cap*ic_cap+-2.37500e-07*ic_cap+4.17000e-05'
+ mcm4m2d_ca_w_1_120_s_0_560 = '-3.84375e-07*ic_cap*ic_cap+-2.37500e-07*ic_cap+4.17000e-05'
+ mcm4m2d_ca_w_1_120_s_0_840 = '-3.84375e-07*ic_cap*ic_cap+-2.37500e-07*ic_cap+4.17000e-05'
+ mcm4m2d_ca_w_1_120_s_1_540 = '-3.84375e-07*ic_cap*ic_cap+-2.37500e-07*ic_cap+4.17000e-05'
+ mcm4m2d_ca_w_1_120_s_3_500 = '-3.84375e-07*ic_cap*ic_cap+-2.37500e-07*ic_cap+4.17000e-05'
+ mcm4m2d_cc_w_0_140_s_0_140 = '-9.18750e-13*ic_cap*ic_cap+-5.25000e-13*ic_cap+1.03000e-10'
+ mcm4m2d_cc_w_0_140_s_0_175 = '-8.46875e-13*ic_cap*ic_cap+-5.87500e-13*ic_cap+1.01000e-10'
+ mcm4m2d_cc_w_0_140_s_0_210 = '-7.75000e-13*ic_cap*ic_cap+-4.25000e-13*ic_cap+9.60000e-11'
+ mcm4m2d_cc_w_0_140_s_0_280 = '-5.68750e-13*ic_cap*ic_cap+-4.00000e-13*ic_cap+8.45000e-11'
+ mcm4m2d_cc_w_0_140_s_0_350 = '-4.53125e-13*ic_cap*ic_cap+-2.62500e-13*ic_cap+7.30000e-11'
+ mcm4m2d_cc_w_0_140_s_0_420 = '-3.15625e-13*ic_cap*ic_cap+-2.12500e-13*ic_cap+6.31000e-11'
+ mcm4m2d_cc_w_0_140_s_0_560 = '-1.62500e-13*ic_cap*ic_cap+-1.25000e-13*ic_cap+4.95000e-11'
+ mcm4m2d_cc_w_0_140_s_0_840 = '-5.31250e-14*ic_cap*ic_cap+-3.75000e-14*ic_cap+3.42000e-11'
+ mcm4m2d_cc_w_0_140_s_1_540 = '5.62500e-14*ic_cap*ic_cap+2.50000e-14*ic_cap+1.64000e-11'
+ mcm4m2d_cc_w_0_140_s_3_500 = '5.03125e-14*ic_cap*ic_cap+3.62500e-14*ic_cap+2.93000e-12'
+ mcm4m2d_cc_w_1_120_s_0_140 = '-7.81250e-13*ic_cap*ic_cap+-3.75000e-13*ic_cap+1.22000e-10'
+ mcm4m2d_cc_w_1_120_s_0_175 = '-7.18750e-13*ic_cap*ic_cap+-3.75000e-13*ic_cap+1.18000e-10'
+ mcm4m2d_cc_w_1_120_s_0_210 = '-5.62500e-13*ic_cap*ic_cap+-2.50000e-13*ic_cap+1.11000e-10'
+ mcm4m2d_cc_w_1_120_s_0_280 = '-4.18750e-13*ic_cap*ic_cap+-2.50000e-13*ic_cap+9.72000e-11'
+ mcm4m2d_cc_w_1_120_s_0_350 = '-3.18750e-13*ic_cap*ic_cap+-2.25000e-13*ic_cap+8.44000e-11'
+ mcm4m2d_cc_w_1_120_s_0_420 = '-2.09375e-13*ic_cap*ic_cap+-1.37500e-13*ic_cap+7.34000e-11'
+ mcm4m2d_cc_w_1_120_s_0_560 = '-7.18750e-14*ic_cap*ic_cap+-6.25000e-14*ic_cap+5.76000e-11'
+ mcm4m2d_cc_w_1_120_s_0_840 = '3.12500e-14*ic_cap*ic_cap+2.50000e-14*ic_cap+3.96000e-11'
+ mcm4m2d_cc_w_1_120_s_1_540 = '1.09375e-13*ic_cap*ic_cap+6.25000e-14*ic_cap+1.93000e-11'
+ mcm4m2d_cc_w_1_120_s_3_500 = '7.31250e-14*ic_cap*ic_cap+5.00000e-14*ic_cap+3.51000e-12'
+ mcm4m2d_cf_w_0_140_s_0_140 = '1.25000e-15*ic_cap*ic_cap+2.89000e-12'
+ mcm4m2d_cf_w_0_140_s_0_175 = '-5.62500e-15*ic_cap*ic_cap+-5.00000e-15*ic_cap+3.60000e-12'
+ mcm4m2d_cf_w_0_140_s_0_210 = '-1.00000e-14*ic_cap*ic_cap+-7.50000e-15*ic_cap+4.32000e-12'
+ mcm4m2d_cf_w_0_140_s_0_280 = '-2.46875e-14*ic_cap*ic_cap+-1.62500e-14*ic_cap+5.73000e-12'
+ mcm4m2d_cf_w_0_140_s_0_350 = '-3.71875e-14*ic_cap*ic_cap+-2.37500e-14*ic_cap+7.10000e-12'
+ mcm4m2d_cf_w_0_140_s_0_420 = '-4.96875e-14*ic_cap*ic_cap+-3.37500e-14*ic_cap+8.52000e-12'
+ mcm4m2d_cf_w_0_140_s_0_560 = '-7.28125e-14*ic_cap*ic_cap+-4.12500e-14*ic_cap+1.11000e-11'
+ mcm4m2d_cf_w_0_140_s_0_840 = '-1.18750e-13*ic_cap*ic_cap+-7.50000e-14*ic_cap+1.59000e-11'
+ mcm4m2d_cf_w_0_140_s_1_540 = '-1.84375e-13*ic_cap*ic_cap+-1.12500e-13*ic_cap+2.51000e-11'
+ mcm4m2d_cf_w_0_140_s_3_500 = '-2.15625e-13*ic_cap*ic_cap+-1.37500e-13*ic_cap+3.60000e-11'
+ mcm4m2d_cf_w_1_120_s_0_140 = '9.37500e-16*ic_cap*ic_cap+-1.25000e-15*ic_cap+2.92000e-12'
+ mcm4m2d_cf_w_1_120_s_0_175 = '-5.93750e-15*ic_cap*ic_cap+-3.75000e-15*ic_cap+3.64000e-12'
+ mcm4m2d_cf_w_1_120_s_0_210 = '-1.21875e-14*ic_cap*ic_cap+-8.75000e-15*ic_cap+4.35000e-12'
+ mcm4m2d_cf_w_1_120_s_0_280 = '-2.50000e-14*ic_cap*ic_cap+-1.75000e-14*ic_cap+5.76000e-12'
+ mcm4m2d_cf_w_1_120_s_0_350 = '-3.81250e-14*ic_cap*ic_cap+-2.50000e-14*ic_cap+7.16000e-12'
+ mcm4m2d_cf_w_1_120_s_0_420 = '-4.87500e-14*ic_cap*ic_cap+-3.50000e-14*ic_cap+8.53000e-12'
+ mcm4m2d_cf_w_1_120_s_0_560 = '-7.53125e-14*ic_cap*ic_cap+-5.12500e-14*ic_cap+1.12000e-11'
+ mcm4m2d_cf_w_1_120_s_0_840 = '-1.18750e-13*ic_cap*ic_cap+-7.50000e-14*ic_cap+1.61000e-11'
+ mcm4m2d_cf_w_1_120_s_1_540 = '-1.81250e-13*ic_cap*ic_cap+-1.25000e-13*ic_cap+2.58000e-11'
+ mcm4m2d_cf_w_1_120_s_3_500 = '-1.93750e-13*ic_cap*ic_cap+-1.25000e-13*ic_cap+3.81000e-11'
+ mcm4m2f_ca_w_0_140_s_0_140 = '-3.62500e-07*ic_cap*ic_cap+-2.25000e-07*ic_cap+3.84000e-05'
+ mcm4m2f_ca_w_0_140_s_0_175 = '-3.62500e-07*ic_cap*ic_cap+-2.25000e-07*ic_cap+3.84000e-05'
+ mcm4m2f_ca_w_0_140_s_0_210 = '-3.62500e-07*ic_cap*ic_cap+-2.25000e-07*ic_cap+3.84000e-05'
+ mcm4m2f_ca_w_0_140_s_0_280 = '-3.62500e-07*ic_cap*ic_cap+-2.25000e-07*ic_cap+3.84000e-05'
+ mcm4m2f_ca_w_0_140_s_0_350 = '-3.62500e-07*ic_cap*ic_cap+-2.25000e-07*ic_cap+3.84000e-05'
+ mcm4m2f_ca_w_0_140_s_0_420 = '-3.62500e-07*ic_cap*ic_cap+-2.25000e-07*ic_cap+3.84000e-05'
+ mcm4m2f_ca_w_0_140_s_0_560 = '-3.62500e-07*ic_cap*ic_cap+-2.25000e-07*ic_cap+3.84000e-05'
+ mcm4m2f_ca_w_0_140_s_0_840 = '-3.62500e-07*ic_cap*ic_cap+-2.25000e-07*ic_cap+3.84000e-05'
+ mcm4m2f_ca_w_0_140_s_1_540 = '-3.62500e-07*ic_cap*ic_cap+-2.25000e-07*ic_cap+3.84000e-05'
+ mcm4m2f_ca_w_0_140_s_3_500 = '-3.62500e-07*ic_cap*ic_cap+-2.25000e-07*ic_cap+3.84000e-05'
+ mcm4m2f_ca_w_1_120_s_0_140 = '-3.62500e-07*ic_cap*ic_cap+-2.25000e-07*ic_cap+3.84000e-05'
+ mcm4m2f_ca_w_1_120_s_0_175 = '-3.62500e-07*ic_cap*ic_cap+-2.25000e-07*ic_cap+3.84000e-05'
+ mcm4m2f_ca_w_1_120_s_0_210 = '-3.62500e-07*ic_cap*ic_cap+-2.25000e-07*ic_cap+3.84000e-05'
+ mcm4m2f_ca_w_1_120_s_0_280 = '-3.62500e-07*ic_cap*ic_cap+-2.25000e-07*ic_cap+3.84000e-05'
+ mcm4m2f_ca_w_1_120_s_0_350 = '-3.62500e-07*ic_cap*ic_cap+-2.25000e-07*ic_cap+3.84000e-05'
+ mcm4m2f_ca_w_1_120_s_0_420 = '-3.62500e-07*ic_cap*ic_cap+-2.25000e-07*ic_cap+3.84000e-05'
+ mcm4m2f_ca_w_1_120_s_0_560 = '-3.62500e-07*ic_cap*ic_cap+-2.25000e-07*ic_cap+3.84000e-05'
+ mcm4m2f_ca_w_1_120_s_0_840 = '-3.62500e-07*ic_cap*ic_cap+-2.25000e-07*ic_cap+3.84000e-05'
+ mcm4m2f_ca_w_1_120_s_1_540 = '-3.62500e-07*ic_cap*ic_cap+-2.25000e-07*ic_cap+3.84000e-05'
+ mcm4m2f_ca_w_1_120_s_3_500 = '-3.62500e-07*ic_cap*ic_cap+-2.25000e-07*ic_cap+3.84000e-05'
+ mcm4m2f_cc_w_0_140_s_0_140 = '-9.46875e-13*ic_cap*ic_cap+-4.87500e-13*ic_cap+1.04000e-10'
+ mcm4m2f_cc_w_0_140_s_0_175 = '-8.84375e-13*ic_cap*ic_cap+-5.87500e-13*ic_cap+1.02000e-10'
+ mcm4m2f_cc_w_0_140_s_0_210 = '-7.75000e-13*ic_cap*ic_cap+-4.25000e-13*ic_cap+9.64000e-11'
+ mcm4m2f_cc_w_0_140_s_0_280 = '-5.71875e-13*ic_cap*ic_cap+-4.12500e-13*ic_cap+8.50000e-11'
+ mcm4m2f_cc_w_0_140_s_0_350 = '-4.62500e-13*ic_cap*ic_cap+-2.75000e-13*ic_cap+7.37000e-11'
+ mcm4m2f_cc_w_0_140_s_0_420 = '-3.34375e-13*ic_cap*ic_cap+-1.62500e-13*ic_cap+6.38000e-11'
+ mcm4m2f_cc_w_0_140_s_0_560 = '-1.81250e-13*ic_cap*ic_cap+-7.50000e-14*ic_cap+5.04000e-11'
+ mcm4m2f_cc_w_0_140_s_0_840 = '-4.68750e-14*ic_cap*ic_cap+-3.75000e-14*ic_cap+3.52000e-11'
+ mcm4m2f_cc_w_0_140_s_1_540 = '5.00000e-14*ic_cap*ic_cap+2.50000e-14*ic_cap+1.76000e-11'
+ mcm4m2f_cc_w_0_140_s_3_500 = '5.62500e-14*ic_cap*ic_cap+4.00000e-14*ic_cap+3.53000e-12'
+ mcm4m2f_cc_w_1_120_s_0_140 = '-7.50000e-13*ic_cap*ic_cap+-5.00000e-13*ic_cap+1.23000e-10'
+ mcm4m2f_cc_w_1_120_s_0_175 = '-7.81250e-13*ic_cap*ic_cap+-3.75000e-13*ic_cap+1.20000e-10'
+ mcm4m2f_cc_w_1_120_s_0_210 = '-5.93750e-13*ic_cap*ic_cap+-3.75000e-13*ic_cap+1.13000e-10'
+ mcm4m2f_cc_w_1_120_s_0_280 = '-4.37500e-13*ic_cap*ic_cap+-3.25000e-13*ic_cap+9.86000e-11'
+ mcm4m2f_cc_w_1_120_s_0_350 = '-3.25000e-13*ic_cap*ic_cap+-2.50000e-13*ic_cap+8.59000e-11'
+ mcm4m2f_cc_w_1_120_s_0_420 = '-2.28125e-13*ic_cap*ic_cap+-1.12500e-13*ic_cap+7.50000e-11'
+ mcm4m2f_cc_w_1_120_s_0_560 = '-7.18750e-14*ic_cap*ic_cap+-6.25000e-14*ic_cap+5.92000e-11'
+ mcm4m2f_cc_w_1_120_s_0_840 = '2.81250e-14*ic_cap*ic_cap+1.25000e-14*ic_cap+4.13000e-11'
+ mcm4m2f_cc_w_1_120_s_1_540 = '1.06250e-13*ic_cap*ic_cap+7.50000e-14*ic_cap+2.09000e-11'
+ mcm4m2f_cc_w_1_120_s_3_500 = '8.15625e-14*ic_cap*ic_cap+6.12500e-14*ic_cap+4.30000e-12'
+ mcm4m2f_cf_w_0_140_s_0_140 = '6.25000e-16*ic_cap*ic_cap+2.66000e-12'
+ mcm4m2f_cf_w_0_140_s_0_175 = '-5.31250e-15*ic_cap*ic_cap+-3.75000e-15*ic_cap+3.31000e-12'
+ mcm4m2f_cf_w_0_140_s_0_210 = '-1.00000e-14*ic_cap*ic_cap+-7.50000e-15*ic_cap+3.98000e-12'
+ mcm4m2f_cf_w_0_140_s_0_280 = '-2.37500e-14*ic_cap*ic_cap+-1.50000e-14*ic_cap+5.28000e-12'
+ mcm4m2f_cf_w_0_140_s_0_350 = '-3.46875e-14*ic_cap*ic_cap+-2.12500e-14*ic_cap+6.53000e-12'
+ mcm4m2f_cf_w_0_140_s_0_420 = '-4.84375e-14*ic_cap*ic_cap+-2.62500e-14*ic_cap+7.86000e-12'
+ mcm4m2f_cf_w_0_140_s_0_560 = '-7.18750e-14*ic_cap*ic_cap+-4.00000e-14*ic_cap+1.03000e-11'
+ mcm4m2f_cf_w_0_140_s_0_840 = '-1.09375e-13*ic_cap*ic_cap+-6.25000e-14*ic_cap+1.47000e-11'
+ mcm4m2f_cf_w_0_140_s_1_540 = '-1.78125e-13*ic_cap*ic_cap+-1.12500e-13*ic_cap+2.35000e-11'
+ mcm4m2f_cf_w_0_140_s_3_500 = '-2.06250e-13*ic_cap*ic_cap+-1.25000e-13*ic_cap+3.44000e-11'
+ mcm4m2f_cf_w_1_120_s_0_175 = '-5.31250e-15*ic_cap*ic_cap+-3.75000e-15*ic_cap+3.34000e-12'
+ mcm4m2f_cf_w_1_120_s_0_210 = '-1.18750e-14*ic_cap*ic_cap+-7.50000e-15*ic_cap+4.00000e-12'
+ mcm4m2f_cf_w_1_120_s_0_280 = '-2.34375e-14*ic_cap*ic_cap+-1.37500e-14*ic_cap+5.30000e-12'
+ mcm4m2f_cf_w_1_120_s_0_350 = '-3.56250e-14*ic_cap*ic_cap+-2.25000e-14*ic_cap+6.58000e-12'
+ mcm4m2f_cf_w_1_120_s_0_420 = '-4.68750e-14*ic_cap*ic_cap+-2.75000e-14*ic_cap+7.85000e-12'
+ mcm4m2f_cf_w_1_120_s_0_560 = '-7.03125e-14*ic_cap*ic_cap+-4.37500e-14*ic_cap+1.03000e-11'
+ mcm4m2f_cf_w_1_120_s_0_840 = '-1.12500e-13*ic_cap*ic_cap+-7.50000e-14*ic_cap+1.49000e-11'
+ mcm4m2f_cf_w_1_120_s_1_540 = '-1.78125e-13*ic_cap*ic_cap+-1.12500e-13*ic_cap+2.42000e-11'
+ mcm4m2f_cf_w_1_120_s_3_500 = '-1.93750e-13*ic_cap*ic_cap+-1.25000e-13*ic_cap+3.66000e-11'
+ mcm4m2l1_ca_w_0_140_s_0_140 = '-6.21875e-07*ic_cap*ic_cap+-3.87500e-07*ic_cap+5.79000e-05'
+ mcm4m2l1_ca_w_0_140_s_0_175 = '-6.21875e-07*ic_cap*ic_cap+-3.87500e-07*ic_cap+5.79000e-05'
+ mcm4m2l1_ca_w_0_140_s_0_210 = '-6.21875e-07*ic_cap*ic_cap+-3.87500e-07*ic_cap+5.79000e-05'
+ mcm4m2l1_ca_w_0_140_s_0_280 = '-6.21875e-07*ic_cap*ic_cap+-3.87500e-07*ic_cap+5.79000e-05'
+ mcm4m2l1_ca_w_0_140_s_0_350 = '-6.21875e-07*ic_cap*ic_cap+-3.87500e-07*ic_cap+5.79000e-05'
+ mcm4m2l1_ca_w_0_140_s_0_420 = '-6.21875e-07*ic_cap*ic_cap+-3.87500e-07*ic_cap+5.79000e-05'
+ mcm4m2l1_ca_w_0_140_s_0_560 = '-6.21875e-07*ic_cap*ic_cap+-3.87500e-07*ic_cap+5.79000e-05'
+ mcm4m2l1_ca_w_0_140_s_0_840 = '-6.21875e-07*ic_cap*ic_cap+-3.87500e-07*ic_cap+5.79000e-05'
+ mcm4m2l1_ca_w_0_140_s_1_540 = '-6.21875e-07*ic_cap*ic_cap+-3.87500e-07*ic_cap+5.79000e-05'
+ mcm4m2l1_ca_w_0_140_s_3_500 = '-6.21875e-07*ic_cap*ic_cap+-3.87500e-07*ic_cap+5.79000e-05'
+ mcm4m2l1_ca_w_1_120_s_0_140 = '-6.21875e-07*ic_cap*ic_cap+-3.87500e-07*ic_cap+5.79000e-05'
+ mcm4m2l1_ca_w_1_120_s_0_175 = '-6.21875e-07*ic_cap*ic_cap+-3.87500e-07*ic_cap+5.79000e-05'
+ mcm4m2l1_ca_w_1_120_s_0_210 = '-6.21875e-07*ic_cap*ic_cap+-3.87500e-07*ic_cap+5.79000e-05'
+ mcm4m2l1_ca_w_1_120_s_0_280 = '-6.21875e-07*ic_cap*ic_cap+-3.87500e-07*ic_cap+5.79000e-05'
+ mcm4m2l1_ca_w_1_120_s_0_350 = '-6.21875e-07*ic_cap*ic_cap+-3.87500e-07*ic_cap+5.79000e-05'
+ mcm4m2l1_ca_w_1_120_s_0_420 = '-6.21875e-07*ic_cap*ic_cap+-3.87500e-07*ic_cap+5.79000e-05'
+ mcm4m2l1_ca_w_1_120_s_0_560 = '-6.21875e-07*ic_cap*ic_cap+-3.87500e-07*ic_cap+5.79000e-05'
+ mcm4m2l1_ca_w_1_120_s_0_840 = '-6.21875e-07*ic_cap*ic_cap+-3.87500e-07*ic_cap+5.79000e-05'
+ mcm4m2l1_ca_w_1_120_s_1_540 = '-6.21875e-07*ic_cap*ic_cap+-3.87500e-07*ic_cap+5.79000e-05'
+ mcm4m2l1_ca_w_1_120_s_3_500 = '-6.21875e-07*ic_cap*ic_cap+-3.87500e-07*ic_cap+5.79000e-05'
+ mcm4m2l1_cc_w_0_140_s_0_140 = '-8.84375e-13*ic_cap*ic_cap+-5.12500e-13*ic_cap+1.01000e-10'
+ mcm4m2l1_cc_w_0_140_s_0_175 = '-8.12500e-13*ic_cap*ic_cap+-5.50000e-13*ic_cap+9.91000e-11'
+ mcm4m2l1_cc_w_0_140_s_0_210 = '-7.06250e-13*ic_cap*ic_cap+-3.75000e-13*ic_cap+9.33000e-11'
+ mcm4m2l1_cc_w_0_140_s_0_280 = '-5.18750e-13*ic_cap*ic_cap+-3.75000e-13*ic_cap+8.16000e-11'
+ mcm4m2l1_cc_w_0_140_s_0_350 = '-3.90625e-13*ic_cap*ic_cap+-2.37500e-13*ic_cap+6.99000e-11'
+ mcm4m2l1_cc_w_0_140_s_0_420 = '-2.96875e-13*ic_cap*ic_cap+-1.87500e-13*ic_cap+5.99000e-11'
+ mcm4m2l1_cc_w_0_140_s_0_560 = '-1.40625e-13*ic_cap*ic_cap+-8.75000e-14*ic_cap+4.60000e-11'
+ mcm4m2l1_cc_w_0_140_s_0_840 = '-6.25000e-15*ic_cap*ic_cap+2.99000e-11'
+ mcm4m2l1_cc_w_0_140_s_1_540 = '8.12500e-14*ic_cap*ic_cap+5.00000e-14*ic_cap+1.24000e-11'
+ mcm4m2l1_cc_w_0_140_s_3_500 = '3.81250e-14*ic_cap*ic_cap+3.00000e-14*ic_cap+1.46000e-12'
+ mcm4m2l1_cc_w_1_120_s_0_140 = '-7.18750e-13*ic_cap*ic_cap+-3.75000e-13*ic_cap+1.16000e-10'
+ mcm4m2l1_cc_w_1_120_s_0_175 = '-7.50000e-13*ic_cap*ic_cap+-2.50000e-13*ic_cap+1.13000e-10'
+ mcm4m2l1_cc_w_1_120_s_0_210 = '-5.59375e-13*ic_cap*ic_cap+-3.37500e-13*ic_cap+1.06000e-10'
+ mcm4m2l1_cc_w_1_120_s_0_280 = '-3.62500e-13*ic_cap*ic_cap+-2.25000e-13*ic_cap+9.13000e-11'
+ mcm4m2l1_cc_w_1_120_s_0_350 = '-2.71875e-13*ic_cap*ic_cap+-1.37500e-13*ic_cap+7.86000e-11'
+ mcm4m2l1_cc_w_1_120_s_0_420 = '-1.46875e-13*ic_cap*ic_cap+-1.12500e-13*ic_cap+6.73000e-11'
+ mcm4m2l1_cc_w_1_120_s_0_560 = '-3.12500e-14*ic_cap*ic_cap+-2.50000e-14*ic_cap+5.17000e-11'
+ mcm4m2l1_cc_w_1_120_s_0_840 = '6.87500e-14*ic_cap*ic_cap+5.00000e-14*ic_cap+3.38000e-11'
+ mcm4m2l1_cc_w_1_120_s_1_540 = '1.15625e-13*ic_cap*ic_cap+8.75000e-14*ic_cap+1.44000e-11'
+ mcm4m2l1_cc_w_1_120_s_3_500 = '5.31250e-14*ic_cap*ic_cap+4.25000e-14*ic_cap+1.71000e-12'
+ mcm4m2l1_cf_w_0_140_s_0_140 = '-4.68750e-15*ic_cap*ic_cap+-6.25000e-15*ic_cap+3.98000e-12'
+ mcm4m2l1_cf_w_0_140_s_0_175 = '-1.53125e-14*ic_cap*ic_cap+-1.12500e-14*ic_cap+4.97000e-12'
+ mcm4m2l1_cf_w_0_140_s_0_210 = '-2.43750e-14*ic_cap*ic_cap+-1.75000e-14*ic_cap+5.97000e-12'
+ mcm4m2l1_cf_w_0_140_s_0_280 = '-4.59375e-14*ic_cap*ic_cap+-3.12500e-14*ic_cap+7.90000e-12'
+ mcm4m2l1_cf_w_0_140_s_0_350 = '-6.56250e-14*ic_cap*ic_cap+-4.50000e-14*ic_cap+9.78000e-12'
+ mcm4m2l1_cf_w_0_140_s_0_420 = '-8.75000e-14*ic_cap*ic_cap+-5.00000e-14*ic_cap+1.17000e-11'
+ mcm4m2l1_cf_w_0_140_s_0_560 = '-1.25000e-13*ic_cap*ic_cap+-7.50000e-14*ic_cap+1.52000e-11'
+ mcm4m2l1_cf_w_0_140_s_0_840 = '-1.81250e-13*ic_cap*ic_cap+-1.25000e-13*ic_cap+2.13000e-11'
+ mcm4m2l1_cf_w_0_140_s_1_540 = '-2.59375e-13*ic_cap*ic_cap+-1.62500e-13*ic_cap+3.21000e-11'
+ mcm4m2l1_cf_w_0_140_s_3_500 = '-2.46875e-13*ic_cap*ic_cap+-1.62500e-13*ic_cap+4.17000e-11'
+ mcm4m2l1_cf_w_1_120_s_0_140 = '-5.00000e-15*ic_cap*ic_cap+-5.00000e-15*ic_cap+4.01000e-12'
+ mcm4m2l1_cf_w_1_120_s_0_175 = '-1.59375e-14*ic_cap*ic_cap+-1.12500e-14*ic_cap+5.01000e-12'
+ mcm4m2l1_cf_w_1_120_s_0_210 = '-2.65625e-14*ic_cap*ic_cap+-1.87500e-14*ic_cap+6.00000e-12'
+ mcm4m2l1_cf_w_1_120_s_0_280 = '-4.65625e-14*ic_cap*ic_cap+-3.12500e-14*ic_cap+7.94000e-12'
+ mcm4m2l1_cf_w_1_120_s_0_350 = '-6.84375e-14*ic_cap*ic_cap+-4.37500e-14*ic_cap+9.87000e-12'
+ mcm4m2l1_cf_w_1_120_s_0_420 = '-8.43750e-14*ic_cap*ic_cap+-6.25000e-14*ic_cap+1.17000e-11'
+ mcm4m2l1_cf_w_1_120_s_0_560 = '-1.18750e-13*ic_cap*ic_cap+-7.50000e-14*ic_cap+1.52000e-11'
+ mcm4m2l1_cf_w_1_120_s_0_840 = '-1.81250e-13*ic_cap*ic_cap+-1.25000e-13*ic_cap+2.16000e-11'
+ mcm4m2l1_cf_w_1_120_s_1_540 = '-2.56250e-13*ic_cap*ic_cap+-1.75000e-13*ic_cap+3.30000e-11'
+ mcm4m2l1_cf_w_1_120_s_3_500 = '-2.21875e-13*ic_cap*ic_cap+-1.62500e-13*ic_cap+4.38000e-11'
+ mcm4m2m1_ca_w_0_140_s_0_140 = '-2.84062e-06*ic_cap*ic_cap+-1.36250e-06*ic_cap+1.49000e-04'
+ mcm4m2m1_ca_w_0_140_s_0_175 = '-2.84062e-06*ic_cap*ic_cap+-1.36250e-06*ic_cap+1.49000e-04'
+ mcm4m2m1_ca_w_0_140_s_0_210 = '-2.84062e-06*ic_cap*ic_cap+-1.36250e-06*ic_cap+1.49000e-04'
+ mcm4m2m1_ca_w_0_140_s_0_280 = '-2.84062e-06*ic_cap*ic_cap+-1.36250e-06*ic_cap+1.49000e-04'
+ mcm4m2m1_ca_w_0_140_s_0_350 = '-2.84062e-06*ic_cap*ic_cap+-1.36250e-06*ic_cap+1.49000e-04'
+ mcm4m2m1_ca_w_0_140_s_0_420 = '-2.84062e-06*ic_cap*ic_cap+-1.36250e-06*ic_cap+1.49000e-04'
+ mcm4m2m1_ca_w_0_140_s_0_560 = '-2.84062e-06*ic_cap*ic_cap+-1.36250e-06*ic_cap+1.49000e-04'
+ mcm4m2m1_ca_w_0_140_s_0_840 = '-2.84062e-06*ic_cap*ic_cap+-1.36250e-06*ic_cap+1.49000e-04'
+ mcm4m2m1_ca_w_0_140_s_1_540 = '-2.84062e-06*ic_cap*ic_cap+-1.36250e-06*ic_cap+1.49000e-04'
+ mcm4m2m1_ca_w_0_140_s_3_500 = '-2.84062e-06*ic_cap*ic_cap+-1.36250e-06*ic_cap+1.49000e-04'
+ mcm4m2m1_ca_w_1_120_s_0_140 = '-2.84062e-06*ic_cap*ic_cap+-1.36250e-06*ic_cap+1.49000e-04'
+ mcm4m2m1_ca_w_1_120_s_0_175 = '-2.84062e-06*ic_cap*ic_cap+-1.36250e-06*ic_cap+1.49000e-04'
+ mcm4m2m1_ca_w_1_120_s_0_210 = '-2.84062e-06*ic_cap*ic_cap+-1.36250e-06*ic_cap+1.49000e-04'
+ mcm4m2m1_ca_w_1_120_s_0_280 = '-2.84062e-06*ic_cap*ic_cap+-1.36250e-06*ic_cap+1.49000e-04'
+ mcm4m2m1_ca_w_1_120_s_0_350 = '-2.84062e-06*ic_cap*ic_cap+-1.36250e-06*ic_cap+1.49000e-04'
+ mcm4m2m1_ca_w_1_120_s_0_420 = '-2.84062e-06*ic_cap*ic_cap+-1.36250e-06*ic_cap+1.49000e-04'
+ mcm4m2m1_ca_w_1_120_s_0_560 = '-2.84062e-06*ic_cap*ic_cap+-1.36250e-06*ic_cap+1.49000e-04'
+ mcm4m2m1_ca_w_1_120_s_0_840 = '-2.84062e-06*ic_cap*ic_cap+-1.36250e-06*ic_cap+1.49000e-04'
+ mcm4m2m1_ca_w_1_120_s_1_540 = '-2.84062e-06*ic_cap*ic_cap+-1.36250e-06*ic_cap+1.49000e-04'
+ mcm4m2m1_ca_w_1_120_s_3_500 = '-2.84062e-06*ic_cap*ic_cap+-1.36250e-06*ic_cap+1.49000e-04'
+ mcm4m2m1_cc_w_0_140_s_0_140 = '-7.40625e-13*ic_cap*ic_cap+-3.37500e-13*ic_cap+9.29000e-11'
+ mcm4m2m1_cc_w_0_140_s_0_175 = '-6.93750e-13*ic_cap*ic_cap+-3.25000e-13*ic_cap+9.05000e-11'
+ mcm4m2m1_cc_w_0_140_s_0_210 = '-5.37500e-13*ic_cap*ic_cap+-3.25000e-13*ic_cap+8.43000e-11'
+ mcm4m2m1_cc_w_0_140_s_0_280 = '-3.43750e-13*ic_cap*ic_cap+-3.00000e-13*ic_cap+7.12000e-11'
+ mcm4m2m1_cc_w_0_140_s_0_350 = '-2.03125e-13*ic_cap*ic_cap+-1.37500e-13*ic_cap+5.89000e-11'
+ mcm4m2m1_cc_w_0_140_s_0_420 = '-1.06250e-13*ic_cap*ic_cap+-1.25000e-13*ic_cap+4.87000e-11'
+ mcm4m2m1_cc_w_0_140_s_0_560 = '1.87500e-14*ic_cap*ic_cap+-2.50000e-14*ic_cap+3.47000e-11'
+ mcm4m2m1_cc_w_0_140_s_0_840 = '9.68750e-14*ic_cap*ic_cap+6.25000e-14*ic_cap+1.95000e-11'
+ mcm4m2m1_cc_w_0_140_s_1_540 = '8.28125e-14*ic_cap*ic_cap+5.37500e-14*ic_cap+5.90000e-12'
+ mcm4m2m1_cc_w_0_140_s_3_500 = '1.51562e-14*ic_cap*ic_cap+9.37500e-15*ic_cap+3.95000e-13'
+ mcm4m2m1_cc_w_1_120_s_0_140 = '-5.37500e-13*ic_cap*ic_cap+-3.50000e-13*ic_cap+1.02000e-10'
+ mcm4m2m1_cc_w_1_120_s_0_175 = '-5.75000e-13*ic_cap*ic_cap+-2.25000e-13*ic_cap+9.96000e-11'
+ mcm4m2m1_cc_w_1_120_s_0_210 = '-4.28125e-13*ic_cap*ic_cap+-2.37500e-13*ic_cap+9.26000e-11'
+ mcm4m2m1_cc_w_1_120_s_0_280 = '-2.53125e-13*ic_cap*ic_cap+-1.37500e-13*ic_cap+7.82000e-11'
+ mcm4m2m1_cc_w_1_120_s_0_350 = '-1.34375e-13*ic_cap*ic_cap+-8.75000e-14*ic_cap+6.51000e-11'
+ mcm4m2m1_cc_w_1_120_s_0_420 = '-3.75000e-14*ic_cap*ic_cap+-5.00000e-14*ic_cap+5.43000e-11'
+ mcm4m2m1_cc_w_1_120_s_0_560 = '7.50000e-14*ic_cap*ic_cap+5.00000e-14*ic_cap+3.91000e-11'
+ mcm4m2m1_cc_w_1_120_s_0_840 = '1.31250e-13*ic_cap*ic_cap+7.50000e-14*ic_cap+2.27000e-11'
+ mcm4m2m1_cc_w_1_120_s_1_540 = '1.13750e-13*ic_cap*ic_cap+7.50000e-14*ic_cap+7.30000e-12'
+ mcm4m2m1_cc_w_1_120_s_3_500 = '1.85938e-14*ic_cap*ic_cap+1.81250e-14*ic_cap+5.30000e-13'
+ mcm4m2m1_cf_w_0_140_s_0_140 = '-9.84375e-14*ic_cap*ic_cap+-4.62500e-14*ic_cap+9.69000e-12'
+ mcm4m2m1_cf_w_0_140_s_0_175 = '-1.42813e-13*ic_cap*ic_cap+-7.12500e-14*ic_cap+1.22000e-11'
+ mcm4m2m1_cf_w_0_140_s_0_210 = '-1.90625e-13*ic_cap*ic_cap+-8.75000e-14*ic_cap+1.47000e-11'
+ mcm4m2m1_cf_w_0_140_s_0_280 = '-2.71875e-13*ic_cap*ic_cap+-1.37500e-13*ic_cap+1.93000e-11'
+ mcm4m2m1_cf_w_0_140_s_0_350 = '-3.46875e-13*ic_cap*ic_cap+-1.62500e-13*ic_cap+2.36000e-11'
+ mcm4m2m1_cf_w_0_140_s_0_420 = '-4.15625e-13*ic_cap*ic_cap+-2.12500e-13*ic_cap+2.76000e-11'
+ mcm4m2m1_cf_w_0_140_s_0_560 = '-4.96875e-13*ic_cap*ic_cap+-2.62500e-13*ic_cap+3.43000e-11'
+ mcm4m2m1_cf_w_0_140_s_0_840 = '-6.09375e-13*ic_cap*ic_cap+-3.12500e-13*ic_cap+4.42000e-11'
+ mcm4m2m1_cf_w_0_140_s_1_540 = '-6.46875e-13*ic_cap*ic_cap+-3.62500e-13*ic_cap+5.59000e-11'
+ mcm4m2m1_cf_w_0_140_s_3_500 = '-6.06250e-13*ic_cap*ic_cap+-3.25000e-13*ic_cap+6.18000e-11'
+ mcm4m2m1_cf_w_1_120_s_0_140 = '-9.65625e-14*ic_cap*ic_cap+-4.62500e-14*ic_cap+9.67000e-12'
+ mcm4m2m1_cf_w_1_120_s_0_175 = '-1.42500e-13*ic_cap*ic_cap+-7.00000e-14*ic_cap+1.22000e-11'
+ mcm4m2m1_cf_w_1_120_s_0_210 = '-1.90625e-13*ic_cap*ic_cap+-8.75000e-14*ic_cap+1.47000e-11'
+ mcm4m2m1_cf_w_1_120_s_0_280 = '-2.71875e-13*ic_cap*ic_cap+-1.37500e-13*ic_cap+1.93000e-11'
+ mcm4m2m1_cf_w_1_120_s_0_350 = '-3.43750e-13*ic_cap*ic_cap+-1.75000e-13*ic_cap+2.36000e-11'
+ mcm4m2m1_cf_w_1_120_s_0_420 = '-4.06250e-13*ic_cap*ic_cap+-2.00000e-13*ic_cap+2.76000e-11'
+ mcm4m2m1_cf_w_1_120_s_0_560 = '-5.03125e-13*ic_cap*ic_cap+-2.62500e-13*ic_cap+3.44000e-11'
+ mcm4m2m1_cf_w_1_120_s_0_840 = '-6.09375e-13*ic_cap*ic_cap+-3.12500e-13*ic_cap+4.46000e-11'
+ mcm4m2m1_cf_w_1_120_s_1_540 = '-6.46875e-13*ic_cap*ic_cap+-3.62500e-13*ic_cap+5.73000e-11'
+ mcm4m2m1_cf_w_1_120_s_3_500 = '-5.81250e-13*ic_cap*ic_cap+-3.25000e-13*ic_cap+6.42000e-11'
+ mcm4m2p1_ca_w_0_140_s_0_140 = '-4.84375e-07*ic_cap*ic_cap+-2.87500e-07*ic_cap+4.56000e-05'
+ mcm4m2p1_ca_w_0_140_s_0_175 = '-4.84375e-07*ic_cap*ic_cap+-2.87500e-07*ic_cap+4.56000e-05'
+ mcm4m2p1_ca_w_0_140_s_0_210 = '-4.84375e-07*ic_cap*ic_cap+-2.87500e-07*ic_cap+4.56000e-05'
+ mcm4m2p1_ca_w_0_140_s_0_280 = '-4.84375e-07*ic_cap*ic_cap+-2.87500e-07*ic_cap+4.56000e-05'
+ mcm4m2p1_ca_w_0_140_s_0_350 = '-4.84375e-07*ic_cap*ic_cap+-2.87500e-07*ic_cap+4.56000e-05'
+ mcm4m2p1_ca_w_0_140_s_0_420 = '-4.84375e-07*ic_cap*ic_cap+-2.87500e-07*ic_cap+4.56000e-05'
+ mcm4m2p1_ca_w_0_140_s_0_560 = '-4.84375e-07*ic_cap*ic_cap+-2.87500e-07*ic_cap+4.56000e-05'
+ mcm4m2p1_ca_w_0_140_s_0_840 = '-4.84375e-07*ic_cap*ic_cap+-2.87500e-07*ic_cap+4.56000e-05'
+ mcm4m2p1_ca_w_0_140_s_1_540 = '-4.84375e-07*ic_cap*ic_cap+-2.87500e-07*ic_cap+4.56000e-05'
+ mcm4m2p1_ca_w_0_140_s_3_500 = '-4.84375e-07*ic_cap*ic_cap+-2.87500e-07*ic_cap+4.56000e-05'
+ mcm4m2p1_ca_w_1_120_s_0_140 = '-4.84375e-07*ic_cap*ic_cap+-2.87500e-07*ic_cap+4.56000e-05'
+ mcm4m2p1_ca_w_1_120_s_0_175 = '-4.84375e-07*ic_cap*ic_cap+-2.87500e-07*ic_cap+4.56000e-05'
+ mcm4m2p1_ca_w_1_120_s_0_210 = '-4.84375e-07*ic_cap*ic_cap+-2.87500e-07*ic_cap+4.56000e-05'
+ mcm4m2p1_ca_w_1_120_s_0_280 = '-4.84375e-07*ic_cap*ic_cap+-2.87500e-07*ic_cap+4.56000e-05'
+ mcm4m2p1_ca_w_1_120_s_0_350 = '-4.84375e-07*ic_cap*ic_cap+-2.87500e-07*ic_cap+4.56000e-05'
+ mcm4m2p1_ca_w_1_120_s_0_420 = '-4.84375e-07*ic_cap*ic_cap+-2.87500e-07*ic_cap+4.56000e-05'
+ mcm4m2p1_ca_w_1_120_s_0_560 = '-4.84375e-07*ic_cap*ic_cap+-2.87500e-07*ic_cap+4.56000e-05'
+ mcm4m2p1_ca_w_1_120_s_0_840 = '-4.84375e-07*ic_cap*ic_cap+-2.87500e-07*ic_cap+4.56000e-05'
+ mcm4m2p1_ca_w_1_120_s_1_540 = '-4.84375e-07*ic_cap*ic_cap+-2.87500e-07*ic_cap+4.56000e-05'
+ mcm4m2p1_ca_w_1_120_s_3_500 = '-4.84375e-07*ic_cap*ic_cap+-2.87500e-07*ic_cap+4.56000e-05'
+ mcm4m2p1_cc_w_0_140_s_0_140 = '-9.28125e-13*ic_cap*ic_cap+-4.87500e-13*ic_cap+1.03000e-10'
+ mcm4m2p1_cc_w_0_140_s_0_175 = '-8.59375e-13*ic_cap*ic_cap+-5.87500e-13*ic_cap+1.01000e-10'
+ mcm4m2p1_cc_w_0_140_s_0_210 = '-7.37500e-13*ic_cap*ic_cap+-4.50000e-13*ic_cap+9.50000e-11'
+ mcm4m2p1_cc_w_0_140_s_0_280 = '-5.46875e-13*ic_cap*ic_cap+-3.87500e-13*ic_cap+8.37000e-11'
+ mcm4m2p1_cc_w_0_140_s_0_350 = '-4.34375e-13*ic_cap*ic_cap+-2.37500e-13*ic_cap+7.23000e-11'
+ mcm4m2p1_cc_w_0_140_s_0_420 = '-3.00000e-13*ic_cap*ic_cap+-2.25000e-13*ic_cap+6.22000e-11'
+ mcm4m2p1_cc_w_0_140_s_0_560 = '-1.59375e-13*ic_cap*ic_cap+-1.37500e-13*ic_cap+4.88000e-11'
+ mcm4m2p1_cc_w_0_140_s_0_840 = '-1.56250e-14*ic_cap*ic_cap+-1.25000e-14*ic_cap+3.29000e-11'
+ mcm4m2p1_cc_w_0_140_s_1_540 = '7.81250e-14*ic_cap*ic_cap+3.75000e-14*ic_cap+1.52000e-11'
+ mcm4m2p1_cc_w_0_140_s_3_500 = '5.65625e-14*ic_cap*ic_cap+3.87500e-14*ic_cap+2.39000e-12'
+ mcm4m2p1_cc_w_1_120_s_0_140 = '-7.18750e-13*ic_cap*ic_cap+-3.75000e-13*ic_cap+1.20000e-10'
+ mcm4m2p1_cc_w_1_120_s_0_175 = '-7.18750e-13*ic_cap*ic_cap+-3.75000e-13*ic_cap+1.17000e-10'
+ mcm4m2p1_cc_w_1_120_s_0_210 = '-5.87500e-13*ic_cap*ic_cap+-3.50000e-13*ic_cap+1.10000e-10'
+ mcm4m2p1_cc_w_1_120_s_0_280 = '-3.96875e-13*ic_cap*ic_cap+-2.87500e-13*ic_cap+9.55000e-11'
+ mcm4m2p1_cc_w_1_120_s_0_350 = '-2.81250e-13*ic_cap*ic_cap+-2.25000e-13*ic_cap+8.27000e-11'
+ mcm4m2p1_cc_w_1_120_s_0_420 = '-1.81250e-13*ic_cap*ic_cap+-1.25000e-13*ic_cap+7.18000e-11'
+ mcm4m2p1_cc_w_1_120_s_0_560 = '-4.68750e-14*ic_cap*ic_cap+-3.75000e-14*ic_cap+5.60000e-11'
+ mcm4m2p1_cc_w_1_120_s_0_840 = '6.87500e-14*ic_cap*ic_cap+5.00000e-14*ic_cap+3.79000e-11'
+ mcm4m2p1_cc_w_1_120_s_1_540 = '1.34375e-13*ic_cap*ic_cap+8.75000e-14*ic_cap+1.78000e-11'
+ mcm4m2p1_cc_w_1_120_s_3_500 = '7.81250e-14*ic_cap*ic_cap+5.50000e-14*ic_cap+2.83000e-12'
+ mcm4m2p1_cf_w_0_140_s_0_140 = '-3.75000e-15*ic_cap*ic_cap+-2.50000e-15*ic_cap+3.16000e-12'
+ mcm4m2p1_cf_w_0_140_s_0_175 = '-1.25000e-14*ic_cap*ic_cap+-7.50000e-15*ic_cap+3.94000e-12'
+ mcm4m2p1_cf_w_0_140_s_0_210 = '-1.90625e-14*ic_cap*ic_cap+-1.12500e-14*ic_cap+4.73000e-12'
+ mcm4m2p1_cf_w_0_140_s_0_280 = '-3.62500e-14*ic_cap*ic_cap+-2.25000e-14*ic_cap+6.26000e-12'
+ mcm4m2p1_cf_w_0_140_s_0_350 = '-5.18750e-14*ic_cap*ic_cap+-3.25000e-14*ic_cap+7.76000e-12'
+ mcm4m2p1_cf_w_0_140_s_0_420 = '-6.75000e-14*ic_cap*ic_cap+-4.00000e-14*ic_cap+9.29000e-12'
+ mcm4m2p1_cf_w_0_140_s_0_560 = '-9.68750e-14*ic_cap*ic_cap+-6.25000e-14*ic_cap+1.21000e-11'
+ mcm4m2p1_cf_w_0_140_s_0_840 = '-1.46875e-13*ic_cap*ic_cap+-8.75000e-14*ic_cap+1.72000e-11'
+ mcm4m2p1_cf_w_0_140_s_1_540 = '-2.28125e-13*ic_cap*ic_cap+-1.37500e-13*ic_cap+2.69000e-11'
+ mcm4m2p1_cf_w_0_140_s_3_500 = '-2.34375e-13*ic_cap*ic_cap+-1.62500e-13*ic_cap+3.75000e-11'
+ mcm4m2p1_cf_w_1_120_s_0_140 = '-5.31250e-15*ic_cap*ic_cap+-3.75000e-15*ic_cap+3.23000e-12'
+ mcm4m2p1_cf_w_1_120_s_0_175 = '-1.25000e-14*ic_cap*ic_cap+-1.00000e-14*ic_cap+4.00000e-12'
+ mcm4m2p1_cf_w_1_120_s_0_210 = '-2.03125e-14*ic_cap*ic_cap+-1.37500e-14*ic_cap+4.77000e-12'
+ mcm4m2p1_cf_w_1_120_s_0_280 = '-3.59375e-14*ic_cap*ic_cap+-2.12500e-14*ic_cap+6.31000e-12'
+ mcm4m2p1_cf_w_1_120_s_0_350 = '-5.21875e-14*ic_cap*ic_cap+-3.37500e-14*ic_cap+7.83000e-12'
+ mcm4m2p1_cf_w_1_120_s_0_420 = '-6.87500e-14*ic_cap*ic_cap+-4.50000e-14*ic_cap+9.33000e-12'
+ mcm4m2p1_cf_w_1_120_s_0_560 = '-9.68750e-14*ic_cap*ic_cap+-6.25000e-14*ic_cap+1.22000e-11'
+ mcm4m2p1_cf_w_1_120_s_0_840 = '-1.46875e-13*ic_cap*ic_cap+-8.75000e-14*ic_cap+1.75000e-11'
+ mcm4m2p1_cf_w_1_120_s_1_540 = '-2.28125e-13*ic_cap*ic_cap+-1.37500e-13*ic_cap+2.78000e-11'
+ mcm4m2p1_cf_w_1_120_s_3_500 = '-2.25000e-13*ic_cap*ic_cap+-1.50000e-13*ic_cap+3.97000e-11'
+ mcm4m3_ca_w_0_300_s_0_300 = '-1.72187e-06*ic_cap*ic_cap+-8.37500e-07*ic_cap+8.85000e-05'
+ mcm4m3_ca_w_0_300_s_0_360 = '-1.72187e-06*ic_cap*ic_cap+-8.37500e-07*ic_cap+8.85000e-05'
+ mcm4m3_ca_w_0_300_s_0_450 = '-1.72187e-06*ic_cap*ic_cap+-8.37500e-07*ic_cap+8.85000e-05'
+ mcm4m3_ca_w_0_300_s_0_600 = '-1.72187e-06*ic_cap*ic_cap+-8.37500e-07*ic_cap+8.85000e-05'
+ mcm4m3_ca_w_0_300_s_0_800 = '-1.72187e-06*ic_cap*ic_cap+-8.37500e-07*ic_cap+8.85000e-05'
+ mcm4m3_ca_w_0_300_s_1_000 = '-1.72187e-06*ic_cap*ic_cap+-8.37500e-07*ic_cap+8.85000e-05'
+ mcm4m3_ca_w_0_300_s_1_200 = '-1.72187e-06*ic_cap*ic_cap+-8.37500e-07*ic_cap+8.85000e-05'
+ mcm4m3_ca_w_0_300_s_2_100 = '-1.72187e-06*ic_cap*ic_cap+-8.37500e-07*ic_cap+8.85000e-05'
+ mcm4m3_ca_w_0_300_s_3_300 = '-1.72187e-06*ic_cap*ic_cap+-8.37500e-07*ic_cap+8.85000e-05'
+ mcm4m3_ca_w_0_300_s_9_000 = '-1.72187e-06*ic_cap*ic_cap+-8.37500e-07*ic_cap+8.85000e-05'
+ mcm4m3_ca_w_2_400_s_0_300 = '-1.72187e-06*ic_cap*ic_cap+-8.37500e-07*ic_cap+8.85000e-05'
+ mcm4m3_ca_w_2_400_s_0_360 = '-1.72187e-06*ic_cap*ic_cap+-8.37500e-07*ic_cap+8.85000e-05'
+ mcm4m3_ca_w_2_400_s_0_450 = '-1.72187e-06*ic_cap*ic_cap+-8.37500e-07*ic_cap+8.85000e-05'
+ mcm4m3_ca_w_2_400_s_0_600 = '-1.72187e-06*ic_cap*ic_cap+-8.37500e-07*ic_cap+8.85000e-05'
+ mcm4m3_ca_w_2_400_s_0_800 = '-1.72187e-06*ic_cap*ic_cap+-8.37500e-07*ic_cap+8.85000e-05'
+ mcm4m3_ca_w_2_400_s_1_000 = '-1.72187e-06*ic_cap*ic_cap+-8.37500e-07*ic_cap+8.85000e-05'
+ mcm4m3_ca_w_2_400_s_1_200 = '-1.72187e-06*ic_cap*ic_cap+-8.37500e-07*ic_cap+8.85000e-05'
+ mcm4m3_ca_w_2_400_s_2_100 = '-1.72187e-06*ic_cap*ic_cap+-8.37500e-07*ic_cap+8.85000e-05'
+ mcm4m3_ca_w_2_400_s_3_300 = '-1.72187e-06*ic_cap*ic_cap+-8.37500e-07*ic_cap+8.85000e-05'
+ mcm4m3_ca_w_2_400_s_9_000 = '-1.72187e-06*ic_cap*ic_cap+-8.37500e-07*ic_cap+8.85000e-05'
+ mcm4m3_cc_w_0_300_s_0_300 = '-6.15625e-13*ic_cap*ic_cap+-3.62500e-13*ic_cap+9.36000e-11'
+ mcm4m3_cc_w_0_300_s_0_360 = '-5.21875e-13*ic_cap*ic_cap+-3.12500e-13*ic_cap+8.61000e-11'
+ mcm4m3_cc_w_0_300_s_0_450 = '-4.18750e-13*ic_cap*ic_cap+-2.50000e-13*ic_cap+7.62000e-11'
+ mcm4m3_cc_w_0_300_s_0_600 = '-2.90625e-13*ic_cap*ic_cap+-1.87500e-13*ic_cap+6.30000e-11'
+ mcm4m3_cc_w_0_300_s_0_800 = '-1.75000e-13*ic_cap*ic_cap+-1.25000e-13*ic_cap+5.05000e-11'
+ mcm4m3_cc_w_0_300_s_1_000 = '-1.09375e-13*ic_cap*ic_cap+-8.75000e-14*ic_cap+4.13000e-11'
+ mcm4m3_cc_w_0_300_s_1_200 = '-7.18750e-14*ic_cap*ic_cap+-6.25000e-14*ic_cap+3.45000e-11'
+ mcm4m3_cc_w_0_300_s_2_100 = '-9.37500e-15*ic_cap*ic_cap+-1.25000e-14*ic_cap+1.80000e-11'
+ mcm4m3_cc_w_0_300_s_3_300 = '3.12500e-15*ic_cap*ic_cap+1.25000e-14*ic_cap+1.01000e-11'
+ mcm4m3_cc_w_0_300_s_9_000 = '4.68750e-15*ic_cap*ic_cap+6.25000e-15*ic_cap+1.90000e-12'
+ mcm4m3_cc_w_2_400_s_0_300 = '-5.93750e-13*ic_cap*ic_cap+-3.75000e-13*ic_cap+1.12000e-10'
+ mcm4m3_cc_w_2_400_s_0_360 = '-5.40625e-13*ic_cap*ic_cap+-3.12500e-13*ic_cap+1.04000e-10'
+ mcm4m3_cc_w_2_400_s_0_450 = '-4.25000e-13*ic_cap*ic_cap+-2.50000e-13*ic_cap+9.29000e-11'
+ mcm4m3_cc_w_2_400_s_0_600 = '-2.93750e-13*ic_cap*ic_cap+-1.75000e-13*ic_cap+7.84000e-11'
+ mcm4m3_cc_w_2_400_s_0_800 = '-1.84375e-13*ic_cap*ic_cap+-1.12500e-13*ic_cap+6.42000e-11'
+ mcm4m3_cc_w_2_400_s_1_000 = '-1.12500e-13*ic_cap*ic_cap+-7.50000e-14*ic_cap+5.38000e-11'
+ mcm4m3_cc_w_2_400_s_1_200 = '-7.50000e-14*ic_cap*ic_cap+-5.00000e-14*ic_cap+4.61000e-11'
+ mcm4m3_cc_w_2_400_s_2_100 = '-9.37500e-15*ic_cap*ic_cap+-1.25000e-14*ic_cap+2.75000e-11'
+ mcm4m3_cc_w_2_400_s_3_300 = '6.25000e-15*ic_cap*ic_cap+1.67000e-11'
+ mcm4m3_cc_w_2_400_s_9_000 = '9.37500e-15*ic_cap*ic_cap+3.95000e-12'
+ mcm4m3_cf_w_0_300_s_0_300 = '-1.46250e-13*ic_cap*ic_cap+-7.50000e-14*ic_cap+1.18000e-11'
+ mcm4m3_cf_w_0_300_s_0_360 = '-1.84375e-13*ic_cap*ic_cap+-8.75000e-14*ic_cap+1.39000e-11'
+ mcm4m3_cf_w_0_300_s_0_450 = '-2.25000e-13*ic_cap*ic_cap+-1.25000e-13*ic_cap+1.67000e-11'
+ mcm4m3_cf_w_0_300_s_0_600 = '-2.93750e-13*ic_cap*ic_cap+-1.50000e-13*ic_cap+2.11000e-11'
+ mcm4m3_cf_w_0_300_s_0_800 = '-3.46875e-13*ic_cap*ic_cap+-1.87500e-13*ic_cap+2.58000e-11'
+ mcm4m3_cf_w_0_300_s_1_000 = '-3.90625e-13*ic_cap*ic_cap+-2.12500e-13*ic_cap+2.99000e-11'
+ mcm4m3_cf_w_0_300_s_1_200 = '-4.21875e-13*ic_cap*ic_cap+-2.37500e-13*ic_cap+3.34000e-11'
+ mcm4m3_cf_w_0_300_s_2_100 = '-4.87500e-13*ic_cap*ic_cap+-2.75000e-13*ic_cap+4.46000e-11'
+ mcm4m3_cf_w_0_300_s_3_300 = '-5.03125e-13*ic_cap*ic_cap+-2.87500e-13*ic_cap+5.12000e-11'
+ mcm4m3_cf_w_0_300_s_9_000 = '-5.09375e-13*ic_cap*ic_cap+-2.87500e-13*ic_cap+5.91000e-11'
+ mcm4m3_cf_w_2_400_s_0_300 = '-1.45000e-13*ic_cap*ic_cap+-7.50000e-14*ic_cap+1.18000e-11'
+ mcm4m3_cf_w_2_400_s_0_360 = '-1.84375e-13*ic_cap*ic_cap+-8.75000e-14*ic_cap+1.39000e-11'
+ mcm4m3_cf_w_2_400_s_0_450 = '-2.31250e-13*ic_cap*ic_cap+-1.25000e-13*ic_cap+1.68000e-11'
+ mcm4m3_cf_w_2_400_s_0_600 = '-2.87500e-13*ic_cap*ic_cap+-1.50000e-13*ic_cap+2.10000e-11'
+ mcm4m3_cf_w_2_400_s_0_800 = '-3.46875e-13*ic_cap*ic_cap+-1.87500e-13*ic_cap+2.59000e-11'
+ mcm4m3_cf_w_2_400_s_1_000 = '-3.90625e-13*ic_cap*ic_cap+-2.12500e-13*ic_cap+3.00000e-11'
+ mcm4m3_cf_w_2_400_s_1_200 = '-4.15625e-13*ic_cap*ic_cap+-2.37500e-13*ic_cap+3.35000e-11'
+ mcm4m3_cf_w_2_400_s_2_100 = '-4.81250e-13*ic_cap*ic_cap+-2.75000e-13*ic_cap+4.46000e-11'
+ mcm4m3_cf_w_2_400_s_3_300 = '-5.06250e-13*ic_cap*ic_cap+-3.00000e-13*ic_cap+5.31000e-11'
+ mcm4m3_cf_w_2_400_s_9_000 = '-5.09375e-13*ic_cap*ic_cap+-2.87500e-13*ic_cap+6.50000e-11'
+ mcm4m3d_ca_w_0_300_s_0_300 = '-1.87812e-06*ic_cap*ic_cap+-9.37500e-07*ic_cap+1.03000e-04'
+ mcm4m3d_ca_w_0_300_s_0_360 = '-1.87812e-06*ic_cap*ic_cap+-9.37500e-07*ic_cap+1.03000e-04'
+ mcm4m3d_ca_w_0_300_s_0_450 = '-1.87812e-06*ic_cap*ic_cap+-9.37500e-07*ic_cap+1.03000e-04'
+ mcm4m3d_ca_w_0_300_s_0_600 = '-1.87812e-06*ic_cap*ic_cap+-9.37500e-07*ic_cap+1.03000e-04'
+ mcm4m3d_ca_w_0_300_s_0_800 = '-1.87812e-06*ic_cap*ic_cap+-9.37500e-07*ic_cap+1.03000e-04'
+ mcm4m3d_ca_w_0_300_s_1_000 = '-1.87812e-06*ic_cap*ic_cap+-9.37500e-07*ic_cap+1.03000e-04'
+ mcm4m3d_ca_w_0_300_s_1_200 = '-1.87812e-06*ic_cap*ic_cap+-9.37500e-07*ic_cap+1.03000e-04'
+ mcm4m3d_ca_w_0_300_s_2_100 = '-1.87812e-06*ic_cap*ic_cap+-9.37500e-07*ic_cap+1.03000e-04'
+ mcm4m3d_ca_w_0_300_s_3_300 = '-1.87812e-06*ic_cap*ic_cap+-9.37500e-07*ic_cap+1.03000e-04'
+ mcm4m3d_ca_w_0_300_s_9_000 = '-1.87812e-06*ic_cap*ic_cap+-9.37500e-07*ic_cap+1.03000e-04'
+ mcm4m3d_ca_w_2_400_s_0_300 = '-1.87812e-06*ic_cap*ic_cap+-9.37500e-07*ic_cap+1.03000e-04'
+ mcm4m3d_ca_w_2_400_s_0_360 = '-1.87812e-06*ic_cap*ic_cap+-9.37500e-07*ic_cap+1.03000e-04'
+ mcm4m3d_ca_w_2_400_s_0_450 = '-1.87812e-06*ic_cap*ic_cap+-9.37500e-07*ic_cap+1.03000e-04'
+ mcm4m3d_ca_w_2_400_s_0_600 = '-1.87812e-06*ic_cap*ic_cap+-9.37500e-07*ic_cap+1.03000e-04'
+ mcm4m3d_ca_w_2_400_s_0_800 = '-1.87812e-06*ic_cap*ic_cap+-9.37500e-07*ic_cap+1.03000e-04'
+ mcm4m3d_ca_w_2_400_s_1_000 = '-1.87812e-06*ic_cap*ic_cap+-9.37500e-07*ic_cap+1.03000e-04'
+ mcm4m3d_ca_w_2_400_s_1_200 = '-1.87812e-06*ic_cap*ic_cap+-9.37500e-07*ic_cap+1.03000e-04'
+ mcm4m3d_ca_w_2_400_s_2_100 = '-1.87812e-06*ic_cap*ic_cap+-9.37500e-07*ic_cap+1.03000e-04'
+ mcm4m3d_ca_w_2_400_s_3_300 = '-1.87812e-06*ic_cap*ic_cap+-9.37500e-07*ic_cap+1.03000e-04'
+ mcm4m3d_ca_w_2_400_s_9_000 = '-1.87812e-06*ic_cap*ic_cap+-9.37500e-07*ic_cap+1.03000e-04'
+ mcm4m3d_cc_w_0_300_s_0_300 = '-5.56250e-13*ic_cap*ic_cap+-3.25000e-13*ic_cap+9.03000e-11'
+ mcm4m3d_cc_w_0_300_s_0_360 = '-4.90625e-13*ic_cap*ic_cap+-3.12500e-13*ic_cap+8.26000e-11'
+ mcm4m3d_cc_w_0_300_s_0_450 = '-3.37500e-13*ic_cap*ic_cap+-2.25000e-13*ic_cap+7.16000e-11'
+ mcm4m3d_cc_w_0_300_s_0_600 = '-2.18750e-13*ic_cap*ic_cap+-1.25000e-13*ic_cap+5.79000e-11'
+ mcm4m3d_cc_w_0_300_s_0_800 = '-9.68750e-14*ic_cap*ic_cap+-6.25000e-14*ic_cap+4.41000e-11'
+ mcm4m3d_cc_w_0_300_s_1_000 = '-3.12500e-14*ic_cap*ic_cap+-5.00000e-14*ic_cap+3.41000e-11'
+ mcm4m3d_cc_w_0_300_s_1_200 = '1.25000e-14*ic_cap*ic_cap+2.68000e-11'
+ mcm4m3d_cc_w_0_300_s_2_100 = '6.56250e-14*ic_cap*ic_cap+3.75000e-14*ic_cap+1.03000e-11'
+ mcm4m3d_cc_w_0_300_s_3_300 = '4.96875e-14*ic_cap*ic_cap+3.62500e-14*ic_cap+3.34000e-12'
+ mcm4m3d_cc_w_0_300_s_9_000 = '3.43750e-15*ic_cap*ic_cap+7.50000e-15*ic_cap+3.00000e-14'
+ mcm4m3d_cc_w_2_400_s_0_300 = '-4.68750e-13*ic_cap*ic_cap+-2.75000e-13*ic_cap+9.75000e-11'
+ mcm4m3d_cc_w_2_400_s_0_360 = '-3.90625e-13*ic_cap*ic_cap+-2.12500e-13*ic_cap+8.91000e-11'
+ mcm4m3d_cc_w_2_400_s_0_450 = '-2.53125e-13*ic_cap*ic_cap+-1.62500e-13*ic_cap+7.76000e-11'
+ mcm4m3d_cc_w_2_400_s_0_600 = '-1.25000e-13*ic_cap*ic_cap+-7.50000e-14*ic_cap+6.27000e-11'
+ mcm4m3d_cc_w_2_400_s_0_800 = '-2.50000e-14*ic_cap*ic_cap+-2.50000e-14*ic_cap+4.80000e-11'
+ mcm4m3d_cc_w_2_400_s_1_000 = '4.06250e-14*ic_cap*ic_cap+1.25000e-14*ic_cap+3.73000e-11'
+ mcm4m3d_cc_w_2_400_s_1_200 = '7.18750e-14*ic_cap*ic_cap+3.75000e-14*ic_cap+2.95000e-11'
+ mcm4m3d_cc_w_2_400_s_2_100 = '1.06250e-13*ic_cap*ic_cap+7.50000e-14*ic_cap+1.18000e-11'
+ mcm4m3d_cc_w_2_400_s_3_300 = '6.96875e-14*ic_cap*ic_cap+4.87500e-14*ic_cap+4.00000e-12'
+ mcm4m3d_cc_w_2_400_s_9_000 = '5.00000e-15*ic_cap*ic_cap+2.50000e-15*ic_cap+3.50000e-14'
+ mcm4m3d_cf_w_0_300_s_0_300 = '-1.34375e-13*ic_cap*ic_cap+-6.25000e-14*ic_cap+1.30000e-11'
+ mcm4m3d_cf_w_0_300_s_0_360 = '-1.71875e-13*ic_cap*ic_cap+-8.75000e-14*ic_cap+1.54000e-11'
+ mcm4m3d_cf_w_0_300_s_0_450 = '-2.15625e-13*ic_cap*ic_cap+-1.12500e-13*ic_cap+1.87000e-11'
+ mcm4m3d_cf_w_0_300_s_0_600 = '-2.81250e-13*ic_cap*ic_cap+-1.50000e-13*ic_cap+2.38000e-11'
+ mcm4m3d_cf_w_0_300_s_0_800 = '-3.46875e-13*ic_cap*ic_cap+-1.87500e-13*ic_cap+2.96000e-11'
+ mcm4m3d_cf_w_0_300_s_1_000 = '-4.00000e-13*ic_cap*ic_cap+-2.25000e-13*ic_cap+3.47000e-11'
+ mcm4m3d_cf_w_0_300_s_1_200 = '-4.31250e-13*ic_cap*ic_cap+-2.50000e-13*ic_cap+3.88000e-11'
+ mcm4m3d_cf_w_0_300_s_2_100 = '-4.90625e-13*ic_cap*ic_cap+-2.87500e-13*ic_cap+5.07000e-11'
+ mcm4m3d_cf_w_0_300_s_3_300 = '-4.90625e-13*ic_cap*ic_cap+-2.87500e-13*ic_cap+5.69000e-11'
+ mcm4m3d_cf_w_0_300_s_9_000 = '-4.40625e-13*ic_cap*ic_cap+-2.62500e-13*ic_cap+6.01000e-11'
+ mcm4m3d_cf_w_2_400_s_0_300 = '-1.34375e-13*ic_cap*ic_cap+-6.25000e-14*ic_cap+1.31000e-11'
+ mcm4m3d_cf_w_2_400_s_0_360 = '-1.65625e-13*ic_cap*ic_cap+-8.75000e-14*ic_cap+1.54000e-11'
+ mcm4m3d_cf_w_2_400_s_0_450 = '-2.15625e-13*ic_cap*ic_cap+-1.12500e-13*ic_cap+1.88000e-11'
+ mcm4m3d_cf_w_2_400_s_0_600 = '-2.81250e-13*ic_cap*ic_cap+-1.50000e-13*ic_cap+2.39000e-11'
+ mcm4m3d_cf_w_2_400_s_0_800 = '-3.46875e-13*ic_cap*ic_cap+-1.87500e-13*ic_cap+2.98000e-11'
+ mcm4m3d_cf_w_2_400_s_1_000 = '-3.96875e-13*ic_cap*ic_cap+-2.12500e-13*ic_cap+3.49000e-11'
+ mcm4m3d_cf_w_2_400_s_1_200 = '-4.25000e-13*ic_cap*ic_cap+-2.50000e-13*ic_cap+3.91000e-11'
+ mcm4m3d_cf_w_2_400_s_2_100 = '-4.78125e-13*ic_cap*ic_cap+-2.87500e-13*ic_cap+5.14000e-11'
+ mcm4m3d_cf_w_2_400_s_3_300 = '-4.68750e-13*ic_cap*ic_cap+-2.75000e-13*ic_cap+5.84000e-11'
+ mcm4m3d_cf_w_2_400_s_9_000 = '-4.03125e-13*ic_cap*ic_cap+-2.37500e-13*ic_cap+6.22000e-11'
+ mcm4m3f_ca_w_0_300_s_0_300 = '-1.84375e-06*ic_cap*ic_cap+-9.25000e-07*ic_cap+1.01000e-04'
+ mcm4m3f_ca_w_0_300_s_0_360 = '-1.84375e-06*ic_cap*ic_cap+-9.25000e-07*ic_cap+1.01000e-04'
+ mcm4m3f_ca_w_0_300_s_0_450 = '-1.84375e-06*ic_cap*ic_cap+-9.25000e-07*ic_cap+1.01000e-04'
+ mcm4m3f_ca_w_0_300_s_0_600 = '-1.84375e-06*ic_cap*ic_cap+-9.25000e-07*ic_cap+1.01000e-04'
+ mcm4m3f_ca_w_0_300_s_0_800 = '-1.84375e-06*ic_cap*ic_cap+-9.25000e-07*ic_cap+1.01000e-04'
+ mcm4m3f_ca_w_0_300_s_1_000 = '-1.84375e-06*ic_cap*ic_cap+-9.25000e-07*ic_cap+1.01000e-04'
+ mcm4m3f_ca_w_0_300_s_1_200 = '-1.84375e-06*ic_cap*ic_cap+-9.25000e-07*ic_cap+1.01000e-04'
+ mcm4m3f_ca_w_0_300_s_2_100 = '-1.84375e-06*ic_cap*ic_cap+-9.25000e-07*ic_cap+1.01000e-04'
+ mcm4m3f_ca_w_0_300_s_3_300 = '-1.84375e-06*ic_cap*ic_cap+-9.25000e-07*ic_cap+1.01000e-04'
+ mcm4m3f_ca_w_0_300_s_9_000 = '-1.84375e-06*ic_cap*ic_cap+-9.25000e-07*ic_cap+1.01000e-04'
+ mcm4m3f_ca_w_2_400_s_0_300 = '-1.84375e-06*ic_cap*ic_cap+-9.25000e-07*ic_cap+1.01000e-04'
+ mcm4m3f_ca_w_2_400_s_0_360 = '-1.84375e-06*ic_cap*ic_cap+-9.25000e-07*ic_cap+1.01000e-04'
+ mcm4m3f_ca_w_2_400_s_0_450 = '-1.84375e-06*ic_cap*ic_cap+-9.25000e-07*ic_cap+1.01000e-04'
+ mcm4m3f_ca_w_2_400_s_0_600 = '-1.84375e-06*ic_cap*ic_cap+-9.25000e-07*ic_cap+1.01000e-04'
+ mcm4m3f_ca_w_2_400_s_0_800 = '-1.84375e-06*ic_cap*ic_cap+-9.25000e-07*ic_cap+1.01000e-04'
+ mcm4m3f_ca_w_2_400_s_1_000 = '-1.84375e-06*ic_cap*ic_cap+-9.25000e-07*ic_cap+1.01000e-04'
+ mcm4m3f_ca_w_2_400_s_1_200 = '-1.84375e-06*ic_cap*ic_cap+-9.25000e-07*ic_cap+1.01000e-04'
+ mcm4m3f_ca_w_2_400_s_2_100 = '-1.84375e-06*ic_cap*ic_cap+-9.25000e-07*ic_cap+1.01000e-04'
+ mcm4m3f_ca_w_2_400_s_3_300 = '-1.84375e-06*ic_cap*ic_cap+-9.25000e-07*ic_cap+1.01000e-04'
+ mcm4m3f_ca_w_2_400_s_9_000 = '-1.84375e-06*ic_cap*ic_cap+-9.25000e-07*ic_cap+1.01000e-04'
+ mcm4m3f_cc_w_0_300_s_0_300 = '-5.59375e-13*ic_cap*ic_cap+-3.37500e-13*ic_cap+9.07000e-11'
+ mcm4m3f_cc_w_0_300_s_0_360 = '-5.00000e-13*ic_cap*ic_cap+-2.75000e-13*ic_cap+8.30000e-11'
+ mcm4m3f_cc_w_0_300_s_0_450 = '-3.37500e-13*ic_cap*ic_cap+-2.50000e-13*ic_cap+7.20000e-11'
+ mcm4m3f_cc_w_0_300_s_0_600 = '-2.25000e-13*ic_cap*ic_cap+-1.25000e-13*ic_cap+5.84000e-11'
+ mcm4m3f_cc_w_0_300_s_0_800 = '-9.37500e-14*ic_cap*ic_cap+-7.50000e-14*ic_cap+4.47000e-11'
+ mcm4m3f_cc_w_0_300_s_1_000 = '-2.50000e-14*ic_cap*ic_cap+-5.00000e-14*ic_cap+3.47000e-11'
+ mcm4m3f_cc_w_0_300_s_1_200 = '2.18750e-14*ic_cap*ic_cap+-1.25000e-14*ic_cap+2.74000e-11'
+ mcm4m3f_cc_w_0_300_s_2_100 = '6.56250e-14*ic_cap*ic_cap+3.75000e-14*ic_cap+1.09000e-11'
+ mcm4m3f_cc_w_0_300_s_3_300 = '5.50000e-14*ic_cap*ic_cap+3.25000e-14*ic_cap+3.74000e-12'
+ mcm4m3f_cc_w_0_300_s_9_000 = '1.09375e-15*ic_cap*ic_cap+5.62500e-15*ic_cap+1.10000e-13'
+ mcm4m3f_cc_w_2_400_s_0_300 = '-4.65625e-13*ic_cap*ic_cap+-2.87500e-13*ic_cap+9.86000e-11'
+ mcm4m3f_cc_w_2_400_s_0_360 = '-3.90625e-13*ic_cap*ic_cap+-2.12500e-13*ic_cap+9.03000e-11'
+ mcm4m3f_cc_w_2_400_s_0_450 = '-2.65625e-13*ic_cap*ic_cap+-1.62500e-13*ic_cap+7.89000e-11'
+ mcm4m3f_cc_w_2_400_s_0_600 = '-1.25000e-13*ic_cap*ic_cap+-7.50000e-14*ic_cap+6.39000e-11'
+ mcm4m3f_cc_w_2_400_s_0_800 = '-2.50000e-14*ic_cap*ic_cap+-2.50000e-14*ic_cap+4.92000e-11'
+ mcm4m3f_cc_w_2_400_s_1_000 = '4.37500e-14*ic_cap*ic_cap+3.85000e-11'
+ mcm4m3f_cc_w_2_400_s_1_200 = '7.18750e-14*ic_cap*ic_cap+3.75000e-14*ic_cap+3.07000e-11'
+ mcm4m3f_cc_w_2_400_s_2_100 = '1.12500e-13*ic_cap*ic_cap+7.50000e-14*ic_cap+1.27000e-11'
+ mcm4m3f_cc_w_2_400_s_3_300 = '8.21875e-14*ic_cap*ic_cap+5.37500e-14*ic_cap+4.61000e-12'
+ mcm4m3f_cc_w_2_400_s_9_000 = '-1.56250e-16*ic_cap*ic_cap+6.25000e-16*ic_cap+1.40000e-13'
+ mcm4m3f_cf_w_0_300_s_0_300 = '-1.37500e-13*ic_cap*ic_cap+-7.50000e-14*ic_cap+1.28000e-11'
+ mcm4m3f_cf_w_0_300_s_0_360 = '-1.71875e-13*ic_cap*ic_cap+-8.75000e-14*ic_cap+1.51000e-11'
+ mcm4m3f_cf_w_0_300_s_0_450 = '-2.15625e-13*ic_cap*ic_cap+-1.12500e-13*ic_cap+1.84000e-11'
+ mcm4m3f_cf_w_0_300_s_0_600 = '-2.81250e-13*ic_cap*ic_cap+-1.50000e-13*ic_cap+2.34000e-11'
+ mcm4m3f_cf_w_0_300_s_0_800 = '-3.46875e-13*ic_cap*ic_cap+-1.87500e-13*ic_cap+2.91000e-11'
+ mcm4m3f_cf_w_0_300_s_1_000 = '-3.93750e-13*ic_cap*ic_cap+-2.25000e-13*ic_cap+3.40000e-11'
+ mcm4m3f_cf_w_0_300_s_1_200 = '-4.31250e-13*ic_cap*ic_cap+-2.50000e-13*ic_cap+3.81000e-11'
+ mcm4m3f_cf_w_0_300_s_2_100 = '-4.87500e-13*ic_cap*ic_cap+-2.75000e-13*ic_cap+4.98000e-11'
+ mcm4m3f_cf_w_0_300_s_3_300 = '-4.90625e-13*ic_cap*ic_cap+-2.87500e-13*ic_cap+5.62000e-11'
+ mcm4m3f_cf_w_0_300_s_9_000 = '-4.34375e-13*ic_cap*ic_cap+-2.62500e-13*ic_cap+5.97000e-11'
+ mcm4m3f_cf_w_2_400_s_0_300 = '-1.37500e-13*ic_cap*ic_cap+-7.50000e-14*ic_cap+1.29000e-11'
+ mcm4m3f_cf_w_2_400_s_0_360 = '-1.71875e-13*ic_cap*ic_cap+-8.75000e-14*ic_cap+1.52000e-11'
+ mcm4m3f_cf_w_2_400_s_0_450 = '-2.09375e-13*ic_cap*ic_cap+-1.12500e-13*ic_cap+1.84000e-11'
+ mcm4m3f_cf_w_2_400_s_0_600 = '-2.75000e-13*ic_cap*ic_cap+-1.50000e-13*ic_cap+2.34000e-11'
+ mcm4m3f_cf_w_2_400_s_0_800 = '-3.40625e-13*ic_cap*ic_cap+-1.87500e-13*ic_cap+2.92000e-11'
+ mcm4m3f_cf_w_2_400_s_1_000 = '-3.93750e-13*ic_cap*ic_cap+-2.25000e-13*ic_cap+3.42000e-11'
+ mcm4m3f_cf_w_2_400_s_1_200 = '-4.21875e-13*ic_cap*ic_cap+-2.37500e-13*ic_cap+3.83000e-11'
+ mcm4m3f_cf_w_2_400_s_2_100 = '-4.78125e-13*ic_cap*ic_cap+-2.87500e-13*ic_cap+5.06000e-11'
+ mcm4m3f_cf_w_2_400_s_3_300 = '-4.71875e-13*ic_cap*ic_cap+-2.87500e-13*ic_cap+5.78000e-11'
+ mcm4m3f_cf_w_2_400_s_9_000 = '-3.96875e-13*ic_cap*ic_cap+-2.37500e-13*ic_cap+6.21000e-11'
+ mcm4m3l1_ca_w_0_300_s_0_300 = '-1.95000e-06*ic_cap*ic_cap+-9.75000e-07*ic_cap+1.09000e-04'
+ mcm4m3l1_ca_w_0_300_s_0_360 = '-1.95000e-06*ic_cap*ic_cap+-9.75000e-07*ic_cap+1.09000e-04'
+ mcm4m3l1_ca_w_0_300_s_0_450 = '-1.95000e-06*ic_cap*ic_cap+-9.75000e-07*ic_cap+1.09000e-04'
+ mcm4m3l1_ca_w_0_300_s_0_600 = '-1.95000e-06*ic_cap*ic_cap+-9.75000e-07*ic_cap+1.09000e-04'
+ mcm4m3l1_ca_w_0_300_s_0_800 = '-1.95000e-06*ic_cap*ic_cap+-9.75000e-07*ic_cap+1.09000e-04'
+ mcm4m3l1_ca_w_0_300_s_1_000 = '-1.95000e-06*ic_cap*ic_cap+-9.75000e-07*ic_cap+1.09000e-04'
+ mcm4m3l1_ca_w_0_300_s_1_200 = '-1.95000e-06*ic_cap*ic_cap+-9.75000e-07*ic_cap+1.09000e-04'
+ mcm4m3l1_ca_w_0_300_s_2_100 = '-1.95000e-06*ic_cap*ic_cap+-9.75000e-07*ic_cap+1.09000e-04'
+ mcm4m3l1_ca_w_0_300_s_3_300 = '-1.95000e-06*ic_cap*ic_cap+-9.75000e-07*ic_cap+1.09000e-04'
+ mcm4m3l1_ca_w_0_300_s_9_000 = '-1.95000e-06*ic_cap*ic_cap+-9.75000e-07*ic_cap+1.09000e-04'
+ mcm4m3l1_ca_w_2_400_s_0_300 = '-1.95000e-06*ic_cap*ic_cap+-9.75000e-07*ic_cap+1.09000e-04'
+ mcm4m3l1_ca_w_2_400_s_0_360 = '-1.95000e-06*ic_cap*ic_cap+-9.75000e-07*ic_cap+1.09000e-04'
+ mcm4m3l1_ca_w_2_400_s_0_450 = '-1.95000e-06*ic_cap*ic_cap+-9.75000e-07*ic_cap+1.09000e-04'
+ mcm4m3l1_ca_w_2_400_s_0_600 = '-1.95000e-06*ic_cap*ic_cap+-9.75000e-07*ic_cap+1.09000e-04'
+ mcm4m3l1_ca_w_2_400_s_0_800 = '-1.95000e-06*ic_cap*ic_cap+-9.75000e-07*ic_cap+1.09000e-04'
+ mcm4m3l1_ca_w_2_400_s_1_000 = '-1.95000e-06*ic_cap*ic_cap+-9.75000e-07*ic_cap+1.09000e-04'
+ mcm4m3l1_ca_w_2_400_s_1_200 = '-1.95000e-06*ic_cap*ic_cap+-9.75000e-07*ic_cap+1.09000e-04'
+ mcm4m3l1_ca_w_2_400_s_2_100 = '-1.95000e-06*ic_cap*ic_cap+-9.75000e-07*ic_cap+1.09000e-04'
+ mcm4m3l1_ca_w_2_400_s_3_300 = '-1.95000e-06*ic_cap*ic_cap+-9.75000e-07*ic_cap+1.09000e-04'
+ mcm4m3l1_ca_w_2_400_s_9_000 = '-1.95000e-06*ic_cap*ic_cap+-9.75000e-07*ic_cap+1.09000e-04'
+ mcm4m3l1_cc_w_0_300_s_0_300 = '-5.50000e-13*ic_cap*ic_cap+-2.75000e-13*ic_cap+8.88000e-11'
+ mcm4m3l1_cc_w_0_300_s_0_360 = '-4.59375e-13*ic_cap*ic_cap+-2.87500e-13*ic_cap+8.08000e-11'
+ mcm4m3l1_cc_w_0_300_s_0_450 = '-3.34375e-13*ic_cap*ic_cap+-2.12500e-13*ic_cap+7.02000e-11'
+ mcm4m3l1_cc_w_0_300_s_0_600 = '-1.93750e-13*ic_cap*ic_cap+-1.00000e-13*ic_cap+5.59000e-11'
+ mcm4m3l1_cc_w_0_300_s_0_800 = '-7.50000e-14*ic_cap*ic_cap+-5.00000e-14*ic_cap+4.19000e-11'
+ mcm4m3l1_cc_w_0_300_s_1_000 = '4.03897e-28*ic_cap*ic_cap+-2.50000e-14*ic_cap+3.17000e-11'
+ mcm4m3l1_cc_w_0_300_s_1_200 = '4.37500e-14*ic_cap*ic_cap+2.50000e-14*ic_cap+2.43000e-11'
+ mcm4m3l1_cc_w_0_300_s_2_100 = '7.62500e-14*ic_cap*ic_cap+4.25000e-14*ic_cap+8.33000e-12'
+ mcm4m3l1_cc_w_0_300_s_3_300 = '4.65625e-14*ic_cap*ic_cap+3.62500e-14*ic_cap+2.24000e-12'
+ mcm4m3l1_cc_w_0_300_s_9_000 = '3.12500e-15*ic_cap*ic_cap+-2.50000e-15*ic_cap+5.00000e-15'
+ mcm4m3l1_cc_w_2_400_s_0_300 = '-4.56250e-13*ic_cap*ic_cap+-2.50000e-13*ic_cap+9.39000e-11'
+ mcm4m3l1_cc_w_2_400_s_0_360 = '-3.53125e-13*ic_cap*ic_cap+-1.87500e-13*ic_cap+8.52000e-11'
+ mcm4m3l1_cc_w_2_400_s_0_450 = '-2.37500e-13*ic_cap*ic_cap+-1.25000e-13*ic_cap+7.39000e-11'
+ mcm4m3l1_cc_w_2_400_s_0_600 = '-1.18750e-13*ic_cap*ic_cap+-5.00000e-14*ic_cap+5.91000e-11'
+ mcm4m3l1_cc_w_2_400_s_0_800 = '-1.25000e-14*ic_cap*ic_cap+4.43000e-11'
+ mcm4m3l1_cc_w_2_400_s_1_000 = '5.00000e-14*ic_cap*ic_cap+2.50000e-14*ic_cap+3.37000e-11'
+ mcm4m3l1_cc_w_2_400_s_1_200 = '8.12500e-14*ic_cap*ic_cap+5.00000e-14*ic_cap+2.60000e-11'
+ mcm4m3l1_cc_w_2_400_s_2_100 = '1.00625e-13*ic_cap*ic_cap+7.50000e-14*ic_cap+9.09000e-12'
+ mcm4m3l1_cc_w_2_400_s_3_300 = '5.68750e-14*ic_cap*ic_cap+4.50000e-14*ic_cap+2.50000e-12'
+ mcm4m3l1_cc_w_2_400_s_9_000 = '3.90625e-15*ic_cap*ic_cap+1.87500e-15*ic_cap'
+ mcm4m3l1_cf_w_0_300_s_0_300 = '-1.43750e-13*ic_cap*ic_cap+-7.50000e-14*ic_cap+1.39000e-11'
+ mcm4m3l1_cf_w_0_300_s_0_360 = '-1.78125e-13*ic_cap*ic_cap+-8.75000e-14*ic_cap+1.64000e-11'
+ mcm4m3l1_cf_w_0_300_s_0_450 = '-2.28125e-13*ic_cap*ic_cap+-1.12500e-13*ic_cap+2.00000e-11'
+ mcm4m3l1_cf_w_0_300_s_0_600 = '-2.93750e-13*ic_cap*ic_cap+-1.50000e-13*ic_cap+2.54000e-11'
+ mcm4m3l1_cf_w_0_300_s_0_800 = '-3.65625e-13*ic_cap*ic_cap+-2.12500e-13*ic_cap+3.17000e-11'
+ mcm4m3l1_cf_w_0_300_s_1_000 = '-4.18750e-13*ic_cap*ic_cap+-2.25000e-13*ic_cap+3.70000e-11'
+ mcm4m3l1_cf_w_0_300_s_1_200 = '-4.50000e-13*ic_cap*ic_cap+-2.75000e-13*ic_cap+4.14000e-11'
+ mcm4m3l1_cf_w_0_300_s_2_100 = '-5.15625e-13*ic_cap*ic_cap+-3.12500e-13*ic_cap+5.35000e-11'
+ mcm4m3l1_cf_w_0_300_s_3_300 = '-4.90625e-13*ic_cap*ic_cap+-2.87500e-13*ic_cap+5.90000e-11'
+ mcm4m3l1_cf_w_0_300_s_9_000 = '-4.53125e-13*ic_cap*ic_cap+-2.62500e-13*ic_cap+6.13000e-11'
+ mcm4m3l1_cf_w_2_400_s_0_300 = '-1.34375e-13*ic_cap*ic_cap+-6.25000e-14*ic_cap+1.39000e-11'
+ mcm4m3l1_cf_w_2_400_s_0_360 = '-1.71875e-13*ic_cap*ic_cap+-8.75000e-14*ic_cap+1.64000e-11'
+ mcm4m3l1_cf_w_2_400_s_0_450 = '-2.18750e-13*ic_cap*ic_cap+-1.25000e-13*ic_cap+2.00000e-11'
+ mcm4m3l1_cf_w_2_400_s_0_600 = '-2.90625e-13*ic_cap*ic_cap+-1.62500e-13*ic_cap+2.55000e-11'
+ mcm4m3l1_cf_w_2_400_s_0_800 = '-3.65625e-13*ic_cap*ic_cap+-2.12500e-13*ic_cap+3.19000e-11'
+ mcm4m3l1_cf_w_2_400_s_1_000 = '-4.15625e-13*ic_cap*ic_cap+-2.37500e-13*ic_cap+3.73000e-11'
+ mcm4m3l1_cf_w_2_400_s_1_200 = '-4.46875e-13*ic_cap*ic_cap+-2.62500e-13*ic_cap+4.17000e-11'
+ mcm4m3l1_cf_w_2_400_s_2_100 = '-5.00000e-13*ic_cap*ic_cap+-3.00000e-13*ic_cap+5.42000e-11'
+ mcm4m3l1_cf_w_2_400_s_3_300 = '-4.71875e-13*ic_cap*ic_cap+-2.87500e-13*ic_cap+6.03000e-11'
+ mcm4m3l1_cf_w_2_400_s_9_000 = '-4.12500e-13*ic_cap*ic_cap+-2.50000e-13*ic_cap+6.27000e-11'
+ mcm4m3m1_ca_w_0_300_s_0_300 = '-2.08750e-06*ic_cap*ic_cap+-1.07500e-06*ic_cap+1.21000e-04'
+ mcm4m3m1_ca_w_0_300_s_0_360 = '-2.08750e-06*ic_cap*ic_cap+-1.07500e-06*ic_cap+1.21000e-04'
+ mcm4m3m1_ca_w_0_300_s_0_450 = '-2.08750e-06*ic_cap*ic_cap+-1.07500e-06*ic_cap+1.21000e-04'
+ mcm4m3m1_ca_w_0_300_s_0_600 = '-2.08750e-06*ic_cap*ic_cap+-1.07500e-06*ic_cap+1.21000e-04'
+ mcm4m3m1_ca_w_0_300_s_0_800 = '-2.08750e-06*ic_cap*ic_cap+-1.07500e-06*ic_cap+1.21000e-04'
+ mcm4m3m1_ca_w_0_300_s_1_000 = '-2.08750e-06*ic_cap*ic_cap+-1.07500e-06*ic_cap+1.21000e-04'
+ mcm4m3m1_ca_w_0_300_s_1_200 = '-2.08750e-06*ic_cap*ic_cap+-1.07500e-06*ic_cap+1.21000e-04'
+ mcm4m3m1_ca_w_0_300_s_2_100 = '-2.08750e-06*ic_cap*ic_cap+-1.07500e-06*ic_cap+1.21000e-04'
+ mcm4m3m1_ca_w_0_300_s_3_300 = '-2.08750e-06*ic_cap*ic_cap+-1.07500e-06*ic_cap+1.21000e-04'
+ mcm4m3m1_ca_w_0_300_s_9_000 = '-2.08750e-06*ic_cap*ic_cap+-1.07500e-06*ic_cap+1.21000e-04'
+ mcm4m3m1_ca_w_2_400_s_0_300 = '-2.08750e-06*ic_cap*ic_cap+-1.07500e-06*ic_cap+1.21000e-04'
+ mcm4m3m1_ca_w_2_400_s_0_360 = '-2.08750e-06*ic_cap*ic_cap+-1.07500e-06*ic_cap+1.21000e-04'
+ mcm4m3m1_ca_w_2_400_s_0_450 = '-2.08750e-06*ic_cap*ic_cap+-1.07500e-06*ic_cap+1.21000e-04'
+ mcm4m3m1_ca_w_2_400_s_0_600 = '-2.08750e-06*ic_cap*ic_cap+-1.07500e-06*ic_cap+1.21000e-04'
+ mcm4m3m1_ca_w_2_400_s_0_800 = '-2.08750e-06*ic_cap*ic_cap+-1.07500e-06*ic_cap+1.21000e-04'
+ mcm4m3m1_ca_w_2_400_s_1_000 = '-2.08750e-06*ic_cap*ic_cap+-1.07500e-06*ic_cap+1.21000e-04'
+ mcm4m3m1_ca_w_2_400_s_1_200 = '-2.08750e-06*ic_cap*ic_cap+-1.07500e-06*ic_cap+1.21000e-04'
+ mcm4m3m1_ca_w_2_400_s_2_100 = '-2.08750e-06*ic_cap*ic_cap+-1.07500e-06*ic_cap+1.21000e-04'
+ mcm4m3m1_ca_w_2_400_s_3_300 = '-2.08750e-06*ic_cap*ic_cap+-1.07500e-06*ic_cap+1.21000e-04'
+ mcm4m3m1_ca_w_2_400_s_9_000 = '-2.08750e-06*ic_cap*ic_cap+-1.07500e-06*ic_cap+1.21000e-04'
+ mcm4m3m1_cc_w_0_300_s_0_300 = '-5.06250e-13*ic_cap*ic_cap+-3.00000e-13*ic_cap+8.60000e-11'
+ mcm4m3m1_cc_w_0_300_s_0_360 = '-4.25000e-13*ic_cap*ic_cap+-2.75000e-13*ic_cap+7.78000e-11'
+ mcm4m3m1_cc_w_0_300_s_0_450 = '-2.96875e-13*ic_cap*ic_cap+-1.87500e-13*ic_cap+6.70000e-11'
+ mcm4m3m1_cc_w_0_300_s_0_600 = '-1.62500e-13*ic_cap*ic_cap+-1.00000e-13*ic_cap+5.24000e-11'
+ mcm4m3m1_cc_w_0_300_s_0_800 = '-3.75000e-14*ic_cap*ic_cap+-5.00000e-14*ic_cap+3.81000e-11'
+ mcm4m3m1_cc_w_0_300_s_1_000 = '2.50000e-14*ic_cap*ic_cap+2.80000e-11'
+ mcm4m3m1_cc_w_0_300_s_1_200 = '7.18750e-14*ic_cap*ic_cap+3.75000e-14*ic_cap+2.06000e-11'
+ mcm4m3m1_cc_w_0_300_s_2_100 = '8.18750e-14*ic_cap*ic_cap+5.25000e-14*ic_cap+5.72000e-12'
+ mcm4m3m1_cc_w_0_300_s_3_300 = '3.46875e-14*ic_cap*ic_cap+2.12500e-14*ic_cap+1.13000e-12'
+ mcm4m3m1_cc_w_0_300_s_9_000 = '-4.68750e-16*ic_cap*ic_cap+-6.25000e-16*ic_cap+3.50000e-14'
+ mcm4m3m1_cc_w_2_400_s_0_300 = '-4.21875e-13*ic_cap*ic_cap+-2.37500e-13*ic_cap+8.85000e-11'
+ mcm4m3m1_cc_w_2_400_s_0_360 = '-3.21875e-13*ic_cap*ic_cap+-1.87500e-13*ic_cap+7.98000e-11'
+ mcm4m3m1_cc_w_2_400_s_0_450 = '-2.15625e-13*ic_cap*ic_cap+-1.37500e-13*ic_cap+6.87000e-11'
+ mcm4m3m1_cc_w_2_400_s_0_600 = '-8.75000e-14*ic_cap*ic_cap+-5.00000e-14*ic_cap+5.38000e-11'
+ mcm4m3m1_cc_w_2_400_s_0_800 = '1.56250e-14*ic_cap*ic_cap+1.25000e-14*ic_cap+3.91000e-11'
+ mcm4m3m1_cc_w_2_400_s_1_000 = '7.50000e-14*ic_cap*ic_cap+5.00000e-14*ic_cap+2.86000e-11'
+ mcm4m3m1_cc_w_2_400_s_1_200 = '9.68750e-14*ic_cap*ic_cap+6.25000e-14*ic_cap+2.13000e-11'
+ mcm4m3m1_cc_w_2_400_s_2_100 = '9.87500e-14*ic_cap*ic_cap+5.75000e-14*ic_cap+5.90000e-12'
+ mcm4m3m1_cc_w_2_400_s_3_300 = '3.75000e-14*ic_cap*ic_cap+2.50000e-14*ic_cap+1.20000e-12'
+ mcm4m3m1_cc_w_2_400_s_9_000 = '-3.12500e-15*ic_cap*ic_cap+5.00000e-14'
+ mcm4m3m1_cf_w_0_300_s_0_300 = '-1.50000e-13*ic_cap*ic_cap+-7.50000e-14*ic_cap+1.56000e-11'
+ mcm4m3m1_cf_w_0_300_s_0_360 = '-1.93750e-13*ic_cap*ic_cap+-1.00000e-13*ic_cap+1.85000e-11'
+ mcm4m3m1_cf_w_0_300_s_0_450 = '-2.46875e-13*ic_cap*ic_cap+-1.37500e-13*ic_cap+2.25000e-11'
+ mcm4m3m1_cf_w_0_300_s_0_600 = '-3.25000e-13*ic_cap*ic_cap+-1.75000e-13*ic_cap+2.86000e-11'
+ mcm4m3m1_cf_w_0_300_s_0_800 = '-4.09375e-13*ic_cap*ic_cap+-2.37500e-13*ic_cap+3.57000e-11'
+ mcm4m3m1_cf_w_0_300_s_1_000 = '-4.62500e-13*ic_cap*ic_cap+-2.75000e-13*ic_cap+4.16000e-11'
+ mcm4m3m1_cf_w_0_300_s_1_200 = '-5.03125e-13*ic_cap*ic_cap+-2.87500e-13*ic_cap+4.64000e-11'
+ mcm4m3m1_cf_w_0_300_s_2_100 = '-5.50000e-13*ic_cap*ic_cap+-3.25000e-13*ic_cap+5.84000e-11'
+ mcm4m3m1_cf_w_0_300_s_3_300 = '-5.06250e-13*ic_cap*ic_cap+-3.25000e-13*ic_cap+6.27000e-11'
+ mcm4m3m1_cf_w_0_300_s_9_000 = '-4.71875e-13*ic_cap*ic_cap+-2.87500e-13*ic_cap+6.39000e-11'
+ mcm4m3m1_cf_w_2_400_s_0_300 = '-1.50000e-13*ic_cap*ic_cap+-7.50000e-14*ic_cap+1.57000e-11'
+ mcm4m3m1_cf_w_2_400_s_0_360 = '-1.93750e-13*ic_cap*ic_cap+-1.00000e-13*ic_cap+1.86000e-11'
+ mcm4m3m1_cf_w_2_400_s_0_450 = '-2.46875e-13*ic_cap*ic_cap+-1.37500e-13*ic_cap+2.26000e-11'
+ mcm4m3m1_cf_w_2_400_s_0_600 = '-3.18750e-13*ic_cap*ic_cap+-1.75000e-13*ic_cap+2.87000e-11'
+ mcm4m3m1_cf_w_2_400_s_0_800 = '-4.03125e-13*ic_cap*ic_cap+-2.37500e-13*ic_cap+3.59000e-11'
+ mcm4m3m1_cf_w_2_400_s_1_000 = '-4.56250e-13*ic_cap*ic_cap+-2.75000e-13*ic_cap+4.18000e-11'
+ mcm4m3m1_cf_w_2_400_s_1_200 = '-5.03125e-13*ic_cap*ic_cap+-2.87500e-13*ic_cap+4.68000e-11'
+ mcm4m3m1_cf_w_2_400_s_2_100 = '-5.34375e-13*ic_cap*ic_cap+-3.37500e-13*ic_cap+5.90000e-11'
+ mcm4m3m1_cf_w_2_400_s_3_300 = '-4.81250e-13*ic_cap*ic_cap+-3.00000e-13*ic_cap+6.35000e-11'
+ mcm4m3m1_cf_w_2_400_s_9_000 = '-4.43750e-13*ic_cap*ic_cap+-2.75000e-13*ic_cap+6.47000e-11'
+ mcm4m3m2_ca_w_0_300_s_0_300 = '-3.00000e-06*ic_cap*ic_cap+-1.50000e-06*ic_cap+1.71000e-04'
+ mcm4m3m2_ca_w_0_300_s_0_360 = '-3.00000e-06*ic_cap*ic_cap+-1.50000e-06*ic_cap+1.71000e-04'
+ mcm4m3m2_ca_w_0_300_s_0_450 = '-3.00000e-06*ic_cap*ic_cap+-1.50000e-06*ic_cap+1.71000e-04'
+ mcm4m3m2_ca_w_0_300_s_0_600 = '-3.00000e-06*ic_cap*ic_cap+-1.50000e-06*ic_cap+1.71000e-04'
+ mcm4m3m2_ca_w_0_300_s_0_800 = '-3.00000e-06*ic_cap*ic_cap+-1.50000e-06*ic_cap+1.71000e-04'
+ mcm4m3m2_ca_w_0_300_s_1_000 = '-3.00000e-06*ic_cap*ic_cap+-1.50000e-06*ic_cap+1.71000e-04'
+ mcm4m3m2_ca_w_0_300_s_1_200 = '-3.00000e-06*ic_cap*ic_cap+-1.50000e-06*ic_cap+1.71000e-04'
+ mcm4m3m2_ca_w_0_300_s_2_100 = '-3.00000e-06*ic_cap*ic_cap+-1.50000e-06*ic_cap+1.71000e-04'
+ mcm4m3m2_ca_w_0_300_s_3_300 = '-3.00000e-06*ic_cap*ic_cap+-1.50000e-06*ic_cap+1.71000e-04'
+ mcm4m3m2_ca_w_0_300_s_9_000 = '-3.00000e-06*ic_cap*ic_cap+-1.50000e-06*ic_cap+1.71000e-04'
+ mcm4m3m2_ca_w_2_400_s_0_300 = '-3.00000e-06*ic_cap*ic_cap+-1.50000e-06*ic_cap+1.71000e-04'
+ mcm4m3m2_ca_w_2_400_s_0_360 = '-3.00000e-06*ic_cap*ic_cap+-1.50000e-06*ic_cap+1.71000e-04'
+ mcm4m3m2_ca_w_2_400_s_0_450 = '-3.00000e-06*ic_cap*ic_cap+-1.50000e-06*ic_cap+1.71000e-04'
+ mcm4m3m2_ca_w_2_400_s_0_600 = '-3.00000e-06*ic_cap*ic_cap+-1.50000e-06*ic_cap+1.71000e-04'
+ mcm4m3m2_ca_w_2_400_s_0_800 = '-3.00000e-06*ic_cap*ic_cap+-1.50000e-06*ic_cap+1.71000e-04'
+ mcm4m3m2_ca_w_2_400_s_1_000 = '-3.00000e-06*ic_cap*ic_cap+-1.50000e-06*ic_cap+1.71000e-04'
+ mcm4m3m2_ca_w_2_400_s_1_200 = '-3.00000e-06*ic_cap*ic_cap+-1.50000e-06*ic_cap+1.71000e-04'
+ mcm4m3m2_ca_w_2_400_s_2_100 = '-3.00000e-06*ic_cap*ic_cap+-1.50000e-06*ic_cap+1.71000e-04'
+ mcm4m3m2_ca_w_2_400_s_3_300 = '-3.00000e-06*ic_cap*ic_cap+-1.50000e-06*ic_cap+1.71000e-04'
+ mcm4m3m2_ca_w_2_400_s_9_000 = '-3.00000e-06*ic_cap*ic_cap+-1.50000e-06*ic_cap+1.71000e-04'
+ mcm4m3m2_cc_w_0_300_s_0_300 = '-4.21875e-13*ic_cap*ic_cap+-2.37500e-13*ic_cap+7.80000e-11'
+ mcm4m3m2_cc_w_0_300_s_0_360 = '-3.37500e-13*ic_cap*ic_cap+-2.00000e-13*ic_cap+6.98000e-11'
+ mcm4m3m2_cc_w_0_300_s_0_450 = '-2.25000e-13*ic_cap*ic_cap+-1.50000e-13*ic_cap+5.89000e-11'
+ mcm4m3m2_cc_w_0_300_s_0_600 = '-9.06250e-14*ic_cap*ic_cap+-6.25000e-14*ic_cap+4.42000e-11'
+ mcm4m3m2_cc_w_0_300_s_0_800 = '1.87500e-14*ic_cap*ic_cap+3.01000e-11'
+ mcm4m3m2_cc_w_0_300_s_1_000 = '7.50000e-14*ic_cap*ic_cap+2.50000e-14*ic_cap+2.03000e-11'
+ mcm4m3m2_cc_w_0_300_s_1_200 = '9.68750e-14*ic_cap*ic_cap+6.25000e-14*ic_cap+1.37000e-11'
+ mcm4m3m2_cc_w_0_300_s_2_100 = '5.75000e-14*ic_cap*ic_cap+4.50000e-14*ic_cap+2.53000e-12'
+ mcm4m3m2_cc_w_0_300_s_3_300 = '1.14063e-14*ic_cap*ic_cap+1.31250e-14*ic_cap+3.70000e-13'
+ mcm4m3m2_cc_w_0_300_s_9_000 = '6.25000e-16*ic_cap*ic_cap+2.50000e-14'
+ mcm4m3m2_cc_w_2_400_s_0_300 = '-3.87500e-13*ic_cap*ic_cap+-2.25000e-13*ic_cap+7.87000e-11'
+ mcm4m3m2_cc_w_2_400_s_0_360 = '-3.03125e-13*ic_cap*ic_cap+-1.62500e-13*ic_cap+7.04000e-11'
+ mcm4m3m2_cc_w_2_400_s_0_450 = '-1.81250e-13*ic_cap*ic_cap+-1.00000e-13*ic_cap+5.91000e-11'
+ mcm4m3m2_cc_w_2_400_s_0_600 = '-6.56250e-14*ic_cap*ic_cap+-3.75000e-14*ic_cap+4.46000e-11'
+ mcm4m3m2_cc_w_2_400_s_0_800 = '3.75000e-14*ic_cap*ic_cap+2.50000e-14*ic_cap+3.03000e-11'
+ mcm4m3m2_cc_w_2_400_s_1_000 = '7.50000e-14*ic_cap*ic_cap+5.00000e-14*ic_cap+2.08000e-11'
+ mcm4m3m2_cc_w_2_400_s_1_200 = '1.06250e-13*ic_cap*ic_cap+7.50000e-14*ic_cap+1.39000e-11'
+ mcm4m3m2_cc_w_2_400_s_2_100 = '5.78125e-14*ic_cap*ic_cap+4.37500e-14*ic_cap+2.55000e-12'
+ mcm4m3m2_cc_w_2_400_s_3_300 = '1.09375e-14*ic_cap*ic_cap+1.87500e-14*ic_cap+3.50000e-13'
+ mcm4m3m2_cc_w_2_400_s_9_000 = '-3.12500e-15*ic_cap*ic_cap+5.00000e-14'
+ mcm4m3m2_cf_w_0_300_s_0_300 = '-2.18750e-13*ic_cap*ic_cap+-1.25000e-13*ic_cap+2.20000e-11'
+ mcm4m3m2_cf_w_0_300_s_0_360 = '-2.71875e-13*ic_cap*ic_cap+-1.37500e-13*ic_cap+2.58000e-11'
+ mcm4m3m2_cf_w_0_300_s_0_450 = '-3.53125e-13*ic_cap*ic_cap+-1.87500e-13*ic_cap+3.13000e-11'
+ mcm4m3m2_cf_w_0_300_s_0_600 = '-4.59375e-13*ic_cap*ic_cap+-2.37500e-13*ic_cap+3.94000e-11'
+ mcm4m3m2_cf_w_0_300_s_0_800 = '-5.59375e-13*ic_cap*ic_cap+-3.12500e-13*ic_cap+4.83000e-11'
+ mcm4m3m2_cf_w_0_300_s_1_000 = '-6.28125e-13*ic_cap*ic_cap+-3.37500e-13*ic_cap+5.54000e-11'
+ mcm4m3m2_cf_w_0_300_s_1_200 = '-6.56250e-13*ic_cap*ic_cap+-3.75000e-13*ic_cap+6.05000e-11'
+ mcm4m3m2_cf_w_0_300_s_2_100 = '-6.53125e-13*ic_cap*ic_cap+-3.87500e-13*ic_cap+7.07000e-11'
+ mcm4m3m2_cf_w_0_300_s_3_300 = '-6.03125e-13*ic_cap*ic_cap+-3.37500e-13*ic_cap+7.29000e-11'
+ mcm4m3m2_cf_w_0_300_s_9_000 = '-6.12500e-13*ic_cap*ic_cap+-3.50000e-13*ic_cap+7.35000e-11'
+ mcm4m3m2_cf_w_2_400_s_0_300 = '-2.21875e-13*ic_cap*ic_cap+-1.12500e-13*ic_cap+2.21000e-11'
+ mcm4m3m2_cf_w_2_400_s_0_360 = '-2.78125e-13*ic_cap*ic_cap+-1.37500e-13*ic_cap+2.60000e-11'
+ mcm4m3m2_cf_w_2_400_s_0_450 = '-3.50000e-13*ic_cap*ic_cap+-2.00000e-13*ic_cap+3.14000e-11'
+ mcm4m3m2_cf_w_2_400_s_0_600 = '-4.56250e-13*ic_cap*ic_cap+-2.50000e-13*ic_cap+3.95000e-11'
+ mcm4m3m2_cf_w_2_400_s_0_800 = '-5.56250e-13*ic_cap*ic_cap+-3.00000e-13*ic_cap+4.85000e-11'
+ mcm4m3m2_cf_w_2_400_s_1_000 = '-6.03125e-13*ic_cap*ic_cap+-3.37500e-13*ic_cap+5.54000e-11'
+ mcm4m3m2_cf_w_2_400_s_1_200 = '-6.34375e-13*ic_cap*ic_cap+-3.62500e-13*ic_cap+6.06000e-11'
+ mcm4m3m2_cf_w_2_400_s_2_100 = '-6.37500e-13*ic_cap*ic_cap+-3.75000e-13*ic_cap+7.12000e-11'
+ mcm4m3m2_cf_w_2_400_s_3_300 = '-5.84375e-13*ic_cap*ic_cap+-3.62500e-13*ic_cap+7.32000e-11'
+ mcm4m3m2_cf_w_2_400_s_9_000 = '-5.87500e-13*ic_cap*ic_cap+-3.75000e-13*ic_cap+7.38000e-11'
+ mcm4m3p1_ca_w_0_300_s_0_300 = '-1.87500e-06*ic_cap*ic_cap+-9.50000e-07*ic_cap+1.04000e-04'
+ mcm4m3p1_ca_w_0_300_s_0_360 = '-1.87500e-06*ic_cap*ic_cap+-9.50000e-07*ic_cap+1.04000e-04'
+ mcm4m3p1_ca_w_0_300_s_0_450 = '-1.87500e-06*ic_cap*ic_cap+-9.50000e-07*ic_cap+1.04000e-04'
+ mcm4m3p1_ca_w_0_300_s_0_600 = '-1.87500e-06*ic_cap*ic_cap+-9.50000e-07*ic_cap+1.04000e-04'
+ mcm4m3p1_ca_w_0_300_s_0_800 = '-1.87500e-06*ic_cap*ic_cap+-9.50000e-07*ic_cap+1.04000e-04'
+ mcm4m3p1_ca_w_0_300_s_1_000 = '-1.87500e-06*ic_cap*ic_cap+-9.50000e-07*ic_cap+1.04000e-04'
+ mcm4m3p1_ca_w_0_300_s_1_200 = '-1.87500e-06*ic_cap*ic_cap+-9.50000e-07*ic_cap+1.04000e-04'
+ mcm4m3p1_ca_w_0_300_s_2_100 = '-1.87500e-06*ic_cap*ic_cap+-9.50000e-07*ic_cap+1.04000e-04'
+ mcm4m3p1_ca_w_0_300_s_3_300 = '-1.87500e-06*ic_cap*ic_cap+-9.50000e-07*ic_cap+1.04000e-04'
+ mcm4m3p1_ca_w_0_300_s_9_000 = '-1.87500e-06*ic_cap*ic_cap+-9.50000e-07*ic_cap+1.04000e-04'
+ mcm4m3p1_ca_w_2_400_s_0_300 = '-1.87500e-06*ic_cap*ic_cap+-9.50000e-07*ic_cap+1.04000e-04'
+ mcm4m3p1_ca_w_2_400_s_0_360 = '-1.87500e-06*ic_cap*ic_cap+-9.50000e-07*ic_cap+1.04000e-04'
+ mcm4m3p1_ca_w_2_400_s_0_450 = '-1.87500e-06*ic_cap*ic_cap+-9.50000e-07*ic_cap+1.04000e-04'
+ mcm4m3p1_ca_w_2_400_s_0_600 = '-1.87500e-06*ic_cap*ic_cap+-9.50000e-07*ic_cap+1.04000e-04'
+ mcm4m3p1_ca_w_2_400_s_0_800 = '-1.87500e-06*ic_cap*ic_cap+-9.50000e-07*ic_cap+1.04000e-04'
+ mcm4m3p1_ca_w_2_400_s_1_000 = '-1.87500e-06*ic_cap*ic_cap+-9.50000e-07*ic_cap+1.04000e-04'
+ mcm4m3p1_ca_w_2_400_s_1_200 = '-1.87500e-06*ic_cap*ic_cap+-9.50000e-07*ic_cap+1.04000e-04'
+ mcm4m3p1_ca_w_2_400_s_2_100 = '-1.87500e-06*ic_cap*ic_cap+-9.50000e-07*ic_cap+1.04000e-04'
+ mcm4m3p1_ca_w_2_400_s_3_300 = '-1.87500e-06*ic_cap*ic_cap+-9.50000e-07*ic_cap+1.04000e-04'
+ mcm4m3p1_ca_w_2_400_s_9_000 = '-1.87500e-06*ic_cap*ic_cap+-9.50000e-07*ic_cap+1.04000e-04'
+ mcm4m3p1_cc_w_0_300_s_0_300 = '-5.56250e-13*ic_cap*ic_cap+-3.50000e-13*ic_cap+8.99000e-11'
+ mcm4m3p1_cc_w_0_300_s_0_360 = '-4.71875e-13*ic_cap*ic_cap+-2.87500e-13*ic_cap+8.20000e-11'
+ mcm4m3p1_cc_w_0_300_s_0_450 = '-3.21875e-13*ic_cap*ic_cap+-2.37500e-13*ic_cap+7.10000e-11'
+ mcm4m3p1_cc_w_0_300_s_0_600 = '-2.06250e-13*ic_cap*ic_cap+-1.25000e-13*ic_cap+5.73000e-11'
+ mcm4m3p1_cc_w_0_300_s_0_800 = '-8.43750e-14*ic_cap*ic_cap+-6.25000e-14*ic_cap+4.35000e-11'
+ mcm4m3p1_cc_w_0_300_s_1_000 = '-3.12500e-15*ic_cap*ic_cap+-1.25000e-14*ic_cap+3.33000e-11'
+ mcm4m3p1_cc_w_0_300_s_1_200 = '3.12500e-14*ic_cap*ic_cap+2.60000e-11'
+ mcm4m3p1_cc_w_0_300_s_2_100 = '7.87500e-14*ic_cap*ic_cap+5.00000e-14*ic_cap+9.64000e-12'
+ mcm4m3p1_cc_w_0_300_s_3_300 = '5.62500e-14*ic_cap*ic_cap+3.50000e-14*ic_cap+2.96000e-12'
+ mcm4m3p1_cc_w_0_300_s_9_000 = '3.90625e-15*ic_cap*ic_cap+3.12500e-15*ic_cap+3.50000e-14'
+ mcm4m3p1_cc_w_2_400_s_0_300 = '-4.50000e-13*ic_cap*ic_cap+-2.75000e-13*ic_cap+9.64000e-11'
+ mcm4m3p1_cc_w_2_400_s_0_360 = '-3.59375e-13*ic_cap*ic_cap+-1.87500e-13*ic_cap+8.78000e-11'
+ mcm4m3p1_cc_w_2_400_s_0_450 = '-2.40625e-13*ic_cap*ic_cap+-1.37500e-13*ic_cap+7.65000e-11'
+ mcm4m3p1_cc_w_2_400_s_0_600 = '-1.09375e-13*ic_cap*ic_cap+-6.25000e-14*ic_cap+6.16000e-11'
+ mcm4m3p1_cc_w_2_400_s_0_800 = '-9.37500e-15*ic_cap*ic_cap+-1.25000e-14*ic_cap+4.69000e-11'
+ mcm4m3p1_cc_w_2_400_s_1_000 = '5.62500e-14*ic_cap*ic_cap+2.50000e-14*ic_cap+3.62000e-11'
+ mcm4m3p1_cc_w_2_400_s_1_200 = '9.68750e-14*ic_cap*ic_cap+6.25000e-14*ic_cap+2.83000e-11'
+ mcm4m3p1_cc_w_2_400_s_2_100 = '1.18750e-13*ic_cap*ic_cap+7.50000e-14*ic_cap+1.09000e-11'
+ mcm4m3p1_cc_w_2_400_s_3_300 = '7.81250e-14*ic_cap*ic_cap+6.00000e-14*ic_cap+3.43000e-12'
+ mcm4m3p1_cc_w_2_400_s_9_000 = '3.28125e-15*ic_cap*ic_cap+3.12500e-15*ic_cap+4.00000e-14'
+ mcm4m3p1_cf_w_0_300_s_0_300 = '-1.43750e-13*ic_cap*ic_cap+-7.50000e-14*ic_cap+1.33000e-11'
+ mcm4m3p1_cf_w_0_300_s_0_360 = '-1.71875e-13*ic_cap*ic_cap+-8.75000e-14*ic_cap+1.56000e-11'
+ mcm4m3p1_cf_w_0_300_s_0_450 = '-2.21875e-13*ic_cap*ic_cap+-1.12500e-13*ic_cap+1.91000e-11'
+ mcm4m3p1_cf_w_0_300_s_0_600 = '-2.93750e-13*ic_cap*ic_cap+-1.50000e-13*ic_cap+2.43000e-11'
+ mcm4m3p1_cf_w_0_300_s_0_800 = '-3.56250e-13*ic_cap*ic_cap+-2.00000e-13*ic_cap+3.02000e-11'
+ mcm4m3p1_cf_w_0_300_s_1_000 = '-4.12500e-13*ic_cap*ic_cap+-2.25000e-13*ic_cap+3.53000e-11'
+ mcm4m3p1_cf_w_0_300_s_1_200 = '-4.46875e-13*ic_cap*ic_cap+-2.62500e-13*ic_cap+3.96000e-11'
+ mcm4m3p1_cf_w_0_300_s_2_100 = '-5.09375e-13*ic_cap*ic_cap+-3.12500e-13*ic_cap+5.15000e-11'
+ mcm4m3p1_cf_w_0_300_s_3_300 = '-4.96875e-13*ic_cap*ic_cap+-2.87500e-13*ic_cap+5.75000e-11'
+ mcm4m3p1_cf_w_0_300_s_9_000 = '-4.50000e-13*ic_cap*ic_cap+-2.75000e-13*ic_cap+6.04000e-11'
+ mcm4m3p1_cf_w_2_400_s_0_300 = '-1.40625e-13*ic_cap*ic_cap+-6.25000e-14*ic_cap+1.34000e-11'
+ mcm4m3p1_cf_w_2_400_s_0_360 = '-1.78125e-13*ic_cap*ic_cap+-8.75000e-14*ic_cap+1.58000e-11'
+ mcm4m3p1_cf_w_2_400_s_0_450 = '-2.25000e-13*ic_cap*ic_cap+-1.25000e-13*ic_cap+1.92000e-11'
+ mcm4m3p1_cf_w_2_400_s_0_600 = '-2.90625e-13*ic_cap*ic_cap+-1.62500e-13*ic_cap+2.44000e-11'
+ mcm4m3p1_cf_w_2_400_s_0_800 = '-3.56250e-13*ic_cap*ic_cap+-2.00000e-13*ic_cap+3.04000e-11'
+ mcm4m3p1_cf_w_2_400_s_1_000 = '-4.06250e-13*ic_cap*ic_cap+-2.25000e-13*ic_cap+3.56000e-11'
+ mcm4m3p1_cf_w_2_400_s_1_200 = '-4.43750e-13*ic_cap*ic_cap+-2.50000e-13*ic_cap+3.99000e-11'
+ mcm4m3p1_cf_w_2_400_s_2_100 = '-4.96875e-13*ic_cap*ic_cap+-2.87500e-13*ic_cap+5.23000e-11'
+ mcm4m3p1_cf_w_2_400_s_3_300 = '-4.71875e-13*ic_cap*ic_cap+-2.87500e-13*ic_cap+5.89000e-11'
+ mcm4m3p1_cf_w_2_400_s_9_000 = '-4.03125e-13*ic_cap*ic_cap+-2.37500e-13*ic_cap+6.23000e-11'
+ mcm4p1_ca_w_0_300_s_0_300 = '-9.06250e-08*ic_cap*ic_cap+-5.75000e-08*ic_cap+1.01000e-05'
+ mcm4p1_ca_w_0_300_s_0_360 = '-9.06250e-08*ic_cap*ic_cap+-5.75000e-08*ic_cap+1.01000e-05'
+ mcm4p1_ca_w_0_300_s_0_450 = '-9.06250e-08*ic_cap*ic_cap+-5.75000e-08*ic_cap+1.01000e-05'
+ mcm4p1_ca_w_0_300_s_0_600 = '-9.06250e-08*ic_cap*ic_cap+-5.75000e-08*ic_cap+1.01000e-05'
+ mcm4p1_ca_w_0_300_s_0_800 = '-9.06250e-08*ic_cap*ic_cap+-5.75000e-08*ic_cap+1.01000e-05'
+ mcm4p1_ca_w_0_300_s_1_000 = '-9.06250e-08*ic_cap*ic_cap+-5.75000e-08*ic_cap+1.01000e-05'
+ mcm4p1_ca_w_0_300_s_1_200 = '-9.06250e-08*ic_cap*ic_cap+-5.75000e-08*ic_cap+1.01000e-05'
+ mcm4p1_ca_w_0_300_s_2_100 = '-9.06250e-08*ic_cap*ic_cap+-5.75000e-08*ic_cap+1.01000e-05'
+ mcm4p1_ca_w_0_300_s_3_300 = '-9.06250e-08*ic_cap*ic_cap+-5.75000e-08*ic_cap+1.01000e-05'
+ mcm4p1_ca_w_0_300_s_9_000 = '-9.06250e-08*ic_cap*ic_cap+-5.75000e-08*ic_cap+1.01000e-05'
+ mcm4p1_ca_w_2_400_s_0_300 = '-9.06250e-08*ic_cap*ic_cap+-5.75000e-08*ic_cap+1.01000e-05'
+ mcm4p1_ca_w_2_400_s_0_360 = '-9.06250e-08*ic_cap*ic_cap+-5.75000e-08*ic_cap+1.01000e-05'
+ mcm4p1_ca_w_2_400_s_0_450 = '-9.06250e-08*ic_cap*ic_cap+-5.75000e-08*ic_cap+1.01000e-05'
+ mcm4p1_ca_w_2_400_s_0_600 = '-9.06250e-08*ic_cap*ic_cap+-5.75000e-08*ic_cap+1.01000e-05'
+ mcm4p1_ca_w_2_400_s_0_800 = '-9.06250e-08*ic_cap*ic_cap+-5.75000e-08*ic_cap+1.01000e-05'
+ mcm4p1_ca_w_2_400_s_1_000 = '-9.06250e-08*ic_cap*ic_cap+-5.75000e-08*ic_cap+1.01000e-05'
+ mcm4p1_ca_w_2_400_s_1_200 = '-9.06250e-08*ic_cap*ic_cap+-5.75000e-08*ic_cap+1.01000e-05'
+ mcm4p1_ca_w_2_400_s_2_100 = '-9.06250e-08*ic_cap*ic_cap+-5.75000e-08*ic_cap+1.01000e-05'
+ mcm4p1_ca_w_2_400_s_3_300 = '-9.06250e-08*ic_cap*ic_cap+-5.75000e-08*ic_cap+1.01000e-05'
+ mcm4p1_ca_w_2_400_s_9_000 = '-9.06250e-08*ic_cap*ic_cap+-5.75000e-08*ic_cap+1.01000e-05'
+ mcm4p1_cc_w_0_300_s_0_300 = '-7.84375e-13*ic_cap*ic_cap+-4.62500e-13*ic_cap+1.07000e-10'
+ mcm4p1_cc_w_0_300_s_0_360 = '-7.53125e-13*ic_cap*ic_cap+-4.37500e-13*ic_cap+1.01000e-10'
+ mcm4p1_cc_w_0_300_s_0_450 = '-6.15625e-13*ic_cap*ic_cap+-3.62500e-13*ic_cap+9.12000e-11'
+ mcm4p1_cc_w_0_300_s_0_600 = '-4.84375e-13*ic_cap*ic_cap+-3.12500e-13*ic_cap+7.90000e-11'
+ mcm4p1_cc_w_0_300_s_0_800 = '-3.53125e-13*ic_cap*ic_cap+-2.37500e-13*ic_cap+6.71000e-11'
+ mcm4p1_cc_w_0_300_s_1_000 = '-2.81250e-13*ic_cap*ic_cap+-1.75000e-13*ic_cap+5.83000e-11'
+ mcm4p1_cc_w_0_300_s_1_200 = '-2.21875e-13*ic_cap*ic_cap+-1.37500e-13*ic_cap+5.16000e-11'
+ mcm4p1_cc_w_0_300_s_2_100 = '-1.00000e-13*ic_cap*ic_cap+-7.50000e-14*ic_cap+3.49000e-11'
+ mcm4p1_cc_w_0_300_s_3_300 = '-3.75000e-14*ic_cap*ic_cap+-2.50000e-14*ic_cap+2.47000e-11'
+ mcm4p1_cc_w_0_300_s_9_000 = '2.15625e-14*ic_cap*ic_cap+1.37500e-14*ic_cap+7.99000e-12'
+ mcm4p1_cc_w_2_400_s_0_300 = '-8.12500e-13*ic_cap*ic_cap+-5.00000e-13*ic_cap+1.35000e-10'
+ mcm4p1_cc_w_2_400_s_0_360 = '-7.18750e-13*ic_cap*ic_cap+-3.75000e-13*ic_cap+1.27000e-10'
+ mcm4p1_cc_w_2_400_s_0_450 = '-5.62500e-13*ic_cap*ic_cap+-2.50000e-13*ic_cap+1.15000e-10'
+ mcm4p1_cc_w_2_400_s_0_600 = '-4.62500e-13*ic_cap*ic_cap+-2.75000e-13*ic_cap+1.01000e-10'
+ mcm4p1_cc_w_2_400_s_0_800 = '-3.15625e-13*ic_cap*ic_cap+-1.87500e-13*ic_cap+8.61000e-11'
+ mcm4p1_cc_w_2_400_s_1_000 = '-2.34375e-13*ic_cap*ic_cap+-1.62500e-13*ic_cap+7.52000e-11'
+ mcm4p1_cc_w_2_400_s_1_200 = '-1.78125e-13*ic_cap*ic_cap+-1.12500e-13*ic_cap+6.70000e-11'
+ mcm4p1_cc_w_2_400_s_2_100 = '-5.93750e-14*ic_cap*ic_cap+-3.75000e-14*ic_cap+4.61000e-11'
+ mcm4p1_cc_w_2_400_s_3_300 = '-6.25000e-15*ic_cap*ic_cap+3.29000e-11'
+ mcm4p1_cc_w_2_400_s_9_000 = '3.75000e-14*ic_cap*ic_cap+2.50000e-14*ic_cap+1.17000e-11'
+ mcm4p1_cf_w_0_300_s_0_300 = '-2.81250e-15*ic_cap*ic_cap+-1.25000e-15*ic_cap+1.50000e-12'
+ mcm4p1_cf_w_0_300_s_0_360 = '-5.62500e-15*ic_cap*ic_cap+-5.00000e-15*ic_cap+1.80000e-12'
+ mcm4p1_cf_w_0_300_s_0_450 = '-9.68750e-15*ic_cap*ic_cap+-6.25000e-15*ic_cap+2.26000e-12'
+ mcm4p1_cf_w_0_300_s_0_600 = '-1.56250e-14*ic_cap*ic_cap+-1.00000e-14*ic_cap+3.01000e-12'
+ mcm4p1_cf_w_0_300_s_0_800 = '-2.40625e-14*ic_cap*ic_cap+-1.62500e-14*ic_cap+3.90000e-12'
+ mcm4p1_cf_w_0_300_s_1_000 = '-3.34375e-14*ic_cap*ic_cap+-2.12500e-14*ic_cap+4.83000e-12'
+ mcm4p1_cf_w_0_300_s_1_200 = '-4.09375e-14*ic_cap*ic_cap+-2.62500e-14*ic_cap+5.73000e-12'
+ mcm4p1_cf_w_0_300_s_2_100 = '-7.15625e-14*ic_cap*ic_cap+-4.62500e-14*ic_cap+9.75000e-12'
+ mcm4p1_cf_w_0_300_s_3_300 = '-1.06250e-13*ic_cap*ic_cap+-7.50000e-14*ic_cap+1.38000e-11'
+ mcm4p1_cf_w_0_300_s_9_000 = '-1.62500e-13*ic_cap*ic_cap+-1.00000e-13*ic_cap+2.53000e-11'
+ mcm4p1_cf_w_2_400_s_0_300 = '-3.12500e-15*ic_cap*ic_cap+-2.50000e-15*ic_cap+1.54000e-12'
+ mcm4p1_cf_w_2_400_s_0_360 = '-6.25000e-15*ic_cap*ic_cap+-5.00000e-15*ic_cap+1.84000e-12'
+ mcm4p1_cf_w_2_400_s_0_450 = '-1.03125e-14*ic_cap*ic_cap+-6.25000e-15*ic_cap+2.28000e-12'
+ mcm4p1_cf_w_2_400_s_0_600 = '-1.68750e-14*ic_cap*ic_cap+-1.00000e-14*ic_cap+3.01000e-12'
+ mcm4p1_cf_w_2_400_s_0_800 = '-2.53125e-14*ic_cap*ic_cap+-1.62500e-14*ic_cap+3.96000e-12'
+ mcm4p1_cf_w_2_400_s_1_000 = '-3.34375e-14*ic_cap*ic_cap+-2.12500e-14*ic_cap+4.89000e-12'
+ mcm4p1_cf_w_2_400_s_1_200 = '-4.15625e-14*ic_cap*ic_cap+-2.62500e-14*ic_cap+5.81000e-12'
+ mcm4p1_cf_w_2_400_s_2_100 = '-7.31250e-14*ic_cap*ic_cap+-4.75000e-14*ic_cap+9.67000e-12'
+ mcm4p1_cf_w_2_400_s_3_300 = '-1.06250e-13*ic_cap*ic_cap+-7.50000e-14*ic_cap+1.42000e-11'
+ mcm4p1_cf_w_2_400_s_9_000 = '-1.62500e-13*ic_cap*ic_cap+-1.00000e-13*ic_cap+2.75000e-11'
+ mcm4p1f_ca_w_0_150_s_0_210 = '-1.48437e-06*ic_cap*ic_cap+-8.37500e-07*ic_cap+1.16000e-04'
+ mcm4p1f_ca_w_0_150_s_0_263 = '-1.48437e-06*ic_cap*ic_cap+-8.37500e-07*ic_cap+1.16000e-04'
+ mcm4p1f_ca_w_0_150_s_0_315 = '-1.48437e-06*ic_cap*ic_cap+-8.37500e-07*ic_cap+1.16000e-04'
+ mcm4p1f_ca_w_0_150_s_0_420 = '-1.48437e-06*ic_cap*ic_cap+-8.37500e-07*ic_cap+1.16000e-04'
+ mcm4p1f_ca_w_0_150_s_0_525 = '-1.48437e-06*ic_cap*ic_cap+-8.37500e-07*ic_cap+1.16000e-04'
+ mcm4p1f_ca_w_0_150_s_0_630 = '-1.48437e-06*ic_cap*ic_cap+-8.37500e-07*ic_cap+1.16000e-04'
+ mcm4p1f_ca_w_0_150_s_0_840 = '-1.48437e-06*ic_cap*ic_cap+-8.37500e-07*ic_cap+1.16000e-04'
+ mcm4p1f_ca_w_0_150_s_1_260 = '-1.48437e-06*ic_cap*ic_cap+-8.37500e-07*ic_cap+1.16000e-04'
+ mcm4p1f_ca_w_0_150_s_2_310 = '-1.48437e-06*ic_cap*ic_cap+-8.37500e-07*ic_cap+1.16000e-04'
+ mcm4p1f_ca_w_0_150_s_5_250 = '-1.48437e-06*ic_cap*ic_cap+-8.37500e-07*ic_cap+1.16000e-04'
+ mcm4p1f_ca_w_1_200_s_0_210 = '-1.48437e-06*ic_cap*ic_cap+-8.37500e-07*ic_cap+1.16000e-04'
+ mcm4p1f_ca_w_1_200_s_0_263 = '-1.48437e-06*ic_cap*ic_cap+-8.37500e-07*ic_cap+1.16000e-04'
+ mcm4p1f_ca_w_1_200_s_0_315 = '-1.48437e-06*ic_cap*ic_cap+-8.37500e-07*ic_cap+1.16000e-04'
+ mcm4p1f_ca_w_1_200_s_0_420 = '-1.48437e-06*ic_cap*ic_cap+-8.37500e-07*ic_cap+1.16000e-04'
+ mcm4p1f_ca_w_1_200_s_0_525 = '-1.48437e-06*ic_cap*ic_cap+-8.37500e-07*ic_cap+1.16000e-04'
+ mcm4p1f_ca_w_1_200_s_0_630 = '-1.48437e-06*ic_cap*ic_cap+-8.37500e-07*ic_cap+1.16000e-04'
+ mcm4p1f_ca_w_1_200_s_0_840 = '-1.48437e-06*ic_cap*ic_cap+-8.37500e-07*ic_cap+1.16000e-04'
+ mcm4p1f_ca_w_1_200_s_1_260 = '-1.48437e-06*ic_cap*ic_cap+-8.37500e-07*ic_cap+1.16000e-04'
+ mcm4p1f_ca_w_1_200_s_2_310 = '-1.48437e-06*ic_cap*ic_cap+-8.37500e-07*ic_cap+1.16000e-04'
+ mcm4p1f_ca_w_1_200_s_5_250 = '-1.48437e-06*ic_cap*ic_cap+-8.37500e-07*ic_cap+1.16000e-04'
+ mcm4p1f_cc_w_0_150_s_0_210 = '-5.62500e-13*ic_cap*ic_cap+-3.25000e-13*ic_cap+7.48000e-11'
+ mcm4p1f_cc_w_0_150_s_0_263 = '-3.59375e-13*ic_cap*ic_cap+-2.12500e-13*ic_cap+6.03000e-11'
+ mcm4p1f_cc_w_0_150_s_0_315 = '-2.53125e-13*ic_cap*ic_cap+-1.37500e-13*ic_cap+5.10000e-11'
+ mcm4p1f_cc_w_0_150_s_0_420 = '-1.25000e-13*ic_cap*ic_cap+-7.50000e-14*ic_cap+3.83000e-11'
+ mcm4p1f_cc_w_0_150_s_0_525 = '-6.56250e-14*ic_cap*ic_cap+-3.75000e-14*ic_cap+3.05000e-11'
+ mcm4p1f_cc_w_0_150_s_0_630 = '-2.81250e-14*ic_cap*ic_cap+-1.25000e-14*ic_cap+2.49000e-11'
+ mcm4p1f_cc_w_0_150_s_0_840 = '9.37500e-15*ic_cap*ic_cap+1.25000e-14*ic_cap+1.74000e-11'
+ mcm4p1f_cc_w_0_150_s_1_260 = '2.90625e-14*ic_cap*ic_cap+2.12500e-14*ic_cap+9.22000e-12'
+ mcm4p1f_cc_w_0_150_s_2_310 = '2.56250e-14*ic_cap*ic_cap+1.75000e-14*ic_cap+2.78000e-12'
+ mcm4p1f_cc_w_0_150_s_5_250 = '6.71875e-15*ic_cap*ic_cap+4.37500e-15*ic_cap+2.45000e-13'
+ mcm4p1f_cc_w_1_200_s_0_210 = '-5.21875e-13*ic_cap*ic_cap+-2.87500e-13*ic_cap+8.87000e-11'
+ mcm4p1f_cc_w_1_200_s_0_263 = '-3.18750e-13*ic_cap*ic_cap+-1.75000e-13*ic_cap+7.30000e-11'
+ mcm4p1f_cc_w_1_200_s_0_315 = '-2.03125e-13*ic_cap*ic_cap+-1.12500e-13*ic_cap+6.24000e-11'
+ mcm4p1f_cc_w_1_200_s_0_420 = '-7.81250e-14*ic_cap*ic_cap+-3.75000e-14*ic_cap+4.83000e-11'
+ mcm4p1f_cc_w_1_200_s_0_525 = '-2.50000e-14*ic_cap*ic_cap+3.93000e-11'
+ mcm4p1f_cc_w_1_200_s_0_630 = '9.37500e-15*ic_cap*ic_cap+1.25000e-14*ic_cap+3.28000e-11'
+ mcm4p1f_cc_w_1_200_s_0_840 = '4.68750e-14*ic_cap*ic_cap+3.75000e-14*ic_cap+2.40000e-11'
+ mcm4p1f_cc_w_1_200_s_1_260 = '6.56250e-14*ic_cap*ic_cap+3.75000e-14*ic_cap+1.42000e-11'
+ mcm4p1f_cc_w_1_200_s_2_310 = '5.31250e-14*ic_cap*ic_cap+2.75000e-14*ic_cap+4.91000e-12'
+ mcm4p1f_cc_w_1_200_s_5_250 = '9.84375e-15*ic_cap*ic_cap+1.31250e-14*ic_cap+4.80000e-13'
+ mcm4p1f_cf_w_0_150_s_0_210 = '-9.56250e-14*ic_cap*ic_cap+-5.75000e-14*ic_cap+1.14000e-11'
+ mcm4p1f_cf_w_0_150_s_0_263 = '-1.25000e-13*ic_cap*ic_cap+-7.50000e-14*ic_cap+1.38000e-11'
+ mcm4p1f_cf_w_0_150_s_0_315 = '-1.53125e-13*ic_cap*ic_cap+-8.75000e-14*ic_cap+1.61000e-11'
+ mcm4p1f_cf_w_0_150_s_0_420 = '-1.93750e-13*ic_cap*ic_cap+-1.00000e-13*ic_cap+2.04000e-11'
+ mcm4p1f_cf_w_0_150_s_0_525 = '-2.28125e-13*ic_cap*ic_cap+-1.37500e-13*ic_cap+2.40000e-11'
+ mcm4p1f_cf_w_0_150_s_0_630 = '-2.56250e-13*ic_cap*ic_cap+-1.50000e-13*ic_cap+2.72000e-11'
+ mcm4p1f_cf_w_0_150_s_0_840 = '-2.87500e-13*ic_cap*ic_cap+-1.75000e-13*ic_cap+3.22000e-11'
+ mcm4p1f_cf_w_0_150_s_1_260 = '-3.09375e-13*ic_cap*ic_cap+-1.87500e-13*ic_cap+3.88000e-11'
+ mcm4p1f_cf_w_0_150_s_2_310 = '-3.09375e-13*ic_cap*ic_cap+-1.87500e-13*ic_cap+4.45000e-11'
+ mcm4p1f_cf_w_0_150_s_5_250 = '-2.93750e-13*ic_cap*ic_cap+-1.75000e-13*ic_cap+4.71000e-11'
+ mcm4p1f_cf_w_1_200_s_0_210 = '-9.46875e-14*ic_cap*ic_cap+-5.37500e-14*ic_cap+1.13000e-11'
+ mcm4p1f_cf_w_1_200_s_0_263 = '-1.21875e-13*ic_cap*ic_cap+-6.25000e-14*ic_cap+1.38000e-11'
+ mcm4p1f_cf_w_1_200_s_0_315 = '-1.46875e-13*ic_cap*ic_cap+-8.75000e-14*ic_cap+1.61000e-11'
+ mcm4p1f_cf_w_1_200_s_0_420 = '-1.90625e-13*ic_cap*ic_cap+-1.12500e-13*ic_cap+2.04000e-11'
+ mcm4p1f_cf_w_1_200_s_0_525 = '-2.28125e-13*ic_cap*ic_cap+-1.37500e-13*ic_cap+2.42000e-11'
+ mcm4p1f_cf_w_1_200_s_0_630 = '-2.53125e-13*ic_cap*ic_cap+-1.37500e-13*ic_cap+2.75000e-11'
+ mcm4p1f_cf_w_1_200_s_0_840 = '-2.87500e-13*ic_cap*ic_cap+-1.75000e-13*ic_cap+3.29000e-11'
+ mcm4p1f_cf_w_1_200_s_1_260 = '-3.09375e-13*ic_cap*ic_cap+-1.87500e-13*ic_cap+4.01000e-11'
+ mcm4p1f_cf_w_1_200_s_2_310 = '-3.12500e-13*ic_cap*ic_cap+-1.75000e-13*ic_cap+4.84000e-11'
+ mcm4p1f_cf_w_1_200_s_5_250 = '-2.78125e-13*ic_cap*ic_cap+-1.62500e-13*ic_cap+5.27000e-11'
+ mcm5d_ca_w_1_600_s_10_000 = '-4.96875e-08*ic_cap*ic_cap+-3.12500e-08*ic_cap+6.88000e-06'
+ mcm5d_ca_w_1_600_s_12_000 = '-4.96875e-08*ic_cap*ic_cap+-3.12500e-08*ic_cap+6.88000e-06'
+ mcm5d_ca_w_1_600_s_1_600 = '-4.96875e-08*ic_cap*ic_cap+-3.12500e-08*ic_cap+6.88000e-06'
+ mcm5d_ca_w_1_600_s_1_700 = '-4.96875e-08*ic_cap*ic_cap+-3.12500e-08*ic_cap+6.88000e-06'
+ mcm5d_ca_w_1_600_s_1_900 = '-4.96875e-08*ic_cap*ic_cap+-3.12500e-08*ic_cap+6.88000e-06'
+ mcm5d_ca_w_1_600_s_2_000 = '-4.96875e-08*ic_cap*ic_cap+-3.12500e-08*ic_cap+6.88000e-06'
+ mcm5d_ca_w_1_600_s_2_400 = '-4.96875e-08*ic_cap*ic_cap+-3.12500e-08*ic_cap+6.88000e-06'
+ mcm5d_ca_w_1_600_s_2_800 = '-4.96875e-08*ic_cap*ic_cap+-3.12500e-08*ic_cap+6.88000e-06'
+ mcm5d_ca_w_1_600_s_3_200 = '-4.96875e-08*ic_cap*ic_cap+-3.12500e-08*ic_cap+6.88000e-06'
+ mcm5d_ca_w_1_600_s_4_800 = '-4.96875e-08*ic_cap*ic_cap+-3.12500e-08*ic_cap+6.88000e-06'
+ mcm5d_ca_w_4_000_s_10_000 = '-4.96875e-08*ic_cap*ic_cap+-3.12500e-08*ic_cap+6.88000e-06'
+ mcm5d_ca_w_4_000_s_12_000 = '-4.96875e-08*ic_cap*ic_cap+-3.12500e-08*ic_cap+6.88000e-06'
+ mcm5d_ca_w_4_000_s_1_600 = '-4.96875e-08*ic_cap*ic_cap+-3.12500e-08*ic_cap+6.88000e-06'
+ mcm5d_ca_w_4_000_s_1_700 = '-4.96875e-08*ic_cap*ic_cap+-3.12500e-08*ic_cap+6.88000e-06'
+ mcm5d_ca_w_4_000_s_1_900 = '-4.96875e-08*ic_cap*ic_cap+-3.12500e-08*ic_cap+6.88000e-06'
+ mcm5d_ca_w_4_000_s_2_000 = '-4.96875e-08*ic_cap*ic_cap+-3.12500e-08*ic_cap+6.88000e-06'
+ mcm5d_ca_w_4_000_s_2_400 = '-4.96875e-08*ic_cap*ic_cap+-3.12500e-08*ic_cap+6.88000e-06'
+ mcm5d_ca_w_4_000_s_2_800 = '-4.96875e-08*ic_cap*ic_cap+-3.12500e-08*ic_cap+6.88000e-06'
+ mcm5d_ca_w_4_000_s_3_200 = '-4.96875e-08*ic_cap*ic_cap+-3.12500e-08*ic_cap+6.88000e-06'
+ mcm5d_ca_w_4_000_s_4_800 = '-4.96875e-08*ic_cap*ic_cap+-3.12500e-08*ic_cap+6.88000e-06'
+ mcm5d_cc_w_1_600_s_10_000 = '6.25000e-15*ic_cap*ic_cap+1.35000e-11'
+ mcm5d_cc_w_1_600_s_12_000 = '1.25000e-14*ic_cap*ic_cap+1.07000e-11'
+ mcm5d_cc_w_1_600_s_1_600 = '-4.75000e-13*ic_cap*ic_cap+-3.25000e-13*ic_cap+7.31000e-11'
+ mcm5d_cc_w_1_600_s_1_700 = '-4.28125e-13*ic_cap*ic_cap+-2.87500e-13*ic_cap+6.95000e-11'
+ mcm5d_cc_w_1_600_s_1_900 = '-3.46875e-13*ic_cap*ic_cap+-2.37500e-13*ic_cap+6.32000e-11'
+ mcm5d_cc_w_1_600_s_2_000 = '-3.15625e-13*ic_cap*ic_cap+-2.12500e-13*ic_cap+6.06000e-11'
+ mcm5d_cc_w_1_600_s_2_400 = '-2.28125e-13*ic_cap*ic_cap+-1.62500e-13*ic_cap+5.22000e-11'
+ mcm5d_cc_w_1_600_s_2_800 = '-1.68750e-13*ic_cap*ic_cap+-1.25000e-13*ic_cap+4.60000e-11'
+ mcm5d_cc_w_1_600_s_3_200 = '-1.34375e-13*ic_cap*ic_cap+-8.75000e-14*ic_cap+4.13000e-11'
+ mcm5d_cc_w_1_600_s_4_800 = '-5.31250e-14*ic_cap*ic_cap+-3.75000e-14*ic_cap+2.91000e-11'
+ mcm5d_cc_w_4_000_s_10_000 = '1.56250e-14*ic_cap*ic_cap+1.25000e-14*ic_cap+1.61000e-11'
+ mcm5d_cc_w_4_000_s_12_000 = '2.18750e-14*ic_cap*ic_cap+1.25000e-14*ic_cap+1.30000e-11'
+ mcm5d_cc_w_4_000_s_1_600 = '-4.28125e-13*ic_cap*ic_cap+-2.87500e-13*ic_cap+7.98000e-11'
+ mcm5d_cc_w_4_000_s_1_700 = '-3.87500e-13*ic_cap*ic_cap+-2.50000e-13*ic_cap+7.59000e-11'
+ mcm5d_cc_w_4_000_s_1_900 = '-3.18750e-13*ic_cap*ic_cap+-2.00000e-13*ic_cap+6.94000e-11'
+ mcm5d_cc_w_4_000_s_2_000 = '-2.84375e-13*ic_cap*ic_cap+-1.87500e-13*ic_cap+6.66000e-11'
+ mcm5d_cc_w_4_000_s_2_400 = '-2.00000e-13*ic_cap*ic_cap+-1.50000e-13*ic_cap+5.77000e-11'
+ mcm5d_cc_w_4_000_s_2_800 = '-1.46875e-13*ic_cap*ic_cap+-1.12500e-13*ic_cap+5.12000e-11'
+ mcm5d_cc_w_4_000_s_3_200 = '-1.12500e-13*ic_cap*ic_cap+-7.50000e-14*ic_cap+4.61000e-11'
+ mcm5d_cc_w_4_000_s_4_800 = '-3.43750e-14*ic_cap*ic_cap+-3.75000e-14*ic_cap+3.30000e-11'
+ mcm5d_cf_w_1_600_s_10_000 = '-1.28125e-13*ic_cap*ic_cap+-8.75000e-14*ic_cap+2.36000e-11'
+ mcm5d_cf_w_1_600_s_12_000 = '-1.37500e-13*ic_cap*ic_cap+-1.00000e-13*ic_cap+2.59000e-11'
+ mcm5d_cf_w_1_600_s_1_600 = '-2.15625e-14*ic_cap*ic_cap+-1.37500e-14*ic_cap+5.31000e-12'
+ mcm5d_cf_w_1_600_s_1_700 = '-2.34375e-14*ic_cap*ic_cap+-1.62500e-14*ic_cap+5.62000e-12'
+ mcm5d_cf_w_1_600_s_1_900 = '-2.81250e-14*ic_cap*ic_cap+-1.75000e-14*ic_cap+6.25000e-12'
+ mcm5d_cf_w_1_600_s_2_000 = '-3.06250e-14*ic_cap*ic_cap+-2.00000e-14*ic_cap+6.56000e-12'
+ mcm5d_cf_w_1_600_s_2_400 = '-3.90625e-14*ic_cap*ic_cap+-2.62500e-14*ic_cap+7.77000e-12'
+ mcm5d_cf_w_1_600_s_2_800 = '-4.75000e-14*ic_cap*ic_cap+-3.00000e-14*ic_cap+8.95000e-12'
+ mcm5d_cf_w_1_600_s_3_200 = '-5.62500e-14*ic_cap*ic_cap+-3.50000e-14*ic_cap+1.01000e-11'
+ mcm5d_cf_w_1_600_s_4_800 = '-8.12500e-14*ic_cap*ic_cap+-5.00000e-14*ic_cap+1.42000e-11'
+ mcm5d_cf_w_4_000_s_10_000 = '-1.31250e-13*ic_cap*ic_cap+-7.50000e-14*ic_cap+2.41000e-11'
+ mcm5d_cf_w_4_000_s_12_000 = '-1.34375e-13*ic_cap*ic_cap+-8.75000e-14*ic_cap+2.65000e-11'
+ mcm5d_cf_w_4_000_s_1_600 = '-2.09375e-14*ic_cap*ic_cap+-1.37500e-14*ic_cap+5.31000e-12'
+ mcm5d_cf_w_4_000_s_1_700 = '-2.34375e-14*ic_cap*ic_cap+-1.37500e-14*ic_cap+5.63000e-12'
+ mcm5d_cf_w_4_000_s_1_900 = '-2.81250e-14*ic_cap*ic_cap+-1.75000e-14*ic_cap+6.26000e-12'
+ mcm5d_cf_w_4_000_s_2_000 = '-3.06250e-14*ic_cap*ic_cap+-2.00000e-14*ic_cap+6.57000e-12'
+ mcm5d_cf_w_4_000_s_2_400 = '-3.90625e-14*ic_cap*ic_cap+-2.62500e-14*ic_cap+7.78000e-12'
+ mcm5d_cf_w_4_000_s_2_800 = '-4.71875e-14*ic_cap*ic_cap+-3.12500e-14*ic_cap+8.97000e-12'
+ mcm5d_cf_w_4_000_s_3_200 = '-5.43750e-14*ic_cap*ic_cap+-3.50000e-14*ic_cap+1.01000e-11'
+ mcm5d_cf_w_4_000_s_4_800 = '-8.12500e-14*ic_cap*ic_cap+-5.00000e-14*ic_cap+1.43000e-11'
+ mcm5f_ca_w_1_600_s_10_000 = '-4.96875e-08*ic_cap*ic_cap+-3.12500e-08*ic_cap+6.48000e-06'
+ mcm5f_ca_w_1_600_s_12_000 = '-4.96875e-08*ic_cap*ic_cap+-3.12500e-08*ic_cap+6.48000e-06'
+ mcm5f_ca_w_1_600_s_1_600 = '-4.96875e-08*ic_cap*ic_cap+-3.12500e-08*ic_cap+6.48000e-06'
+ mcm5f_ca_w_1_600_s_1_700 = '-4.96875e-08*ic_cap*ic_cap+-3.12500e-08*ic_cap+6.48000e-06'
+ mcm5f_ca_w_1_600_s_1_900 = '-4.96875e-08*ic_cap*ic_cap+-3.12500e-08*ic_cap+6.48000e-06'
+ mcm5f_ca_w_1_600_s_2_000 = '-4.96875e-08*ic_cap*ic_cap+-3.12500e-08*ic_cap+6.48000e-06'
+ mcm5f_ca_w_1_600_s_2_400 = '-4.96875e-08*ic_cap*ic_cap+-3.12500e-08*ic_cap+6.48000e-06'
+ mcm5f_ca_w_1_600_s_2_800 = '-4.96875e-08*ic_cap*ic_cap+-3.12500e-08*ic_cap+6.48000e-06'
+ mcm5f_ca_w_1_600_s_3_200 = '-4.96875e-08*ic_cap*ic_cap+-3.12500e-08*ic_cap+6.48000e-06'
+ mcm5f_ca_w_1_600_s_4_800 = '-4.96875e-08*ic_cap*ic_cap+-3.12500e-08*ic_cap+6.48000e-06'
+ mcm5f_ca_w_4_000_s_10_000 = '-4.96875e-08*ic_cap*ic_cap+-3.12500e-08*ic_cap+6.48000e-06'
+ mcm5f_ca_w_4_000_s_12_000 = '-4.96875e-08*ic_cap*ic_cap+-3.12500e-08*ic_cap+6.48000e-06'
+ mcm5f_ca_w_4_000_s_1_600 = '-4.96875e-08*ic_cap*ic_cap+-3.12500e-08*ic_cap+6.48000e-06'
+ mcm5f_ca_w_4_000_s_1_700 = '-4.96875e-08*ic_cap*ic_cap+-3.12500e-08*ic_cap+6.48000e-06'
+ mcm5f_ca_w_4_000_s_1_900 = '-4.96875e-08*ic_cap*ic_cap+-3.12500e-08*ic_cap+6.48000e-06'
+ mcm5f_ca_w_4_000_s_2_000 = '-4.96875e-08*ic_cap*ic_cap+-3.12500e-08*ic_cap+6.48000e-06'
+ mcm5f_ca_w_4_000_s_2_400 = '-4.96875e-08*ic_cap*ic_cap+-3.12500e-08*ic_cap+6.48000e-06'
+ mcm5f_ca_w_4_000_s_2_800 = '-4.96875e-08*ic_cap*ic_cap+-3.12500e-08*ic_cap+6.48000e-06'
+ mcm5f_ca_w_4_000_s_3_200 = '-4.96875e-08*ic_cap*ic_cap+-3.12500e-08*ic_cap+6.48000e-06'
+ mcm5f_ca_w_4_000_s_4_800 = '-4.96875e-08*ic_cap*ic_cap+-3.12500e-08*ic_cap+6.48000e-06'
+ mcm5f_cc_w_1_600_s_10_000 = '1.25000e-14*ic_cap*ic_cap+1.40000e-11'
+ mcm5f_cc_w_1_600_s_12_000 = '1.87500e-14*ic_cap*ic_cap+1.11000e-11'
+ mcm5f_cc_w_1_600_s_1_600 = '-4.68750e-13*ic_cap*ic_cap+-3.25000e-13*ic_cap+7.35000e-11'
+ mcm5f_cc_w_1_600_s_1_700 = '-4.28125e-13*ic_cap*ic_cap+-2.87500e-13*ic_cap+6.99000e-11'
+ mcm5f_cc_w_1_600_s_1_900 = '-3.46875e-13*ic_cap*ic_cap+-2.37500e-13*ic_cap+6.37000e-11'
+ mcm5f_cc_w_1_600_s_2_000 = '-3.15625e-13*ic_cap*ic_cap+-2.12500e-13*ic_cap+6.11000e-11'
+ mcm5f_cc_w_1_600_s_2_400 = '-2.25000e-13*ic_cap*ic_cap+-1.50000e-13*ic_cap+5.27000e-11'
+ mcm5f_cc_w_1_600_s_2_800 = '-1.68750e-13*ic_cap*ic_cap+-1.25000e-13*ic_cap+4.65000e-11'
+ mcm5f_cc_w_1_600_s_3_200 = '-1.34375e-13*ic_cap*ic_cap+-8.75000e-14*ic_cap+4.18000e-11'
+ mcm5f_cc_w_1_600_s_4_800 = '-5.31250e-14*ic_cap*ic_cap+-3.75000e-14*ic_cap+2.97000e-11'
+ mcm5f_cc_w_4_000_s_10_000 = '2.18750e-14*ic_cap*ic_cap+1.25000e-14*ic_cap+1.66000e-11'
+ mcm5f_cc_w_4_000_s_12_000 = '2.81250e-14*ic_cap*ic_cap+1.25000e-14*ic_cap+1.34000e-11'
+ mcm5f_cc_w_4_000_s_1_600 = '-4.31250e-13*ic_cap*ic_cap+-2.75000e-13*ic_cap+8.04000e-11'
+ mcm5f_cc_w_4_000_s_1_700 = '-3.81250e-13*ic_cap*ic_cap+-2.50000e-13*ic_cap+7.64000e-11'
+ mcm5f_cc_w_4_000_s_1_900 = '-3.06250e-13*ic_cap*ic_cap+-2.00000e-13*ic_cap+6.99000e-11'
+ mcm5f_cc_w_4_000_s_2_000 = '-2.81250e-13*ic_cap*ic_cap+-2.00000e-13*ic_cap+6.72000e-11'
+ mcm5f_cc_w_4_000_s_2_400 = '-1.93750e-13*ic_cap*ic_cap+-1.50000e-13*ic_cap+5.83000e-11'
+ mcm5f_cc_w_4_000_s_2_800 = '-1.43750e-13*ic_cap*ic_cap+-1.00000e-13*ic_cap+5.18000e-11'
+ mcm5f_cc_w_4_000_s_3_200 = '-1.09375e-13*ic_cap*ic_cap+-6.25000e-14*ic_cap+4.67000e-11'
+ mcm5f_cc_w_4_000_s_4_800 = '-3.12500e-14*ic_cap*ic_cap+-2.50000e-14*ic_cap+3.36000e-11'
+ mcm5f_cf_w_1_600_s_10_000 = '-1.34375e-13*ic_cap*ic_cap+-8.75000e-14*ic_cap+2.27000e-11'
+ mcm5f_cf_w_1_600_s_12_000 = '-1.43750e-13*ic_cap*ic_cap+-1.00000e-13*ic_cap+2.50000e-11'
+ mcm5f_cf_w_1_600_s_1_600 = '-2.25000e-14*ic_cap*ic_cap+-1.50000e-14*ic_cap+5.01000e-12'
+ mcm5f_cf_w_1_600_s_1_700 = '-2.46875e-14*ic_cap*ic_cap+-1.62500e-14*ic_cap+5.31000e-12'
+ mcm5f_cf_w_1_600_s_1_900 = '-2.90625e-14*ic_cap*ic_cap+-1.87500e-14*ic_cap+5.90000e-12'
+ mcm5f_cf_w_1_600_s_2_000 = '-3.12500e-14*ic_cap*ic_cap+-2.00000e-14*ic_cap+6.19000e-12'
+ mcm5f_cf_w_1_600_s_2_400 = '-3.96875e-14*ic_cap*ic_cap+-2.62500e-14*ic_cap+7.34000e-12'
+ mcm5f_cf_w_1_600_s_2_800 = '-4.87500e-14*ic_cap*ic_cap+-3.00000e-14*ic_cap+8.47000e-12'
+ mcm5f_cf_w_1_600_s_3_200 = '-5.59375e-14*ic_cap*ic_cap+-3.62500e-14*ic_cap+9.54000e-12'
+ mcm5f_cf_w_1_600_s_4_800 = '-8.12500e-14*ic_cap*ic_cap+-5.00000e-14*ic_cap+1.35000e-11'
+ mcm5f_cf_w_4_000_s_10_000 = '-1.34375e-13*ic_cap*ic_cap+-8.75000e-14*ic_cap+2.31000e-11'
+ mcm5f_cf_w_4_000_s_12_000 = '-1.43750e-13*ic_cap*ic_cap+-1.00000e-13*ic_cap+2.56000e-11'
+ mcm5f_cf_w_4_000_s_1_600 = '-2.28125e-14*ic_cap*ic_cap+-1.37500e-14*ic_cap+5.02000e-12'
+ mcm5f_cf_w_4_000_s_1_700 = '-2.50000e-14*ic_cap*ic_cap+-1.50000e-14*ic_cap+5.32000e-12'
+ mcm5f_cf_w_4_000_s_1_900 = '-2.93750e-14*ic_cap*ic_cap+-1.75000e-14*ic_cap+5.91000e-12'
+ mcm5f_cf_w_4_000_s_2_000 = '-3.12500e-14*ic_cap*ic_cap+-2.00000e-14*ic_cap+6.20000e-12'
+ mcm5f_cf_w_4_000_s_2_400 = '-3.96875e-14*ic_cap*ic_cap+-2.62500e-14*ic_cap+7.35000e-12'
+ mcm5f_cf_w_4_000_s_2_800 = '-4.81250e-14*ic_cap*ic_cap+-3.00000e-14*ic_cap+8.48000e-12'
+ mcm5f_cf_w_4_000_s_3_200 = '-5.59375e-14*ic_cap*ic_cap+-3.62500e-14*ic_cap+9.57000e-12'
+ mcm5f_cf_w_4_000_s_4_800 = '-8.43750e-14*ic_cap*ic_cap+-6.25000e-14*ic_cap+1.36000e-11'
+ mcm5l1_ca_w_1_600_s_10_000 = '-5.75000e-08*ic_cap*ic_cap+-3.75000e-08*ic_cap+8.04000e-06'
+ mcm5l1_ca_w_1_600_s_12_000 = '-5.75000e-08*ic_cap*ic_cap+-3.75000e-08*ic_cap+8.04000e-06'
+ mcm5l1_ca_w_1_600_s_1_600 = '-5.75000e-08*ic_cap*ic_cap+-3.75000e-08*ic_cap+8.04000e-06'
+ mcm5l1_ca_w_1_600_s_1_700 = '-5.75000e-08*ic_cap*ic_cap+-3.75000e-08*ic_cap+8.04000e-06'
+ mcm5l1_ca_w_1_600_s_1_900 = '-5.75000e-08*ic_cap*ic_cap+-3.75000e-08*ic_cap+8.04000e-06'
+ mcm5l1_ca_w_1_600_s_2_000 = '-5.75000e-08*ic_cap*ic_cap+-3.75000e-08*ic_cap+8.04000e-06'
+ mcm5l1_ca_w_1_600_s_2_400 = '-5.75000e-08*ic_cap*ic_cap+-3.75000e-08*ic_cap+8.04000e-06'
+ mcm5l1_ca_w_1_600_s_2_800 = '-5.75000e-08*ic_cap*ic_cap+-3.75000e-08*ic_cap+8.04000e-06'
+ mcm5l1_ca_w_1_600_s_3_200 = '-5.75000e-08*ic_cap*ic_cap+-3.75000e-08*ic_cap+8.04000e-06'
+ mcm5l1_ca_w_1_600_s_4_800 = '-5.75000e-08*ic_cap*ic_cap+-3.75000e-08*ic_cap+8.04000e-06'
+ mcm5l1_ca_w_4_000_s_10_000 = '-5.75000e-08*ic_cap*ic_cap+-3.75000e-08*ic_cap+8.04000e-06'
+ mcm5l1_ca_w_4_000_s_12_000 = '-5.75000e-08*ic_cap*ic_cap+-3.75000e-08*ic_cap+8.04000e-06'
+ mcm5l1_ca_w_4_000_s_1_600 = '-5.75000e-08*ic_cap*ic_cap+-3.75000e-08*ic_cap+8.04000e-06'
+ mcm5l1_ca_w_4_000_s_1_700 = '-5.75000e-08*ic_cap*ic_cap+-3.75000e-08*ic_cap+8.04000e-06'
+ mcm5l1_ca_w_4_000_s_1_900 = '-5.75000e-08*ic_cap*ic_cap+-3.75000e-08*ic_cap+8.04000e-06'
+ mcm5l1_ca_w_4_000_s_2_000 = '-5.75000e-08*ic_cap*ic_cap+-3.75000e-08*ic_cap+8.04000e-06'
+ mcm5l1_ca_w_4_000_s_2_400 = '-5.75000e-08*ic_cap*ic_cap+-3.75000e-08*ic_cap+8.04000e-06'
+ mcm5l1_ca_w_4_000_s_2_800 = '-5.75000e-08*ic_cap*ic_cap+-3.75000e-08*ic_cap+8.04000e-06'
+ mcm5l1_ca_w_4_000_s_3_200 = '-5.75000e-08*ic_cap*ic_cap+-3.75000e-08*ic_cap+8.04000e-06'
+ mcm5l1_ca_w_4_000_s_4_800 = '-5.75000e-08*ic_cap*ic_cap+-3.75000e-08*ic_cap+8.04000e-06'
+ mcm5l1_cc_w_1_600_s_10_000 = '6.25000e-15*ic_cap*ic_cap+1.23000e-11'
+ mcm5l1_cc_w_1_600_s_12_000 = '1.00000e-14*ic_cap*ic_cap+5.00000e-15*ic_cap+9.59000e-12'
+ mcm5l1_cc_w_1_600_s_1_600 = '-4.65625e-13*ic_cap*ic_cap+-3.12500e-13*ic_cap+7.19000e-11'
+ mcm5l1_cc_w_1_600_s_1_700 = '-4.12500e-13*ic_cap*ic_cap+-2.75000e-13*ic_cap+6.82000e-11'
+ mcm5l1_cc_w_1_600_s_1_900 = '-3.43750e-13*ic_cap*ic_cap+-2.25000e-13*ic_cap+6.20000e-11'
+ mcm5l1_cc_w_1_600_s_2_000 = '-3.15625e-13*ic_cap*ic_cap+-2.12500e-13*ic_cap+5.94000e-11'
+ mcm5l1_cc_w_1_600_s_2_400 = '-2.25000e-13*ic_cap*ic_cap+-1.50000e-13*ic_cap+5.09000e-11'
+ mcm5l1_cc_w_1_600_s_2_800 = '-1.71875e-13*ic_cap*ic_cap+-1.12500e-13*ic_cap+4.47000e-11'
+ mcm5l1_cc_w_1_600_s_3_200 = '-1.34375e-13*ic_cap*ic_cap+-8.75000e-14*ic_cap+3.99000e-11'
+ mcm5l1_cc_w_1_600_s_4_800 = '-5.31250e-14*ic_cap*ic_cap+-3.75000e-14*ic_cap+2.77000e-11'
+ mcm5l1_cc_w_4_000_s_10_000 = '1.56250e-14*ic_cap*ic_cap+1.25000e-14*ic_cap+1.48000e-11'
+ mcm5l1_cc_w_4_000_s_12_000 = '1.56250e-14*ic_cap*ic_cap+1.25000e-14*ic_cap+1.18000e-11'
+ mcm5l1_cc_w_4_000_s_1_600 = '-4.34375e-13*ic_cap*ic_cap+-2.87500e-13*ic_cap+7.83000e-11'
+ mcm5l1_cc_w_4_000_s_1_700 = '-3.87500e-13*ic_cap*ic_cap+-2.50000e-13*ic_cap+7.44000e-11'
+ mcm5l1_cc_w_4_000_s_1_900 = '-3.12500e-13*ic_cap*ic_cap+-2.00000e-13*ic_cap+6.78000e-11'
+ mcm5l1_cc_w_4_000_s_2_000 = '-2.87500e-13*ic_cap*ic_cap+-2.00000e-13*ic_cap+6.51000e-11'
+ mcm5l1_cc_w_4_000_s_2_400 = '-2.03125e-13*ic_cap*ic_cap+-1.37500e-13*ic_cap+5.62000e-11'
+ mcm5l1_cc_w_4_000_s_2_800 = '-1.50000e-13*ic_cap*ic_cap+-1.00000e-13*ic_cap+4.96000e-11'
+ mcm5l1_cc_w_4_000_s_3_200 = '-1.06250e-13*ic_cap*ic_cap+-7.50000e-14*ic_cap+4.44000e-11'
+ mcm5l1_cc_w_4_000_s_4_800 = '-4.06250e-14*ic_cap*ic_cap+-3.75000e-14*ic_cap+3.15000e-11'
+ mcm5l1_cf_w_1_600_s_10_000 = '-1.37500e-13*ic_cap*ic_cap+-1.00000e-13*ic_cap+2.61000e-11'
+ mcm5l1_cf_w_1_600_s_12_000 = '-1.43750e-13*ic_cap*ic_cap+-1.00000e-13*ic_cap+2.84000e-11'
+ mcm5l1_cf_w_1_600_s_1_600 = '-2.40625e-14*ic_cap*ic_cap+-1.62500e-14*ic_cap+6.16000e-12'
+ mcm5l1_cf_w_1_600_s_1_700 = '-2.65625e-14*ic_cap*ic_cap+-1.87500e-14*ic_cap+6.52000e-12'
+ mcm5l1_cf_w_1_600_s_1_900 = '-3.18750e-14*ic_cap*ic_cap+-2.00000e-14*ic_cap+7.24000e-12'
+ mcm5l1_cf_w_1_600_s_2_000 = '-3.37500e-14*ic_cap*ic_cap+-2.25000e-14*ic_cap+7.59000e-12'
+ mcm5l1_cf_w_1_600_s_2_400 = '-4.37500e-14*ic_cap*ic_cap+-3.00000e-14*ic_cap+8.98000e-12'
+ mcm5l1_cf_w_1_600_s_2_800 = '-5.18750e-14*ic_cap*ic_cap+-3.50000e-14*ic_cap+1.03000e-11'
+ mcm5l1_cf_w_1_600_s_3_200 = '-5.93750e-14*ic_cap*ic_cap+-3.75000e-14*ic_cap+1.16000e-11'
+ mcm5l1_cf_w_1_600_s_4_800 = '-9.06250e-14*ic_cap*ic_cap+-6.25000e-14*ic_cap+1.62000e-11'
+ mcm5l1_cf_w_4_000_s_10_000 = '-1.34375e-13*ic_cap*ic_cap+-8.75000e-14*ic_cap+2.66000e-11'
+ mcm5l1_cf_w_4_000_s_12_000 = '-1.43750e-13*ic_cap*ic_cap+-1.00000e-13*ic_cap+2.91000e-11'
+ mcm5l1_cf_w_4_000_s_1_600 = '-2.40625e-14*ic_cap*ic_cap+-1.62500e-14*ic_cap+6.16000e-12'
+ mcm5l1_cf_w_4_000_s_1_700 = '-2.62500e-14*ic_cap*ic_cap+-1.75000e-14*ic_cap+6.53000e-12'
+ mcm5l1_cf_w_4_000_s_1_900 = '-3.18750e-14*ic_cap*ic_cap+-2.00000e-14*ic_cap+7.25000e-12'
+ mcm5l1_cf_w_4_000_s_2_000 = '-3.40625e-14*ic_cap*ic_cap+-2.12500e-14*ic_cap+7.60000e-12'
+ mcm5l1_cf_w_4_000_s_2_400 = '-4.43750e-14*ic_cap*ic_cap+-3.00000e-14*ic_cap+9.00000e-12'
+ mcm5l1_cf_w_4_000_s_2_800 = '-5.06250e-14*ic_cap*ic_cap+-3.50000e-14*ic_cap+1.03000e-11'
+ mcm5l1_cf_w_4_000_s_3_200 = '-5.93750e-14*ic_cap*ic_cap+-3.75000e-14*ic_cap+1.16000e-11'
+ mcm5l1_cf_w_4_000_s_4_800 = '-9.06250e-14*ic_cap*ic_cap+-6.25000e-14*ic_cap+1.63000e-11'
+ mcm5l1d_ca_w_0_170_s_0_180 = '-6.06250e-07*ic_cap*ic_cap+-3.50000e-07*ic_cap+6.33000e-05'
+ mcm5l1d_ca_w_0_170_s_0_225 = '-6.06250e-07*ic_cap*ic_cap+-3.50000e-07*ic_cap+6.33000e-05'
+ mcm5l1d_ca_w_0_170_s_0_270 = '-6.06250e-07*ic_cap*ic_cap+-3.50000e-07*ic_cap+6.33000e-05'
+ mcm5l1d_ca_w_0_170_s_0_360 = '-6.06250e-07*ic_cap*ic_cap+-3.50000e-07*ic_cap+6.33000e-05'
+ mcm5l1d_ca_w_0_170_s_0_450 = '-6.06250e-07*ic_cap*ic_cap+-3.50000e-07*ic_cap+6.33000e-05'
+ mcm5l1d_ca_w_0_170_s_0_540 = '-6.06250e-07*ic_cap*ic_cap+-3.50000e-07*ic_cap+6.33000e-05'
+ mcm5l1d_ca_w_0_170_s_0_720 = '-6.06250e-07*ic_cap*ic_cap+-3.50000e-07*ic_cap+6.33000e-05'
+ mcm5l1d_ca_w_0_170_s_1_080 = '-6.06250e-07*ic_cap*ic_cap+-3.50000e-07*ic_cap+6.33000e-05'
+ mcm5l1d_ca_w_0_170_s_1_980 = '-6.06250e-07*ic_cap*ic_cap+-3.50000e-07*ic_cap+6.33000e-05'
+ mcm5l1d_ca_w_0_170_s_4_500 = '-6.06250e-07*ic_cap*ic_cap+-3.50000e-07*ic_cap+6.33000e-05'
+ mcm5l1d_ca_w_1_360_s_0_180 = '-6.06250e-07*ic_cap*ic_cap+-3.50000e-07*ic_cap+6.33000e-05'
+ mcm5l1d_ca_w_1_360_s_0_225 = '-6.06250e-07*ic_cap*ic_cap+-3.50000e-07*ic_cap+6.33000e-05'
+ mcm5l1d_ca_w_1_360_s_0_270 = '-6.06250e-07*ic_cap*ic_cap+-3.50000e-07*ic_cap+6.33000e-05'
+ mcm5l1d_ca_w_1_360_s_0_360 = '-6.06250e-07*ic_cap*ic_cap+-3.50000e-07*ic_cap+6.33000e-05'
+ mcm5l1d_ca_w_1_360_s_0_450 = '-6.06250e-07*ic_cap*ic_cap+-3.50000e-07*ic_cap+6.33000e-05'
+ mcm5l1d_ca_w_1_360_s_0_540 = '-6.06250e-07*ic_cap*ic_cap+-3.50000e-07*ic_cap+6.33000e-05'
+ mcm5l1d_ca_w_1_360_s_0_720 = '-6.06250e-07*ic_cap*ic_cap+-3.50000e-07*ic_cap+6.33000e-05'
+ mcm5l1d_ca_w_1_360_s_1_080 = '-6.06250e-07*ic_cap*ic_cap+-3.50000e-07*ic_cap+6.33000e-05'
+ mcm5l1d_ca_w_1_360_s_1_980 = '-6.06250e-07*ic_cap*ic_cap+-3.50000e-07*ic_cap+6.33000e-05'
+ mcm5l1d_ca_w_1_360_s_4_500 = '-6.06250e-07*ic_cap*ic_cap+-3.50000e-07*ic_cap+6.33000e-05'
+ mcm5l1d_cc_w_0_170_s_0_180 = '-7.87500e-13*ic_cap*ic_cap+-5.00000e-13*ic_cap+7.65000e-11'
+ mcm5l1d_cc_w_0_170_s_0_225 = '-5.59375e-13*ic_cap*ic_cap+-3.87500e-13*ic_cap+6.45000e-11'
+ mcm5l1d_cc_w_0_170_s_0_270 = '-4.18750e-13*ic_cap*ic_cap+-3.00000e-13*ic_cap+5.64000e-11'
+ mcm5l1d_cc_w_0_170_s_0_360 = '-2.71875e-13*ic_cap*ic_cap+-1.87500e-13*ic_cap+4.49000e-11'
+ mcm5l1d_cc_w_0_170_s_0_450 = '-1.81250e-13*ic_cap*ic_cap+-1.50000e-13*ic_cap+3.77000e-11'
+ mcm5l1d_cc_w_0_170_s_0_540 = '-1.21875e-13*ic_cap*ic_cap+-1.12500e-13*ic_cap+3.18000e-11'
+ mcm5l1d_cc_w_0_170_s_0_720 = '-5.93750e-14*ic_cap*ic_cap+-6.25000e-14*ic_cap+2.41000e-11'
+ mcm5l1d_cc_w_0_170_s_1_080 = '-3.12500e-15*ic_cap*ic_cap+-1.25000e-14*ic_cap+1.51000e-11'
+ mcm5l1d_cc_w_0_170_s_1_980 = '2.84375e-14*ic_cap*ic_cap+1.12500e-14*ic_cap+5.84000e-12'
+ mcm5l1d_cc_w_0_170_s_4_500 = '1.26562e-14*ic_cap*ic_cap+8.12500e-15*ic_cap+7.85000e-13'
+ mcm5l1d_cc_w_1_360_s_0_180 = '-6.81250e-13*ic_cap*ic_cap+-4.50000e-13*ic_cap+9.23000e-11'
+ mcm5l1d_cc_w_1_360_s_0_225 = '-4.56250e-13*ic_cap*ic_cap+-3.00000e-13*ic_cap+7.91000e-11'
+ mcm5l1d_cc_w_1_360_s_0_270 = '-3.28125e-13*ic_cap*ic_cap+-2.37500e-13*ic_cap+6.98000e-11'
+ mcm5l1d_cc_w_1_360_s_0_360 = '-1.78125e-13*ic_cap*ic_cap+-1.37500e-13*ic_cap+5.68000e-11'
+ mcm5l1d_cc_w_1_360_s_0_450 = '-1.03125e-13*ic_cap*ic_cap+-8.75000e-14*ic_cap+4.81000e-11'
+ mcm5l1d_cc_w_1_360_s_0_540 = '-5.00000e-14*ic_cap*ic_cap+-5.00000e-14*ic_cap+4.16000e-11'
+ mcm5l1d_cc_w_1_360_s_0_720 = '3.12500e-15*ic_cap*ic_cap+-1.25000e-14*ic_cap+3.25000e-11'
+ mcm5l1d_cc_w_1_360_s_1_080 = '5.62500e-14*ic_cap*ic_cap+2.50000e-14*ic_cap+2.14000e-11'
+ mcm5l1d_cc_w_1_360_s_1_980 = '6.25000e-14*ic_cap*ic_cap+2.50000e-14*ic_cap+9.30000e-12'
+ mcm5l1d_cc_w_1_360_s_4_500 = '2.71875e-14*ic_cap*ic_cap+1.62500e-14*ic_cap+1.49000e-12'
+ mcm5l1d_cf_w_0_170_s_0_180 = '-6.87500e-15*ic_cap*ic_cap+-2.50000e-15*ic_cap+5.54000e-12'
+ mcm5l1d_cf_w_0_170_s_0_225 = '-1.96875e-14*ic_cap*ic_cap+-1.12500e-14*ic_cap+6.86000e-12'
+ mcm5l1d_cf_w_0_170_s_0_270 = '-3.28125e-14*ic_cap*ic_cap+-1.87500e-14*ic_cap+8.13000e-12'
+ mcm5l1d_cf_w_0_170_s_0_360 = '-5.78125e-14*ic_cap*ic_cap+-2.87500e-14*ic_cap+1.08000e-11'
+ mcm5l1d_cf_w_0_170_s_0_450 = '-7.81250e-14*ic_cap*ic_cap+-3.75000e-14*ic_cap+1.29000e-11'
+ mcm5l1d_cf_w_0_170_s_0_540 = '-1.03125e-13*ic_cap*ic_cap+-6.25000e-14*ic_cap+1.53000e-11'
+ mcm5l1d_cf_w_0_170_s_0_720 = '-1.31250e-13*ic_cap*ic_cap+-7.50000e-14*ic_cap+1.91000e-11'
+ mcm5l1d_cf_w_0_170_s_1_080 = '-1.78125e-13*ic_cap*ic_cap+-1.12500e-13*ic_cap+2.50000e-11'
+ mcm5l1d_cf_w_0_170_s_1_980 = '-2.09375e-13*ic_cap*ic_cap+-1.37500e-13*ic_cap+3.25000e-11'
+ mcm5l1d_cf_w_0_170_s_4_500 = '-1.96875e-13*ic_cap*ic_cap+-1.37500e-13*ic_cap+3.72000e-11'
+ mcm5l1d_cf_w_1_360_s_0_180 = '-6.87500e-15*ic_cap*ic_cap+-2.50000e-15*ic_cap+5.53000e-12'
+ mcm5l1d_cf_w_1_360_s_0_225 = '-2.00000e-14*ic_cap*ic_cap+-1.00000e-14*ic_cap+6.86000e-12'
+ mcm5l1d_cf_w_1_360_s_0_270 = '-3.21875e-14*ic_cap*ic_cap+-1.62500e-14*ic_cap+8.15000e-12'
+ mcm5l1d_cf_w_1_360_s_0_360 = '-5.34375e-14*ic_cap*ic_cap+-3.12500e-14*ic_cap+1.06000e-11'
+ mcm5l1d_cf_w_1_360_s_0_450 = '-7.81250e-14*ic_cap*ic_cap+-3.75000e-14*ic_cap+1.30000e-11'
+ mcm5l1d_cf_w_1_360_s_0_540 = '-9.68750e-14*ic_cap*ic_cap+-6.25000e-14*ic_cap+1.52000e-11'
+ mcm5l1d_cf_w_1_360_s_0_720 = '-1.31250e-13*ic_cap*ic_cap+-7.50000e-14*ic_cap+1.92000e-11'
+ mcm5l1d_cf_w_1_360_s_1_080 = '-1.68750e-13*ic_cap*ic_cap+-1.00000e-13*ic_cap+2.56000e-11'
+ mcm5l1d_cf_w_1_360_s_1_980 = '-2.00000e-13*ic_cap*ic_cap+-1.25000e-13*ic_cap+3.51000e-11'
+ mcm5l1d_cf_w_1_360_s_4_500 = '-1.71875e-13*ic_cap*ic_cap+-1.12500e-13*ic_cap+4.23000e-11'
+ mcm5l1f_ca_w_0_170_s_0_180 = '-4.68750e-07*ic_cap*ic_cap+-2.75000e-07*ic_cap+4.49000e-05'
+ mcm5l1f_ca_w_0_170_s_0_225 = '-4.68750e-07*ic_cap*ic_cap+-2.75000e-07*ic_cap+4.49000e-05'
+ mcm5l1f_ca_w_0_170_s_0_270 = '-4.68750e-07*ic_cap*ic_cap+-2.75000e-07*ic_cap+4.49000e-05'
+ mcm5l1f_ca_w_0_170_s_0_360 = '-4.68750e-07*ic_cap*ic_cap+-2.75000e-07*ic_cap+4.49000e-05'
+ mcm5l1f_ca_w_0_170_s_0_450 = '-4.68750e-07*ic_cap*ic_cap+-2.75000e-07*ic_cap+4.49000e-05'
+ mcm5l1f_ca_w_0_170_s_0_540 = '-4.68750e-07*ic_cap*ic_cap+-2.75000e-07*ic_cap+4.49000e-05'
+ mcm5l1f_ca_w_0_170_s_0_720 = '-4.68750e-07*ic_cap*ic_cap+-2.75000e-07*ic_cap+4.49000e-05'
+ mcm5l1f_ca_w_0_170_s_1_080 = '-4.68750e-07*ic_cap*ic_cap+-2.75000e-07*ic_cap+4.49000e-05'
+ mcm5l1f_ca_w_0_170_s_1_980 = '-4.68750e-07*ic_cap*ic_cap+-2.75000e-07*ic_cap+4.49000e-05'
+ mcm5l1f_ca_w_0_170_s_4_500 = '-4.68750e-07*ic_cap*ic_cap+-2.75000e-07*ic_cap+4.49000e-05'
+ mcm5l1f_ca_w_1_360_s_0_180 = '-4.68750e-07*ic_cap*ic_cap+-2.75000e-07*ic_cap+4.49000e-05'
+ mcm5l1f_ca_w_1_360_s_0_225 = '-4.68750e-07*ic_cap*ic_cap+-2.75000e-07*ic_cap+4.49000e-05'
+ mcm5l1f_ca_w_1_360_s_0_270 = '-4.68750e-07*ic_cap*ic_cap+-2.75000e-07*ic_cap+4.49000e-05'
+ mcm5l1f_ca_w_1_360_s_0_360 = '-4.68750e-07*ic_cap*ic_cap+-2.75000e-07*ic_cap+4.49000e-05'
+ mcm5l1f_ca_w_1_360_s_0_450 = '-4.68750e-07*ic_cap*ic_cap+-2.75000e-07*ic_cap+4.49000e-05'
+ mcm5l1f_ca_w_1_360_s_0_540 = '-4.68750e-07*ic_cap*ic_cap+-2.75000e-07*ic_cap+4.49000e-05'
+ mcm5l1f_ca_w_1_360_s_0_720 = '-4.68750e-07*ic_cap*ic_cap+-2.75000e-07*ic_cap+4.49000e-05'
+ mcm5l1f_ca_w_1_360_s_1_080 = '-4.68750e-07*ic_cap*ic_cap+-2.75000e-07*ic_cap+4.49000e-05'
+ mcm5l1f_ca_w_1_360_s_1_980 = '-4.68750e-07*ic_cap*ic_cap+-2.75000e-07*ic_cap+4.49000e-05'
+ mcm5l1f_ca_w_1_360_s_4_500 = '-4.68750e-07*ic_cap*ic_cap+-2.75000e-07*ic_cap+4.49000e-05'
+ mcm5l1f_cc_w_0_170_s_0_180 = '-7.84375e-13*ic_cap*ic_cap+-5.12500e-13*ic_cap+7.88000e-11'
+ mcm5l1f_cc_w_0_170_s_0_225 = '-5.81250e-13*ic_cap*ic_cap+-3.75000e-13*ic_cap+6.71000e-11'
+ mcm5l1f_cc_w_0_170_s_0_270 = '-4.31250e-13*ic_cap*ic_cap+-3.00000e-13*ic_cap+5.92000e-11'
+ mcm5l1f_cc_w_0_170_s_0_360 = '-2.87500e-13*ic_cap*ic_cap+-2.00000e-13*ic_cap+4.80000e-11'
+ mcm5l1f_cc_w_0_170_s_0_450 = '-1.90625e-13*ic_cap*ic_cap+-1.62500e-13*ic_cap+4.09000e-11'
+ mcm5l1f_cc_w_0_170_s_0_540 = '-1.34375e-13*ic_cap*ic_cap+-1.12500e-13*ic_cap+3.52000e-11'
+ mcm5l1f_cc_w_0_170_s_0_720 = '-6.87500e-14*ic_cap*ic_cap+-7.50000e-14*ic_cap+2.77000e-11'
+ mcm5l1f_cc_w_0_170_s_1_080 = '-2.50000e-14*ic_cap+1.85000e-11'
+ mcm5l1f_cc_w_0_170_s_1_980 = '4.50000e-14*ic_cap*ic_cap+2.00000e-14*ic_cap+8.13000e-12'
+ mcm5l1f_cc_w_0_170_s_4_500 = '2.34375e-14*ic_cap*ic_cap+1.62500e-14*ic_cap+1.29000e-12'
+ mcm5l1f_cc_w_1_360_s_0_180 = '-6.65625e-13*ic_cap*ic_cap+-4.12500e-13*ic_cap+9.67000e-11'
+ mcm5l1f_cc_w_1_360_s_0_225 = '-4.46875e-13*ic_cap*ic_cap+-2.87500e-13*ic_cap+8.35000e-11'
+ mcm5l1f_cc_w_1_360_s_0_270 = '-3.21875e-13*ic_cap*ic_cap+-2.37500e-13*ic_cap+7.42000e-11'
+ mcm5l1f_cc_w_1_360_s_0_360 = '-1.65625e-13*ic_cap*ic_cap+-1.37500e-13*ic_cap+6.12000e-11'
+ mcm5l1f_cc_w_1_360_s_0_450 = '-8.43750e-14*ic_cap*ic_cap+-8.75000e-14*ic_cap+5.24000e-11'
+ mcm5l1f_cc_w_1_360_s_0_540 = '-3.12500e-14*ic_cap*ic_cap+-5.00000e-14*ic_cap+4.59000e-11'
+ mcm5l1f_cc_w_1_360_s_0_720 = '2.50000e-14*ic_cap*ic_cap+3.67000e-11'
+ mcm5l1f_cc_w_1_360_s_1_080 = '7.81250e-14*ic_cap*ic_cap+3.75000e-14*ic_cap+2.53000e-11'
+ mcm5l1f_cc_w_1_360_s_1_980 = '9.06250e-14*ic_cap*ic_cap+6.25000e-14*ic_cap+1.20000e-11'
+ mcm5l1f_cc_w_1_360_s_4_500 = '4.65625e-14*ic_cap*ic_cap+3.12500e-14*ic_cap+2.14000e-12'
+ mcm5l1f_cf_w_0_170_s_0_180 = '-9.37500e-15*ic_cap*ic_cap+-5.00000e-15*ic_cap+3.98000e-12'
+ mcm5l1f_cf_w_0_170_s_0_225 = '-2.03125e-14*ic_cap*ic_cap+-8.75000e-15*ic_cap+4.94000e-12'
+ mcm5l1f_cf_w_0_170_s_0_270 = '-2.96875e-14*ic_cap*ic_cap+-1.87500e-14*ic_cap+5.86000e-12'
+ mcm5l1f_cf_w_0_170_s_0_360 = '-4.90625e-14*ic_cap*ic_cap+-2.62500e-14*ic_cap+7.86000e-12'
+ mcm5l1f_cf_w_0_170_s_0_450 = '-6.78125e-14*ic_cap*ic_cap+-3.87500e-14*ic_cap+9.44000e-12'
+ mcm5l1f_cf_w_0_170_s_0_540 = '-8.59375e-14*ic_cap*ic_cap+-4.37500e-14*ic_cap+1.13000e-11'
+ mcm5l1f_cf_w_0_170_s_0_720 = '-1.09375e-13*ic_cap*ic_cap+-6.25000e-14*ic_cap+1.43000e-11'
+ mcm5l1f_cf_w_0_170_s_1_080 = '-1.56250e-13*ic_cap*ic_cap+-1.00000e-13*ic_cap+1.94000e-11'
+ mcm5l1f_cf_w_0_170_s_1_980 = '-2.06250e-13*ic_cap*ic_cap+-1.25000e-13*ic_cap+2.70000e-11'
+ mcm5l1f_cf_w_0_170_s_4_500 = '-1.90625e-13*ic_cap*ic_cap+-1.37500e-13*ic_cap+3.31000e-11'
+ mcm5l1f_cf_w_1_360_s_0_180 = '-9.37500e-15*ic_cap*ic_cap+-5.00000e-15*ic_cap+3.97000e-12'
+ mcm5l1f_cf_w_1_360_s_0_225 = '-1.93750e-14*ic_cap*ic_cap+-1.00000e-14*ic_cap+4.93000e-12'
+ mcm5l1f_cf_w_1_360_s_0_270 = '-2.90625e-14*ic_cap*ic_cap+-1.62500e-14*ic_cap+5.87000e-12'
+ mcm5l1f_cf_w_1_360_s_0_360 = '-4.84375e-14*ic_cap*ic_cap+-2.87500e-14*ic_cap+7.72000e-12'
+ mcm5l1f_cf_w_1_360_s_0_450 = '-6.68750e-14*ic_cap*ic_cap+-3.75000e-14*ic_cap+9.51000e-12'
+ mcm5l1f_cf_w_1_360_s_0_540 = '-8.15625e-14*ic_cap*ic_cap+-5.12500e-14*ic_cap+1.12000e-11'
+ mcm5l1f_cf_w_1_360_s_0_720 = '-1.15625e-13*ic_cap*ic_cap+-6.25000e-14*ic_cap+1.44000e-11'
+ mcm5l1f_cf_w_1_360_s_1_080 = '-1.56250e-13*ic_cap*ic_cap+-1.00000e-13*ic_cap+1.98000e-11'
+ mcm5l1f_cf_w_1_360_s_1_980 = '-2.06250e-13*ic_cap*ic_cap+-1.25000e-13*ic_cap+2.90000e-11'
+ mcm5l1f_cf_w_1_360_s_4_500 = '-1.75000e-13*ic_cap*ic_cap+-1.00000e-13*ic_cap+3.76000e-11'
+ mcm5l1p1_ca_w_0_170_s_0_180 = '-1.70000e-06*ic_cap*ic_cap+-8.25000e-07*ic_cap+1.02000e-04'
+ mcm5l1p1_ca_w_0_170_s_0_225 = '-1.70000e-06*ic_cap*ic_cap+-8.25000e-07*ic_cap+1.02000e-04'
+ mcm5l1p1_ca_w_0_170_s_0_270 = '-1.70000e-06*ic_cap*ic_cap+-8.25000e-07*ic_cap+1.02000e-04'
+ mcm5l1p1_ca_w_0_170_s_0_360 = '-1.70000e-06*ic_cap*ic_cap+-8.25000e-07*ic_cap+1.02000e-04'
+ mcm5l1p1_ca_w_0_170_s_0_450 = '-1.70000e-06*ic_cap*ic_cap+-8.25000e-07*ic_cap+1.02000e-04'
+ mcm5l1p1_ca_w_0_170_s_0_540 = '-1.70000e-06*ic_cap*ic_cap+-8.25000e-07*ic_cap+1.02000e-04'
+ mcm5l1p1_ca_w_0_170_s_0_720 = '-1.70000e-06*ic_cap*ic_cap+-8.25000e-07*ic_cap+1.02000e-04'
+ mcm5l1p1_ca_w_0_170_s_1_080 = '-1.70000e-06*ic_cap*ic_cap+-8.25000e-07*ic_cap+1.02000e-04'
+ mcm5l1p1_ca_w_0_170_s_1_980 = '-1.70000e-06*ic_cap*ic_cap+-8.25000e-07*ic_cap+1.02000e-04'
+ mcm5l1p1_ca_w_0_170_s_4_500 = '-1.70000e-06*ic_cap*ic_cap+-8.25000e-07*ic_cap+1.02000e-04'
+ mcm5l1p1_ca_w_1_360_s_0_180 = '-1.70000e-06*ic_cap*ic_cap+-8.25000e-07*ic_cap+1.02000e-04'
+ mcm5l1p1_ca_w_1_360_s_0_225 = '-1.70000e-06*ic_cap*ic_cap+-8.25000e-07*ic_cap+1.02000e-04'
+ mcm5l1p1_ca_w_1_360_s_0_270 = '-1.70000e-06*ic_cap*ic_cap+-8.25000e-07*ic_cap+1.02000e-04'
+ mcm5l1p1_ca_w_1_360_s_0_360 = '-1.70000e-06*ic_cap*ic_cap+-8.25000e-07*ic_cap+1.02000e-04'
+ mcm5l1p1_ca_w_1_360_s_0_450 = '-1.70000e-06*ic_cap*ic_cap+-8.25000e-07*ic_cap+1.02000e-04'
+ mcm5l1p1_ca_w_1_360_s_0_540 = '-1.70000e-06*ic_cap*ic_cap+-8.25000e-07*ic_cap+1.02000e-04'
+ mcm5l1p1_ca_w_1_360_s_0_720 = '-1.70000e-06*ic_cap*ic_cap+-8.25000e-07*ic_cap+1.02000e-04'
+ mcm5l1p1_ca_w_1_360_s_1_080 = '-1.70000e-06*ic_cap*ic_cap+-8.25000e-07*ic_cap+1.02000e-04'
+ mcm5l1p1_ca_w_1_360_s_1_980 = '-1.70000e-06*ic_cap*ic_cap+-8.25000e-07*ic_cap+1.02000e-04'
+ mcm5l1p1_ca_w_1_360_s_4_500 = '-1.70000e-06*ic_cap*ic_cap+-8.25000e-07*ic_cap+1.02000e-04'
+ mcm5l1p1_cc_w_0_170_s_0_180 = '-6.71875e-13*ic_cap*ic_cap+-4.62500e-13*ic_cap+7.21000e-11'
+ mcm5l1p1_cc_w_0_170_s_0_225 = '-4.56250e-13*ic_cap*ic_cap+-3.25000e-13*ic_cap+6.01000e-11'
+ mcm5l1p1_cc_w_0_170_s_0_270 = '-3.09375e-13*ic_cap*ic_cap+-2.37500e-13*ic_cap+5.17000e-11'
+ mcm5l1p1_cc_w_0_170_s_0_360 = '-1.59375e-13*ic_cap*ic_cap+-1.37500e-13*ic_cap+4.00000e-11'
+ mcm5l1p1_cc_w_0_170_s_0_450 = '-7.18750e-14*ic_cap*ic_cap+-8.75000e-14*ic_cap+3.27000e-11'
+ mcm5l1p1_cc_w_0_170_s_0_540 = '-1.87500e-14*ic_cap*ic_cap+-5.00000e-14*ic_cap+2.68000e-11'
+ mcm5l1p1_cc_w_0_170_s_0_720 = '3.75000e-14*ic_cap*ic_cap+1.92000e-11'
+ mcm5l1p1_cc_w_0_170_s_1_080 = '6.87500e-14*ic_cap*ic_cap+2.50000e-14*ic_cap+1.09000e-11'
+ mcm5l1p1_cc_w_0_170_s_1_980 = '5.50000e-14*ic_cap*ic_cap+2.75000e-14*ic_cap+3.61000e-12'
+ mcm5l1p1_cc_w_0_170_s_4_500 = '1.14062e-14*ic_cap*ic_cap+8.37500e-15*ic_cap+4.47000e-13'
+ mcm5l1p1_cc_w_1_360_s_0_180 = '-5.62500e-13*ic_cap*ic_cap+-3.75000e-13*ic_cap+8.63000e-11'
+ mcm5l1p1_cc_w_1_360_s_0_225 = '-3.59375e-13*ic_cap*ic_cap+-2.62500e-13*ic_cap+7.34000e-11'
+ mcm5l1p1_cc_w_1_360_s_0_270 = '-2.21875e-13*ic_cap*ic_cap+-1.87500e-13*ic_cap+6.39000e-11'
+ mcm5l1p1_cc_w_1_360_s_0_360 = '-7.81250e-14*ic_cap*ic_cap+-8.75000e-14*ic_cap+5.11000e-11'
+ mcm5l1p1_cc_w_1_360_s_0_450 = '3.12500e-15*ic_cap*ic_cap+-3.75000e-14*ic_cap+4.24000e-11'
+ mcm5l1p1_cc_w_1_360_s_0_540 = '5.00000e-14*ic_cap*ic_cap+3.60000e-11'
+ mcm5l1p1_cc_w_1_360_s_0_720 = '9.68750e-14*ic_cap*ic_cap+3.75000e-14*ic_cap+2.72000e-11'
+ mcm5l1p1_cc_w_1_360_s_1_080 = '1.21875e-13*ic_cap*ic_cap+6.25000e-14*ic_cap+1.70000e-11'
+ mcm5l1p1_cc_w_1_360_s_1_980 = '9.31250e-14*ic_cap*ic_cap+5.75000e-14*ic_cap+6.69000e-12'
+ mcm5l1p1_cc_w_1_360_s_4_500 = '2.62500e-14*ic_cap*ic_cap+1.62500e-14*ic_cap+9.85000e-13'
+ mcm5l1p1_cf_w_0_170_s_0_180 = '-8.12500e-14*ic_cap*ic_cap+-3.75000e-14*ic_cap+8.78000e-12'
+ mcm5l1p1_cf_w_0_170_s_0_225 = '-1.14687e-13*ic_cap*ic_cap+-5.62500e-14*ic_cap+1.08000e-11'
+ mcm5l1p1_cf_w_0_170_s_0_270 = '-1.43750e-13*ic_cap*ic_cap+-7.50000e-14*ic_cap+1.27000e-11'
+ mcm5l1p1_cf_w_0_170_s_0_360 = '-2.00000e-13*ic_cap*ic_cap+-1.00000e-13*ic_cap+1.66000e-11'
+ mcm5l1p1_cf_w_0_170_s_0_450 = '-2.50000e-13*ic_cap*ic_cap+-1.25000e-13*ic_cap+1.96000e-11'
+ mcm5l1p1_cf_w_0_170_s_0_540 = '-2.87500e-13*ic_cap*ic_cap+-1.50000e-13*ic_cap+2.28000e-11'
+ mcm5l1p1_cf_w_0_170_s_0_720 = '-3.43750e-13*ic_cap*ic_cap+-1.75000e-13*ic_cap+2.76000e-11'
+ mcm5l1p1_cf_w_0_170_s_1_080 = '-3.90625e-13*ic_cap*ic_cap+-2.12500e-13*ic_cap+3.40000e-11'
+ mcm5l1p1_cf_w_0_170_s_1_980 = '-3.87500e-13*ic_cap*ic_cap+-2.25000e-13*ic_cap+4.05000e-11'
+ mcm5l1p1_cf_w_0_170_s_4_500 = '-3.46875e-13*ic_cap*ic_cap+-2.12500e-13*ic_cap+4.35000e-11'
+ mcm5l1p1_cf_w_1_360_s_0_180 = '-8.31250e-14*ic_cap*ic_cap+-4.00000e-14*ic_cap+8.86000e-12'
+ mcm5l1p1_cf_w_1_360_s_0_225 = '-1.16875e-13*ic_cap*ic_cap+-5.50000e-14*ic_cap+1.09000e-11'
+ mcm5l1p1_cf_w_1_360_s_0_270 = '-1.43750e-13*ic_cap*ic_cap+-7.50000e-14*ic_cap+1.28000e-11'
+ mcm5l1p1_cf_w_1_360_s_0_360 = '-2.00000e-13*ic_cap*ic_cap+-1.00000e-13*ic_cap+1.65000e-11'
+ mcm5l1p1_cf_w_1_360_s_0_450 = '-2.43750e-13*ic_cap*ic_cap+-1.25000e-13*ic_cap+1.98000e-11'
+ mcm5l1p1_cf_w_1_360_s_0_540 = '-2.84375e-13*ic_cap*ic_cap+-1.37500e-13*ic_cap+2.28000e-11'
+ mcm5l1p1_cf_w_1_360_s_0_720 = '-3.37500e-13*ic_cap*ic_cap+-1.75000e-13*ic_cap+2.79000e-11'
+ mcm5l1p1_cf_w_1_360_s_1_080 = '-3.96875e-13*ic_cap*ic_cap+-2.12500e-13*ic_cap+3.53000e-11'
+ mcm5l1p1_cf_w_1_360_s_1_980 = '-3.93750e-13*ic_cap*ic_cap+-2.25000e-13*ic_cap+4.41000e-11'
+ mcm5l1p1_cf_w_1_360_s_4_500 = '-3.37500e-13*ic_cap*ic_cap+-2.00000e-13*ic_cap+4.96000e-11'
+ mcm5m1_ca_w_1_600_s_10_000 = '-6.71875e-08*ic_cap*ic_cap+-4.12500e-08*ic_cap+9.50000e-06'
+ mcm5m1_ca_w_1_600_s_12_000 = '-6.71875e-08*ic_cap*ic_cap+-4.12500e-08*ic_cap+9.50000e-06'
+ mcm5m1_ca_w_1_600_s_1_600 = '-6.71875e-08*ic_cap*ic_cap+-4.12500e-08*ic_cap+9.50000e-06'
+ mcm5m1_ca_w_1_600_s_1_700 = '-6.71875e-08*ic_cap*ic_cap+-4.12500e-08*ic_cap+9.50000e-06'
+ mcm5m1_ca_w_1_600_s_1_900 = '-6.71875e-08*ic_cap*ic_cap+-4.12500e-08*ic_cap+9.50000e-06'
+ mcm5m1_ca_w_1_600_s_2_000 = '-6.71875e-08*ic_cap*ic_cap+-4.12500e-08*ic_cap+9.50000e-06'
+ mcm5m1_ca_w_1_600_s_2_400 = '-6.71875e-08*ic_cap*ic_cap+-4.12500e-08*ic_cap+9.50000e-06'
+ mcm5m1_ca_w_1_600_s_2_800 = '-6.71875e-08*ic_cap*ic_cap+-4.12500e-08*ic_cap+9.50000e-06'
+ mcm5m1_ca_w_1_600_s_3_200 = '-6.71875e-08*ic_cap*ic_cap+-4.12500e-08*ic_cap+9.50000e-06'
+ mcm5m1_ca_w_1_600_s_4_800 = '-6.71875e-08*ic_cap*ic_cap+-4.12500e-08*ic_cap+9.50000e-06'
+ mcm5m1_ca_w_4_000_s_10_000 = '-6.71875e-08*ic_cap*ic_cap+-4.12500e-08*ic_cap+9.50000e-06'
+ mcm5m1_ca_w_4_000_s_12_000 = '-6.71875e-08*ic_cap*ic_cap+-4.12500e-08*ic_cap+9.50000e-06'
+ mcm5m1_ca_w_4_000_s_1_600 = '-6.71875e-08*ic_cap*ic_cap+-4.12500e-08*ic_cap+9.50000e-06'
+ mcm5m1_ca_w_4_000_s_1_700 = '-6.71875e-08*ic_cap*ic_cap+-4.12500e-08*ic_cap+9.50000e-06'
+ mcm5m1_ca_w_4_000_s_1_900 = '-6.71875e-08*ic_cap*ic_cap+-4.12500e-08*ic_cap+9.50000e-06'
+ mcm5m1_ca_w_4_000_s_2_000 = '-6.71875e-08*ic_cap*ic_cap+-4.12500e-08*ic_cap+9.50000e-06'
+ mcm5m1_ca_w_4_000_s_2_400 = '-6.71875e-08*ic_cap*ic_cap+-4.12500e-08*ic_cap+9.50000e-06'
+ mcm5m1_ca_w_4_000_s_2_800 = '-6.71875e-08*ic_cap*ic_cap+-4.12500e-08*ic_cap+9.50000e-06'
+ mcm5m1_ca_w_4_000_s_3_200 = '-6.71875e-08*ic_cap*ic_cap+-4.12500e-08*ic_cap+9.50000e-06'
+ mcm5m1_ca_w_4_000_s_4_800 = '-6.71875e-08*ic_cap*ic_cap+-4.12500e-08*ic_cap+9.50000e-06'
+ mcm5m1_cc_w_1_600_s_10_000 = '6.25000e-15*ic_cap*ic_cap+1.10000e-11'
+ mcm5m1_cc_w_1_600_s_12_000 = '8.12500e-15*ic_cap*ic_cap+5.00000e-15*ic_cap+8.51000e-12'
+ mcm5m1_cc_w_1_600_s_1_600 = '-4.53125e-13*ic_cap*ic_cap+-3.12500e-13*ic_cap+7.04000e-11'
+ mcm5m1_cc_w_1_600_s_1_700 = '-4.12500e-13*ic_cap*ic_cap+-2.75000e-13*ic_cap+6.68000e-11'
+ mcm5m1_cc_w_1_600_s_1_900 = '-3.37500e-13*ic_cap*ic_cap+-2.25000e-13*ic_cap+6.05000e-11'
+ mcm5m1_cc_w_1_600_s_2_000 = '-3.06250e-13*ic_cap*ic_cap+-2.25000e-13*ic_cap+5.79000e-11'
+ mcm5m1_cc_w_1_600_s_2_400 = '-2.18750e-13*ic_cap*ic_cap+-1.50000e-13*ic_cap+4.94000e-11'
+ mcm5m1_cc_w_1_600_s_2_800 = '-1.68750e-13*ic_cap*ic_cap+-1.25000e-13*ic_cap+4.32000e-11'
+ mcm5m1_cc_w_1_600_s_3_200 = '-1.34375e-13*ic_cap*ic_cap+-8.75000e-14*ic_cap+3.84000e-11'
+ mcm5m1_cc_w_1_600_s_4_800 = '-5.00000e-14*ic_cap*ic_cap+-5.00000e-14*ic_cap+2.61000e-11'
+ mcm5m1_cc_w_4_000_s_10_000 = '9.37500e-15*ic_cap*ic_cap+1.25000e-14*ic_cap+1.35000e-11'
+ mcm5m1_cc_w_4_000_s_12_000 = '9.37500e-15*ic_cap*ic_cap+1.25000e-14*ic_cap+1.07000e-11'
+ mcm5m1_cc_w_4_000_s_1_600 = '-4.34375e-13*ic_cap*ic_cap+-2.87500e-13*ic_cap+7.66000e-11'
+ mcm5m1_cc_w_4_000_s_1_700 = '-3.87500e-13*ic_cap*ic_cap+-2.50000e-13*ic_cap+7.27000e-11'
+ mcm5m1_cc_w_4_000_s_1_900 = '-3.06250e-13*ic_cap*ic_cap+-2.00000e-13*ic_cap+6.61000e-11'
+ mcm5m1_cc_w_4_000_s_2_000 = '-2.81250e-13*ic_cap*ic_cap+-2.00000e-13*ic_cap+6.33000e-11'
+ mcm5m1_cc_w_4_000_s_2_400 = '-2.03125e-13*ic_cap*ic_cap+-1.37500e-13*ic_cap+5.45000e-11'
+ mcm5m1_cc_w_4_000_s_2_800 = '-1.43750e-13*ic_cap*ic_cap+-1.00000e-13*ic_cap+4.78000e-11'
+ mcm5m1_cc_w_4_000_s_3_200 = '-1.06250e-13*ic_cap*ic_cap+-7.50000e-14*ic_cap+4.27000e-11'
+ mcm5m1_cc_w_4_000_s_4_800 = '-4.06250e-14*ic_cap*ic_cap+-3.75000e-14*ic_cap+2.98000e-11'
+ mcm5m1_cf_w_1_600_s_10_000 = '-1.50000e-13*ic_cap*ic_cap+-1.00000e-13*ic_cap+2.90000e-11'
+ mcm5m1_cf_w_1_600_s_12_000 = '-1.50000e-13*ic_cap*ic_cap+-1.00000e-13*ic_cap+3.11000e-11'
+ mcm5m1_cf_w_1_600_s_1_600 = '-2.68750e-14*ic_cap*ic_cap+-1.75000e-14*ic_cap+7.21000e-12'
+ mcm5m1_cf_w_1_600_s_1_700 = '-3.03125e-14*ic_cap*ic_cap+-1.87500e-14*ic_cap+7.63000e-12'
+ mcm5m1_cf_w_1_600_s_1_900 = '-3.65625e-14*ic_cap*ic_cap+-2.12500e-14*ic_cap+8.47000e-12'
+ mcm5m1_cf_w_1_600_s_2_000 = '-3.90625e-14*ic_cap*ic_cap+-2.37500e-14*ic_cap+8.88000e-12'
+ mcm5m1_cf_w_1_600_s_2_400 = '-5.15625e-14*ic_cap*ic_cap+-3.12500e-14*ic_cap+1.05000e-11'
+ mcm5m1_cf_w_1_600_s_2_800 = '-5.93750e-14*ic_cap*ic_cap+-3.75000e-14*ic_cap+1.20000e-11'
+ mcm5m1_cf_w_1_600_s_3_200 = '-7.18750e-14*ic_cap*ic_cap+-3.75000e-14*ic_cap+1.35000e-11'
+ mcm5m1_cf_w_1_600_s_4_800 = '-1.03125e-13*ic_cap*ic_cap+-6.25000e-14*ic_cap+1.86000e-11'
+ mcm5m1_cf_w_4_000_s_10_000 = '-1.43750e-13*ic_cap*ic_cap+-1.00000e-13*ic_cap+2.95000e-11'
+ mcm5m1_cf_w_4_000_s_12_000 = '-1.46875e-13*ic_cap*ic_cap+-8.75000e-14*ic_cap+3.19000e-11'
+ mcm5m1_cf_w_4_000_s_1_600 = '-2.75000e-14*ic_cap*ic_cap+-1.75000e-14*ic_cap+7.22000e-12'
+ mcm5m1_cf_w_4_000_s_1_700 = '-2.96875e-14*ic_cap*ic_cap+-1.62500e-14*ic_cap+7.64000e-12'
+ mcm5m1_cf_w_4_000_s_1_900 = '-3.53125e-14*ic_cap*ic_cap+-2.12500e-14*ic_cap+8.47000e-12'
+ mcm5m1_cf_w_4_000_s_2_000 = '-3.84375e-14*ic_cap*ic_cap+-2.37500e-14*ic_cap+8.88000e-12'
+ mcm5m1_cf_w_4_000_s_2_400 = '-5.06250e-14*ic_cap*ic_cap+-3.25000e-14*ic_cap+1.05000e-11'
+ mcm5m1_cf_w_4_000_s_2_800 = '-5.93750e-14*ic_cap*ic_cap+-3.75000e-14*ic_cap+1.20000e-11'
+ mcm5m1_cf_w_4_000_s_3_200 = '-6.87500e-14*ic_cap*ic_cap+-5.00000e-14*ic_cap+1.35000e-11'
+ mcm5m1_cf_w_4_000_s_4_800 = '-1.03125e-13*ic_cap*ic_cap+-6.25000e-14*ic_cap+1.87000e-11'
+ mcm5m1d_ca_w_0_140_s_0_140 = '-4.40625e-07*ic_cap*ic_cap+-2.87500e-07*ic_cap+4.31000e-05'
+ mcm5m1d_ca_w_0_140_s_0_175 = '-4.40625e-07*ic_cap*ic_cap+-2.87500e-07*ic_cap+4.31000e-05'
+ mcm5m1d_ca_w_0_140_s_0_210 = '-4.40625e-07*ic_cap*ic_cap+-2.87500e-07*ic_cap+4.31000e-05'
+ mcm5m1d_ca_w_0_140_s_0_280 = '-4.40625e-07*ic_cap*ic_cap+-2.87500e-07*ic_cap+4.31000e-05'
+ mcm5m1d_ca_w_0_140_s_0_350 = '-4.40625e-07*ic_cap*ic_cap+-2.87500e-07*ic_cap+4.31000e-05'
+ mcm5m1d_ca_w_0_140_s_0_420 = '-4.40625e-07*ic_cap*ic_cap+-2.87500e-07*ic_cap+4.31000e-05'
+ mcm5m1d_ca_w_0_140_s_0_560 = '-4.40625e-07*ic_cap*ic_cap+-2.87500e-07*ic_cap+4.31000e-05'
+ mcm5m1d_ca_w_0_140_s_0_840 = '-4.40625e-07*ic_cap*ic_cap+-2.87500e-07*ic_cap+4.31000e-05'
+ mcm5m1d_ca_w_0_140_s_1_540 = '-4.40625e-07*ic_cap*ic_cap+-2.87500e-07*ic_cap+4.31000e-05'
+ mcm5m1d_ca_w_0_140_s_3_500 = '-4.40625e-07*ic_cap*ic_cap+-2.87500e-07*ic_cap+4.31000e-05'
+ mcm5m1d_ca_w_1_120_s_0_140 = '-4.40625e-07*ic_cap*ic_cap+-2.87500e-07*ic_cap+4.31000e-05'
+ mcm5m1d_ca_w_1_120_s_0_175 = '-4.40625e-07*ic_cap*ic_cap+-2.87500e-07*ic_cap+4.31000e-05'
+ mcm5m1d_ca_w_1_120_s_0_210 = '-4.40625e-07*ic_cap*ic_cap+-2.87500e-07*ic_cap+4.31000e-05'
+ mcm5m1d_ca_w_1_120_s_0_280 = '-4.40625e-07*ic_cap*ic_cap+-2.87500e-07*ic_cap+4.31000e-05'
+ mcm5m1d_ca_w_1_120_s_0_350 = '-4.40625e-07*ic_cap*ic_cap+-2.87500e-07*ic_cap+4.31000e-05'
+ mcm5m1d_ca_w_1_120_s_0_420 = '-4.40625e-07*ic_cap*ic_cap+-2.87500e-07*ic_cap+4.31000e-05'
+ mcm5m1d_ca_w_1_120_s_0_560 = '-4.40625e-07*ic_cap*ic_cap+-2.87500e-07*ic_cap+4.31000e-05'
+ mcm5m1d_ca_w_1_120_s_0_840 = '-4.40625e-07*ic_cap*ic_cap+-2.87500e-07*ic_cap+4.31000e-05'
+ mcm5m1d_ca_w_1_120_s_1_540 = '-4.40625e-07*ic_cap*ic_cap+-2.87500e-07*ic_cap+4.31000e-05'
+ mcm5m1d_ca_w_1_120_s_3_500 = '-4.40625e-07*ic_cap*ic_cap+-2.87500e-07*ic_cap+4.31000e-05'
+ mcm5m1d_cc_w_0_140_s_0_140 = '-9.12500e-13*ic_cap*ic_cap+-5.25000e-13*ic_cap+1.03000e-10'
+ mcm5m1d_cc_w_0_140_s_0_175 = '-8.37500e-13*ic_cap*ic_cap+-6.00000e-13*ic_cap+1.01000e-10'
+ mcm5m1d_cc_w_0_140_s_0_210 = '-7.50000e-13*ic_cap*ic_cap+-4.25000e-13*ic_cap+9.56000e-11'
+ mcm5m1d_cc_w_0_140_s_0_280 = '-5.71875e-13*ic_cap*ic_cap+-3.62500e-13*ic_cap+8.45000e-11'
+ mcm5m1d_cc_w_0_140_s_0_350 = '-4.18750e-13*ic_cap*ic_cap+-2.25000e-13*ic_cap+7.26000e-11'
+ mcm5m1d_cc_w_0_140_s_0_420 = '-3.12500e-13*ic_cap*ic_cap+-2.50000e-13*ic_cap+6.30000e-11'
+ mcm5m1d_cc_w_0_140_s_0_560 = '-1.90625e-13*ic_cap*ic_cap+-1.12500e-13*ic_cap+5.00000e-11'
+ mcm5m1d_cc_w_0_140_s_0_840 = '-5.62500e-14*ic_cap*ic_cap+-5.00000e-14*ic_cap+3.48000e-11'
+ mcm5m1d_cc_w_0_140_s_1_540 = '3.75000e-14*ic_cap*ic_cap+2.50000e-14*ic_cap+1.75000e-11'
+ mcm5m1d_cc_w_0_140_s_3_500 = '4.53125e-14*ic_cap*ic_cap+3.37500e-14*ic_cap+3.87000e-12'
+ mcm5m1d_cc_w_1_120_s_0_140 = '-8.12500e-13*ic_cap*ic_cap+-5.00000e-13*ic_cap+1.23000e-10'
+ mcm5m1d_cc_w_1_120_s_0_175 = '-8.12500e-13*ic_cap*ic_cap+-2.50000e-13*ic_cap+1.20000e-10'
+ mcm5m1d_cc_w_1_120_s_0_210 = '-6.25000e-13*ic_cap*ic_cap+-5.00000e-13*ic_cap+1.13000e-10'
+ mcm5m1d_cc_w_1_120_s_0_280 = '-4.59375e-13*ic_cap*ic_cap+-3.12500e-13*ic_cap+9.88000e-11'
+ mcm5m1d_cc_w_1_120_s_0_350 = '-3.59375e-13*ic_cap*ic_cap+-2.62500e-13*ic_cap+8.63000e-11'
+ mcm5m1d_cc_w_1_120_s_0_420 = '-2.25000e-13*ic_cap*ic_cap+-1.75000e-13*ic_cap+7.51000e-11'
+ mcm5m1d_cc_w_1_120_s_0_560 = '-1.06250e-13*ic_cap*ic_cap+-7.50000e-14*ic_cap+5.97000e-11'
+ mcm5m1d_cc_w_1_120_s_0_840 = '1.25000e-14*ic_cap*ic_cap+4.17000e-11'
+ mcm5m1d_cc_w_1_120_s_1_540 = '8.43750e-14*ic_cap*ic_cap+6.25000e-14*ic_cap+2.17000e-11'
+ mcm5m1d_cc_w_1_120_s_3_500 = '6.78125e-14*ic_cap*ic_cap+5.12500e-14*ic_cap+5.18000e-12'
+ mcm5m1d_cf_w_0_140_s_0_140 = '-2.18750e-15*ic_cap*ic_cap+-3.75000e-15*ic_cap+2.99000e-12'
+ mcm5m1d_cf_w_0_140_s_0_175 = '-9.37500e-15*ic_cap*ic_cap+-7.50000e-15*ic_cap+3.73000e-12'
+ mcm5m1d_cf_w_0_140_s_0_210 = '-1.68750e-14*ic_cap*ic_cap+-1.25000e-14*ic_cap+4.49000e-12'
+ mcm5m1d_cf_w_0_140_s_0_280 = '-3.25000e-14*ic_cap*ic_cap+-2.00000e-14*ic_cap+5.95000e-12'
+ mcm5m1d_cf_w_0_140_s_0_350 = '-4.75000e-14*ic_cap*ic_cap+-3.00000e-14*ic_cap+7.38000e-12'
+ mcm5m1d_cf_w_0_140_s_0_420 = '-6.06250e-14*ic_cap*ic_cap+-4.25000e-14*ic_cap+8.82000e-12'
+ mcm5m1d_cf_w_0_140_s_0_560 = '-8.81250e-14*ic_cap*ic_cap+-5.25000e-14*ic_cap+1.15000e-11'
+ mcm5m1d_cf_w_0_140_s_0_840 = '-1.34375e-13*ic_cap*ic_cap+-8.75000e-14*ic_cap+1.64000e-11'
+ mcm5m1d_cf_w_0_140_s_1_540 = '-2.03125e-13*ic_cap*ic_cap+-1.37500e-13*ic_cap+2.56000e-11'
+ mcm5m1d_cf_w_0_140_s_3_500 = '-2.31250e-13*ic_cap*ic_cap+-1.50000e-13*ic_cap+3.66000e-11'
+ mcm5m1d_cf_w_1_120_s_0_140 = '-3.12500e-15*ic_cap*ic_cap+-2.50000e-15*ic_cap+3.06000e-12'
+ mcm5m1d_cf_w_1_120_s_0_175 = '-1.03125e-14*ic_cap*ic_cap+-6.25000e-15*ic_cap+3.80000e-12'
+ mcm5m1d_cf_w_1_120_s_0_210 = '-1.90625e-14*ic_cap*ic_cap+-1.37500e-14*ic_cap+4.55000e-12'
+ mcm5m1d_cf_w_1_120_s_0_280 = '-3.28125e-14*ic_cap*ic_cap+-2.12500e-14*ic_cap+6.01000e-12'
+ mcm5m1d_cf_w_1_120_s_0_350 = '-4.75000e-14*ic_cap*ic_cap+-3.25000e-14*ic_cap+7.45000e-12'
+ mcm5m1d_cf_w_1_120_s_0_420 = '-6.15625e-14*ic_cap*ic_cap+-4.12500e-14*ic_cap+8.86000e-12'
+ mcm5m1d_cf_w_1_120_s_0_560 = '-8.96875e-14*ic_cap*ic_cap+-5.87500e-14*ic_cap+1.16000e-11'
+ mcm5m1d_cf_w_1_120_s_0_840 = '-1.34375e-13*ic_cap*ic_cap+-8.75000e-14*ic_cap+1.66000e-11'
+ mcm5m1d_cf_w_1_120_s_1_540 = '-2.03125e-13*ic_cap*ic_cap+-1.37500e-13*ic_cap+2.63000e-11'
+ mcm5m1d_cf_w_1_120_s_3_500 = '-2.31250e-13*ic_cap*ic_cap+-1.50000e-13*ic_cap+3.92000e-11'
+ mcm5m1f_ca_w_0_140_s_0_140 = '-3.68750e-07*ic_cap*ic_cap+-2.25000e-07*ic_cap+3.53000e-05'
+ mcm5m1f_ca_w_0_140_s_0_175 = '-3.68750e-07*ic_cap*ic_cap+-2.25000e-07*ic_cap+3.53000e-05'
+ mcm5m1f_ca_w_0_140_s_0_210 = '-3.68750e-07*ic_cap*ic_cap+-2.25000e-07*ic_cap+3.53000e-05'
+ mcm5m1f_ca_w_0_140_s_0_280 = '-3.68750e-07*ic_cap*ic_cap+-2.25000e-07*ic_cap+3.53000e-05'
+ mcm5m1f_ca_w_0_140_s_0_350 = '-3.68750e-07*ic_cap*ic_cap+-2.25000e-07*ic_cap+3.53000e-05'
+ mcm5m1f_ca_w_0_140_s_0_420 = '-3.68750e-07*ic_cap*ic_cap+-2.25000e-07*ic_cap+3.53000e-05'
+ mcm5m1f_ca_w_0_140_s_0_560 = '-3.68750e-07*ic_cap*ic_cap+-2.25000e-07*ic_cap+3.53000e-05'
+ mcm5m1f_ca_w_0_140_s_0_840 = '-3.68750e-07*ic_cap*ic_cap+-2.25000e-07*ic_cap+3.53000e-05'
+ mcm5m1f_ca_w_0_140_s_1_540 = '-3.68750e-07*ic_cap*ic_cap+-2.25000e-07*ic_cap+3.53000e-05'
+ mcm5m1f_ca_w_0_140_s_3_500 = '-3.68750e-07*ic_cap*ic_cap+-2.25000e-07*ic_cap+3.53000e-05'
+ mcm5m1f_ca_w_1_120_s_0_140 = '-3.68750e-07*ic_cap*ic_cap+-2.25000e-07*ic_cap+3.53000e-05'
+ mcm5m1f_ca_w_1_120_s_0_175 = '-3.68750e-07*ic_cap*ic_cap+-2.25000e-07*ic_cap+3.53000e-05'
+ mcm5m1f_ca_w_1_120_s_0_210 = '-3.68750e-07*ic_cap*ic_cap+-2.25000e-07*ic_cap+3.53000e-05'
+ mcm5m1f_ca_w_1_120_s_0_280 = '-3.68750e-07*ic_cap*ic_cap+-2.25000e-07*ic_cap+3.53000e-05'
+ mcm5m1f_ca_w_1_120_s_0_350 = '-3.68750e-07*ic_cap*ic_cap+-2.25000e-07*ic_cap+3.53000e-05'
+ mcm5m1f_ca_w_1_120_s_0_420 = '-3.68750e-07*ic_cap*ic_cap+-2.25000e-07*ic_cap+3.53000e-05'
+ mcm5m1f_ca_w_1_120_s_0_560 = '-3.68750e-07*ic_cap*ic_cap+-2.25000e-07*ic_cap+3.53000e-05'
+ mcm5m1f_ca_w_1_120_s_0_840 = '-3.68750e-07*ic_cap*ic_cap+-2.25000e-07*ic_cap+3.53000e-05'
+ mcm5m1f_ca_w_1_120_s_1_540 = '-3.68750e-07*ic_cap*ic_cap+-2.25000e-07*ic_cap+3.53000e-05'
+ mcm5m1f_ca_w_1_120_s_3_500 = '-3.68750e-07*ic_cap*ic_cap+-2.25000e-07*ic_cap+3.53000e-05'
+ mcm5m1f_cc_w_0_140_s_0_140 = '-9.28125e-13*ic_cap*ic_cap+-5.37500e-13*ic_cap+1.04000e-10'
+ mcm5m1f_cc_w_0_140_s_0_175 = '-8.43750e-13*ic_cap*ic_cap+-6.00000e-13*ic_cap+1.02000e-10'
+ mcm5m1f_cc_w_0_140_s_0_210 = '-7.81250e-13*ic_cap*ic_cap+-4.25000e-13*ic_cap+9.71000e-11'
+ mcm5m1f_cc_w_0_140_s_0_280 = '-5.75000e-13*ic_cap*ic_cap+-4.00000e-13*ic_cap+8.58000e-11'
+ mcm5m1f_cc_w_0_140_s_0_350 = '-4.53125e-13*ic_cap*ic_cap+-2.62500e-13*ic_cap+7.46000e-11'
+ mcm5m1f_cc_w_0_140_s_0_420 = '-3.53125e-13*ic_cap*ic_cap+-2.37500e-13*ic_cap+6.50000e-11'
+ mcm5m1f_cc_w_0_140_s_0_560 = '-1.90625e-13*ic_cap*ic_cap+-1.37500e-13*ic_cap+5.17000e-11'
+ mcm5m1f_cc_w_0_140_s_0_840 = '-7.18750e-14*ic_cap*ic_cap+-6.25000e-14*ic_cap+3.70000e-11'
+ mcm5m1f_cc_w_0_140_s_1_540 = '3.43750e-14*ic_cap*ic_cap+1.25000e-14*ic_cap+1.97000e-11'
+ mcm5m1f_cc_w_0_140_s_3_500 = '5.75000e-14*ic_cap*ic_cap+3.75000e-14*ic_cap+4.95000e-12'
+ mcm5m1f_cc_w_1_120_s_0_140 = '-7.50000e-13*ic_cap*ic_cap+-5.00000e-13*ic_cap+1.25000e-10'
+ mcm5m1f_cc_w_1_120_s_0_175 = '-8.12500e-13*ic_cap*ic_cap+-2.50000e-13*ic_cap+1.23000e-10'
+ mcm5m1f_cc_w_1_120_s_0_210 = '-6.56250e-13*ic_cap*ic_cap+-3.75000e-13*ic_cap+1.16000e-10'
+ mcm5m1f_cc_w_1_120_s_0_280 = '-4.93750e-13*ic_cap*ic_cap+-3.25000e-13*ic_cap+1.02000e-10'
+ mcm5m1f_cc_w_1_120_s_0_350 = '-3.68750e-13*ic_cap*ic_cap+-2.25000e-13*ic_cap+8.91000e-11'
+ mcm5m1f_cc_w_1_120_s_0_420 = '-2.65625e-13*ic_cap*ic_cap+-1.37500e-13*ic_cap+7.82000e-11'
+ mcm5m1f_cc_w_1_120_s_0_560 = '-1.09375e-13*ic_cap*ic_cap+-8.75000e-14*ic_cap+6.26000e-11'
+ mcm5m1f_cc_w_1_120_s_0_840 = '6.25000e-15*ic_cap*ic_cap+4.47000e-11'
+ mcm5m1f_cc_w_1_120_s_1_540 = '9.06250e-14*ic_cap*ic_cap+6.25000e-14*ic_cap+2.43000e-11'
+ mcm5m1f_cc_w_1_120_s_3_500 = '8.59375e-14*ic_cap*ic_cap+5.37500e-14*ic_cap+6.46000e-12'
+ mcm5m1f_cf_w_0_140_s_0_140 = '-1.87500e-15*ic_cap*ic_cap+-2.50000e-15*ic_cap+2.45000e-12'
+ mcm5m1f_cf_w_0_140_s_0_175 = '-8.43750e-15*ic_cap*ic_cap+-6.25000e-15*ic_cap+3.06000e-12'
+ mcm5m1f_cf_w_0_140_s_0_210 = '-1.40625e-14*ic_cap*ic_cap+-8.75000e-15*ic_cap+3.68000e-12'
+ mcm5m1f_cf_w_0_140_s_0_280 = '-2.75000e-14*ic_cap*ic_cap+-1.75000e-14*ic_cap+4.88000e-12'
+ mcm5m1f_cf_w_0_140_s_0_350 = '-3.96875e-14*ic_cap*ic_cap+-2.37500e-14*ic_cap+6.06000e-12'
+ mcm5m1f_cf_w_0_140_s_0_420 = '-5.25000e-14*ic_cap*ic_cap+-3.50000e-14*ic_cap+7.28000e-12'
+ mcm5m1f_cf_w_0_140_s_0_560 = '-7.59375e-14*ic_cap*ic_cap+-4.62500e-14*ic_cap+9.53000e-12'
+ mcm5m1f_cf_w_0_140_s_0_840 = '-1.18750e-13*ic_cap*ic_cap+-7.50000e-14*ic_cap+1.37000e-11'
+ mcm5m1f_cf_w_0_140_s_1_540 = '-1.87500e-13*ic_cap*ic_cap+-1.25000e-13*ic_cap+2.20000e-11'
+ mcm5m1f_cf_w_0_140_s_3_500 = '-2.28125e-13*ic_cap*ic_cap+-1.62500e-13*ic_cap+3.32000e-11'
+ mcm5m1f_cf_w_1_120_s_0_140 = '-2.50000e-15*ic_cap*ic_cap+-2.50000e-15*ic_cap+2.49000e-12'
+ mcm5m1f_cf_w_1_120_s_0_175 = '-8.75000e-15*ic_cap*ic_cap+-7.50000e-15*ic_cap+3.10000e-12'
+ mcm5m1f_cf_w_1_120_s_0_210 = '-1.62500e-14*ic_cap*ic_cap+-1.00000e-14*ic_cap+3.72000e-12'
+ mcm5m1f_cf_w_1_120_s_0_280 = '-2.71875e-14*ic_cap*ic_cap+-1.62500e-14*ic_cap+4.92000e-12'
+ mcm5m1f_cf_w_1_120_s_0_350 = '-3.96875e-14*ic_cap*ic_cap+-2.62500e-14*ic_cap+6.11000e-12'
+ mcm5m1f_cf_w_1_120_s_0_420 = '-5.25000e-14*ic_cap*ic_cap+-3.50000e-14*ic_cap+7.29000e-12'
+ mcm5m1f_cf_w_1_120_s_0_560 = '-7.59375e-14*ic_cap*ic_cap+-4.62500e-14*ic_cap+9.56000e-12'
+ mcm5m1f_cf_w_1_120_s_0_840 = '-1.15625e-13*ic_cap*ic_cap+-6.25000e-14*ic_cap+1.38000e-11'
+ mcm5m1f_cf_w_1_120_s_1_540 = '-1.90625e-13*ic_cap*ic_cap+-1.12500e-13*ic_cap+2.26000e-11'
+ mcm5m1f_cf_w_1_120_s_3_500 = '-2.31250e-13*ic_cap*ic_cap+-1.50000e-13*ic_cap+3.55000e-11'
+ mcm5m1l1_ca_w_0_140_s_0_140 = '-2.01875e-06*ic_cap*ic_cap+-1.30000e-06*ic_cap+1.23000e-04'
+ mcm5m1l1_ca_w_0_140_s_0_175 = '-2.01875e-06*ic_cap*ic_cap+-1.30000e-06*ic_cap+1.23000e-04'
+ mcm5m1l1_ca_w_0_140_s_0_210 = '-2.01875e-06*ic_cap*ic_cap+-1.30000e-06*ic_cap+1.23000e-04'
+ mcm5m1l1_ca_w_0_140_s_0_280 = '-2.01875e-06*ic_cap*ic_cap+-1.30000e-06*ic_cap+1.23000e-04'
+ mcm5m1l1_ca_w_0_140_s_0_350 = '-2.01875e-06*ic_cap*ic_cap+-1.30000e-06*ic_cap+1.23000e-04'
+ mcm5m1l1_ca_w_0_140_s_0_420 = '-2.01875e-06*ic_cap*ic_cap+-1.30000e-06*ic_cap+1.23000e-04'
+ mcm5m1l1_ca_w_0_140_s_0_560 = '-2.01875e-06*ic_cap*ic_cap+-1.30000e-06*ic_cap+1.23000e-04'
+ mcm5m1l1_ca_w_0_140_s_0_840 = '-2.01875e-06*ic_cap*ic_cap+-1.30000e-06*ic_cap+1.23000e-04'
+ mcm5m1l1_ca_w_0_140_s_1_540 = '-2.01875e-06*ic_cap*ic_cap+-1.30000e-06*ic_cap+1.23000e-04'
+ mcm5m1l1_ca_w_0_140_s_3_500 = '-2.01875e-06*ic_cap*ic_cap+-1.30000e-06*ic_cap+1.23000e-04'
+ mcm5m1l1_ca_w_1_120_s_0_140 = '-2.01875e-06*ic_cap*ic_cap+-1.30000e-06*ic_cap+1.23000e-04'
+ mcm5m1l1_ca_w_1_120_s_0_175 = '-2.01875e-06*ic_cap*ic_cap+-1.30000e-06*ic_cap+1.23000e-04'
+ mcm5m1l1_ca_w_1_120_s_0_210 = '-2.01875e-06*ic_cap*ic_cap+-1.30000e-06*ic_cap+1.23000e-04'
+ mcm5m1l1_ca_w_1_120_s_0_280 = '-2.01875e-06*ic_cap*ic_cap+-1.30000e-06*ic_cap+1.23000e-04'
+ mcm5m1l1_ca_w_1_120_s_0_350 = '-2.01875e-06*ic_cap*ic_cap+-1.30000e-06*ic_cap+1.23000e-04'
+ mcm5m1l1_ca_w_1_120_s_0_420 = '-2.01875e-06*ic_cap*ic_cap+-1.30000e-06*ic_cap+1.23000e-04'
+ mcm5m1l1_ca_w_1_120_s_0_560 = '-2.01875e-06*ic_cap*ic_cap+-1.30000e-06*ic_cap+1.23000e-04'
+ mcm5m1l1_ca_w_1_120_s_0_840 = '-2.01875e-06*ic_cap*ic_cap+-1.30000e-06*ic_cap+1.23000e-04'
+ mcm5m1l1_ca_w_1_120_s_1_540 = '-2.01875e-06*ic_cap*ic_cap+-1.30000e-06*ic_cap+1.23000e-04'
+ mcm5m1l1_ca_w_1_120_s_3_500 = '-2.01875e-06*ic_cap*ic_cap+-1.30000e-06*ic_cap+1.23000e-04'
+ mcm5m1l1_cc_w_0_140_s_0_140 = '-8.03125e-13*ic_cap*ic_cap+-3.87500e-13*ic_cap+9.56000e-11'
+ mcm5m1l1_cc_w_0_140_s_0_175 = '-7.46875e-13*ic_cap*ic_cap+-4.62500e-13*ic_cap+9.31000e-11'
+ mcm5m1l1_cc_w_0_140_s_0_210 = '-6.09375e-13*ic_cap*ic_cap+-3.37500e-13*ic_cap+8.67000e-11'
+ mcm5m1l1_cc_w_0_140_s_0_280 = '-4.18750e-13*ic_cap*ic_cap+-2.75000e-13*ic_cap+7.45000e-11'
+ mcm5m1l1_cc_w_0_140_s_0_350 = '-2.93750e-13*ic_cap*ic_cap+-2.25000e-13*ic_cap+6.24000e-11'
+ mcm5m1l1_cc_w_0_140_s_0_420 = '-1.84375e-13*ic_cap*ic_cap+-1.12500e-13*ic_cap+5.25000e-11'
+ mcm5m1l1_cc_w_0_140_s_0_560 = '-5.62500e-14*ic_cap*ic_cap+-2.50000e-14*ic_cap+3.86000e-11'
+ mcm5m1l1_cc_w_0_140_s_0_840 = '3.12500e-14*ic_cap*ic_cap+5.00000e-14*ic_cap+2.38000e-11'
+ mcm5m1l1_cc_w_0_140_s_1_540 = '6.34375e-14*ic_cap*ic_cap+4.87500e-14*ic_cap+9.09000e-12'
+ mcm5m1l1_cc_w_0_140_s_3_500 = '2.21875e-14*ic_cap*ic_cap+1.62500e-14*ic_cap+1.36000e-12'
+ mcm5m1l1_cc_w_1_120_s_0_140 = '-6.56250e-13*ic_cap*ic_cap+-2.50000e-13*ic_cap+1.09000e-10'
+ mcm5m1l1_cc_w_1_120_s_0_175 = '-6.65625e-13*ic_cap*ic_cap+-2.37500e-13*ic_cap+1.06000e-10'
+ mcm5m1l1_cc_w_1_120_s_0_210 = '-5.09375e-13*ic_cap*ic_cap+-2.62500e-13*ic_cap+9.89000e-11'
+ mcm5m1l1_cc_w_1_120_s_0_280 = '-3.46875e-13*ic_cap*ic_cap+-1.62500e-13*ic_cap+8.49000e-11'
+ mcm5m1l1_cc_w_1_120_s_0_350 = '-2.46875e-13*ic_cap*ic_cap+-1.37500e-13*ic_cap+7.23000e-11'
+ mcm5m1l1_cc_w_1_120_s_0_420 = '-1.28125e-13*ic_cap*ic_cap+-6.25000e-14*ic_cap+6.11000e-11'
+ mcm5m1l1_cc_w_1_120_s_0_560 = '-1.56250e-14*ic_cap*ic_cap+1.25000e-14*ic_cap+4.62000e-11'
+ mcm5m1l1_cc_w_1_120_s_0_840 = '7.18750e-14*ic_cap*ic_cap+6.25000e-14*ic_cap+2.95000e-11'
+ mcm5m1l1_cc_w_1_120_s_1_540 = '9.37500e-14*ic_cap*ic_cap+7.50000e-14*ic_cap+1.26000e-11'
+ mcm5m1l1_cc_w_1_120_s_3_500 = '3.65625e-14*ic_cap*ic_cap+3.12500e-14*ic_cap+2.20000e-12'
+ mcm5m1l1_cf_w_0_140_s_0_140 = '-6.09375e-14*ic_cap*ic_cap+-4.87500e-14*ic_cap+8.10000e-12'
+ mcm5m1l1_cf_w_0_140_s_0_175 = '-9.34375e-14*ic_cap*ic_cap+-6.87500e-14*ic_cap+1.02000e-11'
+ mcm5m1l1_cf_w_0_140_s_0_210 = '-1.29062e-13*ic_cap*ic_cap+-9.12500e-14*ic_cap+1.23000e-11'
+ mcm5m1l1_cf_w_0_140_s_0_280 = '-1.90625e-13*ic_cap*ic_cap+-1.37500e-13*ic_cap+1.62000e-11'
+ mcm5m1l1_cf_w_0_140_s_0_350 = '-2.40625e-13*ic_cap*ic_cap+-1.62500e-13*ic_cap+1.97000e-11'
+ mcm5m1l1_cf_w_0_140_s_0_420 = '-2.87500e-13*ic_cap*ic_cap+-2.00000e-13*ic_cap+2.31000e-11'
+ mcm5m1l1_cf_w_0_140_s_0_560 = '-3.62500e-13*ic_cap*ic_cap+-2.50000e-13*ic_cap+2.90000e-11'
+ mcm5m1l1_cf_w_0_140_s_0_840 = '-4.59375e-13*ic_cap*ic_cap+-3.12500e-13*ic_cap+3.80000e-11'
+ mcm5m1l1_cf_w_0_140_s_1_540 = '-5.15625e-13*ic_cap*ic_cap+-3.62500e-13*ic_cap+4.98000e-11'
+ mcm5m1l1_cf_w_0_140_s_3_500 = '-4.93750e-13*ic_cap*ic_cap+-3.25000e-13*ic_cap+5.74000e-11'
+ mcm5m1l1_cf_w_1_120_s_0_140 = '-6.37500e-14*ic_cap*ic_cap+-5.25000e-14*ic_cap+8.26000e-12'
+ mcm5m1l1_cf_w_1_120_s_0_175 = '-9.96875e-14*ic_cap*ic_cap+-7.37500e-14*ic_cap+1.04000e-11'
+ mcm5m1l1_cf_w_1_120_s_0_210 = '-1.30313e-13*ic_cap*ic_cap+-9.62500e-14*ic_cap+1.24000e-11'
+ mcm5m1l1_cf_w_1_120_s_0_280 = '-1.90625e-13*ic_cap*ic_cap+-1.37500e-13*ic_cap+1.63000e-11'
+ mcm5m1l1_cf_w_1_120_s_0_350 = '-2.43750e-13*ic_cap*ic_cap+-1.75000e-13*ic_cap+1.99000e-11'
+ mcm5m1l1_cf_w_1_120_s_0_420 = '-2.93750e-13*ic_cap*ic_cap+-2.00000e-13*ic_cap+2.33000e-11'
+ mcm5m1l1_cf_w_1_120_s_0_560 = '-3.62500e-13*ic_cap*ic_cap+-2.50000e-13*ic_cap+2.91000e-11'
+ mcm5m1l1_cf_w_1_120_s_0_840 = '-4.59375e-13*ic_cap*ic_cap+-3.12500e-13*ic_cap+3.83000e-11'
+ mcm5m1l1_cf_w_1_120_s_1_540 = '-5.09375e-13*ic_cap*ic_cap+-3.62500e-13*ic_cap+5.10000e-11'
+ mcm5m1l1_cf_w_1_120_s_3_500 = '-4.87500e-13*ic_cap*ic_cap+-3.50000e-13*ic_cap+6.09000e-11'
+ mcm5m1p1_ca_w_0_140_s_0_140 = '-7.50000e-07*ic_cap*ic_cap+-4.50000e-07*ic_cap+5.44000e-05'
+ mcm5m1p1_ca_w_0_140_s_0_175 = '-7.50000e-07*ic_cap*ic_cap+-4.50000e-07*ic_cap+5.44000e-05'
+ mcm5m1p1_ca_w_0_140_s_0_210 = '-7.50000e-07*ic_cap*ic_cap+-4.50000e-07*ic_cap+5.44000e-05'
+ mcm5m1p1_ca_w_0_140_s_0_280 = '-7.50000e-07*ic_cap*ic_cap+-4.50000e-07*ic_cap+5.44000e-05'
+ mcm5m1p1_ca_w_0_140_s_0_350 = '-7.50000e-07*ic_cap*ic_cap+-4.50000e-07*ic_cap+5.44000e-05'
+ mcm5m1p1_ca_w_0_140_s_0_420 = '-7.50000e-07*ic_cap*ic_cap+-4.50000e-07*ic_cap+5.44000e-05'
+ mcm5m1p1_ca_w_0_140_s_0_560 = '-7.50000e-07*ic_cap*ic_cap+-4.50000e-07*ic_cap+5.44000e-05'
+ mcm5m1p1_ca_w_0_140_s_0_840 = '-7.50000e-07*ic_cap*ic_cap+-4.50000e-07*ic_cap+5.44000e-05'
+ mcm5m1p1_ca_w_0_140_s_1_540 = '-7.50000e-07*ic_cap*ic_cap+-4.50000e-07*ic_cap+5.44000e-05'
+ mcm5m1p1_ca_w_0_140_s_3_500 = '-7.50000e-07*ic_cap*ic_cap+-4.50000e-07*ic_cap+5.44000e-05'
+ mcm5m1p1_ca_w_1_120_s_0_140 = '-7.50000e-07*ic_cap*ic_cap+-4.50000e-07*ic_cap+5.44000e-05'
+ mcm5m1p1_ca_w_1_120_s_0_175 = '-7.50000e-07*ic_cap*ic_cap+-4.50000e-07*ic_cap+5.44000e-05'
+ mcm5m1p1_ca_w_1_120_s_0_210 = '-7.50000e-07*ic_cap*ic_cap+-4.50000e-07*ic_cap+5.44000e-05'
+ mcm5m1p1_ca_w_1_120_s_0_280 = '-7.50000e-07*ic_cap*ic_cap+-4.50000e-07*ic_cap+5.44000e-05'
+ mcm5m1p1_ca_w_1_120_s_0_350 = '-7.50000e-07*ic_cap*ic_cap+-4.50000e-07*ic_cap+5.44000e-05'
+ mcm5m1p1_ca_w_1_120_s_0_420 = '-7.50000e-07*ic_cap*ic_cap+-4.50000e-07*ic_cap+5.44000e-05'
+ mcm5m1p1_ca_w_1_120_s_0_560 = '-7.50000e-07*ic_cap*ic_cap+-4.50000e-07*ic_cap+5.44000e-05'
+ mcm5m1p1_ca_w_1_120_s_0_840 = '-7.50000e-07*ic_cap*ic_cap+-4.50000e-07*ic_cap+5.44000e-05'
+ mcm5m1p1_ca_w_1_120_s_1_540 = '-7.50000e-07*ic_cap*ic_cap+-4.50000e-07*ic_cap+5.44000e-05'
+ mcm5m1p1_ca_w_1_120_s_3_500 = '-7.50000e-07*ic_cap*ic_cap+-4.50000e-07*ic_cap+5.44000e-05'
+ mcm5m1p1_cc_w_0_140_s_0_140 = '-8.93750e-13*ic_cap*ic_cap+-5.00000e-13*ic_cap+1.02000e-10'
+ mcm5m1p1_cc_w_0_140_s_0_175 = '-8.12500e-13*ic_cap*ic_cap+-5.75000e-13*ic_cap+9.98000e-11'
+ mcm5m1p1_cc_w_0_140_s_0_210 = '-7.15625e-13*ic_cap*ic_cap+-4.37500e-13*ic_cap+9.41000e-11'
+ mcm5m1p1_cc_w_0_140_s_0_280 = '-5.31250e-13*ic_cap*ic_cap+-3.00000e-13*ic_cap+8.27000e-11'
+ mcm5m1p1_cc_w_0_140_s_0_350 = '-3.71875e-13*ic_cap*ic_cap+-2.37500e-13*ic_cap+7.09000e-11'
+ mcm5m1p1_cc_w_0_140_s_0_420 = '-2.65625e-13*ic_cap*ic_cap+-2.12500e-13*ic_cap+6.10000e-11'
+ mcm5m1p1_cc_w_0_140_s_0_560 = '-1.31250e-13*ic_cap*ic_cap+-1.00000e-13*ic_cap+4.76000e-11'
+ mcm5m1p1_cc_w_0_140_s_1_540 = '8.12500e-14*ic_cap*ic_cap+5.00000e-14*ic_cap+1.52000e-11'
+ mcm5m1p1_cc_w_0_140_s_3_500 = '5.25000e-14*ic_cap*ic_cap+4.00000e-14*ic_cap+2.95000e-12'
+ mcm5m1p1_cc_w_1_120_s_0_140 = '-7.18750e-13*ic_cap*ic_cap+-3.75000e-13*ic_cap+1.20000e-10'
+ mcm5m1p1_cc_w_1_120_s_0_175 = '-6.87500e-13*ic_cap*ic_cap+-2.50000e-13*ic_cap+1.16000e-10'
+ mcm5m1p1_cc_w_1_120_s_0_210 = '-5.81250e-13*ic_cap*ic_cap+-3.25000e-13*ic_cap+1.10000e-10'
+ mcm5m1p1_cc_w_1_120_s_0_280 = '-3.84375e-13*ic_cap*ic_cap+-2.87500e-13*ic_cap+9.54000e-11'
+ mcm5m1p1_cc_w_1_120_s_0_350 = '-2.62500e-13*ic_cap*ic_cap+-1.50000e-13*ic_cap+8.27000e-11'
+ mcm5m1p1_cc_w_1_120_s_0_420 = '-1.68750e-13*ic_cap*ic_cap+-1.25000e-13*ic_cap+7.19000e-11'
+ mcm5m1p1_cc_w_1_120_s_0_560 = '-2.81250e-14*ic_cap*ic_cap+-3.75000e-14*ic_cap+5.62000e-11'
+ mcm5m1p1_cc_w_1_120_s_0_840 = '6.56250e-14*ic_cap*ic_cap+3.75000e-14*ic_cap+3.86000e-11'
+ mcm5m1p1_cc_w_1_120_s_1_540 = '1.21875e-13*ic_cap*ic_cap+8.75000e-14*ic_cap+1.91000e-11'
+ mcm5m1p1_cc_w_1_120_s_3_500 = '7.78125e-14*ic_cap*ic_cap+5.37500e-14*ic_cap+4.05000e-12'
+ mcm5m1p1_cf_w_0_140_s_0_140 = '-1.87500e-14*ic_cap*ic_cap+-1.25000e-14*ic_cap+3.77000e-12'
+ mcm5m1p1_cf_w_0_140_s_0_175 = '-3.18750e-14*ic_cap*ic_cap+-2.00000e-14*ic_cap+4.71000e-12'
+ mcm5m1p1_cf_w_0_140_s_0_210 = '-4.37500e-14*ic_cap*ic_cap+-2.75000e-14*ic_cap+5.65000e-12'
+ mcm5m1p1_cf_w_0_140_s_0_280 = '-6.90625e-14*ic_cap*ic_cap+-4.37500e-14*ic_cap+7.48000e-12'
+ mcm5m1p1_cf_w_0_140_s_0_350 = '-9.18750e-14*ic_cap*ic_cap+-5.75000e-14*ic_cap+9.24000e-12'
+ mcm5m1p1_cf_w_0_140_s_0_420 = '-1.13750e-13*ic_cap*ic_cap+-7.25000e-14*ic_cap+1.10000e-11'
+ mcm5m1p1_cf_w_0_140_s_0_560 = '-1.56250e-13*ic_cap*ic_cap+-1.00000e-13*ic_cap+1.43000e-11'
+ mcm5m1p1_cf_w_0_140_s_0_840 = '-2.31250e-13*ic_cap*ic_cap+-1.50000e-13*ic_cap+2.01000e-11'
+ mcm5m1p1_cf_w_0_140_s_1_540 = '-3.12500e-13*ic_cap*ic_cap+-2.00000e-13*ic_cap+3.03000e-11'
+ mcm5m1p1_cf_w_0_140_s_3_500 = '-3.18750e-13*ic_cap*ic_cap+-2.00000e-13*ic_cap+4.08000e-11'
+ mcm5m1p1_cf_w_1_120_s_0_140 = '-2.15625e-14*ic_cap*ic_cap+-1.62500e-14*ic_cap+3.92000e-12'
+ mcm5m1p1_cf_w_1_120_s_0_175 = '-3.43750e-14*ic_cap*ic_cap+-2.25000e-14*ic_cap+4.86000e-12'
+ mcm5m1p1_cf_w_1_120_s_0_210 = '-4.68750e-14*ic_cap*ic_cap+-3.00000e-14*ic_cap+5.78000e-12'
+ mcm5m1p1_cf_w_1_120_s_0_280 = '-7.06250e-14*ic_cap*ic_cap+-4.25000e-14*ic_cap+7.61000e-12'
+ mcm5m1p1_cf_w_1_120_s_0_350 = '-9.50000e-14*ic_cap*ic_cap+-6.00000e-14*ic_cap+9.40000e-12'
+ mcm5m1p1_cf_w_1_120_s_0_420 = '-1.21875e-13*ic_cap*ic_cap+-7.25000e-14*ic_cap+1.12000e-11'
+ mcm5m1p1_cf_w_1_120_s_0_560 = '-1.56250e-13*ic_cap*ic_cap+-1.00000e-13*ic_cap+1.44000e-11'
+ mcm5m1p1_cf_w_1_120_s_0_840 = '-2.28125e-13*ic_cap*ic_cap+-1.37500e-13*ic_cap+2.04000e-11'
+ mcm5m1p1_cf_w_1_120_s_1_540 = '-3.25000e-13*ic_cap*ic_cap+-2.00000e-13*ic_cap+3.13000e-11'
+ mcm5m1p1_cf_w_1_120_s_3_500 = '-3.25000e-13*ic_cap*ic_cap+-2.00000e-13*ic_cap+4.36000e-11'
+ mcm5m2_ca_w_1_600_s_10_000 = '-7.50000e-08*ic_cap*ic_cap+-5.00000e-08*ic_cap+1.15000e-05'
+ mcm5m2_ca_w_1_600_s_12_000 = '-7.50000e-08*ic_cap*ic_cap+-5.00000e-08*ic_cap+1.15000e-05'
+ mcm5m2_ca_w_1_600_s_1_600 = '-7.50000e-08*ic_cap*ic_cap+-5.00000e-08*ic_cap+1.15000e-05'
+ mcm5m2_ca_w_1_600_s_1_700 = '-7.50000e-08*ic_cap*ic_cap+-5.00000e-08*ic_cap+1.15000e-05'
+ mcm5m2_ca_w_1_600_s_1_900 = '-7.50000e-08*ic_cap*ic_cap+-5.00000e-08*ic_cap+1.15000e-05'
+ mcm5m2_ca_w_1_600_s_2_000 = '-7.50000e-08*ic_cap*ic_cap+-5.00000e-08*ic_cap+1.15000e-05'
+ mcm5m2_ca_w_1_600_s_2_400 = '-7.50000e-08*ic_cap*ic_cap+-5.00000e-08*ic_cap+1.15000e-05'
+ mcm5m2_ca_w_1_600_s_2_800 = '-7.50000e-08*ic_cap*ic_cap+-5.00000e-08*ic_cap+1.15000e-05'
+ mcm5m2_ca_w_1_600_s_3_200 = '-7.50000e-08*ic_cap*ic_cap+-5.00000e-08*ic_cap+1.15000e-05'
+ mcm5m2_ca_w_1_600_s_4_800 = '-7.50000e-08*ic_cap*ic_cap+-5.00000e-08*ic_cap+1.15000e-05'
+ mcm5m2_ca_w_4_000_s_10_000 = '-7.50000e-08*ic_cap*ic_cap+-5.00000e-08*ic_cap+1.15000e-05'
+ mcm5m2_ca_w_4_000_s_12_000 = '-7.50000e-08*ic_cap*ic_cap+-5.00000e-08*ic_cap+1.15000e-05'
+ mcm5m2_ca_w_4_000_s_1_600 = '-7.50000e-08*ic_cap*ic_cap+-5.00000e-08*ic_cap+1.15000e-05'
+ mcm5m2_ca_w_4_000_s_1_700 = '-7.50000e-08*ic_cap*ic_cap+-5.00000e-08*ic_cap+1.15000e-05'
+ mcm5m2_ca_w_4_000_s_1_900 = '-7.50000e-08*ic_cap*ic_cap+-5.00000e-08*ic_cap+1.15000e-05'
+ mcm5m2_ca_w_4_000_s_2_000 = '-7.50000e-08*ic_cap*ic_cap+-5.00000e-08*ic_cap+1.15000e-05'
+ mcm5m2_ca_w_4_000_s_2_400 = '-7.50000e-08*ic_cap*ic_cap+-5.00000e-08*ic_cap+1.15000e-05'
+ mcm5m2_ca_w_4_000_s_2_800 = '-7.50000e-08*ic_cap*ic_cap+-5.00000e-08*ic_cap+1.15000e-05'
+ mcm5m2_ca_w_4_000_s_3_200 = '-7.50000e-08*ic_cap*ic_cap+-5.00000e-08*ic_cap+1.15000e-05'
+ mcm5m2_ca_w_4_000_s_4_800 = '-7.50000e-08*ic_cap*ic_cap+-5.00000e-08*ic_cap+1.15000e-05'
+ mcm5m2_cc_w_1_600_s_10_000 = '-1.87500e-15*ic_cap*ic_cap+-2.50000e-15*ic_cap+9.75000e-12'
+ mcm5m2_cc_w_1_600_s_12_000 = '1.87500e-15*ic_cap*ic_cap+-2.50000e-15*ic_cap+7.42000e-12'
+ mcm5m2_cc_w_1_600_s_1_600 = '-4.53125e-13*ic_cap*ic_cap+-2.87500e-13*ic_cap+6.87000e-11'
+ mcm5m2_cc_w_1_600_s_1_700 = '-4.12500e-13*ic_cap*ic_cap+-2.75000e-13*ic_cap+6.51000e-11'
+ mcm5m2_cc_w_1_600_s_1_900 = '-3.37500e-13*ic_cap*ic_cap+-2.25000e-13*ic_cap+5.88000e-11'
+ mcm5m2_cc_w_1_600_s_2_000 = '-3.03125e-13*ic_cap*ic_cap+-2.12500e-13*ic_cap+5.61000e-11'
+ mcm5m2_cc_w_1_600_s_2_400 = '-2.25000e-13*ic_cap*ic_cap+-1.50000e-13*ic_cap+4.77000e-11'
+ mcm5m2_cc_w_1_600_s_2_800 = '-1.71875e-13*ic_cap*ic_cap+-1.12500e-13*ic_cap+4.14000e-11'
+ mcm5m2_cc_w_1_600_s_3_200 = '-1.31250e-13*ic_cap*ic_cap+-1.00000e-13*ic_cap+3.65000e-11'
+ mcm5m2_cc_w_1_600_s_4_800 = '-5.31250e-14*ic_cap*ic_cap+-3.75000e-14*ic_cap+2.43000e-11'
+ mcm5m2_cc_w_4_000_s_10_000 = '6.25000e-15*ic_cap*ic_cap+1.21000e-11'
+ mcm5m2_cc_w_4_000_s_12_000 = '1.56250e-15*ic_cap*ic_cap+6.25000e-15*ic_cap+9.55000e-12'
+ mcm5m2_cc_w_4_000_s_1_600 = '-4.31250e-13*ic_cap*ic_cap+-3.00000e-13*ic_cap+7.45000e-11'
+ mcm5m2_cc_w_4_000_s_1_700 = '-3.84375e-13*ic_cap*ic_cap+-2.62500e-13*ic_cap+7.06000e-11'
+ mcm5m2_cc_w_4_000_s_1_900 = '-3.12500e-13*ic_cap*ic_cap+-2.00000e-13*ic_cap+6.41000e-11'
+ mcm5m2_cc_w_4_000_s_2_000 = '-2.84375e-13*ic_cap*ic_cap+-1.87500e-13*ic_cap+6.13000e-11'
+ mcm5m2_cc_w_4_000_s_2_400 = '-2.09375e-13*ic_cap*ic_cap+-1.37500e-13*ic_cap+5.25000e-11'
+ mcm5m2_cc_w_4_000_s_2_800 = '-1.53125e-13*ic_cap*ic_cap+-1.12500e-13*ic_cap+4.59000e-11'
+ mcm5m2_cc_w_4_000_s_3_200 = '-1.12500e-13*ic_cap*ic_cap+-7.50000e-14*ic_cap+4.07000e-11'
+ mcm5m2_cc_w_4_000_s_4_800 = '-4.37500e-14*ic_cap*ic_cap+-2.50000e-14*ic_cap+2.79000e-11'
+ mcm5m2_cf_w_1_600_s_10_000 = '-1.53125e-13*ic_cap*ic_cap+-8.75000e-14*ic_cap+3.23000e-11'
+ mcm5m2_cf_w_1_600_s_12_000 = '-1.56250e-13*ic_cap*ic_cap+-1.00000e-13*ic_cap+3.44000e-11'
+ mcm5m2_cf_w_1_600_s_1_600 = '-2.84375e-14*ic_cap*ic_cap+-1.62500e-14*ic_cap+8.63000e-12'
+ mcm5m2_cf_w_1_600_s_1_700 = '-3.18750e-14*ic_cap*ic_cap+-2.00000e-14*ic_cap+9.13000e-12'
+ mcm5m2_cf_w_1_600_s_1_900 = '-3.78125e-14*ic_cap*ic_cap+-2.37500e-14*ic_cap+1.01000e-11'
+ mcm5m2_cf_w_1_600_s_2_000 = '-4.31250e-14*ic_cap*ic_cap+-2.25000e-14*ic_cap+1.06000e-11'
+ mcm5m2_cf_w_1_600_s_2_400 = '-5.00000e-14*ic_cap*ic_cap+-2.50000e-14*ic_cap+1.24000e-11'
+ mcm5m2_cf_w_1_600_s_2_800 = '-6.56250e-14*ic_cap*ic_cap+-3.75000e-14*ic_cap+1.42000e-11'
+ mcm5m2_cf_w_1_600_s_3_200 = '-7.50000e-14*ic_cap*ic_cap+-5.00000e-14*ic_cap+1.59000e-11'
+ mcm5m2_cf_w_1_600_s_4_800 = '-1.06250e-13*ic_cap*ic_cap+-7.50000e-14*ic_cap+2.16000e-11'
+ mcm5m2_cf_w_4_000_s_10_000 = '-1.46875e-13*ic_cap*ic_cap+-8.75000e-14*ic_cap+3.29000e-11'
+ mcm5m2_cf_w_4_000_s_12_000 = '-1.50000e-13*ic_cap*ic_cap+-1.00000e-13*ic_cap+3.52000e-11'
+ mcm5m2_cf_w_4_000_s_1_600 = '-2.81250e-14*ic_cap*ic_cap+-1.75000e-14*ic_cap+8.63000e-12'
+ mcm5m2_cf_w_4_000_s_1_700 = '-3.12500e-14*ic_cap*ic_cap+-2.00000e-14*ic_cap+9.13000e-12'
+ mcm5m2_cf_w_4_000_s_1_900 = '-3.71875e-14*ic_cap*ic_cap+-2.37500e-14*ic_cap+1.01000e-11'
+ mcm5m2_cf_w_4_000_s_2_000 = '-4.25000e-14*ic_cap*ic_cap+-2.00000e-14*ic_cap+1.06000e-11'
+ mcm5m2_cf_w_4_000_s_2_400 = '-5.62500e-14*ic_cap*ic_cap+-2.50000e-14*ic_cap+1.25000e-11'
+ mcm5m2_cf_w_4_000_s_2_800 = '-6.25000e-14*ic_cap*ic_cap+-5.00000e-14*ic_cap+1.42000e-11'
+ mcm5m2_cf_w_4_000_s_3_200 = '-7.50000e-14*ic_cap*ic_cap+-5.00000e-14*ic_cap+1.59000e-11'
+ mcm5m2_cf_w_4_000_s_4_800 = '-1.06250e-13*ic_cap*ic_cap+-7.50000e-14*ic_cap+2.17000e-11'
+ mcm5m2d_ca_w_0_140_s_0_140 = '-2.90625e-07*ic_cap*ic_cap+-1.87500e-07*ic_cap+3.23000e-05'
+ mcm5m2d_ca_w_0_140_s_0_175 = '-2.90625e-07*ic_cap*ic_cap+-1.87500e-07*ic_cap+3.23000e-05'
+ mcm5m2d_ca_w_0_140_s_0_210 = '-2.90625e-07*ic_cap*ic_cap+-1.87500e-07*ic_cap+3.23000e-05'
+ mcm5m2d_ca_w_0_140_s_0_280 = '-2.90625e-07*ic_cap*ic_cap+-1.87500e-07*ic_cap+3.23000e-05'
+ mcm5m2d_ca_w_0_140_s_0_350 = '-2.90625e-07*ic_cap*ic_cap+-1.87500e-07*ic_cap+3.23000e-05'
+ mcm5m2d_ca_w_0_140_s_0_420 = '-2.90625e-07*ic_cap*ic_cap+-1.87500e-07*ic_cap+3.23000e-05'
+ mcm5m2d_ca_w_0_140_s_0_560 = '-2.90625e-07*ic_cap*ic_cap+-1.87500e-07*ic_cap+3.23000e-05'
+ mcm5m2d_ca_w_0_140_s_0_840 = '-2.90625e-07*ic_cap*ic_cap+-1.87500e-07*ic_cap+3.23000e-05'
+ mcm5m2d_ca_w_0_140_s_1_540 = '-2.90625e-07*ic_cap*ic_cap+-1.87500e-07*ic_cap+3.23000e-05'
+ mcm5m2d_ca_w_0_140_s_3_500 = '-2.90625e-07*ic_cap*ic_cap+-1.87500e-07*ic_cap+3.23000e-05'
+ mcm5m2d_ca_w_1_120_s_0_140 = '-2.90625e-07*ic_cap*ic_cap+-1.87500e-07*ic_cap+3.23000e-05'
+ mcm5m2d_ca_w_1_120_s_0_175 = '-2.90625e-07*ic_cap*ic_cap+-1.87500e-07*ic_cap+3.23000e-05'
+ mcm5m2d_ca_w_1_120_s_0_210 = '-2.90625e-07*ic_cap*ic_cap+-1.87500e-07*ic_cap+3.23000e-05'
+ mcm5m2d_ca_w_1_120_s_0_280 = '-2.90625e-07*ic_cap*ic_cap+-1.87500e-07*ic_cap+3.23000e-05'
+ mcm5m2d_ca_w_1_120_s_0_350 = '-2.90625e-07*ic_cap*ic_cap+-1.87500e-07*ic_cap+3.23000e-05'
+ mcm5m2d_ca_w_1_120_s_0_420 = '-2.90625e-07*ic_cap*ic_cap+-1.87500e-07*ic_cap+3.23000e-05'
+ mcm5m2d_ca_w_1_120_s_0_560 = '-2.90625e-07*ic_cap*ic_cap+-1.87500e-07*ic_cap+3.23000e-05'
+ mcm5m2d_ca_w_1_120_s_0_840 = '-2.90625e-07*ic_cap*ic_cap+-1.87500e-07*ic_cap+3.23000e-05'
+ mcm5m2d_ca_w_1_120_s_1_540 = '-2.90625e-07*ic_cap*ic_cap+-1.87500e-07*ic_cap+3.23000e-05'
+ mcm5m2d_ca_w_1_120_s_3_500 = '-2.90625e-07*ic_cap*ic_cap+-1.87500e-07*ic_cap+3.23000e-05'
+ mcm5m2d_cc_w_0_140_s_0_140 = '-9.59375e-13*ic_cap*ic_cap+-4.62500e-13*ic_cap+1.05000e-10'
+ mcm5m2d_cc_w_0_140_s_0_175 = '-8.43750e-13*ic_cap*ic_cap+-6.50000e-13*ic_cap+1.02000e-10'
+ mcm5m2d_cc_w_0_140_s_0_210 = '-7.71875e-13*ic_cap*ic_cap+-4.62500e-13*ic_cap+9.70000e-11'
+ mcm5m2d_cc_w_0_140_s_0_280 = '-5.90625e-13*ic_cap*ic_cap+-3.62500e-13*ic_cap+8.61000e-11'
+ mcm5m2d_cc_w_0_140_s_0_350 = '-4.59375e-13*ic_cap*ic_cap+-2.62500e-13*ic_cap+7.48000e-11'
+ mcm5m2d_cc_w_0_140_s_0_420 = '-3.40625e-13*ic_cap*ic_cap+-2.37500e-13*ic_cap+6.50000e-11'
+ mcm5m2d_cc_w_0_140_s_0_560 = '-1.96875e-13*ic_cap*ic_cap+-1.37500e-13*ic_cap+5.20000e-11'
+ mcm5m2d_cc_w_0_140_s_0_840 = '-7.81250e-14*ic_cap*ic_cap+-6.25000e-14*ic_cap+3.73000e-11'
+ mcm5m2d_cc_w_0_140_s_1_540 = '3.43750e-14*ic_cap*ic_cap+1.25000e-14*ic_cap+1.99000e-11'
+ mcm5m2d_cc_w_0_140_s_3_500 = '5.40625e-14*ic_cap*ic_cap+3.62500e-14*ic_cap+5.02000e-12'
+ mcm5m2d_cc_w_1_120_s_0_140 = '-8.12500e-13*ic_cap*ic_cap+-5.00000e-13*ic_cap+1.26000e-10'
+ mcm5m2d_cc_w_1_120_s_0_175 = '-8.12500e-13*ic_cap*ic_cap+-2.50000e-13*ic_cap+1.23000e-10'
+ mcm5m2d_cc_w_1_120_s_0_210 = '-6.56250e-13*ic_cap*ic_cap+-3.75000e-13*ic_cap+1.16000e-10'
+ mcm5m2d_cc_w_1_120_s_0_280 = '-5.09375e-13*ic_cap*ic_cap+-3.87500e-13*ic_cap+1.02000e-10'
+ mcm5m2d_cc_w_1_120_s_0_350 = '-3.59375e-13*ic_cap*ic_cap+-2.37500e-13*ic_cap+8.90000e-11'
+ mcm5m2d_cc_w_1_120_s_0_420 = '-2.62500e-13*ic_cap*ic_cap+-1.50000e-13*ic_cap+7.81000e-11'
+ mcm5m2d_cc_w_1_120_s_0_560 = '-1.06250e-13*ic_cap*ic_cap+-7.50000e-14*ic_cap+6.25000e-11'
+ mcm5m2d_cc_w_1_120_s_0_840 = '3.12500e-15*ic_cap*ic_cap+-1.25000e-14*ic_cap+4.46000e-11'
+ mcm5m2d_cc_w_1_120_s_1_540 = '8.43750e-14*ic_cap*ic_cap+6.25000e-14*ic_cap+2.43000e-11'
+ mcm5m2d_cc_w_1_120_s_3_500 = '7.87500e-14*ic_cap*ic_cap+5.50000e-14*ic_cap+6.40000e-12'
+ mcm5m2d_cf_w_0_140_s_0_140 = '1.56250e-15*ic_cap*ic_cap+1.25000e-15*ic_cap+2.25000e-12'
+ mcm5m2d_cf_w_0_140_s_0_175 = '-3.75000e-15*ic_cap*ic_cap+-2.50000e-15*ic_cap+2.81000e-12'
+ mcm5m2d_cf_w_0_140_s_0_210 = '-7.50000e-15*ic_cap*ic_cap+-5.00000e-15*ic_cap+3.37000e-12'
+ mcm5m2d_cf_w_0_140_s_0_280 = '-1.84375e-14*ic_cap*ic_cap+-1.37500e-14*ic_cap+4.48000e-12'
+ mcm5m2d_cf_w_0_140_s_0_350 = '-2.87500e-14*ic_cap*ic_cap+-1.75000e-14*ic_cap+5.57000e-12'
+ mcm5m2d_cf_w_0_140_s_0_420 = '-3.75000e-14*ic_cap*ic_cap+-2.75000e-14*ic_cap+6.67000e-12'
+ mcm5m2d_cf_w_0_140_s_0_560 = '-5.62500e-14*ic_cap*ic_cap+-3.50000e-14*ic_cap+8.75000e-12'
+ mcm5m2d_cf_w_0_140_s_0_840 = '-9.06250e-14*ic_cap*ic_cap+-6.25000e-14*ic_cap+1.26000e-11'
+ mcm5m2d_cf_w_0_140_s_1_540 = '-1.50000e-13*ic_cap*ic_cap+-1.00000e-13*ic_cap+2.05000e-11'
+ mcm5m2d_cf_w_0_140_s_3_500 = '-1.87500e-13*ic_cap*ic_cap+-1.25000e-13*ic_cap+3.15000e-11'
+ mcm5m2d_cf_w_1_120_s_0_140 = '1.25000e-15*ic_cap*ic_cap+2.28000e-12'
+ mcm5m2d_cf_w_1_120_s_0_175 = '-4.37500e-15*ic_cap*ic_cap+-2.50000e-15*ic_cap+2.85000e-12'
+ mcm5m2d_cf_w_1_120_s_0_210 = '-9.06250e-15*ic_cap*ic_cap+-6.25000e-15*ic_cap+3.40000e-12'
+ mcm5m2d_cf_w_1_120_s_0_280 = '-1.90625e-14*ic_cap*ic_cap+-1.37500e-14*ic_cap+4.51000e-12'
+ mcm5m2d_cf_w_1_120_s_0_350 = '-2.87500e-14*ic_cap*ic_cap+-2.00000e-14*ic_cap+5.61000e-12'
+ mcm5m2d_cf_w_1_120_s_0_420 = '-3.87500e-14*ic_cap*ic_cap+-2.50000e-14*ic_cap+6.69000e-12'
+ mcm5m2d_cf_w_1_120_s_0_560 = '-5.71875e-14*ic_cap*ic_cap+-3.62500e-14*ic_cap+8.79000e-12'
+ mcm5m2d_cf_w_1_120_s_0_840 = '-9.37500e-14*ic_cap*ic_cap+-5.00000e-14*ic_cap+1.28000e-11'
+ mcm5m2d_cf_w_1_120_s_1_540 = '-1.56250e-13*ic_cap*ic_cap+-1.00000e-13*ic_cap+2.11000e-11'
+ mcm5m2d_cf_w_1_120_s_3_500 = '-1.93750e-13*ic_cap*ic_cap+-1.25000e-13*ic_cap+3.37000e-11'
+ mcm5m2f_ca_w_0_140_s_0_140 = '-2.71875e-07*ic_cap*ic_cap+-1.62500e-07*ic_cap+2.91000e-05'
+ mcm5m2f_ca_w_0_140_s_0_175 = '-2.71875e-07*ic_cap*ic_cap+-1.62500e-07*ic_cap+2.91000e-05'
+ mcm5m2f_ca_w_0_140_s_0_210 = '-2.71875e-07*ic_cap*ic_cap+-1.62500e-07*ic_cap+2.91000e-05'
+ mcm5m2f_ca_w_0_140_s_0_280 = '-2.71875e-07*ic_cap*ic_cap+-1.62500e-07*ic_cap+2.91000e-05'
+ mcm5m2f_ca_w_0_140_s_0_350 = '-2.71875e-07*ic_cap*ic_cap+-1.62500e-07*ic_cap+2.91000e-05'
+ mcm5m2f_ca_w_0_140_s_0_420 = '-2.71875e-07*ic_cap*ic_cap+-1.62500e-07*ic_cap+2.91000e-05'
+ mcm5m2f_ca_w_0_140_s_0_560 = '-2.71875e-07*ic_cap*ic_cap+-1.62500e-07*ic_cap+2.91000e-05'
+ mcm5m2f_ca_w_0_140_s_0_840 = '-2.71875e-07*ic_cap*ic_cap+-1.62500e-07*ic_cap+2.91000e-05'
+ mcm5m2f_ca_w_0_140_s_1_540 = '-2.71875e-07*ic_cap*ic_cap+-1.62500e-07*ic_cap+2.91000e-05'
+ mcm5m2f_ca_w_0_140_s_3_500 = '-2.71875e-07*ic_cap*ic_cap+-1.62500e-07*ic_cap+2.91000e-05'
+ mcm5m2f_ca_w_1_120_s_0_140 = '-2.71875e-07*ic_cap*ic_cap+-1.62500e-07*ic_cap+2.91000e-05'
+ mcm5m2f_ca_w_1_120_s_0_175 = '-2.71875e-07*ic_cap*ic_cap+-1.62500e-07*ic_cap+2.91000e-05'
+ mcm5m2f_ca_w_1_120_s_0_210 = '-2.71875e-07*ic_cap*ic_cap+-1.62500e-07*ic_cap+2.91000e-05'
+ mcm5m2f_ca_w_1_120_s_0_280 = '-2.71875e-07*ic_cap*ic_cap+-1.62500e-07*ic_cap+2.91000e-05'
+ mcm5m2f_ca_w_1_120_s_0_350 = '-2.71875e-07*ic_cap*ic_cap+-1.62500e-07*ic_cap+2.91000e-05'
+ mcm5m2f_ca_w_1_120_s_0_420 = '-2.71875e-07*ic_cap*ic_cap+-1.62500e-07*ic_cap+2.91000e-05'
+ mcm5m2f_ca_w_1_120_s_0_560 = '-2.71875e-07*ic_cap*ic_cap+-1.62500e-07*ic_cap+2.91000e-05'
+ mcm5m2f_ca_w_1_120_s_0_840 = '-2.71875e-07*ic_cap*ic_cap+-1.62500e-07*ic_cap+2.91000e-05'
+ mcm5m2f_ca_w_1_120_s_1_540 = '-2.71875e-07*ic_cap*ic_cap+-1.62500e-07*ic_cap+2.91000e-05'
+ mcm5m2f_ca_w_1_120_s_3_500 = '-2.71875e-07*ic_cap*ic_cap+-1.62500e-07*ic_cap+2.91000e-05'
+ mcm5m2f_cc_w_0_140_s_0_140 = '-9.40625e-13*ic_cap*ic_cap+-4.87500e-13*ic_cap+1.05000e-10'
+ mcm5m2f_cc_w_0_140_s_0_175 = '-8.87500e-13*ic_cap*ic_cap+-6.75000e-13*ic_cap+1.03000e-10'
+ mcm5m2f_cc_w_0_140_s_0_210 = '-7.62500e-13*ic_cap*ic_cap+-4.50000e-13*ic_cap+9.74000e-11'
+ mcm5m2f_cc_w_0_140_s_0_280 = '-5.96875e-13*ic_cap*ic_cap+-3.62500e-13*ic_cap+8.66000e-11'
+ mcm5m2f_cc_w_0_140_s_0_350 = '-4.65625e-13*ic_cap*ic_cap+-2.62500e-13*ic_cap+7.55000e-11'
+ mcm5m2f_cc_w_0_140_s_0_420 = '-3.59375e-13*ic_cap*ic_cap+-2.62500e-13*ic_cap+6.59000e-11'
+ mcm5m2f_cc_w_0_140_s_0_560 = '-1.90625e-13*ic_cap*ic_cap+-1.37500e-13*ic_cap+5.27000e-11'
+ mcm5m2f_cc_w_0_140_s_0_840 = '-7.81250e-14*ic_cap*ic_cap+-6.25000e-14*ic_cap+3.83000e-11'
+ mcm5m2f_cc_w_0_140_s_1_540 = '2.81250e-14*ic_cap*ic_cap+1.25000e-14*ic_cap+2.12000e-11'
+ mcm5m2f_cc_w_0_140_s_3_500 = '5.84375e-14*ic_cap*ic_cap+3.87500e-14*ic_cap+5.84000e-12'
+ mcm5m2f_cc_w_1_120_s_0_140 = '-8.12500e-13*ic_cap*ic_cap+-5.00000e-13*ic_cap+1.27000e-10'
+ mcm5m2f_cc_w_1_120_s_0_175 = '-8.12500e-13*ic_cap*ic_cap+-2.50000e-13*ic_cap+1.24000e-10'
+ mcm5m2f_cc_w_1_120_s_0_210 = '-5.93750e-13*ic_cap*ic_cap+-3.75000e-13*ic_cap+1.17000e-10'
+ mcm5m2f_cc_w_1_120_s_0_280 = '-4.84375e-13*ic_cap*ic_cap+-3.87500e-13*ic_cap+1.03000e-10'
+ mcm5m2f_cc_w_1_120_s_0_350 = '-3.78125e-13*ic_cap*ic_cap+-2.12500e-13*ic_cap+9.06000e-11'
+ mcm5m2f_cc_w_1_120_s_0_420 = '-2.65625e-13*ic_cap*ic_cap+-1.62500e-13*ic_cap+7.97000e-11'
+ mcm5m2f_cc_w_1_120_s_0_560 = '-1.12500e-13*ic_cap*ic_cap+-7.50000e-14*ic_cap+6.41000e-11'
+ mcm5m2f_cc_w_1_120_s_1_540 = '9.06250e-14*ic_cap*ic_cap+6.25000e-14*ic_cap+2.59000e-11'
+ mcm5m2f_cc_w_1_120_s_3_500 = '9.18750e-14*ic_cap*ic_cap+6.00000e-14*ic_cap+7.36000e-12'
+ mcm5m2f_cf_w_0_140_s_0_140 = '1.25000e-15*ic_cap*ic_cap+2.02000e-12'
+ mcm5m2f_cf_w_0_140_s_0_175 = '-3.75000e-15*ic_cap*ic_cap+-2.50000e-15*ic_cap+2.52000e-12'
+ mcm5m2f_cf_w_0_140_s_0_210 = '-7.18750e-15*ic_cap*ic_cap+-3.75000e-15*ic_cap+3.03000e-12'
+ mcm5m2f_cf_w_0_140_s_0_280 = '-1.75000e-14*ic_cap*ic_cap+-1.25000e-14*ic_cap+4.03000e-12'
+ mcm5m2f_cf_w_0_140_s_0_350 = '-2.65625e-14*ic_cap*ic_cap+-1.62500e-14*ic_cap+5.00000e-12'
+ mcm5m2f_cf_w_0_140_s_0_420 = '-3.59375e-14*ic_cap*ic_cap+-2.37500e-14*ic_cap+6.02000e-12'
+ mcm5m2f_cf_w_0_140_s_0_560 = '-5.15625e-14*ic_cap*ic_cap+-3.12500e-14*ic_cap+7.88000e-12'
+ mcm5m2f_cf_w_0_140_s_0_840 = '-8.28125e-14*ic_cap*ic_cap+-5.62500e-14*ic_cap+1.14000e-11'
+ mcm5m2f_cf_w_0_140_s_1_540 = '-1.46875e-13*ic_cap*ic_cap+-8.75000e-14*ic_cap+1.88000e-11'
+ mcm5m2f_cf_w_0_140_s_3_500 = '-1.87500e-13*ic_cap*ic_cap+-1.25000e-13*ic_cap+2.97000e-11'
+ mcm5m2f_cf_w_1_120_s_0_140 = '9.37500e-16*ic_cap*ic_cap+1.25000e-15*ic_cap+2.04000e-12'
+ mcm5m2f_cf_w_1_120_s_0_175 = '-4.06250e-15*ic_cap*ic_cap+-3.75000e-15*ic_cap+2.55000e-12'
+ mcm5m2f_cf_w_1_120_s_0_210 = '-8.43750e-15*ic_cap*ic_cap+-6.25000e-15*ic_cap+3.05000e-12'
+ mcm5m2f_cf_w_1_120_s_0_280 = '-1.78125e-14*ic_cap*ic_cap+-1.12500e-14*ic_cap+4.05000e-12'
+ mcm5m2f_cf_w_1_120_s_0_350 = '-2.65625e-14*ic_cap*ic_cap+-1.62500e-14*ic_cap+5.03000e-12'
+ mcm5m2f_cf_w_1_120_s_0_420 = '-3.68750e-14*ic_cap*ic_cap+-2.25000e-14*ic_cap+6.03000e-12'
+ mcm5m2f_cf_w_1_120_s_0_560 = '-5.28125e-14*ic_cap*ic_cap+-3.37500e-14*ic_cap+7.91000e-12'
+ mcm5m2f_cf_w_1_120_s_0_840 = '-8.25000e-14*ic_cap*ic_cap+-5.50000e-14*ic_cap+1.15000e-11'
+ mcm5m2f_cf_w_1_120_s_1_540 = '-1.40625e-13*ic_cap*ic_cap+-8.75000e-14*ic_cap+1.92000e-11'
+ mcm5m2f_cf_w_1_120_s_3_500 = '-1.87500e-13*ic_cap*ic_cap+-1.25000e-13*ic_cap+3.17000e-11'
+ mcm5m2l1_ca_w_0_140_s_0_140 = '-5.28125e-07*ic_cap*ic_cap+-3.37500e-07*ic_cap+4.85000e-05'
+ mcm5m2l1_ca_w_0_140_s_0_175 = '-5.28125e-07*ic_cap*ic_cap+-3.37500e-07*ic_cap+4.85000e-05'
+ mcm5m2l1_ca_w_0_140_s_0_210 = '-5.28125e-07*ic_cap*ic_cap+-3.37500e-07*ic_cap+4.85000e-05'
+ mcm5m2l1_ca_w_0_140_s_0_280 = '-5.28125e-07*ic_cap*ic_cap+-3.37500e-07*ic_cap+4.85000e-05'
+ mcm5m2l1_ca_w_0_140_s_0_350 = '-5.28125e-07*ic_cap*ic_cap+-3.37500e-07*ic_cap+4.85000e-05'
+ mcm5m2l1_ca_w_0_140_s_0_420 = '-5.28125e-07*ic_cap*ic_cap+-3.37500e-07*ic_cap+4.85000e-05'
+ mcm5m2l1_ca_w_0_140_s_0_560 = '-5.28125e-07*ic_cap*ic_cap+-3.37500e-07*ic_cap+4.85000e-05'
+ mcm5m2l1_ca_w_0_140_s_0_840 = '-5.28125e-07*ic_cap*ic_cap+-3.37500e-07*ic_cap+4.85000e-05'
+ mcm5m2l1_ca_w_0_140_s_1_540 = '-5.28125e-07*ic_cap*ic_cap+-3.37500e-07*ic_cap+4.85000e-05'
+ mcm5m2l1_ca_w_0_140_s_3_500 = '-5.28125e-07*ic_cap*ic_cap+-3.37500e-07*ic_cap+4.85000e-05'
+ mcm5m2l1_ca_w_1_120_s_0_140 = '-5.28125e-07*ic_cap*ic_cap+-3.37500e-07*ic_cap+4.85000e-05'
+ mcm5m2l1_ca_w_1_120_s_0_175 = '-5.28125e-07*ic_cap*ic_cap+-3.37500e-07*ic_cap+4.85000e-05'
+ mcm5m2l1_ca_w_1_120_s_0_210 = '-5.28125e-07*ic_cap*ic_cap+-3.37500e-07*ic_cap+4.85000e-05'
+ mcm5m2l1_ca_w_1_120_s_0_280 = '-5.28125e-07*ic_cap*ic_cap+-3.37500e-07*ic_cap+4.85000e-05'
+ mcm5m2l1_ca_w_1_120_s_0_350 = '-5.28125e-07*ic_cap*ic_cap+-3.37500e-07*ic_cap+4.85000e-05'
+ mcm5m2l1_ca_w_1_120_s_0_420 = '-5.28125e-07*ic_cap*ic_cap+-3.37500e-07*ic_cap+4.85000e-05'
+ mcm5m2l1_ca_w_1_120_s_0_560 = '-5.28125e-07*ic_cap*ic_cap+-3.37500e-07*ic_cap+4.85000e-05'
+ mcm5m2l1_ca_w_1_120_s_0_840 = '-5.28125e-07*ic_cap*ic_cap+-3.37500e-07*ic_cap+4.85000e-05'
+ mcm5m2l1_ca_w_1_120_s_1_540 = '-5.28125e-07*ic_cap*ic_cap+-3.37500e-07*ic_cap+4.85000e-05'
+ mcm5m2l1_ca_w_1_120_s_3_500 = '-5.28125e-07*ic_cap*ic_cap+-3.37500e-07*ic_cap+4.85000e-05'
+ mcm5m2l1_cc_w_0_140_s_0_140 = '-8.81250e-13*ic_cap*ic_cap+-5.25000e-13*ic_cap+1.02000e-10'
+ mcm5m2l1_cc_w_0_140_s_0_175 = '-8.09375e-13*ic_cap*ic_cap+-5.87500e-13*ic_cap+1.00000e-10'
+ mcm5m2l1_cc_w_0_140_s_0_210 = '-7.37500e-13*ic_cap*ic_cap+-4.50000e-13*ic_cap+9.47000e-11'
+ mcm5m2l1_cc_w_0_140_s_0_280 = '-5.56250e-13*ic_cap*ic_cap+-3.25000e-13*ic_cap+8.34000e-11'
+ mcm5m2l1_cc_w_0_140_s_0_350 = '-3.81250e-13*ic_cap*ic_cap+-2.50000e-13*ic_cap+7.14000e-11'
+ mcm5m2l1_cc_w_0_140_s_0_420 = '-2.75000e-13*ic_cap*ic_cap+-1.75000e-13*ic_cap+6.13000e-11'
+ mcm5m2l1_cc_w_0_140_s_0_560 = '-1.56250e-13*ic_cap*ic_cap+-1.25000e-13*ic_cap+4.83000e-11'
+ mcm5m2l1_cc_w_0_140_s_0_840 = '-2.50000e-14*ic_cap*ic_cap+-2.50000e-14*ic_cap+3.27000e-11'
+ mcm5m2l1_cc_w_0_140_s_1_540 = '5.93750e-14*ic_cap*ic_cap+3.75000e-14*ic_cap+1.56000e-11'
+ mcm5m2l1_cc_w_0_140_s_3_500 = '4.46875e-14*ic_cap*ic_cap+3.37500e-14*ic_cap+2.91000e-12'
+ mcm5m2l1_cc_w_1_120_s_0_140 = '-7.50000e-13*ic_cap*ic_cap+-5.00000e-13*ic_cap+1.20000e-10'
+ mcm5m2l1_cc_w_1_120_s_0_175 = '-7.18750e-13*ic_cap*ic_cap+-3.75000e-13*ic_cap+1.17000e-10'
+ mcm5m2l1_cc_w_1_120_s_0_210 = '-5.84375e-13*ic_cap*ic_cap+-3.37500e-13*ic_cap+1.10000e-10'
+ mcm5m2l1_cc_w_1_120_s_0_280 = '-4.09375e-13*ic_cap*ic_cap+-2.87500e-13*ic_cap+9.58000e-11'
+ mcm5m2l1_cc_w_1_120_s_0_350 = '-2.93750e-13*ic_cap*ic_cap+-2.25000e-13*ic_cap+8.29000e-11'
+ mcm5m2l1_cc_w_1_120_s_0_420 = '-1.78125e-13*ic_cap*ic_cap+-1.37500e-13*ic_cap+7.19000e-11'
+ mcm5m2l1_cc_w_1_120_s_0_560 = '-6.25000e-14*ic_cap*ic_cap+-5.00000e-14*ic_cap+5.65000e-11'
+ mcm5m2l1_cc_w_1_120_s_0_840 = '3.75000e-14*ic_cap*ic_cap+2.50000e-14*ic_cap+3.88000e-11'
+ mcm5m2l1_cc_w_1_120_s_1_540 = '1.00000e-13*ic_cap*ic_cap+7.50000e-14*ic_cap+1.90000e-11'
+ mcm5m2l1_cc_w_1_120_s_3_500 = '6.59375e-14*ic_cap*ic_cap+5.12500e-14*ic_cap+3.81000e-12'
+ mcm5m2l1_cf_w_0_140_s_0_140 = '-4.37500e-15*ic_cap*ic_cap+-5.00000e-15*ic_cap+3.34000e-12'
+ mcm5m2l1_cf_w_0_140_s_0_175 = '-1.37500e-14*ic_cap*ic_cap+-1.00000e-14*ic_cap+4.18000e-12'
+ mcm5m2l1_cf_w_0_140_s_0_210 = '-2.15625e-14*ic_cap*ic_cap+-1.62500e-14*ic_cap+5.02000e-12'
+ mcm5m2l1_cf_w_0_140_s_0_280 = '-4.03125e-14*ic_cap*ic_cap+-2.87500e-14*ic_cap+6.66000e-12'
+ mcm5m2l1_cf_w_0_140_s_0_350 = '-5.71875e-14*ic_cap*ic_cap+-3.87500e-14*ic_cap+8.25000e-12'
+ mcm5m2l1_cf_w_0_140_s_0_420 = '-7.28125e-14*ic_cap*ic_cap+-5.12500e-14*ic_cap+9.85000e-12'
+ mcm5m2l1_cf_w_0_140_s_0_560 = '-1.03125e-13*ic_cap*ic_cap+-6.25000e-14*ic_cap+1.28000e-11'
+ mcm5m2l1_cf_w_0_140_s_0_840 = '-1.56250e-13*ic_cap*ic_cap+-1.00000e-13*ic_cap+1.81000e-11'
+ mcm5m2l1_cf_w_0_140_s_1_540 = '-2.31250e-13*ic_cap*ic_cap+-1.50000e-13*ic_cap+2.80000e-11'
+ mcm5m2l1_cf_w_0_140_s_3_500 = '-2.40625e-13*ic_cap*ic_cap+-1.62500e-13*ic_cap+3.85000e-11'
+ mcm5m2l1_cf_w_1_120_s_0_140 = '-4.37500e-15*ic_cap*ic_cap+-5.00000e-15*ic_cap+3.37000e-12'
+ mcm5m2l1_cf_w_1_120_s_0_175 = '-1.40625e-14*ic_cap*ic_cap+-1.12500e-14*ic_cap+4.22000e-12'
+ mcm5m2l1_cf_w_1_120_s_0_210 = '-2.34375e-14*ic_cap*ic_cap+-1.62500e-14*ic_cap+5.05000e-12'
+ mcm5m2l1_cf_w_1_120_s_0_280 = '-3.96875e-14*ic_cap*ic_cap+-2.62500e-14*ic_cap+6.69000e-12'
+ mcm5m2l1_cf_w_1_120_s_0_350 = '-5.78125e-14*ic_cap*ic_cap+-3.87500e-14*ic_cap+8.30000e-12'
+ mcm5m2l1_cf_w_1_120_s_0_420 = '-7.43750e-14*ic_cap*ic_cap+-5.00000e-14*ic_cap+9.87000e-12'
+ mcm5m2l1_cf_w_1_120_s_0_560 = '-1.06250e-13*ic_cap*ic_cap+-7.50000e-14*ic_cap+1.29000e-11'
+ mcm5m2l1_cf_w_1_120_s_0_840 = '-1.56250e-13*ic_cap*ic_cap+-1.00000e-13*ic_cap+1.83000e-11'
+ mcm5m2l1_cf_w_1_120_s_1_540 = '-2.31250e-13*ic_cap*ic_cap+-1.50000e-13*ic_cap+2.87000e-11'
+ mcm5m2l1_cf_w_1_120_s_3_500 = '-2.34375e-13*ic_cap*ic_cap+-1.62500e-13*ic_cap+4.09000e-11'
+ mcm5m2m1_ca_w_0_140_s_0_140 = '-2.70312e-06*ic_cap*ic_cap+-1.31250e-06*ic_cap+1.39000e-04'
+ mcm5m2m1_ca_w_0_140_s_0_175 = '-2.70312e-06*ic_cap*ic_cap+-1.31250e-06*ic_cap+1.39000e-04'
+ mcm5m2m1_ca_w_0_140_s_0_210 = '-2.70312e-06*ic_cap*ic_cap+-1.31250e-06*ic_cap+1.39000e-04'
+ mcm5m2m1_ca_w_0_140_s_0_280 = '-2.70312e-06*ic_cap*ic_cap+-1.31250e-06*ic_cap+1.39000e-04'
+ mcm5m2m1_ca_w_0_140_s_0_350 = '-2.70312e-06*ic_cap*ic_cap+-1.31250e-06*ic_cap+1.39000e-04'
+ mcm5m2m1_ca_w_0_140_s_0_420 = '-2.70312e-06*ic_cap*ic_cap+-1.31250e-06*ic_cap+1.39000e-04'
+ mcm5m2m1_ca_w_0_140_s_0_560 = '-2.70312e-06*ic_cap*ic_cap+-1.31250e-06*ic_cap+1.39000e-04'
+ mcm5m2m1_ca_w_0_140_s_0_840 = '-2.70312e-06*ic_cap*ic_cap+-1.31250e-06*ic_cap+1.39000e-04'
+ mcm5m2m1_ca_w_0_140_s_1_540 = '-2.70312e-06*ic_cap*ic_cap+-1.31250e-06*ic_cap+1.39000e-04'
+ mcm5m2m1_ca_w_0_140_s_3_500 = '-2.70312e-06*ic_cap*ic_cap+-1.31250e-06*ic_cap+1.39000e-04'
+ mcm5m2m1_ca_w_1_120_s_0_140 = '-2.70312e-06*ic_cap*ic_cap+-1.31250e-06*ic_cap+1.39000e-04'
+ mcm5m2m1_ca_w_1_120_s_0_175 = '-2.70312e-06*ic_cap*ic_cap+-1.31250e-06*ic_cap+1.39000e-04'
+ mcm5m2m1_ca_w_1_120_s_0_210 = '-2.70312e-06*ic_cap*ic_cap+-1.31250e-06*ic_cap+1.39000e-04'
+ mcm5m2m1_ca_w_1_120_s_0_280 = '-2.70312e-06*ic_cap*ic_cap+-1.31250e-06*ic_cap+1.39000e-04'
+ mcm5m2m1_ca_w_1_120_s_0_350 = '-2.70312e-06*ic_cap*ic_cap+-1.31250e-06*ic_cap+1.39000e-04'
+ mcm5m2m1_ca_w_1_120_s_0_420 = '-2.70312e-06*ic_cap*ic_cap+-1.31250e-06*ic_cap+1.39000e-04'
+ mcm5m2m1_ca_w_1_120_s_0_560 = '-2.70312e-06*ic_cap*ic_cap+-1.31250e-06*ic_cap+1.39000e-04'
+ mcm5m2m1_ca_w_1_120_s_0_840 = '-2.70312e-06*ic_cap*ic_cap+-1.31250e-06*ic_cap+1.39000e-04'
+ mcm5m2m1_ca_w_1_120_s_1_540 = '-2.70312e-06*ic_cap*ic_cap+-1.31250e-06*ic_cap+1.39000e-04'
+ mcm5m2m1_ca_w_1_120_s_3_500 = '-2.70312e-06*ic_cap*ic_cap+-1.31250e-06*ic_cap+1.39000e-04'
+ mcm5m2m1_cc_w_0_140_s_0_140 = '-7.71875e-13*ic_cap*ic_cap+-3.37500e-13*ic_cap+9.44000e-11'
+ mcm5m2m1_cc_w_0_140_s_0_175 = '-7.09375e-13*ic_cap*ic_cap+-3.37500e-13*ic_cap+9.18000e-11'
+ mcm5m2m1_cc_w_0_140_s_0_210 = '-5.84375e-13*ic_cap*ic_cap+-3.12500e-13*ic_cap+8.57000e-11'
+ mcm5m2m1_cc_w_0_140_s_0_280 = '-3.53125e-13*ic_cap*ic_cap+-2.62500e-13*ic_cap+7.29000e-11'
+ mcm5m2m1_cc_w_0_140_s_0_350 = '-2.28125e-13*ic_cap*ic_cap+-2.37500e-13*ic_cap+6.06000e-11'
+ mcm5m2m1_cc_w_0_140_s_0_420 = '-1.28125e-13*ic_cap*ic_cap+-1.12500e-13*ic_cap+5.08000e-11'
+ mcm5m2m1_cc_w_0_140_s_0_560 = '-6.25000e-15*ic_cap*ic_cap+-2.50000e-14*ic_cap+3.70000e-11'
+ mcm5m2m1_cc_w_0_140_s_0_840 = '8.12500e-14*ic_cap*ic_cap+2.50000e-14*ic_cap+2.21000e-11'
+ mcm5m2m1_cc_w_0_140_s_1_540 = '7.75000e-14*ic_cap*ic_cap+5.00000e-14*ic_cap+8.08000e-12'
+ mcm5m2m1_cc_w_0_140_s_3_500 = '2.03125e-14*ic_cap*ic_cap+1.62500e-14*ic_cap+1.04000e-12'
+ mcm5m2m1_cc_w_1_120_s_0_140 = '-5.62500e-13*ic_cap*ic_cap+-3.50000e-13*ic_cap+1.06000e-10'
+ mcm5m2m1_cc_w_1_120_s_0_175 = '-5.62500e-13*ic_cap*ic_cap+-2.25000e-13*ic_cap+1.03000e-10'
+ mcm5m2m1_cc_w_1_120_s_0_210 = '-4.56250e-13*ic_cap*ic_cap+-3.00000e-13*ic_cap+9.69000e-11'
+ mcm5m2m1_cc_w_1_120_s_0_280 = '-2.90625e-13*ic_cap*ic_cap+-1.62500e-13*ic_cap+8.26000e-11'
+ mcm5m2m1_cc_w_1_120_s_0_350 = '-1.56250e-13*ic_cap*ic_cap+-1.25000e-13*ic_cap+6.94000e-11'
+ mcm5m2m1_cc_w_1_120_s_0_420 = '-5.93750e-14*ic_cap*ic_cap+-3.75000e-14*ic_cap+5.87000e-11'
+ mcm5m2m1_cc_w_1_120_s_0_560 = '5.31250e-14*ic_cap*ic_cap+1.25000e-14*ic_cap+4.37000e-11'
+ mcm5m2m1_cc_w_1_120_s_0_840 = '1.15625e-13*ic_cap*ic_cap+6.25000e-14*ic_cap+2.73000e-11'
+ mcm5m2m1_cc_w_1_120_s_1_540 = '1.09375e-13*ic_cap*ic_cap+6.25000e-14*ic_cap+1.10000e-11'
+ mcm5m2m1_cc_w_1_120_s_3_500 = '3.56250e-14*ic_cap*ic_cap+2.25000e-14*ic_cap+1.59000e-12'
+ mcm5m2m1_cf_w_0_140_s_0_140 = '-9.87500e-14*ic_cap*ic_cap+-4.50000e-14*ic_cap+9.06000e-12'
+ mcm5m2m1_cf_w_0_140_s_0_175 = '-1.41563e-13*ic_cap*ic_cap+-6.62500e-14*ic_cap+1.14000e-11'
+ mcm5m2m1_cf_w_0_140_s_0_210 = '-1.84375e-13*ic_cap*ic_cap+-8.75000e-14*ic_cap+1.37000e-11'
+ mcm5m2m1_cf_w_0_140_s_0_280 = '-2.68750e-13*ic_cap*ic_cap+-1.25000e-13*ic_cap+1.81000e-11'
+ mcm5m2m1_cf_w_0_140_s_0_350 = '-3.34375e-13*ic_cap*ic_cap+-1.62500e-13*ic_cap+2.20000e-11'
+ mcm5m2m1_cf_w_0_140_s_0_420 = '-4.00000e-13*ic_cap*ic_cap+-2.00000e-13*ic_cap+2.58000e-11'
+ mcm5m2m1_cf_w_0_140_s_0_560 = '-4.81250e-13*ic_cap*ic_cap+-2.50000e-13*ic_cap+3.20000e-11'
+ mcm5m2m1_cf_w_0_140_s_0_840 = '-5.87500e-13*ic_cap*ic_cap+-3.00000e-13*ic_cap+4.14000e-11'
+ mcm5m2m1_cf_w_0_140_s_1_540 = '-6.43750e-13*ic_cap*ic_cap+-3.50000e-13*ic_cap+5.33000e-11'
+ mcm5m2m1_cf_w_0_140_s_3_500 = '-6.18750e-13*ic_cap*ic_cap+-3.25000e-13*ic_cap+6.04000e-11'
+ mcm5m2m1_cf_w_1_120_s_0_140 = '-9.71875e-14*ic_cap*ic_cap+-4.62500e-14*ic_cap+9.04000e-12'
+ mcm5m2m1_cf_w_1_120_s_0_175 = '-1.46875e-13*ic_cap*ic_cap+-6.75000e-14*ic_cap+1.15000e-11'
+ mcm5m2m1_cf_w_1_120_s_0_210 = '-1.84375e-13*ic_cap*ic_cap+-8.75000e-14*ic_cap+1.37000e-11'
+ mcm5m2m1_cf_w_1_120_s_0_280 = '-2.62500e-13*ic_cap*ic_cap+-1.25000e-13*ic_cap+1.80000e-11'
+ mcm5m2m1_cf_w_1_120_s_0_350 = '-3.31250e-13*ic_cap*ic_cap+-1.75000e-13*ic_cap+2.20000e-11'
+ mcm5m2m1_cf_w_1_120_s_0_420 = '-3.93750e-13*ic_cap*ic_cap+-1.75000e-13*ic_cap+2.57000e-11'
+ mcm5m2m1_cf_w_1_120_s_0_560 = '-4.78125e-13*ic_cap*ic_cap+-2.37500e-13*ic_cap+3.20000e-11'
+ mcm5m2m1_cf_w_1_120_s_0_840 = '-5.90625e-13*ic_cap*ic_cap+-3.12500e-13*ic_cap+4.17000e-11'
+ mcm5m2m1_cf_w_1_120_s_1_540 = '-6.46875e-13*ic_cap*ic_cap+-3.62500e-13*ic_cap+5.46000e-11'
+ mcm5m2m1_cf_w_1_120_s_3_500 = '-6.09375e-13*ic_cap*ic_cap+-3.37500e-13*ic_cap+6.38000e-11'
+ mcm5m2p1_ca_w_0_140_s_0_140 = '-3.90625e-07*ic_cap*ic_cap+-2.37500e-07*ic_cap+3.62000e-05'
+ mcm5m2p1_ca_w_0_140_s_0_175 = '-3.90625e-07*ic_cap*ic_cap+-2.37500e-07*ic_cap+3.62000e-05'
+ mcm5m2p1_ca_w_0_140_s_0_210 = '-3.90625e-07*ic_cap*ic_cap+-2.37500e-07*ic_cap+3.62000e-05'
+ mcm5m2p1_ca_w_0_140_s_0_280 = '-3.90625e-07*ic_cap*ic_cap+-2.37500e-07*ic_cap+3.62000e-05'
+ mcm5m2p1_ca_w_0_140_s_0_350 = '-3.90625e-07*ic_cap*ic_cap+-2.37500e-07*ic_cap+3.62000e-05'
+ mcm5m2p1_ca_w_0_140_s_0_420 = '-3.90625e-07*ic_cap*ic_cap+-2.37500e-07*ic_cap+3.62000e-05'
+ mcm5m2p1_ca_w_0_140_s_0_560 = '-3.90625e-07*ic_cap*ic_cap+-2.37500e-07*ic_cap+3.62000e-05'
+ mcm5m2p1_ca_w_0_140_s_0_840 = '-3.90625e-07*ic_cap*ic_cap+-2.37500e-07*ic_cap+3.62000e-05'
+ mcm5m2p1_ca_w_0_140_s_1_540 = '-3.90625e-07*ic_cap*ic_cap+-2.37500e-07*ic_cap+3.62000e-05'
+ mcm5m2p1_ca_w_0_140_s_3_500 = '-3.90625e-07*ic_cap*ic_cap+-2.37500e-07*ic_cap+3.62000e-05'
+ mcm5m2p1_ca_w_1_120_s_0_140 = '-3.90625e-07*ic_cap*ic_cap+-2.37500e-07*ic_cap+3.62000e-05'
+ mcm5m2p1_ca_w_1_120_s_0_175 = '-3.90625e-07*ic_cap*ic_cap+-2.37500e-07*ic_cap+3.62000e-05'
+ mcm5m2p1_ca_w_1_120_s_0_210 = '-3.90625e-07*ic_cap*ic_cap+-2.37500e-07*ic_cap+3.62000e-05'
+ mcm5m2p1_ca_w_1_120_s_0_280 = '-3.90625e-07*ic_cap*ic_cap+-2.37500e-07*ic_cap+3.62000e-05'
+ mcm5m2p1_ca_w_1_120_s_0_350 = '-3.90625e-07*ic_cap*ic_cap+-2.37500e-07*ic_cap+3.62000e-05'
+ mcm5m2p1_ca_w_1_120_s_0_420 = '-3.90625e-07*ic_cap*ic_cap+-2.37500e-07*ic_cap+3.62000e-05'
+ mcm5m2p1_ca_w_1_120_s_0_560 = '-3.90625e-07*ic_cap*ic_cap+-2.37500e-07*ic_cap+3.62000e-05'
+ mcm5m2p1_ca_w_1_120_s_0_840 = '-3.90625e-07*ic_cap*ic_cap+-2.37500e-07*ic_cap+3.62000e-05'
+ mcm5m2p1_ca_w_1_120_s_1_540 = '-3.90625e-07*ic_cap*ic_cap+-2.37500e-07*ic_cap+3.62000e-05'
+ mcm5m2p1_ca_w_1_120_s_3_500 = '-3.90625e-07*ic_cap*ic_cap+-2.37500e-07*ic_cap+3.62000e-05'
+ mcm5m2p1_cc_w_0_140_s_0_140 = '-9.12500e-13*ic_cap*ic_cap+-4.50000e-13*ic_cap+1.04000e-10'
+ mcm5m2p1_cc_w_0_140_s_0_175 = '-8.68750e-13*ic_cap*ic_cap+-6.50000e-13*ic_cap+1.02000e-10'
+ mcm5m2p1_cc_w_0_140_s_0_210 = '-7.53125e-13*ic_cap*ic_cap+-4.62500e-13*ic_cap+9.64000e-11'
+ mcm5m2p1_cc_w_0_140_s_0_280 = '-5.75000e-13*ic_cap*ic_cap+-3.50000e-13*ic_cap+8.54000e-11'
+ mcm5m2p1_cc_w_0_140_s_0_350 = '-4.00000e-13*ic_cap*ic_cap+-2.75000e-13*ic_cap+7.35000e-11'
+ mcm5m2p1_cc_w_0_140_s_0_420 = '-3.21875e-13*ic_cap*ic_cap+-2.37500e-13*ic_cap+6.42000e-11'
+ mcm5m2p1_cc_w_0_140_s_0_560 = '-1.81250e-13*ic_cap*ic_cap+-1.25000e-13*ic_cap+5.11000e-11'
+ mcm5m2p1_cc_w_0_140_s_0_840 = '-5.00000e-14*ic_cap*ic_cap+-5.00000e-14*ic_cap+3.60000e-11'
+ mcm5m2p1_cc_w_0_140_s_1_540 = '5.31250e-14*ic_cap*ic_cap+3.75000e-14*ic_cap+1.87000e-11'
+ mcm5m2p1_cc_w_0_140_s_3_500 = '6.15625e-14*ic_cap*ic_cap+4.37500e-14*ic_cap+4.31000e-12'
+ mcm5m2p1_cc_w_1_120_s_0_140 = '-7.50000e-13*ic_cap*ic_cap+-5.00000e-13*ic_cap+1.24000e-10'
+ mcm5m2p1_cc_w_1_120_s_0_175 = '-6.87500e-13*ic_cap*ic_cap+-2.50000e-13*ic_cap+1.20000e-10'
+ mcm5m2p1_cc_w_1_120_s_0_210 = '-5.93750e-13*ic_cap*ic_cap+-3.75000e-13*ic_cap+1.14000e-10'
+ mcm5m2p1_cc_w_1_120_s_0_280 = '-4.50000e-13*ic_cap*ic_cap+-3.75000e-13*ic_cap+1.00000e-10'
+ mcm5m2p1_cc_w_1_120_s_0_350 = '-3.31250e-13*ic_cap*ic_cap+-2.00000e-13*ic_cap+8.73000e-11'
+ mcm5m2p1_cc_w_1_120_s_0_420 = '-2.15625e-13*ic_cap*ic_cap+-1.37500e-13*ic_cap+7.65000e-11'
+ mcm5m2p1_cc_w_1_120_s_0_560 = '-7.18750e-14*ic_cap*ic_cap+-6.25000e-14*ic_cap+6.08000e-11'
+ mcm5m2p1_cc_w_1_120_s_0_840 = '3.43750e-14*ic_cap*ic_cap+3.75000e-14*ic_cap+4.29000e-11'
+ mcm5m2p1_cc_w_1_120_s_1_540 = '1.15625e-13*ic_cap*ic_cap+6.25000e-14*ic_cap+2.26000e-11'
+ mcm5m2p1_cc_w_1_120_s_3_500 = '9.00000e-14*ic_cap*ic_cap+6.25000e-14*ic_cap+5.47000e-12'
+ mcm5m2p1_cf_w_0_140_s_0_140 = '-3.12500e-15*ic_cap*ic_cap+-2.50000e-15*ic_cap+2.52000e-12'
+ mcm5m2p1_cf_w_0_140_s_0_175 = '-1.06250e-14*ic_cap*ic_cap+-7.50000e-15*ic_cap+3.15000e-12'
+ mcm5m2p1_cf_w_0_140_s_0_210 = '-1.56250e-14*ic_cap*ic_cap+-1.00000e-14*ic_cap+3.78000e-12'
+ mcm5m2p1_cf_w_0_140_s_0_280 = '-3.00000e-14*ic_cap*ic_cap+-2.00000e-14*ic_cap+5.02000e-12'
+ mcm5m2p1_cf_w_0_140_s_0_350 = '-4.34375e-14*ic_cap*ic_cap+-2.62500e-14*ic_cap+6.23000e-12'
+ mcm5m2p1_cf_w_0_140_s_0_420 = '-5.46875e-14*ic_cap*ic_cap+-3.62500e-14*ic_cap+7.45000e-12'
+ mcm5m2p1_cf_w_0_140_s_0_560 = '-7.87500e-14*ic_cap*ic_cap+-4.75000e-14*ic_cap+9.75000e-12'
+ mcm5m2p1_cf_w_0_140_s_0_840 = '-1.25000e-13*ic_cap*ic_cap+-7.50000e-14*ic_cap+1.40000e-11'
+ mcm5m2p1_cf_w_0_140_s_1_540 = '-2.00000e-13*ic_cap*ic_cap+-1.25000e-13*ic_cap+2.25000e-11'
+ mcm5m2p1_cf_w_0_140_s_3_500 = '-2.25000e-13*ic_cap*ic_cap+-1.50000e-13*ic_cap+3.34000e-11'
+ mcm5m2p1_cf_w_1_120_s_0_140 = '-5.00000e-15*ic_cap*ic_cap+-2.50000e-15*ic_cap+2.59000e-12'
+ mcm5m2p1_cf_w_1_120_s_0_175 = '-1.15625e-14*ic_cap*ic_cap+-8.75000e-15*ic_cap+3.22000e-12'
+ mcm5m2p1_cf_w_1_120_s_0_210 = '-1.90625e-14*ic_cap*ic_cap+-1.12500e-14*ic_cap+3.85000e-12'
+ mcm5m2p1_cf_w_1_120_s_0_280 = '-3.06250e-14*ic_cap*ic_cap+-2.00000e-14*ic_cap+5.07000e-12'
+ mcm5m2p1_cf_w_1_120_s_0_350 = '-4.31250e-14*ic_cap*ic_cap+-2.75000e-14*ic_cap+6.28000e-12'
+ mcm5m2p1_cf_w_1_120_s_0_420 = '-5.62500e-14*ic_cap*ic_cap+-3.50000e-14*ic_cap+7.49000e-12'
+ mcm5m2p1_cf_w_1_120_s_0_560 = '-8.06250e-14*ic_cap*ic_cap+-5.00000e-14*ic_cap+9.82000e-12'
+ mcm5m2p1_cf_w_1_120_s_0_840 = '-1.25000e-13*ic_cap*ic_cap+-7.50000e-14*ic_cap+1.42000e-11'
+ mcm5m2p1_cf_w_1_120_s_1_540 = '-1.96875e-13*ic_cap*ic_cap+-1.12500e-13*ic_cap+2.31000e-11'
+ mcm5m2p1_cf_w_1_120_s_3_500 = '-2.31250e-13*ic_cap*ic_cap+-1.50000e-13*ic_cap+3.58000e-11'
+ mcm5m3_ca_w_1_600_s_10_000 = '-1.75000e-07*ic_cap*ic_cap+-1.00000e-07*ic_cap+1.99000e-05'
+ mcm5m3_ca_w_1_600_s_12_000 = '-1.75000e-07*ic_cap*ic_cap+-1.00000e-07*ic_cap+1.99000e-05'
+ mcm5m3_ca_w_1_600_s_1_600 = '-1.75000e-07*ic_cap*ic_cap+-1.00000e-07*ic_cap+1.99000e-05'
+ mcm5m3_ca_w_1_600_s_1_700 = '-1.75000e-07*ic_cap*ic_cap+-1.00000e-07*ic_cap+1.99000e-05'
+ mcm5m3_ca_w_1_600_s_1_900 = '-1.75000e-07*ic_cap*ic_cap+-1.00000e-07*ic_cap+1.99000e-05'
+ mcm5m3_ca_w_1_600_s_2_000 = '-1.75000e-07*ic_cap*ic_cap+-1.00000e-07*ic_cap+1.99000e-05'
+ mcm5m3_ca_w_1_600_s_2_400 = '-1.75000e-07*ic_cap*ic_cap+-1.00000e-07*ic_cap+1.99000e-05'
+ mcm5m3_ca_w_1_600_s_2_800 = '-1.75000e-07*ic_cap*ic_cap+-1.00000e-07*ic_cap+1.99000e-05'
+ mcm5m3_ca_w_1_600_s_3_200 = '-1.75000e-07*ic_cap*ic_cap+-1.00000e-07*ic_cap+1.99000e-05'
+ mcm5m3_ca_w_1_600_s_4_800 = '-1.75000e-07*ic_cap*ic_cap+-1.00000e-07*ic_cap+1.99000e-05'
+ mcm5m3_ca_w_4_000_s_10_000 = '-1.75000e-07*ic_cap*ic_cap+-1.00000e-07*ic_cap+1.99000e-05'
+ mcm5m3_ca_w_4_000_s_12_000 = '-1.75000e-07*ic_cap*ic_cap+-1.00000e-07*ic_cap+1.99000e-05'
+ mcm5m3_ca_w_4_000_s_1_600 = '-1.75000e-07*ic_cap*ic_cap+-1.00000e-07*ic_cap+1.99000e-05'
+ mcm5m3_ca_w_4_000_s_1_700 = '-1.75000e-07*ic_cap*ic_cap+-1.00000e-07*ic_cap+1.99000e-05'
+ mcm5m3_ca_w_4_000_s_1_900 = '-1.75000e-07*ic_cap*ic_cap+-1.00000e-07*ic_cap+1.99000e-05'
+ mcm5m3_ca_w_4_000_s_2_000 = '-1.75000e-07*ic_cap*ic_cap+-1.00000e-07*ic_cap+1.99000e-05'
+ mcm5m3_ca_w_4_000_s_2_400 = '-1.75000e-07*ic_cap*ic_cap+-1.00000e-07*ic_cap+1.99000e-05'
+ mcm5m3_ca_w_4_000_s_2_800 = '-1.75000e-07*ic_cap*ic_cap+-1.00000e-07*ic_cap+1.99000e-05'
+ mcm5m3_ca_w_4_000_s_3_200 = '-1.75000e-07*ic_cap*ic_cap+-1.00000e-07*ic_cap+1.99000e-05'
+ mcm5m3_ca_w_4_000_s_4_800 = '-1.75000e-07*ic_cap*ic_cap+-1.00000e-07*ic_cap+1.99000e-05'
+ mcm5m3_cc_w_1_600_s_10_000 = '1.56250e-15*ic_cap*ic_cap+6.25000e-15*ic_cap+6.90000e-12'
+ mcm5m3_cc_w_1_600_s_12_000 = '1.56250e-15*ic_cap*ic_cap+-6.25000e-15*ic_cap+5.20000e-12'
+ mcm5m3_cc_w_1_600_s_1_600 = '-4.21875e-13*ic_cap*ic_cap+-2.87500e-13*ic_cap+6.33000e-11'
+ mcm5m3_cc_w_1_600_s_1_700 = '-3.78125e-13*ic_cap*ic_cap+-2.37500e-13*ic_cap+5.96000e-11'
+ mcm5m3_cc_w_1_600_s_1_900 = '-3.03125e-13*ic_cap*ic_cap+-2.12500e-13*ic_cap+5.33000e-11'
+ mcm5m3_cc_w_1_600_s_2_000 = '-2.68750e-13*ic_cap*ic_cap+-2.00000e-13*ic_cap+5.06000e-11'
+ mcm5m3_cc_w_1_600_s_2_400 = '-1.90625e-13*ic_cap*ic_cap+-1.37500e-13*ic_cap+4.21000e-11'
+ mcm5m3_cc_w_1_600_s_2_800 = '-1.31250e-13*ic_cap*ic_cap+-1.00000e-13*ic_cap+3.58000e-11'
+ mcm5m3_cc_w_1_600_s_3_200 = '-9.68750e-14*ic_cap*ic_cap+-8.75000e-14*ic_cap+3.11000e-11'
+ mcm5m3_cc_w_1_600_s_4_800 = '-3.12500e-14*ic_cap*ic_cap+-2.50000e-14*ic_cap+1.94000e-11'
+ mcm5m3_cc_w_4_000_s_10_000 = '6.25000e-15*ic_cap*ic_cap+9.15000e-12'
+ mcm5m3_cc_w_4_000_s_12_000 = '3.12500e-15*ic_cap*ic_cap+7.10000e-12'
+ mcm5m3_cc_w_4_000_s_1_600 = '-4.09375e-13*ic_cap*ic_cap+-2.87500e-13*ic_cap+6.86000e-11'
+ mcm5m3_cc_w_4_000_s_1_700 = '-3.59375e-13*ic_cap*ic_cap+-2.37500e-13*ic_cap+6.48000e-11'
+ mcm5m3_cc_w_4_000_s_1_900 = '-2.90625e-13*ic_cap*ic_cap+-1.87500e-13*ic_cap+5.83000e-11'
+ mcm5m3_cc_w_4_000_s_2_000 = '-2.56250e-13*ic_cap*ic_cap+-1.75000e-13*ic_cap+5.55000e-11'
+ mcm5m3_cc_w_4_000_s_2_400 = '-1.75000e-13*ic_cap*ic_cap+-1.25000e-13*ic_cap+4.66000e-11'
+ mcm5m3_cc_w_4_000_s_2_800 = '-1.21875e-13*ic_cap*ic_cap+-8.75000e-14*ic_cap+4.01000e-11'
+ mcm5m3_cc_w_4_000_s_3_200 = '-9.06250e-14*ic_cap*ic_cap+-6.25000e-14*ic_cap+3.52000e-11'
+ mcm5m3_cc_w_4_000_s_4_800 = '-3.12500e-14*ic_cap*ic_cap+-2.50000e-14*ic_cap+2.30000e-11'
+ mcm5m3_cf_w_1_600_s_10_000 = '-2.31250e-13*ic_cap*ic_cap+-1.50000e-13*ic_cap+4.24000e-11'
+ mcm5m3_cf_w_1_600_s_12_000 = '-2.37500e-13*ic_cap*ic_cap+-1.50000e-13*ic_cap+4.41000e-11'
+ mcm5m3_cf_w_1_600_s_1_600 = '-7.50000e-14*ic_cap*ic_cap+-5.00000e-14*ic_cap+1.42000e-11'
+ mcm5m3_cf_w_1_600_s_1_700 = '-8.12500e-14*ic_cap*ic_cap+-5.00000e-14*ic_cap+1.50000e-11'
+ mcm5m3_cf_w_1_600_s_1_900 = '-9.37500e-14*ic_cap*ic_cap+-5.00000e-14*ic_cap+1.65000e-11'
+ mcm5m3_cf_w_1_600_s_2_000 = '-1.00000e-13*ic_cap*ic_cap+-5.00000e-14*ic_cap+1.72000e-11'
+ mcm5m3_cf_w_1_600_s_2_400 = '-1.25000e-13*ic_cap*ic_cap+-7.50000e-14*ic_cap+2.00000e-11'
+ mcm5m3_cf_w_1_600_s_2_800 = '-1.40625e-13*ic_cap*ic_cap+-8.75000e-14*ic_cap+2.25000e-11'
+ mcm5m3_cf_w_1_600_s_3_200 = '-1.59375e-13*ic_cap*ic_cap+-8.75000e-14*ic_cap+2.48000e-11'
+ mcm5m3_cf_w_1_600_s_4_800 = '-2.00000e-13*ic_cap*ic_cap+-1.25000e-13*ic_cap+3.19000e-11'
+ mcm5m3_cf_w_4_000_s_10_000 = '-2.31250e-13*ic_cap*ic_cap+-1.50000e-13*ic_cap+4.33000e-11'
+ mcm5m3_cf_w_4_000_s_12_000 = '-2.37500e-13*ic_cap*ic_cap+-1.50000e-13*ic_cap+4.53000e-11'
+ mcm5m3_cf_w_4_000_s_1_600 = '-7.50000e-14*ic_cap*ic_cap+-5.00000e-14*ic_cap+1.42000e-11'
+ mcm5m3_cf_w_4_000_s_1_700 = '-8.12500e-14*ic_cap*ic_cap+-5.00000e-14*ic_cap+1.50000e-11'
+ mcm5m3_cf_w_4_000_s_1_900 = '-9.37500e-14*ic_cap*ic_cap+-5.00000e-14*ic_cap+1.65000e-11'
+ mcm5m3_cf_w_4_000_s_2_000 = '-1.00000e-13*ic_cap*ic_cap+-5.00000e-14*ic_cap+1.72000e-11'
+ mcm5m3_cf_w_4_000_s_2_400 = '-1.25000e-13*ic_cap*ic_cap+-7.50000e-14*ic_cap+2.00000e-11'
+ mcm5m3_cf_w_4_000_s_2_800 = '-1.40625e-13*ic_cap*ic_cap+-8.75000e-14*ic_cap+2.25000e-11'
+ mcm5m3_cf_w_4_000_s_3_200 = '-1.56250e-13*ic_cap*ic_cap+-1.00000e-13*ic_cap+2.48000e-11'
+ mcm5m3_cf_w_4_000_s_4_800 = '-2.00000e-13*ic_cap*ic_cap+-1.25000e-13*ic_cap+3.21000e-11'
+ mcm5m3d_ca_w_0_300_s_0_300 = '-3.09375e-07*ic_cap*ic_cap+-1.87500e-07*ic_cap+3.40000e-05'
+ mcm5m3d_ca_w_0_300_s_0_360 = '-3.09375e-07*ic_cap*ic_cap+-1.87500e-07*ic_cap+3.40000e-05'
+ mcm5m3d_ca_w_0_300_s_0_450 = '-3.09375e-07*ic_cap*ic_cap+-1.87500e-07*ic_cap+3.40000e-05'
+ mcm5m3d_ca_w_0_300_s_0_600 = '-3.09375e-07*ic_cap*ic_cap+-1.87500e-07*ic_cap+3.40000e-05'
+ mcm5m3d_ca_w_0_300_s_0_800 = '-3.09375e-07*ic_cap*ic_cap+-1.87500e-07*ic_cap+3.40000e-05'
+ mcm5m3d_ca_w_0_300_s_1_000 = '-3.09375e-07*ic_cap*ic_cap+-1.87500e-07*ic_cap+3.40000e-05'
+ mcm5m3d_ca_w_0_300_s_1_200 = '-3.09375e-07*ic_cap*ic_cap+-1.87500e-07*ic_cap+3.40000e-05'
+ mcm5m3d_ca_w_0_300_s_2_100 = '-3.09375e-07*ic_cap*ic_cap+-1.87500e-07*ic_cap+3.40000e-05'
+ mcm5m3d_ca_w_0_300_s_3_300 = '-3.09375e-07*ic_cap*ic_cap+-1.87500e-07*ic_cap+3.40000e-05'
+ mcm5m3d_ca_w_0_300_s_9_000 = '-3.09375e-07*ic_cap*ic_cap+-1.87500e-07*ic_cap+3.40000e-05'
+ mcm5m3d_ca_w_2_400_s_0_300 = '-3.09375e-07*ic_cap*ic_cap+-1.87500e-07*ic_cap+3.40000e-05'
+ mcm5m3d_ca_w_2_400_s_0_360 = '-3.09375e-07*ic_cap*ic_cap+-1.87500e-07*ic_cap+3.40000e-05'
+ mcm5m3d_ca_w_2_400_s_0_450 = '-3.09375e-07*ic_cap*ic_cap+-1.87500e-07*ic_cap+3.40000e-05'
+ mcm5m3d_ca_w_2_400_s_0_600 = '-3.09375e-07*ic_cap*ic_cap+-1.87500e-07*ic_cap+3.40000e-05'
+ mcm5m3d_ca_w_2_400_s_0_800 = '-3.09375e-07*ic_cap*ic_cap+-1.87500e-07*ic_cap+3.40000e-05'
+ mcm5m3d_ca_w_2_400_s_1_000 = '-3.09375e-07*ic_cap*ic_cap+-1.87500e-07*ic_cap+3.40000e-05'
+ mcm5m3d_ca_w_2_400_s_1_200 = '-3.09375e-07*ic_cap*ic_cap+-1.87500e-07*ic_cap+3.40000e-05'
+ mcm5m3d_ca_w_2_400_s_2_100 = '-3.09375e-07*ic_cap*ic_cap+-1.87500e-07*ic_cap+3.40000e-05'
+ mcm5m3d_ca_w_2_400_s_3_300 = '-3.09375e-07*ic_cap*ic_cap+-1.87500e-07*ic_cap+3.40000e-05'
+ mcm5m3d_ca_w_2_400_s_9_000 = '-3.09375e-07*ic_cap*ic_cap+-1.87500e-07*ic_cap+3.40000e-05'
+ mcm5m3d_cc_w_0_300_s_0_300 = '-7.43750e-13*ic_cap*ic_cap+-4.25000e-13*ic_cap+1.01000e-10'
+ mcm5m3d_cc_w_0_300_s_0_360 = '-6.62500e-13*ic_cap*ic_cap+-3.75000e-13*ic_cap+9.37000e-11'
+ mcm5m3d_cc_w_0_300_s_0_450 = '-5.62500e-13*ic_cap*ic_cap+-3.00000e-13*ic_cap+8.39000e-11'
+ mcm5m3d_cc_w_0_300_s_0_600 = '-4.03125e-13*ic_cap*ic_cap+-2.37500e-13*ic_cap+7.03000e-11'
+ mcm5m3d_cc_w_0_300_s_0_800 = '-2.34375e-13*ic_cap*ic_cap+-1.62500e-13*ic_cap+5.64000e-11'
+ mcm5m3d_cc_w_0_300_s_1_000 = '-1.62500e-13*ic_cap*ic_cap+-1.25000e-13*ic_cap+4.64000e-11'
+ mcm5m3d_cc_w_0_300_s_1_200 = '-8.75000e-14*ic_cap*ic_cap+-7.50000e-14*ic_cap+3.85000e-11'
+ mcm5m3d_cc_w_0_300_s_2_100 = '2.18750e-14*ic_cap*ic_cap+1.25000e-14*ic_cap+1.94000e-11'
+ mcm5m3d_cc_w_0_300_s_3_300 = '5.46875e-14*ic_cap*ic_cap+3.37500e-14*ic_cap+8.69000e-12'
+ mcm5m3d_cc_w_0_300_s_9_000 = '9.06250e-15*ic_cap*ic_cap+7.50000e-15*ic_cap+2.80000e-13'
+ mcm5m3d_cc_w_2_400_s_0_300 = '-5.93750e-13*ic_cap*ic_cap+-3.75000e-13*ic_cap+1.13000e-10'
+ mcm5m3d_cc_w_2_400_s_0_360 = '-5.37500e-13*ic_cap*ic_cap+-3.25000e-13*ic_cap+1.05000e-10'
+ mcm5m3d_cc_w_2_400_s_0_450 = '-3.96875e-13*ic_cap*ic_cap+-2.37500e-13*ic_cap+9.32000e-11'
+ mcm5m3d_cc_w_2_400_s_0_600 = '-2.65625e-13*ic_cap*ic_cap+-1.62500e-13*ic_cap+7.81000e-11'
+ mcm5m3d_cc_w_2_400_s_0_800 = '-1.34375e-13*ic_cap*ic_cap+-8.75000e-14*ic_cap+6.28000e-11'
+ mcm5m3d_cc_w_2_400_s_1_000 = '-5.93750e-14*ic_cap*ic_cap+-3.75000e-14*ic_cap+5.15000e-11'
+ mcm5m3d_cc_w_2_400_s_1_200 = '-1.25000e-14*ic_cap*ic_cap+4.30000e-11'
+ mcm5m3d_cc_w_2_400_s_2_100 = '8.12500e-14*ic_cap*ic_cap+5.00000e-14*ic_cap+2.18000e-11'
+ mcm5m3d_cc_w_2_400_s_3_300 = '9.31250e-14*ic_cap*ic_cap+6.25000e-14*ic_cap+9.86000e-12'
+ mcm5m3d_cc_w_2_400_s_9_000 = '1.15625e-14*ic_cap*ic_cap+1.37500e-14*ic_cap+3.20000e-13'
+ mcm5m3d_cf_w_0_300_s_0_300 = '-1.03125e-14*ic_cap*ic_cap+-6.25000e-15*ic_cap+4.94000e-12'
+ mcm5m3d_cf_w_0_300_s_0_360 = '-1.84375e-14*ic_cap*ic_cap+-1.12500e-14*ic_cap+5.91000e-12'
+ mcm5m3d_cf_w_0_300_s_0_450 = '-3.12500e-14*ic_cap*ic_cap+-1.75000e-14*ic_cap+7.38000e-12'
+ mcm5m3d_cf_w_0_300_s_0_600 = '-5.06250e-14*ic_cap*ic_cap+-3.00000e-14*ic_cap+9.72000e-12'
+ mcm5m3d_cf_w_0_300_s_0_800 = '-7.50000e-14*ic_cap*ic_cap+-5.00000e-14*ic_cap+1.26000e-11'
+ mcm5m3d_cf_w_0_300_s_1_000 = '-1.03125e-13*ic_cap*ic_cap+-6.25000e-14*ic_cap+1.54000e-11'
+ mcm5m3d_cf_w_0_300_s_1_200 = '-1.25000e-13*ic_cap*ic_cap+-7.50000e-14*ic_cap+1.81000e-11'
+ mcm5m3d_cf_w_0_300_s_2_100 = '-1.93750e-13*ic_cap*ic_cap+-1.25000e-13*ic_cap+2.77000e-11'
+ mcm5m3d_cf_w_0_300_s_3_300 = '-2.37500e-13*ic_cap*ic_cap+-1.50000e-13*ic_cap+3.55000e-11'
+ mcm5m3d_cf_w_0_300_s_9_000 = '-2.03125e-13*ic_cap*ic_cap+-1.37500e-13*ic_cap+4.31000e-11'
+ mcm5m3d_cf_w_2_400_s_0_300 = '-1.03125e-14*ic_cap*ic_cap+-6.25000e-15*ic_cap+4.99000e-12'
+ mcm5m3d_cf_w_2_400_s_0_360 = '-1.87500e-14*ic_cap*ic_cap+-1.00000e-14*ic_cap+5.96000e-12'
+ mcm5m3d_cf_w_2_400_s_0_450 = '-3.12500e-14*ic_cap*ic_cap+-2.00000e-14*ic_cap+7.39000e-12'
+ mcm5m3d_cf_w_2_400_s_0_600 = '-5.25000e-14*ic_cap*ic_cap+-3.25000e-14*ic_cap+9.73000e-12'
+ mcm5m3d_cf_w_2_400_s_0_800 = '-7.50000e-14*ic_cap*ic_cap+-5.00000e-14*ic_cap+1.27000e-11'
+ mcm5m3d_cf_w_2_400_s_1_000 = '-1.03125e-13*ic_cap*ic_cap+-6.25000e-14*ic_cap+1.56000e-11'
+ mcm5m3d_cf_w_2_400_s_1_200 = '-1.25000e-13*ic_cap*ic_cap+-7.50000e-14*ic_cap+1.83000e-11'
+ mcm5m3d_cf_w_2_400_s_2_100 = '-1.93750e-13*ic_cap*ic_cap+-1.25000e-13*ic_cap+2.83000e-11'
+ mcm5m3d_cf_w_2_400_s_3_300 = '-2.31250e-13*ic_cap*ic_cap+-1.50000e-13*ic_cap+3.69000e-11'
+ mcm5m3d_cf_w_2_400_s_9_000 = '-1.71875e-13*ic_cap*ic_cap+-1.12500e-13*ic_cap+4.56000e-11'
+ mcm5m3f_ca_w_0_300_s_0_300 = '-3.00000e-07*ic_cap*ic_cap+-1.75000e-07*ic_cap+3.24000e-05'
+ mcm5m3f_ca_w_0_300_s_0_360 = '-3.00000e-07*ic_cap*ic_cap+-1.75000e-07*ic_cap+3.24000e-05'
+ mcm5m3f_ca_w_0_300_s_0_450 = '-3.00000e-07*ic_cap*ic_cap+-1.75000e-07*ic_cap+3.24000e-05'
+ mcm5m3f_ca_w_0_300_s_0_600 = '-3.00000e-07*ic_cap*ic_cap+-1.75000e-07*ic_cap+3.24000e-05'
+ mcm5m3f_ca_w_0_300_s_0_800 = '-3.00000e-07*ic_cap*ic_cap+-1.75000e-07*ic_cap+3.24000e-05'
+ mcm5m3f_ca_w_0_300_s_1_000 = '-3.00000e-07*ic_cap*ic_cap+-1.75000e-07*ic_cap+3.24000e-05'
+ mcm5m3f_ca_w_0_300_s_1_200 = '-3.00000e-07*ic_cap*ic_cap+-1.75000e-07*ic_cap+3.24000e-05'
+ mcm5m3f_ca_w_0_300_s_2_100 = '-3.00000e-07*ic_cap*ic_cap+-1.75000e-07*ic_cap+3.24000e-05'
+ mcm5m3f_ca_w_0_300_s_3_300 = '-3.00000e-07*ic_cap*ic_cap+-1.75000e-07*ic_cap+3.24000e-05'
+ mcm5m3f_ca_w_0_300_s_9_000 = '-3.00000e-07*ic_cap*ic_cap+-1.75000e-07*ic_cap+3.24000e-05'
+ mcm5m3f_ca_w_2_400_s_0_300 = '-3.00000e-07*ic_cap*ic_cap+-1.75000e-07*ic_cap+3.24000e-05'
+ mcm5m3f_ca_w_2_400_s_0_360 = '-3.00000e-07*ic_cap*ic_cap+-1.75000e-07*ic_cap+3.24000e-05'
+ mcm5m3f_ca_w_2_400_s_0_450 = '-3.00000e-07*ic_cap*ic_cap+-1.75000e-07*ic_cap+3.24000e-05'
+ mcm5m3f_ca_w_2_400_s_0_600 = '-3.00000e-07*ic_cap*ic_cap+-1.75000e-07*ic_cap+3.24000e-05'
+ mcm5m3f_ca_w_2_400_s_0_800 = '-3.00000e-07*ic_cap*ic_cap+-1.75000e-07*ic_cap+3.24000e-05'
+ mcm5m3f_ca_w_2_400_s_1_000 = '-3.00000e-07*ic_cap*ic_cap+-1.75000e-07*ic_cap+3.24000e-05'
+ mcm5m3f_ca_w_2_400_s_1_200 = '-3.00000e-07*ic_cap*ic_cap+-1.75000e-07*ic_cap+3.24000e-05'
+ mcm5m3f_ca_w_2_400_s_2_100 = '-3.00000e-07*ic_cap*ic_cap+-1.75000e-07*ic_cap+3.24000e-05'
+ mcm5m3f_ca_w_2_400_s_3_300 = '-3.00000e-07*ic_cap*ic_cap+-1.75000e-07*ic_cap+3.24000e-05'
+ mcm5m3f_ca_w_2_400_s_9_000 = '-3.00000e-07*ic_cap*ic_cap+-1.75000e-07*ic_cap+3.24000e-05'
+ mcm5m3f_cc_w_0_300_s_0_300 = '-7.81250e-13*ic_cap*ic_cap+-4.25000e-13*ic_cap+1.02000e-10'
+ mcm5m3f_cc_w_0_300_s_0_360 = '-6.65625e-13*ic_cap*ic_cap+-3.87500e-13*ic_cap+9.41000e-11'
+ mcm5m3f_cc_w_0_300_s_0_450 = '-5.65625e-13*ic_cap*ic_cap+-3.12500e-13*ic_cap+8.44000e-11'
+ mcm5m3f_cc_w_0_300_s_0_600 = '-4.03125e-13*ic_cap*ic_cap+-2.37500e-13*ic_cap+7.08000e-11'
+ mcm5m3f_cc_w_0_300_s_0_800 = '-2.40625e-13*ic_cap*ic_cap+-1.62500e-13*ic_cap+5.71000e-11'
+ mcm5m3f_cc_w_0_300_s_1_000 = '-1.53125e-13*ic_cap*ic_cap+-1.37500e-13*ic_cap+4.70000e-11'
+ mcm5m3f_cc_w_0_300_s_1_200 = '-9.06250e-14*ic_cap*ic_cap+-6.25000e-14*ic_cap+3.92000e-11'
+ mcm5m3f_cc_w_0_300_s_2_100 = '2.18750e-14*ic_cap*ic_cap+1.25000e-14*ic_cap+2.02000e-11'
+ mcm5m3f_cc_w_0_300_s_3_300 = '5.68750e-14*ic_cap*ic_cap+3.75000e-14*ic_cap+9.34000e-12'
+ mcm5m3f_cc_w_0_300_s_9_000 = '1.20312e-14*ic_cap*ic_cap+9.37500e-15*ic_cap+3.50000e-13'
+ mcm5m3f_cc_w_2_400_s_0_300 = '-5.93750e-13*ic_cap*ic_cap+-3.75000e-13*ic_cap+1.14000e-10'
+ mcm5m3f_cc_w_2_400_s_0_360 = '-5.28125e-13*ic_cap*ic_cap+-3.12500e-13*ic_cap+1.06000e-10'
+ mcm5m3f_cc_w_2_400_s_0_450 = '-3.90625e-13*ic_cap*ic_cap+-2.37500e-13*ic_cap+9.43000e-11'
+ mcm5m3f_cc_w_2_400_s_0_600 = '-2.65625e-13*ic_cap*ic_cap+-1.62500e-13*ic_cap+7.93000e-11'
+ mcm5m3f_cc_w_2_400_s_0_800 = '-1.31250e-13*ic_cap*ic_cap+-7.50000e-14*ic_cap+6.40000e-11'
+ mcm5m3f_cc_w_2_400_s_1_000 = '-5.62500e-14*ic_cap*ic_cap+-5.00000e-14*ic_cap+5.27000e-11'
+ mcm5m3f_cc_w_2_400_s_1_200 = '-9.37500e-15*ic_cap*ic_cap+-1.25000e-14*ic_cap+4.42000e-11'
+ mcm5m3f_cc_w_2_400_s_2_100 = '8.75000e-14*ic_cap*ic_cap+5.00000e-14*ic_cap+2.29000e-11'
+ mcm5m3f_cc_w_2_400_s_3_300 = '9.68750e-14*ic_cap*ic_cap+6.25000e-14*ic_cap+1.08000e-11'
+ mcm5m3f_cc_w_2_400_s_9_000 = '1.53125e-14*ic_cap*ic_cap+1.75000e-14*ic_cap+4.15000e-13'
+ mcm5m3f_cf_w_0_300_s_0_300 = '-1.03125e-14*ic_cap*ic_cap+-6.25000e-15*ic_cap+4.70000e-12'
+ mcm5m3f_cf_w_0_300_s_0_360 = '-1.90625e-14*ic_cap*ic_cap+-1.12500e-14*ic_cap+5.63000e-12'
+ mcm5m3f_cf_w_0_300_s_0_450 = '-3.06250e-14*ic_cap*ic_cap+-1.75000e-14*ic_cap+7.03000e-12'
+ mcm5m3f_cf_w_0_300_s_0_600 = '-5.03125e-14*ic_cap*ic_cap+-2.87500e-14*ic_cap+9.28000e-12'
+ mcm5m3f_cf_w_0_300_s_0_800 = '-7.50000e-14*ic_cap*ic_cap+-5.00000e-14*ic_cap+1.20000e-11'
+ mcm5m3f_cf_w_0_300_s_1_000 = '-9.68750e-14*ic_cap*ic_cap+-6.25000e-14*ic_cap+1.47000e-11'
+ mcm5m3f_cf_w_0_300_s_1_200 = '-1.25000e-13*ic_cap*ic_cap+-7.50000e-14*ic_cap+1.73000e-11'
+ mcm5m3f_cf_w_0_300_s_2_100 = '-1.90625e-13*ic_cap*ic_cap+-1.12500e-13*ic_cap+2.66000e-11'
+ mcm5m3f_cf_w_0_300_s_3_300 = '-2.31250e-13*ic_cap*ic_cap+-1.50000e-13*ic_cap+3.43000e-11'
+ mcm5m3f_cf_w_0_300_s_9_000 = '-2.00000e-13*ic_cap*ic_cap+-1.25000e-13*ic_cap+4.24000e-11'
+ mcm5m3f_cf_w_2_400_s_0_300 = '-1.06250e-14*ic_cap*ic_cap+-7.50000e-15*ic_cap+4.75000e-12'
+ mcm5m3f_cf_w_2_400_s_0_360 = '-1.84375e-14*ic_cap*ic_cap+-1.12500e-14*ic_cap+5.67000e-12'
+ mcm5m3f_cf_w_2_400_s_0_450 = '-3.06250e-14*ic_cap*ic_cap+-1.75000e-14*ic_cap+7.03000e-12'
+ mcm5m3f_cf_w_2_400_s_0_600 = '-5.15625e-14*ic_cap*ic_cap+-3.12500e-14*ic_cap+9.27000e-12'
+ mcm5m3f_cf_w_2_400_s_0_800 = '-7.50000e-14*ic_cap*ic_cap+-5.00000e-14*ic_cap+1.21000e-11'
+ mcm5m3f_cf_w_2_400_s_1_000 = '-1.03125e-13*ic_cap*ic_cap+-6.25000e-14*ic_cap+1.49000e-11'
+ mcm5m3f_cf_w_2_400_s_1_200 = '-1.25000e-13*ic_cap*ic_cap+-7.50000e-14*ic_cap+1.75000e-11'
+ mcm5m3f_cf_w_2_400_s_2_100 = '-1.93750e-13*ic_cap*ic_cap+-1.25000e-13*ic_cap+2.72000e-11'
+ mcm5m3f_cf_w_2_400_s_3_300 = '-2.21875e-13*ic_cap*ic_cap+-1.37500e-13*ic_cap+3.56000e-11'
+ mcm5m3f_cf_w_2_400_s_9_000 = '-1.65625e-13*ic_cap*ic_cap+-1.12500e-13*ic_cap+4.50000e-11'
+ mcm5m3l1_ca_w_0_300_s_0_300 = '-3.81250e-07*ic_cap*ic_cap+-2.25000e-07*ic_cap+4.00000e-05'
+ mcm5m3l1_ca_w_0_300_s_0_360 = '-3.81250e-07*ic_cap*ic_cap+-2.25000e-07*ic_cap+4.00000e-05'
+ mcm5m3l1_ca_w_0_300_s_0_450 = '-3.81250e-07*ic_cap*ic_cap+-2.25000e-07*ic_cap+4.00000e-05'
+ mcm5m3l1_ca_w_0_300_s_0_600 = '-3.81250e-07*ic_cap*ic_cap+-2.25000e-07*ic_cap+4.00000e-05'
+ mcm5m3l1_ca_w_0_300_s_0_800 = '-3.81250e-07*ic_cap*ic_cap+-2.25000e-07*ic_cap+4.00000e-05'
+ mcm5m3l1_ca_w_0_300_s_1_000 = '-3.81250e-07*ic_cap*ic_cap+-2.25000e-07*ic_cap+4.00000e-05'
+ mcm5m3l1_ca_w_0_300_s_1_200 = '-3.81250e-07*ic_cap*ic_cap+-2.25000e-07*ic_cap+4.00000e-05'
+ mcm5m3l1_ca_w_0_300_s_2_100 = '-3.81250e-07*ic_cap*ic_cap+-2.25000e-07*ic_cap+4.00000e-05'
+ mcm5m3l1_ca_w_0_300_s_3_300 = '-3.81250e-07*ic_cap*ic_cap+-2.25000e-07*ic_cap+4.00000e-05'
+ mcm5m3l1_ca_w_0_300_s_9_000 = '-3.81250e-07*ic_cap*ic_cap+-2.25000e-07*ic_cap+4.00000e-05'
+ mcm5m3l1_ca_w_2_400_s_0_300 = '-3.81250e-07*ic_cap*ic_cap+-2.25000e-07*ic_cap+4.00000e-05'
+ mcm5m3l1_ca_w_2_400_s_0_360 = '-3.81250e-07*ic_cap*ic_cap+-2.25000e-07*ic_cap+4.00000e-05'
+ mcm5m3l1_ca_w_2_400_s_0_450 = '-3.81250e-07*ic_cap*ic_cap+-2.25000e-07*ic_cap+4.00000e-05'
+ mcm5m3l1_ca_w_2_400_s_0_600 = '-3.81250e-07*ic_cap*ic_cap+-2.25000e-07*ic_cap+4.00000e-05'
+ mcm5m3l1_ca_w_2_400_s_0_800 = '-3.81250e-07*ic_cap*ic_cap+-2.25000e-07*ic_cap+4.00000e-05'
+ mcm5m3l1_ca_w_2_400_s_1_000 = '-3.81250e-07*ic_cap*ic_cap+-2.25000e-07*ic_cap+4.00000e-05'
+ mcm5m3l1_ca_w_2_400_s_1_200 = '-3.81250e-07*ic_cap*ic_cap+-2.25000e-07*ic_cap+4.00000e-05'
+ mcm5m3l1_ca_w_2_400_s_2_100 = '-3.81250e-07*ic_cap*ic_cap+-2.25000e-07*ic_cap+4.00000e-05'
+ mcm5m3l1_ca_w_2_400_s_3_300 = '-3.81250e-07*ic_cap*ic_cap+-2.25000e-07*ic_cap+4.00000e-05'
+ mcm5m3l1_ca_w_2_400_s_9_000 = '-3.81250e-07*ic_cap*ic_cap+-2.25000e-07*ic_cap+4.00000e-05'
+ mcm5m3l1_cc_w_0_300_s_0_300 = '-7.31250e-13*ic_cap*ic_cap+-4.25000e-13*ic_cap+9.96000e-11'
+ mcm5m3l1_cc_w_0_300_s_0_360 = '-6.56250e-13*ic_cap*ic_cap+-3.75000e-13*ic_cap+9.23000e-11'
+ mcm5m3l1_cc_w_0_300_s_0_450 = '-5.28125e-13*ic_cap*ic_cap+-3.37500e-13*ic_cap+8.21000e-11'
+ mcm5m3l1_cc_w_0_300_s_0_600 = '-3.81250e-13*ic_cap*ic_cap+-2.25000e-13*ic_cap+6.83000e-11'
+ mcm5m3l1_cc_w_0_300_s_0_800 = '-2.15625e-13*ic_cap*ic_cap+-1.37500e-13*ic_cap+5.42000e-11'
+ mcm5m3l1_cc_w_0_300_s_1_000 = '-1.40625e-13*ic_cap*ic_cap+-8.75000e-14*ic_cap+4.40000e-11'
+ mcm5m3l1_cc_w_0_300_s_1_200 = '-7.50000e-14*ic_cap*ic_cap+-5.00000e-14*ic_cap+3.61000e-11'
+ mcm5m3l1_cc_w_0_300_s_2_100 = '4.06250e-14*ic_cap*ic_cap+1.25000e-14*ic_cap+1.68000e-11'
+ mcm5m3l1_cc_w_0_300_s_3_300 = '5.84375e-14*ic_cap*ic_cap+3.62500e-14*ic_cap+6.77000e-12'
+ mcm5m3l1_cc_w_0_300_s_9_000 = '4.53125e-15*ic_cap*ic_cap+4.37500e-15*ic_cap+1.55000e-13'
+ mcm5m3l1_cc_w_2_400_s_0_300 = '-5.96875e-13*ic_cap*ic_cap+-3.87500e-13*ic_cap+1.10000e-10'
+ mcm5m3l1_cc_w_2_400_s_0_360 = '-5.00000e-13*ic_cap*ic_cap+-3.00000e-13*ic_cap+1.01000e-10'
+ mcm5m3l1_cc_w_2_400_s_0_450 = '-3.71875e-13*ic_cap*ic_cap+-2.12500e-13*ic_cap+8.94000e-11'
+ mcm5m3l1_cc_w_2_400_s_0_600 = '-2.46875e-13*ic_cap*ic_cap+-1.37500e-13*ic_cap+7.43000e-11'
+ mcm5m3l1_cc_w_2_400_s_0_800 = '-1.18750e-13*ic_cap*ic_cap+-7.50000e-14*ic_cap+5.91000e-11'
+ mcm5m3l1_cc_w_2_400_s_1_000 = '-5.31250e-14*ic_cap*ic_cap+-3.75000e-14*ic_cap+4.79000e-11'
+ mcm5m3l1_cc_w_2_400_s_1_200 = '6.25000e-15*ic_cap*ic_cap+3.93000e-11'
+ mcm5m3l1_cc_w_2_400_s_2_100 = '8.12500e-14*ic_cap*ic_cap+5.00000e-14*ic_cap+1.86000e-11'
+ mcm5m3l1_cc_w_2_400_s_3_300 = '8.46875e-14*ic_cap*ic_cap+5.62500e-14*ic_cap+7.52000e-12'
+ mcm5m3l1_cc_w_2_400_s_9_000 = '6.56250e-15*ic_cap*ic_cap+5.00000e-15*ic_cap+1.65000e-13'
+ mcm5m3l1_cf_w_0_300_s_0_300 = '-1.46875e-14*ic_cap*ic_cap+-8.75000e-15*ic_cap+5.80000e-12'
+ mcm5m3l1_cf_w_0_300_s_0_360 = '-2.40625e-14*ic_cap*ic_cap+-1.62500e-14*ic_cap+6.92000e-12'
+ mcm5m3l1_cf_w_0_300_s_0_450 = '-3.96875e-14*ic_cap*ic_cap+-2.37500e-14*ic_cap+8.63000e-12'
+ mcm5m3l1_cf_w_0_300_s_0_600 = '-5.93750e-14*ic_cap*ic_cap+-3.75000e-14*ic_cap+1.13000e-11'
+ mcm5m3l1_cf_w_0_300_s_0_800 = '-9.68750e-14*ic_cap*ic_cap+-6.25000e-14*ic_cap+1.47000e-11'
+ mcm5m3l1_cf_w_0_300_s_1_000 = '-1.25000e-13*ic_cap*ic_cap+-7.50000e-14*ic_cap+1.79000e-11'
+ mcm5m3l1_cf_w_0_300_s_1_200 = '-1.53125e-13*ic_cap*ic_cap+-8.75000e-14*ic_cap+2.09000e-11'
+ mcm5m3l1_cf_w_0_300_s_2_100 = '-2.28125e-13*ic_cap*ic_cap+-1.37500e-13*ic_cap+3.14000e-11'
+ mcm5m3l1_cf_w_0_300_s_3_300 = '-2.59375e-13*ic_cap*ic_cap+-1.62500e-13*ic_cap+3.92000e-11'
+ mcm5m3l1_cf_w_0_300_s_9_000 = '-2.15625e-13*ic_cap*ic_cap+-1.37500e-13*ic_cap+4.54000e-11'
+ mcm5m3l1_cf_w_2_400_s_0_300 = '-1.37500e-14*ic_cap*ic_cap+-1.00000e-14*ic_cap+5.84000e-12'
+ mcm5m3l1_cf_w_2_400_s_0_360 = '-2.40625e-14*ic_cap*ic_cap+-1.37500e-14*ic_cap+6.97000e-12'
+ mcm5m3l1_cf_w_2_400_s_0_450 = '-4.00000e-14*ic_cap*ic_cap+-2.50000e-14*ic_cap+8.65000e-12'
+ mcm5m3l1_cf_w_2_400_s_0_600 = '-5.93750e-14*ic_cap*ic_cap+-3.75000e-14*ic_cap+1.13000e-11'
+ mcm5m3l1_cf_w_2_400_s_0_800 = '-9.68750e-14*ic_cap*ic_cap+-6.25000e-14*ic_cap+1.48000e-11'
+ mcm5m3l1_cf_w_2_400_s_1_000 = '-1.31250e-13*ic_cap*ic_cap+-7.50000e-14*ic_cap+1.82000e-11'
+ mcm5m3l1_cf_w_2_400_s_1_200 = '-1.50000e-13*ic_cap*ic_cap+-1.00000e-13*ic_cap+2.12000e-11'
+ mcm5m3l1_cf_w_2_400_s_2_100 = '-2.25000e-13*ic_cap*ic_cap+-1.50000e-13*ic_cap+3.21000e-11'
+ mcm5m3l1_cf_w_2_400_s_3_300 = '-2.53125e-13*ic_cap*ic_cap+-1.62500e-13*ic_cap+4.06000e-11'
+ mcm5m3l1_cf_w_2_400_s_9_000 = '-1.81250e-13*ic_cap*ic_cap+-1.25000e-13*ic_cap+4.74000e-11'
+ mcm5m3m1_ca_w_0_300_s_0_300 = '-5.62500e-07*ic_cap*ic_cap+-3.25000e-07*ic_cap+5.27000e-05'
+ mcm5m3m1_ca_w_0_300_s_0_360 = '-5.62500e-07*ic_cap*ic_cap+-3.25000e-07*ic_cap+5.27000e-05'
+ mcm5m3m1_ca_w_0_300_s_0_450 = '-5.62500e-07*ic_cap*ic_cap+-3.25000e-07*ic_cap+5.27000e-05'
+ mcm5m3m1_ca_w_0_300_s_0_600 = '-5.62500e-07*ic_cap*ic_cap+-3.25000e-07*ic_cap+5.27000e-05'
+ mcm5m3m1_ca_w_0_300_s_0_800 = '-5.62500e-07*ic_cap*ic_cap+-3.25000e-07*ic_cap+5.27000e-05'
+ mcm5m3m1_ca_w_0_300_s_1_000 = '-5.62500e-07*ic_cap*ic_cap+-3.25000e-07*ic_cap+5.27000e-05'
+ mcm5m3m1_ca_w_0_300_s_1_200 = '-5.62500e-07*ic_cap*ic_cap+-3.25000e-07*ic_cap+5.27000e-05'
+ mcm5m3m1_ca_w_0_300_s_2_100 = '-5.62500e-07*ic_cap*ic_cap+-3.25000e-07*ic_cap+5.27000e-05'
+ mcm5m3m1_ca_w_0_300_s_3_300 = '-5.62500e-07*ic_cap*ic_cap+-3.25000e-07*ic_cap+5.27000e-05'
+ mcm5m3m1_ca_w_0_300_s_9_000 = '-5.62500e-07*ic_cap*ic_cap+-3.25000e-07*ic_cap+5.27000e-05'
+ mcm5m3m1_ca_w_2_400_s_0_300 = '-5.62500e-07*ic_cap*ic_cap+-3.25000e-07*ic_cap+5.27000e-05'
+ mcm5m3m1_ca_w_2_400_s_0_360 = '-5.62500e-07*ic_cap*ic_cap+-3.25000e-07*ic_cap+5.27000e-05'
+ mcm5m3m1_ca_w_2_400_s_0_450 = '-5.62500e-07*ic_cap*ic_cap+-3.25000e-07*ic_cap+5.27000e-05'
+ mcm5m3m1_ca_w_2_400_s_0_600 = '-5.62500e-07*ic_cap*ic_cap+-3.25000e-07*ic_cap+5.27000e-05'
+ mcm5m3m1_ca_w_2_400_s_0_800 = '-5.62500e-07*ic_cap*ic_cap+-3.25000e-07*ic_cap+5.27000e-05'
+ mcm5m3m1_ca_w_2_400_s_1_000 = '-5.62500e-07*ic_cap*ic_cap+-3.25000e-07*ic_cap+5.27000e-05'
+ mcm5m3m1_ca_w_2_400_s_1_200 = '-5.62500e-07*ic_cap*ic_cap+-3.25000e-07*ic_cap+5.27000e-05'
+ mcm5m3m1_ca_w_2_400_s_2_100 = '-5.62500e-07*ic_cap*ic_cap+-3.25000e-07*ic_cap+5.27000e-05'
+ mcm5m3m1_ca_w_2_400_s_3_300 = '-5.62500e-07*ic_cap*ic_cap+-3.25000e-07*ic_cap+5.27000e-05'
+ mcm5m3m1_ca_w_2_400_s_9_000 = '-5.62500e-07*ic_cap*ic_cap+-3.25000e-07*ic_cap+5.27000e-05'
+ mcm5m3m1_cc_w_0_300_s_0_300 = '-7.12500e-13*ic_cap*ic_cap+-4.00000e-13*ic_cap+9.70000e-11'
+ mcm5m3m1_cc_w_0_300_s_0_360 = '-6.15625e-13*ic_cap*ic_cap+-3.37500e-13*ic_cap+8.92000e-11'
+ mcm5m3m1_cc_w_0_300_s_0_450 = '-5.00000e-13*ic_cap*ic_cap+-2.75000e-13*ic_cap+7.89000e-11'
+ mcm5m3m1_cc_w_0_300_s_0_600 = '-3.28125e-13*ic_cap*ic_cap+-1.87500e-13*ic_cap+6.46000e-11'
+ mcm5m3m1_cc_w_0_300_s_0_800 = '-1.78125e-13*ic_cap*ic_cap+-1.12500e-13*ic_cap+5.04000e-11'
+ mcm5m3m1_cc_w_0_300_s_1_000 = '-9.68750e-14*ic_cap*ic_cap+-8.75000e-14*ic_cap+3.99000e-11'
+ mcm5m3m1_cc_w_0_300_s_1_200 = '-4.68750e-14*ic_cap*ic_cap+-3.75000e-14*ic_cap+3.21000e-11'
+ mcm5m3m1_cc_w_0_300_s_2_100 = '5.31250e-14*ic_cap*ic_cap+1.25000e-14*ic_cap+1.34000e-11'
+ mcm5m3m1_cc_w_0_300_s_3_300 = '5.12500e-14*ic_cap*ic_cap+3.00000e-14*ic_cap+4.63000e-12'
+ mcm5m3m1_cc_w_0_300_s_9_000 = '1.56250e-15*ic_cap*ic_cap+2.50000e-15*ic_cap+7.00000e-14'
+ mcm5m3m1_cc_w_2_400_s_0_300 = '-6.00000e-13*ic_cap*ic_cap+-3.25000e-13*ic_cap+1.05000e-10'
+ mcm5m3m1_cc_w_2_400_s_0_360 = '-4.65625e-13*ic_cap*ic_cap+-2.62500e-13*ic_cap+9.57000e-11'
+ mcm5m3m1_cc_w_2_400_s_0_450 = '-3.56250e-13*ic_cap*ic_cap+-2.00000e-13*ic_cap+8.42000e-11'
+ mcm5m3m1_cc_w_2_400_s_0_600 = '-2.31250e-13*ic_cap*ic_cap+-1.25000e-13*ic_cap+6.91000e-11'
+ mcm5m3m1_cc_w_2_400_s_0_800 = '-1.03125e-13*ic_cap*ic_cap+-6.25000e-14*ic_cap+5.39000e-11'
+ mcm5m3m1_cc_w_2_400_s_1_000 = '-2.18750e-14*ic_cap*ic_cap+-3.75000e-14*ic_cap+4.27000e-11'
+ mcm5m3m1_cc_w_2_400_s_1_200 = '2.81250e-14*ic_cap*ic_cap+1.25000e-14*ic_cap+3.43000e-11'
+ mcm5m3m1_cc_w_2_400_s_2_100 = '9.37500e-14*ic_cap*ic_cap+5.00000e-14*ic_cap+1.45000e-11'
+ mcm5m3m1_cc_w_2_400_s_3_300 = '7.15625e-14*ic_cap*ic_cap+4.87500e-14*ic_cap+5.05000e-12'
+ mcm5m3m1_cc_w_2_400_s_9_000 = '4.06250e-15*ic_cap*ic_cap+1.25000e-15*ic_cap+8.00000e-14'
+ mcm5m3m1_cf_w_0_300_s_0_300 = '-2.84375e-14*ic_cap*ic_cap+-1.62500e-14*ic_cap+7.58000e-12'
+ mcm5m3m1_cf_w_0_300_s_0_360 = '-4.21875e-14*ic_cap*ic_cap+-2.37500e-14*ic_cap+9.02000e-12'
+ mcm5m3m1_cf_w_0_300_s_0_450 = '-6.56250e-14*ic_cap*ic_cap+-3.75000e-14*ic_cap+1.12000e-11'
+ mcm5m3m1_cf_w_0_300_s_0_600 = '-9.37500e-14*ic_cap*ic_cap+-5.00000e-14*ic_cap+1.46000e-11'
+ mcm5m3m1_cf_w_0_300_s_0_800 = '-1.37500e-13*ic_cap*ic_cap+-7.50000e-14*ic_cap+1.88000e-11'
+ mcm5m3m1_cf_w_0_300_s_1_000 = '-1.81250e-13*ic_cap*ic_cap+-1.00000e-13*ic_cap+2.28000e-11'
+ mcm5m3m1_cf_w_0_300_s_1_200 = '-2.09375e-13*ic_cap*ic_cap+-1.12500e-13*ic_cap+2.63000e-11'
+ mcm5m3m1_cf_w_0_300_s_2_100 = '-2.90625e-13*ic_cap*ic_cap+-1.62500e-13*ic_cap+3.79000e-11'
+ mcm5m3m1_cf_w_0_300_s_3_300 = '-3.03125e-13*ic_cap*ic_cap+-1.87500e-13*ic_cap+4.53000e-11'
+ mcm5m3m1_cf_w_0_300_s_9_000 = '-2.59375e-13*ic_cap*ic_cap+-1.62500e-13*ic_cap+4.97000e-11'
+ mcm5m3m1_cf_w_2_400_s_0_300 = '-2.68750e-14*ic_cap*ic_cap+-1.50000e-14*ic_cap+7.59000e-12'
+ mcm5m3m1_cf_w_2_400_s_0_360 = '-4.21875e-14*ic_cap*ic_cap+-2.37500e-14*ic_cap+9.05000e-12'
+ mcm5m3m1_cf_w_2_400_s_0_450 = '-6.56250e-14*ic_cap*ic_cap+-3.75000e-14*ic_cap+1.12000e-11'
+ mcm5m3m1_cf_w_2_400_s_0_600 = '-9.68750e-14*ic_cap*ic_cap+-6.25000e-14*ic_cap+1.46000e-11'
+ mcm5m3m1_cf_w_2_400_s_0_800 = '-1.37500e-13*ic_cap*ic_cap+-7.50000e-14*ic_cap+1.89000e-11'
+ mcm5m3m1_cf_w_2_400_s_1_000 = '-1.78125e-13*ic_cap*ic_cap+-1.12500e-13*ic_cap+2.30000e-11'
+ mcm5m3m1_cf_w_2_400_s_1_200 = '-2.06250e-13*ic_cap*ic_cap+-1.25000e-13*ic_cap+2.66000e-11'
+ mcm5m3m1_cf_w_2_400_s_2_100 = '-2.78125e-13*ic_cap*ic_cap+-1.62500e-13*ic_cap+3.86000e-11'
+ mcm5m3m1_cf_w_2_400_s_3_300 = '-2.81250e-13*ic_cap*ic_cap+-1.75000e-13*ic_cap+4.65000e-11'
+ mcm5m3m1_cf_w_2_400_s_9_000 = '-2.25000e-13*ic_cap*ic_cap+-1.50000e-13*ic_cap+5.13000e-11'
+ mcm5m3m2_ca_w_0_300_s_0_300 = '-1.42500e-06*ic_cap*ic_cap+-7.75000e-07*ic_cap+1.02000e-04'
+ mcm5m3m2_ca_w_0_300_s_0_360 = '-1.42500e-06*ic_cap*ic_cap+-7.75000e-07*ic_cap+1.02000e-04'
+ mcm5m3m2_ca_w_0_300_s_0_450 = '-1.42500e-06*ic_cap*ic_cap+-7.75000e-07*ic_cap+1.02000e-04'
+ mcm5m3m2_ca_w_0_300_s_0_600 = '-1.42500e-06*ic_cap*ic_cap+-7.75000e-07*ic_cap+1.02000e-04'
+ mcm5m3m2_ca_w_0_300_s_0_800 = '-1.42500e-06*ic_cap*ic_cap+-7.75000e-07*ic_cap+1.02000e-04'
+ mcm5m3m2_ca_w_0_300_s_1_000 = '-1.42500e-06*ic_cap*ic_cap+-7.75000e-07*ic_cap+1.02000e-04'
+ mcm5m3m2_ca_w_0_300_s_1_200 = '-1.42500e-06*ic_cap*ic_cap+-7.75000e-07*ic_cap+1.02000e-04'
+ mcm5m3m2_ca_w_0_300_s_2_100 = '-1.42500e-06*ic_cap*ic_cap+-7.75000e-07*ic_cap+1.02000e-04'
+ mcm5m3m2_ca_w_0_300_s_3_300 = '-1.42500e-06*ic_cap*ic_cap+-7.75000e-07*ic_cap+1.02000e-04'
+ mcm5m3m2_ca_w_0_300_s_9_000 = '-1.42500e-06*ic_cap*ic_cap+-7.75000e-07*ic_cap+1.02000e-04'
+ mcm5m3m2_ca_w_2_400_s_0_300 = '-1.42500e-06*ic_cap*ic_cap+-7.75000e-07*ic_cap+1.02000e-04'
+ mcm5m3m2_ca_w_2_400_s_0_360 = '-1.42500e-06*ic_cap*ic_cap+-7.75000e-07*ic_cap+1.02000e-04'
+ mcm5m3m2_ca_w_2_400_s_0_450 = '-1.42500e-06*ic_cap*ic_cap+-7.75000e-07*ic_cap+1.02000e-04'
+ mcm5m3m2_ca_w_2_400_s_0_600 = '-1.42500e-06*ic_cap*ic_cap+-7.75000e-07*ic_cap+1.02000e-04'
+ mcm5m3m2_ca_w_2_400_s_0_800 = '-1.42500e-06*ic_cap*ic_cap+-7.75000e-07*ic_cap+1.02000e-04'
+ mcm5m3m2_ca_w_2_400_s_1_000 = '-1.42500e-06*ic_cap*ic_cap+-7.75000e-07*ic_cap+1.02000e-04'
+ mcm5m3m2_ca_w_2_400_s_1_200 = '-1.42500e-06*ic_cap*ic_cap+-7.75000e-07*ic_cap+1.02000e-04'
+ mcm5m3m2_ca_w_2_400_s_2_100 = '-1.42500e-06*ic_cap*ic_cap+-7.75000e-07*ic_cap+1.02000e-04'
+ mcm5m3m2_ca_w_2_400_s_3_300 = '-1.42500e-06*ic_cap*ic_cap+-7.75000e-07*ic_cap+1.02000e-04'
+ mcm5m3m2_ca_w_2_400_s_9_000 = '-1.42500e-06*ic_cap*ic_cap+-7.75000e-07*ic_cap+1.02000e-04'
+ mcm5m3m2_cc_w_0_300_s_0_300 = '-6.25000e-13*ic_cap*ic_cap+-3.25000e-13*ic_cap+8.92000e-11'
+ mcm5m3m2_cc_w_0_300_s_0_360 = '-5.15625e-13*ic_cap*ic_cap+-2.87500e-13*ic_cap+8.10000e-11'
+ mcm5m3m2_cc_w_0_300_s_0_450 = '-4.03125e-13*ic_cap*ic_cap+-2.37500e-13*ic_cap+7.04000e-11'
+ mcm5m3m2_cc_w_0_300_s_0_600 = '-2.53125e-13*ic_cap*ic_cap+-1.62500e-13*ic_cap+5.62000e-11'
+ mcm5m3m2_cc_w_0_300_s_0_800 = '-1.34375e-13*ic_cap*ic_cap+-1.12500e-13*ic_cap+4.23000e-11'
+ mcm5m3m2_cc_w_0_300_s_1_000 = '-5.00000e-14*ic_cap*ic_cap+-7.50000e-14*ic_cap+3.20000e-11'
+ mcm5m3m2_cc_w_0_300_s_1_200 = '-9.37500e-15*ic_cap*ic_cap+-3.75000e-14*ic_cap+2.46000e-11'
+ mcm5m3m2_cc_w_0_300_s_2_100 = '4.43750e-14*ic_cap*ic_cap+2.25000e-14*ic_cap+8.49000e-12'
+ mcm5m3m2_cc_w_0_300_s_3_300 = '3.50000e-14*ic_cap*ic_cap+2.00000e-14*ic_cap+2.28000e-12'
+ mcm5m3m2_cc_w_0_300_s_9_000 = '-1.25000e-15*ic_cap+5.00000e-14'
+ mcm5m3m2_cc_w_2_400_s_0_300 = '-5.28125e-13*ic_cap*ic_cap+-2.87500e-13*ic_cap+9.45000e-11'
+ mcm5m3m2_cc_w_2_400_s_0_360 = '-4.31250e-13*ic_cap*ic_cap+-2.75000e-13*ic_cap+8.58000e-11'
+ mcm5m3m2_cc_w_2_400_s_0_450 = '-3.15625e-13*ic_cap*ic_cap+-1.87500e-13*ic_cap+7.46000e-11'
+ mcm5m3m2_cc_w_2_400_s_0_600 = '-1.87500e-13*ic_cap*ic_cap+-1.00000e-13*ic_cap+5.96000e-11'
+ mcm5m3m2_cc_w_2_400_s_0_800 = '-7.50000e-14*ic_cap*ic_cap+-5.00000e-14*ic_cap+4.49000e-11'
+ mcm5m3m2_cc_w_2_400_s_1_000 = '-1.25000e-14*ic_cap*ic_cap+-2.50000e-14*ic_cap+3.43000e-11'
+ mcm5m3m2_cc_w_2_400_s_1_200 = '3.43750e-14*ic_cap*ic_cap+1.25000e-14*ic_cap+2.64000e-11'
+ mcm5m3m2_cc_w_2_400_s_2_100 = '6.56250e-14*ic_cap*ic_cap+3.75000e-14*ic_cap+9.40000e-12'
+ mcm5m3m2_cc_w_2_400_s_3_300 = '4.25000e-14*ic_cap*ic_cap+3.00000e-14*ic_cap+2.61000e-12'
+ mcm5m3m2_cc_w_2_400_s_9_000 = '9.37500e-16*ic_cap*ic_cap+3.75000e-15*ic_cap+1.00000e-14'
+ mcm5m3m2_cf_w_0_300_s_0_300 = '-9.37500e-14*ic_cap*ic_cap+-5.00000e-14*ic_cap+1.39000e-11'
+ mcm5m3m2_cf_w_0_300_s_0_360 = '-1.31250e-13*ic_cap*ic_cap+-7.50000e-14*ic_cap+1.65000e-11'
+ mcm5m3m2_cf_w_0_300_s_0_450 = '-1.68750e-13*ic_cap*ic_cap+-1.00000e-13*ic_cap+2.00000e-11'
+ mcm5m3m2_cf_w_0_300_s_0_600 = '-2.25000e-13*ic_cap*ic_cap+-1.25000e-13*ic_cap+2.54000e-11'
+ mcm5m3m2_cf_w_0_300_s_0_800 = '-2.90625e-13*ic_cap*ic_cap+-1.62500e-13*ic_cap+3.16000e-11'
+ mcm5m3m2_cf_w_0_300_s_1_000 = '-3.40625e-13*ic_cap*ic_cap+-1.87500e-13*ic_cap+3.70000e-11'
+ mcm5m3m2_cf_w_0_300_s_1_200 = '-3.75000e-13*ic_cap*ic_cap+-2.25000e-13*ic_cap+4.15000e-11'
+ mcm5m3m2_cf_w_0_300_s_2_100 = '-4.25000e-13*ic_cap*ic_cap+-2.50000e-13*ic_cap+5.35000e-11'
+ mcm5m3m2_cf_w_0_300_s_3_300 = '-4.12500e-13*ic_cap*ic_cap+-2.50000e-13*ic_cap+5.91000e-11'
+ mcm5m3m2_cf_w_0_300_s_9_000 = '-3.96875e-13*ic_cap*ic_cap+-2.37500e-13*ic_cap+6.16000e-11'
+ mcm5m3m2_cf_w_2_400_s_0_300 = '-9.68750e-14*ic_cap*ic_cap+-6.25000e-14*ic_cap+1.40000e-11'
+ mcm5m3m2_cf_w_2_400_s_0_360 = '-1.21875e-13*ic_cap*ic_cap+-6.25000e-14*ic_cap+1.64000e-11'
+ mcm5m3m2_cf_w_2_400_s_0_450 = '-1.68750e-13*ic_cap*ic_cap+-1.00000e-13*ic_cap+2.00000e-11'
+ mcm5m3m2_cf_w_2_400_s_0_600 = '-2.25000e-13*ic_cap*ic_cap+-1.25000e-13*ic_cap+2.54000e-11'
+ mcm5m3m2_cf_w_2_400_s_0_800 = '-2.84375e-13*ic_cap*ic_cap+-1.62500e-13*ic_cap+3.17000e-11'
+ mcm5m3m2_cf_w_2_400_s_1_000 = '-3.34375e-13*ic_cap*ic_cap+-1.87500e-13*ic_cap+3.71000e-11'
+ mcm5m3m2_cf_w_2_400_s_1_200 = '-3.65625e-13*ic_cap*ic_cap+-2.12500e-13*ic_cap+4.16000e-11'
+ mcm5m3m2_cf_w_2_400_s_2_100 = '-4.18750e-13*ic_cap*ic_cap+-2.50000e-13*ic_cap+5.43000e-11'
+ mcm5m3m2_cf_w_2_400_s_3_300 = '-4.00000e-13*ic_cap*ic_cap+-2.50000e-13*ic_cap+6.04000e-11'
+ mcm5m3m2_cf_w_2_400_s_9_000 = '-3.65625e-13*ic_cap*ic_cap+-2.12500e-13*ic_cap+6.30000e-11'
+ mcm5m3p1_ca_w_0_300_s_0_300 = '-3.46875e-07*ic_cap*ic_cap+-2.12500e-07*ic_cap+3.57000e-05'
+ mcm5m3p1_ca_w_0_300_s_0_360 = '-3.46875e-07*ic_cap*ic_cap+-2.12500e-07*ic_cap+3.57000e-05'
+ mcm5m3p1_ca_w_0_300_s_0_450 = '-3.46875e-07*ic_cap*ic_cap+-2.12500e-07*ic_cap+3.57000e-05'
+ mcm5m3p1_ca_w_0_300_s_0_600 = '-3.46875e-07*ic_cap*ic_cap+-2.12500e-07*ic_cap+3.57000e-05'
+ mcm5m3p1_ca_w_0_300_s_0_800 = '-3.46875e-07*ic_cap*ic_cap+-2.12500e-07*ic_cap+3.57000e-05'
+ mcm5m3p1_ca_w_0_300_s_1_000 = '-3.46875e-07*ic_cap*ic_cap+-2.12500e-07*ic_cap+3.57000e-05'
+ mcm5m3p1_ca_w_0_300_s_1_200 = '-3.46875e-07*ic_cap*ic_cap+-2.12500e-07*ic_cap+3.57000e-05'
+ mcm5m3p1_ca_w_0_300_s_2_100 = '-3.46875e-07*ic_cap*ic_cap+-2.12500e-07*ic_cap+3.57000e-05'
+ mcm5m3p1_ca_w_0_300_s_3_300 = '-3.46875e-07*ic_cap*ic_cap+-2.12500e-07*ic_cap+3.57000e-05'
+ mcm5m3p1_ca_w_0_300_s_9_000 = '-3.46875e-07*ic_cap*ic_cap+-2.12500e-07*ic_cap+3.57000e-05'
+ mcm5m3p1_ca_w_2_400_s_0_300 = '-3.46875e-07*ic_cap*ic_cap+-2.12500e-07*ic_cap+3.57000e-05'
+ mcm5m3p1_ca_w_2_400_s_0_360 = '-3.46875e-07*ic_cap*ic_cap+-2.12500e-07*ic_cap+3.57000e-05'
+ mcm5m3p1_ca_w_2_400_s_0_450 = '-3.46875e-07*ic_cap*ic_cap+-2.12500e-07*ic_cap+3.57000e-05'
+ mcm5m3p1_ca_w_2_400_s_0_600 = '-3.46875e-07*ic_cap*ic_cap+-2.12500e-07*ic_cap+3.57000e-05'
+ mcm5m3p1_ca_w_2_400_s_0_800 = '-3.46875e-07*ic_cap*ic_cap+-2.12500e-07*ic_cap+3.57000e-05'
+ mcm5m3p1_ca_w_2_400_s_1_000 = '-3.46875e-07*ic_cap*ic_cap+-2.12500e-07*ic_cap+3.57000e-05'
+ mcm5m3p1_ca_w_2_400_s_1_200 = '-3.46875e-07*ic_cap*ic_cap+-2.12500e-07*ic_cap+3.57000e-05'
+ mcm5m3p1_ca_w_2_400_s_2_100 = '-3.46875e-07*ic_cap*ic_cap+-2.12500e-07*ic_cap+3.57000e-05'
+ mcm5m3p1_ca_w_2_400_s_3_300 = '-3.46875e-07*ic_cap*ic_cap+-2.12500e-07*ic_cap+3.57000e-05'
+ mcm5m3p1_ca_w_2_400_s_9_000 = '-3.46875e-07*ic_cap*ic_cap+-2.12500e-07*ic_cap+3.57000e-05'
+ mcm5m3p1_cc_w_0_300_s_0_300 = '-7.62500e-13*ic_cap*ic_cap+-4.25000e-13*ic_cap+1.01000e-10'
+ mcm5m3p1_cc_w_0_300_s_0_360 = '-6.50000e-13*ic_cap*ic_cap+-3.75000e-13*ic_cap+9.32000e-11'
+ mcm5m3p1_cc_w_0_300_s_0_450 = '-5.21875e-13*ic_cap*ic_cap+-3.37500e-13*ic_cap+8.31000e-11'
+ mcm5m3p1_cc_w_0_300_s_0_600 = '-3.90625e-13*ic_cap*ic_cap+-2.37500e-13*ic_cap+6.97000e-11'
+ mcm5m3p1_cc_w_0_300_s_0_800 = '-2.21875e-13*ic_cap*ic_cap+-1.37500e-13*ic_cap+5.57000e-11'
+ mcm5m3p1_cc_w_0_300_s_1_000 = '-1.37500e-13*ic_cap*ic_cap+-1.25000e-13*ic_cap+4.56000e-11'
+ mcm5m3p1_cc_w_0_300_s_1_200 = '-7.81250e-14*ic_cap*ic_cap+-6.25000e-14*ic_cap+3.78000e-11'
+ mcm5m3p1_cc_w_0_300_s_2_100 = '4.06250e-14*ic_cap*ic_cap+1.25000e-14*ic_cap+1.85000e-11'
+ mcm5m3p1_cc_w_0_300_s_3_300 = '6.34375e-14*ic_cap*ic_cap+3.87500e-14*ic_cap+8.07000e-12'
+ mcm5m3p1_cc_w_0_300_s_9_000 = '9.06250e-15*ic_cap*ic_cap+6.25000e-15*ic_cap+2.20000e-13'
+ mcm5m3p1_cc_w_2_400_s_0_300 = '-5.62500e-13*ic_cap*ic_cap+-2.50000e-13*ic_cap+1.12000e-10'
+ mcm5m3p1_cc_w_2_400_s_0_360 = '-5.34375e-13*ic_cap*ic_cap+-2.87500e-13*ic_cap+1.04000e-10'
+ mcm5m3p1_cc_w_2_400_s_0_450 = '-3.68750e-13*ic_cap*ic_cap+-2.25000e-13*ic_cap+9.20000e-11'
+ mcm5m3p1_cc_w_2_400_s_0_600 = '-2.43750e-13*ic_cap*ic_cap+-1.50000e-13*ic_cap+7.69000e-11'
+ mcm5m3p1_cc_w_2_400_s_0_800 = '-1.06250e-13*ic_cap*ic_cap+-7.50000e-14*ic_cap+6.15000e-11'
+ mcm5m3p1_cc_w_2_400_s_1_000 = '-4.06250e-14*ic_cap*ic_cap+-3.75000e-14*ic_cap+5.03000e-11'
+ mcm5m3p1_cc_w_2_400_s_1_200 = '1.25000e-14*ic_cap*ic_cap+4.18000e-11'
+ mcm5m3p1_cc_w_2_400_s_2_100 = '9.68750e-14*ic_cap*ic_cap+6.25000e-14*ic_cap+2.07000e-11'
+ mcm5m3p1_cc_w_2_400_s_3_300 = '9.93750e-14*ic_cap*ic_cap+6.25000e-14*ic_cap+9.06000e-12'
+ mcm5m3p1_cc_w_2_400_s_9_000 = '1.15625e-14*ic_cap*ic_cap+7.50000e-15*ic_cap+2.35000e-13'
+ mcm5m3p1_cf_w_0_300_s_0_300 = '-1.46875e-14*ic_cap*ic_cap+-8.75000e-15*ic_cap+5.19000e-12'
+ mcm5m3p1_cf_w_0_300_s_0_360 = '-2.43750e-14*ic_cap*ic_cap+-1.50000e-14*ic_cap+6.21000e-12'
+ mcm5m3p1_cf_w_0_300_s_0_450 = '-3.81250e-14*ic_cap*ic_cap+-2.25000e-14*ic_cap+7.74000e-12'
+ mcm5m3p1_cf_w_0_300_s_0_600 = '-6.03125e-14*ic_cap*ic_cap+-3.62500e-14*ic_cap+1.02000e-11'
+ mcm5m3p1_cf_w_0_300_s_0_800 = '-8.75000e-14*ic_cap*ic_cap+-5.00000e-14*ic_cap+1.32000e-11'
+ mcm5m3p1_cf_w_0_300_s_1_000 = '-1.18750e-13*ic_cap*ic_cap+-7.50000e-14*ic_cap+1.62000e-11'
+ mcm5m3p1_cf_w_0_300_s_1_200 = '-1.43750e-13*ic_cap*ic_cap+-7.50000e-14*ic_cap+1.89000e-11'
+ mcm5m3p1_cf_w_0_300_s_2_100 = '-2.21875e-13*ic_cap*ic_cap+-1.37500e-13*ic_cap+2.88000e-11'
+ mcm5m3p1_cf_w_0_300_s_3_300 = '-2.53125e-13*ic_cap*ic_cap+-1.62500e-13*ic_cap+3.66000e-11'
+ mcm5m3p1_cf_w_0_300_s_9_000 = '-2.18750e-13*ic_cap*ic_cap+-1.50000e-13*ic_cap+4.38000e-11'
+ mcm5m3p1_cf_w_2_400_s_0_300 = '-1.59375e-14*ic_cap*ic_cap+-8.75000e-15*ic_cap+5.28000e-12'
+ mcm5m3p1_cf_w_2_400_s_0_360 = '-2.37500e-14*ic_cap*ic_cap+-1.50000e-14*ic_cap+6.28000e-12'
+ mcm5m3p1_cf_w_2_400_s_0_450 = '-3.84375e-14*ic_cap*ic_cap+-2.37500e-14*ic_cap+7.78000e-12'
+ mcm5m3p1_cf_w_2_400_s_0_600 = '-6.06250e-14*ic_cap*ic_cap+-3.75000e-14*ic_cap+1.02000e-11'
+ mcm5m3p1_cf_w_2_400_s_0_800 = '-9.37500e-14*ic_cap*ic_cap+-5.00000e-14*ic_cap+1.34000e-11'
+ mcm5m3p1_cf_w_2_400_s_1_000 = '-1.18750e-13*ic_cap*ic_cap+-7.50000e-14*ic_cap+1.64000e-11'
+ mcm5m3p1_cf_w_2_400_s_1_200 = '-1.43750e-13*ic_cap*ic_cap+-7.50000e-14*ic_cap+1.92000e-11'
+ mcm5m3p1_cf_w_2_400_s_2_100 = '-2.18750e-13*ic_cap*ic_cap+-1.25000e-13*ic_cap+2.95000e-11'
+ mcm5m3p1_cf_w_2_400_s_3_300 = '-2.46875e-13*ic_cap*ic_cap+-1.62500e-13*ic_cap+3.80000e-11'
+ mcm5m3p1_cf_w_2_400_s_9_000 = '-1.78125e-13*ic_cap*ic_cap+-1.12500e-13*ic_cap+4.61000e-11'
+ mcm5m4_ca_w_1_600_s_10_000 = '-1.09687e-06*ic_cap*ic_cap+-5.37500e-07*ic_cap+6.84000e-05'
+ mcm5m4_ca_w_1_600_s_12_000 = '-1.09687e-06*ic_cap*ic_cap+-5.37500e-07*ic_cap+6.84000e-05'
+ mcm5m4_ca_w_1_600_s_1_600 = '-1.09687e-06*ic_cap*ic_cap+-5.37500e-07*ic_cap+6.84000e-05'
+ mcm5m4_ca_w_1_600_s_1_700 = '-1.09687e-06*ic_cap*ic_cap+-5.37500e-07*ic_cap+6.84000e-05'
+ mcm5m4_ca_w_1_600_s_1_900 = '-1.09687e-06*ic_cap*ic_cap+-5.37500e-07*ic_cap+6.84000e-05'
+ mcm5m4_ca_w_1_600_s_2_000 = '-1.09687e-06*ic_cap*ic_cap+-5.37500e-07*ic_cap+6.84000e-05'
+ mcm5m4_ca_w_1_600_s_2_400 = '-1.09687e-06*ic_cap*ic_cap+-5.37500e-07*ic_cap+6.84000e-05'
+ mcm5m4_ca_w_1_600_s_2_800 = '-1.09687e-06*ic_cap*ic_cap+-5.37500e-07*ic_cap+6.84000e-05'
+ mcm5m4_ca_w_1_600_s_3_200 = '-1.09687e-06*ic_cap*ic_cap+-5.37500e-07*ic_cap+6.84000e-05'
+ mcm5m4_ca_w_1_600_s_4_800 = '-1.09687e-06*ic_cap*ic_cap+-5.37500e-07*ic_cap+6.84000e-05'
+ mcm5m4_ca_w_4_000_s_10_000 = '-1.09687e-06*ic_cap*ic_cap+-5.37500e-07*ic_cap+6.84000e-05'
+ mcm5m4_ca_w_4_000_s_12_000 = '-1.09687e-06*ic_cap*ic_cap+-5.37500e-07*ic_cap+6.84000e-05'
+ mcm5m4_ca_w_4_000_s_1_600 = '-1.09687e-06*ic_cap*ic_cap+-5.37500e-07*ic_cap+6.84000e-05'
+ mcm5m4_ca_w_4_000_s_1_700 = '-1.09687e-06*ic_cap*ic_cap+-5.37500e-07*ic_cap+6.84000e-05'
+ mcm5m4_ca_w_4_000_s_1_900 = '-1.09687e-06*ic_cap*ic_cap+-5.37500e-07*ic_cap+6.84000e-05'
+ mcm5m4_ca_w_4_000_s_2_000 = '-1.09687e-06*ic_cap*ic_cap+-5.37500e-07*ic_cap+6.84000e-05'
+ mcm5m4_ca_w_4_000_s_2_400 = '-1.09687e-06*ic_cap*ic_cap+-5.37500e-07*ic_cap+6.84000e-05'
+ mcm5m4_ca_w_4_000_s_2_800 = '-1.09687e-06*ic_cap*ic_cap+-5.37500e-07*ic_cap+6.84000e-05'
+ mcm5m4_ca_w_4_000_s_3_200 = '-1.09687e-06*ic_cap*ic_cap+-5.37500e-07*ic_cap+6.84000e-05'
+ mcm5m4_ca_w_4_000_s_4_800 = '-1.09687e-06*ic_cap*ic_cap+-5.37500e-07*ic_cap+6.84000e-05'
+ mcm5m4_cc_w_1_600_s_12_000 = '1.56250e-15*ic_cap*ic_cap+-6.25000e-15*ic_cap+2.95000e-12'
+ mcm5m4_cc_w_1_600_s_1_600 = '-3.21875e-13*ic_cap*ic_cap+-2.37500e-13*ic_cap+5.05000e-11'
+ mcm5m4_cc_w_1_600_s_1_700 = '-2.81250e-13*ic_cap*ic_cap+-2.00000e-13*ic_cap+4.69000e-11'
+ mcm5m4_cc_w_1_600_s_1_900 = '-2.06250e-13*ic_cap*ic_cap+-1.50000e-13*ic_cap+4.09000e-11'
+ mcm5m4_cc_w_1_600_s_2_000 = '-1.78125e-13*ic_cap*ic_cap+-1.37500e-13*ic_cap+3.84000e-11'
+ mcm5m4_cc_w_1_600_s_2_400 = '-1.09375e-13*ic_cap*ic_cap+-8.75000e-14*ic_cap+3.06000e-11'
+ mcm5m4_cc_w_1_600_s_2_800 = '-6.87500e-14*ic_cap*ic_cap+-5.00000e-14*ic_cap+2.51000e-11'
+ mcm5m4_cc_w_1_600_s_3_200 = '-4.68750e-14*ic_cap*ic_cap+-3.75000e-14*ic_cap+2.11000e-11'
+ mcm5m4_cc_w_1_600_s_4_800 = '-3.12500e-15*ic_cap*ic_cap+-1.25000e-14*ic_cap+1.20000e-11'
+ mcm5m4_cc_w_4_000_s_10_000 = '3.12500e-15*ic_cap*ic_cap+6.00000e-12'
+ mcm5m4_cc_w_4_000_s_12_000 = '4.68750e-15*ic_cap*ic_cap+6.25000e-15*ic_cap+4.60000e-12'
+ mcm5m4_cc_w_4_000_s_1_600 = '-3.12500e-13*ic_cap*ic_cap+-2.25000e-13*ic_cap+5.57000e-11'
+ mcm5m4_cc_w_4_000_s_1_700 = '-2.71875e-13*ic_cap*ic_cap+-1.87500e-13*ic_cap+5.21000e-11'
+ mcm5m4_cc_w_4_000_s_1_900 = '-2.00000e-13*ic_cap*ic_cap+-1.50000e-13*ic_cap+4.59000e-11'
+ mcm5m4_cc_w_4_000_s_2_000 = '-1.71875e-13*ic_cap*ic_cap+-1.37500e-13*ic_cap+4.33000e-11'
+ mcm5m4_cc_w_4_000_s_2_400 = '-1.03125e-13*ic_cap*ic_cap+-8.75000e-14*ic_cap+3.52000e-11'
+ mcm5m4_cc_w_4_000_s_2_800 = '-5.93750e-14*ic_cap*ic_cap+-6.25000e-14*ic_cap+2.95000e-11'
+ mcm5m4_cc_w_4_000_s_3_200 = '-3.43750e-14*ic_cap*ic_cap+-3.75000e-14*ic_cap+2.52000e-11'
+ mcm5m4_cc_w_4_000_s_4_800 = '-3.12500e-15*ic_cap*ic_cap+-1.25000e-14*ic_cap+1.56000e-11'
+ mcm5m4_cf_w_1_600_s_10_000 = '-5.84375e-13*ic_cap*ic_cap+-3.37500e-13*ic_cap+6.96000e-11'
+ mcm5m4_cf_w_1_600_s_12_000 = '-5.84375e-13*ic_cap*ic_cap+-3.37500e-13*ic_cap+7.06000e-11'
+ mcm5m4_cf_w_1_600_s_1_600 = '-4.03125e-13*ic_cap*ic_cap+-2.12500e-13*ic_cap+3.82000e-11'
+ mcm5m4_cf_w_1_600_s_1_700 = '-4.21875e-13*ic_cap*ic_cap+-2.12500e-13*ic_cap+3.97000e-11'
+ mcm5m4_cf_w_1_600_s_1_900 = '-4.43750e-13*ic_cap*ic_cap+-2.25000e-13*ic_cap+4.24000e-11'
+ mcm5m4_cf_w_1_600_s_2_000 = '-4.59375e-13*ic_cap*ic_cap+-2.37500e-13*ic_cap+4.37000e-11'
+ mcm5m4_cf_w_1_600_s_2_400 = '-4.96875e-13*ic_cap*ic_cap+-2.62500e-13*ic_cap+4.81000e-11'
+ mcm5m4_cf_w_1_600_s_2_800 = '-5.21875e-13*ic_cap*ic_cap+-2.87500e-13*ic_cap+5.17000e-11'
+ mcm5m4_cf_w_1_600_s_3_200 = '-5.37500e-13*ic_cap*ic_cap+-3.00000e-13*ic_cap+5.45000e-11'
+ mcm5m4_cf_w_1_600_s_4_800 = '-5.68750e-13*ic_cap*ic_cap+-3.25000e-13*ic_cap+6.19000e-11'
+ mcm5m4_cf_w_4_000_s_10_000 = '-5.78125e-13*ic_cap*ic_cap+-3.37500e-13*ic_cap+7.12000e-11'
+ mcm5m4_cf_w_4_000_s_12_000 = '-5.78125e-13*ic_cap*ic_cap+-3.37500e-13*ic_cap+7.26000e-11'
+ mcm5m4_cf_w_4_000_s_1_600 = '-4.03125e-13*ic_cap*ic_cap+-2.12500e-13*ic_cap+3.82000e-11'
+ mcm5m4_cf_w_4_000_s_1_700 = '-4.21875e-13*ic_cap*ic_cap+-2.12500e-13*ic_cap+3.97000e-11'
+ mcm5m4_cf_w_4_000_s_1_900 = '-4.40625e-13*ic_cap*ic_cap+-2.37500e-13*ic_cap+4.24000e-11'
+ mcm5m4_cf_w_4_000_s_2_000 = '-4.59375e-13*ic_cap*ic_cap+-2.37500e-13*ic_cap+4.37000e-11'
+ mcm5m4_cf_w_4_000_s_2_400 = '-5.00000e-13*ic_cap*ic_cap+-2.75000e-13*ic_cap+4.82000e-11'
+ mcm5m4_cf_w_4_000_s_2_800 = '-5.18750e-13*ic_cap*ic_cap+-2.75000e-13*ic_cap+5.17000e-11'
+ mcm5m4_cf_w_4_000_s_3_200 = '-5.34375e-13*ic_cap*ic_cap+-2.87500e-13*ic_cap+5.46000e-11'
+ mcm5m4_cf_w_4_000_s_4_800 = '-5.68750e-13*ic_cap*ic_cap+-3.25000e-13*ic_cap+6.23000e-11'
+ mcm5m4d_ca_w_0_300_s_0_300 = '-1.17812e-06*ic_cap*ic_cap+-5.87500e-07*ic_cap+7.78000e-05'
+ mcm5m4d_ca_w_0_300_s_0_360 = '-1.17812e-06*ic_cap*ic_cap+-5.87500e-07*ic_cap+7.78000e-05'
+ mcm5m4d_ca_w_0_300_s_0_450 = '-1.17812e-06*ic_cap*ic_cap+-5.87500e-07*ic_cap+7.78000e-05'
+ mcm5m4d_ca_w_0_300_s_0_600 = '-1.17812e-06*ic_cap*ic_cap+-5.87500e-07*ic_cap+7.78000e-05'
+ mcm5m4d_ca_w_0_300_s_0_800 = '-1.17812e-06*ic_cap*ic_cap+-5.87500e-07*ic_cap+7.78000e-05'
+ mcm5m4d_ca_w_0_300_s_1_000 = '-1.17812e-06*ic_cap*ic_cap+-5.87500e-07*ic_cap+7.78000e-05'
+ mcm5m4d_ca_w_0_300_s_1_200 = '-1.17812e-06*ic_cap*ic_cap+-5.87500e-07*ic_cap+7.78000e-05'
+ mcm5m4d_ca_w_0_300_s_2_100 = '-1.17812e-06*ic_cap*ic_cap+-5.87500e-07*ic_cap+7.78000e-05'
+ mcm5m4d_ca_w_0_300_s_3_300 = '-1.17812e-06*ic_cap*ic_cap+-5.87500e-07*ic_cap+7.78000e-05'
+ mcm5m4d_ca_w_0_300_s_9_000 = '-1.17812e-06*ic_cap*ic_cap+-5.87500e-07*ic_cap+7.78000e-05'
+ mcm5m4d_ca_w_2_400_s_0_300 = '-1.17812e-06*ic_cap*ic_cap+-5.87500e-07*ic_cap+7.78000e-05'
+ mcm5m4d_ca_w_2_400_s_0_360 = '-1.17812e-06*ic_cap*ic_cap+-5.87500e-07*ic_cap+7.78000e-05'
+ mcm5m4d_ca_w_2_400_s_0_450 = '-1.17812e-06*ic_cap*ic_cap+-5.87500e-07*ic_cap+7.78000e-05'
+ mcm5m4d_ca_w_2_400_s_0_600 = '-1.17812e-06*ic_cap*ic_cap+-5.87500e-07*ic_cap+7.78000e-05'
+ mcm5m4d_ca_w_2_400_s_0_800 = '-1.17812e-06*ic_cap*ic_cap+-5.87500e-07*ic_cap+7.78000e-05'
+ mcm5m4d_ca_w_2_400_s_1_000 = '-1.17812e-06*ic_cap*ic_cap+-5.87500e-07*ic_cap+7.78000e-05'
+ mcm5m4d_ca_w_2_400_s_1_200 = '-1.17812e-06*ic_cap*ic_cap+-5.87500e-07*ic_cap+7.78000e-05'
+ mcm5m4d_ca_w_2_400_s_2_100 = '-1.17812e-06*ic_cap*ic_cap+-5.87500e-07*ic_cap+7.78000e-05'
+ mcm5m4d_ca_w_2_400_s_3_300 = '-1.17812e-06*ic_cap*ic_cap+-5.87500e-07*ic_cap+7.78000e-05'
+ mcm5m4d_ca_w_2_400_s_9_000 = '-1.17812e-06*ic_cap*ic_cap+-5.87500e-07*ic_cap+7.78000e-05'
+ mcm5m4d_cc_w_0_300_s_0_300 = '-6.18750e-13*ic_cap*ic_cap+-3.50000e-13*ic_cap+9.36000e-11'
+ mcm5m4d_cc_w_0_300_s_0_360 = '-5.56250e-13*ic_cap*ic_cap+-3.25000e-13*ic_cap+8.61000e-11'
+ mcm5m4d_cc_w_0_300_s_0_450 = '-4.28125e-13*ic_cap*ic_cap+-2.87500e-13*ic_cap+7.56000e-11'
+ mcm5m4d_cc_w_0_300_s_0_600 = '-2.81250e-13*ic_cap*ic_cap+-1.75000e-13*ic_cap+6.17000e-11'
+ mcm5m4d_cc_w_0_300_s_0_800 = '-1.65625e-13*ic_cap*ic_cap+-1.12500e-13*ic_cap+4.82000e-11'
+ mcm5m4d_cc_w_0_300_s_1_000 = '-7.81250e-14*ic_cap*ic_cap+-8.75000e-14*ic_cap+3.82000e-11'
+ mcm5m4d_cc_w_0_300_s_1_200 = '-3.12500e-14*ic_cap*ic_cap+-5.00000e-14*ic_cap+3.08000e-11'
+ mcm5m4d_cc_w_0_300_s_2_100 = '3.43750e-14*ic_cap*ic_cap+1.25000e-14*ic_cap+1.35000e-11'
+ mcm5m4d_cc_w_0_300_s_3_300 = '4.34375e-14*ic_cap*ic_cap+2.37500e-14*ic_cap+5.39000e-12'
+ mcm5m4d_cc_w_0_300_s_9_000 = '5.62500e-15*ic_cap*ic_cap+1.25000e-15*ic_cap+1.45000e-13'
+ mcm5m4d_cc_w_2_400_s_0_300 = '-5.62500e-13*ic_cap*ic_cap+-3.25000e-13*ic_cap+1.04000e-10'
+ mcm5m4d_cc_w_2_400_s_0_360 = '-4.53125e-13*ic_cap*ic_cap+-2.87500e-13*ic_cap+9.52000e-11'
+ mcm5m4d_cc_w_2_400_s_0_450 = '-3.37500e-13*ic_cap*ic_cap+-1.75000e-13*ic_cap+8.40000e-11'
+ mcm5m4d_cc_w_2_400_s_0_600 = '-2.06250e-13*ic_cap*ic_cap+-1.25000e-13*ic_cap+6.90000e-11'
+ mcm5m4d_cc_w_2_400_s_0_800 = '-9.37500e-14*ic_cap*ic_cap+-5.00000e-14*ic_cap+5.42000e-11'
+ mcm5m4d_cc_w_2_400_s_1_000 = '-1.56250e-14*ic_cap*ic_cap+-3.75000e-14*ic_cap+4.33000e-11'
+ mcm5m4d_cc_w_2_400_s_1_200 = '2.50000e-14*ic_cap*ic_cap+3.52000e-11'
+ mcm5m4d_cc_w_2_400_s_2_100 = '8.12500e-14*ic_cap*ic_cap+5.00000e-14*ic_cap+1.63000e-11'
+ mcm5m4d_cc_w_2_400_s_3_300 = '6.93750e-14*ic_cap*ic_cap+4.50000e-14*ic_cap+6.86000e-12'
+ mcm5m4d_cc_w_2_400_s_9_000 = '8.12500e-15*ic_cap*ic_cap+1.00000e-14*ic_cap+2.25000e-13'
+ mcm5m4d_cf_w_0_300_s_0_300 = '-7.84375e-14*ic_cap*ic_cap+-3.62500e-14*ic_cap+1.02000e-11'
+ mcm5m4d_cf_w_0_300_s_0_360 = '-1.06250e-13*ic_cap*ic_cap+-5.00000e-14*ic_cap+1.21000e-11'
+ mcm5m4d_cf_w_0_300_s_0_450 = '-1.34375e-13*ic_cap*ic_cap+-6.25000e-14*ic_cap+1.48000e-11'
+ mcm5m4d_cf_w_0_300_s_0_600 = '-1.81250e-13*ic_cap*ic_cap+-1.00000e-13*ic_cap+1.90000e-11'
+ mcm5m4d_cf_w_0_300_s_0_800 = '-2.37500e-13*ic_cap*ic_cap+-1.25000e-13*ic_cap+2.39000e-11'
+ mcm5m4d_cf_w_0_300_s_1_000 = '-2.81250e-13*ic_cap*ic_cap+-1.50000e-13*ic_cap+2.83000e-11'
+ mcm5m4d_cf_w_0_300_s_1_200 = '-3.12500e-13*ic_cap*ic_cap+-1.75000e-13*ic_cap+3.21000e-11'
+ mcm5m4d_cf_w_0_300_s_2_100 = '-3.78125e-13*ic_cap*ic_cap+-2.12500e-13*ic_cap+4.36000e-11'
+ mcm5m4d_cf_w_0_300_s_3_300 = '-3.81250e-13*ic_cap*ic_cap+-2.25000e-13*ic_cap+5.04000e-11'
+ mcm5m4d_cf_w_0_300_s_9_000 = '-3.56250e-13*ic_cap*ic_cap+-2.00000e-13*ic_cap+5.54000e-11'
+ mcm5m4d_cf_w_2_400_s_0_300 = '-7.93750e-14*ic_cap*ic_cap+-3.75000e-14*ic_cap+1.03000e-11'
+ mcm5m4d_cf_w_2_400_s_0_360 = '-1.06250e-13*ic_cap*ic_cap+-5.00000e-14*ic_cap+1.22000e-11'
+ mcm5m4d_cf_w_2_400_s_0_450 = '-1.37500e-13*ic_cap*ic_cap+-7.50000e-14*ic_cap+1.49000e-11'
+ mcm5m4d_cf_w_2_400_s_0_600 = '-1.84375e-13*ic_cap*ic_cap+-8.75000e-14*ic_cap+1.91000e-11'
+ mcm5m4d_cf_w_2_400_s_0_800 = '-2.37500e-13*ic_cap*ic_cap+-1.25000e-13*ic_cap+2.41000e-11'
+ mcm5m4d_cf_w_2_400_s_1_000 = '-2.75000e-13*ic_cap*ic_cap+-1.50000e-13*ic_cap+2.85000e-11'
+ mcm5m4d_cf_w_2_400_s_1_200 = '-3.03125e-13*ic_cap*ic_cap+-1.62500e-13*ic_cap+3.23000e-11'
+ mcm5m4d_cf_w_2_400_s_2_100 = '-3.65625e-13*ic_cap*ic_cap+-2.12500e-13*ic_cap+4.42000e-11'
+ mcm5m4d_cf_w_2_400_s_3_300 = '-3.71875e-13*ic_cap*ic_cap+-2.12500e-13*ic_cap+5.20000e-11'
+ mcm5m4d_cf_w_2_400_s_9_000 = '-3.21875e-13*ic_cap*ic_cap+-1.87500e-13*ic_cap+5.84000e-11'
+ mcm5m4f_ca_w_0_300_s_0_300 = '-1.17188e-06*ic_cap*ic_cap+-5.87500e-07*ic_cap+7.70000e-05'
+ mcm5m4f_ca_w_0_300_s_0_360 = '-1.17188e-06*ic_cap*ic_cap+-5.87500e-07*ic_cap+7.70000e-05'
+ mcm5m4f_ca_w_0_300_s_0_450 = '-1.17188e-06*ic_cap*ic_cap+-5.87500e-07*ic_cap+7.70000e-05'
+ mcm5m4f_ca_w_0_300_s_0_600 = '-1.17188e-06*ic_cap*ic_cap+-5.87500e-07*ic_cap+7.70000e-05'
+ mcm5m4f_ca_w_0_300_s_0_800 = '-1.17188e-06*ic_cap*ic_cap+-5.87500e-07*ic_cap+7.70000e-05'
+ mcm5m4f_ca_w_0_300_s_1_000 = '-1.17188e-06*ic_cap*ic_cap+-5.87500e-07*ic_cap+7.70000e-05'
+ mcm5m4f_ca_w_0_300_s_1_200 = '-1.17188e-06*ic_cap*ic_cap+-5.87500e-07*ic_cap+7.70000e-05'
+ mcm5m4f_ca_w_0_300_s_2_100 = '-1.17188e-06*ic_cap*ic_cap+-5.87500e-07*ic_cap+7.70000e-05'
+ mcm5m4f_ca_w_0_300_s_3_300 = '-1.17188e-06*ic_cap*ic_cap+-5.87500e-07*ic_cap+7.70000e-05'
+ mcm5m4f_ca_w_0_300_s_9_000 = '-1.17188e-06*ic_cap*ic_cap+-5.87500e-07*ic_cap+7.70000e-05'
+ mcm5m4f_ca_w_2_400_s_0_300 = '-1.17188e-06*ic_cap*ic_cap+-5.87500e-07*ic_cap+7.70000e-05'
+ mcm5m4f_ca_w_2_400_s_0_360 = '-1.17188e-06*ic_cap*ic_cap+-5.87500e-07*ic_cap+7.70000e-05'
+ mcm5m4f_ca_w_2_400_s_0_450 = '-1.17188e-06*ic_cap*ic_cap+-5.87500e-07*ic_cap+7.70000e-05'
+ mcm5m4f_ca_w_2_400_s_0_600 = '-1.17188e-06*ic_cap*ic_cap+-5.87500e-07*ic_cap+7.70000e-05'
+ mcm5m4f_ca_w_2_400_s_0_800 = '-1.17188e-06*ic_cap*ic_cap+-5.87500e-07*ic_cap+7.70000e-05'
+ mcm5m4f_ca_w_2_400_s_1_000 = '-1.17188e-06*ic_cap*ic_cap+-5.87500e-07*ic_cap+7.70000e-05'
+ mcm5m4f_ca_w_2_400_s_1_200 = '-1.17188e-06*ic_cap*ic_cap+-5.87500e-07*ic_cap+7.70000e-05'
+ mcm5m4f_ca_w_2_400_s_2_100 = '-1.17188e-06*ic_cap*ic_cap+-5.87500e-07*ic_cap+7.70000e-05'
+ mcm5m4f_ca_w_2_400_s_3_300 = '-1.17188e-06*ic_cap*ic_cap+-5.87500e-07*ic_cap+7.70000e-05'
+ mcm5m4f_ca_w_2_400_s_9_000 = '-1.17188e-06*ic_cap*ic_cap+-5.87500e-07*ic_cap+7.70000e-05'
+ mcm5m4f_cc_w_0_300_s_0_300 = '-6.21875e-13*ic_cap*ic_cap+-3.37500e-13*ic_cap+9.38000e-11'
+ mcm5m4f_cc_w_0_300_s_0_360 = '-5.62500e-13*ic_cap*ic_cap+-3.25000e-13*ic_cap+8.64000e-11'
+ mcm5m4f_cc_w_0_300_s_0_450 = '-4.28125e-13*ic_cap*ic_cap+-2.87500e-13*ic_cap+7.58000e-11'
+ mcm5m4f_cc_w_0_300_s_0_600 = '-2.84375e-13*ic_cap*ic_cap+-1.87500e-13*ic_cap+6.20000e-11'
+ mcm5m4f_cc_w_0_300_s_0_800 = '-1.56250e-13*ic_cap*ic_cap+-1.25000e-13*ic_cap+4.84000e-11'
+ mcm5m4f_cc_w_0_300_s_1_000 = '-7.18750e-14*ic_cap*ic_cap+-8.75000e-14*ic_cap+3.85000e-11'
+ mcm5m4f_cc_w_0_300_s_1_200 = '-3.43750e-14*ic_cap*ic_cap+-3.75000e-14*ic_cap+3.12000e-11'
+ mcm5m4f_cc_w_0_300_s_2_100 = '3.43750e-14*ic_cap*ic_cap+1.25000e-14*ic_cap+1.39000e-11'
+ mcm5m4f_cc_w_0_300_s_3_300 = '4.25000e-14*ic_cap*ic_cap+2.25000e-14*ic_cap+5.70000e-12'
+ mcm5m4f_cc_w_0_300_s_9_000 = '4.21875e-15*ic_cap*ic_cap+6.25000e-16*ic_cap+2.30000e-13'
+ mcm5m4f_cc_w_2_400_s_0_300 = '-5.18750e-13*ic_cap*ic_cap+-3.25000e-13*ic_cap+1.04000e-10'
+ mcm5m4f_cc_w_2_400_s_0_360 = '-4.43750e-13*ic_cap*ic_cap+-2.75000e-13*ic_cap+9.57000e-11'
+ mcm5m4f_cc_w_2_400_s_0_450 = '-3.37500e-13*ic_cap*ic_cap+-1.75000e-13*ic_cap+8.47000e-11'
+ mcm5m4f_cc_w_2_400_s_0_600 = '-2.03125e-13*ic_cap*ic_cap+-1.37500e-13*ic_cap+6.97000e-11'
+ mcm5m4f_cc_w_2_400_s_0_800 = '-9.06250e-14*ic_cap*ic_cap+-6.25000e-14*ic_cap+5.49000e-11'
+ mcm5m4f_cc_w_2_400_s_1_000 = '-1.25000e-14*ic_cap*ic_cap+-2.50000e-14*ic_cap+4.39000e-11'
+ mcm5m4f_cc_w_2_400_s_1_200 = '3.12500e-14*ic_cap*ic_cap+3.59000e-11'
+ mcm5m4f_cc_w_2_400_s_2_100 = '8.12500e-14*ic_cap*ic_cap+5.00000e-14*ic_cap+1.70000e-11'
+ mcm5m4f_cc_w_2_400_s_3_300 = '7.25000e-14*ic_cap*ic_cap+4.25000e-14*ic_cap+7.38000e-12'
+ mcm5m4f_cc_w_2_400_s_9_000 = '5.78125e-15*ic_cap*ic_cap+8.12500e-15*ic_cap+3.05000e-13'
+ mcm5m4f_cf_w_0_300_s_0_300 = '-7.93750e-14*ic_cap*ic_cap+-3.75000e-14*ic_cap+1.01000e-11'
+ mcm5m4f_cf_w_0_300_s_0_360 = '-1.06250e-13*ic_cap*ic_cap+-5.00000e-14*ic_cap+1.20000e-11'
+ mcm5m4f_cf_w_0_300_s_0_450 = '-1.40625e-13*ic_cap*ic_cap+-6.25000e-14*ic_cap+1.47000e-11'
+ mcm5m4f_cf_w_0_300_s_0_600 = '-1.84375e-13*ic_cap*ic_cap+-8.75000e-14*ic_cap+1.88000e-11'
+ mcm5m4f_cf_w_0_300_s_0_800 = '-2.37500e-13*ic_cap*ic_cap+-1.25000e-13*ic_cap+2.37000e-11'
+ mcm5m4f_cf_w_0_300_s_1_000 = '-2.81250e-13*ic_cap*ic_cap+-1.50000e-13*ic_cap+2.80000e-11'
+ mcm5m4f_cf_w_0_300_s_1_200 = '-3.12500e-13*ic_cap*ic_cap+-1.75000e-13*ic_cap+3.17000e-11'
+ mcm5m4f_cf_w_0_300_s_2_100 = '-3.71875e-13*ic_cap*ic_cap+-2.12500e-13*ic_cap+4.31000e-11'
+ mcm5m4f_cf_w_0_300_s_3_300 = '-3.87500e-13*ic_cap*ic_cap+-2.25000e-13*ic_cap+5.01000e-11'
+ mcm5m4f_cf_w_0_300_s_9_000 = '-3.56250e-13*ic_cap*ic_cap+-2.00000e-13*ic_cap+5.53000e-11'
+ mcm5m4f_cf_w_2_400_s_0_300 = '-8.06250e-14*ic_cap*ic_cap+-3.75000e-14*ic_cap+1.02000e-11'
+ mcm5m4f_cf_w_2_400_s_0_360 = '-1.06250e-13*ic_cap*ic_cap+-5.00000e-14*ic_cap+1.21000e-11'
+ mcm5m4f_cf_w_2_400_s_0_450 = '-1.34375e-13*ic_cap*ic_cap+-6.25000e-14*ic_cap+1.47000e-11'
+ mcm5m4f_cf_w_2_400_s_0_600 = '-1.87500e-13*ic_cap*ic_cap+-1.00000e-13*ic_cap+1.89000e-11'
+ mcm5m4f_cf_w_2_400_s_0_800 = '-2.31250e-13*ic_cap*ic_cap+-1.25000e-13*ic_cap+2.38000e-11'
+ mcm5m4f_cf_w_2_400_s_1_000 = '-2.68750e-13*ic_cap*ic_cap+-1.50000e-13*ic_cap+2.81000e-11'
+ mcm5m4f_cf_w_2_400_s_1_200 = '-3.03125e-13*ic_cap*ic_cap+-1.62500e-13*ic_cap+3.19000e-11'
+ mcm5m4f_cf_w_2_400_s_2_100 = '-3.68750e-13*ic_cap*ic_cap+-2.00000e-13*ic_cap+4.38000e-11'
+ mcm5m4f_cf_w_2_400_s_3_300 = '-3.78125e-13*ic_cap*ic_cap+-2.12500e-13*ic_cap+5.17000e-11'
+ mcm5m4f_cf_w_2_400_s_9_000 = '-3.25000e-13*ic_cap*ic_cap+-1.75000e-13*ic_cap+5.85000e-11'
+ mcm5m4l1_ca_w_0_300_s_0_300 = '-1.19375e-06*ic_cap*ic_cap+-6.00000e-07*ic_cap+8.01000e-05'
+ mcm5m4l1_ca_w_0_300_s_0_360 = '-1.19375e-06*ic_cap*ic_cap+-6.00000e-07*ic_cap+8.01000e-05'
+ mcm5m4l1_ca_w_0_300_s_0_450 = '-1.19375e-06*ic_cap*ic_cap+-6.00000e-07*ic_cap+8.01000e-05'
+ mcm5m4l1_ca_w_0_300_s_0_600 = '-1.19375e-06*ic_cap*ic_cap+-6.00000e-07*ic_cap+8.01000e-05'
+ mcm5m4l1_ca_w_0_300_s_0_800 = '-1.19375e-06*ic_cap*ic_cap+-6.00000e-07*ic_cap+8.01000e-05'
+ mcm5m4l1_ca_w_0_300_s_1_000 = '-1.19375e-06*ic_cap*ic_cap+-6.00000e-07*ic_cap+8.01000e-05'
+ mcm5m4l1_ca_w_0_300_s_1_200 = '-1.19375e-06*ic_cap*ic_cap+-6.00000e-07*ic_cap+8.01000e-05'
+ mcm5m4l1_ca_w_0_300_s_2_100 = '-1.19375e-06*ic_cap*ic_cap+-6.00000e-07*ic_cap+8.01000e-05'
+ mcm5m4l1_ca_w_0_300_s_3_300 = '-1.19375e-06*ic_cap*ic_cap+-6.00000e-07*ic_cap+8.01000e-05'
+ mcm5m4l1_ca_w_0_300_s_9_000 = '-1.19375e-06*ic_cap*ic_cap+-6.00000e-07*ic_cap+8.01000e-05'
+ mcm5m4l1_ca_w_2_400_s_0_300 = '-1.19375e-06*ic_cap*ic_cap+-6.00000e-07*ic_cap+8.01000e-05'
+ mcm5m4l1_ca_w_2_400_s_0_360 = '-1.19375e-06*ic_cap*ic_cap+-6.00000e-07*ic_cap+8.01000e-05'
+ mcm5m4l1_ca_w_2_400_s_0_450 = '-1.19375e-06*ic_cap*ic_cap+-6.00000e-07*ic_cap+8.01000e-05'
+ mcm5m4l1_ca_w_2_400_s_0_600 = '-1.19375e-06*ic_cap*ic_cap+-6.00000e-07*ic_cap+8.01000e-05'
+ mcm5m4l1_ca_w_2_400_s_0_800 = '-1.19375e-06*ic_cap*ic_cap+-6.00000e-07*ic_cap+8.01000e-05'
+ mcm5m4l1_ca_w_2_400_s_1_000 = '-1.19375e-06*ic_cap*ic_cap+-6.00000e-07*ic_cap+8.01000e-05'
+ mcm5m4l1_ca_w_2_400_s_1_200 = '-1.19375e-06*ic_cap*ic_cap+-6.00000e-07*ic_cap+8.01000e-05'
+ mcm5m4l1_ca_w_2_400_s_2_100 = '-1.19375e-06*ic_cap*ic_cap+-6.00000e-07*ic_cap+8.01000e-05'
+ mcm5m4l1_ca_w_2_400_s_3_300 = '-1.19375e-06*ic_cap*ic_cap+-6.00000e-07*ic_cap+8.01000e-05'
+ mcm5m4l1_ca_w_2_400_s_9_000 = '-1.19375e-06*ic_cap*ic_cap+-6.00000e-07*ic_cap+8.01000e-05'
+ mcm5m4l1_cc_w_0_300_s_0_300 = '-6.18750e-13*ic_cap*ic_cap+-3.75000e-13*ic_cap+9.30000e-11'
+ mcm5m4l1_cc_w_0_300_s_0_360 = '-5.53125e-13*ic_cap*ic_cap+-3.37500e-13*ic_cap+8.55000e-11'
+ mcm5m4l1_cc_w_0_300_s_0_450 = '-4.21875e-13*ic_cap*ic_cap+-2.62500e-13*ic_cap+7.50000e-11'
+ mcm5m4l1_cc_w_0_300_s_0_600 = '-2.68750e-13*ic_cap*ic_cap+-1.75000e-13*ic_cap+6.08000e-11'
+ mcm5m4l1_cc_w_0_300_s_0_800 = '-1.53125e-13*ic_cap*ic_cap+-1.12500e-13*ic_cap+4.72000e-11'
+ mcm5m4l1_cc_w_0_300_s_1_000 = '-6.87500e-14*ic_cap*ic_cap+-7.50000e-14*ic_cap+3.71000e-11'
+ mcm5m4l1_cc_w_0_300_s_1_200 = '-1.56250e-14*ic_cap*ic_cap+-3.75000e-14*ic_cap+2.96000e-11'
+ mcm5m4l1_cc_w_0_300_s_2_100 = '4.37500e-14*ic_cap*ic_cap+2.50000e-14*ic_cap+1.24000e-11'
+ mcm5m4l1_cc_w_0_300_s_3_300 = '4.09375e-14*ic_cap*ic_cap+2.37500e-14*ic_cap+4.60000e-12'
+ mcm5m4l1_cc_w_0_300_s_9_000 = '3.12500e-16*ic_cap*ic_cap+3.75000e-15*ic_cap+1.60000e-13'
+ mcm5m4l1_cc_w_2_400_s_0_300 = '-5.46875e-13*ic_cap*ic_cap+-3.12500e-13*ic_cap+1.02000e-10'
+ mcm5m4l1_cc_w_2_400_s_0_360 = '-4.46875e-13*ic_cap*ic_cap+-2.62500e-13*ic_cap+9.33000e-11'
+ mcm5m4l1_cc_w_2_400_s_0_450 = '-3.31250e-13*ic_cap*ic_cap+-2.00000e-13*ic_cap+8.20000e-11'
+ mcm5m4l1_cc_w_2_400_s_0_600 = '-1.93750e-13*ic_cap*ic_cap+-1.25000e-13*ic_cap+6.70000e-11'
+ mcm5m4l1_cc_w_2_400_s_0_800 = '-8.43750e-14*ic_cap*ic_cap+-6.25000e-14*ic_cap+5.22000e-11'
+ mcm5m4l1_cc_w_2_400_s_1_000 = '-6.25000e-15*ic_cap*ic_cap+-2.50000e-14*ic_cap+4.12000e-11'
+ mcm5m4l1_cc_w_2_400_s_1_200 = '3.12500e-14*ic_cap*ic_cap+3.32000e-11'
+ mcm5m4l1_cc_w_2_400_s_2_100 = '8.43750e-14*ic_cap*ic_cap+3.75000e-14*ic_cap+1.45000e-11'
+ mcm5m4l1_cc_w_2_400_s_3_300 = '6.84375e-14*ic_cap*ic_cap+4.37500e-14*ic_cap+5.55000e-12'
+ mcm5m4l1_cc_w_2_400_s_9_000 = '6.87500e-15*ic_cap*ic_cap+2.50000e-15*ic_cap+8.50000e-14'
+ mcm5m4l1_cf_w_0_300_s_0_300 = '-7.68750e-14*ic_cap*ic_cap+-3.75000e-14*ic_cap+1.05000e-11'
+ mcm5m4l1_cf_w_0_300_s_0_360 = '-1.06250e-13*ic_cap*ic_cap+-5.00000e-14*ic_cap+1.25000e-11'
+ mcm5m4l1_cf_w_0_300_s_0_450 = '-1.37500e-13*ic_cap*ic_cap+-7.50000e-14*ic_cap+1.53000e-11'
+ mcm5m4l1_cf_w_0_300_s_0_600 = '-1.87500e-13*ic_cap*ic_cap+-1.00000e-13*ic_cap+1.97000e-11'
+ mcm5m4l1_cf_w_0_300_s_0_800 = '-2.43750e-13*ic_cap*ic_cap+-1.25000e-13*ic_cap+2.48000e-11'
+ mcm5m4l1_cf_w_0_300_s_1_000 = '-2.81250e-13*ic_cap*ic_cap+-1.50000e-13*ic_cap+2.92000e-11'
+ mcm5m4l1_cf_w_0_300_s_1_200 = '-3.12500e-13*ic_cap*ic_cap+-1.75000e-13*ic_cap+3.31000e-11'
+ mcm5m4l1_cf_w_0_300_s_2_100 = '-3.81250e-13*ic_cap*ic_cap+-2.25000e-13*ic_cap+4.48000e-11'
+ mcm5m4l1_cf_w_0_300_s_3_300 = '-3.84375e-13*ic_cap*ic_cap+-2.37500e-13*ic_cap+5.15000e-11'
+ mcm5m4l1_cf_w_0_300_s_9_000 = '-3.53125e-13*ic_cap*ic_cap+-2.12500e-13*ic_cap+5.59000e-11'
+ mcm5m4l1_cf_w_2_400_s_0_300 = '-7.78125e-14*ic_cap*ic_cap+-3.87500e-14*ic_cap+1.06000e-11'
+ mcm5m4l1_cf_w_2_400_s_0_360 = '-1.06250e-13*ic_cap*ic_cap+-5.00000e-14*ic_cap+1.26000e-11'
+ mcm5m4l1_cf_w_2_400_s_0_450 = '-1.40625e-13*ic_cap*ic_cap+-6.25000e-14*ic_cap+1.54000e-11'
+ mcm5m4l1_cf_w_2_400_s_0_600 = '-1.84375e-13*ic_cap*ic_cap+-8.75000e-14*ic_cap+1.97000e-11'
+ mcm5m4l1_cf_w_2_400_s_0_800 = '-2.37500e-13*ic_cap*ic_cap+-1.25000e-13*ic_cap+2.49000e-11'
+ mcm5m4l1_cf_w_2_400_s_1_000 = '-2.81250e-13*ic_cap*ic_cap+-1.50000e-13*ic_cap+2.95000e-11'
+ mcm5m4l1_cf_w_2_400_s_1_200 = '-3.09375e-13*ic_cap*ic_cap+-1.62500e-13*ic_cap+3.34000e-11'
+ mcm5m4l1_cf_w_2_400_s_2_100 = '-3.78125e-13*ic_cap*ic_cap+-2.12500e-13*ic_cap+4.56000e-11'
+ mcm5m4l1_cf_w_2_400_s_3_300 = '-3.71875e-13*ic_cap*ic_cap+-2.12500e-13*ic_cap+5.31000e-11'
+ mcm5m4l1_cf_w_2_400_s_9_000 = '-3.21875e-13*ic_cap*ic_cap+-1.87500e-13*ic_cap+5.84000e-11'
+ mcm5m4m1_ca_w_0_300_s_0_300 = '-1.22500e-06*ic_cap*ic_cap+-6.25000e-07*ic_cap+8.35000e-05'
+ mcm5m4m1_ca_w_0_300_s_0_360 = '-1.22500e-06*ic_cap*ic_cap+-6.25000e-07*ic_cap+8.35000e-05'
+ mcm5m4m1_ca_w_0_300_s_0_450 = '-1.22500e-06*ic_cap*ic_cap+-6.25000e-07*ic_cap+8.35000e-05'
+ mcm5m4m1_ca_w_0_300_s_0_600 = '-1.22500e-06*ic_cap*ic_cap+-6.25000e-07*ic_cap+8.35000e-05'
+ mcm5m4m1_ca_w_0_300_s_0_800 = '-1.22500e-06*ic_cap*ic_cap+-6.25000e-07*ic_cap+8.35000e-05'
+ mcm5m4m1_ca_w_0_300_s_1_000 = '-1.22500e-06*ic_cap*ic_cap+-6.25000e-07*ic_cap+8.35000e-05'
+ mcm5m4m1_ca_w_0_300_s_1_200 = '-1.22500e-06*ic_cap*ic_cap+-6.25000e-07*ic_cap+8.35000e-05'
+ mcm5m4m1_ca_w_0_300_s_2_100 = '-1.22500e-06*ic_cap*ic_cap+-6.25000e-07*ic_cap+8.35000e-05'
+ mcm5m4m1_ca_w_0_300_s_3_300 = '-1.22500e-06*ic_cap*ic_cap+-6.25000e-07*ic_cap+8.35000e-05'
+ mcm5m4m1_ca_w_0_300_s_9_000 = '-1.22500e-06*ic_cap*ic_cap+-6.25000e-07*ic_cap+8.35000e-05'
+ mcm5m4m1_ca_w_2_400_s_0_300 = '-1.22500e-06*ic_cap*ic_cap+-6.25000e-07*ic_cap+8.35000e-05'
+ mcm5m4m1_ca_w_2_400_s_0_360 = '-1.22500e-06*ic_cap*ic_cap+-6.25000e-07*ic_cap+8.35000e-05'
+ mcm5m4m1_ca_w_2_400_s_0_450 = '-1.22500e-06*ic_cap*ic_cap+-6.25000e-07*ic_cap+8.35000e-05'
+ mcm5m4m1_ca_w_2_400_s_0_600 = '-1.22500e-06*ic_cap*ic_cap+-6.25000e-07*ic_cap+8.35000e-05'
+ mcm5m4m1_ca_w_2_400_s_0_800 = '-1.22500e-06*ic_cap*ic_cap+-6.25000e-07*ic_cap+8.35000e-05'
+ mcm5m4m1_ca_w_2_400_s_1_000 = '-1.22500e-06*ic_cap*ic_cap+-6.25000e-07*ic_cap+8.35000e-05'
+ mcm5m4m1_ca_w_2_400_s_1_200 = '-1.22500e-06*ic_cap*ic_cap+-6.25000e-07*ic_cap+8.35000e-05'
+ mcm5m4m1_ca_w_2_400_s_2_100 = '-1.22500e-06*ic_cap*ic_cap+-6.25000e-07*ic_cap+8.35000e-05'
+ mcm5m4m1_ca_w_2_400_s_3_300 = '-1.22500e-06*ic_cap*ic_cap+-6.25000e-07*ic_cap+8.35000e-05'
+ mcm5m4m1_ca_w_2_400_s_9_000 = '-1.22500e-06*ic_cap*ic_cap+-6.25000e-07*ic_cap+8.35000e-05'
+ mcm5m4m1_cc_w_0_300_s_0_300 = '-6.09375e-13*ic_cap*ic_cap+-3.37500e-13*ic_cap+9.22000e-11'
+ mcm5m4m1_cc_w_0_300_s_0_360 = '-5.40625e-13*ic_cap*ic_cap+-3.37500e-13*ic_cap+8.45000e-11'
+ mcm5m4m1_cc_w_0_300_s_0_450 = '-4.18750e-13*ic_cap*ic_cap+-2.75000e-13*ic_cap+7.40000e-11'
+ mcm5m4m1_cc_w_0_300_s_0_600 = '-2.59375e-13*ic_cap*ic_cap+-1.87500e-13*ic_cap+5.97000e-11'
+ mcm5m4m1_cc_w_0_300_s_0_800 = '-1.40625e-13*ic_cap*ic_cap+-1.12500e-13*ic_cap+4.59000e-11'
+ mcm5m4m1_cc_w_0_300_s_1_000 = '-5.31250e-14*ic_cap*ic_cap+-6.25000e-14*ic_cap+3.56000e-11'
+ mcm5m4m1_cc_w_0_300_s_1_200 = '-6.25000e-15*ic_cap*ic_cap+-2.50000e-14*ic_cap+2.81000e-11'
+ mcm5m4m1_cc_w_0_300_s_2_100 = '5.31250e-14*ic_cap*ic_cap+1.25000e-14*ic_cap+1.10000e-11'
+ mcm5m4m1_cc_w_0_300_s_3_300 = '4.43750e-14*ic_cap*ic_cap+2.25000e-14*ic_cap+3.61000e-12'
+ mcm5m4m1_cc_w_0_300_s_9_000 = '2.34375e-15*ic_cap*ic_cap+3.12500e-15*ic_cap+5.50000e-14'
+ mcm5m4m1_cc_w_2_400_s_0_300 = '-5.28125e-13*ic_cap*ic_cap+-2.87500e-13*ic_cap+9.94000e-11'
+ mcm5m4m1_cc_w_2_400_s_0_360 = '-4.34375e-13*ic_cap*ic_cap+-2.62500e-13*ic_cap+9.08000e-11'
+ mcm5m4m1_cc_w_2_400_s_0_450 = '-3.15625e-13*ic_cap*ic_cap+-1.87500e-13*ic_cap+7.95000e-11'
+ mcm5m4m1_cc_w_2_400_s_0_600 = '-1.84375e-13*ic_cap*ic_cap+-1.12500e-13*ic_cap+6.45000e-11'
+ mcm5m4m1_cc_w_2_400_s_0_800 = '-6.87500e-14*ic_cap*ic_cap+-5.00000e-14*ic_cap+4.96000e-11'
+ mcm5m4m1_cc_w_2_400_s_1_000 = '-2.50000e-14*ic_cap+3.87000e-11'
+ mcm5m4m1_cc_w_2_400_s_1_200 = '4.37500e-14*ic_cap*ic_cap+3.07000e-11'
+ mcm5m4m1_cc_w_2_400_s_2_100 = '9.37500e-14*ic_cap*ic_cap+5.00000e-14*ic_cap+1.23000e-11'
+ mcm5m4m1_cc_w_2_400_s_3_300 = '5.81250e-14*ic_cap*ic_cap+4.25000e-14*ic_cap+4.21000e-12'
+ mcm5m4m1_cc_w_2_400_s_9_000 = '9.37500e-16*ic_cap*ic_cap+3.75000e-15*ic_cap+9.50000e-14'
+ mcm5m4m1_cf_w_0_300_s_0_300 = '-7.81250e-14*ic_cap*ic_cap+-3.75000e-14*ic_cap+1.10000e-11'
+ mcm5m4m1_cf_w_0_300_s_0_360 = '-1.06250e-13*ic_cap*ic_cap+-5.00000e-14*ic_cap+1.31000e-11'
+ mcm5m4m1_cf_w_0_300_s_0_450 = '-1.40625e-13*ic_cap*ic_cap+-6.25000e-14*ic_cap+1.60000e-11'
+ mcm5m4m1_cf_w_0_300_s_0_600 = '-1.90625e-13*ic_cap*ic_cap+-8.75000e-14*ic_cap+2.06000e-11'
+ mcm5m4m1_cf_w_0_300_s_0_800 = '-2.50000e-13*ic_cap*ic_cap+-1.25000e-13*ic_cap+2.60000e-11'
+ mcm5m4m1_cf_w_0_300_s_1_000 = '-2.93750e-13*ic_cap*ic_cap+-1.50000e-13*ic_cap+3.07000e-11'
+ mcm5m4m1_cf_w_0_300_s_1_200 = '-3.31250e-13*ic_cap*ic_cap+-1.75000e-13*ic_cap+3.48000e-11'
+ mcm5m4m1_cf_w_0_300_s_2_100 = '-3.93750e-13*ic_cap*ic_cap+-2.25000e-13*ic_cap+4.66000e-11'
+ mcm5m4m1_cf_w_0_300_s_3_300 = '-3.90625e-13*ic_cap*ic_cap+-2.37500e-13*ic_cap+5.31000e-11'
+ mcm5m4m1_cf_w_0_300_s_9_000 = '-3.62500e-13*ic_cap*ic_cap+-2.00000e-13*ic_cap+5.67000e-11'
+ mcm5m4m1_cf_w_2_400_s_0_300 = '-7.93750e-14*ic_cap*ic_cap+-3.75000e-14*ic_cap+1.11000e-11'
+ mcm5m4m1_cf_w_2_400_s_0_360 = '-1.00000e-13*ic_cap*ic_cap+-5.00000e-14*ic_cap+1.31000e-11'
+ mcm5m4m1_cf_w_2_400_s_0_450 = '-1.40625e-13*ic_cap*ic_cap+-6.25000e-14*ic_cap+1.61000e-11'
+ mcm5m4m1_cf_w_2_400_s_0_600 = '-1.93750e-13*ic_cap*ic_cap+-1.00000e-13*ic_cap+2.07000e-11'
+ mcm5m4m1_cf_w_2_400_s_0_800 = '-2.46875e-13*ic_cap*ic_cap+-1.37500e-13*ic_cap+2.61000e-11'
+ mcm5m4m1_cf_w_2_400_s_1_000 = '-2.90625e-13*ic_cap*ic_cap+-1.62500e-13*ic_cap+3.09000e-11'
+ mcm5m4m1_cf_w_2_400_s_1_200 = '-3.21875e-13*ic_cap*ic_cap+-1.87500e-13*ic_cap+3.50000e-11'
+ mcm5m4m1_cf_w_2_400_s_2_100 = '-3.81250e-13*ic_cap*ic_cap+-2.25000e-13*ic_cap+4.74000e-11'
+ mcm5m4m1_cf_w_2_400_s_3_300 = '-3.71875e-13*ic_cap*ic_cap+-2.12500e-13*ic_cap+5.45000e-11'
+ mcm5m4m1_cf_w_2_400_s_9_000 = '-3.21875e-13*ic_cap*ic_cap+-1.87500e-13*ic_cap+5.86000e-11'
+ mcm5m4m2_ca_w_0_300_s_0_300 = '-1.26563e-06*ic_cap*ic_cap+-6.37500e-07*ic_cap+8.92000e-05'
+ mcm5m4m2_ca_w_0_300_s_0_360 = '-1.26563e-06*ic_cap*ic_cap+-6.37500e-07*ic_cap+8.92000e-05'
+ mcm5m4m2_ca_w_0_300_s_0_450 = '-1.26563e-06*ic_cap*ic_cap+-6.37500e-07*ic_cap+8.92000e-05'
+ mcm5m4m2_ca_w_0_300_s_0_600 = '-1.26563e-06*ic_cap*ic_cap+-6.37500e-07*ic_cap+8.92000e-05'
+ mcm5m4m2_ca_w_0_300_s_0_800 = '-1.26563e-06*ic_cap*ic_cap+-6.37500e-07*ic_cap+8.92000e-05'
+ mcm5m4m2_ca_w_0_300_s_1_000 = '-1.26563e-06*ic_cap*ic_cap+-6.37500e-07*ic_cap+8.92000e-05'
+ mcm5m4m2_ca_w_0_300_s_1_200 = '-1.26563e-06*ic_cap*ic_cap+-6.37500e-07*ic_cap+8.92000e-05'
+ mcm5m4m2_ca_w_0_300_s_2_100 = '-1.26563e-06*ic_cap*ic_cap+-6.37500e-07*ic_cap+8.92000e-05'
+ mcm5m4m2_ca_w_0_300_s_3_300 = '-1.26563e-06*ic_cap*ic_cap+-6.37500e-07*ic_cap+8.92000e-05'
+ mcm5m4m2_ca_w_0_300_s_9_000 = '-1.26563e-06*ic_cap*ic_cap+-6.37500e-07*ic_cap+8.92000e-05'
+ mcm5m4m2_ca_w_2_400_s_0_300 = '-1.26563e-06*ic_cap*ic_cap+-6.37500e-07*ic_cap+8.92000e-05'
+ mcm5m4m2_ca_w_2_400_s_0_360 = '-1.26563e-06*ic_cap*ic_cap+-6.37500e-07*ic_cap+8.92000e-05'
+ mcm5m4m2_ca_w_2_400_s_0_450 = '-1.26563e-06*ic_cap*ic_cap+-6.37500e-07*ic_cap+8.92000e-05'
+ mcm5m4m2_ca_w_2_400_s_0_600 = '-1.26563e-06*ic_cap*ic_cap+-6.37500e-07*ic_cap+8.92000e-05'
+ mcm5m4m2_ca_w_2_400_s_0_800 = '-1.26563e-06*ic_cap*ic_cap+-6.37500e-07*ic_cap+8.92000e-05'
+ mcm5m4m2_ca_w_2_400_s_1_000 = '-1.26563e-06*ic_cap*ic_cap+-6.37500e-07*ic_cap+8.92000e-05'
+ mcm5m4m2_ca_w_2_400_s_1_200 = '-1.26563e-06*ic_cap*ic_cap+-6.37500e-07*ic_cap+8.92000e-05'
+ mcm5m4m2_ca_w_2_400_s_2_100 = '-1.26563e-06*ic_cap*ic_cap+-6.37500e-07*ic_cap+8.92000e-05'
+ mcm5m4m2_ca_w_2_400_s_3_300 = '-1.26563e-06*ic_cap*ic_cap+-6.37500e-07*ic_cap+8.92000e-05'
+ mcm5m4m2_ca_w_2_400_s_9_000 = '-1.26563e-06*ic_cap*ic_cap+-6.37500e-07*ic_cap+8.92000e-05'
+ mcm5m4m2_cc_w_0_300_s_0_300 = '-6.15625e-13*ic_cap*ic_cap+-3.37500e-13*ic_cap+9.10000e-11'
+ mcm5m4m2_cc_w_0_300_s_0_360 = '-5.31250e-13*ic_cap*ic_cap+-3.25000e-13*ic_cap+8.30000e-11'
+ mcm5m4m2_cc_w_0_300_s_0_450 = '-4.12500e-13*ic_cap*ic_cap+-2.75000e-13*ic_cap+7.24000e-11'
+ mcm5m4m2_cc_w_0_300_s_0_600 = '-2.46875e-13*ic_cap*ic_cap+-1.62500e-13*ic_cap+5.78000e-11'
+ mcm5m4m2_cc_w_0_300_s_0_800 = '-1.28125e-13*ic_cap*ic_cap+-1.12500e-13*ic_cap+4.38000e-11'
+ mcm5m4m2_cc_w_0_300_s_1_000 = '-5.00000e-14*ic_cap*ic_cap+-5.00000e-14*ic_cap+3.35000e-11'
+ mcm5m4m2_cc_w_0_300_s_1_200 = '2.01948e-28*ic_cap*ic_cap+-2.50000e-14*ic_cap+2.59000e-11'
+ mcm5m4m2_cc_w_0_300_s_2_100 = '5.56250e-14*ic_cap*ic_cap+2.25000e-14*ic_cap+9.12000e-12'
+ mcm5m4m2_cc_w_0_300_s_3_300 = '3.68750e-14*ic_cap*ic_cap+2.50000e-14*ic_cap+2.55000e-12'
+ mcm5m4m2_cc_w_0_300_s_9_000 = '1.25000e-15*ic_cap+4.00000e-14'
+ mcm5m4m2_cc_w_2_400_s_0_300 = '-5.28125e-13*ic_cap*ic_cap+-2.87500e-13*ic_cap+9.61000e-11'
+ mcm5m4m2_cc_w_2_400_s_0_360 = '-4.46875e-13*ic_cap*ic_cap+-2.62500e-13*ic_cap+8.77000e-11'
+ mcm5m4m2_cc_w_2_400_s_0_450 = '-3.21875e-13*ic_cap*ic_cap+-1.87500e-13*ic_cap+7.62000e-11'
+ mcm5m4m2_cc_w_2_400_s_0_600 = '-1.87500e-13*ic_cap*ic_cap+-1.25000e-13*ic_cap+6.12000e-11'
+ mcm5m4m2_cc_w_2_400_s_0_800 = '-6.87500e-14*ic_cap*ic_cap+-7.50000e-14*ic_cap+4.63000e-11'
+ mcm5m4m2_cc_w_2_400_s_1_000 = '-2.50000e-14*ic_cap+3.54000e-11'
+ mcm5m4m2_cc_w_2_400_s_1_200 = '4.06250e-14*ic_cap*ic_cap+1.25000e-14*ic_cap+2.75000e-11'
+ mcm5m4m2_cc_w_2_400_s_2_100 = '7.50000e-14*ic_cap*ic_cap+3.75000e-14*ic_cap+9.85000e-12'
+ mcm5m4m2_cc_w_2_400_s_3_300 = '4.65625e-14*ic_cap*ic_cap+3.12500e-14*ic_cap+2.76000e-12'
+ mcm5m4m2_cc_w_2_400_s_9_000 = '2.65625e-15*ic_cap*ic_cap+-6.25000e-16*ic_cap+5.00000e-15'
+ mcm5m4m2_cf_w_0_300_s_0_300 = '-8.43750e-14*ic_cap*ic_cap+-3.75000e-14*ic_cap+1.19000e-11'
+ mcm5m4m2_cf_w_0_300_s_0_360 = '-1.09375e-13*ic_cap*ic_cap+-6.25000e-14*ic_cap+1.41000e-11'
+ mcm5m4m2_cf_w_0_300_s_0_450 = '-1.50000e-13*ic_cap*ic_cap+-7.50000e-14*ic_cap+1.73000e-11'
+ mcm5m4m2_cf_w_0_300_s_0_600 = '-2.00000e-13*ic_cap*ic_cap+-1.00000e-13*ic_cap+2.22000e-11'
+ mcm5m4m2_cf_w_0_300_s_0_800 = '-2.56250e-13*ic_cap*ic_cap+-1.25000e-13*ic_cap+2.79000e-11'
+ mcm5m4m2_cf_w_0_300_s_1_000 = '-3.03125e-13*ic_cap*ic_cap+-1.62500e-13*ic_cap+3.30000e-11'
+ mcm5m4m2_cf_w_0_300_s_1_200 = '-3.40625e-13*ic_cap*ic_cap+-1.87500e-13*ic_cap+3.73000e-11'
+ mcm5m4m2_cf_w_0_300_s_2_100 = '-4.03125e-13*ic_cap*ic_cap+-2.37500e-13*ic_cap+4.94000e-11'
+ mcm5m4m2_cf_w_0_300_s_3_300 = '-3.96875e-13*ic_cap*ic_cap+-2.37500e-13*ic_cap+5.55000e-11'
+ mcm5m4m2_cf_w_0_300_s_9_000 = '-3.65625e-13*ic_cap*ic_cap+-2.12500e-13*ic_cap+5.80000e-11'
+ mcm5m4m2_cf_w_2_400_s_0_300 = '-7.81250e-14*ic_cap*ic_cap+-3.75000e-14*ic_cap+1.19000e-11'
+ mcm5m4m2_cf_w_2_400_s_0_360 = '-1.06250e-13*ic_cap*ic_cap+-5.00000e-14*ic_cap+1.41000e-11'
+ mcm5m4m2_cf_w_2_400_s_0_450 = '-1.43750e-13*ic_cap*ic_cap+-7.50000e-14*ic_cap+1.73000e-11'
+ mcm5m4m2_cf_w_2_400_s_0_600 = '-1.93750e-13*ic_cap*ic_cap+-1.00000e-13*ic_cap+2.22000e-11'
+ mcm5m4m2_cf_w_2_400_s_0_800 = '-2.53125e-13*ic_cap*ic_cap+-1.37500e-13*ic_cap+2.81000e-11'
+ mcm5m4m2_cf_w_2_400_s_1_000 = '-2.96875e-13*ic_cap*ic_cap+-1.62500e-13*ic_cap+3.32000e-11'
+ mcm5m4m2_cf_w_2_400_s_1_200 = '-3.34375e-13*ic_cap*ic_cap+-1.87500e-13*ic_cap+3.76000e-11'
+ mcm5m4m2_cf_w_2_400_s_2_100 = '-3.93750e-13*ic_cap*ic_cap+-2.25000e-13*ic_cap+5.03000e-11'
+ mcm5m4m2_cf_w_2_400_s_3_300 = '-3.75000e-13*ic_cap*ic_cap+-2.25000e-13*ic_cap+5.66000e-11'
+ mcm5m4m2_cf_w_2_400_s_9_000 = '-3.34375e-13*ic_cap*ic_cap+-1.87500e-13*ic_cap+5.94000e-11'
+ mcm5m4m3_ca_w_0_300_s_0_300 = '-2.84375e-06*ic_cap*ic_cap+-1.37500e-06*ic_cap+1.57000e-04'
+ mcm5m4m3_ca_w_0_300_s_0_360 = '-2.84375e-06*ic_cap*ic_cap+-1.37500e-06*ic_cap+1.57000e-04'
+ mcm5m4m3_ca_w_0_300_s_0_450 = '-2.84375e-06*ic_cap*ic_cap+-1.37500e-06*ic_cap+1.57000e-04'
+ mcm5m4m3_ca_w_0_300_s_0_600 = '-2.84375e-06*ic_cap*ic_cap+-1.37500e-06*ic_cap+1.57000e-04'
+ mcm5m4m3_ca_w_0_300_s_0_800 = '-2.84375e-06*ic_cap*ic_cap+-1.37500e-06*ic_cap+1.57000e-04'
+ mcm5m4m3_ca_w_0_300_s_1_000 = '-2.84375e-06*ic_cap*ic_cap+-1.37500e-06*ic_cap+1.57000e-04'
+ mcm5m4m3_ca_w_0_300_s_1_200 = '-2.84375e-06*ic_cap*ic_cap+-1.37500e-06*ic_cap+1.57000e-04'
+ mcm5m4m3_ca_w_0_300_s_2_100 = '-2.84375e-06*ic_cap*ic_cap+-1.37500e-06*ic_cap+1.57000e-04'
+ mcm5m4m3_ca_w_0_300_s_3_300 = '-2.84375e-06*ic_cap*ic_cap+-1.37500e-06*ic_cap+1.57000e-04'
+ mcm5m4m3_ca_w_0_300_s_9_000 = '-2.84375e-06*ic_cap*ic_cap+-1.37500e-06*ic_cap+1.57000e-04'
+ mcm5m4m3_ca_w_2_400_s_0_300 = '-2.84375e-06*ic_cap*ic_cap+-1.37500e-06*ic_cap+1.57000e-04'
+ mcm5m4m3_ca_w_2_400_s_0_360 = '-2.84375e-06*ic_cap*ic_cap+-1.37500e-06*ic_cap+1.57000e-04'
+ mcm5m4m3_ca_w_2_400_s_0_450 = '-2.84375e-06*ic_cap*ic_cap+-1.37500e-06*ic_cap+1.57000e-04'
+ mcm5m4m3_ca_w_2_400_s_0_600 = '-2.84375e-06*ic_cap*ic_cap+-1.37500e-06*ic_cap+1.57000e-04'
+ mcm5m4m3_ca_w_2_400_s_0_800 = '-2.84375e-06*ic_cap*ic_cap+-1.37500e-06*ic_cap+1.57000e-04'
+ mcm5m4m3_ca_w_2_400_s_1_000 = '-2.84375e-06*ic_cap*ic_cap+-1.37500e-06*ic_cap+1.57000e-04'
+ mcm5m4m3_ca_w_2_400_s_1_200 = '-2.84375e-06*ic_cap*ic_cap+-1.37500e-06*ic_cap+1.57000e-04'
+ mcm5m4m3_ca_w_2_400_s_2_100 = '-2.84375e-06*ic_cap*ic_cap+-1.37500e-06*ic_cap+1.57000e-04'
+ mcm5m4m3_ca_w_2_400_s_3_300 = '-2.84375e-06*ic_cap*ic_cap+-1.37500e-06*ic_cap+1.57000e-04'
+ mcm5m4m3_ca_w_2_400_s_9_000 = '-2.84375e-06*ic_cap*ic_cap+-1.37500e-06*ic_cap+1.57000e-04'
+ mcm5m4m3_cc_w_0_300_s_0_300 = '-4.15625e-13*ic_cap*ic_cap+-2.37500e-13*ic_cap+7.96000e-11'
+ mcm5m4m3_cc_w_0_300_s_0_360 = '-3.12500e-13*ic_cap*ic_cap+-2.00000e-13*ic_cap+7.11000e-11'
+ mcm5m4m3_cc_w_0_300_s_0_450 = '-2.15625e-13*ic_cap*ic_cap+-1.37500e-13*ic_cap+6.04000e-11'
+ mcm5m4m3_cc_w_0_300_s_0_600 = '-7.81250e-14*ic_cap*ic_cap+-8.75000e-14*ic_cap+4.57000e-11'
+ mcm5m4m3_cc_w_0_300_s_0_800 = '3.12500e-14*ic_cap*ic_cap+3.16000e-11'
+ mcm5m4m3_cc_w_0_300_s_1_000 = '9.06250e-14*ic_cap*ic_cap+3.75000e-14*ic_cap+2.17000e-11'
+ mcm5m4m3_cc_w_0_300_s_1_200 = '1.15625e-13*ic_cap*ic_cap+6.25000e-14*ic_cap+1.49000e-11'
+ mcm5m4m3_cc_w_0_300_s_2_100 = '7.28125e-14*ic_cap*ic_cap+4.37500e-14*ic_cap+2.94000e-12'
+ mcm5m4m3_cc_w_0_300_s_3_300 = '1.54688e-14*ic_cap*ic_cap+1.18750e-14*ic_cap+4.25000e-13'
+ mcm5m4m3_cc_w_0_300_s_9_000 = '1.40625e-15*ic_cap*ic_cap+5.62500e-15*ic_cap'
+ mcm5m4m3_cc_w_2_400_s_0_300 = '-3.62500e-13*ic_cap*ic_cap+-2.25000e-13*ic_cap+8.05000e-11'
+ mcm5m4m3_cc_w_2_400_s_0_360 = '-2.78125e-13*ic_cap*ic_cap+-1.87500e-13*ic_cap+7.21000e-11'
+ mcm5m4m3_cc_w_2_400_s_0_450 = '-1.59375e-13*ic_cap*ic_cap+-1.37500e-13*ic_cap+6.07000e-11'
+ mcm5m4m3_cc_w_2_400_s_0_600 = '-5.00000e-14*ic_cap*ic_cap+-5.00000e-14*ic_cap+4.63000e-11'
+ mcm5m4m3_cc_w_2_400_s_0_800 = '6.25000e-14*ic_cap*ic_cap+2.50000e-14*ic_cap+3.18000e-11'
+ mcm5m4m3_cc_w_2_400_s_1_000 = '1.12500e-13*ic_cap*ic_cap+5.00000e-14*ic_cap+2.19000e-11'
+ mcm5m4m3_cc_w_2_400_s_1_200 = '1.34375e-13*ic_cap*ic_cap+6.25000e-14*ic_cap+1.50000e-11'
+ mcm5m4m3_cc_w_2_400_s_2_100 = '7.96875e-14*ic_cap*ic_cap+5.62500e-14*ic_cap+2.95000e-12'
+ mcm5m4m3_cc_w_2_400_s_3_300 = '2.03125e-14*ic_cap*ic_cap+6.25000e-15*ic_cap+4.00000e-13'
+ mcm5m4m3_cf_w_0_300_s_0_300 = '-2.28125e-13*ic_cap*ic_cap+-1.12500e-13*ic_cap+2.07000e-11'
+ mcm5m4m3_cf_w_0_300_s_0_360 = '-2.84375e-13*ic_cap*ic_cap+-1.37500e-13*ic_cap+2.43000e-11'
+ mcm5m4m3_cf_w_0_300_s_0_450 = '-3.62500e-13*ic_cap*ic_cap+-1.75000e-13*ic_cap+2.95000e-11'
+ mcm5m4m3_cf_w_0_300_s_0_600 = '-4.68750e-13*ic_cap*ic_cap+-2.50000e-13*ic_cap+3.72000e-11'
+ mcm5m4m3_cf_w_0_300_s_0_800 = '-5.71875e-13*ic_cap*ic_cap+-2.87500e-13*ic_cap+4.58000e-11'
+ mcm5m4m3_cf_w_0_300_s_1_000 = '-6.53125e-13*ic_cap*ic_cap+-3.37500e-13*ic_cap+5.29000e-11'
+ mcm5m4m3_cf_w_0_300_s_1_200 = '-6.96875e-13*ic_cap*ic_cap+-3.62500e-13*ic_cap+5.81000e-11'
+ mcm5m4m3_cf_w_0_300_s_2_100 = '-6.87500e-13*ic_cap*ic_cap+-3.75000e-13*ic_cap+6.87000e-11'
+ mcm5m4m3_cf_w_0_300_s_3_300 = '-6.31250e-13*ic_cap*ic_cap+-3.50000e-13*ic_cap+7.12000e-11'
+ mcm5m4m3_cf_w_0_300_s_9_000 = '-6.12500e-13*ic_cap*ic_cap+-3.25000e-13*ic_cap+7.16000e-11'
+ mcm5m4m3_cf_w_2_400_s_0_300 = '-2.21875e-13*ic_cap*ic_cap+-1.12500e-13*ic_cap+2.07000e-11'
+ mcm5m4m3_cf_w_2_400_s_0_360 = '-2.81250e-13*ic_cap*ic_cap+-1.50000e-13*ic_cap+2.44000e-11'
+ mcm5m4m3_cf_w_2_400_s_0_450 = '-3.53125e-13*ic_cap*ic_cap+-1.87500e-13*ic_cap+2.95000e-11'
+ mcm5m4m3_cf_w_2_400_s_0_600 = '-4.59375e-13*ic_cap*ic_cap+-2.37500e-13*ic_cap+3.72000e-11'
+ mcm5m4m3_cf_w_2_400_s_0_800 = '-5.71875e-13*ic_cap*ic_cap+-2.87500e-13*ic_cap+4.60000e-11'
+ mcm5m4m3_cf_w_2_400_s_1_000 = '-6.28125e-13*ic_cap*ic_cap+-3.37500e-13*ic_cap+5.28000e-11'
+ mcm5m4m3_cf_w_2_400_s_1_200 = '-6.71875e-13*ic_cap*ic_cap+-3.62500e-13*ic_cap+5.81000e-11'
+ mcm5m4m3_cf_w_2_400_s_2_100 = '-6.68750e-13*ic_cap*ic_cap+-3.75000e-13*ic_cap+6.90000e-11'
+ mcm5m4m3_cf_w_2_400_s_3_300 = '-6.15625e-13*ic_cap*ic_cap+-3.37500e-13*ic_cap+7.16000e-11'
+ mcm5m4m3_cf_w_2_400_s_9_000 = '-6.00000e-13*ic_cap*ic_cap+-3.25000e-13*ic_cap+7.21000e-11'
+ mcm5m4p1_ca_w_0_300_s_0_300 = '-1.18750e-06*ic_cap*ic_cap+-6.00000e-07*ic_cap+7.85000e-05'
+ mcm5m4p1_ca_w_0_300_s_0_360 = '-1.18750e-06*ic_cap*ic_cap+-6.00000e-07*ic_cap+7.85000e-05'
+ mcm5m4p1_ca_w_0_300_s_0_450 = '-1.18750e-06*ic_cap*ic_cap+-6.00000e-07*ic_cap+7.85000e-05'
+ mcm5m4p1_ca_w_0_300_s_0_600 = '-1.18750e-06*ic_cap*ic_cap+-6.00000e-07*ic_cap+7.85000e-05'
+ mcm5m4p1_ca_w_0_300_s_0_800 = '-1.18750e-06*ic_cap*ic_cap+-6.00000e-07*ic_cap+7.85000e-05'
+ mcm5m4p1_ca_w_0_300_s_1_000 = '-1.18750e-06*ic_cap*ic_cap+-6.00000e-07*ic_cap+7.85000e-05'
+ mcm5m4p1_ca_w_0_300_s_1_200 = '-1.18750e-06*ic_cap*ic_cap+-6.00000e-07*ic_cap+7.85000e-05'
+ mcm5m4p1_ca_w_0_300_s_2_100 = '-1.18750e-06*ic_cap*ic_cap+-6.00000e-07*ic_cap+7.85000e-05'
+ mcm5m4p1_ca_w_0_300_s_3_300 = '-1.18750e-06*ic_cap*ic_cap+-6.00000e-07*ic_cap+7.85000e-05'
+ mcm5m4p1_ca_w_0_300_s_9_000 = '-1.18750e-06*ic_cap*ic_cap+-6.00000e-07*ic_cap+7.85000e-05'
+ mcm5m4p1_ca_w_2_400_s_0_300 = '-1.18750e-06*ic_cap*ic_cap+-6.00000e-07*ic_cap+7.85000e-05'
+ mcm5m4p1_ca_w_2_400_s_0_360 = '-1.18750e-06*ic_cap*ic_cap+-6.00000e-07*ic_cap+7.85000e-05'
+ mcm5m4p1_ca_w_2_400_s_0_450 = '-1.18750e-06*ic_cap*ic_cap+-6.00000e-07*ic_cap+7.85000e-05'
+ mcm5m4p1_ca_w_2_400_s_0_600 = '-1.18750e-06*ic_cap*ic_cap+-6.00000e-07*ic_cap+7.85000e-05'
+ mcm5m4p1_ca_w_2_400_s_0_800 = '-1.18750e-06*ic_cap*ic_cap+-6.00000e-07*ic_cap+7.85000e-05'
+ mcm5m4p1_ca_w_2_400_s_1_000 = '-1.18750e-06*ic_cap*ic_cap+-6.00000e-07*ic_cap+7.85000e-05'
+ mcm5m4p1_ca_w_2_400_s_1_200 = '-1.18750e-06*ic_cap*ic_cap+-6.00000e-07*ic_cap+7.85000e-05'
+ mcm5m4p1_ca_w_2_400_s_2_100 = '-1.18750e-06*ic_cap*ic_cap+-6.00000e-07*ic_cap+7.85000e-05'
+ mcm5m4p1_ca_w_2_400_s_3_300 = '-1.18750e-06*ic_cap*ic_cap+-6.00000e-07*ic_cap+7.85000e-05'
+ mcm5m4p1_ca_w_2_400_s_9_000 = '-1.18750e-06*ic_cap*ic_cap+-6.00000e-07*ic_cap+7.85000e-05'
+ mcm5m4p1_cc_w_0_300_s_0_300 = '-6.21875e-13*ic_cap*ic_cap+-3.62500e-13*ic_cap+9.34000e-11'
+ mcm5m4p1_cc_w_0_300_s_0_360 = '-5.50000e-13*ic_cap*ic_cap+-3.25000e-13*ic_cap+8.59000e-11'
+ mcm5m4p1_cc_w_0_300_s_0_450 = '-4.25000e-13*ic_cap*ic_cap+-2.75000e-13*ic_cap+7.54000e-11'
+ mcm5m4p1_cc_w_0_300_s_0_600 = '-2.81250e-13*ic_cap*ic_cap+-1.75000e-13*ic_cap+6.15000e-11'
+ mcm5m4p1_cc_w_0_300_s_0_800 = '-1.59375e-13*ic_cap*ic_cap+-1.12500e-13*ic_cap+4.79000e-11'
+ mcm5m4p1_cc_w_0_300_s_1_000 = '-6.56250e-14*ic_cap*ic_cap+-8.75000e-14*ic_cap+3.78000e-11'
+ mcm5m4p1_cc_w_0_300_s_1_200 = '-2.18750e-14*ic_cap*ic_cap+-3.75000e-14*ic_cap+3.04000e-11'
+ mcm5m4p1_cc_w_0_300_s_2_100 = '4.06250e-14*ic_cap*ic_cap+1.25000e-14*ic_cap+1.32000e-11'
+ mcm5m4p1_cc_w_0_300_s_3_300 = '4.68750e-14*ic_cap*ic_cap+2.75000e-14*ic_cap+5.10000e-12'
+ mcm5m4p1_cc_w_0_300_s_9_000 = '4.68750e-15*ic_cap*ic_cap+6.25000e-15*ic_cap+1.45000e-13'
+ mcm5m4p1_cc_w_2_400_s_0_300 = '-5.31250e-13*ic_cap*ic_cap+-3.25000e-13*ic_cap+1.03000e-10'
+ mcm5m4p1_cc_w_2_400_s_0_360 = '-4.43750e-13*ic_cap*ic_cap+-2.50000e-13*ic_cap+9.46000e-11'
+ mcm5m4p1_cc_w_2_400_s_0_450 = '-3.25000e-13*ic_cap*ic_cap+-2.00000e-13*ic_cap+8.33000e-11'
+ mcm5m4p1_cc_w_2_400_s_0_600 = '-1.90625e-13*ic_cap*ic_cap+-1.37500e-13*ic_cap+6.83000e-11'
+ mcm5m4p1_cc_w_2_400_s_0_800 = '-8.12500e-14*ic_cap*ic_cap+-5.00000e-14*ic_cap+5.35000e-11'
+ mcm5m4p1_cc_w_2_400_s_1_000 = '-6.25000e-15*ic_cap*ic_cap+-2.50000e-14*ic_cap+4.26000e-11'
+ mcm5m4p1_cc_w_2_400_s_1_200 = '4.06250e-14*ic_cap*ic_cap+1.25000e-14*ic_cap+3.45000e-11'
+ mcm5m4p1_cc_w_2_400_s_2_100 = '8.75000e-14*ic_cap*ic_cap+5.00000e-14*ic_cap+1.57000e-11'
+ mcm5m4p1_cc_w_2_400_s_3_300 = '7.25000e-14*ic_cap*ic_cap+4.50000e-14*ic_cap+6.43000e-12'
+ mcm5m4p1_cc_w_2_400_s_9_000 = '8.59375e-15*ic_cap*ic_cap+1.31250e-14*ic_cap+1.70000e-13'
+ mcm5m4p1_cf_w_0_300_s_0_300 = '-7.96875e-14*ic_cap*ic_cap+-3.87500e-14*ic_cap+1.03000e-11'
+ mcm5m4p1_cf_w_0_300_s_0_360 = '-1.06250e-13*ic_cap*ic_cap+-5.00000e-14*ic_cap+1.22000e-11'
+ mcm5m4p1_cf_w_0_300_s_0_450 = '-1.40625e-13*ic_cap*ic_cap+-6.25000e-14*ic_cap+1.50000e-11'
+ mcm5m4p1_cf_w_0_300_s_0_600 = '-1.84375e-13*ic_cap*ic_cap+-8.75000e-14*ic_cap+1.92000e-11'
+ mcm5m4p1_cf_w_0_300_s_0_800 = '-2.43750e-13*ic_cap*ic_cap+-1.25000e-13*ic_cap+2.42000e-11'
+ mcm5m4p1_cf_w_0_300_s_1_000 = '-2.84375e-13*ic_cap*ic_cap+-1.62500e-13*ic_cap+2.86000e-11'
+ mcm5m4p1_cf_w_0_300_s_1_200 = '-3.18750e-13*ic_cap*ic_cap+-1.75000e-13*ic_cap+3.24000e-11'
+ mcm5m4p1_cf_w_0_300_s_2_100 = '-3.84375e-13*ic_cap*ic_cap+-2.12500e-13*ic_cap+4.40000e-11'
+ mcm5m4p1_cf_w_0_300_s_3_300 = '-3.90625e-13*ic_cap*ic_cap+-2.37500e-13*ic_cap+5.08000e-11'
+ mcm5m4p1_cf_w_0_300_s_9_000 = '-3.56250e-13*ic_cap*ic_cap+-2.00000e-13*ic_cap+5.56000e-11'
+ mcm5m4p1_cf_w_2_400_s_0_300 = '-8.03125e-14*ic_cap*ic_cap+-3.87500e-14*ic_cap+1.04000e-11'
+ mcm5m4p1_cf_w_2_400_s_0_360 = '-1.06250e-13*ic_cap*ic_cap+-5.00000e-14*ic_cap+1.23000e-11'
+ mcm5m4p1_cf_w_2_400_s_0_450 = '-1.37500e-13*ic_cap*ic_cap+-7.50000e-14*ic_cap+1.50000e-11'
+ mcm5m4p1_cf_w_2_400_s_0_600 = '-1.87500e-13*ic_cap*ic_cap+-1.00000e-13*ic_cap+1.93000e-11'
+ mcm5m4p1_cf_w_2_400_s_0_800 = '-2.43750e-13*ic_cap*ic_cap+-1.25000e-13*ic_cap+2.44000e-11'
+ mcm5m4p1_cf_w_2_400_s_1_000 = '-2.81250e-13*ic_cap*ic_cap+-1.50000e-13*ic_cap+2.88000e-11'
+ mcm5m4p1_cf_w_2_400_s_1_200 = '-3.09375e-13*ic_cap*ic_cap+-1.62500e-13*ic_cap+3.26000e-11'
+ mcm5m4p1_cf_w_2_400_s_2_100 = '-3.78125e-13*ic_cap*ic_cap+-2.12500e-13*ic_cap+4.47000e-11'
+ mcm5m4p1_cf_w_2_400_s_3_300 = '-3.78125e-13*ic_cap*ic_cap+-2.12500e-13*ic_cap+5.24000e-11'
+ mcm5m4p1_cf_w_2_400_s_9_000 = '-3.21875e-13*ic_cap*ic_cap+-1.87500e-13*ic_cap+5.84000e-11'
+ mcm5p1_ca_w_1_600_s_10_000 = '-5.71875e-08*ic_cap*ic_cap+-3.62500e-08*ic_cap+7.26000e-06'
+ mcm5p1_ca_w_1_600_s_12_000 = '-5.71875e-08*ic_cap*ic_cap+-3.62500e-08*ic_cap+7.26000e-06'
+ mcm5p1_ca_w_1_600_s_1_600 = '-5.71875e-08*ic_cap*ic_cap+-3.62500e-08*ic_cap+7.26000e-06'
+ mcm5p1_ca_w_1_600_s_1_700 = '-5.71875e-08*ic_cap*ic_cap+-3.62500e-08*ic_cap+7.26000e-06'
+ mcm5p1_ca_w_1_600_s_1_900 = '-5.71875e-08*ic_cap*ic_cap+-3.62500e-08*ic_cap+7.26000e-06'
+ mcm5p1_ca_w_1_600_s_2_000 = '-5.71875e-08*ic_cap*ic_cap+-3.62500e-08*ic_cap+7.26000e-06'
+ mcm5p1_ca_w_1_600_s_2_400 = '-5.71875e-08*ic_cap*ic_cap+-3.62500e-08*ic_cap+7.26000e-06'
+ mcm5p1_ca_w_1_600_s_2_800 = '-5.71875e-08*ic_cap*ic_cap+-3.62500e-08*ic_cap+7.26000e-06'
+ mcm5p1_ca_w_1_600_s_3_200 = '-5.71875e-08*ic_cap*ic_cap+-3.62500e-08*ic_cap+7.26000e-06'
+ mcm5p1_ca_w_1_600_s_4_800 = '-5.71875e-08*ic_cap*ic_cap+-3.62500e-08*ic_cap+7.26000e-06'
+ mcm5p1_ca_w_4_000_s_10_000 = '-5.71875e-08*ic_cap*ic_cap+-3.62500e-08*ic_cap+7.26000e-06'
+ mcm5p1_ca_w_4_000_s_12_000 = '-5.71875e-08*ic_cap*ic_cap+-3.62500e-08*ic_cap+7.26000e-06'
+ mcm5p1_ca_w_4_000_s_1_600 = '-5.71875e-08*ic_cap*ic_cap+-3.62500e-08*ic_cap+7.26000e-06'
+ mcm5p1_ca_w_4_000_s_1_700 = '-5.71875e-08*ic_cap*ic_cap+-3.62500e-08*ic_cap+7.26000e-06'
+ mcm5p1_ca_w_4_000_s_1_900 = '-5.71875e-08*ic_cap*ic_cap+-3.62500e-08*ic_cap+7.26000e-06'
+ mcm5p1_ca_w_4_000_s_2_000 = '-5.71875e-08*ic_cap*ic_cap+-3.62500e-08*ic_cap+7.26000e-06'
+ mcm5p1_ca_w_4_000_s_2_400 = '-5.71875e-08*ic_cap*ic_cap+-3.62500e-08*ic_cap+7.26000e-06'
+ mcm5p1_ca_w_4_000_s_2_800 = '-5.71875e-08*ic_cap*ic_cap+-3.62500e-08*ic_cap+7.26000e-06'
+ mcm5p1_ca_w_4_000_s_3_200 = '-5.71875e-08*ic_cap*ic_cap+-3.62500e-08*ic_cap+7.26000e-06'
+ mcm5p1_ca_w_4_000_s_4_800 = '-5.71875e-08*ic_cap*ic_cap+-3.62500e-08*ic_cap+7.26000e-06'
+ mcm5p1_cc_w_1_600_s_10_000 = '1.25000e-14*ic_cap*ic_cap+1.31000e-11'
+ mcm5p1_cc_w_1_600_s_12_000 = '1.56250e-14*ic_cap*ic_cap+1.25000e-14*ic_cap+1.03000e-11'
+ mcm5p1_cc_w_1_600_s_1_600 = '-4.62500e-13*ic_cap*ic_cap+-3.00000e-13*ic_cap+7.27000e-11'
+ mcm5p1_cc_w_1_600_s_1_700 = '-4.18750e-13*ic_cap*ic_cap+-2.75000e-13*ic_cap+6.91000e-11'
+ mcm5p1_cc_w_1_600_s_1_900 = '-3.43750e-13*ic_cap*ic_cap+-2.25000e-13*ic_cap+6.28000e-11'
+ mcm5p1_cc_w_1_600_s_2_000 = '-3.09375e-13*ic_cap*ic_cap+-2.12500e-13*ic_cap+6.02000e-11'
+ mcm5p1_cc_w_1_600_s_2_400 = '-2.25000e-13*ic_cap*ic_cap+-1.50000e-13*ic_cap+5.18000e-11'
+ mcm5p1_cc_w_1_600_s_2_800 = '-1.68750e-13*ic_cap*ic_cap+-1.25000e-13*ic_cap+4.56000e-11'
+ mcm5p1_cc_w_1_600_s_3_200 = '-1.28125e-13*ic_cap*ic_cap+-8.75000e-14*ic_cap+4.08000e-11'
+ mcm5p1_cc_w_1_600_s_4_800 = '-4.68750e-14*ic_cap*ic_cap+-3.75000e-14*ic_cap+2.86000e-11'
+ mcm5p1_cc_w_4_000_s_10_000 = '2.50000e-14*ic_cap*ic_cap+2.50000e-14*ic_cap+1.56000e-11'
+ mcm5p1_cc_w_4_000_s_12_000 = '2.18750e-14*ic_cap*ic_cap+1.25000e-14*ic_cap+1.26000e-11'
+ mcm5p1_cc_w_4_000_s_1_600 = '-4.21875e-13*ic_cap*ic_cap+-2.87500e-13*ic_cap+7.93000e-11'
+ mcm5p1_cc_w_4_000_s_1_700 = '-3.81250e-13*ic_cap*ic_cap+-2.50000e-13*ic_cap+7.54000e-11'
+ mcm5p1_cc_w_4_000_s_1_900 = '-3.12500e-13*ic_cap*ic_cap+-2.00000e-13*ic_cap+6.89000e-11'
+ mcm5p1_cc_w_4_000_s_2_000 = '-2.84375e-13*ic_cap*ic_cap+-1.87500e-13*ic_cap+6.62000e-11'
+ mcm5p1_cc_w_4_000_s_2_400 = '-1.87500e-13*ic_cap*ic_cap+-1.25000e-13*ic_cap+5.71000e-11'
+ mcm5p1_cc_w_4_000_s_2_800 = '-1.37500e-13*ic_cap*ic_cap+-1.00000e-13*ic_cap+5.06000e-11'
+ mcm5p1_cc_w_4_000_s_3_200 = '-1.03125e-13*ic_cap*ic_cap+-8.75000e-14*ic_cap+4.55000e-11'
+ mcm5p1_cc_w_4_000_s_4_800 = '-3.12500e-14*ic_cap*ic_cap+-2.50000e-14*ic_cap+3.25000e-11'
+ mcm5p1_cf_w_1_600_s_10_000 = '-1.46875e-13*ic_cap*ic_cap+-8.75000e-14*ic_cap+2.45000e-11'
+ mcm5p1_cf_w_1_600_s_12_000 = '-1.56250e-13*ic_cap*ic_cap+-1.00000e-13*ic_cap+2.68000e-11'
+ mcm5p1_cf_w_1_600_s_1_600 = '-2.56250e-14*ic_cap*ic_cap+-1.75000e-14*ic_cap+5.59000e-12'
+ mcm5p1_cf_w_1_600_s_1_700 = '-2.84375e-14*ic_cap*ic_cap+-1.87500e-14*ic_cap+5.92000e-12'
+ mcm5p1_cf_w_1_600_s_1_900 = '-3.34375e-14*ic_cap*ic_cap+-2.12500e-14*ic_cap+6.58000e-12'
+ mcm5p1_cf_w_1_600_s_2_000 = '-3.65625e-14*ic_cap*ic_cap+-2.37500e-14*ic_cap+6.91000e-12'
+ mcm5p1_cf_w_1_600_s_2_400 = '-4.62500e-14*ic_cap*ic_cap+-3.00000e-14*ic_cap+8.18000e-12'
+ mcm5p1_cf_w_1_600_s_2_800 = '-5.53125e-14*ic_cap*ic_cap+-3.62500e-14*ic_cap+9.41000e-12'
+ mcm5p1_cf_w_1_600_s_3_200 = '-6.43750e-14*ic_cap*ic_cap+-4.00000e-14*ic_cap+1.06000e-11'
+ mcm5p1_cf_w_1_600_s_4_800 = '-9.68750e-14*ic_cap*ic_cap+-6.25000e-14*ic_cap+1.49000e-11'
+ mcm5p1_cf_w_4_000_s_10_000 = '-1.40625e-13*ic_cap*ic_cap+-8.75000e-14*ic_cap+2.49000e-11'
+ mcm5p1_cf_w_4_000_s_12_000 = '-1.50000e-13*ic_cap*ic_cap+-1.00000e-13*ic_cap+2.74000e-11'
+ mcm5p1_cf_w_4_000_s_1_600 = '-2.65625e-14*ic_cap*ic_cap+-1.62500e-14*ic_cap+5.61000e-12'
+ mcm5p1_cf_w_4_000_s_1_700 = '-2.87500e-14*ic_cap*ic_cap+-1.75000e-14*ic_cap+5.94000e-12'
+ mcm5p1_cf_w_4_000_s_1_900 = '-3.34375e-14*ic_cap*ic_cap+-2.12500e-14*ic_cap+6.59000e-12'
+ mcm5p1_cf_w_4_000_s_2_000 = '-3.65625e-14*ic_cap*ic_cap+-2.37500e-14*ic_cap+6.92000e-12'
+ mcm5p1_cf_w_4_000_s_2_400 = '-4.59375e-14*ic_cap*ic_cap+-3.12500e-14*ic_cap+8.19000e-12'
+ mcm5p1_cf_w_4_000_s_2_800 = '-5.53125e-14*ic_cap*ic_cap+-3.62500e-14*ic_cap+9.43000e-12'
+ mcm5p1_cf_w_4_000_s_3_200 = '-6.21875e-14*ic_cap*ic_cap+-4.12500e-14*ic_cap+1.06000e-11'
+ mcm5p1_cf_w_4_000_s_4_800 = '-9.68750e-14*ic_cap*ic_cap+-6.25000e-14*ic_cap+1.50000e-11'
+ mcm5p1f_ca_w_0_150_s_0_210 = '-1.44375e-06*ic_cap*ic_cap+-8.25000e-07*ic_cap+1.13000e-04'
+ mcm5p1f_ca_w_0_150_s_0_263 = '-1.44375e-06*ic_cap*ic_cap+-8.25000e-07*ic_cap+1.13000e-04'
+ mcm5p1f_ca_w_0_150_s_0_315 = '-1.44375e-06*ic_cap*ic_cap+-8.25000e-07*ic_cap+1.13000e-04'
+ mcm5p1f_ca_w_0_150_s_0_420 = '-1.44375e-06*ic_cap*ic_cap+-8.25000e-07*ic_cap+1.13000e-04'
+ mcm5p1f_ca_w_0_150_s_0_525 = '-1.44375e-06*ic_cap*ic_cap+-8.25000e-07*ic_cap+1.13000e-04'
+ mcm5p1f_ca_w_0_150_s_0_630 = '-1.44375e-06*ic_cap*ic_cap+-8.25000e-07*ic_cap+1.13000e-04'
+ mcm5p1f_ca_w_0_150_s_0_840 = '-1.44375e-06*ic_cap*ic_cap+-8.25000e-07*ic_cap+1.13000e-04'
+ mcm5p1f_ca_w_0_150_s_1_260 = '-1.44375e-06*ic_cap*ic_cap+-8.25000e-07*ic_cap+1.13000e-04'
+ mcm5p1f_ca_w_0_150_s_2_310 = '-1.44375e-06*ic_cap*ic_cap+-8.25000e-07*ic_cap+1.13000e-04'
+ mcm5p1f_ca_w_0_150_s_5_250 = '-1.44375e-06*ic_cap*ic_cap+-8.25000e-07*ic_cap+1.13000e-04'
+ mcm5p1f_ca_w_1_200_s_0_210 = '-1.44375e-06*ic_cap*ic_cap+-8.25000e-07*ic_cap+1.13000e-04'
+ mcm5p1f_ca_w_1_200_s_0_263 = '-1.44375e-06*ic_cap*ic_cap+-8.25000e-07*ic_cap+1.13000e-04'
+ mcm5p1f_ca_w_1_200_s_0_315 = '-1.44375e-06*ic_cap*ic_cap+-8.25000e-07*ic_cap+1.13000e-04'
+ mcm5p1f_ca_w_1_200_s_0_420 = '-1.44375e-06*ic_cap*ic_cap+-8.25000e-07*ic_cap+1.13000e-04'
+ mcm5p1f_ca_w_1_200_s_0_525 = '-1.44375e-06*ic_cap*ic_cap+-8.25000e-07*ic_cap+1.13000e-04'
+ mcm5p1f_ca_w_1_200_s_0_630 = '-1.44375e-06*ic_cap*ic_cap+-8.25000e-07*ic_cap+1.13000e-04'
+ mcm5p1f_ca_w_1_200_s_0_840 = '-1.44375e-06*ic_cap*ic_cap+-8.25000e-07*ic_cap+1.13000e-04'
+ mcm5p1f_ca_w_1_200_s_1_260 = '-1.44375e-06*ic_cap*ic_cap+-8.25000e-07*ic_cap+1.13000e-04'
+ mcm5p1f_ca_w_1_200_s_2_310 = '-1.44375e-06*ic_cap*ic_cap+-8.25000e-07*ic_cap+1.13000e-04'
+ mcm5p1f_ca_w_1_200_s_5_250 = '-1.44375e-06*ic_cap*ic_cap+-8.25000e-07*ic_cap+1.13000e-04'
+ mcm5p1f_cc_w_0_150_s_0_210 = '-5.62500e-13*ic_cap*ic_cap+-3.25000e-13*ic_cap+7.51000e-11'
+ mcm5p1f_cc_w_0_150_s_0_263 = '-3.65625e-13*ic_cap*ic_cap+-2.12500e-13*ic_cap+6.08000e-11'
+ mcm5p1f_cc_w_0_150_s_0_315 = '-2.56250e-13*ic_cap*ic_cap+-1.50000e-13*ic_cap+5.15000e-11'
+ mcm5p1f_cc_w_0_150_s_0_420 = '-1.34375e-13*ic_cap*ic_cap+-8.75000e-14*ic_cap+3.89000e-11'
+ mcm5p1f_cc_w_0_150_s_0_525 = '-7.50000e-14*ic_cap*ic_cap+-5.00000e-14*ic_cap+3.12000e-11'
+ mcm5p1f_cc_w_0_150_s_0_630 = '-3.12500e-14*ic_cap*ic_cap+-2.50000e-14*ic_cap+2.56000e-11'
+ mcm5p1f_cc_w_0_150_s_0_840 = '6.25000e-15*ic_cap*ic_cap+1.81000e-11'
+ mcm5p1f_cc_w_0_150_s_1_260 = '2.31250e-14*ic_cap*ic_cap+2.50000e-14*ic_cap+9.93000e-12'
+ mcm5p1f_cc_w_0_150_s_2_310 = '2.21875e-14*ic_cap*ic_cap+1.62500e-14*ic_cap+3.34000e-12'
+ mcm5p1f_cc_w_0_150_s_5_250 = '2.90625e-15*ic_cap*ic_cap+4.37500e-15*ic_cap+4.63000e-13'
+ mcm5p1f_cc_w_1_200_s_0_210 = '-5.34375e-13*ic_cap*ic_cap+-3.12500e-13*ic_cap+9.02000e-11'
+ mcm5p1f_cc_w_1_200_s_0_263 = '-3.34375e-13*ic_cap*ic_cap+-1.87500e-13*ic_cap+7.46000e-11'
+ mcm5p1f_cc_w_1_200_s_0_315 = '-2.25000e-13*ic_cap*ic_cap+-1.25000e-13*ic_cap+6.41000e-11'
+ mcm5p1f_cc_w_1_200_s_0_420 = '-1.03125e-13*ic_cap*ic_cap+-6.25000e-14*ic_cap+5.02000e-11'
+ mcm5p1f_cc_w_1_200_s_0_525 = '-3.75000e-14*ic_cap*ic_cap+-2.50000e-14*ic_cap+4.11000e-11'
+ mcm5p1f_cc_w_1_200_s_0_630 = '-9.37500e-15*ic_cap*ic_cap+-1.25000e-14*ic_cap+3.47000e-11'
+ mcm5p1f_cc_w_1_200_s_0_840 = '2.81250e-14*ic_cap*ic_cap+3.75000e-14*ic_cap+2.59000e-11'
+ mcm5p1f_cc_w_1_200_s_1_260 = '4.68750e-14*ic_cap*ic_cap+3.75000e-14*ic_cap+1.60000e-11'
+ mcm5p1f_cc_w_1_200_s_2_310 = '4.37500e-14*ic_cap*ic_cap+3.00000e-14*ic_cap+6.20000e-12'
+ mcm5p1f_cc_w_1_200_s_5_250 = '1.59375e-14*ic_cap*ic_cap+1.12500e-14*ic_cap+8.40000e-13'
+ mcm5p1f_cf_w_0_150_s_0_210 = '-9.37500e-14*ic_cap*ic_cap+-5.25000e-14*ic_cap+1.11000e-11'
+ mcm5p1f_cf_w_0_150_s_0_263 = '-1.18750e-13*ic_cap*ic_cap+-7.50000e-14*ic_cap+1.34000e-11'
+ mcm5p1f_cf_w_0_150_s_0_315 = '-1.46875e-13*ic_cap*ic_cap+-8.75000e-14*ic_cap+1.57000e-11'
+ mcm5p1f_cf_w_0_150_s_0_420 = '-1.90625e-13*ic_cap*ic_cap+-1.12500e-13*ic_cap+1.99000e-11'
+ mcm5p1f_cf_w_0_150_s_0_525 = '-2.21875e-13*ic_cap*ic_cap+-1.37500e-13*ic_cap+2.34000e-11'
+ mcm5p1f_cf_w_0_150_s_0_630 = '-2.50000e-13*ic_cap*ic_cap+-1.50000e-13*ic_cap+2.65000e-11'
+ mcm5p1f_cf_w_0_150_s_0_840 = '-2.84375e-13*ic_cap*ic_cap+-1.62500e-13*ic_cap+3.15000e-11'
+ mcm5p1f_cf_w_0_150_s_1_260 = '-3.03125e-13*ic_cap*ic_cap+-1.87500e-13*ic_cap+3.81000e-11'
+ mcm5p1f_cf_w_0_150_s_2_310 = '-3.09375e-13*ic_cap*ic_cap+-1.87500e-13*ic_cap+4.40000e-11'
+ mcm5p1f_cf_w_0_150_s_5_250 = '-2.93750e-13*ic_cap*ic_cap+-1.75000e-13*ic_cap+4.69000e-11'
+ mcm5p1f_cf_w_1_200_s_0_210 = '-9.18750e-14*ic_cap*ic_cap+-5.25000e-14*ic_cap+1.10000e-11'
+ mcm5p1f_cf_w_1_200_s_0_263 = '-1.18750e-13*ic_cap*ic_cap+-7.50000e-14*ic_cap+1.34000e-11'
+ mcm5p1f_cf_w_1_200_s_0_315 = '-1.43750e-13*ic_cap*ic_cap+-7.50000e-14*ic_cap+1.57000e-11'
+ mcm5p1f_cf_w_1_200_s_0_420 = '-1.81250e-13*ic_cap*ic_cap+-1.00000e-13*ic_cap+1.98000e-11'
+ mcm5p1f_cf_w_1_200_s_0_525 = '-2.18750e-13*ic_cap*ic_cap+-1.25000e-13*ic_cap+2.35000e-11'
+ mcm5p1f_cf_w_1_200_s_0_630 = '-2.40625e-13*ic_cap*ic_cap+-1.37500e-13*ic_cap+2.67000e-11'
+ mcm5p1f_cf_w_1_200_s_0_840 = '-2.78125e-13*ic_cap*ic_cap+-1.62500e-13*ic_cap+3.21000e-11'
+ mcm5p1f_cf_w_1_200_s_1_260 = '-3.09375e-13*ic_cap*ic_cap+-1.87500e-13*ic_cap+3.94000e-11'
+ mcm5p1f_cf_w_1_200_s_2_310 = '-3.09375e-13*ic_cap*ic_cap+-1.87500e-13*ic_cap+4.79000e-11'
+ mcm5p1f_cf_w_1_200_s_5_250 = '-2.87500e-13*ic_cap*ic_cap+-1.75000e-13*ic_cap+5.31000e-11'
+ mcp1f_ca_w_0_150_s_0_210 = '-1.40313e-06*ic_cap*ic_cap+-7.87500e-07*ic_cap+1.06000e-04'
+ mcp1f_ca_w_0_150_s_0_263 = '-1.40313e-06*ic_cap*ic_cap+-7.87500e-07*ic_cap+1.06000e-04'
+ mcp1f_ca_w_0_150_s_0_315 = '-1.40313e-06*ic_cap*ic_cap+-7.87500e-07*ic_cap+1.06000e-04'
+ mcp1f_ca_w_0_150_s_0_420 = '-1.40313e-06*ic_cap*ic_cap+-7.87500e-07*ic_cap+1.06000e-04'
+ mcp1f_ca_w_0_150_s_0_525 = '-1.40313e-06*ic_cap*ic_cap+-7.87500e-07*ic_cap+1.06000e-04'
+ mcp1f_ca_w_0_150_s_0_630 = '-1.40313e-06*ic_cap*ic_cap+-7.87500e-07*ic_cap+1.06000e-04'
+ mcp1f_ca_w_0_150_s_0_840 = '-1.40313e-06*ic_cap*ic_cap+-7.87500e-07*ic_cap+1.06000e-04'
+ mcp1f_ca_w_0_150_s_1_260 = '-1.40313e-06*ic_cap*ic_cap+-7.87500e-07*ic_cap+1.06000e-04'
+ mcp1f_ca_w_0_150_s_2_310 = '-1.40313e-06*ic_cap*ic_cap+-7.87500e-07*ic_cap+1.06000e-04'
+ mcp1f_ca_w_0_150_s_5_250 = '-1.40313e-06*ic_cap*ic_cap+-7.87500e-07*ic_cap+1.06000e-04'
+ mcp1f_ca_w_1_200_s_0_210 = '-1.40313e-06*ic_cap*ic_cap+-7.87500e-07*ic_cap+1.06000e-04'
+ mcp1f_ca_w_1_200_s_0_263 = '-1.40313e-06*ic_cap*ic_cap+-7.87500e-07*ic_cap+1.06000e-04'
+ mcp1f_ca_w_1_200_s_0_315 = '-1.40313e-06*ic_cap*ic_cap+-7.87500e-07*ic_cap+1.06000e-04'
+ mcp1f_ca_w_1_200_s_0_420 = '-1.40313e-06*ic_cap*ic_cap+-7.87500e-07*ic_cap+1.06000e-04'
+ mcp1f_ca_w_1_200_s_0_525 = '-1.40313e-06*ic_cap*ic_cap+-7.87500e-07*ic_cap+1.06000e-04'
+ mcp1f_ca_w_1_200_s_0_630 = '-1.40313e-06*ic_cap*ic_cap+-7.87500e-07*ic_cap+1.06000e-04'
+ mcp1f_ca_w_1_200_s_0_840 = '-1.40313e-06*ic_cap*ic_cap+-7.87500e-07*ic_cap+1.06000e-04'
+ mcp1f_ca_w_1_200_s_1_260 = '-1.40313e-06*ic_cap*ic_cap+-7.87500e-07*ic_cap+1.06000e-04'
+ mcp1f_ca_w_1_200_s_2_310 = '-1.40313e-06*ic_cap*ic_cap+-7.87500e-07*ic_cap+1.06000e-04'
+ mcp1f_ca_w_1_200_s_5_250 = '-1.40313e-06*ic_cap*ic_cap+-7.87500e-07*ic_cap+1.06000e-04'
+ mcp1f_cc_w_0_150_s_0_210 = '-5.81250e-13*ic_cap*ic_cap+-3.25000e-13*ic_cap+7.62000e-11'
+ mcp1f_cc_w_0_150_s_0_263 = '-3.78125e-13*ic_cap*ic_cap+-2.12500e-13*ic_cap+6.19000e-11'
+ mcp1f_cc_w_0_150_s_0_315 = '-2.59375e-13*ic_cap*ic_cap+-1.62500e-13*ic_cap+5.27000e-11'
+ mcp1f_cc_w_0_150_s_0_420 = '-1.46875e-13*ic_cap*ic_cap+-8.75000e-14*ic_cap+4.04000e-11'
+ mcp1f_cc_w_0_150_s_0_525 = '-8.43750e-14*ic_cap*ic_cap+-6.25000e-14*ic_cap+3.29000e-11'
+ mcp1f_cc_w_0_150_s_0_630 = '-4.68750e-14*ic_cap*ic_cap+-3.75000e-14*ic_cap+2.76000e-11'
+ mcp1f_cc_w_0_150_s_0_840 = '-1.25000e-14*ic_cap*ic_cap+2.03000e-11'
+ mcp1f_cc_w_0_150_s_1_260 = '1.56250e-14*ic_cap*ic_cap+1.25000e-14*ic_cap+1.18000e-11'
+ mcp1f_cc_w_0_150_s_2_310 = '1.53125e-14*ic_cap*ic_cap+8.75000e-15*ic_cap+5.10000e-12'
+ mcp1f_cc_w_0_150_s_5_250 = '2.81250e-15*ic_cap*ic_cap+1.25000e-15*ic_cap+1.20000e-12'
+ mcp1f_cc_w_1_200_s_0_210 = '-5.68750e-13*ic_cap*ic_cap+-3.00000e-13*ic_cap+9.44000e-11'
+ mcp1f_cc_w_1_200_s_0_263 = '-3.65625e-13*ic_cap*ic_cap+-2.12500e-13*ic_cap+7.89000e-11'
+ mcp1f_cc_w_1_200_s_0_315 = '-2.62500e-13*ic_cap*ic_cap+-1.50000e-13*ic_cap+6.86000e-11'
+ mcp1f_cc_w_1_200_s_0_420 = '-1.37500e-13*ic_cap*ic_cap+-7.50000e-14*ic_cap+5.49000e-11'
+ mcp1f_cc_w_1_200_s_0_525 = '-8.43750e-14*ic_cap*ic_cap+-3.75000e-14*ic_cap+4.61000e-11'
+ mcp1f_cc_w_1_200_s_0_630 = '-4.68750e-14*ic_cap*ic_cap+-3.75000e-14*ic_cap+3.98000e-11'
+ mcp1f_cc_w_1_200_s_0_840 = '-1.25000e-14*ic_cap*ic_cap+3.12000e-11'
+ mcp1f_cc_w_1_200_s_1_260 = '9.37500e-15*ic_cap*ic_cap+1.25000e-14*ic_cap+2.14000e-11'
+ mcp1f_cc_w_1_200_s_2_310 = '1.56250e-14*ic_cap*ic_cap+1.25000e-14*ic_cap+1.08000e-11'
+ mcp1f_cc_w_1_200_s_5_250 = '1.09375e-14*ic_cap*ic_cap+6.25000e-15*ic_cap+3.40000e-12'
+ mcp1f_cf_w_0_150_s_0_210 = '-8.87500e-14*ic_cap*ic_cap+-5.00000e-14*ic_cap+1.03000e-11'
+ mcp1f_cf_w_0_150_s_0_263 = '-1.15625e-13*ic_cap*ic_cap+-6.25000e-14*ic_cap+1.25000e-11'
+ mcp1f_cf_w_0_150_s_0_315 = '-1.37500e-13*ic_cap*ic_cap+-7.50000e-14*ic_cap+1.45000e-11'
+ mcp1f_cf_w_0_150_s_0_420 = '-1.81250e-13*ic_cap*ic_cap+-1.00000e-13*ic_cap+1.85000e-11'
+ mcp1f_cf_w_0_150_s_0_525 = '-2.06250e-13*ic_cap*ic_cap+-1.25000e-13*ic_cap+2.17000e-11'
+ mcp1f_cf_w_0_150_s_0_630 = '-2.34375e-13*ic_cap*ic_cap+-1.37500e-13*ic_cap+2.46000e-11'
+ mcp1f_cf_w_0_150_s_0_840 = '-2.68750e-13*ic_cap*ic_cap+-1.50000e-13*ic_cap+2.94000e-11'
+ mcp1f_cf_w_0_150_s_1_260 = '-2.96875e-13*ic_cap*ic_cap+-1.87500e-13*ic_cap+3.62000e-11'
+ mcp1f_cf_w_0_150_s_2_310 = '-3.06250e-13*ic_cap*ic_cap+-1.75000e-13*ic_cap+4.24000e-11'
+ mcp1f_cf_w_0_150_s_5_250 = '-2.93750e-13*ic_cap*ic_cap+-1.75000e-13*ic_cap+4.63000e-11'
+ mcp1f_cf_w_1_200_s_0_210 = '-8.65625e-14*ic_cap*ic_cap+-4.87500e-14*ic_cap+1.02000e-11'
+ mcp1f_cf_w_1_200_s_0_263 = '-1.15625e-13*ic_cap*ic_cap+-6.25000e-14*ic_cap+1.25000e-11'
+ mcp1f_cf_w_1_200_s_0_315 = '-1.40625e-13*ic_cap*ic_cap+-8.75000e-14*ic_cap+1.46000e-11'
+ mcp1f_cf_w_1_200_s_0_420 = '-1.75000e-13*ic_cap*ic_cap+-1.00000e-13*ic_cap+1.84000e-11'
+ mcp1f_cf_w_1_200_s_0_525 = '-2.12500e-13*ic_cap*ic_cap+-1.25000e-13*ic_cap+2.19000e-11'
+ mcp1f_cf_w_1_200_s_0_630 = '-2.34375e-13*ic_cap*ic_cap+-1.37500e-13*ic_cap+2.49000e-11'
+ mcp1f_cf_w_1_200_s_0_840 = '-2.62500e-13*ic_cap*ic_cap+-1.50000e-13*ic_cap+2.99000e-11'
+ mcp1f_cf_w_1_200_s_1_260 = '-2.93750e-13*ic_cap*ic_cap+-1.75000e-13*ic_cap+3.71000e-11'
+ mcp1f_cf_w_1_200_s_2_310 = '-3.09375e-13*ic_cap*ic_cap+-1.87500e-13*ic_cap+4.64000e-11'
+ mcp1f_cf_w_1_200_s_5_250 = '-3.06250e-13*ic_cap*ic_cap+-1.75000e-13*ic_cap+5.36000e-11'
+ mcrdld_ca_w_10_000_s_10_000 = '-2.28125e-08*ic_cap*ic_cap+-1.37500e-08*ic_cap+2.63000e-06'
+ mcrdld_ca_w_10_000_s_12_000 = '-2.28125e-08*ic_cap*ic_cap+-1.37500e-08*ic_cap+2.63000e-06'
+ mcrdld_ca_w_10_000_s_30_000 = '-2.28125e-08*ic_cap*ic_cap+-1.37500e-08*ic_cap+2.63000e-06'
+ mcrdld_ca_w_10_000_s_5_000 = '-2.28125e-08*ic_cap*ic_cap+-1.37500e-08*ic_cap+2.63000e-06'
+ mcrdld_ca_w_10_000_s_8_000 = '-2.28125e-08*ic_cap*ic_cap+-1.37500e-08*ic_cap+2.63000e-06'
+ mcrdld_ca_w_40_000_s_10_000 = '-2.28125e-08*ic_cap*ic_cap+-1.37500e-08*ic_cap+2.63000e-06'
+ mcrdld_ca_w_40_000_s_12_000 = '-2.28125e-08*ic_cap*ic_cap+-1.37500e-08*ic_cap+2.63000e-06'
+ mcrdld_ca_w_40_000_s_30_000 = '-2.28125e-08*ic_cap*ic_cap+-1.37500e-08*ic_cap+2.63000e-06'
+ mcrdld_ca_w_40_000_s_5_000 = '-2.28125e-08*ic_cap*ic_cap+-1.37500e-08*ic_cap+2.63000e-06'
+ mcrdld_ca_w_40_000_s_8_000 = '-2.28125e-08*ic_cap*ic_cap+-1.37500e-08*ic_cap+2.63000e-06'
+ mcrdld_cc_w_10_000_s_10_000 = '-2.43750e-13*ic_cap*ic_cap+-1.50000e-13*ic_cap+3.18000e-11'
+ mcrdld_cc_w_10_000_s_12_000 = '-1.96875e-13*ic_cap*ic_cap+-1.37500e-13*ic_cap+2.78000e-11'
+ mcrdld_cc_w_10_000_s_30_000 = '-6.25000e-14*ic_cap*ic_cap+-5.00000e-14*ic_cap+1.22000e-11'
+ mcrdld_cc_w_10_000_s_5_000 = '-5.68750e-13*ic_cap*ic_cap+-3.50000e-13*ic_cap+5.14000e-11'
+ mcrdld_cc_w_10_000_s_8_000 = '-3.18750e-13*ic_cap*ic_cap+-2.00000e-13*ic_cap+3.73000e-11'
+ mcrdld_cc_w_40_000_s_10_000 = '-2.43750e-13*ic_cap*ic_cap+-1.50000e-13*ic_cap+4.17000e-11'
+ mcrdld_cc_w_40_000_s_12_000 = '-1.90625e-13*ic_cap*ic_cap+-1.37500e-13*ic_cap+3.72000e-11'
+ mcrdld_cc_w_40_000_s_30_000 = '-6.25000e-14*ic_cap*ic_cap+-5.00000e-14*ic_cap+1.94000e-11'
+ mcrdld_cc_w_40_000_s_5_000 = '-5.65625e-13*ic_cap*ic_cap+-3.37500e-13*ic_cap+6.27000e-11'
+ mcrdld_cc_w_40_000_s_8_000 = '-3.12500e-13*ic_cap*ic_cap+-2.00000e-13*ic_cap+4.76000e-11'
+ mcrdld_cf_w_10_000_s_10_000 = '-4.06250e-14*ic_cap*ic_cap+-3.75000e-14*ic_cap+1.11000e-11'
+ mcrdld_cf_w_10_000_s_12_000 = '-5.31250e-14*ic_cap*ic_cap+-3.75000e-14*ic_cap+1.28000e-11'
+ mcrdld_cf_w_10_000_s_30_000 = '-1.28125e-13*ic_cap*ic_cap+-8.75000e-14*ic_cap+2.31000e-11'
+ mcrdld_cf_w_10_000_s_5_000 = '3.12500e-16*ic_cap*ic_cap+-1.25000e-15*ic_cap+6.11000e-12'
+ mcrdld_cf_w_10_000_s_8_000 = '-2.62500e-14*ic_cap*ic_cap+-1.75000e-14*ic_cap+9.23000e-12'
+ mcrdld_cf_w_40_000_s_10_000 = '-4.06250e-14*ic_cap*ic_cap+-3.75000e-14*ic_cap+1.12000e-11'
+ mcrdld_cf_w_40_000_s_12_000 = '-5.93750e-14*ic_cap*ic_cap+-3.75000e-14*ic_cap+1.30000e-11'
+ mcrdld_cf_w_40_000_s_30_000 = '-1.21875e-13*ic_cap*ic_cap+-8.75000e-14*ic_cap+2.38000e-11'
+ mcrdld_cf_w_40_000_s_5_000 = '-1.87500e-15*ic_cap*ic_cap+-2.50000e-15*ic_cap+6.23000e-12'
+ mcrdld_cf_w_40_000_s_8_000 = '-2.84375e-14*ic_cap*ic_cap+-1.87500e-14*ic_cap+9.36000e-12'
+ mcrdlf_ca_w_10_000_s_10_000 = '-2.28125e-08*ic_cap*ic_cap+-1.37500e-08*ic_cap+2.57000e-06'
+ mcrdlf_ca_w_10_000_s_12_000 = '-2.28125e-08*ic_cap*ic_cap+-1.37500e-08*ic_cap+2.57000e-06'
+ mcrdlf_ca_w_10_000_s_30_000 = '-2.28125e-08*ic_cap*ic_cap+-1.37500e-08*ic_cap+2.57000e-06'
+ mcrdlf_ca_w_10_000_s_5_000 = '-2.28125e-08*ic_cap*ic_cap+-1.37500e-08*ic_cap+2.57000e-06'
+ mcrdlf_ca_w_10_000_s_8_000 = '-2.28125e-08*ic_cap*ic_cap+-1.37500e-08*ic_cap+2.57000e-06'
+ mcrdlf_ca_w_40_000_s_10_000 = '-2.28125e-08*ic_cap*ic_cap+-1.37500e-08*ic_cap+2.57000e-06'
+ mcrdlf_ca_w_40_000_s_12_000 = '-2.28125e-08*ic_cap*ic_cap+-1.37500e-08*ic_cap+2.57000e-06'
+ mcrdlf_ca_w_40_000_s_30_000 = '-2.28125e-08*ic_cap*ic_cap+-1.37500e-08*ic_cap+2.57000e-06'
+ mcrdlf_ca_w_40_000_s_5_000 = '-2.28125e-08*ic_cap*ic_cap+-1.37500e-08*ic_cap+2.57000e-06'
+ mcrdlf_ca_w_40_000_s_8_000 = '-2.28125e-08*ic_cap*ic_cap+-1.37500e-08*ic_cap+2.57000e-06'
+ mcrdlf_cc_w_10_000_s_10_000 = '-2.40625e-13*ic_cap*ic_cap+-1.62500e-13*ic_cap+3.20000e-11'
+ mcrdlf_cc_w_10_000_s_12_000 = '-1.93750e-13*ic_cap*ic_cap+-1.25000e-13*ic_cap+2.80000e-11'
+ mcrdlf_cc_w_10_000_s_30_000 = '-5.93750e-14*ic_cap*ic_cap+-3.75000e-14*ic_cap+1.23000e-11'
+ mcrdlf_cc_w_10_000_s_5_000 = '-5.68750e-13*ic_cap*ic_cap+-3.50000e-13*ic_cap+5.16000e-11'
+ mcrdlf_cc_w_10_000_s_8_000 = '-3.18750e-13*ic_cap*ic_cap+-2.00000e-13*ic_cap+3.75000e-11'
+ mcrdlf_cc_w_40_000_s_10_000 = '-2.50000e-13*ic_cap*ic_cap+-1.50000e-13*ic_cap+4.20000e-11'
+ mcrdlf_cc_w_40_000_s_12_000 = '-1.90625e-13*ic_cap*ic_cap+-1.12500e-13*ic_cap+3.74000e-11'
+ mcrdlf_cc_w_40_000_s_30_000 = '-5.93750e-14*ic_cap*ic_cap+-3.75000e-14*ic_cap+1.95000e-11'
+ mcrdlf_cc_w_40_000_s_5_000 = '-5.62500e-13*ic_cap*ic_cap+-3.50000e-13*ic_cap+6.29000e-11'
+ mcrdlf_cc_w_40_000_s_8_000 = '-3.18750e-13*ic_cap*ic_cap+-2.00000e-13*ic_cap+4.79000e-11'
+ mcrdlf_cf_w_10_000_s_10_000 = '-4.37500e-14*ic_cap*ic_cap+-2.50000e-14*ic_cap+1.09000e-11'
+ mcrdlf_cf_w_10_000_s_12_000 = '-5.93750e-14*ic_cap*ic_cap+-3.75000e-14*ic_cap+1.26000e-11'
+ mcrdlf_cf_w_10_000_s_30_000 = '-1.28125e-13*ic_cap*ic_cap+-8.75000e-14*ic_cap+2.28000e-11'
+ mcrdlf_cf_w_10_000_s_5_000 = '6.25000e-16*ic_cap*ic_cap+5.97000e-12'
+ mcrdlf_cf_w_10_000_s_8_000 = '-2.65625e-14*ic_cap*ic_cap+-1.87500e-14*ic_cap+9.04000e-12'
+ mcrdlf_cf_w_40_000_s_10_000 = '-4.37500e-14*ic_cap*ic_cap+-2.50000e-14*ic_cap+1.10000e-11'
+ mcrdlf_cf_w_40_000_s_12_000 = '-5.31250e-14*ic_cap*ic_cap+-3.75000e-14*ic_cap+1.27000e-11'
+ mcrdlf_cf_w_40_000_s_30_000 = '-1.21875e-13*ic_cap*ic_cap+-8.75000e-14*ic_cap+2.35000e-11'
+ mcrdlf_cf_w_40_000_s_5_000 = '-1.56250e-15*ic_cap*ic_cap+-1.25000e-15*ic_cap+6.08000e-12'
+ mcrdlf_cf_w_40_000_s_8_000 = '-2.87500e-14*ic_cap*ic_cap+-1.75000e-14*ic_cap+9.16000e-12'
+ mcrdll1_ca_w_10_000_s_10_000 = '-2.43750e-08*ic_cap*ic_cap+-1.50000e-08*ic_cap+2.78000e-06'
+ mcrdll1_ca_w_10_000_s_12_000 = '-2.43750e-08*ic_cap*ic_cap+-1.50000e-08*ic_cap+2.78000e-06'
+ mcrdll1_ca_w_10_000_s_30_000 = '-2.43750e-08*ic_cap*ic_cap+-1.50000e-08*ic_cap+2.78000e-06'
+ mcrdll1_ca_w_10_000_s_5_000 = '-2.43750e-08*ic_cap*ic_cap+-1.50000e-08*ic_cap+2.78000e-06'
+ mcrdll1_ca_w_10_000_s_8_000 = '-2.43750e-08*ic_cap*ic_cap+-1.50000e-08*ic_cap+2.78000e-06'
+ mcrdll1_ca_w_40_000_s_10_000 = '-2.43750e-08*ic_cap*ic_cap+-1.50000e-08*ic_cap+2.78000e-06'
+ mcrdll1_ca_w_40_000_s_12_000 = '-2.43750e-08*ic_cap*ic_cap+-1.50000e-08*ic_cap+2.78000e-06'
+ mcrdll1_ca_w_40_000_s_30_000 = '-2.43750e-08*ic_cap*ic_cap+-1.50000e-08*ic_cap+2.78000e-06'
+ mcrdll1_ca_w_40_000_s_5_000 = '-2.43750e-08*ic_cap*ic_cap+-1.50000e-08*ic_cap+2.78000e-06'
+ mcrdll1_ca_w_40_000_s_8_000 = '-2.43750e-08*ic_cap*ic_cap+-1.50000e-08*ic_cap+2.78000e-06'
+ mcrdll1_cc_w_10_000_s_10_000 = '-2.40625e-13*ic_cap*ic_cap+-1.62500e-13*ic_cap+3.13000e-11'
+ mcrdll1_cc_w_10_000_s_12_000 = '-2.00000e-13*ic_cap*ic_cap+-1.25000e-13*ic_cap+2.74000e-11'
+ mcrdll1_cc_w_10_000_s_30_000 = '-5.93750e-14*ic_cap*ic_cap+-3.75000e-14*ic_cap+1.18000e-11'
+ mcrdll1_cc_w_10_000_s_5_000 = '-5.65625e-13*ic_cap*ic_cap+-3.37500e-13*ic_cap+5.09000e-11'
+ mcrdll1_cc_w_10_000_s_8_000 = '-3.18750e-13*ic_cap*ic_cap+-2.00000e-13*ic_cap+3.68000e-11'
+ mcrdll1_cc_w_40_000_s_10_000 = '-2.43750e-13*ic_cap*ic_cap+-1.50000e-13*ic_cap+4.12000e-11'
+ mcrdll1_cc_w_40_000_s_12_000 = '-1.93750e-13*ic_cap*ic_cap+-1.25000e-13*ic_cap+3.68000e-11'
+ mcrdll1_cc_w_40_000_s_30_000 = '-6.25000e-14*ic_cap*ic_cap+-5.00000e-14*ic_cap+1.90000e-11'
+ mcrdll1_cc_w_40_000_s_5_000 = '-5.65625e-13*ic_cap*ic_cap+-3.37500e-13*ic_cap+6.22000e-11'
+ mcrdll1_cc_w_40_000_s_8_000 = '-3.21875e-13*ic_cap*ic_cap+-1.87500e-13*ic_cap+4.72000e-11'
+ mcrdll1_cf_w_10_000_s_10_000 = '-4.37500e-14*ic_cap*ic_cap+-2.50000e-14*ic_cap+1.16000e-11'
+ mcrdll1_cf_w_10_000_s_12_000 = '-5.93750e-14*ic_cap*ic_cap+-3.75000e-14*ic_cap+1.34000e-11'
+ mcrdll1_cf_w_10_000_s_30_000 = '-1.34375e-13*ic_cap*ic_cap+-8.75000e-14*ic_cap+2.38000e-11'
+ mcrdll1_cf_w_10_000_s_5_000 = '1.25000e-15*ic_cap*ic_cap+6.41000e-12'
+ mcrdll1_cf_w_10_000_s_8_000 = '-2.71875e-14*ic_cap*ic_cap+-1.87500e-14*ic_cap+9.67000e-12'
+ mcrdll1_cf_w_40_000_s_10_000 = '-4.06250e-14*ic_cap*ic_cap+-3.75000e-14*ic_cap+1.17000e-11'
+ mcrdll1_cf_w_40_000_s_12_000 = '-5.31250e-14*ic_cap*ic_cap+-3.75000e-14*ic_cap+1.35000e-11'
+ mcrdll1_cf_w_40_000_s_30_000 = '-1.18750e-13*ic_cap*ic_cap+-7.50000e-14*ic_cap+2.45000e-11'
+ mcrdll1_cf_w_40_000_s_5_000 = '1.87500e-15*ic_cap*ic_cap+-2.50000e-15*ic_cap+6.49000e-12'
+ mcrdll1_cf_w_40_000_s_8_000 = '-2.65625e-14*ic_cap*ic_cap+-1.87500e-14*ic_cap+9.76000e-12'
+ mcrdll1d_ca_w_0_170_s_0_180 = '-5.68750e-07*ic_cap*ic_cap+-3.25000e-07*ic_cap+5.80000e-05'
+ mcrdll1d_ca_w_0_170_s_0_225 = '-5.68750e-07*ic_cap*ic_cap+-3.25000e-07*ic_cap+5.80000e-05'
+ mcrdll1d_ca_w_0_170_s_0_270 = '-5.68750e-07*ic_cap*ic_cap+-3.25000e-07*ic_cap+5.80000e-05'
+ mcrdll1d_ca_w_0_170_s_0_360 = '-5.68750e-07*ic_cap*ic_cap+-3.25000e-07*ic_cap+5.80000e-05'
+ mcrdll1d_ca_w_0_170_s_0_450 = '-5.68750e-07*ic_cap*ic_cap+-3.25000e-07*ic_cap+5.80000e-05'
+ mcrdll1d_ca_w_0_170_s_0_540 = '-5.68750e-07*ic_cap*ic_cap+-3.25000e-07*ic_cap+5.80000e-05'
+ mcrdll1d_ca_w_0_170_s_0_720 = '-5.68750e-07*ic_cap*ic_cap+-3.25000e-07*ic_cap+5.80000e-05'
+ mcrdll1d_ca_w_0_170_s_1_080 = '-5.68750e-07*ic_cap*ic_cap+-3.25000e-07*ic_cap+5.80000e-05'
+ mcrdll1d_ca_w_0_170_s_1_980 = '-5.68750e-07*ic_cap*ic_cap+-3.25000e-07*ic_cap+5.80000e-05'
+ mcrdll1d_ca_w_0_170_s_4_500 = '-5.68750e-07*ic_cap*ic_cap+-3.25000e-07*ic_cap+5.80000e-05'
+ mcrdll1d_ca_w_1_360_s_0_180 = '-5.68750e-07*ic_cap*ic_cap+-3.25000e-07*ic_cap+5.80000e-05'
+ mcrdll1d_ca_w_1_360_s_0_225 = '-5.68750e-07*ic_cap*ic_cap+-3.25000e-07*ic_cap+5.80000e-05'
+ mcrdll1d_ca_w_1_360_s_0_270 = '-5.68750e-07*ic_cap*ic_cap+-3.25000e-07*ic_cap+5.80000e-05'
+ mcrdll1d_ca_w_1_360_s_0_360 = '-5.68750e-07*ic_cap*ic_cap+-3.25000e-07*ic_cap+5.80000e-05'
+ mcrdll1d_ca_w_1_360_s_0_450 = '-5.68750e-07*ic_cap*ic_cap+-3.25000e-07*ic_cap+5.80000e-05'
+ mcrdll1d_ca_w_1_360_s_0_540 = '-5.68750e-07*ic_cap*ic_cap+-3.25000e-07*ic_cap+5.80000e-05'
+ mcrdll1d_ca_w_1_360_s_0_720 = '-5.68750e-07*ic_cap*ic_cap+-3.25000e-07*ic_cap+5.80000e-05'
+ mcrdll1d_ca_w_1_360_s_1_080 = '-5.68750e-07*ic_cap*ic_cap+-3.25000e-07*ic_cap+5.80000e-05'
+ mcrdll1d_ca_w_1_360_s_1_980 = '-5.68750e-07*ic_cap*ic_cap+-3.25000e-07*ic_cap+5.80000e-05'
+ mcrdll1d_ca_w_1_360_s_4_500 = '-5.68750e-07*ic_cap*ic_cap+-3.25000e-07*ic_cap+5.80000e-05'
+ mcrdll1d_cc_w_0_170_s_0_180 = '-7.84375e-13*ic_cap*ic_cap+-5.12500e-13*ic_cap+7.71000e-11'
+ mcrdll1d_cc_w_0_170_s_0_225 = '-5.68750e-13*ic_cap*ic_cap+-3.75000e-13*ic_cap+6.53000e-11'
+ mcrdll1d_cc_w_0_170_s_0_270 = '-4.25000e-13*ic_cap*ic_cap+-3.00000e-13*ic_cap+5.73000e-11'
+ mcrdll1d_cc_w_0_170_s_0_360 = '-2.81250e-13*ic_cap*ic_cap+-2.00000e-13*ic_cap+4.60000e-11'
+ mcrdll1d_cc_w_0_170_s_0_450 = '-1.87500e-13*ic_cap*ic_cap+-1.50000e-13*ic_cap+3.89000e-11'
+ mcrdll1d_cc_w_0_170_s_0_540 = '-1.40625e-13*ic_cap*ic_cap+-1.12500e-13*ic_cap+3.32000e-11'
+ mcrdll1d_cc_w_0_170_s_0_720 = '-7.18750e-14*ic_cap*ic_cap+-6.25000e-14*ic_cap+2.56000e-11'
+ mcrdll1d_cc_w_0_170_s_1_080 = '-1.25000e-14*ic_cap*ic_cap+-2.50000e-14*ic_cap+1.67000e-11'
+ mcrdll1d_cc_w_0_170_s_1_980 = '2.12500e-14*ic_cap*ic_cap+7.50000e-15*ic_cap+7.48000e-12'
+ mcrdll1d_cc_w_0_170_s_4_500 = '1.37500e-14*ic_cap*ic_cap+7.50000e-15*ic_cap+1.61000e-12'
+ mcrdll1d_cc_w_1_360_s_0_180 = '-6.93750e-13*ic_cap*ic_cap+-4.50000e-13*ic_cap+9.55000e-11'
+ mcrdll1d_cc_w_1_360_s_0_225 = '-4.81250e-13*ic_cap*ic_cap+-3.25000e-13*ic_cap+8.26000e-11'
+ mcrdll1d_cc_w_1_360_s_0_270 = '-3.43750e-13*ic_cap*ic_cap+-2.50000e-13*ic_cap+7.32000e-11'
+ mcrdll1d_cc_w_1_360_s_0_360 = '-2.06250e-13*ic_cap*ic_cap+-1.50000e-13*ic_cap+6.05000e-11'
+ mcrdll1d_cc_w_1_360_s_0_450 = '-1.25000e-13*ic_cap*ic_cap+-1.00000e-13*ic_cap+5.19000e-11'
+ mcrdll1d_cc_w_1_360_s_0_540 = '-7.50000e-14*ic_cap*ic_cap+-7.50000e-14*ic_cap+4.55000e-11'
+ mcrdll1d_cc_w_1_360_s_0_720 = '-1.87500e-14*ic_cap*ic_cap+-2.50000e-14*ic_cap+3.65000e-11'
+ mcrdll1d_cc_w_1_360_s_1_080 = '3.75000e-14*ic_cap*ic_cap+2.56000e-11'
+ mcrdll1d_cc_w_1_360_s_1_980 = '5.62500e-14*ic_cap*ic_cap+2.50000e-14*ic_cap+1.31000e-11'
+ mcrdll1d_cc_w_1_360_s_4_500 = '3.25000e-14*ic_cap*ic_cap+2.50000e-14*ic_cap+3.58000e-12'
+ mcrdll1d_cf_w_0_170_s_0_180 = '-8.12500e-15*ic_cap*ic_cap+-2.50000e-15*ic_cap+5.08000e-12'
+ mcrdll1d_cf_w_0_170_s_0_225 = '-2.09375e-14*ic_cap*ic_cap+-8.75000e-15*ic_cap+6.29000e-12'
+ mcrdll1d_cf_w_0_170_s_0_270 = '-3.12500e-14*ic_cap*ic_cap+-1.50000e-14*ic_cap+7.44000e-12'
+ mcrdll1d_cf_w_0_170_s_0_360 = '-5.50000e-14*ic_cap*ic_cap+-2.75000e-14*ic_cap+9.92000e-12'
+ mcrdll1d_cf_w_0_170_s_0_450 = '-7.81250e-14*ic_cap*ic_cap+-3.75000e-14*ic_cap+1.19000e-11'
+ mcrdll1d_cf_w_0_170_s_0_540 = '-9.37500e-14*ic_cap*ic_cap+-5.00000e-14*ic_cap+1.41000e-11'
+ mcrdll1d_cf_w_0_170_s_0_720 = '-1.25000e-13*ic_cap*ic_cap+-7.50000e-14*ic_cap+1.77000e-11'
+ mcrdll1d_cf_w_0_170_s_1_080 = '-1.68750e-13*ic_cap*ic_cap+-1.00000e-13*ic_cap+2.34000e-11'
+ mcrdll1d_cf_w_0_170_s_1_980 = '-2.06250e-13*ic_cap*ic_cap+-1.25000e-13*ic_cap+3.09000e-11'
+ mcrdll1d_cf_w_0_170_s_4_500 = '-2.03125e-13*ic_cap*ic_cap+-1.37500e-13*ic_cap+3.64000e-11'
+ mcrdll1d_cf_w_1_360_s_0_180 = '-8.43750e-15*ic_cap*ic_cap+-3.75000e-15*ic_cap+5.08000e-12'
+ mcrdll1d_cf_w_1_360_s_0_225 = '-2.06250e-14*ic_cap*ic_cap+-1.00000e-14*ic_cap+6.29000e-12'
+ mcrdll1d_cf_w_1_360_s_0_270 = '-3.15625e-14*ic_cap*ic_cap+-1.62500e-14*ic_cap+7.47000e-12'
+ mcrdll1d_cf_w_1_360_s_0_360 = '-5.34375e-14*ic_cap*ic_cap+-2.87500e-14*ic_cap+9.77000e-12'
+ mcrdll1d_cf_w_1_360_s_0_450 = '-7.18750e-14*ic_cap*ic_cap+-3.75000e-14*ic_cap+1.19000e-11'
+ mcrdll1d_cf_w_1_360_s_0_540 = '-9.37500e-14*ic_cap*ic_cap+-5.00000e-14*ic_cap+1.40000e-11'
+ mcrdll1d_cf_w_1_360_s_0_720 = '-1.28125e-13*ic_cap*ic_cap+-6.25000e-14*ic_cap+1.78000e-11'
+ mcrdll1d_cf_w_1_360_s_1_080 = '-1.68750e-13*ic_cap*ic_cap+-1.00000e-13*ic_cap+2.39000e-11'
+ mcrdll1d_cf_w_1_360_s_1_980 = '-2.00000e-13*ic_cap*ic_cap+-1.25000e-13*ic_cap+3.34000e-11'
+ mcrdll1d_cf_w_1_360_s_4_500 = '-1.93750e-13*ic_cap*ic_cap+-1.25000e-13*ic_cap+4.22000e-11'
+ mcrdll1f_ca_w_0_170_s_0_180 = '-4.40625e-07*ic_cap*ic_cap+-2.37500e-07*ic_cap+3.97000e-05'
+ mcrdll1f_ca_w_0_170_s_0_225 = '-4.40625e-07*ic_cap*ic_cap+-2.37500e-07*ic_cap+3.97000e-05'
+ mcrdll1f_ca_w_0_170_s_0_270 = '-4.40625e-07*ic_cap*ic_cap+-2.37500e-07*ic_cap+3.97000e-05'
+ mcrdll1f_ca_w_0_170_s_0_360 = '-4.40625e-07*ic_cap*ic_cap+-2.37500e-07*ic_cap+3.97000e-05'
+ mcrdll1f_ca_w_0_170_s_0_450 = '-4.40625e-07*ic_cap*ic_cap+-2.37500e-07*ic_cap+3.97000e-05'
+ mcrdll1f_ca_w_0_170_s_0_540 = '-4.40625e-07*ic_cap*ic_cap+-2.37500e-07*ic_cap+3.97000e-05'
+ mcrdll1f_ca_w_0_170_s_0_720 = '-4.40625e-07*ic_cap*ic_cap+-2.37500e-07*ic_cap+3.97000e-05'
+ mcrdll1f_ca_w_0_170_s_1_080 = '-4.40625e-07*ic_cap*ic_cap+-2.37500e-07*ic_cap+3.97000e-05'
+ mcrdll1f_ca_w_0_170_s_1_980 = '-4.40625e-07*ic_cap*ic_cap+-2.37500e-07*ic_cap+3.97000e-05'
+ mcrdll1f_ca_w_0_170_s_4_500 = '-4.40625e-07*ic_cap*ic_cap+-2.37500e-07*ic_cap+3.97000e-05'
+ mcrdll1f_ca_w_1_360_s_0_180 = '-4.40625e-07*ic_cap*ic_cap+-2.37500e-07*ic_cap+3.97000e-05'
+ mcrdll1f_ca_w_1_360_s_0_225 = '-4.40625e-07*ic_cap*ic_cap+-2.37500e-07*ic_cap+3.97000e-05'
+ mcrdll1f_ca_w_1_360_s_0_270 = '-4.40625e-07*ic_cap*ic_cap+-2.37500e-07*ic_cap+3.97000e-05'
+ mcrdll1f_ca_w_1_360_s_0_360 = '-4.40625e-07*ic_cap*ic_cap+-2.37500e-07*ic_cap+3.97000e-05'
+ mcrdll1f_ca_w_1_360_s_0_450 = '-4.40625e-07*ic_cap*ic_cap+-2.37500e-07*ic_cap+3.97000e-05'
+ mcrdll1f_ca_w_1_360_s_0_540 = '-4.40625e-07*ic_cap*ic_cap+-2.37500e-07*ic_cap+3.97000e-05'
+ mcrdll1f_ca_w_1_360_s_0_720 = '-4.40625e-07*ic_cap*ic_cap+-2.37500e-07*ic_cap+3.97000e-05'
+ mcrdll1f_ca_w_1_360_s_1_080 = '-4.40625e-07*ic_cap*ic_cap+-2.37500e-07*ic_cap+3.97000e-05'
+ mcrdll1f_ca_w_1_360_s_1_980 = '-4.40625e-07*ic_cap*ic_cap+-2.37500e-07*ic_cap+3.97000e-05'
+ mcrdll1f_ca_w_1_360_s_4_500 = '-4.40625e-07*ic_cap*ic_cap+-2.37500e-07*ic_cap+3.97000e-05'
+ mcrdll1f_cc_w_0_170_s_0_180 = '-7.96875e-13*ic_cap*ic_cap+-5.12500e-13*ic_cap+7.95000e-11'
+ mcrdll1f_cc_w_0_170_s_0_225 = '-5.78125e-13*ic_cap*ic_cap+-3.87500e-13*ic_cap+6.78000e-11'
+ mcrdll1f_cc_w_0_170_s_0_270 = '-4.40625e-13*ic_cap*ic_cap+-3.12500e-13*ic_cap+6.01000e-11'
+ mcrdll1f_cc_w_0_170_s_0_360 = '-3.00000e-13*ic_cap*ic_cap+-2.25000e-13*ic_cap+4.91000e-11'
+ mcrdll1f_cc_w_0_170_s_0_450 = '-2.00000e-13*ic_cap*ic_cap+-1.50000e-13*ic_cap+4.22000e-11'
+ mcrdll1f_cc_w_0_170_s_0_540 = '-1.43750e-13*ic_cap*ic_cap+-1.25000e-13*ic_cap+3.66000e-11'
+ mcrdll1f_cc_w_0_170_s_0_720 = '-7.50000e-14*ic_cap*ic_cap+-7.50000e-14*ic_cap+2.92000e-11'
+ mcrdll1f_cc_w_0_170_s_1_080 = '-1.25000e-14*ic_cap*ic_cap+-2.50000e-14*ic_cap+2.03000e-11'
+ mcrdll1f_cc_w_0_170_s_1_980 = '4.06250e-14*ic_cap*ic_cap+1.25000e-14*ic_cap+1.02000e-11'
+ mcrdll1f_cc_w_0_170_s_4_500 = '2.78125e-14*ic_cap*ic_cap+1.62500e-14*ic_cap+2.50000e-12'
+ mcrdll1f_cc_w_1_360_s_0_180 = '-6.84375e-13*ic_cap*ic_cap+-4.37500e-13*ic_cap+1.00000e-10'
+ mcrdll1f_cc_w_1_360_s_0_225 = '-4.65625e-13*ic_cap*ic_cap+-3.12500e-13*ic_cap+8.69000e-11'
+ mcrdll1f_cc_w_1_360_s_0_270 = '-3.31250e-13*ic_cap*ic_cap+-2.25000e-13*ic_cap+7.76000e-11'
+ mcrdll1f_cc_w_1_360_s_0_360 = '-1.90625e-13*ic_cap*ic_cap+-1.37500e-13*ic_cap+6.49000e-11'
+ mcrdll1f_cc_w_1_360_s_0_450 = '-1.09375e-13*ic_cap*ic_cap+-8.75000e-14*ic_cap+5.63000e-11'
+ mcrdll1f_cc_w_1_360_s_0_540 = '-5.31250e-14*ic_cap*ic_cap+-6.25000e-14*ic_cap+4.98000e-11'
+ mcrdll1f_cc_w_1_360_s_0_720 = '4.03897e-28*ic_cap*ic_cap+-2.50000e-14*ic_cap+4.08000e-11'
+ mcrdll1f_cc_w_1_360_s_1_080 = '5.00000e-14*ic_cap*ic_cap+2.50000e-14*ic_cap+2.98000e-11'
+ mcrdll1f_cc_w_1_360_s_1_980 = '8.12500e-14*ic_cap*ic_cap+5.00000e-14*ic_cap+1.63000e-11'
+ mcrdll1f_cc_w_1_360_s_4_500 = '5.43750e-14*ic_cap*ic_cap+3.75000e-14*ic_cap+4.82000e-12'
+ mcrdll1f_cf_w_0_170_s_0_180 = '-1.06250e-14*ic_cap*ic_cap+-5.00000e-15*ic_cap+3.51000e-12'
+ mcrdll1f_cf_w_0_170_s_0_225 = '-2.00000e-14*ic_cap*ic_cap+-1.00000e-14*ic_cap+4.35000e-12'
+ mcrdll1f_cf_w_0_170_s_0_270 = '-2.90625e-14*ic_cap*ic_cap+-1.62500e-14*ic_cap+5.18000e-12'
+ mcrdll1f_cf_w_0_170_s_0_360 = '-4.78125e-14*ic_cap*ic_cap+-2.62500e-14*ic_cap+6.97000e-12'
+ mcrdll1f_cf_w_0_170_s_0_450 = '-6.50000e-14*ic_cap*ic_cap+-3.50000e-14*ic_cap+8.36000e-12'
+ mcrdll1f_cf_w_0_170_s_0_540 = '-8.31250e-14*ic_cap*ic_cap+-4.50000e-14*ic_cap+1.01000e-11'
+ mcrdll1f_cf_w_0_170_s_0_720 = '-1.03125e-13*ic_cap*ic_cap+-6.25000e-14*ic_cap+1.28000e-11'
+ mcrdll1f_cf_w_0_170_s_1_080 = '-1.53125e-13*ic_cap*ic_cap+-8.75000e-14*ic_cap+1.76000e-11'
+ mcrdll1f_cf_w_0_170_s_1_980 = '-2.06250e-13*ic_cap*ic_cap+-1.25000e-13*ic_cap+2.49000e-11'
+ mcrdll1f_cf_w_0_170_s_4_500 = '-2.03125e-13*ic_cap*ic_cap+-1.37500e-13*ic_cap+3.18000e-11'
+ mcrdll1f_cf_w_1_360_s_0_180 = '-1.06250e-14*ic_cap*ic_cap+-5.00000e-15*ic_cap+3.51000e-12'
+ mcrdll1f_cf_w_1_360_s_0_225 = '-2.00000e-14*ic_cap*ic_cap+-1.00000e-14*ic_cap+4.36000e-12'
+ mcrdll1f_cf_w_1_360_s_0_270 = '-2.87500e-14*ic_cap*ic_cap+-1.50000e-14*ic_cap+5.19000e-12'
+ mcrdll1f_cf_w_1_360_s_0_360 = '-4.62500e-14*ic_cap*ic_cap+-2.75000e-14*ic_cap+6.83000e-12'
+ mcrdll1f_cf_w_1_360_s_0_450 = '-6.37500e-14*ic_cap*ic_cap+-3.50000e-14*ic_cap+8.42000e-12'
+ mcrdll1f_cf_w_1_360_s_0_540 = '-7.93750e-14*ic_cap*ic_cap+-4.25000e-14*ic_cap+9.94000e-12'
+ mcrdll1f_cf_w_1_360_s_0_720 = '-1.09375e-13*ic_cap*ic_cap+-6.25000e-14*ic_cap+1.28000e-11'
+ mcrdll1f_cf_w_1_360_s_1_080 = '-1.53125e-13*ic_cap*ic_cap+-8.75000e-14*ic_cap+1.78000e-11'
+ mcrdll1f_cf_w_1_360_s_1_980 = '-2.06250e-13*ic_cap*ic_cap+-1.25000e-13*ic_cap+2.67000e-11'
+ mcrdll1f_cf_w_1_360_s_4_500 = '-2.00000e-13*ic_cap*ic_cap+-1.25000e-13*ic_cap+3.66000e-11'
+ mcrdll1p1_ca_w_0_170_s_0_180 = '-1.67813e-06*ic_cap*ic_cap+-8.12500e-07*ic_cap+9.69000e-05'
+ mcrdll1p1_ca_w_0_170_s_0_225 = '-1.67813e-06*ic_cap*ic_cap+-8.12500e-07*ic_cap+9.69000e-05'
+ mcrdll1p1_ca_w_0_170_s_0_270 = '-1.67813e-06*ic_cap*ic_cap+-8.12500e-07*ic_cap+9.69000e-05'
+ mcrdll1p1_ca_w_0_170_s_0_360 = '-1.67813e-06*ic_cap*ic_cap+-8.12500e-07*ic_cap+9.69000e-05'
+ mcrdll1p1_ca_w_0_170_s_0_450 = '-1.67813e-06*ic_cap*ic_cap+-8.12500e-07*ic_cap+9.69000e-05'
+ mcrdll1p1_ca_w_0_170_s_0_540 = '-1.67813e-06*ic_cap*ic_cap+-8.12500e-07*ic_cap+9.69000e-05'
+ mcrdll1p1_ca_w_0_170_s_0_720 = '-1.67813e-06*ic_cap*ic_cap+-8.12500e-07*ic_cap+9.69000e-05'
+ mcrdll1p1_ca_w_0_170_s_1_080 = '-1.67813e-06*ic_cap*ic_cap+-8.12500e-07*ic_cap+9.69000e-05'
+ mcrdll1p1_ca_w_0_170_s_1_980 = '-1.67813e-06*ic_cap*ic_cap+-8.12500e-07*ic_cap+9.69000e-05'
+ mcrdll1p1_ca_w_0_170_s_4_500 = '-1.67813e-06*ic_cap*ic_cap+-8.12500e-07*ic_cap+9.69000e-05'
+ mcrdll1p1_ca_w_1_360_s_0_180 = '-1.67813e-06*ic_cap*ic_cap+-8.12500e-07*ic_cap+9.69000e-05'
+ mcrdll1p1_ca_w_1_360_s_0_225 = '-1.67813e-06*ic_cap*ic_cap+-8.12500e-07*ic_cap+9.69000e-05'
+ mcrdll1p1_ca_w_1_360_s_0_270 = '-1.67813e-06*ic_cap*ic_cap+-8.12500e-07*ic_cap+9.69000e-05'
+ mcrdll1p1_ca_w_1_360_s_0_360 = '-1.67813e-06*ic_cap*ic_cap+-8.12500e-07*ic_cap+9.69000e-05'
+ mcrdll1p1_ca_w_1_360_s_0_450 = '-1.67813e-06*ic_cap*ic_cap+-8.12500e-07*ic_cap+9.69000e-05'
+ mcrdll1p1_ca_w_1_360_s_0_540 = '-1.67813e-06*ic_cap*ic_cap+-8.12500e-07*ic_cap+9.69000e-05'
+ mcrdll1p1_ca_w_1_360_s_0_720 = '-1.67813e-06*ic_cap*ic_cap+-8.12500e-07*ic_cap+9.69000e-05'
+ mcrdll1p1_ca_w_1_360_s_1_080 = '-1.67813e-06*ic_cap*ic_cap+-8.12500e-07*ic_cap+9.69000e-05'
+ mcrdll1p1_ca_w_1_360_s_1_980 = '-1.67813e-06*ic_cap*ic_cap+-8.12500e-07*ic_cap+9.69000e-05'
+ mcrdll1p1_ca_w_1_360_s_4_500 = '-1.67813e-06*ic_cap*ic_cap+-8.12500e-07*ic_cap+9.69000e-05'
+ mcrdll1p1_cc_w_0_170_s_0_180 = '-6.81250e-13*ic_cap*ic_cap+-4.75000e-13*ic_cap+7.29000e-11'
+ mcrdll1p1_cc_w_0_170_s_0_225 = '-4.62500e-13*ic_cap*ic_cap+-3.25000e-13*ic_cap+6.09000e-11'
+ mcrdll1p1_cc_w_0_170_s_0_270 = '-3.18750e-13*ic_cap*ic_cap+-2.50000e-13*ic_cap+5.27000e-11'
+ mcrdll1p1_cc_w_0_170_s_0_360 = '-1.68750e-13*ic_cap*ic_cap+-1.50000e-13*ic_cap+4.10000e-11'
+ mcrdll1p1_cc_w_0_170_s_0_450 = '-8.12500e-14*ic_cap*ic_cap+-1.00000e-13*ic_cap+3.39000e-11'
+ mcrdll1p1_cc_w_0_170_s_0_540 = '-2.81250e-14*ic_cap*ic_cap+-6.25000e-14*ic_cap+2.80000e-11'
+ mcrdll1p1_cc_w_0_170_s_0_720 = '3.12500e-14*ic_cap*ic_cap+-2.50000e-14*ic_cap+2.05000e-11'
+ mcrdll1p1_cc_w_0_170_s_1_080 = '7.18750e-14*ic_cap*ic_cap+1.25000e-14*ic_cap+1.21000e-11'
+ mcrdll1p1_cc_w_0_170_s_1_980 = '5.62500e-14*ic_cap*ic_cap+2.50000e-14*ic_cap+4.79000e-12'
+ mcrdll1p1_cc_w_0_170_s_4_500 = '1.65000e-14*ic_cap*ic_cap+8.75000e-15*ic_cap+9.61000e-13'
+ mcrdll1p1_cc_w_1_360_s_0_180 = '-5.90625e-13*ic_cap*ic_cap+-3.87500e-13*ic_cap+8.97000e-11'
+ mcrdll1p1_cc_w_1_360_s_0_225 = '-3.65625e-13*ic_cap*ic_cap+-2.62500e-13*ic_cap+7.67000e-11'
+ mcrdll1p1_cc_w_1_360_s_0_270 = '-2.40625e-13*ic_cap*ic_cap+-1.87500e-13*ic_cap+6.74000e-11'
+ mcrdll1p1_cc_w_1_360_s_0_360 = '-9.37500e-14*ic_cap*ic_cap+-1.00000e-13*ic_cap+5.46000e-11'
+ mcrdll1p1_cc_w_1_360_s_0_450 = '-1.87500e-14*ic_cap*ic_cap+-5.00000e-14*ic_cap+4.61000e-11'
+ mcrdll1p1_cc_w_1_360_s_0_540 = '2.81250e-14*ic_cap*ic_cap+-1.25000e-14*ic_cap+3.98000e-11'
+ mcrdll1p1_cc_w_1_360_s_0_720 = '7.50000e-14*ic_cap*ic_cap+2.50000e-14*ic_cap+3.11000e-11'
+ mcrdll1p1_cc_w_1_360_s_1_080 = '1.06250e-13*ic_cap*ic_cap+5.00000e-14*ic_cap+2.09000e-11'
+ mcrdll1p1_cc_w_1_360_s_1_980 = '9.00000e-14*ic_cap*ic_cap+6.25000e-14*ic_cap+9.91000e-12'
+ mcrdll1p1_cc_w_1_360_s_4_500 = '3.53125e-14*ic_cap*ic_cap+3.12500e-14*ic_cap+2.56000e-12'
+ mcrdll1p1_cf_w_0_170_s_0_180 = '-8.21875e-14*ic_cap*ic_cap+-3.87500e-14*ic_cap+8.32000e-12'
+ mcrdll1p1_cf_w_0_170_s_0_225 = '-1.13125e-13*ic_cap*ic_cap+-5.50000e-14*ic_cap+1.02000e-11'
+ mcrdll1p1_cf_w_0_170_s_0_270 = '-1.41563e-13*ic_cap*ic_cap+-6.62500e-14*ic_cap+1.20000e-11'
+ mcrdll1p1_cf_w_0_170_s_0_360 = '-2.06250e-13*ic_cap*ic_cap+-1.00000e-13*ic_cap+1.58000e-11'
+ mcrdll1p1_cf_w_0_170_s_0_450 = '-2.43750e-13*ic_cap*ic_cap+-1.25000e-13*ic_cap+1.86000e-11'
+ mcrdll1p1_cf_w_0_170_s_0_540 = '-2.84375e-13*ic_cap*ic_cap+-1.37500e-13*ic_cap+2.17000e-11'
+ mcrdll1p1_cf_w_0_170_s_0_720 = '-3.37500e-13*ic_cap*ic_cap+-1.75000e-13*ic_cap+2.64000e-11'
+ mcrdll1p1_cf_w_0_170_s_1_080 = '-3.90625e-13*ic_cap*ic_cap+-2.12500e-13*ic_cap+3.28000e-11'
+ mcrdll1p1_cf_w_0_170_s_1_980 = '-3.93750e-13*ic_cap*ic_cap+-2.25000e-13*ic_cap+3.95000e-11'
+ mcrdll1p1_cf_w_0_170_s_4_500 = '-3.59375e-13*ic_cap*ic_cap+-2.12500e-13*ic_cap+4.32000e-11'
+ mcrdll1p1_cf_w_1_360_s_0_180 = '-8.43750e-14*ic_cap*ic_cap+-3.75000e-14*ic_cap+8.41000e-12'
+ mcrdll1p1_cf_w_1_360_s_0_225 = '-1.14375e-13*ic_cap*ic_cap+-5.25000e-14*ic_cap+1.03000e-11'
+ mcrdll1p1_cf_w_1_360_s_0_270 = '-1.47812e-13*ic_cap*ic_cap+-6.62500e-14*ic_cap+1.22000e-11'
+ mcrdll1p1_cf_w_1_360_s_0_360 = '-1.96875e-13*ic_cap*ic_cap+-8.75000e-14*ic_cap+1.56000e-11'
+ mcrdll1p1_cf_w_1_360_s_0_450 = '-2.43750e-13*ic_cap*ic_cap+-1.25000e-13*ic_cap+1.88000e-11'
+ mcrdll1p1_cf_w_1_360_s_0_540 = '-2.81250e-13*ic_cap*ic_cap+-1.50000e-13*ic_cap+2.17000e-11'
+ mcrdll1p1_cf_w_1_360_s_0_720 = '-3.43750e-13*ic_cap*ic_cap+-1.75000e-13*ic_cap+2.67000e-11'
+ mcrdll1p1_cf_w_1_360_s_1_080 = '-3.96875e-13*ic_cap*ic_cap+-2.12500e-13*ic_cap+3.39000e-11'
+ mcrdll1p1_cf_w_1_360_s_1_980 = '-4.15625e-13*ic_cap*ic_cap+-2.37500e-13*ic_cap+4.34000e-11'
+ mcrdll1p1_cf_w_1_360_s_4_500 = '-3.71875e-13*ic_cap*ic_cap+-2.12500e-13*ic_cap+5.04000e-11'
+ mcrdlm1_ca_w_10_000_s_10_000 = '-2.56250e-08*ic_cap*ic_cap+-1.50000e-08*ic_cap+2.93000e-06'
+ mcrdlm1_ca_w_10_000_s_12_000 = '-2.56250e-08*ic_cap*ic_cap+-1.50000e-08*ic_cap+2.93000e-06'
+ mcrdlm1_ca_w_10_000_s_30_000 = '-2.56250e-08*ic_cap*ic_cap+-1.50000e-08*ic_cap+2.93000e-06'
+ mcrdlm1_ca_w_10_000_s_5_000 = '-2.56250e-08*ic_cap*ic_cap+-1.50000e-08*ic_cap+2.93000e-06'
+ mcrdlm1_ca_w_10_000_s_8_000 = '-2.56250e-08*ic_cap*ic_cap+-1.50000e-08*ic_cap+2.93000e-06'
+ mcrdlm1_ca_w_40_000_s_10_000 = '-2.56250e-08*ic_cap*ic_cap+-1.50000e-08*ic_cap+2.93000e-06'
+ mcrdlm1_ca_w_40_000_s_12_000 = '-2.56250e-08*ic_cap*ic_cap+-1.50000e-08*ic_cap+2.93000e-06'
+ mcrdlm1_ca_w_40_000_s_30_000 = '-2.56250e-08*ic_cap*ic_cap+-1.50000e-08*ic_cap+2.93000e-06'
+ mcrdlm1_ca_w_40_000_s_5_000 = '-2.56250e-08*ic_cap*ic_cap+-1.50000e-08*ic_cap+2.93000e-06'
+ mcrdlm1_ca_w_40_000_s_8_000 = '-2.56250e-08*ic_cap*ic_cap+-1.50000e-08*ic_cap+2.93000e-06'
+ mcrdlm1_cc_w_10_000_s_10_000 = '-2.40625e-13*ic_cap*ic_cap+-1.62500e-13*ic_cap+3.09000e-11'
+ mcrdlm1_cc_w_10_000_s_12_000 = '-1.93750e-13*ic_cap*ic_cap+-1.25000e-13*ic_cap+2.69000e-11'
+ mcrdlm1_cc_w_10_000_s_30_000 = '-5.93750e-14*ic_cap*ic_cap+-3.75000e-14*ic_cap+1.15000e-11'
+ mcrdlm1_cc_w_10_000_s_5_000 = '-5.59375e-13*ic_cap*ic_cap+-3.37500e-13*ic_cap+5.04000e-11'
+ mcrdlm1_cc_w_10_000_s_8_000 = '-3.12500e-13*ic_cap*ic_cap+-2.00000e-13*ic_cap+3.63000e-11'
+ mcrdlm1_cc_w_40_000_s_10_000 = '-2.50000e-13*ic_cap*ic_cap+-1.50000e-13*ic_cap+4.08000e-11'
+ mcrdlm1_cc_w_40_000_s_12_000 = '-2.00000e-13*ic_cap*ic_cap+-1.25000e-13*ic_cap+3.64000e-11'
+ mcrdlm1_cc_w_40_000_s_30_000 = '-5.93750e-14*ic_cap*ic_cap+-3.75000e-14*ic_cap+1.86000e-11'
+ mcrdlm1_cc_w_40_000_s_5_000 = '-5.65625e-13*ic_cap*ic_cap+-3.37500e-13*ic_cap+6.17000e-11'
+ mcrdlm1_cc_w_40_000_s_8_000 = '-3.18750e-13*ic_cap*ic_cap+-2.00000e-13*ic_cap+4.67000e-11'
+ mcrdlm1_cf_w_10_000_s_10_000 = '-4.37500e-14*ic_cap*ic_cap+-2.50000e-14*ic_cap+1.21000e-11'
+ mcrdlm1_cf_w_10_000_s_12_000 = '-5.93750e-14*ic_cap*ic_cap+-3.75000e-14*ic_cap+1.40000e-11'
+ mcrdlm1_cf_w_10_000_s_30_000 = '-1.34375e-13*ic_cap*ic_cap+-8.75000e-14*ic_cap+2.45000e-11'
+ mcrdlm1_cf_w_10_000_s_5_000 = '1.25000e-15*ic_cap*ic_cap+6.73000e-12'
+ mcrdlm1_cf_w_10_000_s_8_000 = '-2.71875e-14*ic_cap*ic_cap+-1.87500e-14*ic_cap+1.01000e-11'
+ mcrdlm1_cf_w_40_000_s_10_000 = '-4.37500e-14*ic_cap*ic_cap+-2.50000e-14*ic_cap+1.22000e-11'
+ mcrdlm1_cf_w_40_000_s_12_000 = '-5.93750e-14*ic_cap*ic_cap+-3.75000e-14*ic_cap+1.41000e-11'
+ mcrdlm1_cf_w_40_000_s_30_000 = '-1.28125e-13*ic_cap*ic_cap+-8.75000e-14*ic_cap+2.53000e-11'
+ mcrdlm1_cf_w_40_000_s_5_000 = '3.12500e-16*ic_cap*ic_cap+-1.25000e-15*ic_cap+6.82000e-12'
+ mcrdlm1_cf_w_40_000_s_8_000 = '-2.78125e-14*ic_cap*ic_cap+-2.12500e-14*ic_cap+1.02000e-11'
+ mcrdlm1d_ca_w_0_140_s_0_140 = '-3.96875e-07*ic_cap*ic_cap+-2.62500e-07*ic_cap+3.65000e-05'
+ mcrdlm1d_ca_w_0_140_s_0_175 = '-3.96875e-07*ic_cap*ic_cap+-2.62500e-07*ic_cap+3.65000e-05'
+ mcrdlm1d_ca_w_0_140_s_0_210 = '-3.96875e-07*ic_cap*ic_cap+-2.62500e-07*ic_cap+3.65000e-05'
+ mcrdlm1d_ca_w_0_140_s_0_280 = '-3.96875e-07*ic_cap*ic_cap+-2.62500e-07*ic_cap+3.65000e-05'
+ mcrdlm1d_ca_w_0_140_s_0_350 = '-3.96875e-07*ic_cap*ic_cap+-2.62500e-07*ic_cap+3.65000e-05'
+ mcrdlm1d_ca_w_0_140_s_0_420 = '-3.96875e-07*ic_cap*ic_cap+-2.62500e-07*ic_cap+3.65000e-05'
+ mcrdlm1d_ca_w_0_140_s_0_560 = '-3.96875e-07*ic_cap*ic_cap+-2.62500e-07*ic_cap+3.65000e-05'
+ mcrdlm1d_ca_w_0_140_s_0_840 = '-3.96875e-07*ic_cap*ic_cap+-2.62500e-07*ic_cap+3.65000e-05'
+ mcrdlm1d_ca_w_0_140_s_1_540 = '-3.96875e-07*ic_cap*ic_cap+-2.62500e-07*ic_cap+3.65000e-05'
+ mcrdlm1d_ca_w_0_140_s_3_500 = '-3.96875e-07*ic_cap*ic_cap+-2.62500e-07*ic_cap+3.65000e-05'
+ mcrdlm1d_ca_w_1_120_s_0_140 = '-3.96875e-07*ic_cap*ic_cap+-2.62500e-07*ic_cap+3.65000e-05'
+ mcrdlm1d_ca_w_1_120_s_0_175 = '-3.96875e-07*ic_cap*ic_cap+-2.62500e-07*ic_cap+3.65000e-05'
+ mcrdlm1d_ca_w_1_120_s_0_210 = '-3.96875e-07*ic_cap*ic_cap+-2.62500e-07*ic_cap+3.65000e-05'
+ mcrdlm1d_ca_w_1_120_s_0_280 = '-3.96875e-07*ic_cap*ic_cap+-2.62500e-07*ic_cap+3.65000e-05'
+ mcrdlm1d_ca_w_1_120_s_0_350 = '-3.96875e-07*ic_cap*ic_cap+-2.62500e-07*ic_cap+3.65000e-05'
+ mcrdlm1d_ca_w_1_120_s_0_420 = '-3.96875e-07*ic_cap*ic_cap+-2.62500e-07*ic_cap+3.65000e-05'
+ mcrdlm1d_ca_w_1_120_s_0_560 = '-3.96875e-07*ic_cap*ic_cap+-2.62500e-07*ic_cap+3.65000e-05'
+ mcrdlm1d_ca_w_1_120_s_0_840 = '-3.96875e-07*ic_cap*ic_cap+-2.62500e-07*ic_cap+3.65000e-05'
+ mcrdlm1d_ca_w_1_120_s_1_540 = '-3.96875e-07*ic_cap*ic_cap+-2.62500e-07*ic_cap+3.65000e-05'
+ mcrdlm1d_ca_w_1_120_s_3_500 = '-3.96875e-07*ic_cap*ic_cap+-2.62500e-07*ic_cap+3.65000e-05'
+ mcrdlm1d_cc_w_0_140_s_0_140 = '-9.28125e-13*ic_cap*ic_cap+-5.12500e-13*ic_cap+1.04000e-10'
+ mcrdlm1d_cc_w_0_140_s_0_175 = '-8.96875e-13*ic_cap*ic_cap+-5.37500e-13*ic_cap+1.02000e-10'
+ mcrdlm1d_cc_w_0_140_s_0_210 = '-7.81250e-13*ic_cap*ic_cap+-4.00000e-13*ic_cap+9.66000e-11'
+ mcrdlm1d_cc_w_0_140_s_0_280 = '-5.78125e-13*ic_cap*ic_cap+-3.62500e-13*ic_cap+8.55000e-11'
+ mcrdlm1d_cc_w_0_140_s_0_350 = '-4.46875e-13*ic_cap*ic_cap+-2.62500e-13*ic_cap+7.40000e-11'
+ mcrdlm1d_cc_w_0_140_s_0_420 = '-3.53125e-13*ic_cap*ic_cap+-2.12500e-13*ic_cap+6.49000e-11'
+ mcrdlm1d_cc_w_0_140_s_0_560 = '-1.93750e-13*ic_cap*ic_cap+-1.25000e-13*ic_cap+5.17000e-11'
+ mcrdlm1d_cc_w_0_140_s_0_840 = '-6.87500e-14*ic_cap*ic_cap+-5.00000e-14*ic_cap+3.72000e-11'
+ mcrdlm1d_cc_w_0_140_s_1_540 = '1.56250e-14*ic_cap*ic_cap+1.25000e-14*ic_cap+2.08000e-11'
+ mcrdlm1d_cc_w_0_140_s_3_500 = '4.81250e-14*ic_cap*ic_cap+3.25000e-14*ic_cap+6.54000e-12'
+ mcrdlm1d_cc_w_1_120_s_0_140 = '-7.81250e-13*ic_cap*ic_cap+-3.75000e-13*ic_cap+1.26000e-10'
+ mcrdlm1d_cc_w_1_120_s_0_175 = '-7.81250e-13*ic_cap*ic_cap+-3.75000e-13*ic_cap+1.23000e-10'
+ mcrdlm1d_cc_w_1_120_s_0_210 = '-5.93750e-13*ic_cap*ic_cap+-3.75000e-13*ic_cap+1.16000e-10'
+ mcrdlm1d_cc_w_1_120_s_0_280 = '-5.21875e-13*ic_cap*ic_cap+-3.87500e-13*ic_cap+1.03000e-10'
+ mcrdlm1d_cc_w_1_120_s_0_350 = '-3.78125e-13*ic_cap*ic_cap+-2.12500e-13*ic_cap+9.03000e-11'
+ mcrdlm1d_cc_w_1_120_s_0_420 = '-2.84375e-13*ic_cap*ic_cap+-1.87500e-13*ic_cap+7.95000e-11'
+ mcrdlm1d_cc_w_1_120_s_0_560 = '-1.31250e-13*ic_cap*ic_cap+-7.50000e-14*ic_cap+6.41000e-11'
+ mcrdlm1d_cc_w_1_120_s_0_840 = '-2.18750e-14*ic_cap*ic_cap+-1.25000e-14*ic_cap+4.68000e-11'
+ mcrdlm1d_cc_w_1_120_s_1_540 = '6.25000e-14*ic_cap*ic_cap+5.00000e-14*ic_cap+2.72000e-11'
+ mcrdlm1d_cc_w_1_120_s_3_500 = '7.12500e-14*ic_cap*ic_cap+5.00000e-14*ic_cap+9.66000e-12'
+ mcrdlm1d_cf_w_0_140_s_0_140 = '-3.75000e-15*ic_cap*ic_cap+-5.00000e-15*ic_cap+2.53000e-12'
+ mcrdlm1d_cf_w_0_140_s_0_175 = '-1.03125e-14*ic_cap*ic_cap+-8.75000e-15*ic_cap+3.16000e-12'
+ mcrdlm1d_cf_w_0_140_s_0_210 = '-1.71875e-14*ic_cap*ic_cap+-1.37500e-14*ic_cap+3.80000e-12'
+ mcrdlm1d_cf_w_0_140_s_0_280 = '-3.09375e-14*ic_cap*ic_cap+-2.12500e-14*ic_cap+5.04000e-12'
+ mcrdlm1d_cf_w_0_140_s_0_350 = '-4.43750e-14*ic_cap*ic_cap+-3.00000e-14*ic_cap+6.25000e-12'
+ mcrdlm1d_cf_w_0_140_s_0_420 = '-5.81250e-14*ic_cap*ic_cap+-3.75000e-14*ic_cap+7.49000e-12'
+ mcrdlm1d_cf_w_0_140_s_0_560 = '-8.06250e-14*ic_cap*ic_cap+-5.50000e-14*ic_cap+9.74000e-12'
+ mcrdlm1d_cf_w_0_140_s_0_840 = '-1.25000e-13*ic_cap*ic_cap+-7.50000e-14*ic_cap+1.39000e-11'
+ mcrdlm1d_cf_w_0_140_s_1_540 = '-1.93750e-13*ic_cap*ic_cap+-1.25000e-13*ic_cap+2.22000e-11'
+ mcrdlm1d_cf_w_0_140_s_3_500 = '-2.28125e-13*ic_cap*ic_cap+-1.62500e-13*ic_cap+3.32000e-11'
+ mcrdlm1d_cf_w_1_120_s_0_140 = '-5.62500e-15*ic_cap*ic_cap+-5.00000e-15*ic_cap+2.61000e-12'
+ mcrdlm1d_cf_w_1_120_s_0_175 = '-1.18750e-14*ic_cap*ic_cap+-1.00000e-14*ic_cap+3.24000e-12'
+ mcrdlm1d_cf_w_1_120_s_0_210 = '-1.90625e-14*ic_cap*ic_cap+-1.37500e-14*ic_cap+3.87000e-12'
+ mcrdlm1d_cf_w_1_120_s_0_280 = '-3.25000e-14*ic_cap*ic_cap+-2.25000e-14*ic_cap+5.12000e-12'
+ mcrdlm1d_cf_w_1_120_s_0_350 = '-4.59375e-14*ic_cap*ic_cap+-3.12500e-14*ic_cap+6.34000e-12'
+ mcrdlm1d_cf_w_1_120_s_0_420 = '-5.81250e-14*ic_cap*ic_cap+-4.00000e-14*ic_cap+7.53000e-12'
+ mcrdlm1d_cf_w_1_120_s_0_560 = '-8.21875e-14*ic_cap*ic_cap+-5.62500e-14*ic_cap+9.83000e-12'
+ mcrdlm1d_cf_w_1_120_s_0_840 = '-1.25000e-13*ic_cap*ic_cap+-7.50000e-14*ic_cap+1.41000e-11'
+ mcrdlm1d_cf_w_1_120_s_1_540 = '-1.90625e-13*ic_cap*ic_cap+-1.37500e-13*ic_cap+2.27000e-11'
+ mcrdlm1d_cf_w_1_120_s_3_500 = '-2.37500e-13*ic_cap*ic_cap+-1.75000e-13*ic_cap+3.56000e-11'
+ mcrdlm1f_ca_w_0_140_s_0_140 = '-3.25000e-07*ic_cap*ic_cap+-2.00000e-07*ic_cap+2.87000e-05'
+ mcrdlm1f_ca_w_0_140_s_0_175 = '-3.25000e-07*ic_cap*ic_cap+-2.00000e-07*ic_cap+2.87000e-05'
+ mcrdlm1f_ca_w_0_140_s_0_210 = '-3.25000e-07*ic_cap*ic_cap+-2.00000e-07*ic_cap+2.87000e-05'
+ mcrdlm1f_ca_w_0_140_s_0_280 = '-3.25000e-07*ic_cap*ic_cap+-2.00000e-07*ic_cap+2.87000e-05'
+ mcrdlm1f_ca_w_0_140_s_0_350 = '-3.25000e-07*ic_cap*ic_cap+-2.00000e-07*ic_cap+2.87000e-05'
+ mcrdlm1f_ca_w_0_140_s_0_420 = '-3.25000e-07*ic_cap*ic_cap+-2.00000e-07*ic_cap+2.87000e-05'
+ mcrdlm1f_ca_w_0_140_s_0_560 = '-3.25000e-07*ic_cap*ic_cap+-2.00000e-07*ic_cap+2.87000e-05'
+ mcrdlm1f_ca_w_0_140_s_0_840 = '-3.25000e-07*ic_cap*ic_cap+-2.00000e-07*ic_cap+2.87000e-05'
+ mcrdlm1f_ca_w_0_140_s_1_540 = '-3.25000e-07*ic_cap*ic_cap+-2.00000e-07*ic_cap+2.87000e-05'
+ mcrdlm1f_ca_w_0_140_s_3_500 = '-3.25000e-07*ic_cap*ic_cap+-2.00000e-07*ic_cap+2.87000e-05'
+ mcrdlm1f_ca_w_1_120_s_0_140 = '-3.25000e-07*ic_cap*ic_cap+-2.00000e-07*ic_cap+2.87000e-05'
+ mcrdlm1f_ca_w_1_120_s_0_175 = '-3.25000e-07*ic_cap*ic_cap+-2.00000e-07*ic_cap+2.87000e-05'
+ mcrdlm1f_ca_w_1_120_s_0_210 = '-3.25000e-07*ic_cap*ic_cap+-2.00000e-07*ic_cap+2.87000e-05'
+ mcrdlm1f_ca_w_1_120_s_0_280 = '-3.25000e-07*ic_cap*ic_cap+-2.00000e-07*ic_cap+2.87000e-05'
+ mcrdlm1f_ca_w_1_120_s_0_350 = '-3.25000e-07*ic_cap*ic_cap+-2.00000e-07*ic_cap+2.87000e-05'
+ mcrdlm1f_ca_w_1_120_s_0_420 = '-3.25000e-07*ic_cap*ic_cap+-2.00000e-07*ic_cap+2.87000e-05'
+ mcrdlm1f_ca_w_1_120_s_0_560 = '-3.25000e-07*ic_cap*ic_cap+-2.00000e-07*ic_cap+2.87000e-05'
+ mcrdlm1f_ca_w_1_120_s_0_840 = '-3.25000e-07*ic_cap*ic_cap+-2.00000e-07*ic_cap+2.87000e-05'
+ mcrdlm1f_ca_w_1_120_s_1_540 = '-3.25000e-07*ic_cap*ic_cap+-2.00000e-07*ic_cap+2.87000e-05'
+ mcrdlm1f_ca_w_1_120_s_3_500 = '-3.25000e-07*ic_cap*ic_cap+-2.00000e-07*ic_cap+2.87000e-05'
+ mcrdlm1f_cc_w_0_140_s_0_140 = '-9.43750e-13*ic_cap*ic_cap+-5.25000e-13*ic_cap+1.05000e-10'
+ mcrdlm1f_cc_w_0_140_s_0_175 = '-8.96875e-13*ic_cap*ic_cap+-5.12500e-13*ic_cap+1.03000e-10'
+ mcrdlm1f_cc_w_0_140_s_0_210 = '-7.90625e-13*ic_cap*ic_cap+-4.12500e-13*ic_cap+9.77000e-11'
+ mcrdlm1f_cc_w_0_140_s_0_280 = '-5.84375e-13*ic_cap*ic_cap+-3.37500e-13*ic_cap+8.68000e-11'
+ mcrdlm1f_cc_w_0_140_s_0_350 = '-4.56250e-13*ic_cap*ic_cap+-2.75000e-13*ic_cap+7.54000e-11'
+ mcrdlm1f_cc_w_0_140_s_0_420 = '-3.65625e-13*ic_cap*ic_cap+-2.37500e-13*ic_cap+6.65000e-11'
+ mcrdlm1f_cc_w_0_140_s_0_560 = '-2.09375e-13*ic_cap*ic_cap+-1.37500e-13*ic_cap+5.36000e-11'
+ mcrdlm1f_cc_w_0_140_s_0_840 = '-9.06250e-14*ic_cap*ic_cap+-6.25000e-14*ic_cap+3.94000e-11'
+ mcrdlm1f_cc_w_0_140_s_1_540 = '2.18750e-14*ic_cap*ic_cap+1.25000e-14*ic_cap+2.30000e-11'
+ mcrdlm1f_cc_w_0_140_s_3_500 = '6.12500e-14*ic_cap*ic_cap+3.75000e-14*ic_cap+8.05000e-12'
+ mcrdlm1f_cc_w_1_120_s_0_140 = '-8.12500e-13*ic_cap*ic_cap+-5.00000e-13*ic_cap+1.29000e-10'
+ mcrdlm1f_cc_w_1_120_s_0_175 = '-7.50000e-13*ic_cap*ic_cap+-2.50000e-13*ic_cap+1.25000e-10'
+ mcrdlm1f_cc_w_1_120_s_0_210 = '-6.25000e-13*ic_cap*ic_cap+-5.00000e-13*ic_cap+1.19000e-10'
+ mcrdlm1f_cc_w_1_120_s_0_280 = '-4.78125e-13*ic_cap*ic_cap+-3.87500e-13*ic_cap+1.05000e-10'
+ mcrdlm1f_cc_w_1_120_s_0_350 = '-3.84375e-13*ic_cap*ic_cap+-2.37500e-13*ic_cap+9.30000e-11'
+ mcrdlm1f_cc_w_1_120_s_0_420 = '-2.65625e-13*ic_cap*ic_cap+-2.12500e-13*ic_cap+8.20000e-11'
+ mcrdlm1f_cc_w_1_120_s_0_560 = '-1.31250e-13*ic_cap*ic_cap+-1.00000e-13*ic_cap+6.69000e-11'
+ mcrdlm1f_cc_w_1_120_s_0_840 = '-2.18750e-14*ic_cap*ic_cap+-1.25000e-14*ic_cap+4.96000e-11'
+ mcrdlm1f_cc_w_1_120_s_1_540 = '7.18750e-14*ic_cap*ic_cap+3.75000e-14*ic_cap+2.99000e-11'
+ mcrdlm1f_cc_w_1_120_s_3_500 = '9.06250e-14*ic_cap*ic_cap+6.25000e-14*ic_cap+1.14000e-11'
+ mcrdlm1f_cf_w_0_140_s_0_140 = '-4.37500e-15*ic_cap*ic_cap+-2.50000e-15*ic_cap+2.00000e-12'
+ mcrdlm1f_cf_w_0_140_s_0_175 = '-9.68750e-15*ic_cap*ic_cap+-6.25000e-15*ic_cap+2.49000e-12'
+ mcrdlm1f_cf_w_0_140_s_0_210 = '-1.53125e-14*ic_cap*ic_cap+-1.12500e-14*ic_cap+3.00000e-12'
+ mcrdlm1f_cf_w_0_140_s_0_280 = '-2.68750e-14*ic_cap*ic_cap+-1.75000e-14*ic_cap+3.98000e-12'
+ mcrdlm1f_cf_w_0_140_s_0_350 = '-3.78125e-14*ic_cap*ic_cap+-2.37500e-14*ic_cap+4.94000e-12'
+ mcrdlm1f_cf_w_0_140_s_0_420 = '-4.93750e-14*ic_cap*ic_cap+-3.00000e-14*ic_cap+5.94000e-12'
+ mcrdlm1f_cf_w_0_140_s_0_560 = '-6.90625e-14*ic_cap*ic_cap+-4.62500e-14*ic_cap+7.76000e-12'
+ mcrdlm1f_cf_w_0_140_s_0_840 = '-1.07188e-13*ic_cap*ic_cap+-6.62500e-14*ic_cap+1.12000e-11'
+ mcrdlm1f_cf_w_0_140_s_1_540 = '-1.71875e-13*ic_cap*ic_cap+-1.12500e-13*ic_cap+1.83000e-11'
+ mcrdlm1f_cf_w_0_140_s_3_500 = '-2.28125e-13*ic_cap*ic_cap+-1.62500e-13*ic_cap+2.92000e-11'
+ mcrdlm1f_cf_w_1_120_s_0_140 = '-4.68750e-15*ic_cap*ic_cap+-3.75000e-15*ic_cap+2.04000e-12'
+ mcrdlm1f_cf_w_1_120_s_0_175 = '-1.03125e-14*ic_cap*ic_cap+-6.25000e-15*ic_cap+2.54000e-12'
+ mcrdlm1f_cf_w_1_120_s_0_210 = '-1.65625e-14*ic_cap*ic_cap+-1.12500e-14*ic_cap+3.04000e-12'
+ mcrdlm1f_cf_w_1_120_s_0_280 = '-2.75000e-14*ic_cap*ic_cap+-1.75000e-14*ic_cap+4.03000e-12'
+ mcrdlm1f_cf_w_1_120_s_0_350 = '-3.84375e-14*ic_cap*ic_cap+-2.37500e-14*ic_cap+5.00000e-12'
+ mcrdlm1f_cf_w_1_120_s_0_420 = '-4.87500e-14*ic_cap*ic_cap+-3.00000e-14*ic_cap+5.95000e-12'
+ mcrdlm1f_cf_w_1_120_s_0_560 = '-7.00000e-14*ic_cap*ic_cap+-4.50000e-14*ic_cap+7.81000e-12'
+ mcrdlm1f_cf_w_1_120_s_0_840 = '-1.06563e-13*ic_cap*ic_cap+-6.62500e-14*ic_cap+1.13000e-11'
+ mcrdlm1f_cf_w_1_120_s_1_540 = '-1.78125e-13*ic_cap*ic_cap+-1.12500e-13*ic_cap+1.88000e-11'
+ mcrdlm1f_cf_w_1_120_s_3_500 = '-2.37500e-13*ic_cap*ic_cap+-1.50000e-13*ic_cap+3.12000e-11'
+ mcrdlm1l1_ca_w_0_140_s_0_140 = '-2.01250e-06*ic_cap*ic_cap+-1.27500e-06*ic_cap+1.17000e-04'
+ mcrdlm1l1_ca_w_0_140_s_0_175 = '-2.01250e-06*ic_cap*ic_cap+-1.27500e-06*ic_cap+1.17000e-04'
+ mcrdlm1l1_ca_w_0_140_s_0_210 = '-2.01250e-06*ic_cap*ic_cap+-1.27500e-06*ic_cap+1.17000e-04'
+ mcrdlm1l1_ca_w_0_140_s_0_280 = '-2.01250e-06*ic_cap*ic_cap+-1.27500e-06*ic_cap+1.17000e-04'
+ mcrdlm1l1_ca_w_0_140_s_0_350 = '-2.01250e-06*ic_cap*ic_cap+-1.27500e-06*ic_cap+1.17000e-04'
+ mcrdlm1l1_ca_w_0_140_s_0_420 = '-2.01250e-06*ic_cap*ic_cap+-1.27500e-06*ic_cap+1.17000e-04'
+ mcrdlm1l1_ca_w_0_140_s_0_560 = '-2.01250e-06*ic_cap*ic_cap+-1.27500e-06*ic_cap+1.17000e-04'
+ mcrdlm1l1_ca_w_0_140_s_0_840 = '-2.01250e-06*ic_cap*ic_cap+-1.27500e-06*ic_cap+1.17000e-04'
+ mcrdlm1l1_ca_w_0_140_s_1_540 = '-2.01250e-06*ic_cap*ic_cap+-1.27500e-06*ic_cap+1.17000e-04'
+ mcrdlm1l1_ca_w_0_140_s_3_500 = '-2.01250e-06*ic_cap*ic_cap+-1.27500e-06*ic_cap+1.17000e-04'
+ mcrdlm1l1_ca_w_1_120_s_0_140 = '-2.01250e-06*ic_cap*ic_cap+-1.27500e-06*ic_cap+1.17000e-04'
+ mcrdlm1l1_ca_w_1_120_s_0_175 = '-2.01250e-06*ic_cap*ic_cap+-1.27500e-06*ic_cap+1.17000e-04'
+ mcrdlm1l1_ca_w_1_120_s_0_210 = '-2.01250e-06*ic_cap*ic_cap+-1.27500e-06*ic_cap+1.17000e-04'
+ mcrdlm1l1_ca_w_1_120_s_0_280 = '-2.01250e-06*ic_cap*ic_cap+-1.27500e-06*ic_cap+1.17000e-04'
+ mcrdlm1l1_ca_w_1_120_s_0_350 = '-2.01250e-06*ic_cap*ic_cap+-1.27500e-06*ic_cap+1.17000e-04'
+ mcrdlm1l1_ca_w_1_120_s_0_420 = '-2.01250e-06*ic_cap*ic_cap+-1.27500e-06*ic_cap+1.17000e-04'
+ mcrdlm1l1_ca_w_1_120_s_0_560 = '-2.01250e-06*ic_cap*ic_cap+-1.27500e-06*ic_cap+1.17000e-04'
+ mcrdlm1l1_ca_w_1_120_s_0_840 = '-2.01250e-06*ic_cap*ic_cap+-1.27500e-06*ic_cap+1.17000e-04'
+ mcrdlm1l1_ca_w_1_120_s_1_540 = '-2.01250e-06*ic_cap*ic_cap+-1.27500e-06*ic_cap+1.17000e-04'
+ mcrdlm1l1_ca_w_1_120_s_3_500 = '-2.01250e-06*ic_cap*ic_cap+-1.27500e-06*ic_cap+1.17000e-04'
+ mcrdlm1l1_cc_w_0_140_s_0_140 = '-7.75000e-13*ic_cap*ic_cap+-4.00000e-13*ic_cap+9.58000e-11'
+ mcrdlm1l1_cc_w_0_140_s_0_175 = '-7.00000e-13*ic_cap*ic_cap+-4.50000e-13*ic_cap+9.30000e-11'
+ mcrdlm1l1_cc_w_0_140_s_0_210 = '-5.96875e-13*ic_cap*ic_cap+-3.37500e-13*ic_cap+8.74000e-11'
+ mcrdlm1l1_cc_w_0_140_s_0_280 = '-4.06250e-13*ic_cap*ic_cap+-3.00000e-13*ic_cap+7.52000e-11'
+ mcrdlm1l1_cc_w_0_140_s_0_350 = '-3.25000e-13*ic_cap*ic_cap+-1.75000e-13*ic_cap+6.40000e-11'
+ mcrdlm1l1_cc_w_0_140_s_0_420 = '-1.90625e-13*ic_cap*ic_cap+-8.75000e-14*ic_cap+5.38000e-11'
+ mcrdlm1l1_cc_w_0_140_s_0_560 = '-6.87500e-14*ic_cap*ic_cap+-5.00000e-14*ic_cap+4.04000e-11'
+ mcrdlm1l1_cc_w_0_140_s_0_840 = '1.87500e-14*ic_cap*ic_cap+2.50000e-14*ic_cap+2.60000e-11'
+ mcrdlm1l1_cc_w_0_140_s_1_540 = '5.31250e-14*ic_cap*ic_cap+3.75000e-14*ic_cap+1.14000e-11'
+ mcrdlm1l1_cc_w_0_140_s_3_500 = '2.96875e-14*ic_cap*ic_cap+2.37500e-14*ic_cap+2.65000e-12'
+ mcrdlm1l1_cc_w_1_120_s_0_140 = '-6.56250e-13*ic_cap*ic_cap+-1.25000e-13*ic_cap+1.12000e-10'
+ mcrdlm1l1_cc_w_1_120_s_0_175 = '-6.40625e-13*ic_cap*ic_cap+-3.12500e-13*ic_cap+1.09000e-10'
+ mcrdlm1l1_cc_w_1_120_s_0_210 = '-5.71875e-13*ic_cap*ic_cap+-3.12500e-13*ic_cap+1.03000e-10'
+ mcrdlm1l1_cc_w_1_120_s_0_280 = '-3.87500e-13*ic_cap*ic_cap+-2.25000e-13*ic_cap+8.88000e-11'
+ mcrdlm1l1_cc_w_1_120_s_0_350 = '-2.31250e-13*ic_cap*ic_cap+-1.50000e-13*ic_cap+7.58000e-11'
+ mcrdlm1l1_cc_w_1_120_s_0_420 = '-1.59375e-13*ic_cap*ic_cap+-6.25000e-14*ic_cap+6.55000e-11'
+ mcrdlm1l1_cc_w_1_120_s_0_560 = '-4.06250e-14*ic_cap*ic_cap+1.25000e-14*ic_cap+5.06000e-11'
+ mcrdlm1l1_cc_w_1_120_s_0_840 = '5.62500e-14*ic_cap*ic_cap+5.00000e-14*ic_cap+3.41000e-11'
+ mcrdlm1l1_cc_w_1_120_s_1_540 = '8.12500e-14*ic_cap*ic_cap+5.00000e-14*ic_cap+1.72000e-11'
+ mcrdlm1l1_cc_w_1_120_s_3_500 = '4.18750e-14*ic_cap*ic_cap+4.00000e-14*ic_cap+5.02000e-12'
+ mcrdlm1l1_cf_w_0_140_s_0_140 = '-6.28125e-14*ic_cap*ic_cap+-5.12500e-14*ic_cap+7.64000e-12'
+ mcrdlm1l1_cf_w_0_140_s_0_175 = '-9.65625e-14*ic_cap*ic_cap+-7.12500e-14*ic_cap+9.66000e-12'
+ mcrdlm1l1_cf_w_0_140_s_0_210 = '-1.27813e-13*ic_cap*ic_cap+-9.62500e-14*ic_cap+1.16000e-11'
+ mcrdlm1l1_cf_w_0_140_s_0_280 = '-1.90625e-13*ic_cap*ic_cap+-1.37500e-13*ic_cap+1.53000e-11'
+ mcrdlm1l1_cf_w_0_140_s_0_350 = '-2.40625e-13*ic_cap*ic_cap+-1.62500e-13*ic_cap+1.86000e-11'
+ mcrdlm1l1_cf_w_0_140_s_0_420 = '-2.87500e-13*ic_cap*ic_cap+-2.00000e-13*ic_cap+2.18000e-11'
+ mcrdlm1l1_cf_w_0_140_s_0_560 = '-3.56250e-13*ic_cap*ic_cap+-2.50000e-13*ic_cap+2.73000e-11'
+ mcrdlm1l1_cf_w_0_140_s_0_840 = '-4.50000e-13*ic_cap*ic_cap+-3.00000e-13*ic_cap+3.58000e-11'
+ mcrdlm1l1_cf_w_0_140_s_1_540 = '-5.09375e-13*ic_cap*ic_cap+-3.62500e-13*ic_cap+4.74000e-11'
+ mcrdlm1l1_cf_w_0_140_s_3_500 = '-5.00000e-13*ic_cap*ic_cap+-3.50000e-13*ic_cap+5.60000e-11'
+ mcrdlm1l1_cf_w_1_120_s_0_140 = '-6.53125e-14*ic_cap*ic_cap+-5.37500e-14*ic_cap+7.79000e-12'
+ mcrdlm1l1_cf_w_1_120_s_0_175 = '-9.96875e-14*ic_cap*ic_cap+-7.62500e-14*ic_cap+9.81000e-12'
+ mcrdlm1l1_cf_w_1_120_s_0_210 = '-1.30000e-13*ic_cap*ic_cap+-9.50000e-14*ic_cap+1.17000e-11'
+ mcrdlm1l1_cf_w_1_120_s_0_280 = '-1.90625e-13*ic_cap*ic_cap+-1.37500e-13*ic_cap+1.54000e-11'
+ mcrdlm1l1_cf_w_1_120_s_0_350 = '-2.43750e-13*ic_cap*ic_cap+-1.75000e-13*ic_cap+1.88000e-11'
+ mcrdlm1l1_cf_w_1_120_s_0_420 = '-2.87500e-13*ic_cap*ic_cap+-2.00000e-13*ic_cap+2.19000e-11'
+ mcrdlm1l1_cf_w_1_120_s_0_560 = '-3.59375e-13*ic_cap*ic_cap+-2.37500e-13*ic_cap+2.74000e-11'
+ mcrdlm1l1_cf_w_1_120_s_0_840 = '-4.50000e-13*ic_cap*ic_cap+-3.25000e-13*ic_cap+3.61000e-11'
+ mcrdlm1l1_cf_w_1_120_s_1_540 = '-5.15625e-13*ic_cap*ic_cap+-3.62500e-13*ic_cap+4.86000e-11'
+ mcrdlm1l1_cf_w_1_120_s_3_500 = '-5.06250e-13*ic_cap*ic_cap+-3.50000e-13*ic_cap+6.00000e-11'
+ mcrdlm1p1_ca_w_0_140_s_0_140 = '-7.09375e-07*ic_cap*ic_cap+-4.12500e-07*ic_cap+4.78000e-05'
+ mcrdlm1p1_ca_w_0_140_s_0_175 = '-7.09375e-07*ic_cap*ic_cap+-4.12500e-07*ic_cap+4.78000e-05'
+ mcrdlm1p1_ca_w_0_140_s_0_210 = '-7.09375e-07*ic_cap*ic_cap+-4.12500e-07*ic_cap+4.78000e-05'
+ mcrdlm1p1_ca_w_0_140_s_0_280 = '-7.09375e-07*ic_cap*ic_cap+-4.12500e-07*ic_cap+4.78000e-05'
+ mcrdlm1p1_ca_w_0_140_s_0_350 = '-7.09375e-07*ic_cap*ic_cap+-4.12500e-07*ic_cap+4.78000e-05'
+ mcrdlm1p1_ca_w_0_140_s_0_420 = '-7.09375e-07*ic_cap*ic_cap+-4.12500e-07*ic_cap+4.78000e-05'
+ mcrdlm1p1_ca_w_0_140_s_0_560 = '-7.09375e-07*ic_cap*ic_cap+-4.12500e-07*ic_cap+4.78000e-05'
+ mcrdlm1p1_ca_w_0_140_s_0_840 = '-7.09375e-07*ic_cap*ic_cap+-4.12500e-07*ic_cap+4.78000e-05'
+ mcrdlm1p1_ca_w_0_140_s_1_540 = '-7.09375e-07*ic_cap*ic_cap+-4.12500e-07*ic_cap+4.78000e-05'
+ mcrdlm1p1_ca_w_0_140_s_3_500 = '-7.09375e-07*ic_cap*ic_cap+-4.12500e-07*ic_cap+4.78000e-05'
+ mcrdlm1p1_ca_w_1_120_s_0_140 = '-7.09375e-07*ic_cap*ic_cap+-4.12500e-07*ic_cap+4.78000e-05'
+ mcrdlm1p1_ca_w_1_120_s_0_175 = '-7.09375e-07*ic_cap*ic_cap+-4.12500e-07*ic_cap+4.78000e-05'
+ mcrdlm1p1_ca_w_1_120_s_0_210 = '-7.09375e-07*ic_cap*ic_cap+-4.12500e-07*ic_cap+4.78000e-05'
+ mcrdlm1p1_ca_w_1_120_s_0_280 = '-7.09375e-07*ic_cap*ic_cap+-4.12500e-07*ic_cap+4.78000e-05'
+ mcrdlm1p1_ca_w_1_120_s_0_350 = '-7.09375e-07*ic_cap*ic_cap+-4.12500e-07*ic_cap+4.78000e-05'
+ mcrdlm1p1_ca_w_1_120_s_0_420 = '-7.09375e-07*ic_cap*ic_cap+-4.12500e-07*ic_cap+4.78000e-05'
+ mcrdlm1p1_ca_w_1_120_s_0_560 = '-7.09375e-07*ic_cap*ic_cap+-4.12500e-07*ic_cap+4.78000e-05'
+ mcrdlm1p1_ca_w_1_120_s_0_840 = '-7.09375e-07*ic_cap*ic_cap+-4.12500e-07*ic_cap+4.78000e-05'
+ mcrdlm1p1_ca_w_1_120_s_1_540 = '-7.09375e-07*ic_cap*ic_cap+-4.12500e-07*ic_cap+4.78000e-05'
+ mcrdlm1p1_ca_w_1_120_s_3_500 = '-7.09375e-07*ic_cap*ic_cap+-4.12500e-07*ic_cap+4.78000e-05'
+ mcrdlm1p1_cc_w_0_140_s_0_140 = '-9.15625e-13*ic_cap*ic_cap+-5.12500e-13*ic_cap+1.03000e-10'
+ mcrdlm1p1_cc_w_0_140_s_0_175 = '-8.84375e-13*ic_cap*ic_cap+-5.37500e-13*ic_cap+1.01000e-10'
+ mcrdlm1p1_cc_w_0_140_s_0_210 = '-7.37500e-13*ic_cap*ic_cap+-3.75000e-13*ic_cap+9.50000e-11'
+ mcrdlm1p1_cc_w_0_140_s_0_280 = '-5.31250e-13*ic_cap*ic_cap+-3.50000e-13*ic_cap+8.37000e-11'
+ mcrdlm1p1_cc_w_0_140_s_0_350 = '-3.96875e-13*ic_cap*ic_cap+-2.37500e-13*ic_cap+7.21000e-11'
+ mcrdlm1p1_cc_w_0_140_s_0_420 = '-2.87500e-13*ic_cap*ic_cap+-1.75000e-13*ic_cap+6.25000e-11'
+ mcrdlm1p1_cc_w_0_140_s_0_560 = '-1.37500e-13*ic_cap*ic_cap+-1.00000e-13*ic_cap+4.94000e-11'
+ mcrdlm1p1_cc_w_0_140_s_0_840 = '-2.18750e-14*ic_cap*ic_cap+-1.25000e-14*ic_cap+3.47000e-11'
+ mcrdlm1p1_cc_w_0_140_s_1_540 = '7.50000e-14*ic_cap*ic_cap+5.00000e-14*ic_cap+1.81000e-11'
+ mcrdlm1p1_cc_w_0_140_s_3_500 = '6.09375e-14*ic_cap*ic_cap+4.62500e-14*ic_cap+5.22000e-12'
+ mcrdlm1p1_cc_w_1_120_s_0_140 = '-7.18750e-13*ic_cap*ic_cap+-3.75000e-13*ic_cap+1.23000e-10'
+ mcrdlm1p1_cc_w_1_120_s_0_175 = '-7.18750e-13*ic_cap*ic_cap+-3.75000e-13*ic_cap+1.20000e-10'
+ mcrdlm1p1_cc_w_1_120_s_0_210 = '-5.62500e-13*ic_cap*ic_cap+-2.50000e-13*ic_cap+1.13000e-10'
+ mcrdlm1p1_cc_w_1_120_s_0_280 = '-4.28125e-13*ic_cap*ic_cap+-3.37500e-13*ic_cap+9.92000e-11'
+ mcrdlm1p1_cc_w_1_120_s_0_350 = '-2.75000e-13*ic_cap*ic_cap+-1.75000e-13*ic_cap+8.63000e-11'
+ mcrdlm1p1_cc_w_1_120_s_0_420 = '-1.90625e-13*ic_cap*ic_cap+-1.12500e-13*ic_cap+7.59000e-11'
+ mcrdlm1p1_cc_w_1_120_s_0_560 = '-7.18750e-14*ic_cap*ic_cap+-3.75000e-14*ic_cap+6.08000e-11'
+ mcrdlm1p1_cc_w_1_120_s_0_840 = '5.00000e-14*ic_cap*ic_cap+2.50000e-14*ic_cap+4.35000e-11'
+ mcrdlm1p1_cc_w_1_120_s_1_540 = '1.06250e-13*ic_cap*ic_cap+7.50000e-14*ic_cap+2.44000e-11'
+ mcrdlm1p1_cc_w_1_120_s_3_500 = '9.09375e-14*ic_cap*ic_cap+6.62500e-14*ic_cap+8.04000e-12'
+ mcrdlm1p1_cf_w_0_140_s_0_140 = '-2.03125e-14*ic_cap*ic_cap+-1.37500e-14*ic_cap+3.31000e-12'
+ mcrdlm1p1_cf_w_0_140_s_0_175 = '-3.21875e-14*ic_cap*ic_cap+-2.12500e-14*ic_cap+4.13000e-12'
+ mcrdlm1p1_cf_w_0_140_s_0_210 = '-4.43750e-14*ic_cap*ic_cap+-2.75000e-14*ic_cap+4.96000e-12'
+ mcrdlm1p1_cf_w_0_140_s_0_280 = '-6.78125e-14*ic_cap*ic_cap+-4.12500e-14*ic_cap+6.57000e-12'
+ mcrdlm1p1_cf_w_0_140_s_0_350 = '-9.09375e-14*ic_cap*ic_cap+-5.62500e-14*ic_cap+8.13000e-12'
+ mcrdlm1p1_cf_w_0_140_s_0_420 = '-1.12812e-13*ic_cap*ic_cap+-6.62500e-14*ic_cap+9.69000e-12'
+ mcrdlm1p1_cf_w_0_140_s_0_560 = '-1.48437e-13*ic_cap*ic_cap+-9.37500e-14*ic_cap+1.25000e-11'
+ mcrdlm1p1_cf_w_0_140_s_0_840 = '-2.18750e-13*ic_cap*ic_cap+-1.25000e-13*ic_cap+1.77000e-11'
+ mcrdlm1p1_cf_w_0_140_s_1_540 = '-3.06250e-13*ic_cap*ic_cap+-2.00000e-13*ic_cap+2.71000e-11'
+ mcrdlm1p1_cf_w_0_140_s_3_500 = '-3.28125e-13*ic_cap*ic_cap+-2.12500e-13*ic_cap+3.80000e-11'
+ mcrdlm1p1_cf_w_1_120_s_0_140 = '-2.31250e-14*ic_cap*ic_cap+-1.50000e-14*ic_cap+3.46000e-12'
+ mcrdlm1p1_cf_w_1_120_s_0_175 = '-3.50000e-14*ic_cap*ic_cap+-2.25000e-14*ic_cap+4.29000e-12'
+ mcrdlm1p1_cf_w_1_120_s_0_210 = '-4.81250e-14*ic_cap*ic_cap+-2.75000e-14*ic_cap+5.11000e-12'
+ mcrdlm1p1_cf_w_1_120_s_0_280 = '-7.09375e-14*ic_cap*ic_cap+-4.37500e-14*ic_cap+6.72000e-12'
+ mcrdlm1p1_cf_w_1_120_s_0_350 = '-9.28125e-14*ic_cap*ic_cap+-5.62500e-14*ic_cap+8.28000e-12'
+ mcrdlm1p1_cf_w_1_120_s_0_420 = '-1.14375e-13*ic_cap*ic_cap+-7.00000e-14*ic_cap+9.81000e-12'
+ mcrdlm1p1_cf_w_1_120_s_0_560 = '-1.54688e-13*ic_cap*ic_cap+-9.37500e-14*ic_cap+1.27000e-11'
+ mcrdlm1p1_cf_w_1_120_s_0_840 = '-2.18750e-13*ic_cap*ic_cap+-1.25000e-13*ic_cap+1.79000e-11'
+ mcrdlm1p1_cf_w_1_120_s_1_540 = '-3.15625e-13*ic_cap*ic_cap+-1.87500e-13*ic_cap+2.79000e-11'
+ mcrdlm1p1_cf_w_1_120_s_3_500 = '-3.37500e-13*ic_cap*ic_cap+-2.25000e-13*ic_cap+4.07000e-11'
+ mcrdlm2_ca_w_10_000_s_10_000 = '-2.71875e-08*ic_cap*ic_cap+-1.62500e-08*ic_cap+3.10000e-06'
+ mcrdlm2_ca_w_10_000_s_12_000 = '-2.71875e-08*ic_cap*ic_cap+-1.62500e-08*ic_cap+3.10000e-06'
+ mcrdlm2_ca_w_10_000_s_30_000 = '-2.71875e-08*ic_cap*ic_cap+-1.62500e-08*ic_cap+3.10000e-06'
+ mcrdlm2_ca_w_10_000_s_5_000 = '-2.71875e-08*ic_cap*ic_cap+-1.62500e-08*ic_cap+3.10000e-06'
+ mcrdlm2_ca_w_10_000_s_8_000 = '-2.71875e-08*ic_cap*ic_cap+-1.62500e-08*ic_cap+3.10000e-06'
+ mcrdlm2_ca_w_40_000_s_10_000 = '-2.71875e-08*ic_cap*ic_cap+-1.62500e-08*ic_cap+3.10000e-06'
+ mcrdlm2_ca_w_40_000_s_12_000 = '-2.71875e-08*ic_cap*ic_cap+-1.62500e-08*ic_cap+3.10000e-06'
+ mcrdlm2_ca_w_40_000_s_30_000 = '-2.71875e-08*ic_cap*ic_cap+-1.62500e-08*ic_cap+3.10000e-06'
+ mcrdlm2_ca_w_40_000_s_5_000 = '-2.71875e-08*ic_cap*ic_cap+-1.62500e-08*ic_cap+3.10000e-06'
+ mcrdlm2_ca_w_40_000_s_8_000 = '-2.71875e-08*ic_cap*ic_cap+-1.62500e-08*ic_cap+3.10000e-06'
+ mcrdlm2_cc_w_10_000_s_10_000 = '-2.40625e-13*ic_cap*ic_cap+-1.62500e-13*ic_cap+3.04000e-11'
+ mcrdlm2_cc_w_10_000_s_12_000 = '-2.00000e-13*ic_cap*ic_cap+-1.25000e-13*ic_cap+2.65000e-11'
+ mcrdlm2_cc_w_10_000_s_30_000 = '-6.25000e-14*ic_cap*ic_cap+-5.00000e-14*ic_cap+1.12000e-11'
+ mcrdlm2_cc_w_10_000_s_5_000 = '-5.56250e-13*ic_cap*ic_cap+-3.50000e-13*ic_cap+4.99000e-11'
+ mcrdlm2_cc_w_10_000_s_8_000 = '-3.18750e-13*ic_cap*ic_cap+-2.00000e-13*ic_cap+3.59000e-11'
+ mcrdlm2_cc_w_40_000_s_10_000 = '-2.43750e-13*ic_cap*ic_cap+-1.50000e-13*ic_cap+4.03000e-11'
+ mcrdlm2_cc_w_40_000_s_12_000 = '-1.87500e-13*ic_cap*ic_cap+-1.25000e-13*ic_cap+3.58000e-11'
+ mcrdlm2_cc_w_40_000_s_30_000 = '-5.93750e-14*ic_cap*ic_cap+-3.75000e-14*ic_cap+1.83000e-11'
+ mcrdlm2_cc_w_40_000_s_5_000 = '-5.65625e-13*ic_cap*ic_cap+-3.37500e-13*ic_cap+6.12000e-11'
+ mcrdlm2_cc_w_40_000_s_8_000 = '-3.21875e-13*ic_cap*ic_cap+-2.12500e-13*ic_cap+4.62000e-11'
+ mcrdlm2_cf_w_10_000_s_10_000 = '-4.68750e-14*ic_cap*ic_cap+-3.75000e-14*ic_cap+1.27000e-11'
+ mcrdlm2_cf_w_10_000_s_12_000 = '-6.56250e-14*ic_cap*ic_cap+-3.75000e-14*ic_cap+1.46000e-11'
+ mcrdlm2_cf_w_10_000_s_30_000 = '-1.37500e-13*ic_cap*ic_cap+-1.00000e-13*ic_cap+2.52000e-11'
+ mcrdlm2_cf_w_10_000_s_5_000 = '1.25000e-15*ic_cap*ic_cap+7.07000e-12'
+ mcrdlm2_cf_w_10_000_s_8_000 = '-2.81250e-14*ic_cap*ic_cap+-1.25000e-14*ic_cap+1.06000e-11'
+ mcrdlm2_cf_w_40_000_s_10_000 = '-4.68750e-14*ic_cap*ic_cap+-3.75000e-14*ic_cap+1.28000e-11'
+ mcrdlm2_cf_w_40_000_s_12_000 = '-5.93750e-14*ic_cap*ic_cap+-3.75000e-14*ic_cap+1.47000e-11'
+ mcrdlm2_cf_w_40_000_s_30_000 = '-1.25000e-13*ic_cap*ic_cap+-7.50000e-14*ic_cap+2.60000e-11'
+ mcrdlm2_cf_w_40_000_s_5_000 = '1.87500e-15*ic_cap*ic_cap+-2.50000e-15*ic_cap+7.14000e-12'
+ mcrdlm2_cf_w_40_000_s_8_000 = '-3.12500e-14*ic_cap*ic_cap+-2.50000e-14*ic_cap+1.07000e-11'
+ mcrdlm2d_ca_w_0_140_s_0_140 = '-2.40625e-07*ic_cap*ic_cap+-1.62500e-07*ic_cap+2.39000e-05'
+ mcrdlm2d_ca_w_0_140_s_0_175 = '-2.40625e-07*ic_cap*ic_cap+-1.62500e-07*ic_cap+2.39000e-05'
+ mcrdlm2d_ca_w_0_140_s_0_210 = '-2.40625e-07*ic_cap*ic_cap+-1.62500e-07*ic_cap+2.39000e-05'
+ mcrdlm2d_ca_w_0_140_s_0_280 = '-2.40625e-07*ic_cap*ic_cap+-1.62500e-07*ic_cap+2.39000e-05'
+ mcrdlm2d_ca_w_0_140_s_0_350 = '-2.40625e-07*ic_cap*ic_cap+-1.62500e-07*ic_cap+2.39000e-05'
+ mcrdlm2d_ca_w_0_140_s_0_420 = '-2.40625e-07*ic_cap*ic_cap+-1.62500e-07*ic_cap+2.39000e-05'
+ mcrdlm2d_ca_w_0_140_s_0_560 = '-2.40625e-07*ic_cap*ic_cap+-1.62500e-07*ic_cap+2.39000e-05'
+ mcrdlm2d_ca_w_0_140_s_0_840 = '-2.40625e-07*ic_cap*ic_cap+-1.62500e-07*ic_cap+2.39000e-05'
+ mcrdlm2d_ca_w_0_140_s_1_540 = '-2.40625e-07*ic_cap*ic_cap+-1.62500e-07*ic_cap+2.39000e-05'
+ mcrdlm2d_ca_w_0_140_s_3_500 = '-2.40625e-07*ic_cap*ic_cap+-1.62500e-07*ic_cap+2.39000e-05'
+ mcrdlm2d_ca_w_1_120_s_0_140 = '-2.40625e-07*ic_cap*ic_cap+-1.62500e-07*ic_cap+2.39000e-05'
+ mcrdlm2d_ca_w_1_120_s_0_175 = '-2.40625e-07*ic_cap*ic_cap+-1.62500e-07*ic_cap+2.39000e-05'
+ mcrdlm2d_ca_w_1_120_s_0_210 = '-2.40625e-07*ic_cap*ic_cap+-1.62500e-07*ic_cap+2.39000e-05'
+ mcrdlm2d_ca_w_1_120_s_0_280 = '-2.40625e-07*ic_cap*ic_cap+-1.62500e-07*ic_cap+2.39000e-05'
+ mcrdlm2d_ca_w_1_120_s_0_350 = '-2.40625e-07*ic_cap*ic_cap+-1.62500e-07*ic_cap+2.39000e-05'
+ mcrdlm2d_ca_w_1_120_s_0_420 = '-2.40625e-07*ic_cap*ic_cap+-1.62500e-07*ic_cap+2.39000e-05'
+ mcrdlm2d_ca_w_1_120_s_0_560 = '-2.40625e-07*ic_cap*ic_cap+-1.62500e-07*ic_cap+2.39000e-05'
+ mcrdlm2d_ca_w_1_120_s_0_840 = '-2.40625e-07*ic_cap*ic_cap+-1.62500e-07*ic_cap+2.39000e-05'
+ mcrdlm2d_ca_w_1_120_s_1_540 = '-2.40625e-07*ic_cap*ic_cap+-1.62500e-07*ic_cap+2.39000e-05'
+ mcrdlm2d_ca_w_1_120_s_3_500 = '-2.40625e-07*ic_cap*ic_cap+-1.62500e-07*ic_cap+2.39000e-05'
+ mcrdlm2d_cc_w_0_140_s_0_140 = '-9.21875e-13*ic_cap*ic_cap+-5.37500e-13*ic_cap+1.05000e-10'
+ mcrdlm2d_cc_w_0_140_s_0_175 = '-9.43750e-13*ic_cap*ic_cap+-5.50000e-13*ic_cap+1.04000e-10'
+ mcrdlm2d_cc_w_0_140_s_0_210 = '-7.96875e-13*ic_cap*ic_cap+-4.12500e-13*ic_cap+9.82000e-11'
+ mcrdlm2d_cc_w_0_140_s_0_280 = '-6.09375e-13*ic_cap*ic_cap+-2.62500e-13*ic_cap+8.74000e-11'
+ mcrdlm2d_cc_w_0_140_s_0_350 = '-4.59375e-13*ic_cap*ic_cap+-2.87500e-13*ic_cap+7.60000e-11'
+ mcrdlm2d_cc_w_0_140_s_0_420 = '-3.71875e-13*ic_cap*ic_cap+-2.37500e-13*ic_cap+6.72000e-11'
+ mcrdlm2d_cc_w_0_140_s_0_560 = '-2.03125e-13*ic_cap*ic_cap+-1.37500e-13*ic_cap+5.42000e-11'
+ mcrdlm2d_cc_w_0_140_s_0_840 = '-8.43750e-14*ic_cap*ic_cap+-6.25000e-14*ic_cap+4.02000e-11'
+ mcrdlm2d_cc_w_0_140_s_1_540 = '1.25000e-14*ic_cap*ic_cap+2.42000e-11'
+ mcrdlm2d_cc_w_0_140_s_3_500 = '5.65625e-14*ic_cap*ic_cap+3.37500e-14*ic_cap+9.06000e-12'
+ mcrdlm2d_cc_w_1_120_s_0_140 = '-7.81250e-13*ic_cap*ic_cap+-3.75000e-13*ic_cap+1.30000e-10'
+ mcrdlm2d_cc_w_1_120_s_0_175 = '-7.18750e-13*ic_cap*ic_cap+-3.75000e-13*ic_cap+1.26000e-10'
+ mcrdlm2d_cc_w_1_120_s_0_210 = '-6.25000e-13*ic_cap*ic_cap+-5.00000e-13*ic_cap+1.20000e-10'
+ mcrdlm2d_cc_w_1_120_s_0_280 = '-4.78125e-13*ic_cap*ic_cap+-3.87500e-13*ic_cap+1.06000e-10'
+ mcrdlm2d_cc_w_1_120_s_0_350 = '-3.90625e-13*ic_cap*ic_cap+-2.37500e-13*ic_cap+9.41000e-11'
+ mcrdlm2d_cc_w_1_120_s_0_420 = '-2.65625e-13*ic_cap*ic_cap+-2.12500e-13*ic_cap+8.30000e-11'
+ mcrdlm2d_cc_w_1_120_s_0_560 = '-1.46875e-13*ic_cap*ic_cap+-8.75000e-14*ic_cap+6.81000e-11'
+ mcrdlm2d_cc_w_1_120_s_0_840 = '-1.87500e-14*ic_cap*ic_cap+-2.50000e-14*ic_cap+5.07000e-11'
+ mcrdlm2d_cc_w_1_120_s_1_540 = '6.56250e-14*ic_cap*ic_cap+3.75000e-14*ic_cap+3.12000e-11'
+ mcrdlm2d_cc_w_1_120_s_3_500 = '8.43750e-14*ic_cap*ic_cap+6.25000e-14*ic_cap+1.26000e-11'
+ mcrdlm2d_cf_w_0_140_s_0_140 = '-9.37500e-16*ic_cap*ic_cap+-1.25000e-15*ic_cap+1.67000e-12'
+ mcrdlm2d_cf_w_0_140_s_0_175 = '-5.00000e-15*ic_cap*ic_cap+-5.00000e-15*ic_cap+2.08000e-12'
+ mcrdlm2d_cf_w_0_140_s_0_210 = '-9.37500e-15*ic_cap*ic_cap+-7.50000e-15*ic_cap+2.51000e-12'
+ mcrdlm2d_cf_w_0_140_s_0_280 = '-1.81250e-14*ic_cap*ic_cap+-1.25000e-14*ic_cap+3.33000e-12'
+ mcrdlm2d_cf_w_0_140_s_0_350 = '-2.65625e-14*ic_cap*ic_cap+-1.62500e-14*ic_cap+4.14000e-12'
+ mcrdlm2d_cf_w_0_140_s_0_420 = '-3.53125e-14*ic_cap*ic_cap+-2.12500e-14*ic_cap+4.98000e-12'
+ mcrdlm2d_cf_w_0_140_s_0_560 = '-4.87500e-14*ic_cap*ic_cap+-3.25000e-14*ic_cap+6.50000e-12'
+ mcrdlm2d_cf_w_0_140_s_0_840 = '-7.84375e-14*ic_cap*ic_cap+-4.87500e-14*ic_cap+9.43000e-12'
+ mcrdlm2d_cf_w_0_140_s_1_540 = '-1.31250e-13*ic_cap*ic_cap+-7.50000e-14*ic_cap+1.57000e-11'
+ mcrdlm2d_cf_w_0_140_s_3_500 = '-1.87500e-13*ic_cap*ic_cap+-1.25000e-13*ic_cap+2.61000e-11'
+ mcrdlm2d_cf_w_1_120_s_0_140 = '-1.87500e-15*ic_cap*ic_cap+-2.50000e-15*ic_cap+1.71000e-12'
+ mcrdlm2d_cf_w_1_120_s_0_175 = '-5.93750e-15*ic_cap*ic_cap+-3.75000e-15*ic_cap+2.13000e-12'
+ mcrdlm2d_cf_w_1_120_s_0_210 = '-1.06250e-14*ic_cap*ic_cap+-7.50000e-15*ic_cap+2.55000e-12'
+ mcrdlm2d_cf_w_1_120_s_0_280 = '-1.87500e-14*ic_cap*ic_cap+-1.25000e-14*ic_cap+3.37000e-12'
+ mcrdlm2d_cf_w_1_120_s_0_350 = '-2.71875e-14*ic_cap*ic_cap+-1.87500e-14*ic_cap+4.19000e-12'
+ mcrdlm2d_cf_w_1_120_s_0_420 = '-3.50000e-14*ic_cap*ic_cap+-2.25000e-14*ic_cap+4.99000e-12'
+ mcrdlm2d_cf_w_1_120_s_0_560 = '-5.06250e-14*ic_cap*ic_cap+-3.25000e-14*ic_cap+6.56000e-12'
+ mcrdlm2d_cf_w_1_120_s_0_840 = '-7.81250e-14*ic_cap*ic_cap+-5.00000e-14*ic_cap+9.53000e-12'
+ mcrdlm2d_cf_w_1_120_s_1_540 = '-1.34375e-13*ic_cap*ic_cap+-8.75000e-14*ic_cap+1.61000e-11'
+ mcrdlm2d_cf_w_1_120_s_3_500 = '-1.93750e-13*ic_cap*ic_cap+-1.25000e-13*ic_cap+2.78000e-11'
+ mcrdlm2f_ca_w_0_140_s_0_140 = '-2.15625e-07*ic_cap*ic_cap+-1.37500e-07*ic_cap+2.06000e-05'
+ mcrdlm2f_ca_w_0_140_s_0_175 = '-2.15625e-07*ic_cap*ic_cap+-1.37500e-07*ic_cap+2.06000e-05'
+ mcrdlm2f_ca_w_0_140_s_0_210 = '-2.15625e-07*ic_cap*ic_cap+-1.37500e-07*ic_cap+2.06000e-05'
+ mcrdlm2f_ca_w_0_140_s_0_280 = '-2.15625e-07*ic_cap*ic_cap+-1.37500e-07*ic_cap+2.06000e-05'
+ mcrdlm2f_ca_w_0_140_s_0_350 = '-2.15625e-07*ic_cap*ic_cap+-1.37500e-07*ic_cap+2.06000e-05'
+ mcrdlm2f_ca_w_0_140_s_0_420 = '-2.15625e-07*ic_cap*ic_cap+-1.37500e-07*ic_cap+2.06000e-05'
+ mcrdlm2f_ca_w_0_140_s_0_560 = '-2.15625e-07*ic_cap*ic_cap+-1.37500e-07*ic_cap+2.06000e-05'
+ mcrdlm2f_ca_w_0_140_s_0_840 = '-2.15625e-07*ic_cap*ic_cap+-1.37500e-07*ic_cap+2.06000e-05'
+ mcrdlm2f_ca_w_0_140_s_1_540 = '-2.15625e-07*ic_cap*ic_cap+-1.37500e-07*ic_cap+2.06000e-05'
+ mcrdlm2f_ca_w_0_140_s_3_500 = '-2.15625e-07*ic_cap*ic_cap+-1.37500e-07*ic_cap+2.06000e-05'
+ mcrdlm2f_ca_w_1_120_s_0_140 = '-2.15625e-07*ic_cap*ic_cap+-1.37500e-07*ic_cap+2.06000e-05'
+ mcrdlm2f_ca_w_1_120_s_0_175 = '-2.15625e-07*ic_cap*ic_cap+-1.37500e-07*ic_cap+2.06000e-05'
+ mcrdlm2f_ca_w_1_120_s_0_210 = '-2.15625e-07*ic_cap*ic_cap+-1.37500e-07*ic_cap+2.06000e-05'
+ mcrdlm2f_ca_w_1_120_s_0_280 = '-2.15625e-07*ic_cap*ic_cap+-1.37500e-07*ic_cap+2.06000e-05'
+ mcrdlm2f_ca_w_1_120_s_0_350 = '-2.15625e-07*ic_cap*ic_cap+-1.37500e-07*ic_cap+2.06000e-05'
+ mcrdlm2f_ca_w_1_120_s_0_420 = '-2.15625e-07*ic_cap*ic_cap+-1.37500e-07*ic_cap+2.06000e-05'
+ mcrdlm2f_ca_w_1_120_s_0_560 = '-2.15625e-07*ic_cap*ic_cap+-1.37500e-07*ic_cap+2.06000e-05'
+ mcrdlm2f_ca_w_1_120_s_0_840 = '-2.15625e-07*ic_cap*ic_cap+-1.37500e-07*ic_cap+2.06000e-05'
+ mcrdlm2f_ca_w_1_120_s_1_540 = '-2.15625e-07*ic_cap*ic_cap+-1.37500e-07*ic_cap+2.06000e-05'
+ mcrdlm2f_ca_w_1_120_s_3_500 = '-2.15625e-07*ic_cap*ic_cap+-1.37500e-07*ic_cap+2.06000e-05'
+ mcrdlm2f_cc_w_0_140_s_0_140 = '-9.62500e-13*ic_cap*ic_cap+-5.25000e-13*ic_cap+1.06000e-10'
+ mcrdlm2f_cc_w_0_140_s_0_175 = '-9.28125e-13*ic_cap*ic_cap+-5.37500e-13*ic_cap+1.04000e-10'
+ mcrdlm2f_cc_w_0_140_s_0_210 = '-8.00000e-13*ic_cap*ic_cap+-4.25000e-13*ic_cap+9.87000e-11'
+ mcrdlm2f_cc_w_0_140_s_0_280 = '-6.15625e-13*ic_cap*ic_cap+-3.12500e-13*ic_cap+8.79000e-11'
+ mcrdlm2f_cc_w_0_140_s_0_350 = '-4.43750e-13*ic_cap*ic_cap+-3.50000e-13*ic_cap+7.66000e-11'
+ mcrdlm2f_cc_w_0_140_s_0_420 = '-3.90625e-13*ic_cap*ic_cap+-1.87500e-13*ic_cap+6.79000e-11'
+ mcrdlm2f_cc_w_0_140_s_0_560 = '-2.12500e-13*ic_cap*ic_cap+-1.50000e-13*ic_cap+5.51000e-11'
+ mcrdlm2f_cc_w_0_140_s_0_840 = '-9.37500e-14*ic_cap*ic_cap+-7.50000e-14*ic_cap+4.14000e-11'
+ mcrdlm2f_cc_w_0_140_s_1_540 = '6.25000e-15*ic_cap*ic_cap+2.56000e-11'
+ mcrdlm2f_cc_w_0_140_s_3_500 = '6.56250e-14*ic_cap*ic_cap+3.75000e-14*ic_cap+1.02000e-11'
+ mcrdlm2f_cc_w_1_120_s_0_140 = '-8.43750e-13*ic_cap*ic_cap+-3.75000e-13*ic_cap+1.32000e-10'
+ mcrdlm2f_cc_w_1_120_s_0_175 = '-7.81250e-13*ic_cap*ic_cap+-3.75000e-13*ic_cap+1.28000e-10'
+ mcrdlm2f_cc_w_1_120_s_0_210 = '-6.87500e-13*ic_cap*ic_cap+-5.00000e-13*ic_cap+1.22000e-10'
+ mcrdlm2f_cc_w_1_120_s_0_280 = '-5.28125e-13*ic_cap*ic_cap+-3.62500e-13*ic_cap+1.08000e-10'
+ mcrdlm2f_cc_w_1_120_s_0_350 = '-3.65625e-13*ic_cap*ic_cap+-2.37500e-13*ic_cap+9.52000e-11'
+ mcrdlm2f_cc_w_1_120_s_0_420 = '-2.71875e-13*ic_cap*ic_cap+-2.37500e-13*ic_cap+8.46000e-11'
+ mcrdlm2f_cc_w_1_120_s_0_560 = '-1.53125e-13*ic_cap*ic_cap+-1.12500e-13*ic_cap+6.97000e-11'
+ mcrdlm2f_cc_w_1_120_s_0_840 = '-2.50000e-14*ic_cap*ic_cap+-2.50000e-14*ic_cap+5.25000e-11'
+ mcrdlm2f_cc_w_1_120_s_1_540 = '6.56250e-14*ic_cap*ic_cap+3.75000e-14*ic_cap+3.30000e-11'
+ mcrdlm2f_cc_w_1_120_s_3_500 = '1.00000e-13*ic_cap*ic_cap+7.50000e-14*ic_cap+1.39000e-11'
+ mcrdlm2f_cf_w_0_140_s_0_140 = '-1.56250e-15*ic_cap*ic_cap+-1.25000e-15*ic_cap+1.44000e-12'
+ mcrdlm2f_cf_w_0_140_s_0_175 = '-5.31250e-15*ic_cap*ic_cap+-3.75000e-15*ic_cap+1.80000e-12'
+ mcrdlm2f_cf_w_0_140_s_0_210 = '-8.43750e-15*ic_cap*ic_cap+-6.25000e-15*ic_cap+2.16000e-12'
+ mcrdlm2f_cf_w_0_140_s_0_280 = '-1.68750e-14*ic_cap*ic_cap+-1.00000e-14*ic_cap+2.88000e-12'
+ mcrdlm2f_cf_w_0_140_s_0_350 = '-2.46875e-14*ic_cap*ic_cap+-1.62500e-14*ic_cap+3.58000e-12'
+ mcrdlm2f_cf_w_0_140_s_0_420 = '-3.21875e-14*ic_cap*ic_cap+-2.12500e-14*ic_cap+4.31000e-12'
+ mcrdlm2f_cf_w_0_140_s_0_560 = '-4.50000e-14*ic_cap*ic_cap+-3.00000e-14*ic_cap+5.64000e-12'
+ mcrdlm2f_cf_w_0_140_s_0_840 = '-7.18750e-14*ic_cap*ic_cap+-4.50000e-14*ic_cap+8.21000e-12'
+ mcrdlm2f_cf_w_0_140_s_1_540 = '-1.25000e-13*ic_cap*ic_cap+-7.50000e-14*ic_cap+1.39000e-11'
+ mcrdlm2f_cf_w_0_140_s_3_500 = '-1.87500e-13*ic_cap*ic_cap+-1.25000e-13*ic_cap+2.38000e-11'
+ mcrdlm2f_cf_w_1_120_s_0_140 = '-2.50000e-15*ic_cap*ic_cap+-2.50000e-15*ic_cap+1.48000e-12'
+ mcrdlm2f_cf_w_1_120_s_0_175 = '-6.25000e-15*ic_cap*ic_cap+-5.00000e-15*ic_cap+1.84000e-12'
+ mcrdlm2f_cf_w_1_120_s_0_210 = '-1.03125e-14*ic_cap*ic_cap+-6.25000e-15*ic_cap+2.20000e-12'
+ mcrdlm2f_cf_w_1_120_s_0_280 = '-1.78125e-14*ic_cap*ic_cap+-1.12500e-14*ic_cap+2.91000e-12'
+ mcrdlm2f_cf_w_1_120_s_0_350 = '-2.53125e-14*ic_cap*ic_cap+-1.62500e-14*ic_cap+3.62000e-12'
+ mcrdlm2f_cf_w_1_120_s_0_420 = '-3.28125e-14*ic_cap*ic_cap+-2.12500e-14*ic_cap+4.32000e-12'
+ mcrdlm2f_cf_w_1_120_s_0_560 = '-4.68750e-14*ic_cap*ic_cap+-3.00000e-14*ic_cap+5.68000e-12'
+ mcrdlm2f_cf_w_1_120_s_0_840 = '-7.28125e-14*ic_cap*ic_cap+-4.62500e-14*ic_cap+8.31000e-12'
+ mcrdlm2f_cf_w_1_120_s_1_540 = '-1.31250e-13*ic_cap*ic_cap+-7.50000e-14*ic_cap+1.42000e-11'
+ mcrdlm2f_cf_w_1_120_s_3_500 = '-1.93750e-13*ic_cap*ic_cap+-1.25000e-13*ic_cap+2.53000e-11'
+ mcrdlm2l1_ca_w_0_140_s_0_140 = '-4.78125e-07*ic_cap*ic_cap+-3.12500e-07*ic_cap+4.01000e-05'
+ mcrdlm2l1_ca_w_0_140_s_0_175 = '-4.78125e-07*ic_cap*ic_cap+-3.12500e-07*ic_cap+4.01000e-05'
+ mcrdlm2l1_ca_w_0_140_s_0_210 = '-4.78125e-07*ic_cap*ic_cap+-3.12500e-07*ic_cap+4.01000e-05'
+ mcrdlm2l1_ca_w_0_140_s_0_280 = '-4.78125e-07*ic_cap*ic_cap+-3.12500e-07*ic_cap+4.01000e-05'
+ mcrdlm2l1_ca_w_0_140_s_0_350 = '-4.78125e-07*ic_cap*ic_cap+-3.12500e-07*ic_cap+4.01000e-05'
+ mcrdlm2l1_ca_w_0_140_s_0_420 = '-4.78125e-07*ic_cap*ic_cap+-3.12500e-07*ic_cap+4.01000e-05'
+ mcrdlm2l1_ca_w_0_140_s_0_560 = '-4.78125e-07*ic_cap*ic_cap+-3.12500e-07*ic_cap+4.01000e-05'
+ mcrdlm2l1_ca_w_0_140_s_0_840 = '-4.78125e-07*ic_cap*ic_cap+-3.12500e-07*ic_cap+4.01000e-05'
+ mcrdlm2l1_ca_w_0_140_s_1_540 = '-4.78125e-07*ic_cap*ic_cap+-3.12500e-07*ic_cap+4.01000e-05'
+ mcrdlm2l1_ca_w_0_140_s_3_500 = '-4.78125e-07*ic_cap*ic_cap+-3.12500e-07*ic_cap+4.01000e-05'
+ mcrdlm2l1_ca_w_1_120_s_0_140 = '-4.78125e-07*ic_cap*ic_cap+-3.12500e-07*ic_cap+4.01000e-05'
+ mcrdlm2l1_ca_w_1_120_s_0_175 = '-4.78125e-07*ic_cap*ic_cap+-3.12500e-07*ic_cap+4.01000e-05'
+ mcrdlm2l1_ca_w_1_120_s_0_210 = '-4.78125e-07*ic_cap*ic_cap+-3.12500e-07*ic_cap+4.01000e-05'
+ mcrdlm2l1_ca_w_1_120_s_0_280 = '-4.78125e-07*ic_cap*ic_cap+-3.12500e-07*ic_cap+4.01000e-05'
+ mcrdlm2l1_ca_w_1_120_s_0_350 = '-4.78125e-07*ic_cap*ic_cap+-3.12500e-07*ic_cap+4.01000e-05'
+ mcrdlm2l1_ca_w_1_120_s_0_420 = '-4.78125e-07*ic_cap*ic_cap+-3.12500e-07*ic_cap+4.01000e-05'
+ mcrdlm2l1_ca_w_1_120_s_0_560 = '-4.78125e-07*ic_cap*ic_cap+-3.12500e-07*ic_cap+4.01000e-05'
+ mcrdlm2l1_ca_w_1_120_s_0_840 = '-4.78125e-07*ic_cap*ic_cap+-3.12500e-07*ic_cap+4.01000e-05'
+ mcrdlm2l1_ca_w_1_120_s_1_540 = '-4.78125e-07*ic_cap*ic_cap+-3.12500e-07*ic_cap+4.01000e-05'
+ mcrdlm2l1_ca_w_1_120_s_3_500 = '-4.78125e-07*ic_cap*ic_cap+-3.12500e-07*ic_cap+4.01000e-05'
+ mcrdlm2l1_cc_w_0_140_s_0_140 = '-8.87500e-13*ic_cap*ic_cap+-5.25000e-13*ic_cap+1.03000e-10'
+ mcrdlm2l1_cc_w_0_140_s_0_175 = '-8.53125e-13*ic_cap*ic_cap+-5.37500e-13*ic_cap+1.01000e-10'
+ mcrdlm2l1_cc_w_0_140_s_0_210 = '-7.62500e-13*ic_cap*ic_cap+-4.00000e-13*ic_cap+9.59000e-11'
+ mcrdlm2l1_cc_w_0_140_s_0_280 = '-5.68750e-13*ic_cap*ic_cap+-3.25000e-13*ic_cap+8.47000e-11'
+ mcrdlm2l1_cc_w_0_140_s_0_350 = '-4.25000e-13*ic_cap*ic_cap+-2.50000e-13*ic_cap+7.32000e-11'
+ mcrdlm2l1_cc_w_0_140_s_0_420 = '-3.06250e-13*ic_cap*ic_cap+-1.75000e-13*ic_cap+6.35000e-11'
+ mcrdlm2l1_cc_w_0_140_s_0_560 = '-1.71875e-13*ic_cap*ic_cap+-1.37500e-13*ic_cap+5.06000e-11'
+ mcrdlm2l1_cc_w_0_140_s_0_840 = '-4.06250e-14*ic_cap*ic_cap+-3.75000e-14*ic_cap+3.58000e-11'
+ mcrdlm2l1_cc_w_0_140_s_1_540 = '4.06250e-14*ic_cap*ic_cap+3.75000e-14*ic_cap+1.95000e-11'
+ mcrdlm2l1_cc_w_0_140_s_3_500 = '5.03125e-14*ic_cap*ic_cap+3.87500e-14*ic_cap+5.89000e-12'
+ mcrdlm2l1_cc_w_1_120_s_0_140 = '-7.18750e-13*ic_cap*ic_cap+-3.75000e-13*ic_cap+1.24000e-10'
+ mcrdlm2l1_cc_w_1_120_s_0_175 = '-7.18750e-13*ic_cap*ic_cap+-3.75000e-13*ic_cap+1.21000e-10'
+ mcrdlm2l1_cc_w_1_120_s_0_210 = '-6.25000e-13*ic_cap*ic_cap+-2.50000e-13*ic_cap+1.15000e-10'
+ mcrdlm2l1_cc_w_1_120_s_0_280 = '-4.78125e-13*ic_cap*ic_cap+-3.37500e-13*ic_cap+1.01000e-10'
+ mcrdlm2l1_cc_w_1_120_s_0_350 = '-3.09375e-13*ic_cap*ic_cap+-1.87500e-13*ic_cap+8.78000e-11'
+ mcrdlm2l1_cc_w_1_120_s_0_420 = '-2.12500e-13*ic_cap*ic_cap+-1.50000e-13*ic_cap+7.71000e-11'
+ mcrdlm2l1_cc_w_1_120_s_0_560 = '-9.37500e-14*ic_cap*ic_cap+-7.50000e-14*ic_cap+6.20000e-11'
+ mcrdlm2l1_cc_w_1_120_s_0_840 = '9.37500e-15*ic_cap*ic_cap+1.25000e-14*ic_cap+4.49000e-11'
+ mcrdlm2l1_cc_w_1_120_s_1_540 = '7.81250e-14*ic_cap*ic_cap+6.25000e-14*ic_cap+2.57000e-11'
+ mcrdlm2l1_cc_w_1_120_s_3_500 = '7.75000e-14*ic_cap*ic_cap+5.00000e-14*ic_cap+8.76000e-12'
+ mcrdlm2l1_cf_w_0_140_s_0_140 = '-7.18750e-15*ic_cap*ic_cap+-6.25000e-15*ic_cap+2.76000e-12'
+ mcrdlm2l1_cf_w_0_140_s_0_175 = '-1.50000e-14*ic_cap*ic_cap+-1.25000e-14*ic_cap+3.45000e-12'
+ mcrdlm2l1_cf_w_0_140_s_0_210 = '-2.31250e-14*ic_cap*ic_cap+-1.75000e-14*ic_cap+4.15000e-12'
+ mcrdlm2l1_cf_w_0_140_s_0_280 = '-3.93750e-14*ic_cap*ic_cap+-3.00000e-14*ic_cap+5.51000e-12'
+ mcrdlm2l1_cf_w_0_140_s_0_350 = '-5.56250e-14*ic_cap*ic_cap+-3.75000e-14*ic_cap+6.83000e-12'
+ mcrdlm2l1_cf_w_0_140_s_0_420 = '-7.09375e-14*ic_cap*ic_cap+-4.62500e-14*ic_cap+8.16000e-12'
+ mcrdlm2l1_cf_w_0_140_s_0_560 = '-9.75000e-14*ic_cap*ic_cap+-6.50000e-14*ic_cap+1.06000e-11'
+ mcrdlm2l1_cf_w_0_140_s_0_840 = '-1.46875e-13*ic_cap*ic_cap+-8.75000e-14*ic_cap+1.51000e-11'
+ mcrdlm2l1_cf_w_0_140_s_1_540 = '-2.15625e-13*ic_cap*ic_cap+-1.37500e-13*ic_cap+2.37000e-11'
+ mcrdlm2l1_cf_w_0_140_s_3_500 = '-2.50000e-13*ic_cap*ic_cap+-1.75000e-13*ic_cap+3.47000e-11'
+ mcrdlm2l1_cf_w_1_120_s_0_140 = '-7.81250e-15*ic_cap*ic_cap+-6.25000e-15*ic_cap+2.80000e-12'
+ mcrdlm2l1_cf_w_1_120_s_0_175 = '-1.59375e-14*ic_cap*ic_cap+-1.12500e-14*ic_cap+3.50000e-12'
+ mcrdlm2l1_cf_w_1_120_s_0_210 = '-2.43750e-14*ic_cap*ic_cap+-1.75000e-14*ic_cap+4.19000e-12'
+ mcrdlm2l1_cf_w_1_120_s_0_280 = '-4.03125e-14*ic_cap*ic_cap+-2.87500e-14*ic_cap+5.55000e-12'
+ mcrdlm2l1_cf_w_1_120_s_0_350 = '-5.56250e-14*ic_cap*ic_cap+-3.75000e-14*ic_cap+6.88000e-12'
+ mcrdlm2l1_cf_w_1_120_s_0_420 = '-7.03125e-14*ic_cap*ic_cap+-4.87500e-14*ic_cap+8.17000e-12'
+ mcrdlm2l1_cf_w_1_120_s_0_560 = '-1.00312e-13*ic_cap*ic_cap+-6.62500e-14*ic_cap+1.07000e-11'
+ mcrdlm2l1_cf_w_1_120_s_0_840 = '-1.43750e-13*ic_cap*ic_cap+-1.00000e-13*ic_cap+1.52000e-11'
+ mcrdlm2l1_cf_w_1_120_s_1_540 = '-2.18750e-13*ic_cap*ic_cap+-1.50000e-13*ic_cap+2.43000e-11'
+ mcrdlm2l1_cf_w_1_120_s_3_500 = '-2.50000e-13*ic_cap*ic_cap+-1.75000e-13*ic_cap+3.70000e-11'
+ mcrdlm2m1_ca_w_0_140_s_0_140 = '-2.68125e-06*ic_cap*ic_cap+-1.27500e-06*ic_cap+1.31000e-04'
+ mcrdlm2m1_ca_w_0_140_s_0_175 = '-2.68125e-06*ic_cap*ic_cap+-1.27500e-06*ic_cap+1.31000e-04'
+ mcrdlm2m1_ca_w_0_140_s_0_210 = '-2.68125e-06*ic_cap*ic_cap+-1.27500e-06*ic_cap+1.31000e-04'
+ mcrdlm2m1_ca_w_0_140_s_0_280 = '-2.68125e-06*ic_cap*ic_cap+-1.27500e-06*ic_cap+1.31000e-04'
+ mcrdlm2m1_ca_w_0_140_s_0_350 = '-2.68125e-06*ic_cap*ic_cap+-1.27500e-06*ic_cap+1.31000e-04'
+ mcrdlm2m1_ca_w_0_140_s_0_420 = '-2.68125e-06*ic_cap*ic_cap+-1.27500e-06*ic_cap+1.31000e-04'
+ mcrdlm2m1_ca_w_0_140_s_0_560 = '-2.68125e-06*ic_cap*ic_cap+-1.27500e-06*ic_cap+1.31000e-04'
+ mcrdlm2m1_ca_w_0_140_s_0_840 = '-2.68125e-06*ic_cap*ic_cap+-1.27500e-06*ic_cap+1.31000e-04'
+ mcrdlm2m1_ca_w_0_140_s_1_540 = '-2.68125e-06*ic_cap*ic_cap+-1.27500e-06*ic_cap+1.31000e-04'
+ mcrdlm2m1_ca_w_0_140_s_3_500 = '-2.68125e-06*ic_cap*ic_cap+-1.27500e-06*ic_cap+1.31000e-04'
+ mcrdlm2m1_ca_w_1_120_s_0_140 = '-2.68125e-06*ic_cap*ic_cap+-1.27500e-06*ic_cap+1.31000e-04'
+ mcrdlm2m1_ca_w_1_120_s_0_175 = '-2.68125e-06*ic_cap*ic_cap+-1.27500e-06*ic_cap+1.31000e-04'
+ mcrdlm2m1_ca_w_1_120_s_0_210 = '-2.68125e-06*ic_cap*ic_cap+-1.27500e-06*ic_cap+1.31000e-04'
+ mcrdlm2m1_ca_w_1_120_s_0_280 = '-2.68125e-06*ic_cap*ic_cap+-1.27500e-06*ic_cap+1.31000e-04'
+ mcrdlm2m1_ca_w_1_120_s_0_350 = '-2.68125e-06*ic_cap*ic_cap+-1.27500e-06*ic_cap+1.31000e-04'
+ mcrdlm2m1_ca_w_1_120_s_0_420 = '-2.68125e-06*ic_cap*ic_cap+-1.27500e-06*ic_cap+1.31000e-04'
+ mcrdlm2m1_ca_w_1_120_s_0_560 = '-2.68125e-06*ic_cap*ic_cap+-1.27500e-06*ic_cap+1.31000e-04'
+ mcrdlm2m1_ca_w_1_120_s_0_840 = '-2.68125e-06*ic_cap*ic_cap+-1.27500e-06*ic_cap+1.31000e-04'
+ mcrdlm2m1_ca_w_1_120_s_1_540 = '-2.68125e-06*ic_cap*ic_cap+-1.27500e-06*ic_cap+1.31000e-04'
+ mcrdlm2m1_ca_w_1_120_s_3_500 = '-2.68125e-06*ic_cap*ic_cap+-1.27500e-06*ic_cap+1.31000e-04'
+ mcrdlm2m1_cc_w_0_140_s_0_140 = '-7.28125e-13*ic_cap*ic_cap+-3.87500e-13*ic_cap+9.48000e-11'
+ mcrdlm2m1_cc_w_0_140_s_0_175 = '-6.50000e-13*ic_cap*ic_cap+-4.50000e-13*ic_cap+9.20000e-11'
+ mcrdlm2m1_cc_w_0_140_s_0_210 = '-5.25000e-13*ic_cap*ic_cap+-3.25000e-13*ic_cap+8.60000e-11'
+ mcrdlm2m1_cc_w_0_140_s_0_280 = '-3.46875e-13*ic_cap*ic_cap+-2.62500e-13*ic_cap+7.41000e-11'
+ mcrdlm2m1_cc_w_0_140_s_0_350 = '-2.50000e-13*ic_cap*ic_cap+-2.00000e-13*ic_cap+6.26000e-11'
+ mcrdlm2m1_cc_w_0_140_s_0_420 = '-1.46875e-13*ic_cap*ic_cap+-1.37500e-13*ic_cap+5.25000e-11'
+ mcrdlm2m1_cc_w_0_140_s_0_560 = '-2.18750e-14*ic_cap*ic_cap+-3.75000e-14*ic_cap+3.93000e-11'
+ mcrdlm2m1_cc_w_0_140_s_0_840 = '6.25000e-14*ic_cap*ic_cap+2.50000e-14*ic_cap+2.49000e-11'
+ mcrdlm2m1_cc_w_0_140_s_1_540 = '7.50000e-14*ic_cap*ic_cap+5.00000e-14*ic_cap+1.08000e-11'
+ mcrdlm2m1_cc_w_0_140_s_3_500 = '3.09375e-14*ic_cap*ic_cap+2.62500e-14*ic_cap+2.50000e-12'
+ mcrdlm2m1_cc_w_1_120_s_0_140 = '-6.25000e-13*ic_cap*ic_cap+-2.50000e-13*ic_cap+1.11000e-10'
+ mcrdlm2m1_cc_w_1_120_s_0_175 = '-6.00000e-13*ic_cap*ic_cap+-2.75000e-13*ic_cap+1.08000e-10'
+ mcrdlm2m1_cc_w_1_120_s_0_210 = '-5.31250e-13*ic_cap*ic_cap+-3.25000e-13*ic_cap+1.02000e-10'
+ mcrdlm2m1_cc_w_1_120_s_0_280 = '-3.34375e-13*ic_cap*ic_cap+-2.12500e-13*ic_cap+8.75000e-11'
+ mcrdlm2m1_cc_w_1_120_s_0_350 = '-1.75000e-13*ic_cap*ic_cap+-1.50000e-13*ic_cap+7.44000e-11'
+ mcrdlm2m1_cc_w_1_120_s_0_420 = '-1.03125e-13*ic_cap*ic_cap+-6.25000e-14*ic_cap+6.42000e-11'
+ mcrdlm2m1_cc_w_1_120_s_0_560 = '9.37500e-15*ic_cap*ic_cap+-1.25000e-14*ic_cap+4.93000e-11'
+ mcrdlm2m1_cc_w_1_120_s_0_840 = '9.06250e-14*ic_cap*ic_cap+3.75000e-14*ic_cap+3.31000e-11'
+ mcrdlm2m1_cc_w_1_120_s_1_540 = '1.03125e-13*ic_cap*ic_cap+6.25000e-14*ic_cap+1.65000e-11'
+ mcrdlm2m1_cc_w_1_120_s_3_500 = '5.09375e-14*ic_cap*ic_cap+3.37500e-14*ic_cap+4.73000e-12'
+ mcrdlm2m1_cf_w_0_140_s_0_140 = '-9.96875e-14*ic_cap*ic_cap+-4.87500e-14*ic_cap+8.45000e-12'
+ mcrdlm2m1_cf_w_0_140_s_0_175 = '-1.44687e-13*ic_cap*ic_cap+-6.62500e-14*ic_cap+1.07000e-11'
+ mcrdlm2m1_cf_w_0_140_s_0_210 = '-1.90625e-13*ic_cap*ic_cap+-8.75000e-14*ic_cap+1.29000e-11'
+ mcrdlm2m1_cf_w_0_140_s_0_280 = '-2.65625e-13*ic_cap*ic_cap+-1.37500e-13*ic_cap+1.69000e-11'
+ mcrdlm2m1_cf_w_0_140_s_0_350 = '-3.34375e-13*ic_cap*ic_cap+-1.62500e-13*ic_cap+2.06000e-11'
+ mcrdlm2m1_cf_w_0_140_s_0_420 = '-3.90625e-13*ic_cap*ic_cap+-1.87500e-13*ic_cap+2.40000e-11'
+ mcrdlm2m1_cf_w_0_140_s_0_560 = '-4.87500e-13*ic_cap*ic_cap+-2.50000e-13*ic_cap+3.00000e-11'
+ mcrdlm2m1_cf_w_0_140_s_0_840 = '-5.81250e-13*ic_cap*ic_cap+-3.00000e-13*ic_cap+3.87000e-11'
+ mcrdlm2m1_cf_w_0_140_s_1_540 = '-6.46875e-13*ic_cap*ic_cap+-3.62500e-13*ic_cap+5.05000e-11'
+ mcrdlm2m1_cf_w_0_140_s_3_500 = '-6.21875e-13*ic_cap*ic_cap+-3.37500e-13*ic_cap+5.87000e-11'
+ mcrdlm2m1_cf_w_1_120_s_0_140 = '-9.84375e-14*ic_cap*ic_cap+-4.87500e-14*ic_cap+8.46000e-12'
+ mcrdlm2m1_cf_w_1_120_s_0_175 = '-1.43750e-13*ic_cap*ic_cap+-7.00000e-14*ic_cap+1.07000e-11'
+ mcrdlm2m1_cf_w_1_120_s_0_210 = '-1.90625e-13*ic_cap*ic_cap+-8.75000e-14*ic_cap+1.29000e-11'
+ mcrdlm2m1_cf_w_1_120_s_0_280 = '-2.65625e-13*ic_cap*ic_cap+-1.37500e-13*ic_cap+1.69000e-11'
+ mcrdlm2m1_cf_w_1_120_s_0_350 = '-3.40625e-13*ic_cap*ic_cap+-1.62500e-13*ic_cap+2.07000e-11'
+ mcrdlm2m1_cf_w_1_120_s_0_420 = '-3.87500e-13*ic_cap*ic_cap+-2.00000e-13*ic_cap+2.40000e-11'
+ mcrdlm2m1_cf_w_1_120_s_0_560 = '-4.78125e-13*ic_cap*ic_cap+-2.37500e-13*ic_cap+2.99000e-11'
+ mcrdlm2m1_cf_w_1_120_s_0_840 = '-5.84375e-13*ic_cap*ic_cap+-3.12500e-13*ic_cap+3.90000e-11'
+ mcrdlm2m1_cf_w_1_120_s_1_540 = '-6.50000e-13*ic_cap*ic_cap+-3.50000e-13*ic_cap+5.16000e-11'
+ mcrdlm2m1_cf_w_1_120_s_3_500 = '-6.43750e-13*ic_cap*ic_cap+-3.25000e-13*ic_cap+6.29000e-11'
+ mcrdlm2p1_ca_w_0_140_s_0_140 = '-3.40625e-07*ic_cap*ic_cap+-2.12500e-07*ic_cap+2.78000e-05'
+ mcrdlm2p1_ca_w_0_140_s_0_175 = '-3.40625e-07*ic_cap*ic_cap+-2.12500e-07*ic_cap+2.78000e-05'
+ mcrdlm2p1_ca_w_0_140_s_0_210 = '-3.40625e-07*ic_cap*ic_cap+-2.12500e-07*ic_cap+2.78000e-05'
+ mcrdlm2p1_ca_w_0_140_s_0_280 = '-3.40625e-07*ic_cap*ic_cap+-2.12500e-07*ic_cap+2.78000e-05'
+ mcrdlm2p1_ca_w_0_140_s_0_350 = '-3.40625e-07*ic_cap*ic_cap+-2.12500e-07*ic_cap+2.78000e-05'
+ mcrdlm2p1_ca_w_0_140_s_0_420 = '-3.40625e-07*ic_cap*ic_cap+-2.12500e-07*ic_cap+2.78000e-05'
+ mcrdlm2p1_ca_w_0_140_s_0_560 = '-3.40625e-07*ic_cap*ic_cap+-2.12500e-07*ic_cap+2.78000e-05'
+ mcrdlm2p1_ca_w_0_140_s_0_840 = '-3.40625e-07*ic_cap*ic_cap+-2.12500e-07*ic_cap+2.78000e-05'
+ mcrdlm2p1_ca_w_0_140_s_1_540 = '-3.40625e-07*ic_cap*ic_cap+-2.12500e-07*ic_cap+2.78000e-05'
+ mcrdlm2p1_ca_w_0_140_s_3_500 = '-3.40625e-07*ic_cap*ic_cap+-2.12500e-07*ic_cap+2.78000e-05'
+ mcrdlm2p1_ca_w_1_120_s_0_140 = '-3.40625e-07*ic_cap*ic_cap+-2.12500e-07*ic_cap+2.78000e-05'
+ mcrdlm2p1_ca_w_1_120_s_0_175 = '-3.40625e-07*ic_cap*ic_cap+-2.12500e-07*ic_cap+2.78000e-05'
+ mcrdlm2p1_ca_w_1_120_s_0_210 = '-3.40625e-07*ic_cap*ic_cap+-2.12500e-07*ic_cap+2.78000e-05'
+ mcrdlm2p1_ca_w_1_120_s_0_280 = '-3.40625e-07*ic_cap*ic_cap+-2.12500e-07*ic_cap+2.78000e-05'
+ mcrdlm2p1_ca_w_1_120_s_0_350 = '-3.40625e-07*ic_cap*ic_cap+-2.12500e-07*ic_cap+2.78000e-05'
+ mcrdlm2p1_ca_w_1_120_s_0_420 = '-3.40625e-07*ic_cap*ic_cap+-2.12500e-07*ic_cap+2.78000e-05'
+ mcrdlm2p1_ca_w_1_120_s_0_560 = '-3.40625e-07*ic_cap*ic_cap+-2.12500e-07*ic_cap+2.78000e-05'
+ mcrdlm2p1_ca_w_1_120_s_0_840 = '-3.40625e-07*ic_cap*ic_cap+-2.12500e-07*ic_cap+2.78000e-05'
+ mcrdlm2p1_ca_w_1_120_s_1_540 = '-3.40625e-07*ic_cap*ic_cap+-2.12500e-07*ic_cap+2.78000e-05'
+ mcrdlm2p1_ca_w_1_120_s_3_500 = '-3.40625e-07*ic_cap*ic_cap+-2.12500e-07*ic_cap+2.78000e-05'
+ mcrdlm2p1_cc_w_0_140_s_0_140 = '-9.40625e-13*ic_cap*ic_cap+-5.37500e-13*ic_cap+1.05000e-10'
+ mcrdlm2p1_cc_w_0_140_s_0_175 = '-9.09375e-13*ic_cap*ic_cap+-5.37500e-13*ic_cap+1.03000e-10'
+ mcrdlm2p1_cc_w_0_140_s_0_210 = '-7.78125e-13*ic_cap*ic_cap+-4.12500e-13*ic_cap+9.76000e-11'
+ mcrdlm2p1_cc_w_0_140_s_0_280 = '-6.00000e-13*ic_cap*ic_cap+-2.75000e-13*ic_cap+8.67000e-11'
+ mcrdlm2p1_cc_w_0_140_s_0_350 = '-4.50000e-13*ic_cap*ic_cap+-2.75000e-13*ic_cap+7.54000e-11'
+ mcrdlm2p1_cc_w_0_140_s_0_420 = '-3.62500e-13*ic_cap*ic_cap+-1.75000e-13*ic_cap+6.64000e-11'
+ mcrdlm2p1_cc_w_0_140_s_0_560 = '-1.90625e-13*ic_cap*ic_cap+-1.37500e-13*ic_cap+5.33000e-11'
+ mcrdlm2p1_cc_w_0_140_s_0_840 = '-5.93750e-14*ic_cap*ic_cap+-6.25000e-14*ic_cap+3.90000e-11'
+ mcrdlm2p1_cc_w_0_140_s_1_540 = '4.06250e-14*ic_cap*ic_cap+1.25000e-14*ic_cap+2.28000e-11'
+ mcrdlm2p1_cc_w_0_140_s_3_500 = '7.12500e-14*ic_cap*ic_cap+4.50000e-14*ic_cap+8.01000e-12'
+ mcrdlm2p1_cc_w_1_120_s_0_140 = '-8.12500e-13*ic_cap*ic_cap+-5.00000e-13*ic_cap+1.29000e-10'
+ mcrdlm2p1_cc_w_1_120_s_0_175 = '-7.18750e-13*ic_cap*ic_cap+-3.75000e-13*ic_cap+1.25000e-10'
+ mcrdlm2p1_cc_w_1_120_s_0_210 = '-6.56250e-13*ic_cap*ic_cap+-3.75000e-13*ic_cap+1.19000e-10'
+ mcrdlm2p1_cc_w_1_120_s_0_280 = '-4.81250e-13*ic_cap*ic_cap+-3.75000e-13*ic_cap+1.05000e-10'
+ mcrdlm2p1_cc_w_1_120_s_0_350 = '-3.68750e-13*ic_cap*ic_cap+-2.00000e-13*ic_cap+9.25000e-11'
+ mcrdlm2p1_cc_w_1_120_s_0_420 = '-2.40625e-13*ic_cap*ic_cap+-1.87500e-13*ic_cap+8.15000e-11'
+ mcrdlm2p1_cc_w_1_120_s_0_560 = '-1.03125e-13*ic_cap*ic_cap+-6.25000e-14*ic_cap+6.62000e-11'
+ mcrdlm2p1_cc_w_1_120_s_0_840 = '3.12500e-15*ic_cap*ic_cap+-1.25000e-14*ic_cap+4.91000e-11'
+ mcrdlm2p1_cc_w_1_120_s_1_540 = '1.00000e-13*ic_cap*ic_cap+5.00000e-14*ic_cap+2.95000e-11'
+ mcrdlm2p1_cc_w_1_120_s_3_500 = '1.03125e-13*ic_cap*ic_cap+6.25000e-14*ic_cap+1.13000e-11'
+ mcrdlm2p1_cf_w_0_140_s_0_140 = '-5.93750e-15*ic_cap*ic_cap+-3.75000e-15*ic_cap+1.94000e-12'
+ mcrdlm2p1_cf_w_0_140_s_0_175 = '-1.15625e-14*ic_cap*ic_cap+-8.75000e-15*ic_cap+2.42000e-12'
+ mcrdlm2p1_cf_w_0_140_s_0_210 = '-1.75000e-14*ic_cap*ic_cap+-1.25000e-14*ic_cap+2.91000e-12'
+ mcrdlm2p1_cf_w_0_140_s_0_280 = '-2.96875e-14*ic_cap*ic_cap+-1.87500e-14*ic_cap+3.86000e-12'
+ mcrdlm2p1_cf_w_0_140_s_0_350 = '-4.06250e-14*ic_cap*ic_cap+-2.50000e-14*ic_cap+4.79000e-12'
+ mcrdlm2p1_cf_w_0_140_s_0_420 = '-5.21875e-14*ic_cap*ic_cap+-3.37500e-14*ic_cap+5.76000e-12'
+ mcrdlm2p1_cf_w_0_140_s_0_560 = '-7.34375e-14*ic_cap*ic_cap+-4.37500e-14*ic_cap+7.53000e-12'
+ mcrdlm2p1_cf_w_0_140_s_0_840 = '-1.14062e-13*ic_cap*ic_cap+-6.62500e-14*ic_cap+1.09000e-11'
+ mcrdlm2p1_cf_w_0_140_s_1_540 = '-1.78125e-13*ic_cap*ic_cap+-1.12500e-13*ic_cap+1.78000e-11'
+ mcrdlm2p1_cf_w_0_140_s_3_500 = '-2.40625e-13*ic_cap*ic_cap+-1.62500e-13*ic_cap+2.86000e-11'
+ mcrdlm2p1_cf_w_1_120_s_0_140 = '-7.81250e-15*ic_cap*ic_cap+-6.25000e-15*ic_cap+2.02000e-12'
+ mcrdlm2p1_cf_w_1_120_s_0_175 = '-1.28125e-14*ic_cap*ic_cap+-8.75000e-15*ic_cap+2.49000e-12'
+ mcrdlm2p1_cf_w_1_120_s_0_210 = '-1.87500e-14*ic_cap*ic_cap+-1.25000e-14*ic_cap+2.97000e-12'
+ mcrdlm2p1_cf_w_1_120_s_0_280 = '-3.00000e-14*ic_cap*ic_cap+-2.00000e-14*ic_cap+3.92000e-12'
+ mcrdlm2p1_cf_w_1_120_s_0_350 = '-4.15625e-14*ic_cap*ic_cap+-2.62500e-14*ic_cap+4.87000e-12'
+ mcrdlm2p1_cf_w_1_120_s_0_420 = '-5.25000e-14*ic_cap*ic_cap+-3.25000e-14*ic_cap+5.79000e-12'
+ mcrdlm2p1_cf_w_1_120_s_0_560 = '-7.43750e-14*ic_cap*ic_cap+-4.50000e-14*ic_cap+7.60000e-12'
+ mcrdlm2p1_cf_w_1_120_s_0_840 = '-1.12813e-13*ic_cap*ic_cap+-6.87500e-14*ic_cap+1.10000e-11'
+ mcrdlm2p1_cf_w_1_120_s_1_540 = '-1.78125e-13*ic_cap*ic_cap+-1.12500e-13*ic_cap+1.82000e-11'
+ mcrdlm2p1_cf_w_1_120_s_3_500 = '-2.40625e-13*ic_cap*ic_cap+-1.62500e-13*ic_cap+3.04000e-11'
+ mcrdlm3_ca_w_10_000_s_10_000 = '-3.25000e-08*ic_cap*ic_cap+-2.00000e-08*ic_cap+3.50000e-06'
+ mcrdlm3_ca_w_10_000_s_12_000 = '-3.25000e-08*ic_cap*ic_cap+-2.00000e-08*ic_cap+3.50000e-06'
+ mcrdlm3_ca_w_10_000_s_30_000 = '-3.25000e-08*ic_cap*ic_cap+-2.00000e-08*ic_cap+3.50000e-06'
+ mcrdlm3_ca_w_10_000_s_5_000 = '-3.25000e-08*ic_cap*ic_cap+-2.00000e-08*ic_cap+3.50000e-06'
+ mcrdlm3_ca_w_10_000_s_8_000 = '-3.25000e-08*ic_cap*ic_cap+-2.00000e-08*ic_cap+3.50000e-06'
+ mcrdlm3_ca_w_40_000_s_10_000 = '-3.25000e-08*ic_cap*ic_cap+-2.00000e-08*ic_cap+3.50000e-06'
+ mcrdlm3_ca_w_40_000_s_12_000 = '-3.25000e-08*ic_cap*ic_cap+-2.00000e-08*ic_cap+3.50000e-06'
+ mcrdlm3_ca_w_40_000_s_30_000 = '-3.25000e-08*ic_cap*ic_cap+-2.00000e-08*ic_cap+3.50000e-06'
+ mcrdlm3_ca_w_40_000_s_5_000 = '-3.25000e-08*ic_cap*ic_cap+-2.00000e-08*ic_cap+3.50000e-06'
+ mcrdlm3_ca_w_40_000_s_8_000 = '-3.25000e-08*ic_cap*ic_cap+-2.00000e-08*ic_cap+3.50000e-06'
+ mcrdlm3_cc_w_10_000_s_10_000 = '-2.37500e-13*ic_cap*ic_cap+-1.50000e-13*ic_cap+2.95000e-11'
+ mcrdlm3_cc_w_10_000_s_12_000 = '-1.87500e-13*ic_cap*ic_cap+-1.25000e-13*ic_cap+2.55000e-11'
+ mcrdlm3_cc_w_10_000_s_30_000 = '-6.31250e-14*ic_cap*ic_cap+-4.00000e-14*ic_cap+1.06000e-11'
+ mcrdlm3_cc_w_10_000_s_5_000 = '-5.53125e-13*ic_cap*ic_cap+-3.37500e-13*ic_cap+4.89000e-11'
+ mcrdlm3_cc_w_10_000_s_8_000 = '-3.12500e-13*ic_cap*ic_cap+-2.00000e-13*ic_cap+3.49000e-11'
+ mcrdlm3_cc_w_40_000_s_10_000 = '-2.37500e-13*ic_cap*ic_cap+-1.50000e-13*ic_cap+3.93000e-11'
+ mcrdlm3_cc_w_40_000_s_12_000 = '-1.93750e-13*ic_cap*ic_cap+-1.25000e-13*ic_cap+3.50000e-11'
+ mcrdlm3_cc_w_40_000_s_30_000 = '-6.25000e-14*ic_cap*ic_cap+-5.00000e-14*ic_cap+1.77000e-11'
+ mcrdlm3_cc_w_40_000_s_5_000 = '-5.59375e-13*ic_cap*ic_cap+-3.37500e-13*ic_cap+6.02000e-11'
+ mcrdlm3_cc_w_40_000_s_8_000 = '-3.12500e-13*ic_cap*ic_cap+-2.00000e-13*ic_cap+4.52000e-11'
+ mcrdlm3_cf_w_10_000_s_10_000 = '-5.93750e-14*ic_cap*ic_cap+-3.75000e-14*ic_cap+1.39000e-11'
+ mcrdlm3_cf_w_10_000_s_12_000 = '-7.50000e-14*ic_cap*ic_cap+-5.00000e-14*ic_cap+1.59000e-11'
+ mcrdlm3_cf_w_10_000_s_30_000 = '-1.50000e-13*ic_cap*ic_cap+-1.00000e-13*ic_cap+2.67000e-11'
+ mcrdlm3_cf_w_10_000_s_5_000 = '-6.25000e-15*ic_cap*ic_cap+-2.50000e-15*ic_cap+7.87000e-12'
+ mcrdlm3_cf_w_10_000_s_8_000 = '-4.37500e-14*ic_cap*ic_cap+-2.50000e-14*ic_cap+1.17000e-11'
+ mcrdlm3_cf_w_40_000_s_10_000 = '-6.56250e-14*ic_cap*ic_cap+-3.75000e-14*ic_cap+1.40000e-11'
+ mcrdlm3_cf_w_40_000_s_12_000 = '-7.81250e-14*ic_cap*ic_cap+-3.75000e-14*ic_cap+1.60000e-11'
+ mcrdlm3_cf_w_40_000_s_30_000 = '-1.53125e-13*ic_cap*ic_cap+-8.75000e-14*ic_cap+2.77000e-11'
+ mcrdlm3_cf_w_40_000_s_5_000 = '-1.28125e-14*ic_cap*ic_cap+1.25000e-15*ic_cap+7.93000e-12'
+ mcrdlm3_cf_w_40_000_s_8_000 = '-5.00000e-14*ic_cap*ic_cap+-2.50000e-14*ic_cap+1.18000e-11'
+ mcrdlm3d_ca_w_0_300_s_0_300 = '-1.71875e-07*ic_cap*ic_cap+-1.12500e-07*ic_cap+1.77000e-05'
+ mcrdlm3d_ca_w_0_300_s_0_360 = '-1.71875e-07*ic_cap*ic_cap+-1.12500e-07*ic_cap+1.77000e-05'
+ mcrdlm3d_ca_w_0_300_s_0_450 = '-1.71875e-07*ic_cap*ic_cap+-1.12500e-07*ic_cap+1.77000e-05'
+ mcrdlm3d_ca_w_0_300_s_0_600 = '-1.71875e-07*ic_cap*ic_cap+-1.12500e-07*ic_cap+1.77000e-05'
+ mcrdlm3d_ca_w_0_300_s_0_800 = '-1.71875e-07*ic_cap*ic_cap+-1.12500e-07*ic_cap+1.77000e-05'
+ mcrdlm3d_ca_w_0_300_s_1_000 = '-1.71875e-07*ic_cap*ic_cap+-1.12500e-07*ic_cap+1.77000e-05'
+ mcrdlm3d_ca_w_0_300_s_1_200 = '-1.71875e-07*ic_cap*ic_cap+-1.12500e-07*ic_cap+1.77000e-05'
+ mcrdlm3d_ca_w_0_300_s_2_100 = '-1.71875e-07*ic_cap*ic_cap+-1.12500e-07*ic_cap+1.77000e-05'
+ mcrdlm3d_ca_w_0_300_s_3_300 = '-1.71875e-07*ic_cap*ic_cap+-1.12500e-07*ic_cap+1.77000e-05'
+ mcrdlm3d_ca_w_0_300_s_9_000 = '-1.71875e-07*ic_cap*ic_cap+-1.12500e-07*ic_cap+1.77000e-05'
+ mcrdlm3d_ca_w_2_400_s_0_300 = '-1.71875e-07*ic_cap*ic_cap+-1.12500e-07*ic_cap+1.77000e-05'
+ mcrdlm3d_ca_w_2_400_s_0_360 = '-1.71875e-07*ic_cap*ic_cap+-1.12500e-07*ic_cap+1.77000e-05'
+ mcrdlm3d_ca_w_2_400_s_0_450 = '-1.71875e-07*ic_cap*ic_cap+-1.12500e-07*ic_cap+1.77000e-05'
+ mcrdlm3d_ca_w_2_400_s_0_600 = '-1.71875e-07*ic_cap*ic_cap+-1.12500e-07*ic_cap+1.77000e-05'
+ mcrdlm3d_ca_w_2_400_s_0_800 = '-1.71875e-07*ic_cap*ic_cap+-1.12500e-07*ic_cap+1.77000e-05'
+ mcrdlm3d_ca_w_2_400_s_1_000 = '-1.71875e-07*ic_cap*ic_cap+-1.12500e-07*ic_cap+1.77000e-05'
+ mcrdlm3d_ca_w_2_400_s_1_200 = '-1.71875e-07*ic_cap*ic_cap+-1.12500e-07*ic_cap+1.77000e-05'
+ mcrdlm3d_ca_w_2_400_s_2_100 = '-1.71875e-07*ic_cap*ic_cap+-1.12500e-07*ic_cap+1.77000e-05'
+ mcrdlm3d_ca_w_2_400_s_3_300 = '-1.71875e-07*ic_cap*ic_cap+-1.12500e-07*ic_cap+1.77000e-05'
+ mcrdlm3d_ca_w_2_400_s_9_000 = '-1.71875e-07*ic_cap*ic_cap+-1.12500e-07*ic_cap+1.77000e-05'
+ mcrdlm3d_cc_w_0_300_s_0_300 = '-7.53125e-13*ic_cap*ic_cap+-4.37500e-13*ic_cap+1.05000e-10'
+ mcrdlm3d_cc_w_0_300_s_0_360 = '-7.00000e-13*ic_cap*ic_cap+-4.25000e-13*ic_cap+9.83000e-11'
+ mcrdlm3d_cc_w_0_300_s_0_450 = '-5.90625e-13*ic_cap*ic_cap+-3.62500e-13*ic_cap+8.86000e-11'
+ mcrdlm3d_cc_w_0_300_s_0_600 = '-4.46875e-13*ic_cap*ic_cap+-2.62500e-13*ic_cap+7.58000e-11'
+ mcrdlm3d_cc_w_0_300_s_0_800 = '-2.93750e-13*ic_cap*ic_cap+-2.25000e-13*ic_cap+6.31000e-11'
+ mcrdlm3d_cc_w_0_300_s_1_000 = '-2.06250e-13*ic_cap*ic_cap+-1.50000e-13*ic_cap+5.37000e-11'
+ mcrdlm3d_cc_w_0_300_s_1_200 = '-1.50000e-13*ic_cap*ic_cap+-1.00000e-13*ic_cap+4.67000e-11'
+ mcrdlm3d_cc_w_0_300_s_2_100 = '-3.12500e-14*ic_cap*ic_cap+-2.50000e-14*ic_cap+2.87000e-11'
+ mcrdlm3d_cc_w_0_300_s_3_300 = '2.81250e-14*ic_cap*ic_cap+1.25000e-14*ic_cap+1.78000e-11'
+ mcrdlm3d_cc_w_0_300_s_9_000 = '3.62500e-14*ic_cap*ic_cap+2.50000e-14*ic_cap+2.89000e-12'
+ mcrdlm3d_cc_w_2_400_s_0_300 = '-6.56250e-13*ic_cap*ic_cap+-3.75000e-13*ic_cap+1.26000e-10'
+ mcrdlm3d_cc_w_2_400_s_0_360 = '-5.93750e-13*ic_cap*ic_cap+-3.75000e-13*ic_cap+1.18000e-10'
+ mcrdlm3d_cc_w_2_400_s_0_450 = '-4.75000e-13*ic_cap*ic_cap+-4.00000e-13*ic_cap+1.07000e-10'
+ mcrdlm3d_cc_w_2_400_s_0_600 = '-3.37500e-13*ic_cap*ic_cap+-2.00000e-13*ic_cap+9.19000e-11'
+ mcrdlm3d_cc_w_2_400_s_0_800 = '-2.00000e-13*ic_cap*ic_cap+-1.25000e-13*ic_cap+7.69000e-11'
+ mcrdlm3d_cc_w_2_400_s_1_000 = '-1.28125e-13*ic_cap*ic_cap+-8.75000e-14*ic_cap+6.59000e-11'
+ mcrdlm3d_cc_w_2_400_s_1_200 = '-7.18750e-14*ic_cap*ic_cap+-6.25000e-14*ic_cap+5.75000e-11'
+ mcrdlm3d_cc_w_2_400_s_2_100 = '3.12500e-14*ic_cap*ic_cap+2.50000e-14*ic_cap+3.62000e-11'
+ mcrdlm3d_cc_w_2_400_s_3_300 = '7.81250e-14*ic_cap*ic_cap+3.75000e-14*ic_cap+2.27000e-11'
+ mcrdlm3d_cc_w_2_400_s_9_000 = '5.84375e-14*ic_cap*ic_cap+3.87500e-14*ic_cap+4.01000e-12'
+ mcrdlm3d_cf_w_0_300_s_0_300 = '-6.25000e-15*ic_cap*ic_cap+-5.00000e-15*ic_cap+2.61000e-12'
+ mcrdlm3d_cf_w_0_300_s_0_360 = '-1.12500e-14*ic_cap*ic_cap+-7.50000e-15*ic_cap+3.13000e-12'
+ mcrdlm3d_cf_w_0_300_s_0_450 = '-1.81250e-14*ic_cap*ic_cap+-1.25000e-14*ic_cap+3.92000e-12'
+ mcrdlm3d_cf_w_0_300_s_0_600 = '-3.00000e-14*ic_cap*ic_cap+-1.75000e-14*ic_cap+5.21000e-12'
+ mcrdlm3d_cf_w_0_300_s_0_800 = '-4.56250e-14*ic_cap*ic_cap+-3.00000e-14*ic_cap+6.76000e-12'
+ mcrdlm3d_cf_w_0_300_s_1_000 = '-6.00000e-14*ic_cap*ic_cap+-3.75000e-14*ic_cap+8.33000e-12'
+ mcrdlm3d_cf_w_0_300_s_1_200 = '-7.34375e-14*ic_cap*ic_cap+-4.62500e-14*ic_cap+9.85000e-12'
+ mcrdlm3d_cf_w_0_300_s_2_100 = '-1.25000e-13*ic_cap*ic_cap+-7.50000e-14*ic_cap+1.62000e-11'
+ mcrdlm3d_cf_w_0_300_s_3_300 = '-1.65625e-13*ic_cap*ic_cap+-1.12500e-13*ic_cap+2.21000e-11'
+ mcrdlm3d_cf_w_0_300_s_9_000 = '-1.93750e-13*ic_cap*ic_cap+-1.25000e-13*ic_cap+3.39000e-11'
+ mcrdlm3d_cf_w_2_400_s_0_300 = '-7.50000e-15*ic_cap*ic_cap+-5.00000e-15*ic_cap+2.67000e-12'
+ mcrdlm3d_cf_w_2_400_s_0_360 = '-1.21875e-14*ic_cap*ic_cap+-8.75000e-15*ic_cap+3.18000e-12'
+ mcrdlm3d_cf_w_2_400_s_0_450 = '-1.90625e-14*ic_cap*ic_cap+-1.37500e-14*ic_cap+3.94000e-12'
+ mcrdlm3d_cf_w_2_400_s_0_600 = '-3.12500e-14*ic_cap*ic_cap+-2.00000e-14*ic_cap+5.20000e-12'
+ mcrdlm3d_cf_w_2_400_s_0_800 = '-4.56250e-14*ic_cap*ic_cap+-3.00000e-14*ic_cap+6.83000e-12'
+ mcrdlm3d_cf_w_2_400_s_1_000 = '-6.09375e-14*ic_cap*ic_cap+-3.87500e-14*ic_cap+8.43000e-12'
+ mcrdlm3d_cf_w_2_400_s_1_200 = '-7.43750e-14*ic_cap*ic_cap+-4.75000e-14*ic_cap+9.97000e-12'
+ mcrdlm3d_cf_w_2_400_s_2_100 = '-1.25000e-13*ic_cap*ic_cap+-7.50000e-14*ic_cap+1.62000e-11'
+ mcrdlm3d_cf_w_2_400_s_3_300 = '-1.71875e-13*ic_cap*ic_cap+-1.12500e-13*ic_cap+2.29000e-11'
+ mcrdlm3d_cf_w_2_400_s_9_000 = '-1.87500e-13*ic_cap*ic_cap+-1.25000e-13*ic_cap+3.71000e-11'
+ mcrdlm3f_ca_w_0_300_s_0_300 = '-1.62500e-07*ic_cap*ic_cap+-1.00000e-07*ic_cap+1.61000e-05'
+ mcrdlm3f_ca_w_0_300_s_0_360 = '-1.62500e-07*ic_cap*ic_cap+-1.00000e-07*ic_cap+1.61000e-05'
+ mcrdlm3f_ca_w_0_300_s_0_450 = '-1.62500e-07*ic_cap*ic_cap+-1.00000e-07*ic_cap+1.61000e-05'
+ mcrdlm3f_ca_w_0_300_s_0_600 = '-1.62500e-07*ic_cap*ic_cap+-1.00000e-07*ic_cap+1.61000e-05'
+ mcrdlm3f_ca_w_0_300_s_0_800 = '-1.62500e-07*ic_cap*ic_cap+-1.00000e-07*ic_cap+1.61000e-05'
+ mcrdlm3f_ca_w_0_300_s_1_000 = '-1.62500e-07*ic_cap*ic_cap+-1.00000e-07*ic_cap+1.61000e-05'
+ mcrdlm3f_ca_w_0_300_s_1_200 = '-1.62500e-07*ic_cap*ic_cap+-1.00000e-07*ic_cap+1.61000e-05'
+ mcrdlm3f_ca_w_0_300_s_2_100 = '-1.62500e-07*ic_cap*ic_cap+-1.00000e-07*ic_cap+1.61000e-05'
+ mcrdlm3f_ca_w_0_300_s_3_300 = '-1.62500e-07*ic_cap*ic_cap+-1.00000e-07*ic_cap+1.61000e-05'
+ mcrdlm3f_ca_w_0_300_s_9_000 = '-1.62500e-07*ic_cap*ic_cap+-1.00000e-07*ic_cap+1.61000e-05'
+ mcrdlm3f_ca_w_2_400_s_0_300 = '-1.62500e-07*ic_cap*ic_cap+-1.00000e-07*ic_cap+1.61000e-05'
+ mcrdlm3f_ca_w_2_400_s_0_360 = '-1.62500e-07*ic_cap*ic_cap+-1.00000e-07*ic_cap+1.61000e-05'
+ mcrdlm3f_ca_w_2_400_s_0_450 = '-1.62500e-07*ic_cap*ic_cap+-1.00000e-07*ic_cap+1.61000e-05'
+ mcrdlm3f_ca_w_2_400_s_0_600 = '-1.62500e-07*ic_cap*ic_cap+-1.00000e-07*ic_cap+1.61000e-05'
+ mcrdlm3f_ca_w_2_400_s_0_800 = '-1.62500e-07*ic_cap*ic_cap+-1.00000e-07*ic_cap+1.61000e-05'
+ mcrdlm3f_ca_w_2_400_s_1_000 = '-1.62500e-07*ic_cap*ic_cap+-1.00000e-07*ic_cap+1.61000e-05'
+ mcrdlm3f_ca_w_2_400_s_1_200 = '-1.62500e-07*ic_cap*ic_cap+-1.00000e-07*ic_cap+1.61000e-05'
+ mcrdlm3f_ca_w_2_400_s_2_100 = '-1.62500e-07*ic_cap*ic_cap+-1.00000e-07*ic_cap+1.61000e-05'
+ mcrdlm3f_ca_w_2_400_s_3_300 = '-1.62500e-07*ic_cap*ic_cap+-1.00000e-07*ic_cap+1.61000e-05'
+ mcrdlm3f_ca_w_2_400_s_9_000 = '-1.62500e-07*ic_cap*ic_cap+-1.00000e-07*ic_cap+1.61000e-05'
+ mcrdlm3f_cc_w_0_300_s_0_300 = '-8.03125e-13*ic_cap*ic_cap+-4.37500e-13*ic_cap+1.06000e-10'
+ mcrdlm3f_cc_w_0_300_s_0_360 = '-7.00000e-13*ic_cap*ic_cap+-4.25000e-13*ic_cap+9.87000e-11'
+ mcrdlm3f_cc_w_0_300_s_0_450 = '-5.96875e-13*ic_cap*ic_cap+-3.62500e-13*ic_cap+8.91000e-11'
+ mcrdlm3f_cc_w_0_300_s_0_600 = '-4.46875e-13*ic_cap*ic_cap+-2.62500e-13*ic_cap+7.63000e-11'
+ mcrdlm3f_cc_w_0_300_s_0_800 = '-3.00000e-13*ic_cap*ic_cap+-2.25000e-13*ic_cap+6.38000e-11'
+ mcrdlm3f_cc_w_0_300_s_1_000 = '-2.12500e-13*ic_cap*ic_cap+-1.50000e-13*ic_cap+5.45000e-11'
+ mcrdlm3f_cc_w_0_300_s_1_200 = '-1.53125e-13*ic_cap*ic_cap+-1.12500e-13*ic_cap+4.75000e-11'
+ mcrdlm3f_cc_w_0_300_s_2_100 = '-2.81250e-14*ic_cap*ic_cap+-3.75000e-14*ic_cap+2.96000e-11'
+ mcrdlm3f_cc_w_0_300_s_3_300 = '3.12500e-14*ic_cap*ic_cap+2.50000e-14*ic_cap+1.87000e-11'
+ mcrdlm3f_cc_w_0_300_s_9_000 = '4.15625e-14*ic_cap*ic_cap+2.87500e-14*ic_cap+3.26000e-12'
+ mcrdlm3f_cc_w_2_400_s_0_300 = '-7.18750e-13*ic_cap*ic_cap+-3.75000e-13*ic_cap+1.28000e-10'
+ mcrdlm3f_cc_w_2_400_s_0_360 = '-5.93750e-13*ic_cap*ic_cap+-3.75000e-13*ic_cap+1.19000e-10'
+ mcrdlm3f_cc_w_2_400_s_0_450 = '-4.68750e-13*ic_cap*ic_cap+-3.75000e-13*ic_cap+1.08000e-10'
+ mcrdlm3f_cc_w_2_400_s_0_600 = '-3.37500e-13*ic_cap*ic_cap+-2.00000e-13*ic_cap+9.31000e-11'
+ mcrdlm3f_cc_w_2_400_s_0_800 = '-1.96875e-13*ic_cap*ic_cap+-1.37500e-13*ic_cap+7.81000e-11'
+ mcrdlm3f_cc_w_2_400_s_1_000 = '-1.28125e-13*ic_cap*ic_cap+-8.75000e-14*ic_cap+6.72000e-11'
+ mcrdlm3f_cc_w_2_400_s_1_200 = '-6.56250e-14*ic_cap*ic_cap+-6.25000e-14*ic_cap+5.87000e-11'
+ mcrdlm3f_cc_w_2_400_s_2_100 = '4.37500e-14*ic_cap*ic_cap+2.50000e-14*ic_cap+3.74000e-11'
+ mcrdlm3f_cc_w_2_400_s_3_300 = '8.12500e-14*ic_cap*ic_cap+5.00000e-14*ic_cap+2.39000e-11'
+ mcrdlm3f_cc_w_2_400_s_9_000 = '6.71875e-14*ic_cap*ic_cap+5.12500e-14*ic_cap+4.48000e-12'
+ mcrdlm3f_cf_w_0_300_s_0_300 = '-6.87500e-15*ic_cap*ic_cap+-5.00000e-15*ic_cap+2.38000e-12'
+ mcrdlm3f_cf_w_0_300_s_0_360 = '-1.12500e-14*ic_cap*ic_cap+-7.50000e-15*ic_cap+2.85000e-12'
+ mcrdlm3f_cf_w_0_300_s_0_450 = '-1.84375e-14*ic_cap*ic_cap+-1.12500e-14*ic_cap+3.58000e-12'
+ mcrdlm3f_cf_w_0_300_s_0_600 = '-2.93750e-14*ic_cap*ic_cap+-1.75000e-14*ic_cap+4.76000e-12'
+ mcrdlm3f_cf_w_0_300_s_0_800 = '-4.37500e-14*ic_cap*ic_cap+-2.75000e-14*ic_cap+6.17000e-12'
+ mcrdlm3f_cf_w_0_300_s_1_000 = '-5.78125e-14*ic_cap*ic_cap+-3.62500e-14*ic_cap+7.62000e-12'
+ mcrdlm3f_cf_w_0_300_s_1_200 = '-7.09375e-14*ic_cap*ic_cap+-4.37500e-14*ic_cap+9.03000e-12'
+ mcrdlm3f_cf_w_0_300_s_2_100 = '-1.18750e-13*ic_cap*ic_cap+-7.50000e-14*ic_cap+1.49000e-11'
+ mcrdlm3f_cf_w_0_300_s_3_300 = '-1.62500e-13*ic_cap*ic_cap+-1.00000e-13*ic_cap+2.06000e-11'
+ mcrdlm3f_cf_w_0_300_s_9_000 = '-1.93750e-13*ic_cap*ic_cap+-1.25000e-13*ic_cap+3.25000e-11'
+ mcrdlm3f_cf_w_2_400_s_0_300 = '-8.12500e-15*ic_cap*ic_cap+-5.00000e-15*ic_cap+2.43000e-12'
+ mcrdlm3f_cf_w_2_400_s_0_360 = '-1.18750e-14*ic_cap*ic_cap+-7.50000e-15*ic_cap+2.89000e-12'
+ mcrdlm3f_cf_w_2_400_s_0_450 = '-1.90625e-14*ic_cap*ic_cap+-1.12500e-14*ic_cap+3.59000e-12'
+ mcrdlm3f_cf_w_2_400_s_0_600 = '-3.03125e-14*ic_cap*ic_cap+-1.87500e-14*ic_cap+4.74000e-12'
+ mcrdlm3f_cf_w_2_400_s_0_800 = '-4.46875e-14*ic_cap*ic_cap+-2.87500e-14*ic_cap+6.24000e-12'
+ mcrdlm3f_cf_w_2_400_s_1_000 = '-5.87500e-14*ic_cap*ic_cap+-3.75000e-14*ic_cap+7.71000e-12'
+ mcrdlm3f_cf_w_2_400_s_1_200 = '-7.18750e-14*ic_cap*ic_cap+-4.50000e-14*ic_cap+9.13000e-12'
+ mcrdlm3f_cf_w_2_400_s_2_100 = '-1.25000e-13*ic_cap*ic_cap+-7.50000e-14*ic_cap+1.50000e-11'
+ mcrdlm3f_cf_w_2_400_s_3_300 = '-1.65625e-13*ic_cap*ic_cap+-1.12500e-13*ic_cap+2.13000e-11'
+ mcrdlm3f_cf_w_2_400_s_9_000 = '-1.93750e-13*ic_cap*ic_cap+-1.25000e-13*ic_cap+3.56000e-11'
+ mcrdlm3l1_ca_w_0_300_s_0_300 = '-2.43750e-07*ic_cap*ic_cap+-1.50000e-07*ic_cap+2.37000e-05'
+ mcrdlm3l1_ca_w_0_300_s_0_360 = '-2.43750e-07*ic_cap*ic_cap+-1.50000e-07*ic_cap+2.37000e-05'
+ mcrdlm3l1_ca_w_0_300_s_0_450 = '-2.43750e-07*ic_cap*ic_cap+-1.50000e-07*ic_cap+2.37000e-05'
+ mcrdlm3l1_ca_w_0_300_s_0_600 = '-2.43750e-07*ic_cap*ic_cap+-1.50000e-07*ic_cap+2.37000e-05'
+ mcrdlm3l1_ca_w_0_300_s_0_800 = '-2.43750e-07*ic_cap*ic_cap+-1.50000e-07*ic_cap+2.37000e-05'
+ mcrdlm3l1_ca_w_0_300_s_1_000 = '-2.43750e-07*ic_cap*ic_cap+-1.50000e-07*ic_cap+2.37000e-05'
+ mcrdlm3l1_ca_w_0_300_s_1_200 = '-2.43750e-07*ic_cap*ic_cap+-1.50000e-07*ic_cap+2.37000e-05'
+ mcrdlm3l1_ca_w_0_300_s_2_100 = '-2.43750e-07*ic_cap*ic_cap+-1.50000e-07*ic_cap+2.37000e-05'
+ mcrdlm3l1_ca_w_0_300_s_3_300 = '-2.43750e-07*ic_cap*ic_cap+-1.50000e-07*ic_cap+2.37000e-05'
+ mcrdlm3l1_ca_w_0_300_s_9_000 = '-2.43750e-07*ic_cap*ic_cap+-1.50000e-07*ic_cap+2.37000e-05'
+ mcrdlm3l1_ca_w_2_400_s_0_300 = '-2.43750e-07*ic_cap*ic_cap+-1.50000e-07*ic_cap+2.37000e-05'
+ mcrdlm3l1_ca_w_2_400_s_0_360 = '-2.43750e-07*ic_cap*ic_cap+-1.50000e-07*ic_cap+2.37000e-05'
+ mcrdlm3l1_ca_w_2_400_s_0_450 = '-2.43750e-07*ic_cap*ic_cap+-1.50000e-07*ic_cap+2.37000e-05'
+ mcrdlm3l1_ca_w_2_400_s_0_600 = '-2.43750e-07*ic_cap*ic_cap+-1.50000e-07*ic_cap+2.37000e-05'
+ mcrdlm3l1_ca_w_2_400_s_0_800 = '-2.43750e-07*ic_cap*ic_cap+-1.50000e-07*ic_cap+2.37000e-05'
+ mcrdlm3l1_ca_w_2_400_s_1_000 = '-2.43750e-07*ic_cap*ic_cap+-1.50000e-07*ic_cap+2.37000e-05'
+ mcrdlm3l1_ca_w_2_400_s_1_200 = '-2.43750e-07*ic_cap*ic_cap+-1.50000e-07*ic_cap+2.37000e-05'
+ mcrdlm3l1_ca_w_2_400_s_2_100 = '-2.43750e-07*ic_cap*ic_cap+-1.50000e-07*ic_cap+2.37000e-05'
+ mcrdlm3l1_ca_w_2_400_s_3_300 = '-2.43750e-07*ic_cap*ic_cap+-1.50000e-07*ic_cap+2.37000e-05'
+ mcrdlm3l1_ca_w_2_400_s_9_000 = '-2.43750e-07*ic_cap*ic_cap+-1.50000e-07*ic_cap+2.37000e-05'
+ mcrdlm3l1_cc_w_0_300_s_0_300 = '-7.68750e-13*ic_cap*ic_cap+-4.25000e-13*ic_cap+1.04000e-10'
+ mcrdlm3l1_cc_w_0_300_s_0_360 = '-6.90625e-13*ic_cap*ic_cap+-4.37500e-13*ic_cap+9.68000e-11'
+ mcrdlm3l1_cc_w_0_300_s_0_450 = '-5.50000e-13*ic_cap*ic_cap+-3.00000e-13*ic_cap+8.67000e-11'
+ mcrdlm3l1_cc_w_0_300_s_0_600 = '-4.21875e-13*ic_cap*ic_cap+-2.62500e-13*ic_cap+7.38000e-11'
+ mcrdlm3l1_cc_w_0_300_s_0_800 = '-2.78125e-13*ic_cap*ic_cap+-2.12500e-13*ic_cap+6.09000e-11'
+ mcrdlm3l1_cc_w_0_300_s_1_000 = '-1.87500e-13*ic_cap*ic_cap+-1.25000e-13*ic_cap+5.13000e-11'
+ mcrdlm3l1_cc_w_0_300_s_1_200 = '-1.28125e-13*ic_cap*ic_cap+-8.75000e-14*ic_cap+4.41000e-11'
+ mcrdlm3l1_cc_w_0_300_s_2_100 = '-1.56250e-14*ic_cap*ic_cap+-1.25000e-14*ic_cap+2.59000e-11'
+ mcrdlm3l1_cc_w_0_300_s_3_300 = '3.75000e-14*ic_cap*ic_cap+2.50000e-14*ic_cap+1.51000e-11'
+ mcrdlm3l1_cc_w_0_300_s_9_000 = '2.68750e-14*ic_cap*ic_cap+2.00000e-14*ic_cap+2.07000e-12'
+ mcrdlm3l1_cc_w_2_400_s_0_300 = '-6.56250e-13*ic_cap*ic_cap+-3.75000e-13*ic_cap+1.23000e-10'
+ mcrdlm3l1_cc_w_2_400_s_0_360 = '-5.62500e-13*ic_cap*ic_cap+-2.50000e-13*ic_cap+1.14000e-10'
+ mcrdlm3l1_cc_w_2_400_s_0_450 = '-4.59375e-13*ic_cap*ic_cap+-2.87500e-13*ic_cap+1.03000e-10'
+ mcrdlm3l1_cc_w_2_400_s_0_600 = '-3.25000e-13*ic_cap*ic_cap+-1.75000e-13*ic_cap+8.82000e-11'
+ mcrdlm3l1_cc_w_2_400_s_0_800 = '-1.84375e-13*ic_cap*ic_cap+-1.12500e-13*ic_cap+7.31000e-11'
+ mcrdlm3l1_cc_w_2_400_s_1_000 = '-1.18750e-13*ic_cap*ic_cap+-7.50000e-14*ic_cap+6.22000e-11'
+ mcrdlm3l1_cc_w_2_400_s_1_200 = '-5.62500e-14*ic_cap*ic_cap+-5.00000e-14*ic_cap+5.38000e-11'
+ mcrdlm3l1_cc_w_2_400_s_2_100 = '3.75000e-14*ic_cap*ic_cap+2.50000e-14*ic_cap+3.28000e-11'
+ mcrdlm3l1_cc_w_2_400_s_3_300 = '7.50000e-14*ic_cap*ic_cap+5.00000e-14*ic_cap+1.97000e-11'
+ mcrdlm3l1_cc_w_2_400_s_9_000 = '4.56250e-14*ic_cap*ic_cap+3.00000e-14*ic_cap+3.00000e-12'
+ mcrdlm3l1_cf_w_0_300_s_0_300 = '-1.06250e-14*ic_cap*ic_cap+-7.50000e-15*ic_cap+3.47000e-12'
+ mcrdlm3l1_cf_w_0_300_s_0_360 = '-1.75000e-14*ic_cap*ic_cap+-1.25000e-14*ic_cap+4.15000e-12'
+ mcrdlm3l1_cf_w_0_300_s_0_450 = '-2.71875e-14*ic_cap*ic_cap+-1.87500e-14*ic_cap+5.18000e-12'
+ mcrdlm3l1_cf_w_0_300_s_0_600 = '-4.28125e-14*ic_cap*ic_cap+-2.87500e-14*ic_cap+6.84000e-12'
+ mcrdlm3l1_cf_w_0_300_s_0_800 = '-6.34375e-14*ic_cap*ic_cap+-4.12500e-14*ic_cap+8.86000e-12'
+ mcrdlm3l1_cf_w_0_300_s_1_000 = '-8.56250e-14*ic_cap*ic_cap+-5.00000e-14*ic_cap+1.09000e-11'
+ mcrdlm3l1_cf_w_0_300_s_1_200 = '-1.03125e-13*ic_cap*ic_cap+-6.25000e-14*ic_cap+1.28000e-11'
+ mcrdlm3l1_cf_w_0_300_s_2_100 = '-1.62500e-13*ic_cap*ic_cap+-1.00000e-13*ic_cap+2.04000e-11'
+ mcrdlm3l1_cf_w_0_300_s_3_300 = '-2.03125e-13*ic_cap*ic_cap+-1.37500e-13*ic_cap+2.70000e-11'
+ mcrdlm3l1_cf_w_0_300_s_9_000 = '-2.09375e-13*ic_cap*ic_cap+-1.37500e-13*ic_cap+3.80000e-11'
+ mcrdlm3l1_cf_w_2_400_s_0_300 = '-1.12500e-14*ic_cap*ic_cap+-7.50000e-15*ic_cap+3.52000e-12'
+ mcrdlm3l1_cf_w_2_400_s_0_360 = '-1.84375e-14*ic_cap*ic_cap+-1.37500e-14*ic_cap+4.20000e-12'
+ mcrdlm3l1_cf_w_2_400_s_0_450 = '-2.81250e-14*ic_cap*ic_cap+-2.00000e-14*ic_cap+5.20000e-12'
+ mcrdlm3l1_cf_w_2_400_s_0_600 = '-4.37500e-14*ic_cap*ic_cap+-2.75000e-14*ic_cap+6.83000e-12'
+ mcrdlm3l1_cf_w_2_400_s_0_800 = '-6.37500e-14*ic_cap*ic_cap+-4.25000e-14*ic_cap+8.94000e-12'
+ mcrdlm3l1_cf_w_2_400_s_1_000 = '-8.40625e-14*ic_cap*ic_cap+-5.37500e-14*ic_cap+1.10000e-11'
+ mcrdlm3l1_cf_w_2_400_s_1_200 = '-1.00000e-13*ic_cap*ic_cap+-7.50000e-14*ic_cap+1.29000e-11'
+ mcrdlm3l1_cf_w_2_400_s_2_100 = '-1.59375e-13*ic_cap*ic_cap+-1.12500e-13*ic_cap+2.05000e-11'
+ mcrdlm3l1_cf_w_2_400_s_3_300 = '-2.03125e-13*ic_cap*ic_cap+-1.37500e-13*ic_cap+2.80000e-11'
+ mcrdlm3l1_cf_w_2_400_s_9_000 = '-1.96875e-13*ic_cap*ic_cap+-1.37500e-13*ic_cap+4.15000e-11'
+ mcrdlm3m1_ca_w_0_300_s_0_300 = '-4.21875e-07*ic_cap*ic_cap+-2.37500e-07*ic_cap+3.64000e-05'
+ mcrdlm3m1_ca_w_0_300_s_0_360 = '-4.21875e-07*ic_cap*ic_cap+-2.37500e-07*ic_cap+3.64000e-05'
+ mcrdlm3m1_ca_w_0_300_s_0_450 = '-4.21875e-07*ic_cap*ic_cap+-2.37500e-07*ic_cap+3.64000e-05'
+ mcrdlm3m1_ca_w_0_300_s_0_600 = '-4.21875e-07*ic_cap*ic_cap+-2.37500e-07*ic_cap+3.64000e-05'
+ mcrdlm3m1_ca_w_0_300_s_0_800 = '-4.21875e-07*ic_cap*ic_cap+-2.37500e-07*ic_cap+3.64000e-05'
+ mcrdlm3m1_ca_w_0_300_s_1_000 = '-4.21875e-07*ic_cap*ic_cap+-2.37500e-07*ic_cap+3.64000e-05'
+ mcrdlm3m1_ca_w_0_300_s_1_200 = '-4.21875e-07*ic_cap*ic_cap+-2.37500e-07*ic_cap+3.64000e-05'
+ mcrdlm3m1_ca_w_0_300_s_2_100 = '-4.21875e-07*ic_cap*ic_cap+-2.37500e-07*ic_cap+3.64000e-05'
+ mcrdlm3m1_ca_w_0_300_s_3_300 = '-4.21875e-07*ic_cap*ic_cap+-2.37500e-07*ic_cap+3.64000e-05'
+ mcrdlm3m1_ca_w_0_300_s_9_000 = '-4.21875e-07*ic_cap*ic_cap+-2.37500e-07*ic_cap+3.64000e-05'
+ mcrdlm3m1_ca_w_2_400_s_0_300 = '-4.21875e-07*ic_cap*ic_cap+-2.37500e-07*ic_cap+3.64000e-05'
+ mcrdlm3m1_ca_w_2_400_s_0_360 = '-4.21875e-07*ic_cap*ic_cap+-2.37500e-07*ic_cap+3.64000e-05'
+ mcrdlm3m1_ca_w_2_400_s_0_450 = '-4.21875e-07*ic_cap*ic_cap+-2.37500e-07*ic_cap+3.64000e-05'
+ mcrdlm3m1_ca_w_2_400_s_0_600 = '-4.21875e-07*ic_cap*ic_cap+-2.37500e-07*ic_cap+3.64000e-05'
+ mcrdlm3m1_ca_w_2_400_s_0_800 = '-4.21875e-07*ic_cap*ic_cap+-2.37500e-07*ic_cap+3.64000e-05'
+ mcrdlm3m1_ca_w_2_400_s_1_000 = '-4.21875e-07*ic_cap*ic_cap+-2.37500e-07*ic_cap+3.64000e-05'
+ mcrdlm3m1_ca_w_2_400_s_1_200 = '-4.21875e-07*ic_cap*ic_cap+-2.37500e-07*ic_cap+3.64000e-05'
+ mcrdlm3m1_ca_w_2_400_s_2_100 = '-4.21875e-07*ic_cap*ic_cap+-2.37500e-07*ic_cap+3.64000e-05'
+ mcrdlm3m1_ca_w_2_400_s_3_300 = '-4.21875e-07*ic_cap*ic_cap+-2.37500e-07*ic_cap+3.64000e-05'
+ mcrdlm3m1_ca_w_2_400_s_9_000 = '-4.21875e-07*ic_cap*ic_cap+-2.37500e-07*ic_cap+3.64000e-05'
+ mcrdlm3m1_cc_w_0_300_s_0_300 = '-7.28125e-13*ic_cap*ic_cap+-4.37500e-13*ic_cap+1.01000e-10'
+ mcrdlm3m1_cc_w_0_300_s_0_360 = '-6.46875e-13*ic_cap*ic_cap+-4.12500e-13*ic_cap+9.37000e-11'
+ mcrdlm3m1_cc_w_0_300_s_0_450 = '-5.18750e-13*ic_cap*ic_cap+-3.00000e-13*ic_cap+8.35000e-11'
+ mcrdlm3m1_cc_w_0_300_s_0_600 = '-3.75000e-13*ic_cap*ic_cap+-2.25000e-13*ic_cap+7.01000e-11'
+ mcrdlm3m1_cc_w_0_300_s_0_800 = '-2.40625e-13*ic_cap*ic_cap+-1.87500e-13*ic_cap+5.70000e-11'
+ mcrdlm3m1_cc_w_0_300_s_1_000 = '-1.53125e-13*ic_cap*ic_cap+-1.12500e-13*ic_cap+4.73000e-11'
+ mcrdlm3m1_cc_w_0_300_s_1_200 = '-1.00000e-13*ic_cap*ic_cap+-7.50000e-14*ic_cap+4.00000e-11'
+ mcrdlm3m1_cc_w_0_300_s_2_100 = '6.25000e-15*ic_cap*ic_cap+2.17000e-11'
+ mcrdlm3m1_cc_w_0_300_s_3_300 = '3.75000e-14*ic_cap*ic_cap+2.50000e-14*ic_cap+1.18000e-11'
+ mcrdlm3m1_cc_w_0_300_s_9_000 = '2.06250e-14*ic_cap*ic_cap+1.25000e-14*ic_cap+1.31000e-12'
+ mcrdlm3m1_cc_w_2_400_s_0_300 = '-5.93750e-13*ic_cap*ic_cap+-3.75000e-13*ic_cap+1.17000e-10'
+ mcrdlm3m1_cc_w_2_400_s_0_360 = '-5.40625e-13*ic_cap*ic_cap+-4.12500e-13*ic_cap+1.09000e-10'
+ mcrdlm3m1_cc_w_2_400_s_0_450 = '-4.50000e-13*ic_cap*ic_cap+-2.75000e-13*ic_cap+9.80000e-11'
+ mcrdlm3m1_cc_w_2_400_s_0_600 = '-3.00000e-13*ic_cap*ic_cap+-1.75000e-13*ic_cap+8.29000e-11'
+ mcrdlm3m1_cc_w_2_400_s_0_800 = '-1.68750e-13*ic_cap*ic_cap+-1.00000e-13*ic_cap+6.80000e-11'
+ mcrdlm3m1_cc_w_2_400_s_1_000 = '-9.06250e-14*ic_cap*ic_cap+-6.25000e-14*ic_cap+5.70000e-11'
+ mcrdlm3m1_cc_w_2_400_s_1_200 = '-4.68750e-14*ic_cap*ic_cap+-3.75000e-14*ic_cap+4.88000e-11'
+ mcrdlm3m1_cc_w_2_400_s_2_100 = '4.37500e-14*ic_cap*ic_cap+2.50000e-14*ic_cap+2.82000e-11'
+ mcrdlm3m1_cc_w_2_400_s_3_300 = '6.87500e-14*ic_cap*ic_cap+5.00000e-14*ic_cap+1.61000e-11'
+ mcrdlm3m1_cc_w_2_400_s_9_000 = '2.87500e-14*ic_cap*ic_cap+2.25000e-14*ic_cap+2.13000e-12'
+ mcrdlm3m1_cf_w_0_300_s_0_300 = '-2.40625e-14*ic_cap*ic_cap+-1.37500e-14*ic_cap+5.24000e-12'
+ mcrdlm3m1_cf_w_0_300_s_0_360 = '-3.56250e-14*ic_cap*ic_cap+-2.00000e-14*ic_cap+6.25000e-12'
+ mcrdlm3m1_cf_w_0_300_s_0_450 = '-5.15625e-14*ic_cap*ic_cap+-2.87500e-14*ic_cap+7.74000e-12'
+ mcrdlm3m1_cf_w_0_300_s_0_600 = '-7.46875e-14*ic_cap*ic_cap+-4.37500e-14*ic_cap+1.01000e-11'
+ mcrdlm3m1_cf_w_0_300_s_0_800 = '-1.06250e-13*ic_cap*ic_cap+-5.00000e-14*ic_cap+1.30000e-11'
+ mcrdlm3m1_cf_w_0_300_s_1_000 = '-1.37500e-13*ic_cap*ic_cap+-7.50000e-14*ic_cap+1.58000e-11'
+ mcrdlm3m1_cf_w_0_300_s_1_200 = '-1.59375e-13*ic_cap*ic_cap+-8.75000e-14*ic_cap+1.83000e-11'
+ mcrdlm3m1_cf_w_0_300_s_2_100 = '-2.25000e-13*ic_cap*ic_cap+-1.25000e-13*ic_cap+2.77000e-11'
+ mcrdlm3m1_cf_w_0_300_s_3_300 = '-2.65625e-13*ic_cap*ic_cap+-1.62500e-13*ic_cap+3.49000e-11'
+ mcrdlm3m1_cf_w_0_300_s_9_000 = '-2.56250e-13*ic_cap*ic_cap+-1.75000e-13*ic_cap+4.43000e-11'
+ mcrdlm3m1_cf_w_2_400_s_0_300 = '-2.37500e-14*ic_cap*ic_cap+-1.50000e-14*ic_cap+5.26000e-12'
+ mcrdlm3m1_cf_w_2_400_s_0_360 = '-3.56250e-14*ic_cap*ic_cap+-2.00000e-14*ic_cap+6.27000e-12'
+ mcrdlm3m1_cf_w_2_400_s_0_450 = '-5.12500e-14*ic_cap*ic_cap+-3.00000e-14*ic_cap+7.74000e-12'
+ mcrdlm3m1_cf_w_2_400_s_0_600 = '-7.65625e-14*ic_cap*ic_cap+-4.37500e-14*ic_cap+1.01000e-11'
+ mcrdlm3m1_cf_w_2_400_s_0_800 = '-1.09375e-13*ic_cap*ic_cap+-6.25000e-14*ic_cap+1.31000e-11'
+ mcrdlm3m1_cf_w_2_400_s_1_000 = '-1.34375e-13*ic_cap*ic_cap+-8.75000e-14*ic_cap+1.59000e-11'
+ mcrdlm3m1_cf_w_2_400_s_1_200 = '-1.59375e-13*ic_cap*ic_cap+-8.75000e-14*ic_cap+1.85000e-11'
+ mcrdlm3m1_cf_w_2_400_s_2_100 = '-2.28125e-13*ic_cap*ic_cap+-1.37500e-13*ic_cap+2.79000e-11'
+ mcrdlm3m1_cf_w_2_400_s_3_300 = '-2.59375e-13*ic_cap*ic_cap+-1.62500e-13*ic_cap+3.61000e-11'
+ mcrdlm3m1_cf_w_2_400_s_9_000 = '-2.43750e-13*ic_cap*ic_cap+-1.50000e-13*ic_cap+4.82000e-11'
+ mcrdlm3m2_ca_w_0_300_s_0_300 = '-1.28750e-06*ic_cap*ic_cap+-7.00000e-07*ic_cap+8.57000e-05'
+ mcrdlm3m2_ca_w_0_300_s_0_360 = '-1.28750e-06*ic_cap*ic_cap+-7.00000e-07*ic_cap+8.57000e-05'
+ mcrdlm3m2_ca_w_0_300_s_0_450 = '-1.28750e-06*ic_cap*ic_cap+-7.00000e-07*ic_cap+8.57000e-05'
+ mcrdlm3m2_ca_w_0_300_s_0_600 = '-1.28750e-06*ic_cap*ic_cap+-7.00000e-07*ic_cap+8.57000e-05'
+ mcrdlm3m2_ca_w_0_300_s_0_800 = '-1.28750e-06*ic_cap*ic_cap+-7.00000e-07*ic_cap+8.57000e-05'
+ mcrdlm3m2_ca_w_0_300_s_1_000 = '-1.28750e-06*ic_cap*ic_cap+-7.00000e-07*ic_cap+8.57000e-05'
+ mcrdlm3m2_ca_w_0_300_s_1_200 = '-1.28750e-06*ic_cap*ic_cap+-7.00000e-07*ic_cap+8.57000e-05'
+ mcrdlm3m2_ca_w_0_300_s_2_100 = '-1.28750e-06*ic_cap*ic_cap+-7.00000e-07*ic_cap+8.57000e-05'
+ mcrdlm3m2_ca_w_0_300_s_3_300 = '-1.28750e-06*ic_cap*ic_cap+-7.00000e-07*ic_cap+8.57000e-05'
+ mcrdlm3m2_ca_w_0_300_s_9_000 = '-1.28750e-06*ic_cap*ic_cap+-7.00000e-07*ic_cap+8.57000e-05'
+ mcrdlm3m2_ca_w_2_400_s_0_300 = '-1.28750e-06*ic_cap*ic_cap+-7.00000e-07*ic_cap+8.57000e-05'
+ mcrdlm3m2_ca_w_2_400_s_0_360 = '-1.28750e-06*ic_cap*ic_cap+-7.00000e-07*ic_cap+8.57000e-05'
+ mcrdlm3m2_ca_w_2_400_s_0_450 = '-1.28750e-06*ic_cap*ic_cap+-7.00000e-07*ic_cap+8.57000e-05'
+ mcrdlm3m2_ca_w_2_400_s_0_600 = '-1.28750e-06*ic_cap*ic_cap+-7.00000e-07*ic_cap+8.57000e-05'
+ mcrdlm3m2_ca_w_2_400_s_0_800 = '-1.28750e-06*ic_cap*ic_cap+-7.00000e-07*ic_cap+8.57000e-05'
+ mcrdlm3m2_ca_w_2_400_s_1_000 = '-1.28750e-06*ic_cap*ic_cap+-7.00000e-07*ic_cap+8.57000e-05'
+ mcrdlm3m2_ca_w_2_400_s_1_200 = '-1.28750e-06*ic_cap*ic_cap+-7.00000e-07*ic_cap+8.57000e-05'
+ mcrdlm3m2_ca_w_2_400_s_2_100 = '-1.28750e-06*ic_cap*ic_cap+-7.00000e-07*ic_cap+8.57000e-05'
+ mcrdlm3m2_ca_w_2_400_s_3_300 = '-1.28750e-06*ic_cap*ic_cap+-7.00000e-07*ic_cap+8.57000e-05'
+ mcrdlm3m2_ca_w_2_400_s_9_000 = '-1.28750e-06*ic_cap*ic_cap+-7.00000e-07*ic_cap+8.57000e-05'
+ mcrdlm3m2_cc_w_0_300_s_0_300 = '-6.31250e-13*ic_cap*ic_cap+-3.75000e-13*ic_cap+9.31000e-11'
+ mcrdlm3m2_cc_w_0_300_s_0_360 = '-5.68750e-13*ic_cap*ic_cap+-3.25000e-13*ic_cap+8.55000e-11'
+ mcrdlm3m2_cc_w_0_300_s_0_450 = '-4.37500e-13*ic_cap*ic_cap+-2.50000e-13*ic_cap+7.53000e-11'
+ mcrdlm3m2_cc_w_0_300_s_0_600 = '-3.06250e-13*ic_cap*ic_cap+-1.75000e-13*ic_cap+6.18000e-11'
+ mcrdlm3m2_cc_w_0_300_s_0_800 = '-1.87500e-13*ic_cap*ic_cap+-1.25000e-13*ic_cap+4.88000e-11'
+ mcrdlm3m2_cc_w_0_300_s_1_000 = '-1.12500e-13*ic_cap*ic_cap+-1.00000e-13*ic_cap+3.92000e-11'
+ mcrdlm3m2_cc_w_0_300_s_1_200 = '-6.87500e-14*ic_cap*ic_cap+-5.00000e-14*ic_cap+3.23000e-11'
+ mcrdlm3m2_cc_w_0_300_s_3_300 = '2.03125e-14*ic_cap*ic_cap+8.75000e-15*ic_cap+7.64000e-12'
+ mcrdlm3m2_cc_w_0_300_s_9_000 = '6.00000e-15*ic_cap*ic_cap+5.50000e-15*ic_cap+7.65000e-13'
+ mcrdlm3m2_cc_w_2_400_s_0_300 = '-5.68750e-13*ic_cap*ic_cap+-3.25000e-13*ic_cap+1.07000e-10'
+ mcrdlm3m2_cc_w_2_400_s_0_360 = '-5.21875e-13*ic_cap*ic_cap+-3.12500e-13*ic_cap+9.93000e-11'
+ mcrdlm3m2_cc_w_2_400_s_0_450 = '-4.00000e-13*ic_cap*ic_cap+-2.50000e-13*ic_cap+8.82000e-11'
+ mcrdlm3m2_cc_w_2_400_s_0_600 = '-2.56250e-13*ic_cap*ic_cap+-1.50000e-13*ic_cap+7.34000e-11'
+ mcrdlm3m2_cc_w_2_400_s_0_800 = '-1.43750e-13*ic_cap*ic_cap+-1.00000e-13*ic_cap+5.89000e-11'
+ mcrdlm3m2_cc_w_2_400_s_1_000 = '-7.18750e-14*ic_cap*ic_cap+-6.25000e-14*ic_cap+4.84000e-11'
+ mcrdlm3m2_cc_w_2_400_s_1_200 = '-2.81250e-14*ic_cap*ic_cap+-1.25000e-14*ic_cap+4.05000e-11'
+ mcrdlm3m2_cc_w_2_400_s_2_100 = '3.43750e-14*ic_cap*ic_cap+1.25000e-14*ic_cap+2.19000e-11'
+ mcrdlm3m2_cc_w_2_400_s_3_300 = '3.75000e-14*ic_cap*ic_cap+2.50000e-14*ic_cap+1.18000e-11'
+ mcrdlm3m2_cc_w_2_400_s_9_000 = '2.12500e-14*ic_cap*ic_cap+1.50000e-14*ic_cap+1.27000e-12'
+ mcrdlm3m2_cf_w_0_300_s_0_300 = '-9.28125e-14*ic_cap*ic_cap+-4.62500e-14*ic_cap+1.16000e-11'
+ mcrdlm3m2_cf_w_0_300_s_0_360 = '-1.15625e-13*ic_cap*ic_cap+-6.25000e-14*ic_cap+1.36000e-11'
+ mcrdlm3m2_cf_w_0_300_s_0_450 = '-1.53125e-13*ic_cap*ic_cap+-8.75000e-14*ic_cap+1.65000e-11'
+ mcrdlm3m2_cf_w_0_300_s_0_600 = '-2.03125e-13*ic_cap*ic_cap+-1.12500e-13*ic_cap+2.09000e-11'
+ mcrdlm3m2_cf_w_0_300_s_0_800 = '-2.56250e-13*ic_cap*ic_cap+-1.50000e-13*ic_cap+2.59000e-11'
+ mcrdlm3m2_cf_w_0_300_s_1_000 = '-2.93750e-13*ic_cap*ic_cap+-1.75000e-13*ic_cap+3.02000e-11'
+ mcrdlm3m2_cf_w_0_300_s_1_200 = '-3.21875e-13*ic_cap*ic_cap+-1.87500e-13*ic_cap+3.38000e-11'
+ mcrdlm3m2_cf_w_0_300_s_2_100 = '-3.78125e-13*ic_cap*ic_cap+-2.37500e-13*ic_cap+4.52000e-11'
+ mcrdlm3m2_cf_w_0_300_s_3_300 = '-3.90625e-13*ic_cap*ic_cap+-2.37500e-13*ic_cap+5.18000e-11'
+ mcrdlm3m2_cf_w_0_300_s_9_000 = '-3.84375e-13*ic_cap*ic_cap+-2.37500e-13*ic_cap+5.84000e-11'
+ mcrdlm3m2_cf_w_2_400_s_0_300 = '-8.87500e-14*ic_cap*ic_cap+-5.50000e-14*ic_cap+1.16000e-11'
+ mcrdlm3m2_cf_w_2_400_s_0_360 = '-1.21875e-13*ic_cap*ic_cap+-6.25000e-14*ic_cap+1.37000e-11'
+ mcrdlm3m2_cf_w_2_400_s_0_450 = '-1.53125e-13*ic_cap*ic_cap+-8.75000e-14*ic_cap+1.65000e-11'
+ mcrdlm3m2_cf_w_2_400_s_0_600 = '-2.03125e-13*ic_cap*ic_cap+-1.12500e-13*ic_cap+2.09000e-11'
+ mcrdlm3m2_cf_w_2_400_s_0_800 = '-2.53125e-13*ic_cap*ic_cap+-1.37500e-13*ic_cap+2.59000e-11'
+ mcrdlm3m2_cf_w_2_400_s_1_000 = '-2.93750e-13*ic_cap*ic_cap+-1.75000e-13*ic_cap+3.03000e-11'
+ mcrdlm3m2_cf_w_2_400_s_1_200 = '-3.12500e-13*ic_cap*ic_cap+-1.75000e-13*ic_cap+3.39000e-11'
+ mcrdlm3m2_cf_w_2_400_s_2_100 = '-3.68750e-13*ic_cap*ic_cap+-2.25000e-13*ic_cap+4.54000e-11'
+ mcrdlm3m2_cf_w_2_400_s_3_300 = '-3.84375e-13*ic_cap*ic_cap+-2.37500e-13*ic_cap+5.36000e-11'
+ mcrdlm3m2_cf_w_2_400_s_9_000 = '-3.75000e-13*ic_cap*ic_cap+-2.25000e-13*ic_cap+6.34000e-11'
+ mcrdlm3p1_ca_w_0_300_s_0_300 = '-2.12500e-07*ic_cap*ic_cap+-1.25000e-07*ic_cap+1.94000e-05'
+ mcrdlm3p1_ca_w_0_300_s_0_360 = '-2.12500e-07*ic_cap*ic_cap+-1.25000e-07*ic_cap+1.94000e-05'
+ mcrdlm3p1_ca_w_0_300_s_0_450 = '-2.12500e-07*ic_cap*ic_cap+-1.25000e-07*ic_cap+1.94000e-05'
+ mcrdlm3p1_ca_w_0_300_s_0_600 = '-2.12500e-07*ic_cap*ic_cap+-1.25000e-07*ic_cap+1.94000e-05'
+ mcrdlm3p1_ca_w_0_300_s_0_800 = '-2.12500e-07*ic_cap*ic_cap+-1.25000e-07*ic_cap+1.94000e-05'
+ mcrdlm3p1_ca_w_0_300_s_1_000 = '-2.12500e-07*ic_cap*ic_cap+-1.25000e-07*ic_cap+1.94000e-05'
+ mcrdlm3p1_ca_w_0_300_s_1_200 = '-2.12500e-07*ic_cap*ic_cap+-1.25000e-07*ic_cap+1.94000e-05'
+ mcrdlm3p1_ca_w_0_300_s_2_100 = '-2.12500e-07*ic_cap*ic_cap+-1.25000e-07*ic_cap+1.94000e-05'
+ mcrdlm3p1_ca_w_0_300_s_3_300 = '-2.12500e-07*ic_cap*ic_cap+-1.25000e-07*ic_cap+1.94000e-05'
+ mcrdlm3p1_ca_w_0_300_s_9_000 = '-2.12500e-07*ic_cap*ic_cap+-1.25000e-07*ic_cap+1.94000e-05'
+ mcrdlm3p1_ca_w_2_400_s_0_300 = '-2.12500e-07*ic_cap*ic_cap+-1.25000e-07*ic_cap+1.94000e-05'
+ mcrdlm3p1_ca_w_2_400_s_0_360 = '-2.12500e-07*ic_cap*ic_cap+-1.25000e-07*ic_cap+1.94000e-05'
+ mcrdlm3p1_ca_w_2_400_s_0_450 = '-2.12500e-07*ic_cap*ic_cap+-1.25000e-07*ic_cap+1.94000e-05'
+ mcrdlm3p1_ca_w_2_400_s_0_600 = '-2.12500e-07*ic_cap*ic_cap+-1.25000e-07*ic_cap+1.94000e-05'
+ mcrdlm3p1_ca_w_2_400_s_0_800 = '-2.12500e-07*ic_cap*ic_cap+-1.25000e-07*ic_cap+1.94000e-05'
+ mcrdlm3p1_ca_w_2_400_s_1_000 = '-2.12500e-07*ic_cap*ic_cap+-1.25000e-07*ic_cap+1.94000e-05'
+ mcrdlm3p1_ca_w_2_400_s_1_200 = '-2.12500e-07*ic_cap*ic_cap+-1.25000e-07*ic_cap+1.94000e-05'
+ mcrdlm3p1_ca_w_2_400_s_2_100 = '-2.12500e-07*ic_cap*ic_cap+-1.25000e-07*ic_cap+1.94000e-05'
+ mcrdlm3p1_ca_w_2_400_s_3_300 = '-2.12500e-07*ic_cap*ic_cap+-1.25000e-07*ic_cap+1.94000e-05'
+ mcrdlm3p1_ca_w_2_400_s_9_000 = '-2.12500e-07*ic_cap*ic_cap+-1.25000e-07*ic_cap+1.94000e-05'
+ mcrdlm3p1_cc_w_0_300_s_0_300 = '-7.71875e-13*ic_cap*ic_cap+-4.37500e-13*ic_cap+1.05000e-10'
+ mcrdlm3p1_cc_w_0_300_s_0_360 = '-7.03125e-13*ic_cap*ic_cap+-4.37500e-13*ic_cap+9.79000e-11'
+ mcrdlm3p1_cc_w_0_300_s_0_450 = '-5.81250e-13*ic_cap*ic_cap+-3.50000e-13*ic_cap+8.81000e-11'
+ mcrdlm3p1_cc_w_0_300_s_0_600 = '-4.28125e-13*ic_cap*ic_cap+-2.62500e-13*ic_cap+7.51000e-11'
+ mcrdlm3p1_cc_w_0_300_s_0_800 = '-2.81250e-13*ic_cap*ic_cap+-2.00000e-13*ic_cap+6.24000e-11'
+ mcrdlm3p1_cc_w_0_300_s_1_000 = '-1.90625e-13*ic_cap*ic_cap+-1.37500e-13*ic_cap+5.30000e-11'
+ mcrdlm3p1_cc_w_0_300_s_1_200 = '-1.31250e-13*ic_cap*ic_cap+-1.00000e-13*ic_cap+4.59000e-11'
+ mcrdlm3p1_cc_w_0_300_s_2_100 = '-9.37500e-15*ic_cap*ic_cap+-1.25000e-14*ic_cap+2.77000e-11'
+ mcrdlm3p1_cc_w_0_300_s_3_300 = '4.37500e-14*ic_cap*ic_cap+2.50000e-14*ic_cap+1.69000e-11'
+ mcrdlm3p1_cc_w_0_300_s_9_000 = '3.84375e-14*ic_cap*ic_cap+2.62500e-14*ic_cap+2.58000e-12'
+ mcrdlm3p1_cc_w_2_400_s_0_300 = '-6.56250e-13*ic_cap*ic_cap+-3.75000e-13*ic_cap+1.25000e-10'
+ mcrdlm3p1_cc_w_2_400_s_0_360 = '-5.93750e-13*ic_cap*ic_cap+-3.75000e-13*ic_cap+1.17000e-10'
+ mcrdlm3p1_cc_w_2_400_s_0_450 = '-4.75000e-13*ic_cap*ic_cap+-3.25000e-13*ic_cap+1.06000e-10'
+ mcrdlm3p1_cc_w_2_400_s_0_600 = '-3.15625e-13*ic_cap*ic_cap+-1.87500e-13*ic_cap+9.07000e-11'
+ mcrdlm3p1_cc_w_2_400_s_0_800 = '-1.78125e-13*ic_cap*ic_cap+-1.12500e-13*ic_cap+7.57000e-11'
+ mcrdlm3p1_cc_w_2_400_s_1_000 = '-1.03125e-13*ic_cap*ic_cap+-8.75000e-14*ic_cap+6.46000e-11'
+ mcrdlm3p1_cc_w_2_400_s_1_200 = '-4.06250e-14*ic_cap*ic_cap+-3.75000e-14*ic_cap+5.62000e-11'
+ mcrdlm3p1_cc_w_2_400_s_2_100 = '4.68750e-14*ic_cap*ic_cap+3.75000e-14*ic_cap+3.51000e-11'
+ mcrdlm3p1_cc_w_2_400_s_3_300 = '8.43750e-14*ic_cap*ic_cap+6.25000e-14*ic_cap+2.18000e-11'
+ mcrdlm3p1_cc_w_2_400_s_9_000 = '5.81250e-14*ic_cap*ic_cap+4.25000e-14*ic_cap+3.67000e-12'
+ mcrdlm3p1_cf_w_0_300_s_0_300 = '-1.12500e-14*ic_cap*ic_cap+-7.50000e-15*ic_cap+2.87000e-12'
+ mcrdlm3p1_cf_w_0_300_s_0_360 = '-1.68750e-14*ic_cap*ic_cap+-1.00000e-14*ic_cap+3.43000e-12'
+ mcrdlm3p1_cf_w_0_300_s_0_450 = '-2.56250e-14*ic_cap*ic_cap+-1.50000e-14*ic_cap+4.29000e-12'
+ mcrdlm3p1_cf_w_0_300_s_0_600 = '-4.03125e-14*ic_cap*ic_cap+-2.37500e-14*ic_cap+5.70000e-12'
+ mcrdlm3p1_cf_w_0_300_s_0_800 = '-5.87500e-14*ic_cap*ic_cap+-3.75000e-14*ic_cap+7.37000e-12'
+ mcrdlm3p1_cf_w_0_300_s_1_000 = '-7.50000e-14*ic_cap*ic_cap+-4.75000e-14*ic_cap+9.07000e-12'
+ mcrdlm3p1_cf_w_0_300_s_1_200 = '-9.09375e-14*ic_cap*ic_cap+-5.62500e-14*ic_cap+1.07000e-11'
+ mcrdlm3p1_cf_w_0_300_s_2_100 = '-1.46875e-13*ic_cap*ic_cap+-8.75000e-14*ic_cap+1.74000e-11'
+ mcrdlm3p1_cf_w_0_300_s_3_300 = '-1.93750e-13*ic_cap*ic_cap+-1.25000e-13*ic_cap+2.36000e-11'
+ mcrdlm3p1_cf_w_0_300_s_9_000 = '-2.15625e-13*ic_cap*ic_cap+-1.37500e-13*ic_cap+3.52000e-11'
+ mcrdlm3p1_cf_w_2_400_s_0_300 = '-1.21875e-14*ic_cap*ic_cap+-8.75000e-15*ic_cap+2.95000e-12'
+ mcrdlm3p1_cf_w_2_400_s_0_360 = '-1.78125e-14*ic_cap*ic_cap+-1.12500e-14*ic_cap+3.50000e-12'
+ mcrdlm3p1_cf_w_2_400_s_0_450 = '-2.75000e-14*ic_cap*ic_cap+-1.75000e-14*ic_cap+4.35000e-12'
+ mcrdlm3p1_cf_w_2_400_s_0_600 = '-4.06250e-14*ic_cap*ic_cap+-2.50000e-14*ic_cap+5.70000e-12'
+ mcrdlm3p1_cf_w_2_400_s_0_800 = '-5.93750e-14*ic_cap*ic_cap+-3.75000e-14*ic_cap+7.48000e-12'
+ mcrdlm3p1_cf_w_2_400_s_1_000 = '-7.68750e-14*ic_cap*ic_cap+-4.75000e-14*ic_cap+9.21000e-12'
+ mcrdlm3p1_cf_w_2_400_s_1_200 = '-9.50000e-14*ic_cap*ic_cap+-5.75000e-14*ic_cap+1.09000e-11'
+ mcrdlm3p1_cf_w_2_400_s_2_100 = '-1.50000e-13*ic_cap*ic_cap+-1.00000e-13*ic_cap+1.75000e-11'
+ mcrdlm3p1_cf_w_2_400_s_3_300 = '-2.00000e-13*ic_cap*ic_cap+-1.25000e-13*ic_cap+2.45000e-11'
+ mcrdlm3p1_cf_w_2_400_s_9_000 = '-2.15625e-13*ic_cap*ic_cap+-1.37500e-13*ic_cap+3.86000e-11'
+ mcrdlm4_ca_w_10_000_s_10_000 = '-3.90625e-08*ic_cap*ic_cap+-2.37500e-08*ic_cap+4.00000e-06'
+ mcrdlm4_ca_w_10_000_s_12_000 = '-3.90625e-08*ic_cap*ic_cap+-2.37500e-08*ic_cap+4.00000e-06'
+ mcrdlm4_ca_w_10_000_s_30_000 = '-3.90625e-08*ic_cap*ic_cap+-2.37500e-08*ic_cap+4.00000e-06'
+ mcrdlm4_ca_w_10_000_s_5_000 = '-3.90625e-08*ic_cap*ic_cap+-2.37500e-08*ic_cap+4.00000e-06'
+ mcrdlm4_ca_w_10_000_s_8_000 = '-3.90625e-08*ic_cap*ic_cap+-2.37500e-08*ic_cap+4.00000e-06'
+ mcrdlm4_ca_w_40_000_s_10_000 = '-3.90625e-08*ic_cap*ic_cap+-2.37500e-08*ic_cap+4.00000e-06'
+ mcrdlm4_ca_w_40_000_s_12_000 = '-3.90625e-08*ic_cap*ic_cap+-2.37500e-08*ic_cap+4.00000e-06'
+ mcrdlm4_ca_w_40_000_s_30_000 = '-3.90625e-08*ic_cap*ic_cap+-2.37500e-08*ic_cap+4.00000e-06'
+ mcrdlm4_ca_w_40_000_s_5_000 = '-3.90625e-08*ic_cap*ic_cap+-2.37500e-08*ic_cap+4.00000e-06'
+ mcrdlm4_ca_w_40_000_s_8_000 = '-3.90625e-08*ic_cap*ic_cap+-2.37500e-08*ic_cap+4.00000e-06'
+ mcrdlm4_cc_w_10_000_s_10_000 = '-2.34375e-13*ic_cap*ic_cap+-1.37500e-13*ic_cap+2.85000e-11'
+ mcrdlm4_cc_w_10_000_s_12_000 = '-1.81250e-13*ic_cap*ic_cap+-1.25000e-13*ic_cap+2.45000e-11'
+ mcrdlm4_cc_w_10_000_s_30_000 = '-6.34375e-14*ic_cap*ic_cap+-3.87500e-14*ic_cap+9.97000e-12'
+ mcrdlm4_cc_w_10_000_s_5_000 = '-5.43750e-13*ic_cap*ic_cap+-3.25000e-13*ic_cap+4.78000e-11'
+ mcrdlm4_cc_w_10_000_s_8_000 = '-3.00000e-13*ic_cap*ic_cap+-2.00000e-13*ic_cap+3.38000e-11'
+ mcrdlm4_cc_w_40_000_s_10_000 = '-2.34375e-13*ic_cap*ic_cap+-1.62500e-13*ic_cap+3.83000e-11'
+ mcrdlm4_cc_w_40_000_s_12_000 = '-1.90625e-13*ic_cap*ic_cap+-1.12500e-13*ic_cap+3.40000e-11'
+ mcrdlm4_cc_w_40_000_s_30_000 = '-5.93750e-14*ic_cap*ic_cap+-3.75000e-14*ic_cap+1.70000e-11'
+ mcrdlm4_cc_w_40_000_s_5_000 = '-5.50000e-13*ic_cap*ic_cap+-3.25000e-13*ic_cap+5.90000e-11'
+ mcrdlm4_cc_w_40_000_s_8_000 = '-3.03125e-13*ic_cap*ic_cap+-1.87500e-13*ic_cap+4.41000e-11'
+ mcrdlm4_cf_w_10_000_s_10_000 = '-7.18750e-14*ic_cap*ic_cap+-3.75000e-14*ic_cap+1.54000e-11'
+ mcrdlm4_cf_w_10_000_s_12_000 = '-8.75000e-14*ic_cap*ic_cap+-5.00000e-14*ic_cap+1.75000e-11'
+ mcrdlm4_cf_w_10_000_s_30_000 = '-1.62500e-13*ic_cap*ic_cap+-1.00000e-13*ic_cap+2.84000e-11'
+ mcrdlm4_cf_w_10_000_s_5_000 = '-8.75000e-15*ic_cap*ic_cap+-5.00000e-15*ic_cap+8.79000e-12'
+ mcrdlm4_cf_w_10_000_s_8_000 = '-5.00000e-14*ic_cap*ic_cap+-2.50000e-14*ic_cap+1.30000e-11'
+ mcrdlm4_cf_w_40_000_s_10_000 = '-6.56250e-14*ic_cap*ic_cap+-3.75000e-14*ic_cap+1.53000e-11'
+ mcrdlm4_cf_w_40_000_s_12_000 = '-8.75000e-14*ic_cap*ic_cap+-5.00000e-14*ic_cap+1.75000e-11'
+ mcrdlm4_cf_w_40_000_s_30_000 = '-1.62500e-13*ic_cap*ic_cap+-1.00000e-13*ic_cap+2.94000e-11'
+ mcrdlm4_cf_w_40_000_s_5_000 = '-9.68750e-15*ic_cap*ic_cap+-1.25000e-15*ic_cap+8.71000e-12'
+ mcrdlm4_cf_w_40_000_s_8_000 = '-5.00000e-14*ic_cap*ic_cap+-2.50000e-14*ic_cap+1.29000e-11'
+ mcrdlm4d_ca_w_0_300_s_0_300 = '-1.18750e-07*ic_cap*ic_cap+-7.50000e-08*ic_cap+1.34000e-05'
+ mcrdlm4d_ca_w_0_300_s_0_360 = '-1.18750e-07*ic_cap*ic_cap+-7.50000e-08*ic_cap+1.34000e-05'
+ mcrdlm4d_ca_w_0_300_s_0_450 = '-1.18750e-07*ic_cap*ic_cap+-7.50000e-08*ic_cap+1.34000e-05'
+ mcrdlm4d_ca_w_0_300_s_0_600 = '-1.18750e-07*ic_cap*ic_cap+-7.50000e-08*ic_cap+1.34000e-05'
+ mcrdlm4d_ca_w_0_300_s_0_800 = '-1.18750e-07*ic_cap*ic_cap+-7.50000e-08*ic_cap+1.34000e-05'
+ mcrdlm4d_ca_w_0_300_s_1_000 = '-1.18750e-07*ic_cap*ic_cap+-7.50000e-08*ic_cap+1.34000e-05'
+ mcrdlm4d_ca_w_0_300_s_1_200 = '-1.18750e-07*ic_cap*ic_cap+-7.50000e-08*ic_cap+1.34000e-05'
+ mcrdlm4d_ca_w_0_300_s_2_100 = '-1.18750e-07*ic_cap*ic_cap+-7.50000e-08*ic_cap+1.34000e-05'
+ mcrdlm4d_ca_w_0_300_s_3_300 = '-1.18750e-07*ic_cap*ic_cap+-7.50000e-08*ic_cap+1.34000e-05'
+ mcrdlm4d_ca_w_0_300_s_9_000 = '-1.18750e-07*ic_cap*ic_cap+-7.50000e-08*ic_cap+1.34000e-05'
+ mcrdlm4d_ca_w_2_400_s_0_300 = '-1.18750e-07*ic_cap*ic_cap+-7.50000e-08*ic_cap+1.34000e-05'
+ mcrdlm4d_ca_w_2_400_s_0_360 = '-1.18750e-07*ic_cap*ic_cap+-7.50000e-08*ic_cap+1.34000e-05'
+ mcrdlm4d_ca_w_2_400_s_0_450 = '-1.18750e-07*ic_cap*ic_cap+-7.50000e-08*ic_cap+1.34000e-05'
+ mcrdlm4d_ca_w_2_400_s_0_600 = '-1.18750e-07*ic_cap*ic_cap+-7.50000e-08*ic_cap+1.34000e-05'
+ mcrdlm4d_ca_w_2_400_s_0_800 = '-1.18750e-07*ic_cap*ic_cap+-7.50000e-08*ic_cap+1.34000e-05'
+ mcrdlm4d_ca_w_2_400_s_1_000 = '-1.18750e-07*ic_cap*ic_cap+-7.50000e-08*ic_cap+1.34000e-05'
+ mcrdlm4d_ca_w_2_400_s_1_200 = '-1.18750e-07*ic_cap*ic_cap+-7.50000e-08*ic_cap+1.34000e-05'
+ mcrdlm4d_ca_w_2_400_s_2_100 = '-1.18750e-07*ic_cap*ic_cap+-7.50000e-08*ic_cap+1.34000e-05'
+ mcrdlm4d_ca_w_2_400_s_3_300 = '-1.18750e-07*ic_cap*ic_cap+-7.50000e-08*ic_cap+1.34000e-05'
+ mcrdlm4d_ca_w_2_400_s_9_000 = '-1.18750e-07*ic_cap*ic_cap+-7.50000e-08*ic_cap+1.34000e-05'
+ mcrdlm4d_cc_w_0_300_s_0_300 = '-8.15625e-13*ic_cap*ic_cap+-4.37500e-13*ic_cap+1.07000e-10'
+ mcrdlm4d_cc_w_0_300_s_0_360 = '-7.25000e-13*ic_cap*ic_cap+-4.00000e-13*ic_cap+9.98000e-11'
+ mcrdlm4d_cc_w_0_300_s_0_450 = '-6.50000e-13*ic_cap*ic_cap+-4.00000e-13*ic_cap+9.07000e-11'
+ mcrdlm4d_cc_w_0_300_s_0_600 = '-4.78125e-13*ic_cap*ic_cap+-2.87500e-13*ic_cap+7.78000e-11'
+ mcrdlm4d_cc_w_0_300_s_0_800 = '-3.53125e-13*ic_cap*ic_cap+-2.37500e-13*ic_cap+6.58000e-11'
+ mcrdlm4d_cc_w_0_300_s_1_000 = '-2.68750e-13*ic_cap*ic_cap+-1.75000e-13*ic_cap+5.66000e-11'
+ mcrdlm4d_cc_w_0_300_s_1_200 = '-2.06250e-13*ic_cap*ic_cap+-1.50000e-13*ic_cap+4.97000e-11'
+ mcrdlm4d_cc_w_0_300_s_2_100 = '-7.50000e-14*ic_cap*ic_cap+-5.00000e-14*ic_cap+3.19000e-11'
+ mcrdlm4d_cc_w_0_300_s_3_300 = '-3.12500e-15*ic_cap*ic_cap+-1.25000e-14*ic_cap+2.07000e-11'
+ mcrdlm4d_cc_w_0_300_s_9_000 = '3.75000e-14*ic_cap*ic_cap+2.25000e-14*ic_cap+3.82000e-12'
+ mcrdlm4d_cc_w_2_400_s_0_300 = '-7.50000e-13*ic_cap*ic_cap+-5.00000e-13*ic_cap+1.31000e-10'
+ mcrdlm4d_cc_w_2_400_s_0_360 = '-7.18750e-13*ic_cap*ic_cap+-3.75000e-13*ic_cap+1.23000e-10'
+ mcrdlm4d_cc_w_2_400_s_0_450 = '-5.93750e-13*ic_cap*ic_cap+-3.75000e-13*ic_cap+1.12000e-10'
+ mcrdlm4d_cc_w_2_400_s_0_600 = '-4.21875e-13*ic_cap*ic_cap+-2.62500e-13*ic_cap+9.68000e-11'
+ mcrdlm4d_cc_w_2_400_s_0_800 = '-2.71875e-13*ic_cap*ic_cap+-1.62500e-13*ic_cap+8.15000e-11'
+ mcrdlm4d_cc_w_2_400_s_1_000 = '-2.03125e-13*ic_cap*ic_cap+-1.62500e-13*ic_cap+7.05000e-11'
+ mcrdlm4d_cc_w_2_400_s_1_200 = '-1.40625e-13*ic_cap*ic_cap+-1.12500e-13*ic_cap+6.20000e-11'
+ mcrdlm4d_cc_w_2_400_s_2_100 = '-1.25000e-14*ic_cap*ic_cap+-2.50000e-14*ic_cap+4.01000e-11'
+ mcrdlm4d_cc_w_2_400_s_3_300 = '4.68750e-14*ic_cap*ic_cap+1.25000e-14*ic_cap+2.59000e-11'
+ mcrdlm4d_cc_w_2_400_s_9_000 = '6.18750e-14*ic_cap*ic_cap+4.50000e-14*ic_cap+4.98000e-12'
+ mcrdlm4d_cf_w_0_300_s_0_300 = '-2.50000e-15*ic_cap*ic_cap+-2.50000e-15*ic_cap+1.98000e-12'
+ mcrdlm4d_cf_w_0_300_s_0_360 = '-5.93750e-15*ic_cap*ic_cap+-3.75000e-15*ic_cap+2.38000e-12'
+ mcrdlm4d_cf_w_0_300_s_0_450 = '-1.12500e-14*ic_cap*ic_cap+-7.50000e-15*ic_cap+3.00000e-12'
+ mcrdlm4d_cf_w_0_300_s_0_600 = '-2.06250e-14*ic_cap*ic_cap+-1.25000e-14*ic_cap+4.02000e-12'
+ mcrdlm4d_cf_w_0_300_s_0_800 = '-3.09375e-14*ic_cap*ic_cap+-1.87500e-14*ic_cap+5.19000e-12'
+ mcrdlm4d_cf_w_0_300_s_1_000 = '-4.15625e-14*ic_cap*ic_cap+-2.62500e-14*ic_cap+6.42000e-12'
+ mcrdlm4d_cf_w_0_300_s_1_200 = '-5.15625e-14*ic_cap*ic_cap+-3.12500e-14*ic_cap+7.63000e-12'
+ mcrdlm4d_cf_w_0_300_s_2_100 = '-9.06250e-14*ic_cap*ic_cap+-6.25000e-14*ic_cap+1.28000e-11'
+ mcrdlm4d_cf_w_0_300_s_3_300 = '-1.34375e-13*ic_cap*ic_cap+-8.75000e-14*ic_cap+1.80000e-11'
+ mcrdlm4d_cf_w_0_300_s_9_000 = '-1.78125e-13*ic_cap*ic_cap+-1.12500e-13*ic_cap+3.02000e-11'
+ mcrdlm4d_cf_w_2_400_s_0_300 = '-2.81250e-15*ic_cap*ic_cap+-1.25000e-15*ic_cap+2.01000e-12'
+ mcrdlm4d_cf_w_2_400_s_0_360 = '-6.56250e-15*ic_cap*ic_cap+-3.75000e-15*ic_cap+2.41000e-12'
+ mcrdlm4d_cf_w_2_400_s_0_450 = '-1.18750e-14*ic_cap*ic_cap+-7.50000e-15*ic_cap+3.00000e-12'
+ mcrdlm4d_cf_w_2_400_s_0_600 = '-2.03125e-14*ic_cap*ic_cap+-1.12500e-14*ic_cap+3.97000e-12'
+ mcrdlm4d_cf_w_2_400_s_0_800 = '-3.09375e-14*ic_cap*ic_cap+-1.87500e-14*ic_cap+5.24000e-12'
+ mcrdlm4d_cf_w_2_400_s_1_000 = '-4.18750e-14*ic_cap*ic_cap+-2.50000e-14*ic_cap+6.49000e-12'
+ mcrdlm4d_cf_w_2_400_s_1_200 = '-5.18750e-14*ic_cap*ic_cap+-3.25000e-14*ic_cap+7.71000e-12'
+ mcrdlm4d_cf_w_2_400_s_2_100 = '-9.06250e-14*ic_cap*ic_cap+-6.25000e-14*ic_cap+1.28000e-11'
+ mcrdlm4d_cf_w_2_400_s_3_300 = '-1.34375e-13*ic_cap*ic_cap+-8.75000e-14*ic_cap+1.86000e-11'
+ mcrdlm4d_cf_w_2_400_s_9_000 = '-1.81250e-13*ic_cap*ic_cap+-1.25000e-13*ic_cap+3.31000e-11'
+ mcrdlm4f_ca_w_0_300_s_0_300 = '-1.15625e-07*ic_cap*ic_cap+-6.25000e-08*ic_cap+1.27000e-05'
+ mcrdlm4f_ca_w_0_300_s_0_360 = '-1.15625e-07*ic_cap*ic_cap+-6.25000e-08*ic_cap+1.27000e-05'
+ mcrdlm4f_ca_w_0_300_s_0_450 = '-1.15625e-07*ic_cap*ic_cap+-6.25000e-08*ic_cap+1.27000e-05'
+ mcrdlm4f_ca_w_0_300_s_0_600 = '-1.15625e-07*ic_cap*ic_cap+-6.25000e-08*ic_cap+1.27000e-05'
+ mcrdlm4f_ca_w_0_300_s_0_800 = '-1.15625e-07*ic_cap*ic_cap+-6.25000e-08*ic_cap+1.27000e-05'
+ mcrdlm4f_ca_w_0_300_s_1_000 = '-1.15625e-07*ic_cap*ic_cap+-6.25000e-08*ic_cap+1.27000e-05'
+ mcrdlm4f_ca_w_0_300_s_1_200 = '-1.15625e-07*ic_cap*ic_cap+-6.25000e-08*ic_cap+1.27000e-05'
+ mcrdlm4f_ca_w_0_300_s_2_100 = '-1.15625e-07*ic_cap*ic_cap+-6.25000e-08*ic_cap+1.27000e-05'
+ mcrdlm4f_ca_w_0_300_s_3_300 = '-1.15625e-07*ic_cap*ic_cap+-6.25000e-08*ic_cap+1.27000e-05'
+ mcrdlm4f_ca_w_0_300_s_9_000 = '-1.15625e-07*ic_cap*ic_cap+-6.25000e-08*ic_cap+1.27000e-05'
+ mcrdlm4f_ca_w_2_400_s_0_300 = '-1.15625e-07*ic_cap*ic_cap+-6.25000e-08*ic_cap+1.27000e-05'
+ mcrdlm4f_ca_w_2_400_s_0_360 = '-1.15625e-07*ic_cap*ic_cap+-6.25000e-08*ic_cap+1.27000e-05'
+ mcrdlm4f_ca_w_2_400_s_0_450 = '-1.15625e-07*ic_cap*ic_cap+-6.25000e-08*ic_cap+1.27000e-05'
+ mcrdlm4f_ca_w_2_400_s_0_600 = '-1.15625e-07*ic_cap*ic_cap+-6.25000e-08*ic_cap+1.27000e-05'
+ mcrdlm4f_ca_w_2_400_s_0_800 = '-1.15625e-07*ic_cap*ic_cap+-6.25000e-08*ic_cap+1.27000e-05'
+ mcrdlm4f_ca_w_2_400_s_1_000 = '-1.15625e-07*ic_cap*ic_cap+-6.25000e-08*ic_cap+1.27000e-05'
+ mcrdlm4f_ca_w_2_400_s_1_200 = '-1.15625e-07*ic_cap*ic_cap+-6.25000e-08*ic_cap+1.27000e-05'
+ mcrdlm4f_ca_w_2_400_s_2_100 = '-1.15625e-07*ic_cap*ic_cap+-6.25000e-08*ic_cap+1.27000e-05'
+ mcrdlm4f_ca_w_2_400_s_3_300 = '-1.15625e-07*ic_cap*ic_cap+-6.25000e-08*ic_cap+1.27000e-05'
+ mcrdlm4f_ca_w_2_400_s_9_000 = '-1.15625e-07*ic_cap*ic_cap+-6.25000e-08*ic_cap+1.27000e-05'
+ mcrdlm4f_cc_w_0_300_s_0_300 = '-8.03125e-13*ic_cap*ic_cap+-4.37500e-13*ic_cap+1.07000e-10'
+ mcrdlm4f_cc_w_0_300_s_0_360 = '-7.21875e-13*ic_cap*ic_cap+-4.12500e-13*ic_cap+1.00000e-10'
+ mcrdlm4f_cc_w_0_300_s_0_450 = '-6.50000e-13*ic_cap*ic_cap+-4.00000e-13*ic_cap+9.09000e-11'
+ mcrdlm4f_cc_w_0_300_s_0_600 = '-4.75000e-13*ic_cap*ic_cap+-3.00000e-13*ic_cap+7.80000e-11'
+ mcrdlm4f_cc_w_0_300_s_0_800 = '-3.56250e-13*ic_cap*ic_cap+-2.50000e-13*ic_cap+6.61000e-11'
+ mcrdlm4f_cc_w_0_300_s_1_000 = '-2.68750e-13*ic_cap*ic_cap+-1.75000e-13*ic_cap+5.70000e-11'
+ mcrdlm4f_cc_w_0_300_s_1_200 = '-2.03125e-13*ic_cap*ic_cap+-1.62500e-13*ic_cap+5.01000e-11'
+ mcrdlm4f_cc_w_0_300_s_2_100 = '-7.81250e-14*ic_cap*ic_cap+-6.25000e-14*ic_cap+3.25000e-11'
+ mcrdlm4f_cc_w_0_300_s_3_300 = '-6.25000e-15*ic_cap*ic_cap+2.13000e-11'
+ mcrdlm4f_cc_w_0_300_s_9_000 = '4.25000e-14*ic_cap*ic_cap+2.75000e-14*ic_cap+4.11000e-12'
+ mcrdlm4f_cc_w_2_400_s_0_300 = '-7.81250e-13*ic_cap*ic_cap+-3.75000e-13*ic_cap+1.32000e-10'
+ mcrdlm4f_cc_w_2_400_s_0_360 = '-7.18750e-13*ic_cap*ic_cap+-3.75000e-13*ic_cap+1.24000e-10'
+ mcrdlm4f_cc_w_2_400_s_0_450 = '-5.93750e-13*ic_cap*ic_cap+-3.75000e-13*ic_cap+1.13000e-10'
+ mcrdlm4f_cc_w_2_400_s_0_600 = '-4.18750e-13*ic_cap*ic_cap+-2.50000e-13*ic_cap+9.74000e-11'
+ mcrdlm4f_cc_w_2_400_s_0_800 = '-2.81250e-13*ic_cap*ic_cap+-1.75000e-13*ic_cap+8.23000e-11'
+ mcrdlm4f_cc_w_2_400_s_1_000 = '-1.96875e-13*ic_cap*ic_cap+-1.62500e-13*ic_cap+7.12000e-11'
+ mcrdlm4f_cc_w_2_400_s_1_200 = '-1.37500e-13*ic_cap*ic_cap+-1.25000e-13*ic_cap+6.27000e-11'
+ mcrdlm4f_cc_w_2_400_s_2_100 = '-1.25000e-14*ic_cap*ic_cap+-2.50000e-14*ic_cap+4.09000e-11'
+ mcrdlm4f_cc_w_2_400_s_3_300 = '5.00000e-14*ic_cap*ic_cap+2.50000e-14*ic_cap+2.67000e-11'
+ mcrdlm4f_cc_w_2_400_s_9_000 = '6.93750e-14*ic_cap*ic_cap+4.50000e-14*ic_cap+5.36000e-12'
+ mcrdlm4f_cf_w_0_300_s_0_300 = '-3.75000e-15*ic_cap*ic_cap+-2.50000e-15*ic_cap+1.88000e-12'
+ mcrdlm4f_cf_w_0_300_s_0_360 = '-6.56250e-15*ic_cap*ic_cap+-3.75000e-15*ic_cap+2.25000e-12'
+ mcrdlm4f_cf_w_0_300_s_0_450 = '-1.18750e-14*ic_cap*ic_cap+-7.50000e-15*ic_cap+2.84000e-12'
+ mcrdlm4f_cf_w_0_300_s_0_600 = '-2.06250e-14*ic_cap*ic_cap+-1.25000e-14*ic_cap+3.80000e-12'
+ mcrdlm4f_cf_w_0_300_s_0_800 = '-3.06250e-14*ic_cap*ic_cap+-2.00000e-14*ic_cap+4.91000e-12'
+ mcrdlm4f_cf_w_0_300_s_1_000 = '-4.18750e-14*ic_cap*ic_cap+-2.50000e-14*ic_cap+6.09000e-12'
+ mcrdlm4f_cf_w_0_300_s_1_200 = '-5.15625e-14*ic_cap*ic_cap+-3.37500e-14*ic_cap+7.24000e-12'
+ mcrdlm4f_cf_w_0_300_s_2_100 = '-9.06250e-14*ic_cap*ic_cap+-6.25000e-14*ic_cap+1.22000e-11'
+ mcrdlm4f_cf_w_0_300_s_3_300 = '-1.34375e-13*ic_cap*ic_cap+-8.75000e-14*ic_cap+1.72000e-11'
+ mcrdlm4f_cf_w_0_300_s_9_000 = '-1.81250e-13*ic_cap*ic_cap+-1.25000e-13*ic_cap+2.94000e-11'
+ mcrdlm4f_cf_w_2_400_s_0_300 = '-3.12500e-15*ic_cap*ic_cap+-2.50000e-15*ic_cap+1.90000e-12'
+ mcrdlm4f_cf_w_2_400_s_0_360 = '-6.87500e-15*ic_cap*ic_cap+-5.00000e-15*ic_cap+2.28000e-12'
+ mcrdlm4f_cf_w_2_400_s_0_450 = '-1.18750e-14*ic_cap*ic_cap+-7.50000e-15*ic_cap+2.83000e-12'
+ mcrdlm4f_cf_w_2_400_s_0_600 = '-2.00000e-14*ic_cap*ic_cap+-1.25000e-14*ic_cap+3.75000e-12'
+ mcrdlm4f_cf_w_2_400_s_0_800 = '-3.09375e-14*ic_cap*ic_cap+-1.87500e-14*ic_cap+4.96000e-12'
+ mcrdlm4f_cf_w_2_400_s_1_000 = '-4.09375e-14*ic_cap*ic_cap+-2.62500e-14*ic_cap+6.14000e-12'
+ mcrdlm4f_cf_w_2_400_s_1_200 = '-5.18750e-14*ic_cap*ic_cap+-3.25000e-14*ic_cap+7.31000e-12'
+ mcrdlm4f_cf_w_2_400_s_2_100 = '-9.37500e-14*ic_cap*ic_cap+-5.00000e-14*ic_cap+1.22000e-11'
+ mcrdlm4f_cf_w_2_400_s_3_300 = '-1.34375e-13*ic_cap*ic_cap+-8.75000e-14*ic_cap+1.78000e-11'
+ mcrdlm4f_cf_w_2_400_s_9_000 = '-1.87500e-13*ic_cap*ic_cap+-1.25000e-13*ic_cap+3.22000e-11'
+ mcrdlm4l1_ca_w_0_300_s_0_300 = '-1.34375e-07*ic_cap*ic_cap+-8.75000e-08*ic_cap+1.57000e-05'
+ mcrdlm4l1_ca_w_0_300_s_0_360 = '-1.34375e-07*ic_cap*ic_cap+-8.75000e-08*ic_cap+1.57000e-05'
+ mcrdlm4l1_ca_w_0_300_s_0_450 = '-1.34375e-07*ic_cap*ic_cap+-8.75000e-08*ic_cap+1.57000e-05'
+ mcrdlm4l1_ca_w_0_300_s_0_600 = '-1.34375e-07*ic_cap*ic_cap+-8.75000e-08*ic_cap+1.57000e-05'
+ mcrdlm4l1_ca_w_0_300_s_0_800 = '-1.34375e-07*ic_cap*ic_cap+-8.75000e-08*ic_cap+1.57000e-05'
+ mcrdlm4l1_ca_w_0_300_s_1_000 = '-1.34375e-07*ic_cap*ic_cap+-8.75000e-08*ic_cap+1.57000e-05'
+ mcrdlm4l1_ca_w_0_300_s_1_200 = '-1.34375e-07*ic_cap*ic_cap+-8.75000e-08*ic_cap+1.57000e-05'
+ mcrdlm4l1_ca_w_0_300_s_2_100 = '-1.34375e-07*ic_cap*ic_cap+-8.75000e-08*ic_cap+1.57000e-05'
+ mcrdlm4l1_ca_w_0_300_s_3_300 = '-1.34375e-07*ic_cap*ic_cap+-8.75000e-08*ic_cap+1.57000e-05'
+ mcrdlm4l1_ca_w_0_300_s_9_000 = '-1.34375e-07*ic_cap*ic_cap+-8.75000e-08*ic_cap+1.57000e-05'
+ mcrdlm4l1_ca_w_2_400_s_0_300 = '-1.34375e-07*ic_cap*ic_cap+-8.75000e-08*ic_cap+1.57000e-05'
+ mcrdlm4l1_ca_w_2_400_s_0_360 = '-1.34375e-07*ic_cap*ic_cap+-8.75000e-08*ic_cap+1.57000e-05'
+ mcrdlm4l1_ca_w_2_400_s_0_450 = '-1.34375e-07*ic_cap*ic_cap+-8.75000e-08*ic_cap+1.57000e-05'
+ mcrdlm4l1_ca_w_2_400_s_0_600 = '-1.34375e-07*ic_cap*ic_cap+-8.75000e-08*ic_cap+1.57000e-05'
+ mcrdlm4l1_ca_w_2_400_s_0_800 = '-1.34375e-07*ic_cap*ic_cap+-8.75000e-08*ic_cap+1.57000e-05'
+ mcrdlm4l1_ca_w_2_400_s_1_000 = '-1.34375e-07*ic_cap*ic_cap+-8.75000e-08*ic_cap+1.57000e-05'
+ mcrdlm4l1_ca_w_2_400_s_1_200 = '-1.34375e-07*ic_cap*ic_cap+-8.75000e-08*ic_cap+1.57000e-05'
+ mcrdlm4l1_ca_w_2_400_s_2_100 = '-1.34375e-07*ic_cap*ic_cap+-8.75000e-08*ic_cap+1.57000e-05'
+ mcrdlm4l1_ca_w_2_400_s_3_300 = '-1.34375e-07*ic_cap*ic_cap+-8.75000e-08*ic_cap+1.57000e-05'
+ mcrdlm4l1_ca_w_2_400_s_9_000 = '-1.34375e-07*ic_cap*ic_cap+-8.75000e-08*ic_cap+1.57000e-05'
+ mcrdlm4l1_cc_w_0_300_s_0_300 = '-7.84375e-13*ic_cap*ic_cap+-4.37500e-13*ic_cap+1.06000e-10'
+ mcrdlm4l1_cc_w_0_300_s_0_360 = '-7.21875e-13*ic_cap*ic_cap+-4.12500e-13*ic_cap+9.92000e-11'
+ mcrdlm4l1_cc_w_0_300_s_0_450 = '-6.28125e-13*ic_cap*ic_cap+-3.87500e-13*ic_cap+8.98000e-11'
+ mcrdlm4l1_cc_w_0_300_s_0_600 = '-4.78125e-13*ic_cap*ic_cap+-2.87500e-13*ic_cap+7.71000e-11'
+ mcrdlm4l1_cc_w_0_300_s_0_800 = '-3.34375e-13*ic_cap*ic_cap+-2.12500e-13*ic_cap+6.47000e-11'
+ mcrdlm4l1_cc_w_0_300_s_1_000 = '-2.62500e-13*ic_cap*ic_cap+-1.75000e-13*ic_cap+5.55000e-11'
+ mcrdlm4l1_cc_w_0_300_s_1_200 = '-2.06250e-13*ic_cap*ic_cap+-1.25000e-13*ic_cap+4.86000e-11'
+ mcrdlm4l1_cc_w_0_300_s_2_100 = '-6.56250e-14*ic_cap*ic_cap+-6.25000e-14*ic_cap+3.04000e-11'
+ mcrdlm4l1_cc_w_0_300_s_9_000 = '3.31250e-14*ic_cap*ic_cap+2.00000e-14*ic_cap+3.08000e-12'
+ mcrdlm4l1_cc_w_2_400_s_0_300 = '-7.50000e-13*ic_cap*ic_cap+-5.00000e-13*ic_cap+1.29000e-10'
+ mcrdlm4l1_cc_w_2_400_s_0_360 = '-6.56250e-13*ic_cap*ic_cap+-3.75000e-13*ic_cap+1.21000e-10'
+ mcrdlm4l1_cc_w_2_400_s_0_450 = '-5.78125e-13*ic_cap*ic_cap+-3.12500e-13*ic_cap+1.10000e-10'
+ mcrdlm4l1_cc_w_2_400_s_0_600 = '-4.00000e-13*ic_cap*ic_cap+-2.50000e-13*ic_cap+9.46000e-11'
+ mcrdlm4l1_cc_w_2_400_s_0_800 = '-2.71875e-13*ic_cap*ic_cap+-1.62500e-13*ic_cap+7.96000e-11'
+ mcrdlm4l1_cc_w_2_400_s_1_000 = '-1.90625e-13*ic_cap*ic_cap+-1.37500e-13*ic_cap+6.84000e-11'
+ mcrdlm4l1_cc_w_2_400_s_1_200 = '-1.25000e-13*ic_cap*ic_cap+-1.00000e-13*ic_cap+5.98000e-11'
+ mcrdlm4l1_cc_w_2_400_s_2_100 = '-9.37500e-15*ic_cap*ic_cap+-1.25000e-14*ic_cap+3.80000e-11'
+ mcrdlm4l1_cc_w_2_400_s_3_300 = '5.00000e-14*ic_cap*ic_cap+2.50000e-14*ic_cap+2.39000e-11'
+ mcrdlm4l1_cc_w_2_400_s_9_000 = '5.34375e-14*ic_cap*ic_cap+3.87500e-14*ic_cap+4.05000e-12'
+ mcrdlm4l1_cf_w_0_300_s_0_300 = '-3.12500e-15*ic_cap*ic_cap+-2.50000e-15*ic_cap+2.32000e-12'
+ mcrdlm4l1_cf_w_0_300_s_0_360 = '-6.87500e-15*ic_cap*ic_cap+-5.00000e-15*ic_cap+2.78000e-12'
+ mcrdlm4l1_cf_w_0_300_s_0_450 = '-1.25000e-14*ic_cap*ic_cap+-7.50000e-15*ic_cap+3.49000e-12'
+ mcrdlm4l1_cf_w_0_300_s_0_600 = '-2.31250e-14*ic_cap*ic_cap+-1.50000e-14*ic_cap+4.67000e-12'
+ mcrdlm4l1_cf_w_0_300_s_0_800 = '-3.53125e-14*ic_cap*ic_cap+-2.12500e-14*ic_cap+6.04000e-12'
+ mcrdlm4l1_cf_w_0_300_s_1_000 = '-4.81250e-14*ic_cap*ic_cap+-3.00000e-14*ic_cap+7.46000e-12'
+ mcrdlm4l1_cf_w_0_300_s_1_200 = '-6.03125e-14*ic_cap*ic_cap+-3.62500e-14*ic_cap+8.84000e-12'
+ mcrdlm4l1_cf_w_0_300_s_2_100 = '-1.03125e-13*ic_cap*ic_cap+-6.25000e-14*ic_cap+1.46000e-11'
+ mcrdlm4l1_cf_w_0_300_s_3_300 = '-1.43750e-13*ic_cap*ic_cap+-1.00000e-13*ic_cap+2.03000e-11'
+ mcrdlm4l1_cf_w_0_300_s_9_000 = '-1.87500e-13*ic_cap*ic_cap+-1.25000e-13*ic_cap+3.25000e-11'
+ mcrdlm4l1_cf_w_2_400_s_0_300 = '-3.12500e-15*ic_cap*ic_cap+-2.50000e-15*ic_cap+2.34000e-12'
+ mcrdlm4l1_cf_w_2_400_s_0_360 = '-7.18750e-15*ic_cap*ic_cap+-6.25000e-15*ic_cap+2.80000e-12'
+ mcrdlm4l1_cf_w_2_400_s_0_450 = '-1.34375e-14*ic_cap*ic_cap+-8.75000e-15*ic_cap+3.49000e-12'
+ mcrdlm4l1_cf_w_2_400_s_0_600 = '-2.28125e-14*ic_cap*ic_cap+-1.62500e-14*ic_cap+4.61000e-12'
+ mcrdlm4l1_cf_w_2_400_s_0_800 = '-3.50000e-14*ic_cap*ic_cap+-2.25000e-14*ic_cap+6.08000e-12'
+ mcrdlm4l1_cf_w_2_400_s_1_000 = '-4.84375e-14*ic_cap*ic_cap+-3.12500e-14*ic_cap+7.53000e-12'
+ mcrdlm4l1_cf_w_2_400_s_1_200 = '-5.93750e-14*ic_cap*ic_cap+-4.00000e-14*ic_cap+8.92000e-12'
+ mcrdlm4l1_cf_w_2_400_s_2_100 = '-1.03125e-13*ic_cap*ic_cap+-6.25000e-14*ic_cap+1.47000e-11'
+ mcrdlm4l1_cf_w_2_400_s_3_300 = '-1.50000e-13*ic_cap*ic_cap+-1.00000e-13*ic_cap+2.11000e-11'
+ mcrdlm4l1_cf_w_2_400_s_9_000 = '-1.81250e-13*ic_cap*ic_cap+-1.25000e-13*ic_cap+3.55000e-11'
+ mcrdlm4m1_ca_w_0_300_s_0_300 = '-1.68750e-07*ic_cap*ic_cap+-1.00000e-07*ic_cap+1.91000e-05'
+ mcrdlm4m1_ca_w_0_300_s_0_360 = '-1.68750e-07*ic_cap*ic_cap+-1.00000e-07*ic_cap+1.91000e-05'
+ mcrdlm4m1_ca_w_0_300_s_0_450 = '-1.68750e-07*ic_cap*ic_cap+-1.00000e-07*ic_cap+1.91000e-05'
+ mcrdlm4m1_ca_w_0_300_s_0_600 = '-1.68750e-07*ic_cap*ic_cap+-1.00000e-07*ic_cap+1.91000e-05'
+ mcrdlm4m1_ca_w_0_300_s_0_800 = '-1.68750e-07*ic_cap*ic_cap+-1.00000e-07*ic_cap+1.91000e-05'
+ mcrdlm4m1_ca_w_0_300_s_1_000 = '-1.68750e-07*ic_cap*ic_cap+-1.00000e-07*ic_cap+1.91000e-05'
+ mcrdlm4m1_ca_w_0_300_s_1_200 = '-1.68750e-07*ic_cap*ic_cap+-1.00000e-07*ic_cap+1.91000e-05'
+ mcrdlm4m1_ca_w_0_300_s_2_100 = '-1.68750e-07*ic_cap*ic_cap+-1.00000e-07*ic_cap+1.91000e-05'
+ mcrdlm4m1_ca_w_0_300_s_3_300 = '-1.68750e-07*ic_cap*ic_cap+-1.00000e-07*ic_cap+1.91000e-05'
+ mcrdlm4m1_ca_w_0_300_s_9_000 = '-1.68750e-07*ic_cap*ic_cap+-1.00000e-07*ic_cap+1.91000e-05'
+ mcrdlm4m1_ca_w_2_400_s_0_300 = '-1.68750e-07*ic_cap*ic_cap+-1.00000e-07*ic_cap+1.91000e-05'
+ mcrdlm4m1_ca_w_2_400_s_0_360 = '-1.68750e-07*ic_cap*ic_cap+-1.00000e-07*ic_cap+1.91000e-05'
+ mcrdlm4m1_ca_w_2_400_s_0_450 = '-1.68750e-07*ic_cap*ic_cap+-1.00000e-07*ic_cap+1.91000e-05'
+ mcrdlm4m1_ca_w_2_400_s_0_600 = '-1.68750e-07*ic_cap*ic_cap+-1.00000e-07*ic_cap+1.91000e-05'
+ mcrdlm4m1_ca_w_2_400_s_0_800 = '-1.68750e-07*ic_cap*ic_cap+-1.00000e-07*ic_cap+1.91000e-05'
+ mcrdlm4m1_ca_w_2_400_s_1_000 = '-1.68750e-07*ic_cap*ic_cap+-1.00000e-07*ic_cap+1.91000e-05'
+ mcrdlm4m1_ca_w_2_400_s_1_200 = '-1.68750e-07*ic_cap*ic_cap+-1.00000e-07*ic_cap+1.91000e-05'
+ mcrdlm4m1_ca_w_2_400_s_2_100 = '-1.68750e-07*ic_cap*ic_cap+-1.00000e-07*ic_cap+1.91000e-05'
+ mcrdlm4m1_ca_w_2_400_s_3_300 = '-1.68750e-07*ic_cap*ic_cap+-1.00000e-07*ic_cap+1.91000e-05'
+ mcrdlm4m1_ca_w_2_400_s_9_000 = '-1.68750e-07*ic_cap*ic_cap+-1.00000e-07*ic_cap+1.91000e-05'
+ mcrdlm4m1_cc_w_0_300_s_0_300 = '-8.31250e-13*ic_cap*ic_cap+-4.50000e-13*ic_cap+1.06000e-10'
+ mcrdlm4m1_cc_w_0_300_s_0_360 = '-7.12500e-13*ic_cap*ic_cap+-4.00000e-13*ic_cap+9.83000e-11'
+ mcrdlm4m1_cc_w_0_300_s_0_450 = '-6.21875e-13*ic_cap*ic_cap+-3.62500e-13*ic_cap+8.89000e-11'
+ mcrdlm4m1_cc_w_0_300_s_0_600 = '-4.78125e-13*ic_cap*ic_cap+-2.87500e-13*ic_cap+7.61000e-11'
+ mcrdlm4m1_cc_w_0_300_s_0_800 = '-3.28125e-13*ic_cap*ic_cap+-2.12500e-13*ic_cap+6.34000e-11'
+ mcrdlm4m1_cc_w_0_300_s_1_000 = '-2.53125e-13*ic_cap*ic_cap+-1.62500e-13*ic_cap+5.41000e-11'
+ mcrdlm4m1_cc_w_0_300_s_1_200 = '-1.87500e-13*ic_cap*ic_cap+-1.50000e-13*ic_cap+4.69000e-11'
+ mcrdlm4m1_cc_w_0_300_s_2_100 = '-5.62500e-14*ic_cap*ic_cap+-5.00000e-14*ic_cap+2.85000e-11'
+ mcrdlm4m1_cc_w_0_300_s_3_300 = '6.25000e-15*ic_cap*ic_cap+1.72000e-11'
+ mcrdlm4m1_cc_w_0_300_s_9_000 = '2.53125e-14*ic_cap*ic_cap+1.87500e-14*ic_cap+2.40000e-12'
+ mcrdlm4m1_cc_w_2_400_s_0_300 = '-7.18750e-13*ic_cap*ic_cap+-3.75000e-13*ic_cap+1.27000e-10'
+ mcrdlm4m1_cc_w_2_400_s_0_360 = '-6.87500e-13*ic_cap*ic_cap+-5.00000e-13*ic_cap+1.19000e-10'
+ mcrdlm4m1_cc_w_2_400_s_0_450 = '-5.34375e-13*ic_cap*ic_cap+-3.12500e-13*ic_cap+1.07000e-10'
+ mcrdlm4m1_cc_w_2_400_s_0_600 = '-3.96875e-13*ic_cap*ic_cap+-2.37500e-13*ic_cap+9.22000e-11'
+ mcrdlm4m1_cc_w_2_400_s_0_800 = '-2.65625e-13*ic_cap*ic_cap+-1.62500e-13*ic_cap+7.71000e-11'
+ mcrdlm4m1_cc_w_2_400_s_1_000 = '-1.75000e-13*ic_cap*ic_cap+-1.25000e-13*ic_cap+6.58000e-11'
+ mcrdlm4m1_cc_w_2_400_s_1_200 = '-1.28125e-13*ic_cap*ic_cap+-8.75000e-14*ic_cap+5.74000e-11'
+ mcrdlm4m1_cc_w_2_400_s_2_100 = '-9.37500e-15*ic_cap*ic_cap+-1.25000e-14*ic_cap+3.55000e-11'
+ mcrdlm4m1_cc_w_2_400_s_3_300 = '5.00000e-14*ic_cap*ic_cap+2.50000e-14*ic_cap+2.16000e-11'
+ mcrdlm4m1_cc_w_2_400_s_9_000 = '4.31250e-14*ic_cap*ic_cap+3.50000e-14*ic_cap+3.19000e-12'
+ mcrdlm4m1_cf_w_0_300_s_0_300 = '-4.37500e-15*ic_cap*ic_cap+-2.50000e-15*ic_cap+2.81000e-12'
+ mcrdlm4m1_cf_w_0_300_s_0_360 = '-8.75000e-15*ic_cap*ic_cap+-5.00000e-15*ic_cap+3.36000e-12'
+ mcrdlm4m1_cf_w_0_300_s_0_450 = '-1.59375e-14*ic_cap*ic_cap+-8.75000e-15*ic_cap+4.22000e-12'
+ mcrdlm4m1_cf_w_0_300_s_0_600 = '-2.71875e-14*ic_cap*ic_cap+-1.62500e-14*ic_cap+5.60000e-12'
+ mcrdlm4m1_cf_w_0_300_s_0_800 = '-4.21875e-14*ic_cap*ic_cap+-2.37500e-14*ic_cap+7.26000e-12'
+ mcrdlm4m1_cf_w_0_300_s_1_000 = '-5.87500e-14*ic_cap*ic_cap+-3.25000e-14*ic_cap+8.94000e-12'
+ mcrdlm4m1_cf_w_0_300_s_1_200 = '-7.40625e-14*ic_cap*ic_cap+-4.37500e-14*ic_cap+1.06000e-11'
+ mcrdlm4m1_cf_w_0_300_s_2_100 = '-1.18750e-13*ic_cap*ic_cap+-7.50000e-14*ic_cap+1.72000e-11'
+ mcrdlm4m1_cf_w_0_300_s_3_300 = '-1.68750e-13*ic_cap*ic_cap+-1.00000e-13*ic_cap+2.35000e-11'
+ mcrdlm4m1_cf_w_0_300_s_9_000 = '-1.93750e-13*ic_cap*ic_cap+-1.25000e-13*ic_cap+3.53000e-11'
+ mcrdlm4m1_cf_w_2_400_s_0_300 = '-4.37500e-15*ic_cap*ic_cap+-2.50000e-15*ic_cap+2.83000e-12'
+ mcrdlm4m1_cf_w_2_400_s_0_360 = '-9.37500e-15*ic_cap*ic_cap+-5.00000e-15*ic_cap+3.38000e-12'
+ mcrdlm4m1_cf_w_2_400_s_0_450 = '-1.62500e-14*ic_cap*ic_cap+-1.00000e-14*ic_cap+4.20000e-12'
+ mcrdlm4m1_cf_w_2_400_s_0_600 = '-2.78125e-14*ic_cap*ic_cap+-1.62500e-14*ic_cap+5.55000e-12'
+ mcrdlm4m1_cf_w_2_400_s_0_800 = '-4.21875e-14*ic_cap*ic_cap+-2.62500e-14*ic_cap+7.30000e-12'
+ mcrdlm4m1_cf_w_2_400_s_1_000 = '-5.78125e-14*ic_cap*ic_cap+-3.37500e-14*ic_cap+9.03000e-12'
+ mcrdlm4m1_cf_w_2_400_s_1_200 = '-7.34375e-14*ic_cap*ic_cap+-4.37500e-14*ic_cap+1.07000e-11'
+ mcrdlm4m1_cf_w_2_400_s_2_100 = '-1.18750e-13*ic_cap*ic_cap+-7.50000e-14*ic_cap+1.73000e-11'
+ mcrdlm4m1_cf_w_2_400_s_3_300 = '-1.62500e-13*ic_cap*ic_cap+-1.00000e-13*ic_cap+2.43000e-11'
+ mcrdlm4m1_cf_w_2_400_s_9_000 = '-1.84375e-13*ic_cap*ic_cap+-1.12500e-13*ic_cap+3.85000e-11'
+ mcrdlm4m2_ca_w_0_300_s_0_300 = '-2.12500e-07*ic_cap*ic_cap+-1.25000e-07*ic_cap+2.49000e-05'
+ mcrdlm4m2_ca_w_0_300_s_0_360 = '-2.12500e-07*ic_cap*ic_cap+-1.25000e-07*ic_cap+2.49000e-05'
+ mcrdlm4m2_ca_w_0_300_s_0_450 = '-2.12500e-07*ic_cap*ic_cap+-1.25000e-07*ic_cap+2.49000e-05'
+ mcrdlm4m2_ca_w_0_300_s_0_600 = '-2.12500e-07*ic_cap*ic_cap+-1.25000e-07*ic_cap+2.49000e-05'
+ mcrdlm4m2_ca_w_0_300_s_0_800 = '-2.12500e-07*ic_cap*ic_cap+-1.25000e-07*ic_cap+2.49000e-05'
+ mcrdlm4m2_ca_w_0_300_s_1_000 = '-2.12500e-07*ic_cap*ic_cap+-1.25000e-07*ic_cap+2.49000e-05'
+ mcrdlm4m2_ca_w_0_300_s_1_200 = '-2.12500e-07*ic_cap*ic_cap+-1.25000e-07*ic_cap+2.49000e-05'
+ mcrdlm4m2_ca_w_0_300_s_2_100 = '-2.12500e-07*ic_cap*ic_cap+-1.25000e-07*ic_cap+2.49000e-05'
+ mcrdlm4m2_ca_w_0_300_s_3_300 = '-2.12500e-07*ic_cap*ic_cap+-1.25000e-07*ic_cap+2.49000e-05'
+ mcrdlm4m2_ca_w_0_300_s_9_000 = '-2.12500e-07*ic_cap*ic_cap+-1.25000e-07*ic_cap+2.49000e-05'
+ mcrdlm4m2_ca_w_2_400_s_0_300 = '-2.12500e-07*ic_cap*ic_cap+-1.25000e-07*ic_cap+2.49000e-05'
+ mcrdlm4m2_ca_w_2_400_s_0_360 = '-2.12500e-07*ic_cap*ic_cap+-1.25000e-07*ic_cap+2.49000e-05'
+ mcrdlm4m2_ca_w_2_400_s_0_450 = '-2.12500e-07*ic_cap*ic_cap+-1.25000e-07*ic_cap+2.49000e-05'
+ mcrdlm4m2_ca_w_2_400_s_0_600 = '-2.12500e-07*ic_cap*ic_cap+-1.25000e-07*ic_cap+2.49000e-05'
+ mcrdlm4m2_ca_w_2_400_s_0_800 = '-2.12500e-07*ic_cap*ic_cap+-1.25000e-07*ic_cap+2.49000e-05'
+ mcrdlm4m2_ca_w_2_400_s_1_000 = '-2.12500e-07*ic_cap*ic_cap+-1.25000e-07*ic_cap+2.49000e-05'
+ mcrdlm4m2_ca_w_2_400_s_1_200 = '-2.12500e-07*ic_cap*ic_cap+-1.25000e-07*ic_cap+2.49000e-05'
+ mcrdlm4m2_ca_w_2_400_s_2_100 = '-2.12500e-07*ic_cap*ic_cap+-1.25000e-07*ic_cap+2.49000e-05'
+ mcrdlm4m2_ca_w_2_400_s_3_300 = '-2.12500e-07*ic_cap*ic_cap+-1.25000e-07*ic_cap+2.49000e-05'
+ mcrdlm4m2_ca_w_2_400_s_9_000 = '-2.12500e-07*ic_cap*ic_cap+-1.25000e-07*ic_cap+2.49000e-05'
+ mcrdlm4m2_cc_w_0_300_s_0_300 = '-7.93750e-13*ic_cap*ic_cap+-4.75000e-13*ic_cap+1.04000e-10'
+ mcrdlm4m2_cc_w_0_300_s_0_360 = '-6.93750e-13*ic_cap*ic_cap+-3.75000e-13*ic_cap+9.66000e-11'
+ mcrdlm4m2_cc_w_0_300_s_0_450 = '-6.06250e-13*ic_cap*ic_cap+-3.50000e-13*ic_cap+8.72000e-11'
+ mcrdlm4m2_cc_w_0_300_s_0_600 = '-4.65625e-13*ic_cap*ic_cap+-2.62500e-13*ic_cap+7.42000e-11'
+ mcrdlm4m2_cc_w_0_300_s_0_800 = '-3.15625e-13*ic_cap*ic_cap+-2.12500e-13*ic_cap+6.13000e-11'
+ mcrdlm4m2_cc_w_0_300_s_1_000 = '-2.43750e-13*ic_cap*ic_cap+-1.50000e-13*ic_cap+5.18000e-11'
+ mcrdlm4m2_cc_w_0_300_s_1_200 = '-1.78125e-13*ic_cap*ic_cap+-1.37500e-13*ic_cap+4.45000e-11'
+ mcrdlm4m2_cc_w_0_300_s_2_100 = '-5.93750e-14*ic_cap*ic_cap+-3.75000e-14*ic_cap+2.60000e-11'
+ mcrdlm4m2_cc_w_0_300_s_3_300 = '6.25000e-15*ic_cap*ic_cap+1.48000e-11'
+ mcrdlm4m2_cc_w_0_300_s_9_000 = '1.84375e-14*ic_cap*ic_cap+8.75000e-15*ic_cap+1.71000e-12'
+ mcrdlm4m2_cc_w_2_400_s_0_300 = '-7.81250e-13*ic_cap*ic_cap+-3.75000e-13*ic_cap+1.24000e-10'
+ mcrdlm4m2_cc_w_2_400_s_0_360 = '-6.56250e-13*ic_cap*ic_cap+-3.75000e-13*ic_cap+1.15000e-10'
+ mcrdlm4m2_cc_w_2_400_s_0_450 = '-5.53125e-13*ic_cap*ic_cap+-3.37500e-13*ic_cap+1.04000e-10'
+ mcrdlm4m2_cc_w_2_400_s_0_600 = '-3.96875e-13*ic_cap*ic_cap+-2.37500e-13*ic_cap+8.88000e-11'
+ mcrdlm4m2_cc_w_2_400_s_0_800 = '-2.62500e-13*ic_cap*ic_cap+-1.75000e-13*ic_cap+7.37000e-11'
+ mcrdlm4m2_cc_w_2_400_s_1_000 = '-1.87500e-13*ic_cap*ic_cap+-1.25000e-13*ic_cap+6.26000e-11'
+ mcrdlm4m2_cc_w_2_400_s_1_200 = '-1.25000e-13*ic_cap*ic_cap+-7.50000e-14*ic_cap+5.40000e-11'
+ mcrdlm4m2_cc_w_2_400_s_2_100 = '-1.56250e-14*ic_cap*ic_cap+-1.25000e-14*ic_cap+3.24000e-11'
+ mcrdlm4m2_cc_w_2_400_s_3_300 = '3.75000e-14*ic_cap*ic_cap+2.50000e-14*ic_cap+1.89000e-11'
+ mcrdlm4m2_cc_w_2_400_s_9_000 = '3.12500e-14*ic_cap*ic_cap+2.25000e-14*ic_cap+2.37000e-12'
+ mcrdlm4m2_cf_w_0_300_s_0_300 = '-3.75000e-15*ic_cap*ic_cap+-2.50000e-15*ic_cap+3.63000e-12'
+ mcrdlm4m2_cf_w_0_300_s_0_360 = '-9.68750e-15*ic_cap*ic_cap+-6.25000e-15*ic_cap+4.34000e-12'
+ mcrdlm4m2_cf_w_0_300_s_0_450 = '-1.84375e-14*ic_cap*ic_cap+-1.12500e-14*ic_cap+5.42000e-12'
+ mcrdlm4m2_cf_w_0_300_s_0_600 = '-3.25000e-14*ic_cap*ic_cap+-2.00000e-14*ic_cap+7.17000e-12'
+ mcrdlm4m2_cf_w_0_300_s_0_800 = '-5.00000e-14*ic_cap*ic_cap+-3.00000e-14*ic_cap+9.27000e-12'
+ mcrdlm4m2_cf_w_0_300_s_1_000 = '-7.18750e-14*ic_cap*ic_cap+-3.75000e-14*ic_cap+1.14000e-11'
+ mcrdlm4m2_cf_w_0_300_s_1_200 = '-8.12500e-14*ic_cap*ic_cap+-5.00000e-14*ic_cap+1.33000e-11'
+ mcrdlm4m2_cf_w_0_300_s_2_100 = '-1.40625e-13*ic_cap*ic_cap+-8.75000e-14*ic_cap+2.12000e-11'
+ mcrdlm4m2_cf_w_0_300_s_3_300 = '-1.84375e-13*ic_cap*ic_cap+-1.12500e-13*ic_cap+2.81000e-11'
+ mcrdlm4m2_cf_w_0_300_s_9_000 = '-2.00000e-13*ic_cap*ic_cap+-1.25000e-13*ic_cap+3.91000e-11'
+ mcrdlm4m2_cf_w_2_400_s_0_300 = '-3.75000e-15*ic_cap*ic_cap+-2.50000e-15*ic_cap+3.65000e-12'
+ mcrdlm4m2_cf_w_2_400_s_0_360 = '-1.00000e-14*ic_cap*ic_cap+-5.00000e-15*ic_cap+4.36000e-12'
+ mcrdlm4m2_cf_w_2_400_s_0_450 = '-1.81250e-14*ic_cap*ic_cap+-1.25000e-14*ic_cap+5.41000e-12'
+ mcrdlm4m2_cf_w_2_400_s_0_600 = '-3.25000e-14*ic_cap*ic_cap+-2.00000e-14*ic_cap+7.12000e-12'
+ mcrdlm4m2_cf_w_2_400_s_0_800 = '-5.03125e-14*ic_cap*ic_cap+-3.12500e-14*ic_cap+9.33000e-12'
+ mcrdlm4m2_cf_w_2_400_s_1_000 = '-7.18750e-14*ic_cap*ic_cap+-3.75000e-14*ic_cap+1.15000e-11'
+ mcrdlm4m2_cf_w_2_400_s_1_200 = '-8.43750e-14*ic_cap*ic_cap+-6.25000e-14*ic_cap+1.35000e-11'
+ mcrdlm4m2_cf_w_2_400_s_2_100 = '-1.40625e-13*ic_cap*ic_cap+-8.75000e-14*ic_cap+2.14000e-11'
+ mcrdlm4m2_cf_w_2_400_s_3_300 = '-1.78125e-13*ic_cap*ic_cap+-1.12500e-13*ic_cap+2.91000e-11'
+ mcrdlm4m2_cf_w_2_400_s_9_000 = '-1.87500e-13*ic_cap*ic_cap+-1.25000e-13*ic_cap+4.26000e-11'
+ mcrdlm4m3_ca_w_0_300_s_0_300 = '-1.75938e-06*ic_cap*ic_cap+-8.62500e-07*ic_cap+9.25000e-05'
+ mcrdlm4m3_ca_w_0_300_s_0_360 = '-1.75938e-06*ic_cap*ic_cap+-8.62500e-07*ic_cap+9.25000e-05'
+ mcrdlm4m3_ca_w_0_300_s_0_450 = '-1.75938e-06*ic_cap*ic_cap+-8.62500e-07*ic_cap+9.25000e-05'
+ mcrdlm4m3_ca_w_0_300_s_0_600 = '-1.75938e-06*ic_cap*ic_cap+-8.62500e-07*ic_cap+9.25000e-05'
+ mcrdlm4m3_ca_w_0_300_s_0_800 = '-1.75938e-06*ic_cap*ic_cap+-8.62500e-07*ic_cap+9.25000e-05'
+ mcrdlm4m3_ca_w_0_300_s_1_000 = '-1.75938e-06*ic_cap*ic_cap+-8.62500e-07*ic_cap+9.25000e-05'
+ mcrdlm4m3_ca_w_0_300_s_1_200 = '-1.75938e-06*ic_cap*ic_cap+-8.62500e-07*ic_cap+9.25000e-05'
+ mcrdlm4m3_ca_w_0_300_s_2_100 = '-1.75938e-06*ic_cap*ic_cap+-8.62500e-07*ic_cap+9.25000e-05'
+ mcrdlm4m3_ca_w_0_300_s_3_300 = '-1.75938e-06*ic_cap*ic_cap+-8.62500e-07*ic_cap+9.25000e-05'
+ mcrdlm4m3_ca_w_0_300_s_9_000 = '-1.75938e-06*ic_cap*ic_cap+-8.62500e-07*ic_cap+9.25000e-05'
+ mcrdlm4m3_ca_w_2_400_s_0_300 = '-1.75938e-06*ic_cap*ic_cap+-8.62500e-07*ic_cap+9.25000e-05'
+ mcrdlm4m3_ca_w_2_400_s_0_360 = '-1.75938e-06*ic_cap*ic_cap+-8.62500e-07*ic_cap+9.25000e-05'
+ mcrdlm4m3_ca_w_2_400_s_0_450 = '-1.75938e-06*ic_cap*ic_cap+-8.62500e-07*ic_cap+9.25000e-05'
+ mcrdlm4m3_ca_w_2_400_s_0_600 = '-1.75938e-06*ic_cap*ic_cap+-8.62500e-07*ic_cap+9.25000e-05'
+ mcrdlm4m3_ca_w_2_400_s_0_800 = '-1.75938e-06*ic_cap*ic_cap+-8.62500e-07*ic_cap+9.25000e-05'
+ mcrdlm4m3_ca_w_2_400_s_1_000 = '-1.75938e-06*ic_cap*ic_cap+-8.62500e-07*ic_cap+9.25000e-05'
+ mcrdlm4m3_ca_w_2_400_s_1_200 = '-1.75938e-06*ic_cap*ic_cap+-8.62500e-07*ic_cap+9.25000e-05'
+ mcrdlm4m3_ca_w_2_400_s_2_100 = '-1.75938e-06*ic_cap*ic_cap+-8.62500e-07*ic_cap+9.25000e-05'
+ mcrdlm4m3_ca_w_2_400_s_3_300 = '-1.75938e-06*ic_cap*ic_cap+-8.62500e-07*ic_cap+9.25000e-05'
+ mcrdlm4m3_ca_w_2_400_s_9_000 = '-1.75938e-06*ic_cap*ic_cap+-8.62500e-07*ic_cap+9.25000e-05'
+ mcrdlm4m3_cc_w_0_300_s_0_300 = '-6.15625e-13*ic_cap*ic_cap+-3.62500e-13*ic_cap+9.29000e-11'
+ mcrdlm4m3_cc_w_0_300_s_0_360 = '-4.90625e-13*ic_cap*ic_cap+-2.87500e-13*ic_cap+8.49000e-11'
+ mcrdlm4m3_cc_w_0_300_s_0_450 = '-4.06250e-13*ic_cap*ic_cap+-2.50000e-13*ic_cap+7.50000e-11'
+ mcrdlm4m3_cc_w_0_300_s_0_600 = '-2.71875e-13*ic_cap*ic_cap+-1.62500e-13*ic_cap+6.16000e-11'
+ mcrdlm4m3_cc_w_0_300_s_0_800 = '-1.65625e-13*ic_cap*ic_cap+-1.12500e-13*ic_cap+4.89000e-11'
+ mcrdlm4m3_cc_w_0_300_s_1_000 = '-9.37500e-14*ic_cap*ic_cap+-7.50000e-14*ic_cap+3.94000e-11'
+ mcrdlm4m3_cc_w_0_300_s_1_200 = '-4.68750e-14*ic_cap*ic_cap+-3.75000e-14*ic_cap+3.23000e-11'
+ mcrdlm4m3_cc_w_0_300_s_2_100 = '9.37500e-15*ic_cap*ic_cap+1.25000e-14*ic_cap+1.56000e-11'
+ mcrdlm4m3_cc_w_0_300_s_3_300 = '2.59375e-14*ic_cap*ic_cap+1.62500e-14*ic_cap+7.52000e-12'
+ mcrdlm4m3_cc_w_0_300_s_9_000 = '5.96875e-15*ic_cap*ic_cap+7.37500e-15*ic_cap+5.95000e-13'
+ mcrdlm4m3_cc_w_2_400_s_0_300 = '-6.43750e-13*ic_cap*ic_cap+-3.00000e-13*ic_cap+1.09000e-10'
+ mcrdlm4m3_cc_w_2_400_s_0_360 = '-4.90625e-13*ic_cap*ic_cap+-2.62500e-13*ic_cap+9.95000e-11'
+ mcrdlm4m3_cc_w_2_400_s_0_450 = '-3.87500e-13*ic_cap*ic_cap+-2.25000e-13*ic_cap+8.85000e-11'
+ mcrdlm4m3_cc_w_2_400_s_0_600 = '-2.50000e-13*ic_cap*ic_cap+-1.50000e-13*ic_cap+7.37000e-11'
+ mcrdlm4m3_cc_w_2_400_s_0_800 = '-1.40625e-13*ic_cap*ic_cap+-8.75000e-14*ic_cap+5.92000e-11'
+ mcrdlm4m3_cc_w_2_400_s_1_000 = '-5.93750e-14*ic_cap*ic_cap+-6.25000e-14*ic_cap+4.84000e-11'
+ mcrdlm4m3_cc_w_2_400_s_1_200 = '-2.50000e-14*ic_cap*ic_cap+-2.50000e-14*ic_cap+4.06000e-11'
+ mcrdlm4m3_cc_w_2_400_s_2_100 = '3.75000e-14*ic_cap*ic_cap+2.50000e-14*ic_cap+2.16000e-11'
+ mcrdlm4m3_cc_w_2_400_s_3_300 = '5.00000e-14*ic_cap*ic_cap+2.50000e-14*ic_cap+1.11000e-11'
+ mcrdlm4m3_cc_w_2_400_s_9_000 = '1.75000e-14*ic_cap*ic_cap+1.37500e-14*ic_cap+9.05000e-13'
+ mcrdlm4m3_cf_w_0_300_s_0_300 = '-1.49063e-13*ic_cap*ic_cap+-7.12500e-14*ic_cap+1.24000e-11'
+ mcrdlm4m3_cf_w_0_300_s_0_360 = '-1.87500e-13*ic_cap*ic_cap+-1.00000e-13*ic_cap+1.46000e-11'
+ mcrdlm4m3_cf_w_0_300_s_0_450 = '-2.34375e-13*ic_cap*ic_cap+-1.12500e-13*ic_cap+1.77000e-11'
+ mcrdlm4m3_cf_w_0_300_s_0_600 = '-3.00000e-13*ic_cap*ic_cap+-1.50000e-13*ic_cap+2.23000e-11'
+ mcrdlm4m3_cf_w_0_300_s_0_800 = '-3.62500e-13*ic_cap*ic_cap+-2.00000e-13*ic_cap+2.74000e-11'
+ mcrdlm4m3_cf_w_0_300_s_1_000 = '-4.12500e-13*ic_cap*ic_cap+-2.25000e-13*ic_cap+3.19000e-11'
+ mcrdlm4m3_cf_w_0_300_s_1_200 = '-4.43750e-13*ic_cap*ic_cap+-2.50000e-13*ic_cap+3.56000e-11'
+ mcrdlm4m3_cf_w_0_300_s_2_100 = '-5.03125e-13*ic_cap*ic_cap+-2.87500e-13*ic_cap+4.70000e-11'
+ mcrdlm4m3_cf_w_0_300_s_3_300 = '-5.21875e-13*ic_cap*ic_cap+-3.12500e-13*ic_cap+5.39000e-11'
+ mcrdlm4m3_cf_w_0_300_s_9_000 = '-5.06250e-13*ic_cap*ic_cap+-3.00000e-13*ic_cap+6.04000e-11'
+ mcrdlm4m3_cf_w_2_400_s_0_300 = '-1.45313e-13*ic_cap*ic_cap+-8.12500e-14*ic_cap+1.24000e-11'
+ mcrdlm4m3_cf_w_2_400_s_0_360 = '-1.84375e-13*ic_cap*ic_cap+-8.75000e-14*ic_cap+1.46000e-11'
+ mcrdlm4m3_cf_w_2_400_s_0_450 = '-2.34375e-13*ic_cap*ic_cap+-1.12500e-13*ic_cap+1.77000e-11'
+ mcrdlm4m3_cf_w_2_400_s_0_600 = '-3.00000e-13*ic_cap*ic_cap+-1.50000e-13*ic_cap+2.23000e-11'
+ mcrdlm4m3_cf_w_2_400_s_0_800 = '-3.62500e-13*ic_cap*ic_cap+-2.00000e-13*ic_cap+2.75000e-11'
+ mcrdlm4m3_cf_w_2_400_s_1_000 = '-4.09375e-13*ic_cap*ic_cap+-2.12500e-13*ic_cap+3.20000e-11'
+ mcrdlm4m3_cf_w_2_400_s_1_200 = '-4.40625e-13*ic_cap*ic_cap+-2.37500e-13*ic_cap+3.58000e-11'
+ mcrdlm4m3_cf_w_2_400_s_2_100 = '-5.03125e-13*ic_cap*ic_cap+-2.87500e-13*ic_cap+4.75000e-11'
+ mcrdlm4m3_cf_w_2_400_s_3_300 = '-5.25000e-13*ic_cap*ic_cap+-3.00000e-13*ic_cap+5.59000e-11'
+ mcrdlm4m3_cf_w_2_400_s_9_000 = '-4.96875e-13*ic_cap*ic_cap+-2.87500e-13*ic_cap+6.53000e-11'
+ mcrdlm4p1_ca_w_0_300_s_0_300 = '-1.31250e-07*ic_cap*ic_cap+-7.50000e-08*ic_cap+1.41000e-05'
+ mcrdlm4p1_ca_w_0_300_s_0_360 = '-1.31250e-07*ic_cap*ic_cap+-7.50000e-08*ic_cap+1.41000e-05'
+ mcrdlm4p1_ca_w_0_300_s_0_450 = '-1.31250e-07*ic_cap*ic_cap+-7.50000e-08*ic_cap+1.41000e-05'
+ mcrdlm4p1_ca_w_0_300_s_0_600 = '-1.31250e-07*ic_cap*ic_cap+-7.50000e-08*ic_cap+1.41000e-05'
+ mcrdlm4p1_ca_w_0_300_s_0_800 = '-1.31250e-07*ic_cap*ic_cap+-7.50000e-08*ic_cap+1.41000e-05'
+ mcrdlm4p1_ca_w_0_300_s_1_000 = '-1.31250e-07*ic_cap*ic_cap+-7.50000e-08*ic_cap+1.41000e-05'
+ mcrdlm4p1_ca_w_0_300_s_1_200 = '-1.31250e-07*ic_cap*ic_cap+-7.50000e-08*ic_cap+1.41000e-05'
+ mcrdlm4p1_ca_w_0_300_s_2_100 = '-1.31250e-07*ic_cap*ic_cap+-7.50000e-08*ic_cap+1.41000e-05'
+ mcrdlm4p1_ca_w_0_300_s_3_300 = '-1.31250e-07*ic_cap*ic_cap+-7.50000e-08*ic_cap+1.41000e-05'
+ mcrdlm4p1_ca_w_0_300_s_9_000 = '-1.31250e-07*ic_cap*ic_cap+-7.50000e-08*ic_cap+1.41000e-05'
+ mcrdlm4p1_ca_w_2_400_s_0_300 = '-1.31250e-07*ic_cap*ic_cap+-7.50000e-08*ic_cap+1.41000e-05'
+ mcrdlm4p1_ca_w_2_400_s_0_360 = '-1.31250e-07*ic_cap*ic_cap+-7.50000e-08*ic_cap+1.41000e-05'
+ mcrdlm4p1_ca_w_2_400_s_0_450 = '-1.31250e-07*ic_cap*ic_cap+-7.50000e-08*ic_cap+1.41000e-05'
+ mcrdlm4p1_ca_w_2_400_s_0_600 = '-1.31250e-07*ic_cap*ic_cap+-7.50000e-08*ic_cap+1.41000e-05'
+ mcrdlm4p1_ca_w_2_400_s_0_800 = '-1.31250e-07*ic_cap*ic_cap+-7.50000e-08*ic_cap+1.41000e-05'
+ mcrdlm4p1_ca_w_2_400_s_1_000 = '-1.31250e-07*ic_cap*ic_cap+-7.50000e-08*ic_cap+1.41000e-05'
+ mcrdlm4p1_ca_w_2_400_s_1_200 = '-1.31250e-07*ic_cap*ic_cap+-7.50000e-08*ic_cap+1.41000e-05'
+ mcrdlm4p1_ca_w_2_400_s_2_100 = '-1.31250e-07*ic_cap*ic_cap+-7.50000e-08*ic_cap+1.41000e-05'
+ mcrdlm4p1_ca_w_2_400_s_3_300 = '-1.31250e-07*ic_cap*ic_cap+-7.50000e-08*ic_cap+1.41000e-05'
+ mcrdlm4p1_ca_w_2_400_s_9_000 = '-1.31250e-07*ic_cap*ic_cap+-7.50000e-08*ic_cap+1.41000e-05'
+ mcrdlm4p1_cc_w_0_300_s_0_300 = '-8.21875e-13*ic_cap*ic_cap+-4.37500e-13*ic_cap+1.07000e-10'
+ mcrdlm4p1_cc_w_0_300_s_0_360 = '-7.18750e-13*ic_cap*ic_cap+-4.00000e-13*ic_cap+9.96000e-11'
+ mcrdlm4p1_cc_w_0_300_s_0_450 = '-6.34375e-13*ic_cap*ic_cap+-3.87500e-13*ic_cap+9.03000e-11'
+ mcrdlm4p1_cc_w_0_300_s_0_600 = '-4.68750e-13*ic_cap*ic_cap+-3.00000e-13*ic_cap+7.75000e-11'
+ mcrdlm4p1_cc_w_0_300_s_0_800 = '-3.46875e-13*ic_cap*ic_cap+-2.37500e-13*ic_cap+6.54000e-11'
+ mcrdlm4p1_cc_w_0_300_s_1_000 = '-2.65625e-13*ic_cap*ic_cap+-1.87500e-13*ic_cap+5.63000e-11'
+ mcrdlm4p1_cc_w_0_300_s_1_200 = '-2.00000e-13*ic_cap*ic_cap+-1.50000e-13*ic_cap+4.93000e-11'
+ mcrdlm4p1_cc_w_0_300_s_2_100 = '-6.25000e-14*ic_cap*ic_cap+-5.00000e-14*ic_cap+3.14000e-11'
+ mcrdlm4p1_cc_w_0_300_s_9_000 = '3.96875e-14*ic_cap*ic_cap+2.62500e-14*ic_cap+3.56000e-12'
+ mcrdlm4p1_cc_w_2_400_s_0_300 = '-7.81250e-13*ic_cap*ic_cap+-3.75000e-13*ic_cap+1.31000e-10'
+ mcrdlm4p1_cc_w_2_400_s_0_360 = '-6.56250e-13*ic_cap*ic_cap+-3.75000e-13*ic_cap+1.22000e-10'
+ mcrdlm4p1_cc_w_2_400_s_0_450 = '-5.62500e-13*ic_cap*ic_cap+-2.50000e-13*ic_cap+1.11000e-10'
+ mcrdlm4p1_cc_w_2_400_s_0_600 = '-4.09375e-13*ic_cap*ic_cap+-2.37500e-13*ic_cap+9.61000e-11'
+ mcrdlm4p1_cc_w_2_400_s_0_800 = '-2.65625e-13*ic_cap*ic_cap+-1.62500e-13*ic_cap+8.09000e-11'
+ mcrdlm4p1_cc_w_2_400_s_1_000 = '-1.81250e-13*ic_cap*ic_cap+-1.50000e-13*ic_cap+6.97000e-11'
+ mcrdlm4p1_cc_w_2_400_s_1_200 = '-1.28125e-13*ic_cap*ic_cap+-1.12500e-13*ic_cap+6.13000e-11'
+ mcrdlm4p1_cc_w_2_400_s_2_100 = '-3.12500e-15*ic_cap*ic_cap+-1.25000e-14*ic_cap+3.94000e-11'
+ mcrdlm4p1_cc_w_2_400_s_3_300 = '5.62500e-14*ic_cap*ic_cap+2.50000e-14*ic_cap+2.52000e-11'
+ mcrdlm4p1_cc_w_2_400_s_9_000 = '6.46875e-14*ic_cap*ic_cap+4.37500e-14*ic_cap+4.65000e-12'
+ mcrdlm4p1_cf_w_0_300_s_0_300 = '-4.37500e-15*ic_cap*ic_cap+-2.50000e-15*ic_cap+2.09000e-12'
+ mcrdlm4p1_cf_w_0_300_s_0_360 = '-8.12500e-15*ic_cap*ic_cap+-5.00000e-15*ic_cap+2.51000e-12'
+ mcrdlm4p1_cf_w_0_300_s_0_450 = '-1.40625e-14*ic_cap*ic_cap+-8.75000e-15*ic_cap+3.16000e-12'
+ mcrdlm4p1_cf_w_0_300_s_0_600 = '-2.43750e-14*ic_cap*ic_cap+-1.50000e-14*ic_cap+4.23000e-12'
+ mcrdlm4p1_cf_w_0_300_s_0_800 = '-3.59375e-14*ic_cap*ic_cap+-2.37500e-14*ic_cap+5.46000e-12'
+ mcrdlm4p1_cf_w_0_300_s_1_000 = '-4.84375e-14*ic_cap*ic_cap+-2.87500e-14*ic_cap+6.76000e-12'
+ mcrdlm4p1_cf_w_0_300_s_1_200 = '-5.87500e-14*ic_cap*ic_cap+-3.50000e-14*ic_cap+8.01000e-12'
+ mcrdlm4p1_cf_w_0_300_s_2_100 = '-1.03125e-13*ic_cap*ic_cap+-6.25000e-14*ic_cap+1.34000e-11'
+ mcrdlm4p1_cf_w_0_300_s_3_300 = '-1.50000e-13*ic_cap*ic_cap+-1.00000e-13*ic_cap+1.88000e-11'
+ mcrdlm4p1_cf_w_0_300_s_9_000 = '-1.84375e-13*ic_cap*ic_cap+-1.37500e-13*ic_cap+3.09000e-11'
+ mcrdlm4p1_cf_w_2_400_s_0_300 = '-4.68750e-15*ic_cap*ic_cap+-3.75000e-15*ic_cap+2.13000e-12'
+ mcrdlm4p1_cf_w_2_400_s_0_360 = '-9.06250e-15*ic_cap*ic_cap+-6.25000e-15*ic_cap+2.55000e-12'
+ mcrdlm4p1_cf_w_2_400_s_0_450 = '-1.46875e-14*ic_cap*ic_cap+-8.75000e-15*ic_cap+3.17000e-12'
+ mcrdlm4p1_cf_w_2_400_s_0_600 = '-2.37500e-14*ic_cap*ic_cap+-1.50000e-14*ic_cap+4.18000e-12'
+ mcrdlm4p1_cf_w_2_400_s_0_800 = '-3.59375e-14*ic_cap*ic_cap+-2.37500e-14*ic_cap+5.52000e-12'
+ mcrdlm4p1_cf_w_2_400_s_1_000 = '-4.81250e-14*ic_cap*ic_cap+-3.00000e-14*ic_cap+6.83000e-12'
+ mcrdlm4p1_cf_w_2_400_s_1_200 = '-5.96875e-14*ic_cap*ic_cap+-3.87500e-14*ic_cap+8.11000e-12'
+ mcrdlm4p1_cf_w_2_400_s_2_100 = '-1.03125e-13*ic_cap*ic_cap+-6.25000e-14*ic_cap+1.34000e-11'
+ mcrdlm4p1_cf_w_2_400_s_3_300 = '-1.46875e-13*ic_cap*ic_cap+-8.75000e-14*ic_cap+1.94000e-11'
+ mcrdlm4p1_cf_w_2_400_s_9_000 = '-1.93750e-13*ic_cap*ic_cap+-1.25000e-13*ic_cap+3.39000e-11'
+ mcrdlm5_ca_w_10_000_s_10_000 = '-6.31250e-08*ic_cap*ic_cap+-3.75000e-08*ic_cap+5.44000e-06'
+ mcrdlm5_ca_w_10_000_s_12_000 = '-6.31250e-08*ic_cap*ic_cap+-3.75000e-08*ic_cap+5.44000e-06'
+ mcrdlm5_ca_w_10_000_s_30_000 = '-6.31250e-08*ic_cap*ic_cap+-3.75000e-08*ic_cap+5.44000e-06'
+ mcrdlm5_ca_w_10_000_s_5_000 = '-6.31250e-08*ic_cap*ic_cap+-3.75000e-08*ic_cap+5.44000e-06'
+ mcrdlm5_ca_w_10_000_s_8_000 = '-6.31250e-08*ic_cap*ic_cap+-3.75000e-08*ic_cap+5.44000e-06'
+ mcrdlm5_ca_w_40_000_s_10_000 = '-6.31250e-08*ic_cap*ic_cap+-3.75000e-08*ic_cap+5.44000e-06'
+ mcrdlm5_ca_w_40_000_s_12_000 = '-6.31250e-08*ic_cap*ic_cap+-3.75000e-08*ic_cap+5.44000e-06'
+ mcrdlm5_ca_w_40_000_s_30_000 = '-6.31250e-08*ic_cap*ic_cap+-3.75000e-08*ic_cap+5.44000e-06'
+ mcrdlm5_ca_w_40_000_s_5_000 = '-6.31250e-08*ic_cap*ic_cap+-3.75000e-08*ic_cap+5.44000e-06'
+ mcrdlm5_ca_w_40_000_s_8_000 = '-6.31250e-08*ic_cap*ic_cap+-3.75000e-08*ic_cap+5.44000e-06'
+ mcrdlm5_cc_w_10_000_s_10_000 = '-2.18750e-13*ic_cap*ic_cap+-1.50000e-13*ic_cap+2.63000e-11'
+ mcrdlm5_cc_w_10_000_s_12_000 = '-1.75000e-13*ic_cap*ic_cap+-1.25000e-13*ic_cap+2.25000e-11'
+ mcrdlm5_cc_w_10_000_s_30_000 = '-5.53125e-14*ic_cap*ic_cap+-4.62500e-14*ic_cap+8.70000e-12'
+ mcrdlm5_cc_w_10_000_s_5_000 = '-5.25000e-13*ic_cap*ic_cap+-3.25000e-13*ic_cap+4.54000e-11'
+ mcrdlm5_cc_w_10_000_s_8_000 = '-2.90625e-13*ic_cap*ic_cap+-1.87500e-13*ic_cap+3.16000e-11'
+ mcrdlm5_cc_w_40_000_s_10_000 = '-2.25000e-13*ic_cap*ic_cap+-1.50000e-13*ic_cap+3.62000e-11'
+ mcrdlm5_cc_w_40_000_s_12_000 = '-1.78125e-13*ic_cap*ic_cap+-1.12500e-13*ic_cap+3.20000e-11'
+ mcrdlm5_cc_w_40_000_s_30_000 = '-5.62500e-14*ic_cap*ic_cap+-5.00000e-14*ic_cap+1.57000e-11'
+ mcrdlm5_cc_w_40_000_s_5_000 = '-5.40625e-13*ic_cap*ic_cap+-3.37500e-13*ic_cap+5.67000e-11'
+ mcrdlm5_cc_w_40_000_s_8_000 = '-2.93750e-13*ic_cap*ic_cap+-2.00000e-13*ic_cap+4.19000e-11'
+ mcrdlm5_cf_w_10_000_s_10_000 = '-1.09375e-13*ic_cap*ic_cap+-6.25000e-14*ic_cap+1.92000e-11'
+ mcrdlm5_cf_w_10_000_s_12_000 = '-1.28125e-13*ic_cap*ic_cap+-8.75000e-14*ic_cap+2.15000e-11'
+ mcrdlm5_cf_w_10_000_s_30_000 = '-2.15625e-13*ic_cap*ic_cap+-1.37500e-13*ic_cap+3.26000e-11'
+ mcrdlm5_cf_w_10_000_s_5_000 = '-2.81250e-14*ic_cap*ic_cap+-1.25000e-14*ic_cap+1.14000e-11'
+ mcrdlm5_cf_w_10_000_s_8_000 = '-8.12500e-14*ic_cap*ic_cap+-5.00000e-14*ic_cap+1.64000e-11'
+ mcrdlm5_cf_w_40_000_s_10_000 = '-1.09375e-13*ic_cap*ic_cap+-6.25000e-14*ic_cap+1.92000e-11'
+ mcrdlm5_cf_w_40_000_s_12_000 = '-1.31250e-13*ic_cap*ic_cap+-7.50000e-14*ic_cap+2.16000e-11'
+ mcrdlm5_cf_w_40_000_s_30_000 = '-2.00000e-13*ic_cap*ic_cap+-1.25000e-13*ic_cap+3.38000e-11'
+ mcrdlm5_cf_w_40_000_s_5_000 = '-3.43750e-14*ic_cap*ic_cap+-1.25000e-14*ic_cap+1.14000e-11'
+ mcrdlm5_cf_w_40_000_s_8_000 = '-8.75000e-14*ic_cap*ic_cap+-5.00000e-14*ic_cap+1.64000e-11'
+ mcrdlm5d_ca_w_1_600_s_10_000 = '-1.15625e-07*ic_cap*ic_cap+-6.25000e-08*ic_cap+1.24000e-05'
+ mcrdlm5d_ca_w_1_600_s_12_000 = '-1.15625e-07*ic_cap*ic_cap+-6.25000e-08*ic_cap+1.24000e-05'
+ mcrdlm5d_ca_w_1_600_s_1_600 = '-1.15625e-07*ic_cap*ic_cap+-6.25000e-08*ic_cap+1.24000e-05'
+ mcrdlm5d_ca_w_1_600_s_1_700 = '-1.15625e-07*ic_cap*ic_cap+-6.25000e-08*ic_cap+1.24000e-05'
+ mcrdlm5d_ca_w_1_600_s_1_900 = '-1.15625e-07*ic_cap*ic_cap+-6.25000e-08*ic_cap+1.24000e-05'
+ mcrdlm5d_ca_w_1_600_s_2_000 = '-1.15625e-07*ic_cap*ic_cap+-6.25000e-08*ic_cap+1.24000e-05'
+ mcrdlm5d_ca_w_1_600_s_2_400 = '-1.15625e-07*ic_cap*ic_cap+-6.25000e-08*ic_cap+1.24000e-05'
+ mcrdlm5d_ca_w_1_600_s_2_800 = '-1.15625e-07*ic_cap*ic_cap+-6.25000e-08*ic_cap+1.24000e-05'
+ mcrdlm5d_ca_w_1_600_s_3_200 = '-1.15625e-07*ic_cap*ic_cap+-6.25000e-08*ic_cap+1.24000e-05'
+ mcrdlm5d_ca_w_1_600_s_4_800 = '-1.15625e-07*ic_cap*ic_cap+-6.25000e-08*ic_cap+1.24000e-05'
+ mcrdlm5d_ca_w_4_000_s_10_000 = '-1.15625e-07*ic_cap*ic_cap+-6.25000e-08*ic_cap+1.24000e-05'
+ mcrdlm5d_ca_w_4_000_s_12_000 = '-1.15625e-07*ic_cap*ic_cap+-6.25000e-08*ic_cap+1.24000e-05'
+ mcrdlm5d_ca_w_4_000_s_1_600 = '-1.15625e-07*ic_cap*ic_cap+-6.25000e-08*ic_cap+1.24000e-05'
+ mcrdlm5d_ca_w_4_000_s_1_700 = '-1.15625e-07*ic_cap*ic_cap+-6.25000e-08*ic_cap+1.24000e-05'
+ mcrdlm5d_ca_w_4_000_s_1_900 = '-1.15625e-07*ic_cap*ic_cap+-6.25000e-08*ic_cap+1.24000e-05'
+ mcrdlm5d_ca_w_4_000_s_2_000 = '-1.15625e-07*ic_cap*ic_cap+-6.25000e-08*ic_cap+1.24000e-05'
+ mcrdlm5d_ca_w_4_000_s_2_400 = '-1.15625e-07*ic_cap*ic_cap+-6.25000e-08*ic_cap+1.24000e-05'
+ mcrdlm5d_ca_w_4_000_s_2_800 = '-1.15625e-07*ic_cap*ic_cap+-6.25000e-08*ic_cap+1.24000e-05'
+ mcrdlm5d_ca_w_4_000_s_3_200 = '-1.15625e-07*ic_cap*ic_cap+-6.25000e-08*ic_cap+1.24000e-05'
+ mcrdlm5d_ca_w_4_000_s_4_800 = '-1.15625e-07*ic_cap*ic_cap+-6.25000e-08*ic_cap+1.24000e-05'
+ mcrdlm5d_cc_w_1_600_s_10_000 = '5.46875e-14*ic_cap*ic_cap+3.62500e-14*ic_cap+4.51000e-12'
+ mcrdlm5d_cc_w_1_600_s_12_000 = '4.50000e-14*ic_cap*ic_cap+3.00000e-14*ic_cap+2.62000e-12'
+ mcrdlm5d_cc_w_1_600_s_1_600 = '-3.96875e-13*ic_cap*ic_cap+-2.62500e-13*ic_cap+6.64000e-11'
+ mcrdlm5d_cc_w_1_600_s_1_700 = '-3.43750e-13*ic_cap*ic_cap+-2.50000e-13*ic_cap+6.25000e-11'
+ mcrdlm5d_cc_w_1_600_s_1_900 = '-2.68750e-13*ic_cap*ic_cap+-1.75000e-13*ic_cap+5.60000e-11'
+ mcrdlm5d_cc_w_1_600_s_2_000 = '-2.31250e-13*ic_cap*ic_cap+-1.75000e-13*ic_cap+5.32000e-11'
+ mcrdlm5d_cc_w_1_600_s_2_400 = '-1.37500e-13*ic_cap*ic_cap+-1.25000e-13*ic_cap+4.42000e-11'
+ mcrdlm5d_cc_w_1_600_s_2_800 = '-8.75000e-14*ic_cap*ic_cap+-7.50000e-14*ic_cap+3.77000e-11'
+ mcrdlm5d_cc_w_1_600_s_3_200 = '-4.68750e-14*ic_cap*ic_cap+-3.75000e-14*ic_cap+3.25000e-11'
+ mcrdlm5d_cc_w_1_600_s_4_800 = '2.81250e-14*ic_cap*ic_cap+1.25000e-14*ic_cap+1.94000e-11'
+ mcrdlm5d_cc_w_4_000_s_10_000 = '6.71875e-14*ic_cap*ic_cap+4.12500e-14*ic_cap+4.75000e-12'
+ mcrdlm5d_cc_w_4_000_s_12_000 = '5.21875e-14*ic_cap*ic_cap+3.87500e-14*ic_cap+2.79000e-12'
+ mcrdlm5d_cc_w_4_000_s_1_600 = '-3.43750e-13*ic_cap*ic_cap+-2.25000e-13*ic_cap+6.93000e-11'
+ mcrdlm5d_cc_w_4_000_s_1_700 = '-2.96875e-13*ic_cap*ic_cap+-2.12500e-13*ic_cap+6.54000e-11'
+ mcrdlm5d_cc_w_4_000_s_1_900 = '-2.18750e-13*ic_cap*ic_cap+-1.50000e-13*ic_cap+5.86000e-11'
+ mcrdlm5d_cc_w_4_000_s_2_000 = '-1.90625e-13*ic_cap*ic_cap+-1.37500e-13*ic_cap+5.57000e-11'
+ mcrdlm5d_cc_w_4_000_s_2_400 = '-1.00000e-13*ic_cap*ic_cap+-7.50000e-14*ic_cap+4.63000e-11'
+ mcrdlm5d_cc_w_4_000_s_2_800 = '-5.31250e-14*ic_cap*ic_cap+-3.75000e-14*ic_cap+3.94000e-11'
+ mcrdlm5d_cc_w_4_000_s_3_200 = '-1.25000e-14*ic_cap*ic_cap+-2.50000e-14*ic_cap+3.40000e-11'
+ mcrdlm5d_cc_w_4_000_s_4_800 = '5.93750e-14*ic_cap*ic_cap+3.75000e-14*ic_cap+2.03000e-11'
+ mcrdlm5d_cf_w_1_600_s_10_000 = '-2.18750e-13*ic_cap*ic_cap+-1.50000e-13*ic_cap+3.49000e-11'
+ mcrdlm5d_cf_w_1_600_s_12_000 = '-2.09375e-13*ic_cap*ic_cap+-1.37500e-13*ic_cap+3.66000e-11'
+ mcrdlm5d_cf_w_1_600_s_1_600 = '-5.84375e-14*ic_cap*ic_cap+-3.37500e-14*ic_cap+9.43000e-12'
+ mcrdlm5d_cf_w_1_600_s_1_700 = '-6.28125e-14*ic_cap*ic_cap+-3.62500e-14*ic_cap+9.98000e-12'
+ mcrdlm5d_cf_w_1_600_s_1_900 = '-7.43750e-14*ic_cap*ic_cap+-4.75000e-14*ic_cap+1.11000e-11'
+ mcrdlm5d_cf_w_1_600_s_2_000 = '-7.81250e-14*ic_cap*ic_cap+-3.75000e-14*ic_cap+1.16000e-11'
+ mcrdlm5d_cf_w_1_600_s_2_400 = '-9.68750e-14*ic_cap*ic_cap+-6.25000e-14*ic_cap+1.37000e-11'
+ mcrdlm5d_cf_w_1_600_s_2_800 = '-1.15625e-13*ic_cap*ic_cap+-6.25000e-14*ic_cap+1.57000e-11'
+ mcrdlm5d_cf_w_1_600_s_3_200 = '-1.34375e-13*ic_cap*ic_cap+-8.75000e-14*ic_cap+1.76000e-11'
+ mcrdlm5d_cf_w_1_600_s_4_800 = '-1.84375e-13*ic_cap*ic_cap+-1.12500e-13*ic_cap+2.40000e-11'
+ mcrdlm5d_cf_w_4_000_s_10_000 = '-2.09375e-13*ic_cap*ic_cap+-1.37500e-13*ic_cap+3.55000e-11'
+ mcrdlm5d_cf_w_4_000_s_12_000 = '-2.00000e-13*ic_cap*ic_cap+-1.25000e-13*ic_cap+3.73000e-11'
+ mcrdlm5d_cf_w_4_000_s_1_600 = '-5.75000e-14*ic_cap*ic_cap+-3.50000e-14*ic_cap+9.42000e-12'
+ mcrdlm5d_cf_w_4_000_s_1_700 = '-6.25000e-14*ic_cap*ic_cap+-3.75000e-14*ic_cap+9.98000e-12'
+ mcrdlm5d_cf_w_4_000_s_1_900 = '-7.37500e-14*ic_cap*ic_cap+-4.50000e-14*ic_cap+1.11000e-11'
+ mcrdlm5d_cf_w_4_000_s_2_000 = '-7.50000e-14*ic_cap*ic_cap+-5.00000e-14*ic_cap+1.16000e-11'
+ mcrdlm5d_cf_w_4_000_s_2_400 = '-9.68750e-14*ic_cap*ic_cap+-6.25000e-14*ic_cap+1.37000e-11'
+ mcrdlm5d_cf_w_4_000_s_2_800 = '-1.12500e-13*ic_cap*ic_cap+-7.50000e-14*ic_cap+1.57000e-11'
+ mcrdlm5d_cf_w_4_000_s_3_200 = '-1.28125e-13*ic_cap*ic_cap+-8.75000e-14*ic_cap+1.76000e-11'
+ mcrdlm5d_cf_w_4_000_s_4_800 = '-1.78125e-13*ic_cap*ic_cap+-1.12500e-13*ic_cap+2.41000e-11'
+ mcrdlm5f_ca_w_1_600_s_10_000 = '-1.16875e-07*ic_cap*ic_cap+-6.75000e-08*ic_cap+1.20000e-05'
+ mcrdlm5f_ca_w_1_600_s_12_000 = '-1.16875e-07*ic_cap*ic_cap+-6.75000e-08*ic_cap+1.20000e-05'
+ mcrdlm5f_ca_w_1_600_s_1_600 = '-1.16875e-07*ic_cap*ic_cap+-6.75000e-08*ic_cap+1.20000e-05'
+ mcrdlm5f_ca_w_1_600_s_1_700 = '-1.16875e-07*ic_cap*ic_cap+-6.75000e-08*ic_cap+1.20000e-05'
+ mcrdlm5f_ca_w_1_600_s_1_900 = '-1.16875e-07*ic_cap*ic_cap+-6.75000e-08*ic_cap+1.20000e-05'
+ mcrdlm5f_ca_w_1_600_s_2_000 = '-1.16875e-07*ic_cap*ic_cap+-6.75000e-08*ic_cap+1.20000e-05'
+ mcrdlm5f_ca_w_1_600_s_2_400 = '-1.16875e-07*ic_cap*ic_cap+-6.75000e-08*ic_cap+1.20000e-05'
+ mcrdlm5f_ca_w_1_600_s_2_800 = '-1.16875e-07*ic_cap*ic_cap+-6.75000e-08*ic_cap+1.20000e-05'
+ mcrdlm5f_ca_w_1_600_s_3_200 = '-1.16875e-07*ic_cap*ic_cap+-6.75000e-08*ic_cap+1.20000e-05'
+ mcrdlm5f_ca_w_1_600_s_4_800 = '-1.16875e-07*ic_cap*ic_cap+-6.75000e-08*ic_cap+1.20000e-05'
+ mcrdlm5f_ca_w_4_000_s_10_000 = '-1.16875e-07*ic_cap*ic_cap+-6.75000e-08*ic_cap+1.20000e-05'
+ mcrdlm5f_ca_w_4_000_s_12_000 = '-1.16875e-07*ic_cap*ic_cap+-6.75000e-08*ic_cap+1.20000e-05'
+ mcrdlm5f_ca_w_4_000_s_1_600 = '-1.16875e-07*ic_cap*ic_cap+-6.75000e-08*ic_cap+1.20000e-05'
+ mcrdlm5f_ca_w_4_000_s_1_700 = '-1.16875e-07*ic_cap*ic_cap+-6.75000e-08*ic_cap+1.20000e-05'
+ mcrdlm5f_ca_w_4_000_s_1_900 = '-1.16875e-07*ic_cap*ic_cap+-6.75000e-08*ic_cap+1.20000e-05'
+ mcrdlm5f_ca_w_4_000_s_2_000 = '-1.16875e-07*ic_cap*ic_cap+-6.75000e-08*ic_cap+1.20000e-05'
+ mcrdlm5f_ca_w_4_000_s_2_400 = '-1.16875e-07*ic_cap*ic_cap+-6.75000e-08*ic_cap+1.20000e-05'
+ mcrdlm5f_ca_w_4_000_s_2_800 = '-1.16875e-07*ic_cap*ic_cap+-6.75000e-08*ic_cap+1.20000e-05'
+ mcrdlm5f_ca_w_4_000_s_3_200 = '-1.16875e-07*ic_cap*ic_cap+-6.75000e-08*ic_cap+1.20000e-05'
+ mcrdlm5f_ca_w_4_000_s_4_800 = '-1.16875e-07*ic_cap*ic_cap+-6.75000e-08*ic_cap+1.20000e-05'
+ mcrdlm5f_cc_w_1_600_s_10_000 = '5.84375e-14*ic_cap*ic_cap+3.87500e-14*ic_cap+4.80000e-12'
+ mcrdlm5f_cc_w_1_600_s_12_000 = '4.87500e-14*ic_cap*ic_cap+3.25000e-14*ic_cap+2.83000e-12'
+ mcrdlm5f_cc_w_1_600_s_1_600 = '-4.00000e-13*ic_cap*ic_cap+-2.75000e-13*ic_cap+6.69000e-11'
+ mcrdlm5f_cc_w_1_600_s_1_700 = '-3.50000e-13*ic_cap*ic_cap+-2.50000e-13*ic_cap+6.30000e-11'
+ mcrdlm5f_cc_w_1_600_s_1_900 = '-2.71875e-13*ic_cap*ic_cap+-1.87500e-13*ic_cap+5.65000e-11'
+ mcrdlm5f_cc_w_1_600_s_2_000 = '-2.37500e-13*ic_cap*ic_cap+-1.75000e-13*ic_cap+5.37000e-11'
+ mcrdlm5f_cc_w_1_600_s_2_400 = '-1.43750e-13*ic_cap*ic_cap+-1.00000e-13*ic_cap+4.48000e-11'
+ mcrdlm5f_cc_w_1_600_s_2_800 = '-8.75000e-14*ic_cap*ic_cap+-7.50000e-14*ic_cap+3.82000e-11'
+ mcrdlm5f_cc_w_1_600_s_3_200 = '-4.68750e-14*ic_cap*ic_cap+-3.75000e-14*ic_cap+3.30000e-11'
+ mcrdlm5f_cc_w_1_600_s_4_800 = '2.81250e-14*ic_cap*ic_cap+1.25000e-14*ic_cap+1.99000e-11'
+ mcrdlm5f_cc_w_4_000_s_10_000 = '7.12500e-14*ic_cap*ic_cap+4.75000e-14*ic_cap+5.08000e-12'
+ mcrdlm5f_cc_w_4_000_s_12_000 = '5.65625e-14*ic_cap*ic_cap+3.87500e-14*ic_cap+3.03000e-12'
+ mcrdlm5f_cc_w_4_000_s_1_600 = '-3.43750e-13*ic_cap*ic_cap+-2.25000e-13*ic_cap+6.99000e-11'
+ mcrdlm5f_cc_w_4_000_s_1_700 = '-2.87500e-13*ic_cap*ic_cap+-2.00000e-13*ic_cap+6.59000e-11'
+ mcrdlm5f_cc_w_4_000_s_1_900 = '-2.09375e-13*ic_cap*ic_cap+-1.37500e-13*ic_cap+5.91000e-11'
+ mcrdlm5f_cc_w_4_000_s_2_000 = '-1.81250e-13*ic_cap*ic_cap+-1.25000e-13*ic_cap+5.62000e-11'
+ mcrdlm5f_cc_w_4_000_s_2_400 = '-9.68750e-14*ic_cap*ic_cap+-8.75000e-14*ic_cap+4.69000e-11'
+ mcrdlm5f_cc_w_4_000_s_2_800 = '-4.68750e-14*ic_cap*ic_cap+-3.75000e-14*ic_cap+4.00000e-11'
+ mcrdlm5f_cc_w_4_000_s_3_200 = '-1.56250e-14*ic_cap*ic_cap+-1.25000e-14*ic_cap+3.47000e-11'
+ mcrdlm5f_cc_w_4_000_s_4_800 = '5.62500e-14*ic_cap*ic_cap+2.50000e-14*ic_cap+2.09000e-11'
+ mcrdlm5f_cf_w_1_600_s_10_000 = '-2.21875e-13*ic_cap*ic_cap+-1.37500e-13*ic_cap+3.43000e-11'
+ mcrdlm5f_cf_w_1_600_s_12_000 = '-2.21875e-13*ic_cap*ic_cap+-1.37500e-13*ic_cap+3.61000e-11'
+ mcrdlm5f_cf_w_1_600_s_1_600 = '-5.87500e-14*ic_cap*ic_cap+-3.50000e-14*ic_cap+9.13000e-12'
+ mcrdlm5f_cf_w_1_600_s_1_700 = '-6.43750e-14*ic_cap*ic_cap+-3.75000e-14*ic_cap+9.67000e-12'
+ mcrdlm5f_cf_w_1_600_s_1_900 = '-7.28125e-14*ic_cap*ic_cap+-4.37500e-14*ic_cap+1.07000e-11'
+ mcrdlm5f_cf_w_1_600_s_2_000 = '-7.56250e-14*ic_cap*ic_cap+-5.25000e-14*ic_cap+1.12000e-11'
+ mcrdlm5f_cf_w_1_600_s_2_400 = '-1.00000e-13*ic_cap*ic_cap+-5.00000e-14*ic_cap+1.33000e-11'
+ mcrdlm5f_cf_w_1_600_s_2_800 = '-1.15625e-13*ic_cap*ic_cap+-6.25000e-14*ic_cap+1.52000e-11'
+ mcrdlm5f_cf_w_1_600_s_3_200 = '-1.31250e-13*ic_cap*ic_cap+-7.50000e-14*ic_cap+1.70000e-11'
+ mcrdlm5f_cf_w_1_600_s_4_800 = '-1.78125e-13*ic_cap*ic_cap+-1.12500e-13*ic_cap+2.33000e-11'
+ mcrdlm5f_cf_w_4_000_s_10_000 = '-2.15625e-13*ic_cap*ic_cap+-1.37500e-13*ic_cap+3.49000e-11'
+ mcrdlm5f_cf_w_4_000_s_12_000 = '-2.09375e-13*ic_cap*ic_cap+-1.37500e-13*ic_cap+3.68000e-11'
+ mcrdlm5f_cf_w_4_000_s_1_600 = '-5.87500e-14*ic_cap*ic_cap+-3.50000e-14*ic_cap+9.13000e-12'
+ mcrdlm5f_cf_w_4_000_s_1_700 = '-6.37500e-14*ic_cap*ic_cap+-3.75000e-14*ic_cap+9.67000e-12'
+ mcrdlm5f_cf_w_4_000_s_1_900 = '-7.18750e-14*ic_cap*ic_cap+-4.50000e-14*ic_cap+1.07000e-11'
+ mcrdlm5f_cf_w_4_000_s_2_000 = '-8.06250e-14*ic_cap*ic_cap+-4.75000e-14*ic_cap+1.13000e-11'
+ mcrdlm5f_cf_w_4_000_s_2_400 = '-9.68750e-14*ic_cap*ic_cap+-6.25000e-14*ic_cap+1.33000e-11'
+ mcrdlm5f_cf_w_4_000_s_2_800 = '-1.12500e-13*ic_cap*ic_cap+-7.50000e-14*ic_cap+1.52000e-11'
+ mcrdlm5f_cf_w_4_000_s_3_200 = '-1.31250e-13*ic_cap*ic_cap+-7.50000e-14*ic_cap+1.71000e-11'
+ mcrdlm5f_cf_w_4_000_s_4_800 = '-1.78125e-13*ic_cap*ic_cap+-1.12500e-13*ic_cap+2.35000e-11'
+ mcrdlm5l1_ca_w_1_600_s_10_000 = '-1.18750e-07*ic_cap*ic_cap+-7.50000e-08*ic_cap+1.35000e-05'
+ mcrdlm5l1_ca_w_1_600_s_12_000 = '-1.18750e-07*ic_cap*ic_cap+-7.50000e-08*ic_cap+1.35000e-05'
+ mcrdlm5l1_ca_w_1_600_s_1_600 = '-1.18750e-07*ic_cap*ic_cap+-7.50000e-08*ic_cap+1.35000e-05'
+ mcrdlm5l1_ca_w_1_600_s_1_700 = '-1.18750e-07*ic_cap*ic_cap+-7.50000e-08*ic_cap+1.35000e-05'
+ mcrdlm5l1_ca_w_1_600_s_1_900 = '-1.18750e-07*ic_cap*ic_cap+-7.50000e-08*ic_cap+1.35000e-05'
+ mcrdlm5l1_ca_w_1_600_s_2_000 = '-1.18750e-07*ic_cap*ic_cap+-7.50000e-08*ic_cap+1.35000e-05'
+ mcrdlm5l1_ca_w_1_600_s_2_400 = '-1.18750e-07*ic_cap*ic_cap+-7.50000e-08*ic_cap+1.35000e-05'
+ mcrdlm5l1_ca_w_1_600_s_2_800 = '-1.18750e-07*ic_cap*ic_cap+-7.50000e-08*ic_cap+1.35000e-05'
+ mcrdlm5l1_ca_w_1_600_s_3_200 = '-1.18750e-07*ic_cap*ic_cap+-7.50000e-08*ic_cap+1.35000e-05'
+ mcrdlm5l1_ca_w_1_600_s_4_800 = '-1.18750e-07*ic_cap*ic_cap+-7.50000e-08*ic_cap+1.35000e-05'
+ mcrdlm5l1_ca_w_4_000_s_10_000 = '-1.18750e-07*ic_cap*ic_cap+-7.50000e-08*ic_cap+1.35000e-05'
+ mcrdlm5l1_ca_w_4_000_s_12_000 = '-1.18750e-07*ic_cap*ic_cap+-7.50000e-08*ic_cap+1.35000e-05'
+ mcrdlm5l1_ca_w_4_000_s_1_600 = '-1.18750e-07*ic_cap*ic_cap+-7.50000e-08*ic_cap+1.35000e-05'
+ mcrdlm5l1_ca_w_4_000_s_1_700 = '-1.18750e-07*ic_cap*ic_cap+-7.50000e-08*ic_cap+1.35000e-05'
+ mcrdlm5l1_ca_w_4_000_s_1_900 = '-1.18750e-07*ic_cap*ic_cap+-7.50000e-08*ic_cap+1.35000e-05'
+ mcrdlm5l1_ca_w_4_000_s_2_000 = '-1.18750e-07*ic_cap*ic_cap+-7.50000e-08*ic_cap+1.35000e-05'
+ mcrdlm5l1_ca_w_4_000_s_2_400 = '-1.18750e-07*ic_cap*ic_cap+-7.50000e-08*ic_cap+1.35000e-05'
+ mcrdlm5l1_ca_w_4_000_s_2_800 = '-1.18750e-07*ic_cap*ic_cap+-7.50000e-08*ic_cap+1.35000e-05'
+ mcrdlm5l1_ca_w_4_000_s_3_200 = '-1.18750e-07*ic_cap*ic_cap+-7.50000e-08*ic_cap+1.35000e-05'
+ mcrdlm5l1_ca_w_4_000_s_4_800 = '-1.18750e-07*ic_cap*ic_cap+-7.50000e-08*ic_cap+1.35000e-05'
+ mcrdlm5l1_cc_w_1_600_s_10_000 = '5.15625e-14*ic_cap*ic_cap+3.12500e-14*ic_cap+3.79000e-12'
+ mcrdlm5l1_cc_w_1_600_s_12_000 = '3.81250e-14*ic_cap*ic_cap+2.50000e-14*ic_cap+2.14000e-12'
+ mcrdlm5l1_cc_w_1_600_s_1_600 = '-3.90625e-13*ic_cap*ic_cap+-2.87500e-13*ic_cap+6.52000e-11'
+ mcrdlm5l1_cc_w_1_600_s_1_700 = '-3.40625e-13*ic_cap*ic_cap+-2.37500e-13*ic_cap+6.13000e-11'
+ mcrdlm5l1_cc_w_1_600_s_1_900 = '-2.71875e-13*ic_cap*ic_cap+-1.87500e-13*ic_cap+5.49000e-11'
+ mcrdlm5l1_cc_w_1_600_s_2_000 = '-2.37500e-13*ic_cap*ic_cap+-1.75000e-13*ic_cap+5.21000e-11'
+ mcrdlm5l1_cc_w_1_600_s_2_400 = '-1.43750e-13*ic_cap*ic_cap+-1.00000e-13*ic_cap+4.30000e-11'
+ mcrdlm5l1_cc_w_1_600_s_2_800 = '-8.43750e-14*ic_cap*ic_cap+-6.25000e-14*ic_cap+3.64000e-11'
+ mcrdlm5l1_cc_w_1_600_s_3_200 = '-4.68750e-14*ic_cap*ic_cap+-3.75000e-14*ic_cap+3.12000e-11'
+ mcrdlm5l1_cc_w_1_600_s_4_800 = '3.12500e-14*ic_cap*ic_cap+1.81000e-11'
+ mcrdlm5l1_cc_w_4_000_s_10_000 = '5.93750e-14*ic_cap*ic_cap+3.50000e-14*ic_cap+4.01000e-12'
+ mcrdlm5l1_cc_w_4_000_s_12_000 = '4.31250e-14*ic_cap*ic_cap+3.50000e-14*ic_cap+2.28000e-12'
+ mcrdlm5l1_cc_w_4_000_s_1_600 = '-3.34375e-13*ic_cap*ic_cap+-2.12500e-13*ic_cap+6.77000e-11'
+ mcrdlm5l1_cc_w_4_000_s_1_700 = '-2.90625e-13*ic_cap*ic_cap+-1.87500e-13*ic_cap+6.37000e-11'
+ mcrdlm5l1_cc_w_4_000_s_1_900 = '-2.15625e-13*ic_cap*ic_cap+-1.62500e-13*ic_cap+5.70000e-11'
+ mcrdlm5l1_cc_w_4_000_s_2_000 = '-1.87500e-13*ic_cap*ic_cap+-1.25000e-13*ic_cap+5.41000e-11'
+ mcrdlm5l1_cc_w_4_000_s_2_400 = '-1.06250e-13*ic_cap*ic_cap+-7.50000e-14*ic_cap+4.48000e-11'
+ mcrdlm5l1_cc_w_4_000_s_2_800 = '-4.06250e-14*ic_cap*ic_cap+-3.75000e-14*ic_cap+3.78000e-11'
+ mcrdlm5l1_cc_w_4_000_s_3_200 = '-1.56250e-14*ic_cap*ic_cap+-1.25000e-14*ic_cap+3.25000e-11'
+ mcrdlm5l1_cc_w_4_000_s_4_800 = '5.31250e-14*ic_cap*ic_cap+3.75000e-14*ic_cap+1.89000e-11'
+ mcrdlm5l1_cf_w_1_600_s_10_000 = '-2.21875e-13*ic_cap*ic_cap+-1.37500e-13*ic_cap+3.66000e-11'
+ mcrdlm5l1_cf_w_1_600_s_12_000 = '-2.15625e-13*ic_cap*ic_cap+-1.37500e-13*ic_cap+3.82000e-11'
+ mcrdlm5l1_cf_w_1_600_s_1_600 = '-6.21875e-14*ic_cap*ic_cap+-3.62500e-14*ic_cap+1.03000e-11'
+ mcrdlm5l1_cf_w_1_600_s_1_700 = '-6.71875e-14*ic_cap*ic_cap+-4.12500e-14*ic_cap+1.09000e-11'
+ mcrdlm5l1_cf_w_1_600_s_1_900 = '-7.50000e-14*ic_cap*ic_cap+-5.00000e-14*ic_cap+1.20000e-11'
+ mcrdlm5l1_cf_w_1_600_s_2_000 = '-8.12500e-14*ic_cap*ic_cap+-5.00000e-14*ic_cap+1.26000e-11'
+ mcrdlm5l1_cf_w_1_600_s_2_400 = '-1.03125e-13*ic_cap*ic_cap+-6.25000e-14*ic_cap+1.49000e-11'
+ mcrdlm5l1_cf_w_1_600_s_2_800 = '-1.18750e-13*ic_cap*ic_cap+-7.50000e-14*ic_cap+1.70000e-11'
+ mcrdlm5l1_cf_w_1_600_s_3_200 = '-1.34375e-13*ic_cap*ic_cap+-8.75000e-14*ic_cap+1.90000e-11'
+ mcrdlm5l1_cf_w_1_600_s_4_800 = '-1.90625e-13*ic_cap*ic_cap+-1.12500e-13*ic_cap+2.58000e-11'
+ mcrdlm5l1_cf_w_4_000_s_10_000 = '-2.09375e-13*ic_cap*ic_cap+-1.37500e-13*ic_cap+3.72000e-11'
+ mcrdlm5l1_cf_w_4_000_s_12_000 = '-2.03125e-13*ic_cap*ic_cap+-1.37500e-13*ic_cap+3.89000e-11'
+ mcrdlm5l1_cf_w_4_000_s_1_600 = '-6.21875e-14*ic_cap*ic_cap+-3.62500e-14*ic_cap+1.03000e-11'
+ mcrdlm5l1_cf_w_4_000_s_1_700 = '-6.75000e-14*ic_cap*ic_cap+-4.00000e-14*ic_cap+1.09000e-11'
+ mcrdlm5l1_cf_w_4_000_s_1_900 = '-7.81250e-14*ic_cap*ic_cap+-3.75000e-14*ic_cap+1.21000e-11'
+ mcrdlm5l1_cf_w_4_000_s_2_000 = '-8.12500e-14*ic_cap*ic_cap+-5.00000e-14*ic_cap+1.26000e-11'
+ mcrdlm5l1_cf_w_4_000_s_2_400 = '-1.03125e-13*ic_cap*ic_cap+-6.25000e-14*ic_cap+1.49000e-11'
+ mcrdlm5l1_cf_w_4_000_s_2_800 = '-1.18750e-13*ic_cap*ic_cap+-7.50000e-14*ic_cap+1.70000e-11'
+ mcrdlm5l1_cf_w_4_000_s_3_200 = '-1.37500e-13*ic_cap*ic_cap+-7.50000e-14*ic_cap+1.91000e-11'
+ mcrdlm5l1_cf_w_4_000_s_4_800 = '-1.81250e-13*ic_cap*ic_cap+-1.25000e-13*ic_cap+2.59000e-11'
+ mcrdlm5m1_ca_w_1_600_s_10_000 = '-1.31250e-07*ic_cap*ic_cap+-7.50000e-08*ic_cap+1.50000e-05'
+ mcrdlm5m1_ca_w_1_600_s_12_000 = '-1.31250e-07*ic_cap*ic_cap+-7.50000e-08*ic_cap+1.50000e-05'
+ mcrdlm5m1_ca_w_1_600_s_1_600 = '-1.31250e-07*ic_cap*ic_cap+-7.50000e-08*ic_cap+1.50000e-05'
+ mcrdlm5m1_ca_w_1_600_s_1_700 = '-1.31250e-07*ic_cap*ic_cap+-7.50000e-08*ic_cap+1.50000e-05'
+ mcrdlm5m1_ca_w_1_600_s_1_900 = '-1.31250e-07*ic_cap*ic_cap+-7.50000e-08*ic_cap+1.50000e-05'
+ mcrdlm5m1_ca_w_1_600_s_2_000 = '-1.31250e-07*ic_cap*ic_cap+-7.50000e-08*ic_cap+1.50000e-05'
+ mcrdlm5m1_ca_w_1_600_s_2_400 = '-1.31250e-07*ic_cap*ic_cap+-7.50000e-08*ic_cap+1.50000e-05'
+ mcrdlm5m1_ca_w_1_600_s_2_800 = '-1.31250e-07*ic_cap*ic_cap+-7.50000e-08*ic_cap+1.50000e-05'
+ mcrdlm5m1_ca_w_1_600_s_3_200 = '-1.31250e-07*ic_cap*ic_cap+-7.50000e-08*ic_cap+1.50000e-05'
+ mcrdlm5m1_ca_w_1_600_s_4_800 = '-1.31250e-07*ic_cap*ic_cap+-7.50000e-08*ic_cap+1.50000e-05'
+ mcrdlm5m1_ca_w_4_000_s_10_000 = '-1.31250e-07*ic_cap*ic_cap+-7.50000e-08*ic_cap+1.50000e-05'
+ mcrdlm5m1_ca_w_4_000_s_12_000 = '-1.31250e-07*ic_cap*ic_cap+-7.50000e-08*ic_cap+1.50000e-05'
+ mcrdlm5m1_ca_w_4_000_s_1_600 = '-1.31250e-07*ic_cap*ic_cap+-7.50000e-08*ic_cap+1.50000e-05'
+ mcrdlm5m1_ca_w_4_000_s_1_700 = '-1.31250e-07*ic_cap*ic_cap+-7.50000e-08*ic_cap+1.50000e-05'
+ mcrdlm5m1_ca_w_4_000_s_1_900 = '-1.31250e-07*ic_cap*ic_cap+-7.50000e-08*ic_cap+1.50000e-05'
+ mcrdlm5m1_ca_w_4_000_s_2_000 = '-1.31250e-07*ic_cap*ic_cap+-7.50000e-08*ic_cap+1.50000e-05'
+ mcrdlm5m1_ca_w_4_000_s_2_400 = '-1.31250e-07*ic_cap*ic_cap+-7.50000e-08*ic_cap+1.50000e-05'
+ mcrdlm5m1_ca_w_4_000_s_2_800 = '-1.31250e-07*ic_cap*ic_cap+-7.50000e-08*ic_cap+1.50000e-05'
+ mcrdlm5m1_ca_w_4_000_s_3_200 = '-1.31250e-07*ic_cap*ic_cap+-7.50000e-08*ic_cap+1.50000e-05'
+ mcrdlm5m1_ca_w_4_000_s_4_800 = '-1.31250e-07*ic_cap*ic_cap+-7.50000e-08*ic_cap+1.50000e-05'
+ mcrdlm5m1_cc_w_1_600_s_10_000 = '4.68750e-14*ic_cap*ic_cap+2.75000e-14*ic_cap+3.12000e-12'
+ mcrdlm5m1_cc_w_1_600_s_12_000 = '3.46875e-14*ic_cap*ic_cap+2.12500e-14*ic_cap+1.66000e-12'
+ mcrdlm5m1_cc_w_1_600_s_1_600 = '-3.90625e-13*ic_cap*ic_cap+-2.87500e-13*ic_cap+6.39000e-11'
+ mcrdlm5m1_cc_w_1_600_s_1_700 = '-3.40625e-13*ic_cap*ic_cap+-2.37500e-13*ic_cap+5.99000e-11'
+ mcrdlm5m1_cc_w_1_600_s_1_900 = '-2.68750e-13*ic_cap*ic_cap+-1.75000e-13*ic_cap+5.35000e-11'
+ mcrdlm5m1_cc_w_1_600_s_2_000 = '-2.31250e-13*ic_cap*ic_cap+-1.75000e-13*ic_cap+5.06000e-11'
+ mcrdlm5m1_cc_w_1_600_s_2_400 = '-1.34375e-13*ic_cap*ic_cap+-8.75000e-14*ic_cap+4.15000e-11'
+ mcrdlm5m1_cc_w_1_600_s_2_800 = '-8.12500e-14*ic_cap*ic_cap+-7.50000e-14*ic_cap+3.49000e-11'
+ mcrdlm5m1_cc_w_1_600_s_3_200 = '-4.68750e-14*ic_cap*ic_cap+-3.75000e-14*ic_cap+2.97000e-11'
+ mcrdlm5m1_cc_w_1_600_s_4_800 = '3.12500e-14*ic_cap*ic_cap+2.50000e-14*ic_cap+1.67000e-11'
+ mcrdlm5m1_cc_w_4_000_s_10_000 = '5.25000e-14*ic_cap*ic_cap+3.75000e-14*ic_cap+3.30000e-12'
+ mcrdlm5m1_cc_w_4_000_s_12_000 = '3.87500e-14*ic_cap*ic_cap+2.50000e-14*ic_cap+1.76000e-12'
+ mcrdlm5m1_cc_w_4_000_s_1_600 = '-3.34375e-13*ic_cap*ic_cap+-2.12500e-13*ic_cap+6.60000e-11'
+ mcrdlm5m1_cc_w_4_000_s_1_700 = '-2.93750e-13*ic_cap*ic_cap+-2.00000e-13*ic_cap+6.21000e-11'
+ mcrdlm5m1_cc_w_4_000_s_1_900 = '-2.18750e-13*ic_cap*ic_cap+-1.50000e-13*ic_cap+5.53000e-11'
+ mcrdlm5m1_cc_w_4_000_s_2_000 = '-1.87500e-13*ic_cap*ic_cap+-1.50000e-13*ic_cap+5.24000e-11'
+ mcrdlm5m1_cc_w_4_000_s_2_400 = '-1.09375e-13*ic_cap*ic_cap+-8.75000e-14*ic_cap+4.32000e-11'
+ mcrdlm5m1_cc_w_4_000_s_2_800 = '-4.37500e-14*ic_cap*ic_cap+-2.50000e-14*ic_cap+3.61000e-11'
+ mcrdlm5m1_cc_w_4_000_s_3_200 = '-9.37500e-15*ic_cap*ic_cap+-1.25000e-14*ic_cap+3.07000e-11'
+ mcrdlm5m1_cc_w_4_000_s_4_800 = '5.00000e-14*ic_cap*ic_cap+2.50000e-14*ic_cap+1.74000e-11'
+ mcrdlm5m1_cf_w_1_600_s_10_000 = '-2.18750e-13*ic_cap*ic_cap+-1.50000e-13*ic_cap+3.85000e-11'
+ mcrdlm5m1_cf_w_1_600_s_12_000 = '-2.18750e-13*ic_cap*ic_cap+-1.50000e-13*ic_cap+4.00000e-11'
+ mcrdlm5m1_cf_w_1_600_s_1_600 = '-5.93750e-14*ic_cap*ic_cap+-3.75000e-14*ic_cap+1.13000e-11'
+ mcrdlm5m1_cf_w_1_600_s_1_700 = '-7.18750e-14*ic_cap*ic_cap+-3.75000e-14*ic_cap+1.20000e-11'
+ mcrdlm5m1_cf_w_1_600_s_1_900 = '-8.12500e-14*ic_cap*ic_cap+-5.00000e-14*ic_cap+1.33000e-11'
+ mcrdlm5m1_cf_w_1_600_s_2_000 = '-8.75000e-14*ic_cap*ic_cap+-5.00000e-14*ic_cap+1.39000e-11'
+ mcrdlm5m1_cf_w_1_600_s_2_400 = '-1.03125e-13*ic_cap*ic_cap+-6.25000e-14*ic_cap+1.63000e-11'
+ mcrdlm5m1_cf_w_1_600_s_2_800 = '-1.25000e-13*ic_cap*ic_cap+-7.50000e-14*ic_cap+1.86000e-11'
+ mcrdlm5m1_cf_w_1_600_s_3_200 = '-1.46875e-13*ic_cap*ic_cap+-8.75000e-14*ic_cap+2.08000e-11'
+ mcrdlm5m1_cf_w_1_600_s_4_800 = '-1.96875e-13*ic_cap*ic_cap+-1.12500e-13*ic_cap+2.79000e-11'
+ mcrdlm5m1_cf_w_4_000_s_10_000 = '-2.12500e-13*ic_cap*ic_cap+-1.25000e-13*ic_cap+3.91000e-11'
+ mcrdlm5m1_cf_w_4_000_s_12_000 = '-2.03125e-13*ic_cap*ic_cap+-1.37500e-13*ic_cap+4.06000e-11'
+ mcrdlm5m1_cf_w_4_000_s_1_600 = '-5.93750e-14*ic_cap*ic_cap+-3.75000e-14*ic_cap+1.13000e-11'
+ mcrdlm5m1_cf_w_4_000_s_1_700 = '-7.18750e-14*ic_cap*ic_cap+-3.75000e-14*ic_cap+1.20000e-11'
+ mcrdlm5m1_cf_w_4_000_s_1_900 = '-8.12500e-14*ic_cap*ic_cap+-5.00000e-14*ic_cap+1.33000e-11'
+ mcrdlm5m1_cf_w_4_000_s_2_000 = '-8.75000e-14*ic_cap*ic_cap+-5.00000e-14*ic_cap+1.39000e-11'
+ mcrdlm5m1_cf_w_4_000_s_2_400 = '-1.09375e-13*ic_cap*ic_cap+-6.25000e-14*ic_cap+1.64000e-11'
+ mcrdlm5m1_cf_w_4_000_s_2_800 = '-1.25000e-13*ic_cap*ic_cap+-7.50000e-14*ic_cap+1.87000e-11'
+ mcrdlm5m1_cf_w_4_000_s_3_200 = '-1.46875e-13*ic_cap*ic_cap+-8.75000e-14*ic_cap+2.09000e-11'
+ mcrdlm5m1_cf_w_4_000_s_4_800 = '-1.93750e-13*ic_cap*ic_cap+-1.25000e-13*ic_cap+2.81000e-11'
+ mcrdlm5m2_ca_w_1_600_s_10_000 = '-1.40625e-07*ic_cap*ic_cap+-8.75000e-08*ic_cap+1.70000e-05'
+ mcrdlm5m2_ca_w_1_600_s_12_000 = '-1.40625e-07*ic_cap*ic_cap+-8.75000e-08*ic_cap+1.70000e-05'
+ mcrdlm5m2_ca_w_1_600_s_1_600 = '-1.40625e-07*ic_cap*ic_cap+-8.75000e-08*ic_cap+1.70000e-05'
+ mcrdlm5m2_ca_w_1_600_s_1_700 = '-1.40625e-07*ic_cap*ic_cap+-8.75000e-08*ic_cap+1.70000e-05'
+ mcrdlm5m2_ca_w_1_600_s_1_900 = '-1.40625e-07*ic_cap*ic_cap+-8.75000e-08*ic_cap+1.70000e-05'
+ mcrdlm5m2_ca_w_1_600_s_2_000 = '-1.40625e-07*ic_cap*ic_cap+-8.75000e-08*ic_cap+1.70000e-05'
+ mcrdlm5m2_ca_w_1_600_s_2_400 = '-1.40625e-07*ic_cap*ic_cap+-8.75000e-08*ic_cap+1.70000e-05'
+ mcrdlm5m2_ca_w_1_600_s_2_800 = '-1.40625e-07*ic_cap*ic_cap+-8.75000e-08*ic_cap+1.70000e-05'
+ mcrdlm5m2_ca_w_1_600_s_3_200 = '-1.40625e-07*ic_cap*ic_cap+-8.75000e-08*ic_cap+1.70000e-05'
+ mcrdlm5m2_ca_w_1_600_s_4_800 = '-1.40625e-07*ic_cap*ic_cap+-8.75000e-08*ic_cap+1.70000e-05'
+ mcrdlm5m2_ca_w_4_000_s_10_000 = '-1.40625e-07*ic_cap*ic_cap+-8.75000e-08*ic_cap+1.70000e-05'
+ mcrdlm5m2_ca_w_4_000_s_12_000 = '-1.40625e-07*ic_cap*ic_cap+-8.75000e-08*ic_cap+1.70000e-05'
+ mcrdlm5m2_ca_w_4_000_s_1_600 = '-1.40625e-07*ic_cap*ic_cap+-8.75000e-08*ic_cap+1.70000e-05'
+ mcrdlm5m2_ca_w_4_000_s_1_700 = '-1.40625e-07*ic_cap*ic_cap+-8.75000e-08*ic_cap+1.70000e-05'
+ mcrdlm5m2_ca_w_4_000_s_1_900 = '-1.40625e-07*ic_cap*ic_cap+-8.75000e-08*ic_cap+1.70000e-05'
+ mcrdlm5m2_ca_w_4_000_s_2_000 = '-1.40625e-07*ic_cap*ic_cap+-8.75000e-08*ic_cap+1.70000e-05'
+ mcrdlm5m2_ca_w_4_000_s_2_400 = '-1.40625e-07*ic_cap*ic_cap+-8.75000e-08*ic_cap+1.70000e-05'
+ mcrdlm5m2_ca_w_4_000_s_2_800 = '-1.40625e-07*ic_cap*ic_cap+-8.75000e-08*ic_cap+1.70000e-05'
+ mcrdlm5m2_ca_w_4_000_s_3_200 = '-1.40625e-07*ic_cap*ic_cap+-8.75000e-08*ic_cap+1.70000e-05'
+ mcrdlm5m2_ca_w_4_000_s_4_800 = '-1.40625e-07*ic_cap*ic_cap+-8.75000e-08*ic_cap+1.70000e-05'
+ mcrdlm5m2_cc_w_1_600_s_10_000 = '3.87500e-14*ic_cap*ic_cap+2.00000e-14*ic_cap+2.48000e-12'
+ mcrdlm5m2_cc_w_1_600_s_12_000 = '2.68750e-14*ic_cap*ic_cap+1.25000e-14*ic_cap+1.27000e-12'
+ mcrdlm5m2_cc_w_1_600_s_1_600 = '-3.93750e-13*ic_cap*ic_cap+-2.75000e-13*ic_cap+6.22000e-11'
+ mcrdlm5m2_cc_w_1_600_s_1_700 = '-3.46875e-13*ic_cap*ic_cap+-2.37500e-13*ic_cap+5.83000e-11'
+ mcrdlm5m2_cc_w_1_600_s_1_900 = '-2.62500e-13*ic_cap*ic_cap+-1.75000e-13*ic_cap+5.17000e-11'
+ mcrdlm5m2_cc_w_1_600_s_2_000 = '-2.25000e-13*ic_cap*ic_cap+-1.75000e-13*ic_cap+4.88000e-11'
+ mcrdlm5m2_cc_w_1_600_s_2_400 = '-1.34375e-13*ic_cap*ic_cap+-1.12500e-13*ic_cap+3.98000e-11'
+ mcrdlm5m2_cc_w_1_600_s_2_800 = '-7.81250e-14*ic_cap*ic_cap+-6.25000e-14*ic_cap+3.31000e-11'
+ mcrdlm5m2_cc_w_1_600_s_3_200 = '-4.37500e-14*ic_cap*ic_cap+-5.00000e-14*ic_cap+2.79000e-11'
+ mcrdlm5m2_cc_w_1_600_s_4_800 = '2.81250e-14*ic_cap*ic_cap+1.25000e-14*ic_cap+1.51000e-11'
+ mcrdlm5m2_cc_w_4_000_s_10_000 = '4.62500e-14*ic_cap*ic_cap+3.00000e-14*ic_cap+2.60000e-12'
+ mcrdlm5m2_cc_w_4_000_s_12_000 = '3.15625e-14*ic_cap*ic_cap+2.62500e-14*ic_cap+1.32000e-12'
+ mcrdlm5m2_cc_w_4_000_s_1_600 = '-3.40625e-13*ic_cap*ic_cap+-2.12500e-13*ic_cap+6.41000e-11'
+ mcrdlm5m2_cc_w_4_000_s_1_700 = '-2.93750e-13*ic_cap*ic_cap+-2.00000e-13*ic_cap+6.01000e-11'
+ mcrdlm5m2_cc_w_4_000_s_1_900 = '-2.18750e-13*ic_cap*ic_cap+-1.50000e-13*ic_cap+5.33000e-11'
+ mcrdlm5m2_cc_w_4_000_s_2_000 = '-1.84375e-13*ic_cap*ic_cap+-1.37500e-13*ic_cap+5.03000e-11'
+ mcrdlm5m2_cc_w_4_000_s_2_400 = '-1.06250e-13*ic_cap*ic_cap+-7.50000e-14*ic_cap+4.11000e-11'
+ mcrdlm5m2_cc_w_4_000_s_2_800 = '-5.31250e-14*ic_cap*ic_cap+-3.75000e-14*ic_cap+3.42000e-11'
+ mcrdlm5m2_cc_w_4_000_s_3_200 = '-1.87500e-14*ic_cap*ic_cap+-2.50000e-14*ic_cap+2.89000e-11'
+ mcrdlm5m2_cc_w_4_000_s_4_800 = '5.00000e-14*ic_cap*ic_cap+2.50000e-14*ic_cap+1.57000e-11'
+ mcrdlm5m2_cf_w_1_600_s_10_000 = '-2.21875e-13*ic_cap*ic_cap+-1.37500e-13*ic_cap+4.09000e-11'
+ mcrdlm5m2_cf_w_1_600_s_12_000 = '-2.15625e-13*ic_cap*ic_cap+-1.37500e-13*ic_cap+4.21000e-11'
+ mcrdlm5m2_cf_w_1_600_s_1_600 = '-6.56250e-14*ic_cap*ic_cap+-3.75000e-14*ic_cap+1.27000e-11'
+ mcrdlm5m2_cf_w_1_600_s_1_700 = '-7.18750e-14*ic_cap*ic_cap+-3.75000e-14*ic_cap+1.35000e-11'
+ mcrdlm5m2_cf_w_1_600_s_1_900 = '-8.12500e-14*ic_cap*ic_cap+-5.00000e-14*ic_cap+1.49000e-11'
+ mcrdlm5m2_cf_w_1_600_s_2_000 = '-8.75000e-14*ic_cap*ic_cap+-5.00000e-14*ic_cap+1.56000e-11'
+ mcrdlm5m2_cf_w_1_600_s_2_400 = '-1.12500e-13*ic_cap*ic_cap+-7.50000e-14*ic_cap+1.83000e-11'
+ mcrdlm5m2_cf_w_1_600_s_2_800 = '-1.31250e-13*ic_cap*ic_cap+-7.50000e-14*ic_cap+2.08000e-11'
+ mcrdlm5m2_cf_w_1_600_s_3_200 = '-1.46875e-13*ic_cap*ic_cap+-8.75000e-14*ic_cap+2.31000e-11'
+ mcrdlm5m2_cf_w_1_600_s_4_800 = '-2.00000e-13*ic_cap*ic_cap+-1.25000e-13*ic_cap+3.06000e-11'
+ mcrdlm5m2_cf_w_4_000_s_10_000 = '-2.09375e-13*ic_cap*ic_cap+-1.37500e-13*ic_cap+4.14000e-11'
+ mcrdlm5m2_cf_w_4_000_s_12_000 = '-2.00000e-13*ic_cap*ic_cap+-1.25000e-13*ic_cap+4.27000e-11'
+ mcrdlm5m2_cf_w_4_000_s_1_600 = '-6.56250e-14*ic_cap*ic_cap+-3.75000e-14*ic_cap+1.27000e-11'
+ mcrdlm5m2_cf_w_4_000_s_1_700 = '-7.18750e-14*ic_cap*ic_cap+-3.75000e-14*ic_cap+1.35000e-11'
+ mcrdlm5m2_cf_w_4_000_s_1_900 = '-8.12500e-14*ic_cap*ic_cap+-5.00000e-14*ic_cap+1.49000e-11'
+ mcrdlm5m2_cf_w_4_000_s_2_000 = '-8.75000e-14*ic_cap*ic_cap+-5.00000e-14*ic_cap+1.56000e-11'
+ mcrdlm5m2_cf_w_4_000_s_2_400 = '-1.09375e-13*ic_cap*ic_cap+-6.25000e-14*ic_cap+1.83000e-11'
+ mcrdlm5m2_cf_w_4_000_s_2_800 = '-1.28125e-13*ic_cap*ic_cap+-8.75000e-14*ic_cap+2.08000e-11'
+ mcrdlm5m2_cf_w_4_000_s_3_200 = '-1.50000e-13*ic_cap*ic_cap+-1.00000e-13*ic_cap+2.32000e-11'
+ mcrdlm5m2_cf_w_4_000_s_4_800 = '-1.96875e-13*ic_cap*ic_cap+-1.12500e-13*ic_cap+3.08000e-11'
+ mcrdlm5m3_ca_w_1_600_s_10_000 = '-2.34375e-07*ic_cap*ic_cap+-1.37500e-07*ic_cap+2.53000e-05'
+ mcrdlm5m3_ca_w_1_600_s_12_000 = '-2.34375e-07*ic_cap*ic_cap+-1.37500e-07*ic_cap+2.53000e-05'
+ mcrdlm5m3_ca_w_1_600_s_1_600 = '-2.34375e-07*ic_cap*ic_cap+-1.37500e-07*ic_cap+2.53000e-05'
+ mcrdlm5m3_ca_w_1_600_s_1_700 = '-2.34375e-07*ic_cap*ic_cap+-1.37500e-07*ic_cap+2.53000e-05'
+ mcrdlm5m3_ca_w_1_600_s_1_900 = '-2.34375e-07*ic_cap*ic_cap+-1.37500e-07*ic_cap+2.53000e-05'
+ mcrdlm5m3_ca_w_1_600_s_2_000 = '-2.34375e-07*ic_cap*ic_cap+-1.37500e-07*ic_cap+2.53000e-05'
+ mcrdlm5m3_ca_w_1_600_s_2_400 = '-2.34375e-07*ic_cap*ic_cap+-1.37500e-07*ic_cap+2.53000e-05'
+ mcrdlm5m3_ca_w_1_600_s_2_800 = '-2.34375e-07*ic_cap*ic_cap+-1.37500e-07*ic_cap+2.53000e-05'
+ mcrdlm5m3_ca_w_1_600_s_3_200 = '-2.34375e-07*ic_cap*ic_cap+-1.37500e-07*ic_cap+2.53000e-05'
+ mcrdlm5m3_ca_w_1_600_s_4_800 = '-2.34375e-07*ic_cap*ic_cap+-1.37500e-07*ic_cap+2.53000e-05'
+ mcrdlm5m3_ca_w_4_000_s_10_000 = '-2.34375e-07*ic_cap*ic_cap+-1.37500e-07*ic_cap+2.53000e-05'
+ mcrdlm5m3_ca_w_4_000_s_12_000 = '-2.34375e-07*ic_cap*ic_cap+-1.37500e-07*ic_cap+2.53000e-05'
+ mcrdlm5m3_ca_w_4_000_s_1_600 = '-2.34375e-07*ic_cap*ic_cap+-1.37500e-07*ic_cap+2.53000e-05'
+ mcrdlm5m3_ca_w_4_000_s_1_700 = '-2.34375e-07*ic_cap*ic_cap+-1.37500e-07*ic_cap+2.53000e-05'
+ mcrdlm5m3_ca_w_4_000_s_1_900 = '-2.34375e-07*ic_cap*ic_cap+-1.37500e-07*ic_cap+2.53000e-05'
+ mcrdlm5m3_ca_w_4_000_s_2_000 = '-2.34375e-07*ic_cap*ic_cap+-1.37500e-07*ic_cap+2.53000e-05'
+ mcrdlm5m3_ca_w_4_000_s_2_400 = '-2.34375e-07*ic_cap*ic_cap+-1.37500e-07*ic_cap+2.53000e-05'
+ mcrdlm5m3_ca_w_4_000_s_2_800 = '-2.34375e-07*ic_cap*ic_cap+-1.37500e-07*ic_cap+2.53000e-05'
+ mcrdlm5m3_ca_w_4_000_s_3_200 = '-2.34375e-07*ic_cap*ic_cap+-1.37500e-07*ic_cap+2.53000e-05'
+ mcrdlm5m3_ca_w_4_000_s_4_800 = '-2.34375e-07*ic_cap*ic_cap+-1.37500e-07*ic_cap+2.53000e-05'
+ mcrdlm5m3_cc_w_1_600_s_10_000 = '3.00000e-14*ic_cap*ic_cap+1.75000e-14*ic_cap+1.26000e-12'
+ mcrdlm5m3_cc_w_1_600_s_12_000 = '1.81250e-14*ic_cap*ic_cap+1.00000e-14*ic_cap+5.70000e-13'
+ mcrdlm5m3_cc_w_1_600_s_1_600 = '-3.53125e-13*ic_cap*ic_cap+-2.37500e-13*ic_cap+5.67000e-11'
+ mcrdlm5m3_cc_w_1_600_s_1_700 = '-3.06250e-13*ic_cap*ic_cap+-2.00000e-13*ic_cap+5.28000e-11'
+ mcrdlm5m3_cc_w_1_600_s_1_900 = '-2.28125e-13*ic_cap*ic_cap+-1.62500e-13*ic_cap+4.62000e-11'
+ mcrdlm5m3_cc_w_1_600_s_2_000 = '-1.93750e-13*ic_cap*ic_cap+-1.50000e-13*ic_cap+4.34000e-11'
+ mcrdlm5m3_cc_w_1_600_s_2_400 = '-1.03125e-13*ic_cap*ic_cap+-8.75000e-14*ic_cap+3.44000e-11'
+ mcrdlm5m3_cc_w_1_600_s_2_800 = '-5.62500e-14*ic_cap*ic_cap+-5.00000e-14*ic_cap+2.79000e-11'
+ mcrdlm5m3_cc_w_1_600_s_3_200 = '-2.18750e-14*ic_cap*ic_cap+-1.25000e-14*ic_cap+2.29000e-11'
+ mcrdlm5m3_cc_w_1_600_s_4_800 = '4.06250e-14*ic_cap*ic_cap+1.25000e-14*ic_cap+1.10000e-11'
+ mcrdlm5m3_cc_w_4_000_s_10_000 = '3.46875e-14*ic_cap*ic_cap+2.37500e-14*ic_cap+1.33000e-12'
+ mcrdlm5m3_cc_w_4_000_s_12_000 = '1.96875e-14*ic_cap*ic_cap+1.00000e-14*ic_cap+6.30000e-13'
+ mcrdlm5m3_cc_w_4_000_s_1_600 = '-3.15625e-13*ic_cap*ic_cap+-2.12500e-13*ic_cap+5.82000e-11'
+ mcrdlm5m3_cc_w_4_000_s_1_700 = '-2.65625e-13*ic_cap*ic_cap+-1.87500e-13*ic_cap+5.42000e-11'
+ mcrdlm5m3_cc_w_4_000_s_1_900 = '-1.93750e-13*ic_cap*ic_cap+-1.25000e-13*ic_cap+4.75000e-11'
+ mcrdlm5m3_cc_w_4_000_s_2_000 = '-1.62500e-13*ic_cap*ic_cap+-1.25000e-13*ic_cap+4.46000e-11'
+ mcrdlm5m3_cc_w_4_000_s_2_400 = '-7.18750e-14*ic_cap*ic_cap+-6.25000e-14*ic_cap+3.53000e-11'
+ mcrdlm5m3_cc_w_4_000_s_2_800 = '-2.50000e-14*ic_cap*ic_cap+-2.50000e-14*ic_cap+2.87000e-11'
+ mcrdlm5m3_cc_w_4_000_s_3_200 = '6.25000e-15*ic_cap*ic_cap+2.36000e-11'
+ mcrdlm5m3_cc_w_4_000_s_4_800 = '6.56250e-14*ic_cap*ic_cap+3.75000e-14*ic_cap+1.14000e-11'
+ mcrdlm5m3_cf_w_1_600_s_10_000 = '-2.81250e-13*ic_cap*ic_cap+-1.75000e-13*ic_cap+4.85000e-11'
+ mcrdlm5m3_cf_w_1_600_s_12_000 = '-2.71875e-13*ic_cap*ic_cap+-1.62500e-13*ic_cap+4.92000e-11'
+ mcrdlm5m3_cf_w_1_600_s_1_600 = '-1.12500e-13*ic_cap*ic_cap+-7.50000e-14*ic_cap+1.83000e-11'
+ mcrdlm5m3_cf_w_1_600_s_1_700 = '-1.25000e-13*ic_cap*ic_cap+-7.50000e-14*ic_cap+1.93000e-11'
+ mcrdlm5m3_cf_w_1_600_s_1_900 = '-1.37500e-13*ic_cap*ic_cap+-7.50000e-14*ic_cap+2.12000e-11'
+ mcrdlm5m3_cf_w_1_600_s_2_000 = '-1.53125e-13*ic_cap*ic_cap+-8.75000e-14*ic_cap+2.22000e-11'
+ mcrdlm5m3_cf_w_1_600_s_2_400 = '-1.84375e-13*ic_cap*ic_cap+-1.12500e-13*ic_cap+2.57000e-11'
+ mcrdlm5m3_cf_w_1_600_s_2_800 = '-2.06250e-13*ic_cap*ic_cap+-1.25000e-13*ic_cap+2.88000e-11'
+ mcrdlm5m3_cf_w_1_600_s_3_200 = '-2.28125e-13*ic_cap*ic_cap+-1.37500e-13*ic_cap+3.16000e-11'
+ mcrdlm5m3_cf_w_1_600_s_4_800 = '-2.75000e-13*ic_cap*ic_cap+-1.75000e-13*ic_cap+3.98000e-11'
+ mcrdlm5m3_cf_w_4_000_s_10_000 = '-2.68750e-13*ic_cap*ic_cap+-1.75000e-13*ic_cap+4.90000e-11'
+ mcrdlm5m3_cf_w_4_000_s_12_000 = '-2.53125e-13*ic_cap*ic_cap+-1.62500e-13*ic_cap+4.97000e-11'
+ mcrdlm5m3_cf_w_4_000_s_1_600 = '-1.12500e-13*ic_cap*ic_cap+-7.50000e-14*ic_cap+1.83000e-11'
+ mcrdlm5m3_cf_w_4_000_s_1_700 = '-1.25000e-13*ic_cap*ic_cap+-7.50000e-14*ic_cap+1.93000e-11'
+ mcrdlm5m3_cf_w_4_000_s_1_900 = '-1.37500e-13*ic_cap*ic_cap+-7.50000e-14*ic_cap+2.12000e-11'
+ mcrdlm5m3_cf_w_4_000_s_2_000 = '-1.50000e-13*ic_cap*ic_cap+-7.50000e-14*ic_cap+2.22000e-11'
+ mcrdlm5m3_cf_w_4_000_s_2_400 = '-1.78125e-13*ic_cap*ic_cap+-1.12500e-13*ic_cap+2.57000e-11'
+ mcrdlm5m3_cf_w_4_000_s_2_800 = '-2.06250e-13*ic_cap*ic_cap+-1.25000e-13*ic_cap+2.89000e-11'
+ mcrdlm5m3_cf_w_4_000_s_3_200 = '-2.28125e-13*ic_cap*ic_cap+-1.37500e-13*ic_cap+3.17000e-11'
+ mcrdlm5m3_cf_w_4_000_s_4_800 = '-2.71875e-13*ic_cap*ic_cap+-1.62500e-13*ic_cap+4.00000e-11'
+ mcrdlm5m4_ca_w_1_600_s_10_000 = '-1.16250e-06*ic_cap*ic_cap+-5.75000e-07*ic_cap+7.39000e-05'
+ mcrdlm5m4_ca_w_1_600_s_12_000 = '-1.16250e-06*ic_cap*ic_cap+-5.75000e-07*ic_cap+7.39000e-05'
+ mcrdlm5m4_ca_w_1_600_s_1_600 = '-1.16250e-06*ic_cap*ic_cap+-5.75000e-07*ic_cap+7.39000e-05'
+ mcrdlm5m4_ca_w_1_600_s_1_700 = '-1.16250e-06*ic_cap*ic_cap+-5.75000e-07*ic_cap+7.39000e-05'
+ mcrdlm5m4_ca_w_1_600_s_1_900 = '-1.16250e-06*ic_cap*ic_cap+-5.75000e-07*ic_cap+7.39000e-05'
+ mcrdlm5m4_ca_w_1_600_s_2_000 = '-1.16250e-06*ic_cap*ic_cap+-5.75000e-07*ic_cap+7.39000e-05'
+ mcrdlm5m4_ca_w_1_600_s_2_400 = '-1.16250e-06*ic_cap*ic_cap+-5.75000e-07*ic_cap+7.39000e-05'
+ mcrdlm5m4_ca_w_1_600_s_2_800 = '-1.16250e-06*ic_cap*ic_cap+-5.75000e-07*ic_cap+7.39000e-05'
+ mcrdlm5m4_ca_w_1_600_s_3_200 = '-1.16250e-06*ic_cap*ic_cap+-5.75000e-07*ic_cap+7.39000e-05'
+ mcrdlm5m4_ca_w_1_600_s_4_800 = '-1.16250e-06*ic_cap*ic_cap+-5.75000e-07*ic_cap+7.39000e-05'
+ mcrdlm5m4_ca_w_4_000_s_10_000 = '-1.16250e-06*ic_cap*ic_cap+-5.75000e-07*ic_cap+7.39000e-05'
+ mcrdlm5m4_ca_w_4_000_s_12_000 = '-1.16250e-06*ic_cap*ic_cap+-5.75000e-07*ic_cap+7.39000e-05'
+ mcrdlm5m4_ca_w_4_000_s_1_600 = '-1.16250e-06*ic_cap*ic_cap+-5.75000e-07*ic_cap+7.39000e-05'
+ mcrdlm5m4_ca_w_4_000_s_1_700 = '-1.16250e-06*ic_cap*ic_cap+-5.75000e-07*ic_cap+7.39000e-05'
+ mcrdlm5m4_ca_w_4_000_s_1_900 = '-1.16250e-06*ic_cap*ic_cap+-5.75000e-07*ic_cap+7.39000e-05'
+ mcrdlm5m4_ca_w_4_000_s_2_000 = '-1.16250e-06*ic_cap*ic_cap+-5.75000e-07*ic_cap+7.39000e-05'
+ mcrdlm5m4_ca_w_4_000_s_2_400 = '-1.16250e-06*ic_cap*ic_cap+-5.75000e-07*ic_cap+7.39000e-05'
+ mcrdlm5m4_ca_w_4_000_s_2_800 = '-1.16250e-06*ic_cap*ic_cap+-5.75000e-07*ic_cap+7.39000e-05'
+ mcrdlm5m4_ca_w_4_000_s_3_200 = '-1.16250e-06*ic_cap*ic_cap+-5.75000e-07*ic_cap+7.39000e-05'
+ mcrdlm5m4_ca_w_4_000_s_4_800 = '-1.16250e-06*ic_cap*ic_cap+-5.75000e-07*ic_cap+7.39000e-05'
+ mcrdlm5m4_cc_w_1_600_s_10_000 = '1.29688e-14*ic_cap*ic_cap+5.62500e-15*ic_cap+4.30000e-13'
+ mcrdlm5m4_cc_w_1_600_s_12_000 = '7.50000e-15*ic_cap*ic_cap+-1.25000e-15*ic_cap+1.80000e-13'
+ mcrdlm5m4_cc_w_1_600_s_1_600 = '-2.53125e-13*ic_cap*ic_cap+-1.87500e-13*ic_cap+4.40000e-11'
+ mcrdlm5m4_cc_w_1_600_s_1_700 = '-2.09375e-13*ic_cap*ic_cap+-1.62500e-13*ic_cap+4.03000e-11'
+ mcrdlm5m4_cc_w_1_600_s_1_900 = '-1.34375e-13*ic_cap*ic_cap+-1.12500e-13*ic_cap+3.40000e-11'
+ mcrdlm5m4_cc_w_1_600_s_2_000 = '-1.12500e-13*ic_cap*ic_cap+-1.00000e-13*ic_cap+3.15000e-11'
+ mcrdlm5m4_cc_w_1_600_s_2_400 = '-3.12500e-14*ic_cap*ic_cap+-5.00000e-14*ic_cap+2.33000e-11'
+ mcrdlm5m4_cc_w_1_600_s_2_800 = '9.37500e-15*ic_cap*ic_cap+-1.25000e-14*ic_cap+1.77000e-11'
+ mcrdlm5m4_cc_w_1_600_s_3_200 = '3.12500e-14*ic_cap*ic_cap+2.01948e-28*ic_cap+1.37000e-11'
+ mcrdlm5m4_cc_w_1_600_s_4_800 = '4.62500e-14*ic_cap*ic_cap+2.75000e-14*ic_cap+5.39000e-12'
+ mcrdlm5m4_cc_w_4_000_s_10_000 = '2.00000e-14*ic_cap*ic_cap+1.00000e-14*ic_cap+4.45000e-13'
+ mcrdlm5m4_cc_w_4_000_s_12_000 = '1.15625e-14*ic_cap*ic_cap+2.50000e-15*ic_cap+1.80000e-13'
+ mcrdlm5m4_cc_w_4_000_s_1_600 = '-2.25000e-13*ic_cap*ic_cap+-1.50000e-13*ic_cap+4.55000e-11'
+ mcrdlm5m4_cc_w_4_000_s_1_700 = '-1.75000e-13*ic_cap*ic_cap+-1.50000e-13*ic_cap+4.16000e-11'
+ mcrdlm5m4_cc_w_4_000_s_1_900 = '-1.03125e-13*ic_cap*ic_cap+-8.75000e-14*ic_cap+3.53000e-11'
+ mcrdlm5m4_cc_w_4_000_s_2_000 = '-6.87500e-14*ic_cap*ic_cap+-5.00000e-14*ic_cap+3.25000e-11'
+ mcrdlm5m4_cc_w_4_000_s_2_400 = '-6.25000e-15*ic_cap*ic_cap+-2.50000e-14*ic_cap+2.43000e-11'
+ mcrdlm5m4_cc_w_4_000_s_2_800 = '3.12500e-14*ic_cap*ic_cap+1.86000e-11'
+ mcrdlm5m4_cc_w_4_000_s_3_200 = '5.31250e-14*ic_cap*ic_cap+1.25000e-14*ic_cap+1.44000e-11'
+ mcrdlm5m4_cc_w_4_000_s_4_800 = '6.06250e-14*ic_cap*ic_cap+4.00000e-14*ic_cap+5.85000e-12'
+ mcrdlm5m4_cf_w_1_600_s_10_000 = '-6.00000e-13*ic_cap*ic_cap+-3.50000e-13*ic_cap+7.23000e-11'
+ mcrdlm5m4_cf_w_1_600_s_12_000 = '-5.90625e-13*ic_cap*ic_cap+-3.37500e-13*ic_cap+7.25000e-11'
+ mcrdlm5m4_cf_w_1_600_s_1_600 = '-4.34375e-13*ic_cap*ic_cap+-2.37500e-13*ic_cap+4.21000e-11'
+ mcrdlm5m4_cf_w_1_600_s_1_700 = '-4.53125e-13*ic_cap*ic_cap+-2.37500e-13*ic_cap+4.38000e-11'
+ mcrdlm5m4_cf_w_1_600_s_1_900 = '-4.93750e-13*ic_cap*ic_cap+-2.75000e-13*ic_cap+4.70000e-11'
+ mcrdlm5m4_cf_w_1_600_s_2_000 = '-5.06250e-13*ic_cap*ic_cap+-2.75000e-13*ic_cap+4.84000e-11'
+ mcrdlm5m4_cf_w_1_600_s_2_400 = '-5.53125e-13*ic_cap*ic_cap+-2.87500e-13*ic_cap+5.34000e-11'
+ mcrdlm5m4_cf_w_1_600_s_2_800 = '-5.81250e-13*ic_cap*ic_cap+-3.25000e-13*ic_cap+5.73000e-11'
+ mcrdlm5m4_cf_w_1_600_s_3_200 = '-5.96875e-13*ic_cap*ic_cap+-3.37500e-13*ic_cap+6.03000e-11'
+ mcrdlm5m4_cf_w_1_600_s_4_800 = '-6.18750e-13*ic_cap*ic_cap+-3.50000e-13*ic_cap+6.74000e-11'
+ mcrdlm5m4_cf_w_4_000_s_10_000 = '-5.75000e-13*ic_cap*ic_cap+-3.25000e-13*ic_cap+7.29000e-11'
+ mcrdlm5m4_cf_w_4_000_s_12_000 = '-5.68750e-13*ic_cap*ic_cap+-3.25000e-13*ic_cap+7.32000e-11'
+ mcrdlm5m4_cf_w_4_000_s_1_600 = '-4.37500e-13*ic_cap*ic_cap+-2.25000e-13*ic_cap+4.22000e-11'
+ mcrdlm5m4_cf_w_4_000_s_1_700 = '-4.59375e-13*ic_cap*ic_cap+-2.37500e-13*ic_cap+4.39000e-11'
+ mcrdlm5m4_cf_w_4_000_s_1_900 = '-4.90625e-13*ic_cap*ic_cap+-2.62500e-13*ic_cap+4.70000e-11'
+ mcrdlm5m4_cf_w_4_000_s_2_000 = '-4.96875e-13*ic_cap*ic_cap+-2.62500e-13*ic_cap+4.83000e-11'
+ mcrdlm5m4_cf_w_4_000_s_2_400 = '-5.43750e-13*ic_cap*ic_cap+-3.00000e-13*ic_cap+5.33000e-11'
+ mcrdlm5m4_cf_w_4_000_s_2_800 = '-5.78125e-13*ic_cap*ic_cap+-3.12500e-13*ic_cap+5.73000e-11'
+ mcrdlm5m4_cf_w_4_000_s_3_200 = '-6.00000e-13*ic_cap*ic_cap+-3.25000e-13*ic_cap+6.05000e-11'
+ mcrdlm5m4_cf_w_4_000_s_4_800 = '-6.12500e-13*ic_cap*ic_cap+-3.50000e-13*ic_cap+6.77000e-11'
+ mcrdlm5p1_ca_w_1_600_s_10_000 = '-1.18750e-07*ic_cap*ic_cap+-7.50000e-08*ic_cap+1.27000e-05'
+ mcrdlm5p1_ca_w_1_600_s_12_000 = '-1.18750e-07*ic_cap*ic_cap+-7.50000e-08*ic_cap+1.27000e-05'
+ mcrdlm5p1_ca_w_1_600_s_1_600 = '-1.18750e-07*ic_cap*ic_cap+-7.50000e-08*ic_cap+1.27000e-05'
+ mcrdlm5p1_ca_w_1_600_s_1_700 = '-1.18750e-07*ic_cap*ic_cap+-7.50000e-08*ic_cap+1.27000e-05'
+ mcrdlm5p1_ca_w_1_600_s_1_900 = '-1.18750e-07*ic_cap*ic_cap+-7.50000e-08*ic_cap+1.27000e-05'
+ mcrdlm5p1_ca_w_1_600_s_2_000 = '-1.18750e-07*ic_cap*ic_cap+-7.50000e-08*ic_cap+1.27000e-05'
+ mcrdlm5p1_ca_w_1_600_s_2_400 = '-1.18750e-07*ic_cap*ic_cap+-7.50000e-08*ic_cap+1.27000e-05'
+ mcrdlm5p1_ca_w_1_600_s_2_800 = '-1.18750e-07*ic_cap*ic_cap+-7.50000e-08*ic_cap+1.27000e-05'
+ mcrdlm5p1_ca_w_1_600_s_3_200 = '-1.18750e-07*ic_cap*ic_cap+-7.50000e-08*ic_cap+1.27000e-05'
+ mcrdlm5p1_ca_w_1_600_s_4_800 = '-1.18750e-07*ic_cap*ic_cap+-7.50000e-08*ic_cap+1.27000e-05'
+ mcrdlm5p1_ca_w_4_000_s_10_000 = '-1.18750e-07*ic_cap*ic_cap+-7.50000e-08*ic_cap+1.27000e-05'
+ mcrdlm5p1_ca_w_4_000_s_12_000 = '-1.18750e-07*ic_cap*ic_cap+-7.50000e-08*ic_cap+1.27000e-05'
+ mcrdlm5p1_ca_w_4_000_s_1_600 = '-1.18750e-07*ic_cap*ic_cap+-7.50000e-08*ic_cap+1.27000e-05'
+ mcrdlm5p1_ca_w_4_000_s_1_700 = '-1.18750e-07*ic_cap*ic_cap+-7.50000e-08*ic_cap+1.27000e-05'
+ mcrdlm5p1_ca_w_4_000_s_1_900 = '-1.18750e-07*ic_cap*ic_cap+-7.50000e-08*ic_cap+1.27000e-05'
+ mcrdlm5p1_ca_w_4_000_s_2_000 = '-1.18750e-07*ic_cap*ic_cap+-7.50000e-08*ic_cap+1.27000e-05'
+ mcrdlm5p1_ca_w_4_000_s_2_400 = '-1.18750e-07*ic_cap*ic_cap+-7.50000e-08*ic_cap+1.27000e-05'
+ mcrdlm5p1_ca_w_4_000_s_2_800 = '-1.18750e-07*ic_cap*ic_cap+-7.50000e-08*ic_cap+1.27000e-05'
+ mcrdlm5p1_ca_w_4_000_s_3_200 = '-1.18750e-07*ic_cap*ic_cap+-7.50000e-08*ic_cap+1.27000e-05'
+ mcrdlm5p1_ca_w_4_000_s_4_800 = '-1.18750e-07*ic_cap*ic_cap+-7.50000e-08*ic_cap+1.27000e-05'
+ mcrdlm5p1_cc_w_1_600_s_10_000 = '5.71875e-14*ic_cap*ic_cap+3.62500e-14*ic_cap+4.25000e-12'
+ mcrdlm5p1_cc_w_1_600_s_12_000 = '4.56250e-14*ic_cap*ic_cap+3.00000e-14*ic_cap+2.44000e-12'
+ mcrdlm5p1_cc_w_1_600_s_1_600 = '-3.93750e-13*ic_cap*ic_cap+-2.50000e-13*ic_cap+6.60000e-11'
+ mcrdlm5p1_cc_w_1_600_s_1_700 = '-3.40625e-13*ic_cap*ic_cap+-2.37500e-13*ic_cap+6.21000e-11'
+ mcrdlm5p1_cc_w_1_600_s_1_900 = '-2.68750e-13*ic_cap*ic_cap+-1.75000e-13*ic_cap+5.57000e-11'
+ mcrdlm5p1_cc_w_1_600_s_2_000 = '-2.31250e-13*ic_cap*ic_cap+-1.75000e-13*ic_cap+5.29000e-11'
+ mcrdlm5p1_cc_w_1_600_s_2_400 = '-1.37500e-13*ic_cap*ic_cap+-1.00000e-13*ic_cap+4.38000e-11'
+ mcrdlm5p1_cc_w_1_600_s_2_800 = '-8.43750e-14*ic_cap*ic_cap+-6.25000e-14*ic_cap+3.73000e-11'
+ mcrdlm5p1_cc_w_1_600_s_3_200 = '-4.37500e-14*ic_cap*ic_cap+-2.50000e-14*ic_cap+3.21000e-11'
+ mcrdlm5p1_cc_w_1_600_s_4_800 = '3.43750e-14*ic_cap*ic_cap+1.25000e-14*ic_cap+1.90000e-11'
+ mcrdlm5p1_cc_w_4_000_s_10_000 = '6.96875e-14*ic_cap*ic_cap+4.62500e-14*ic_cap+4.47000e-12'
+ mcrdlm5p1_cc_w_4_000_s_12_000 = '5.37500e-14*ic_cap*ic_cap+3.25000e-14*ic_cap+2.57000e-12'
+ mcrdlm5p1_cc_w_4_000_s_1_600 = '-3.37500e-13*ic_cap*ic_cap+-2.25000e-13*ic_cap+6.88000e-11'
+ mcrdlm5p1_cc_w_4_000_s_1_700 = '-2.84375e-13*ic_cap*ic_cap+-1.87500e-13*ic_cap+6.47000e-11'
+ mcrdlm5p1_cc_w_4_000_s_1_900 = '-2.09375e-13*ic_cap*ic_cap+-1.62500e-13*ic_cap+5.80000e-11'
+ mcrdlm5p1_cc_w_4_000_s_2_000 = '-1.78125e-13*ic_cap*ic_cap+-1.37500e-13*ic_cap+5.51000e-11'
+ mcrdlm5p1_cc_w_4_000_s_2_400 = '-1.00000e-13*ic_cap*ic_cap+-7.50000e-14*ic_cap+4.59000e-11'
+ mcrdlm5p1_cc_w_4_000_s_2_800 = '-4.06250e-14*ic_cap*ic_cap+-3.75000e-14*ic_cap+3.89000e-11'
+ mcrdlm5p1_cc_w_4_000_s_3_200 = '-6.25000e-15*ic_cap*ic_cap+3.35000e-11'
+ mcrdlm5p1_cc_w_4_000_s_4_800 = '6.56250e-14*ic_cap*ic_cap+3.75000e-14*ic_cap+1.98000e-11'
+ mcrdlm5p1_cf_w_1_600_s_10_000 = '-2.28125e-13*ic_cap*ic_cap+-1.37500e-13*ic_cap+3.55000e-11'
+ mcrdlm5p1_cf_w_1_600_s_12_000 = '-2.21875e-13*ic_cap*ic_cap+-1.37500e-13*ic_cap+3.72000e-11'
+ mcrdlm5p1_cf_w_1_600_s_1_600 = '-6.21875e-14*ic_cap*ic_cap+-3.87500e-14*ic_cap+9.71000e-12'
+ mcrdlm5p1_cf_w_1_600_s_1_700 = '-6.90625e-14*ic_cap*ic_cap+-4.37500e-14*ic_cap+1.03000e-11'
+ mcrdlm5p1_cf_w_1_600_s_1_900 = '-7.96875e-14*ic_cap*ic_cap+-4.37500e-14*ic_cap+1.14000e-11'
+ mcrdlm5p1_cf_w_1_600_s_2_000 = '-8.12500e-14*ic_cap*ic_cap+-5.00000e-14*ic_cap+1.19000e-11'
+ mcrdlm5p1_cf_w_1_600_s_2_400 = '-1.03125e-13*ic_cap*ic_cap+-6.25000e-14*ic_cap+1.41000e-11'
+ mcrdlm5p1_cf_w_1_600_s_2_800 = '-1.18750e-13*ic_cap*ic_cap+-7.50000e-14*ic_cap+1.61000e-11'
+ mcrdlm5p1_cf_w_1_600_s_3_200 = '-1.40625e-13*ic_cap*ic_cap+-8.75000e-14*ic_cap+1.81000e-11'
+ mcrdlm5p1_cf_w_1_600_s_4_800 = '-1.90625e-13*ic_cap*ic_cap+-1.12500e-13*ic_cap+2.46000e-11'
+ mcrdlm5p1_cf_w_4_000_s_10_000 = '-2.18750e-13*ic_cap*ic_cap+-1.50000e-13*ic_cap+3.61000e-11'
+ mcrdlm5p1_cf_w_4_000_s_12_000 = '-2.09375e-13*ic_cap*ic_cap+-1.37500e-13*ic_cap+3.79000e-11'
+ mcrdlm5p1_cf_w_4_000_s_1_600 = '-6.25000e-14*ic_cap*ic_cap+-3.75000e-14*ic_cap+9.71000e-12'
+ mcrdlm5p1_cf_w_4_000_s_1_700 = '-6.93750e-14*ic_cap*ic_cap+-3.75000e-14*ic_cap+1.03000e-11'
+ mcrdlm5p1_cf_w_4_000_s_1_900 = '-7.90625e-14*ic_cap*ic_cap+-4.12500e-14*ic_cap+1.14000e-11'
+ mcrdlm5p1_cf_w_4_000_s_2_000 = '-8.75000e-14*ic_cap*ic_cap+-5.00000e-14*ic_cap+1.20000e-11'
+ mcrdlm5p1_cf_w_4_000_s_2_400 = '-1.03125e-13*ic_cap*ic_cap+-6.25000e-14*ic_cap+1.41000e-11'
+ mcrdlm5p1_cf_w_4_000_s_2_800 = '-1.25000e-13*ic_cap*ic_cap+-7.50000e-14*ic_cap+1.62000e-11'
+ mcrdlm5p1_cf_w_4_000_s_3_200 = '-1.37500e-13*ic_cap*ic_cap+-7.50000e-14*ic_cap+1.81000e-11'
+ mcrdlm5p1_cf_w_4_000_s_4_800 = '-1.84375e-13*ic_cap*ic_cap+-1.12500e-13*ic_cap+2.47000e-11'
+ mcrdlp1_ca_w_10_000_s_10_000 = '-2.37500e-08*ic_cap*ic_cap+-1.50000e-08*ic_cap+2.68000e-06'
+ mcrdlp1_ca_w_10_000_s_12_000 = '-2.37500e-08*ic_cap*ic_cap+-1.50000e-08*ic_cap+2.68000e-06'
+ mcrdlp1_ca_w_10_000_s_30_000 = '-2.37500e-08*ic_cap*ic_cap+-1.50000e-08*ic_cap+2.68000e-06'
+ mcrdlp1_ca_w_10_000_s_5_000 = '-2.37500e-08*ic_cap*ic_cap+-1.50000e-08*ic_cap+2.68000e-06'
+ mcrdlp1_ca_w_10_000_s_8_000 = '-2.37500e-08*ic_cap*ic_cap+-1.50000e-08*ic_cap+2.68000e-06'
+ mcrdlp1_ca_w_40_000_s_10_000 = '-2.37500e-08*ic_cap*ic_cap+-1.50000e-08*ic_cap+2.68000e-06'
+ mcrdlp1_ca_w_40_000_s_12_000 = '-2.37500e-08*ic_cap*ic_cap+-1.50000e-08*ic_cap+2.68000e-06'
+ mcrdlp1_ca_w_40_000_s_30_000 = '-2.37500e-08*ic_cap*ic_cap+-1.50000e-08*ic_cap+2.68000e-06'
+ mcrdlp1_ca_w_40_000_s_5_000 = '-2.37500e-08*ic_cap*ic_cap+-1.50000e-08*ic_cap+2.68000e-06'
+ mcrdlp1_ca_w_40_000_s_8_000 = '-2.37500e-08*ic_cap*ic_cap+-1.50000e-08*ic_cap+2.68000e-06'
+ mcrdlp1_cc_w_10_000_s_10_000 = '-2.37500e-13*ic_cap*ic_cap+-1.50000e-13*ic_cap+3.16000e-11'
+ mcrdlp1_cc_w_10_000_s_12_000 = '-1.90625e-13*ic_cap*ic_cap+-1.37500e-13*ic_cap+2.76000e-11'
+ mcrdlp1_cc_w_10_000_s_30_000 = '-6.25000e-14*ic_cap*ic_cap+-5.00000e-14*ic_cap+1.21000e-11'
+ mcrdlp1_cc_w_10_000_s_5_000 = '-5.62500e-13*ic_cap*ic_cap+-3.50000e-13*ic_cap+5.12000e-11'
+ mcrdlp1_cc_w_10_000_s_8_000 = '-3.15625e-13*ic_cap*ic_cap+-1.87500e-13*ic_cap+3.71000e-11'
+ mcrdlp1_cc_w_40_000_s_10_000 = '-2.40625e-13*ic_cap*ic_cap+-1.62500e-13*ic_cap+4.15000e-11'
+ mcrdlp1_cc_w_40_000_s_12_000 = '-1.93750e-13*ic_cap*ic_cap+-1.25000e-13*ic_cap+3.71000e-11'
+ mcrdlp1_cc_w_40_000_s_30_000 = '-5.93750e-14*ic_cap*ic_cap+-3.75000e-14*ic_cap+1.92000e-11'
+ mcrdlp1_cc_w_40_000_s_5_000 = '-5.62500e-13*ic_cap*ic_cap+-3.50000e-13*ic_cap+6.25000e-11'
+ mcrdlp1_cc_w_40_000_s_8_000 = '-3.15625e-13*ic_cap*ic_cap+-2.12500e-13*ic_cap+4.75000e-11'
+ mcrdlp1_cf_w_10_000_s_10_000 = '-4.37500e-14*ic_cap*ic_cap+-2.50000e-14*ic_cap+1.13000e-11'
+ mcrdlp1_cf_w_10_000_s_12_000 = '-6.56250e-14*ic_cap*ic_cap+-3.75000e-14*ic_cap+1.31000e-11'
+ mcrdlp1_cf_w_10_000_s_30_000 = '-1.34375e-13*ic_cap*ic_cap+-8.75000e-14*ic_cap+2.34000e-11'
+ mcrdlp1_cf_w_10_000_s_5_000 = '-3.12500e-16*ic_cap*ic_cap+-1.25000e-15*ic_cap+6.21000e-12'
+ mcrdlp1_cf_w_10_000_s_8_000 = '-2.81250e-14*ic_cap*ic_cap+-1.75000e-14*ic_cap+9.38000e-12'
+ mcrdlp1_cf_w_40_000_s_10_000 = '-5.00000e-14*ic_cap*ic_cap+-2.50000e-14*ic_cap+1.15000e-11'
+ mcrdlp1_cf_w_40_000_s_12_000 = '-5.93750e-14*ic_cap*ic_cap+-3.75000e-14*ic_cap+1.32000e-11'
+ mcrdlp1_cf_w_40_000_s_30_000 = '-1.28125e-13*ic_cap*ic_cap+-8.75000e-14*ic_cap+2.41000e-11'
+ mcrdlp1_cf_w_40_000_s_5_000 = '-3.43750e-15*ic_cap*ic_cap+-1.25000e-15*ic_cap+6.36000e-12'
+ mcrdlp1_cf_w_40_000_s_8_000 = '-3.15625e-14*ic_cap*ic_cap+-2.12500e-14*ic_cap+9.54000e-12'
+ mcrdlp1f_ca_w_0_150_s_0_210 = '-1.44688e-06*ic_cap*ic_cap+-7.87500e-07*ic_cap+1.09000e-04'
+ mcrdlp1f_ca_w_0_150_s_0_263 = '-1.44688e-06*ic_cap*ic_cap+-7.87500e-07*ic_cap+1.09000e-04'
+ mcrdlp1f_ca_w_0_150_s_0_315 = '-1.44688e-06*ic_cap*ic_cap+-7.87500e-07*ic_cap+1.09000e-04'
+ mcrdlp1f_ca_w_0_150_s_0_420 = '-1.44688e-06*ic_cap*ic_cap+-7.87500e-07*ic_cap+1.09000e-04'
+ mcrdlp1f_ca_w_0_150_s_0_525 = '-1.44688e-06*ic_cap*ic_cap+-7.87500e-07*ic_cap+1.09000e-04'
+ mcrdlp1f_ca_w_0_150_s_0_630 = '-1.44688e-06*ic_cap*ic_cap+-7.87500e-07*ic_cap+1.09000e-04'
+ mcrdlp1f_ca_w_0_150_s_0_840 = '-1.44688e-06*ic_cap*ic_cap+-7.87500e-07*ic_cap+1.09000e-04'
+ mcrdlp1f_ca_w_0_150_s_1_260 = '-1.44688e-06*ic_cap*ic_cap+-7.87500e-07*ic_cap+1.09000e-04'
+ mcrdlp1f_ca_w_0_150_s_2_310 = '-1.44688e-06*ic_cap*ic_cap+-7.87500e-07*ic_cap+1.09000e-04'
+ mcrdlp1f_ca_w_0_150_s_5_250 = '-1.44688e-06*ic_cap*ic_cap+-7.87500e-07*ic_cap+1.09000e-04'
+ mcrdlp1f_ca_w_1_200_s_0_210 = '-1.44688e-06*ic_cap*ic_cap+-7.87500e-07*ic_cap+1.09000e-04'
+ mcrdlp1f_ca_w_1_200_s_0_263 = '-1.44688e-06*ic_cap*ic_cap+-7.87500e-07*ic_cap+1.09000e-04'
+ mcrdlp1f_ca_w_1_200_s_0_315 = '-1.44688e-06*ic_cap*ic_cap+-7.87500e-07*ic_cap+1.09000e-04'
+ mcrdlp1f_ca_w_1_200_s_0_420 = '-1.44688e-06*ic_cap*ic_cap+-7.87500e-07*ic_cap+1.09000e-04'
+ mcrdlp1f_ca_w_1_200_s_0_525 = '-1.44688e-06*ic_cap*ic_cap+-7.87500e-07*ic_cap+1.09000e-04'
+ mcrdlp1f_ca_w_1_200_s_0_630 = '-1.44688e-06*ic_cap*ic_cap+-7.87500e-07*ic_cap+1.09000e-04'
+ mcrdlp1f_ca_w_1_200_s_0_840 = '-1.44688e-06*ic_cap*ic_cap+-7.87500e-07*ic_cap+1.09000e-04'
+ mcrdlp1f_ca_w_1_200_s_1_260 = '-1.44688e-06*ic_cap*ic_cap+-7.87500e-07*ic_cap+1.09000e-04'
+ mcrdlp1f_ca_w_1_200_s_2_310 = '-1.44688e-06*ic_cap*ic_cap+-7.87500e-07*ic_cap+1.09000e-04'
+ mcrdlp1f_ca_w_1_200_s_5_250 = '-1.44688e-06*ic_cap*ic_cap+-7.87500e-07*ic_cap+1.09000e-04'
+ mcrdlp1f_cc_w_0_150_s_0_210 = '-5.62500e-13*ic_cap*ic_cap+-3.25000e-13*ic_cap+7.57000e-11'
+ mcrdlp1f_cc_w_0_150_s_0_263 = '-3.71875e-13*ic_cap*ic_cap+-2.12500e-13*ic_cap+6.15000e-11'
+ mcrdlp1f_cc_w_0_150_s_0_315 = '-2.62500e-13*ic_cap*ic_cap+-1.50000e-13*ic_cap+5.24000e-11'
+ mcrdlp1f_cc_w_0_150_s_0_420 = '-1.37500e-13*ic_cap*ic_cap+-7.50000e-14*ic_cap+3.98000e-11'
+ mcrdlp1f_cc_w_0_150_s_0_525 = '-8.12500e-14*ic_cap*ic_cap+-5.00000e-14*ic_cap+3.23000e-11'
+ mcrdlp1f_cc_w_0_150_s_0_630 = '-4.37500e-14*ic_cap*ic_cap+-2.50000e-14*ic_cap+2.69000e-11'
+ mcrdlp1f_cc_w_0_150_s_0_840 = '-6.25000e-15*ic_cap*ic_cap+1.95000e-11'
+ mcrdlp1f_cc_w_0_150_s_1_260 = '1.87500e-14*ic_cap*ic_cap+1.11000e-11'
+ mcrdlp1f_cc_w_0_150_s_2_310 = '1.78125e-14*ic_cap*ic_cap+1.37500e-14*ic_cap+4.42000e-12'
+ mcrdlp1f_cc_w_0_150_s_5_250 = '4.09375e-15*ic_cap*ic_cap+4.62500e-15*ic_cap+8.77000e-13'
+ mcrdlp1f_cc_w_1_200_s_0_210 = '-5.59375e-13*ic_cap*ic_cap+-3.12500e-13*ic_cap+9.30000e-11'
+ mcrdlp1f_cc_w_1_200_s_0_263 = '-3.50000e-13*ic_cap*ic_cap+-2.00000e-13*ic_cap+7.73000e-11'
+ mcrdlp1f_cc_w_1_200_s_0_315 = '-2.40625e-13*ic_cap*ic_cap+-1.37500e-13*ic_cap+6.69000e-11'
+ mcrdlp1f_cc_w_1_200_s_0_420 = '-1.21875e-13*ic_cap*ic_cap+-6.25000e-14*ic_cap+5.31000e-11'
+ mcrdlp1f_cc_w_1_200_s_0_525 = '-5.93750e-14*ic_cap*ic_cap+-3.75000e-14*ic_cap+4.42000e-11'
+ mcrdlp1f_cc_w_1_200_s_0_630 = '-2.81250e-14*ic_cap*ic_cap+-1.25000e-14*ic_cap+3.79000e-11'
+ mcrdlp1f_cc_w_1_200_s_0_840 = '3.12500e-15*ic_cap*ic_cap+1.25000e-14*ic_cap+2.92000e-11'
+ mcrdlp1f_cc_w_1_200_s_1_260 = '3.12500e-14*ic_cap*ic_cap+2.50000e-14*ic_cap+1.93000e-11'
+ mcrdlp1f_cc_w_1_200_s_2_310 = '3.53125e-14*ic_cap*ic_cap+2.87500e-14*ic_cap+8.91000e-12'
+ mcrdlp1f_cc_w_1_200_s_5_250 = '1.78125e-14*ic_cap*ic_cap+8.75000e-15*ic_cap+2.15000e-12'
+ mcrdlp1f_cf_w_0_150_s_0_210 = '-9.15625e-14*ic_cap*ic_cap+-5.12500e-14*ic_cap+1.06000e-11'
+ mcrdlp1f_cf_w_0_150_s_0_263 = '-1.15625e-13*ic_cap*ic_cap+-6.25000e-14*ic_cap+1.28000e-11'
+ mcrdlp1f_cf_w_0_150_s_0_315 = '-1.43750e-13*ic_cap*ic_cap+-7.50000e-14*ic_cap+1.50000e-11'
+ mcrdlp1f_cf_w_0_150_s_0_420 = '-1.84375e-13*ic_cap*ic_cap+-1.12500e-13*ic_cap+1.90000e-11'
+ mcrdlp1f_cf_w_0_150_s_0_525 = '-2.18750e-13*ic_cap*ic_cap+-1.25000e-13*ic_cap+2.24000e-11'
+ mcrdlp1f_cf_w_0_150_s_0_630 = '-2.40625e-13*ic_cap*ic_cap+-1.37500e-13*ic_cap+2.53000e-11'
+ mcrdlp1f_cf_w_0_150_s_0_840 = '-2.71875e-13*ic_cap*ic_cap+-1.62500e-13*ic_cap+3.02000e-11'
+ mcrdlp1f_cf_w_0_150_s_1_260 = '-3.00000e-13*ic_cap*ic_cap+-1.75000e-13*ic_cap+3.69000e-11'
+ mcrdlp1f_cf_w_0_150_s_2_310 = '-3.03125e-13*ic_cap*ic_cap+-1.87500e-13*ic_cap+4.30000e-11'
+ mcrdlp1f_cf_w_0_150_s_5_250 = '-2.93750e-13*ic_cap*ic_cap+-1.75000e-13*ic_cap+4.65000e-11'
+ mcrdlp1f_cf_w_1_200_s_0_210 = '-8.93750e-14*ic_cap*ic_cap+-5.00000e-14*ic_cap+1.05000e-11'
+ mcrdlp1f_cf_w_1_200_s_0_263 = '-1.15625e-13*ic_cap*ic_cap+-6.25000e-14*ic_cap+1.28000e-11'
+ mcrdlp1f_cf_w_1_200_s_0_315 = '-1.40625e-13*ic_cap*ic_cap+-8.75000e-14*ic_cap+1.50000e-11'
+ mcrdlp1f_cf_w_1_200_s_0_420 = '-1.81250e-13*ic_cap*ic_cap+-1.00000e-13*ic_cap+1.90000e-11'
+ mcrdlp1f_cf_w_1_200_s_0_525 = '-2.12500e-13*ic_cap*ic_cap+-1.25000e-13*ic_cap+2.25000e-11'
+ mcrdlp1f_cf_w_1_200_s_0_630 = '-2.40625e-13*ic_cap*ic_cap+-1.37500e-13*ic_cap+2.56000e-11'
+ mcrdlp1f_cf_w_1_200_s_0_840 = '-2.71875e-13*ic_cap*ic_cap+-1.62500e-13*ic_cap+3.08000e-11'
+ mcrdlp1f_cf_w_1_200_s_1_260 = '-3.00000e-13*ic_cap*ic_cap+-1.75000e-13*ic_cap+3.80000e-11'
+ mcrdlp1f_cf_w_1_200_s_2_310 = '-3.15625e-13*ic_cap*ic_cap+-1.87500e-13*ic_cap+4.71000e-11'
+ mcrdlp1f_cf_w_1_200_s_5_250 = '-2.93750e-13*ic_cap*ic_cap+-1.75000e-13*ic_cap+5.35000e-11'
+ sky130_fd_pr__nfet_20v0_nvt__hvvsat_mult = '2.48546e-02*hvn_saturation*hvn_saturation+-5.96510e-02*hvn_saturation+1.00000e-18'
+ sky130_fd_pr__nfet_20v0_nvt__k2_diff = '2.67500e-04*hvn_bodyeffect*hvn_bodyeffect+-1.23650e-01'
+ sky130_fd_pr__nfet_20v0_nvt__rdrift_mult = '9.42313e-03*nfet_20v0_nvt*nfet_20v0_nvt+1.17758e-01*nfet_20v0_nvt+7.26100e-01'
+ sky130_fd_pr__nfet_20v0_nvt__vth0_diff = '1.63812e-04*hvntvn_threshold*hvntvn_threshold+3.39563e-02*hvntvn_threshold+3.06540e-02'
+ sky130_fd_pr__nfet_20v0_nvt_iso__hvvsat_mult = '2.48544e-02*hvn_saturation*hvn_saturation+-5.96505e-02*hvn_saturation+1.00000e-18'
+ sky130_fd_pr__nfet_20v0_nvt_iso__rdrift_mult = '2.07703e-02*nfet_20v0_nvt_iso*nfet_20v0_nvt_iso+1.69501e-01*nfet_20v0_nvt_iso+8.20770e-01'
+ sky130_fd_pr__nfet_20v0_nvt_iso__vth0_diff = '2.00325e-04*hvntvn_threshold*hvntvn_threshold+3.47038e-02*hvntvn_threshold+4.46980e-03'
+ sky130_fd_pr__nfet_20v0__ajunction_mult = '8.57188e-04*hvn_diode*hvn_diode+1.47809e-01*hvn_diode+9.95050e-01'
+ sky130_fd_pr__nfet_20v0__dlc_diff = '-4.33125e-09*poly_cd'
+ sky130_fd_pr__nfet_20v0__dwc_diff = '8.04375e-09*ndiff_cd'
+ sky130_fd_pr__nfet_20v0__hvvsat_mult = '1.77529e-02*hvn_saturation*hvn_saturation+-4.26070e-02*hvn_saturation+1.00000e-18'
+ sky130_fd_pr__nfet_20v0__k2_diff = '5.62500e-07*hvn_bodyeffect*hvn_bodyeffect+4.02000e-04*hvn_bodyeffect+-2.74000e-02'
+ sky130_fd_pr__nfet_20v0__lint_diff = '-4.33125e-09*poly_cd'
+ sky130_fd_pr__nfet_20v0__overlap_mult = '6.37187e-03*hvtox*hvtox+-2.25000e-01*hvtox+8.98050e-01'
+ sky130_fd_pr__nfet_20v0__pjunction_mult = '1.53313e-03*hvn_diode*hvn_diode+1.40267e-01*hvn_diode+1.01440e+00'
+ sky130_fd_pr__nfet_20v0__rdrift_mult = '1.18628e-02*nfet_20v0*nfet_20v0+1.65219e-01*nfet_20v0+9.69820e-01'
+ sky130_fd_pr__nfet_20v0__toxe_mult = '1.50000e-02*hvtox+1.00000e+00'
+ sky130_fd_pr__nfet_20v0__vth0_diff = '5.06875e-05*hvn_threshold*hvn_threshold+3.60338e-02*hvn_threshold+3.48240e-02'
+ sky130_fd_pr__nfet_20v0__wint_diff = '8.04375e-09*ndiff_cd'
+ sky130_fd_pr__nfet_20v0_iso__hvvsat_mult = '2.48546e-02*hvn_saturation*hvn_saturation+-5.96511e-02*hvn_saturation+1.00000e-18'
+ sky130_fd_pr__nfet_20v0_iso__k2_diff = '6.75000e-06*hvn_bodyeffect*hvn_bodyeffect+7.95000e-05*hvn_bodyeffect+-1.98730e-02'
+ sky130_fd_pr__nfet_20v0_iso__rdrift_mult = '2.61019e-02*nfet_20v0_iso*nfet_20v0_iso+2.62590e-01*nfet_20v0_iso+9.16610e-01'
+ sky130_fd_pr__nfet_20v0_iso__vth0_diff = '9.62000e-05*hvn_threshold*hvn_threshold+3.58925e-02*hvn_threshold+-1.23920e-03'
+ n20zvtvh1defet_js_mult_pmc = '2.81250e-01*n20zvtvh1defet*n20zvtvh1defet+-1.12500e+00*n20zvtvh1defet+1.00000e+00'
+ sky130_fd_pr__nfet_20v0_zvt__agidl_diff = '1.40625e-16*hvn_subvt*hvn_subvt+-5.62500e-16*hvn_subvt'
+ sky130_fd_pr__nfet_20v0_zvt__ags_diff = '4.64219e-02*hvn_saturation*hvn_saturation+1.85688e-01*hvn_saturation'
+ sky130_fd_pr__nfet_20v0_zvt__keta_diff = '5.85125e-03*hvn_bodyeffect*hvn_bodyeffect+2.34050e-02*hvn_bodyeffect'
+ sky130_fd_pr__nfet_20v0_zvt__rdrift_mult = '4.43304e-02*nfet_20v0_zvt*nfet_20v0_zvt+2.53678e-01*nfet_20v0_zvt+1.00000e+00'
+ sky130_fd_pr__nfet_20v0_zvt__u0_diff = '4.88469e-03*hvn_mobility*hvn_mobility+-1.95388e-02*hvn_mobility'
+ sky130_fd_pr__nfet_20v0_zvt__vth0_diff = '1.07719e-03*hvn_threshold*hvn_threshold+9.52125e-03*hvn_threshold'
+ sky130_fd_pr__nfet_g5v0d10v5__a0_diff_1 = '6.72069e-04*hvn_saturation*hvn_saturation+-2.19321e-02*hvn_saturation+-2.15260e-03'
+ sky130_fd_pr__nfet_g5v0d10v5__a0_diff_10 = '1.21613e-05*hvn_saturation*hvn_saturation+-8.96250e-04*hvn_saturation+-4.36880e-04'
+ sky130_fd_pr__nfet_g5v0d10v5__a0_diff_14 = '6.05656e-04*hvn_saturation*hvn_saturation+-1.46919e-02*hvn_saturation+-2.46390e-02'
+ sky130_fd_pr__nfet_g5v0d10v5__a0_diff_16 = '4.10975e-04*hvn_saturation*hvn_saturation+-9.08413e-03*hvn_saturation+-4.94610e-03'
+ sky130_fd_pr__nfet_g5v0d10v5__a0_diff_17 = '8.95844e-05*hvn_saturation*hvn_saturation+-2.41271e-03*hvn_saturation+-3.59950e-03'
+ sky130_fd_pr__nfet_g5v0d10v5__a0_diff_18 = '3.29313e-05*hvn_saturation*hvn_saturation+-1.54642e-03*hvn_saturation+-5.30120e-03'
+ sky130_fd_pr__nfet_g5v0d10v5__a0_diff_19 = '8.70062e-06*hvn_saturation*hvn_saturation+-7.34127e-04*hvn_saturation+-2.91810e-03'
+ sky130_fd_pr__nfet_g5v0d10v5__a0_diff_22 = '3.97156e-04*hvn_saturation*hvn_saturation+-9.17438e-03*hvn_saturation+-1.08900e-02'
+ sky130_fd_pr__nfet_g5v0d10v5__a0_diff_23 = '5.20947e-05*hvn_saturation*hvn_saturation+-1.92030e-03*hvn_saturation+-8.23330e-03'
+ sky130_fd_pr__nfet_g5v0d10v5__a0_diff_24 = '3.68000e-05*hvn_saturation*hvn_saturation+-1.81113e-03*hvn_saturation+-6.09830e-03'
+ sky130_fd_pr__nfet_g5v0d10v5__a0_diff_25 = '4.13962e-05*hvn_saturation*hvn_saturation+-9.06360e-04*hvn_saturation+-3.75040e-03'
+ sky130_fd_pr__nfet_g5v0d10v5__a0_diff_29 = '3.32619e-04*hvn_saturation*hvn_saturation+-6.99413e-03*hvn_saturation+-5.35540e-03'
+ sky130_fd_pr__nfet_g5v0d10v5__a0_diff_3 = '5.05131e-04*hvn_saturation*hvn_saturation+-9.02875e-03*hvn_saturation+-2.94110e-03'
+ sky130_fd_pr__nfet_g5v0d10v5__a0_diff_30 = '6.13406e-05*hvn_saturation*hvn_saturation+-1.94814e-03*hvn_saturation+-6.72890e-03'
+ sky130_fd_pr__nfet_g5v0d10v5__a0_diff_31 = '3.23156e-05*hvn_saturation*hvn_saturation+-1.65566e-03*hvn_saturation+-4.90340e-03'
+ sky130_fd_pr__nfet_g5v0d10v5__a0_diff_32 = '2.24562e-06*hvn_saturation*hvn_saturation+-5.95357e-04*hvn_saturation+-2.75110e-03'
+ sky130_fd_pr__nfet_g5v0d10v5__a0_diff_4 = '8.43906e-05*hvn_saturation*hvn_saturation+-1.66329e-03*hvn_saturation+-6.99810e-03'
+ sky130_fd_pr__nfet_g5v0d10v5__a0_diff_5 = '2.14063e-05*hvn_saturation*hvn_saturation+-1.15555e-03*hvn_saturation+-2.72390e-03'
+ sky130_fd_pr__nfet_g5v0d10v5__a0_diff_7 = '-1.96365e-02*hvn_saturation*hvn_saturation+6.96438e-02*hvn_saturation+-7.16120e-03'
+ sky130_fd_pr__nfet_g5v0d10v5__a0_diff_8 = '8.52594e-05*hvn_saturation*hvn_saturation+-2.17589e-03*hvn_saturation+-3.47460e-03'
+ sky130_fd_pr__nfet_g5v0d10v5__a0_diff_9 = '3.60938e-06*hvn_saturation*hvn_saturation+-2.53291e-03*hvn_saturation+-3.36410e-03'
+ sky130_fd_pr__nfet_g5v0d10v5__ags_diff_1 = '1.35350e-04*hvn_saturation*hvn_saturation+4.30075e-02*hvn_saturation+-1.91560e-03'
+ sky130_fd_pr__nfet_g5v0d10v5__ags_diff_10 = '-4.76375e-05*hvn_saturation*hvn_saturation+4.66388e-03*hvn_saturation+-1.28630e-03'
+ sky130_fd_pr__nfet_g5v0d10v5__ags_diff_14 = '-2.45562e-04*hvn_saturation*hvn_saturation+3.10073e-02*hvn_saturation+4.32900e-02'
+ sky130_fd_pr__nfet_g5v0d10v5__ags_diff_16 = '-4.68637e-04*hvn_saturation*hvn_saturation+2.68212e-02*hvn_saturation+6.99320e-03'
+ sky130_fd_pr__nfet_g5v0d10v5__ags_diff_17 = '-1.51556e-04*hvn_saturation*hvn_saturation+1.19976e-02*hvn_saturation+3.07540e-03'
+ sky130_fd_pr__nfet_g5v0d10v5__ags_diff_18 = '-7.44375e-05*hvn_saturation*hvn_saturation+7.31975e-03*hvn_saturation+1.51430e-02'
+ sky130_fd_pr__nfet_g5v0d10v5__ags_diff_19 = '-5.88094e-05*hvn_saturation*hvn_saturation+2.96951e-03*hvn_saturation+3.47790e-03'
+ sky130_fd_pr__nfet_g5v0d10v5__ags_diff_22 = '-4.83031e-04*hvn_saturation*hvn_saturation+2.67519e-02*hvn_saturation+2.12210e-02'
+ sky130_fd_pr__nfet_g5v0d10v5__ags_diff_23 = '-1.42062e-04*hvn_saturation*hvn_saturation+8.65450e-03*hvn_saturation+2.25240e-02'
+ sky130_fd_pr__nfet_g5v0d10v5__ags_diff_24 = '-7.59437e-05*hvn_saturation*hvn_saturation+5.63025e-03*hvn_saturation+9.92010e-03'
+ sky130_fd_pr__nfet_g5v0d10v5__ags_diff_25 = '-5.81312e-05*hvn_saturation*hvn_saturation+2.57448e-03*hvn_saturation+5.77920e-03'
+ sky130_fd_pr__nfet_g5v0d10v5__ags_diff_29 = '-4.85944e-04*hvn_saturation*hvn_saturation+2.24673e-02*hvn_saturation+5.52110e-03'
+ sky130_fd_pr__nfet_g5v0d10v5__ags_diff_3 = '-5.13800e-04*hvn_saturation*hvn_saturation+2.62098e-02*hvn_saturation+-2.55020e-03'
+ sky130_fd_pr__nfet_g5v0d10v5__ags_diff_30 = '-1.35563e-04*hvn_saturation*hvn_saturation+9.24350e-03*hvn_saturation+1.58990e-02'
+ sky130_fd_pr__nfet_g5v0d10v5__ags_diff_31 = '-8.28750e-05*hvn_saturation*hvn_saturation+5.27850e-03*hvn_saturation+5.64400e-03'
+ sky130_fd_pr__nfet_g5v0d10v5__ags_diff_32 = '-5.62188e-05*hvn_saturation*hvn_saturation+1.86803e-03*hvn_saturation+1.98780e-03'
+ sky130_fd_pr__nfet_g5v0d10v5__ags_diff_4 = '-1.59031e-04*hvn_saturation*hvn_saturation+8.33962e-03*hvn_saturation+1.60720e-02'
+ sky130_fd_pr__nfet_g5v0d10v5__ags_diff_5 = '-5.76313e-05*hvn_saturation*hvn_saturation+6.67213e-03*hvn_saturation+9.26560e-03'
+ sky130_fd_pr__nfet_g5v0d10v5__ags_diff_7 = '-1.34756e-02*hvn_saturation*hvn_saturation+8.12613e-02*hvn_saturation+2.41410e-03'
+ sky130_fd_pr__nfet_g5v0d10v5__ags_diff_8 = '-1.60131e-04*hvn_saturation*hvn_saturation+1.10753e-02*hvn_saturation+1.77710e-03'
+ sky130_fd_pr__nfet_g5v0d10v5__ags_diff_9 = '3.00563e-05*hvn_saturation*hvn_saturation+1.52411e-02*hvn_saturation+9.50360e-03'
+ sky130_fd_pr__nfet_g5v0d10v5__ajunction_mult = '9.37500e-07*hvn_diode*hvn_diode+4.43837e-02*hvn_diode+9.95050e-01'
+ sky130_fd_pr__nfet_g5v0d10v5__b0_diff_35 = '2.77681e-09*hvn_saturation*hvn_saturation+-4.63263e-08*hvn_saturation+3.95160e-08'
+ sky130_fd_pr__nfet_g5v0d10v5__b0_diff_36 = '5.92463e-10*hvn_saturation*hvn_saturation+-1.28888e-08*hvn_saturation+-1.43040e-09'
+ sky130_fd_pr__nfet_g5v0d10v5__b0_diff_37 = '1.10325e-09*hvn_saturation*hvn_saturation+-2.22053e-08*hvn_saturation+-1.12960e-08'
+ sky130_fd_pr__nfet_g5v0d10v5__b0_diff_38 = '7.33937e-10*hvn_saturation*hvn_saturation+-1.33922e-08*hvn_saturation+-1.64620e-08'
+ sky130_fd_pr__nfet_g5v0d10v5__b0_diff_39 = '7.91794e-10*hvn_saturation*hvn_saturation+-1.07699e-08*hvn_saturation+1.65480e-09'
+ sky130_fd_pr__nfet_g5v0d10v5__b0_diff_43 = '2.80731e-09*hvn_saturation*hvn_saturation+-5.92512e-08*hvn_saturation+-3.10920e-08'
+ sky130_fd_pr__nfet_g5v0d10v5__b0_diff_44 = '1.12531e-09*hvn_saturation*hvn_saturation+-2.75295e-08*hvn_saturation+-7.73300e-09'
+ sky130_fd_pr__nfet_g5v0d10v5__b0_diff_45 = '1.12575e-09*hvn_saturation*hvn_saturation+-4.60225e-08*hvn_saturation+-4.24020e-08'
+ sky130_fd_pr__nfet_g5v0d10v5__b1_diff_35 = '9.75425e-11*hvn_saturation*hvn_saturation+1.13855e-09*hvn_saturation+5.72020e-10'
+ sky130_fd_pr__nfet_g5v0d10v5__b1_diff_36 = '6.29250e-11*hvn_saturation*hvn_saturation+-1.89400e-11*hvn_saturation+-6.57050e-10'
+ sky130_fd_pr__nfet_g5v0d10v5__b1_diff_37 = '-9.72500e-11*hvn_saturation*hvn_saturation+5.91875e-10*hvn_saturation+2.34120e-09'
+ sky130_fd_pr__nfet_g5v0d10v5__b1_diff_38 = '-7.46359e-11*hvn_saturation*hvn_saturation+5.44040e-10*hvn_saturation+-2.76660e-11'
+ sky130_fd_pr__nfet_g5v0d10v5__b1_diff_39 = '1.02879e-09*hvn_saturation*hvn_saturation+-4.22780e-09*hvn_saturation+3.47080e-10'
+ sky130_fd_pr__nfet_g5v0d10v5__b1_diff_43 = '7.27934e-11*hvn_saturation*hvn_saturation+-1.35581e-10*hvn_saturation+1.52480e-10'
+ sky130_fd_pr__nfet_g5v0d10v5__b1_diff_44 = '-3.24369e-11*hvn_saturation*hvn_saturation+1.00455e-10*hvn_saturation+7.14180e-10'
+ sky130_fd_pr__nfet_g5v0d10v5__b1_diff_45 = '-3.56531e-12*hvn_saturation*hvn_saturation+1.11429e-10*hvn_saturation+3.42160e-10'
+ sky130_fd_pr__nfet_g5v0d10v5__dlc_diff = '-4.33125e-09*poly_cd'
+ sky130_fd_pr__nfet_g5v0d10v5__dwc_diff = '8.04375e-09*diff_cd'
+ sky130_fd_pr__nfet_g5v0d10v5__k2_diff_0 = '7.47250e-05*hvn_bodyeffect*hvn_bodyeffect+-2.81925e-04*hvn_bodyeffect+-4.06730e-03'
+ sky130_fd_pr__nfet_g5v0d10v5__k2_diff_1 = '7.09375e-06*hvn_bodyeffect*hvn_bodyeffect+-5.62800e-04*hvn_bodyeffect+4.13810e-03'
+ sky130_fd_pr__nfet_g5v0d10v5__k2_diff_10 = '-3.25000e-06*hvn_bodyeffect*hvn_bodyeffect+3.78250e-04*hvn_bodyeffect+-1.17680e-02'
+ sky130_fd_pr__nfet_g5v0d10v5__k2_diff_11 = '9.21187e-05*hvn_bodyeffect*hvn_bodyeffect+-1.20142e-03*hvn_bodyeffect+5.75240e-03'
+ sky130_fd_pr__nfet_g5v0d10v5__k2_diff_12 = '1.98603e-05*hvn_bodyeffect*hvn_bodyeffect+-1.38954e-04*hvn_bodyeffect+-5.84930e-04'
+ sky130_fd_pr__nfet_g5v0d10v5__k2_diff_13 = '4.15625e-06*hvn_bodyeffect*hvn_bodyeffect+-7.95750e-05*hvn_bodyeffect+-4.00790e-03'
+ sky130_fd_pr__nfet_g5v0d10v5__k2_diff_14 = '5.90000e-06*hvn_bodyeffect*hvn_bodyeffect+-4.82875e-04*hvn_bodyeffect+3.89160e-03'
+ sky130_fd_pr__nfet_g5v0d10v5__k2_diff_15 = '5.16031e-05*hvn_bodyeffect*hvn_bodyeffect+5.98913e-04*hvn_bodyeffect+-5.04340e-03'
+ sky130_fd_pr__nfet_g5v0d10v5__k2_diff_16 = '8.15625e-06*hvn_bodyeffect*hvn_bodyeffect+-5.96375e-04*hvn_bodyeffect+-5.48090e-03'
+ sky130_fd_pr__nfet_g5v0d10v5__k2_diff_17 = '5.28125e-06*hvn_bodyeffect*hvn_bodyeffect+-3.89875e-04*hvn_bodyeffect+-1.39660e-02'
+ sky130_fd_pr__nfet_g5v0d10v5__k2_diff_18 = '5.40625e-06*hvn_bodyeffect*hvn_bodyeffect+-3.72375e-04*hvn_bodyeffect+-1.85650e-02'
+ sky130_fd_pr__nfet_g5v0d10v5__k2_diff_19 = '3.78125e-06*hvn_bodyeffect*hvn_bodyeffect+-2.39875e-04*hvn_bodyeffect+-2.02800e-02'
+ sky130_fd_pr__nfet_g5v0d10v5__k2_diff_2 = '1.02894e-04*hvn_bodyeffect*hvn_bodyeffect+-1.09700e-04*hvn_bodyeffect+-4.62100e-03'
+ sky130_fd_pr__nfet_g5v0d10v5__k2_diff_20 = '7.74563e-05*hvn_bodyeffect*hvn_bodyeffect+-3.08350e-04*hvn_bodyeffect+-1.15350e-03'
+ sky130_fd_pr__nfet_g5v0d10v5__k2_diff_21 = '1.55562e-05*hvn_bodyeffect*hvn_bodyeffect+5.81250e-05*hvn_bodyeffect+-4.25180e-03'
+ sky130_fd_pr__nfet_g5v0d10v5__k2_diff_22 = '8.95312e-06*hvn_bodyeffect*hvn_bodyeffect+-6.68037e-04*hvn_bodyeffect+5.08750e-03'
+ sky130_fd_pr__nfet_g5v0d10v5__k2_diff_23 = '5.33125e-06*hvn_bodyeffect*hvn_bodyeffect+-4.05875e-04*hvn_bodyeffect+-4.77300e-03'
+ sky130_fd_pr__nfet_g5v0d10v5__k2_diff_24 = '8.30000e-06*hvn_bodyeffect*hvn_bodyeffect+-5.66175e-04*hvn_bodyeffect+-9.10710e-03'
+ sky130_fd_pr__nfet_g5v0d10v5__k2_diff_25 = '3.36250e-06*hvn_bodyeffect*hvn_bodyeffect+-2.16700e-04*hvn_bodyeffect+-1.07550e-02'
+ sky130_fd_pr__nfet_g5v0d10v5__k2_diff_26 = '4.41250e-05*hvn_bodyeffect*hvn_bodyeffect+9.23325e-04*hvn_bodyeffect+-2.55850e-03'
+ sky130_fd_pr__nfet_g5v0d10v5__k2_diff_27 = '3.25125e-05*hvn_bodyeffect*hvn_bodyeffect+-5.72250e-05*hvn_bodyeffect+2.83010e-03'
+ sky130_fd_pr__nfet_g5v0d10v5__k2_diff_28 = '2.19844e-05*hvn_bodyeffect*hvn_bodyeffect+-6.95262e-04*hvn_bodyeffect+7.47220e-03'
+ sky130_fd_pr__nfet_g5v0d10v5__k2_diff_29 = '5.25000e-06*hvn_bodyeffect*hvn_bodyeffect+-4.04075e-04*hvn_bodyeffect+5.16790e-03'
+ sky130_fd_pr__nfet_g5v0d10v5__k2_diff_3 = '3.60938e-06*hvn_bodyeffect*hvn_bodyeffect+-2.31688e-04*hvn_bodyeffect+-3.45700e-03'
+ sky130_fd_pr__nfet_g5v0d10v5__k2_diff_30 = '3.67813e-06*hvn_bodyeffect*hvn_bodyeffect+-3.17788e-04*hvn_bodyeffect+-4.45540e-03'
+ sky130_fd_pr__nfet_g5v0d10v5__k2_diff_31 = '3.52500e-06*hvn_bodyeffect*hvn_bodyeffect+-2.53775e-04*hvn_bodyeffect+-9.10030e-03'
+ sky130_fd_pr__nfet_g5v0d10v5__k2_diff_32 = '4.09063e-06*hvn_bodyeffect*hvn_bodyeffect+-2.91113e-04*hvn_bodyeffect+-1.04880e-02'
+ sky130_fd_pr__nfet_g5v0d10v5__k2_diff_33 = '6.44478e-05*hvn_bodyeffect*hvn_bodyeffect+5.09866e-04*hvn_bodyeffect+-3.90410e-03'
+ sky130_fd_pr__nfet_g5v0d10v5__k2_diff_34 = '8.86875e-06*hvn_bodyeffect*hvn_bodyeffect+-5.74000e-04*hvn_bodyeffect+7.24290e-03'
+ sky130_fd_pr__nfet_g5v0d10v5__k2_diff_35 = '-5.02500e-06*hvn_bodyeffect*hvn_bodyeffect+2.15860e-03*hvn_bodyeffect+-4.43320e-03'
+ sky130_fd_pr__nfet_g5v0d10v5__k2_diff_36 = '-1.07625e-05*hvn_bodyeffect*hvn_bodyeffect+2.51013e-03*hvn_bodyeffect+-7.64730e-03'
+ sky130_fd_pr__nfet_g5v0d10v5__k2_diff_37 = '-4.45313e-05*hvn_bodyeffect*hvn_bodyeffect+3.21803e-03*hvn_bodyeffect+-6.06140e-03'
+ sky130_fd_pr__nfet_g5v0d10v5__k2_diff_38 = '-1.31469e-05*hvn_bodyeffect*hvn_bodyeffect+2.66701e-03*hvn_bodyeffect+-5.27760e-03'
+ sky130_fd_pr__nfet_g5v0d10v5__k2_diff_39 = '-1.76688e-05*hvn_bodyeffect*hvn_bodyeffect+2.95490e-03*hvn_bodyeffect+-8.06770e-03'
+ sky130_fd_pr__nfet_g5v0d10v5__k2_diff_4 = '9.68750e-07*hvn_bodyeffect*hvn_bodyeffect+-7.36250e-05*hvn_bodyeffect+-1.26690e-02'
+ sky130_fd_pr__nfet_g5v0d10v5__k2_diff_40 = '1.02106e-04*hvn_bodyeffect*hvn_bodyeffect+-4.77350e-05*hvn_bodyeffect+-6.53330e-04'
+ sky130_fd_pr__nfet_g5v0d10v5__k2_diff_41 = '1.08906e-05*hvn_bodyeffect*hvn_bodyeffect+2.39024e-03*hvn_bodyeffect+-6.55530e-03'
+ sky130_fd_pr__nfet_g5v0d10v5__k2_diff_42 = '-1.48750e-05*hvn_bodyeffect*hvn_bodyeffect+3.01000e-03*hvn_bodyeffect+-1.06280e-02'
+ sky130_fd_pr__nfet_g5v0d10v5__k2_diff_43 = '4.37500e-07*hvn_bodyeffect*hvn_bodyeffect+3.07425e-04*hvn_bodyeffect+-2.38730e-03'
+ sky130_fd_pr__nfet_g5v0d10v5__k2_diff_44 = '-9.61563e-06*hvn_bodyeffect*hvn_bodyeffect+9.61763e-04*hvn_bodyeffect+-9.15210e-03'
+ sky130_fd_pr__nfet_g5v0d10v5__k2_diff_45 = '-1.73750e-05*hvn_bodyeffect*hvn_bodyeffect+1.17925e-03*hvn_bodyeffect+-1.30790e-02'
+ sky130_fd_pr__nfet_g5v0d10v5__k2_diff_46 = '9.30331e-05*hvn_bodyeffect*hvn_bodyeffect+-7.46963e-04*hvn_bodyeffect+-9.03280e-04'
+ sky130_fd_pr__nfet_g5v0d10v5__k2_diff_47 = '3.98438e-07*hvn_bodyeffect*hvn_bodyeffect+3.53151e-04*hvn_bodyeffect+5.47120e-04'
+ sky130_fd_pr__nfet_g5v0d10v5__k2_diff_48 = '1.36953e-05*hvn_bodyeffect*hvn_bodyeffect+5.07219e-04*hvn_bodyeffect+1.86390e-03'
+ sky130_fd_pr__nfet_g5v0d10v5__k2_diff_5 = '2.65625e-06*hvn_bodyeffect*hvn_bodyeffect+-1.58375e-04*hvn_bodyeffect+-1.64010e-02'
+ sky130_fd_pr__nfet_g5v0d10v5__k2_diff_6 = '9.01237e-05*hvn_bodyeffect*hvn_bodyeffect+-1.12295e-03*hvn_bodyeffect+2.69350e-03'
+ sky130_fd_pr__nfet_g5v0d10v5__k2_diff_7 = '-4.52750e-05*hvn_bodyeffect*hvn_bodyeffect+4.53250e-05*hvn_bodyeffect+6.64270e-03'
+ sky130_fd_pr__nfet_g5v0d10v5__k2_diff_8 = '-6.62500e-06*hvn_bodyeffect*hvn_bodyeffect+4.94500e-04*hvn_bodyeffect+-1.60860e-02'
+ sky130_fd_pr__nfet_g5v0d10v5__k2_diff_9 = '-5.68438e-06*hvn_bodyeffect*hvn_bodyeffect+4.10037e-04*hvn_bodyeffect+-9.78190e-03'
+ sky130_fd_pr__nfet_g5v0d10v5__lint_diff = '-4.33125e-09*poly_cd'
+ sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_0 = '-2.89969e-04*hvn_subvt*hvn_subvt+4.64249e-02*hvn_subvt+2.08090e-01'
+ sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_1 = '-9.71875e-05*hvn_subvt*hvn_subvt+1.53863e-02*hvn_subvt+2.88340e-01'
+ sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_10 = '6.20312e-04*hvn_subvt*hvn_subvt+-1.79287e-02*hvn_subvt+5.42610e-01'
+ sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_11 = '7.18438e-04*hvn_subvt*hvn_subvt+-5.21838e-02*hvn_subvt+5.07110e-01'
+ sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_12 = '6.93438e-04*hvn_subvt*hvn_subvt+-4.23913e-02*hvn_subvt+4.56740e-01'
+ sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_13 = '5.26563e-04*hvn_subvt*hvn_subvt+-1.54587e-02*hvn_subvt+4.51360e-01'
+ sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_14 = '-8.46875e-05*hvn_subvt*hvn_subvt+1.62163e-02*hvn_subvt+2.87850e-01'
+ sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_15 = '-2.22500e-04*hvn_subvt*hvn_subvt+5.97250e-02*hvn_subvt+1.69520e-01'
+ sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_16 = '5.90625e-05*hvn_subvt*hvn_subvt+4.44375e-03*hvn_subvt+3.34880e-01'
+ sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_17 = '-6.09375e-05*hvn_subvt*hvn_subvt+1.14962e-02*hvn_subvt+3.52290e-01'
+ sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_18 = '7.31250e-05*hvn_subvt*hvn_subvt+1.32000e-03*hvn_subvt+3.95460e-01'
+ sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_19 = '1.93750e-05*hvn_subvt*hvn_subvt+5.36500e-03*hvn_subvt+4.49450e-01'
+ sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_2 = '-1.18237e-03*hvn_subvt*hvn_subvt+4.17620e-02*hvn_subvt+1.98860e-01'
+ sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_20 = '3.35313e-04*hvn_subvt*hvn_subvt+-2.04138e-02*hvn_subvt+3.28460e-01'
+ sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_21 = '2.19063e-04*hvn_subvt*hvn_subvt+-1.74375e-03*hvn_subvt+2.96770e-01'
+ sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_22 = '-6.87500e-05*hvn_subvt*hvn_subvt+1.18250e-02*hvn_subvt+3.00100e-01'
+ sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_23 = '-2.15625e-05*hvn_subvt*hvn_subvt+6.50875e-03*hvn_subvt+3.43330e-01'
+ sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_24 = '1.34375e-05*hvn_subvt*hvn_subvt+3.96625e-03*hvn_subvt+3.87060e-01'
+ sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_25 = '-3.28125e-05*hvn_subvt*hvn_subvt+8.54375e-03*hvn_subvt+4.46960e-01'
+ sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_26 = '1.34688e-04*hvn_subvt*hvn_subvt+-7.56250e-04*hvn_subvt+2.60880e-01'
+ sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_27 = '-2.63125e-04*hvn_subvt*hvn_subvt+1.16250e-03*hvn_subvt+2.72160e-01'
+ sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_28 = '-1.81875e-04*hvn_subvt*hvn_subvt+1.18650e-02*hvn_subvt+2.97170e-01'
+ sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_29 = '-5.87500e-05*hvn_subvt*hvn_subvt+1.01925e-02*hvn_subvt+2.85520e-01'
+ sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_3 = '3.04375e-04*hvn_subvt*hvn_subvt+-1.04175e-02*hvn_subvt+4.05030e-01'
+ sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_30 = '-1.25000e-05*hvn_subvt*hvn_subvt+6.63500e-03*hvn_subvt+3.27400e-01'
+ sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_31 = '-3.56250e-05*hvn_subvt*hvn_subvt+7.74250e-03*hvn_subvt+3.75610e-01'
+ sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_32 = '-5.18750e-05*hvn_subvt*hvn_subvt+9.95500e-03*hvn_subvt+4.24180e-01'
+ sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_33 = '-1.48437e-04*hvn_subvt*hvn_subvt+3.00262e-02*hvn_subvt+2.29790e-01'
+ sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_34 = '-1.43750e-05*hvn_subvt*hvn_subvt+1.14125e-02*hvn_subvt+2.80640e-01'
+ sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_35 = '7.68438e-04*hvn_subvt*hvn_subvt+3.44137e-02*hvn_subvt+4.49640e-01'
+ sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_36 = '2.71562e-03*hvn_subvt*hvn_subvt+-4.52125e-02*hvn_subvt+7.29180e-01'
+ sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_37 = '1.67469e-03*hvn_subvt*hvn_subvt+7.47125e-03*hvn_subvt+4.85030e-01'
+ sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_38 = '8.69375e-04*hvn_subvt*hvn_subvt+4.58750e-03*hvn_subvt+5.45160e-01'
+ sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_39 = '1.67531e-03*hvn_subvt*hvn_subvt+-2.09238e-02*hvn_subvt+6.18840e-01'
+ sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_4 = '1.77500e-04*hvn_subvt*hvn_subvt+-2.18500e-03*hvn_subvt+4.09770e-01'
+ sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_40 = '1.39312e-03*hvn_subvt*hvn_subvt+-2.41550e-02*hvn_subvt+5.08070e-01'
+ sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_41 = '1.42625e-03*hvn_subvt*hvn_subvt+-4.97500e-04*hvn_subvt+4.47840e-01'
+ sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_42 = '1.58781e-03*hvn_subvt*hvn_subvt+1.46187e-02*hvn_subvt+4.67940e-01'
+ sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_43 = '5.31250e-04*hvn_subvt*hvn_subvt+-7.13250e-03*hvn_subvt+4.67470e-01'
+ sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_44 = '4.79687e-04*hvn_subvt*hvn_subvt+-2.84375e-03*hvn_subvt+4.92520e-01'
+ sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_45 = '6.41563e-04*hvn_subvt*hvn_subvt+-1.74763e-02*hvn_subvt+5.27920e-01'
+ sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_46 = '5.97188e-04*hvn_subvt*hvn_subvt+-3.66163e-02*hvn_subvt+5.26700e-01'
+ sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_47 = '7.61563e-04*hvn_subvt*hvn_subvt+-2.75288e-02*hvn_subvt+4.83060e-01'
+ sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_48 = '9.12812e-04*hvn_subvt*hvn_subvt+-4.68262e-02*hvn_subvt+5.03590e-01'
+ sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_5 = '2.91562e-04*hvn_subvt*hvn_subvt+-1.13687e-02*hvn_subvt+4.43440e-01'
+ sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_6 = '5.48125e-04*hvn_subvt*hvn_subvt+-3.87775e-02*hvn_subvt+4.66140e-01'
+ sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_7 = '7.56875e-04*hvn_subvt*hvn_subvt+-1.52300e-02*hvn_subvt+4.40780e-01'
+ sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_8 = '4.17187e-04*hvn_subvt*hvn_subvt+-1.34262e-02*hvn_subvt+4.50850e-01'
+ sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_9 = '3.82813e-04*hvn_subvt*hvn_subvt+-5.41375e-03*hvn_subvt+4.75000e-01'
+ sky130_fd_pr__nfet_g5v0d10v5__overlap_mult = '2.36250e-04*hvtox*hvtox+3.48425e-02*hvtox+8.98050e-01'
+ sky130_fd_pr__nfet_g5v0d10v5__pjunction_mult = '1.87500e-06*hvn_diode*hvn_diode+5.91425e-02*hvn_diode+1.01440e+00'
+ sky130_fd_pr__rf_nfet_g5v0d10v5_b__ajunction_mult = '9.37500e-07*hvn_diode*hvn_diode+4.43837e-02*hvn_diode+9.95050e-01'
+ sky130_fd_pr__rf_nfet_g5v0d10v5_b__dlc_diff = '-4.33125e-09*poly_cd'
+ sky130_fd_pr__rf_nfet_g5v0d10v5_b__lint_diff = '-4.33125e-09*poly_cd'
+ sky130_fd_pr__rf_nfet_g5v0d10v5_b__overlap_mult = '2.36250e-04*hvtox*hvtox+3.48425e-02*hvtox+8.98050e-01'
+ sky130_fd_pr__rf_nfet_g5v0d10v5_b__pjunction_mult = '1.87500e-06*hvn_diode*hvn_diode+5.91425e-02*hvn_diode+1.01440e+00'
+ sky130_fd_pr__rf_nfet_g5v0d10v5_b__rbpb_mult = '5.00000e-02*hvn_bodyeffect+1.00000e+00'
+ sky130_fd_pr__rf_nfet_g5v0d10v5_b__rshg_diff = '1.75000e+00*ic_res'
+ sky130_fd_pr__rf_nfet_g5v0d10v5_b__toxe_mult = '1.50000e-02*hvtox+1.00000e+00'
+ sky130_fd_pr__rf_nfet_g5v0d10v5_b__wint_diff = '8.04375e-09*diff_cd'
+ sky130_fd_pr__rf_nfet_g5v0d10v5_b__xgw_diff = '1.60625e-08*diff_cd'
+ sky130_fd_pr__rf_nfet_g5v0d10v5_bM10__k2_diff_0 = '6.73731e-05*hvn_bodyeffect*hvn_bodyeffect+1.44721e-03*hvn_bodyeffect+5.94980e-04'
+ sky130_fd_pr__rf_nfet_g5v0d10v5_bM10__k2_diff_1 = '4.82875e-05*hvn_bodyeffect*hvn_bodyeffect+2.60342e-03*hvn_bodyeffect+-6.80590e-03'
+ sky130_fd_pr__rf_nfet_g5v0d10v5_bM10__k2_diff_2 = '5.88812e-05*hvn_bodyeffect*hvn_bodyeffect+1.91960e-03*hvn_bodyeffect+-1.71730e-03'
+ sky130_fd_pr__rf_nfet_g5v0d10v5_bM10__u0_diff_0 = '-7.68594e-05*hvn_mobility*hvn_mobility+1.74013e-04*hvn_mobility+-1.64490e-03'
+ sky130_fd_pr__rf_nfet_g5v0d10v5_bM10__u0_diff_1 = '-6.29875e-05*hvn_mobility*hvn_mobility+3.40150e-04*hvn_mobility+-2.93900e-03'
+ sky130_fd_pr__rf_nfet_g5v0d10v5_bM10__u0_diff_2 = '-1.05841e-04*hvn_mobility*hvn_mobility+-8.23638e-04*hvn_mobility+-4.10540e-03'
+ sky130_fd_pr__rf_nfet_g5v0d10v5_bM10__vsat_diff_0 = '-1.58063e+01*hvn_saturation*hvn_saturation+2.77575e+03*hvn_saturation+1.10090e+03'
+ sky130_fd_pr__rf_nfet_g5v0d10v5_bM10__vsat_diff_1 = '-1.25478e+02*hvn_saturation*hvn_saturation+1.14561e+03*hvn_saturation+-3.86290e+03'
+ sky130_fd_pr__rf_nfet_g5v0d10v5_bM10__vsat_diff_2 = '1.89456e+02*hvn_saturation*hvn_saturation+3.27588e+03*hvn_saturation+-5.55680e+03'
+ sky130_fd_pr__rf_nfet_g5v0d10v5_bM10__vth0_diff_0 = '-1.66438e-04*hvn_threshold*hvn_threshold+1.97085e-02*hvn_threshold+-1.50750e-02'
+ sky130_fd_pr__rf_nfet_g5v0d10v5_bM10__vth0_diff_1 = '-1.62219e-04*hvn_threshold*hvn_threshold+1.69419e-02*hvn_threshold+-1.26710e-02'
+ sky130_fd_pr__rf_nfet_g5v0d10v5_bM10__vth0_diff_2 = '-1.69625e-04*hvn_threshold*hvn_threshold+1.76940e-02*hvn_threshold+-2.21230e-02'
+ sky130_fd_pr__rf_nfet_g5v0d10v5_bM02__k2_diff_0 = '6.49969e-05*hvn_bodyeffect*hvn_bodyeffect+1.48076e-03*hvn_bodyeffect+1.31270e-03'
+ sky130_fd_pr__rf_nfet_g5v0d10v5_bM02__k2_diff_1 = '4.33569e-05*hvn_bodyeffect*hvn_bodyeffect+2.97512e-03*hvn_bodyeffect+-5.34210e-04'
+ sky130_fd_pr__rf_nfet_g5v0d10v5_bM02__u0_diff_0 = '-7.58844e-05*hvn_mobility*hvn_mobility+2.36187e-04*hvn_mobility+-2.96850e-03'
+ sky130_fd_pr__rf_nfet_g5v0d10v5_bM02__u0_diff_1 = '-5.67477e-05*hvn_mobility*hvn_mobility+5.00359e-04*hvn_mobility+-1.01150e-03'
+ sky130_fd_pr__rf_nfet_g5v0d10v5_bM02__vsat_diff_0 = '-1.05934e+02*hvn_saturation*hvn_saturation+1.86891e+03*hvn_saturation+-3.50340e+03'
+ sky130_fd_pr__rf_nfet_g5v0d10v5_bM02__vsat_diff_1 = '-1.37866e+02*hvn_saturation*hvn_saturation+1.07262e+03*hvn_saturation+3.23350e+02'
+ sky130_fd_pr__rf_nfet_g5v0d10v5_bM02__vth0_diff_0 = '-1.63406e-04*hvn_threshold*hvn_threshold+1.97464e-02*hvn_threshold+-1.52620e-02'
+ sky130_fd_pr__rf_nfet_g5v0d10v5_bM02__vth0_diff_1 = '-1.63219e-04*hvn_threshold*hvn_threshold+1.69772e-02*hvn_threshold+-2.53650e-03'
+ sky130_fd_pr__rf_nfet_g5v0d10v5_bM04__k2_diff_0 = '6.42844e-05*hvn_bodyeffect*hvn_bodyeffect+1.50469e-03*hvn_bodyeffect+1.01730e-03'
+ sky130_fd_pr__rf_nfet_g5v0d10v5_bM04__k2_diff_1 = '4.41862e-05*hvn_bodyeffect*hvn_bodyeffect+2.84487e-03*hvn_bodyeffect+-5.78480e-04'
+ sky130_fd_pr__rf_nfet_g5v0d10v5_bM04__k2_diff_2 = '5.32719e-05*hvn_bodyeffect*hvn_bodyeffect+2.20489e-03*hvn_bodyeffect+-1.51370e-03'
+ sky130_fd_pr__rf_nfet_g5v0d10v5_bM04__u0_diff_0 = '-7.63000e-05*hvn_mobility*hvn_mobility+2.03675e-04*hvn_mobility+-3.12710e-03'
+ sky130_fd_pr__rf_nfet_g5v0d10v5_bM04__u0_diff_1 = '-5.58209e-05*hvn_mobility*hvn_mobility+4.70666e-04*hvn_mobility+-1.39930e-03'
+ sky130_fd_pr__rf_nfet_g5v0d10v5_bM04__u0_diff_2 = '-6.19250e-05*hvn_mobility*hvn_mobility+3.00125e-04*hvn_mobility+-3.00200e-03'
+ sky130_fd_pr__rf_nfet_g5v0d10v5_bM04__vsat_diff_0 = '-8.86719e+01*hvn_saturation*hvn_saturation+1.90121e+03*hvn_saturation+-3.94640e+03'
+ sky130_fd_pr__rf_nfet_g5v0d10v5_bM04__vsat_diff_1 = '-1.36300e+02*hvn_saturation*hvn_saturation+1.00510e+03*hvn_saturation+-1.84170e+03'
+ sky130_fd_pr__rf_nfet_g5v0d10v5_bM04__vsat_diff_2 = '-1.28133e+02*hvn_saturation*hvn_saturation+1.10697e+03*hvn_saturation+-2.99490e+03'
+ sky130_fd_pr__rf_nfet_g5v0d10v5_bM04__vth0_diff_0 = '-1.63094e-04*hvn_threshold*hvn_threshold+1.96286e-02*hvn_threshold+-2.45260e-02'
+ sky130_fd_pr__rf_nfet_g5v0d10v5_bM04__vth0_diff_1 = '-1.60731e-04*hvn_threshold*hvn_threshold+1.69806e-02*hvn_threshold+-9.99980e-03'
+ sky130_fd_pr__rf_nfet_g5v0d10v5_bM04__vth0_diff_2 = '-1.61125e-04*hvn_threshold*hvn_threshold+1.79651e-02*hvn_threshold+-8.21650e-03'
+ sky130_fd_pr__nfet_g5v0d10v5__toxe_mult = '1.50000e-02*hvtox+1.00000e+00'
+ sky130_fd_pr__nfet_g5v0d10v5__u0_diff_0 = '-8.24500e-06*hvn_mobility*hvn_mobility+9.28155e-04*hvn_mobility+4.51800e-03'
+ sky130_fd_pr__nfet_g5v0d10v5__u0_diff_1 = '-1.04884e-05*hvn_mobility*hvn_mobility+3.44494e-04*hvn_mobility+8.19840e-04'
+ sky130_fd_pr__nfet_g5v0d10v5__u0_diff_10 = '-2.09728e-05*hvn_mobility*hvn_mobility+-1.26125e-06*hvn_mobility+-3.02860e-04'
+ sky130_fd_pr__nfet_g5v0d10v5__u0_diff_11 = '-5.71222e-05*hvn_mobility*hvn_mobility+2.79756e-04*hvn_mobility+5.01580e-04'
+ sky130_fd_pr__nfet_g5v0d10v5__u0_diff_12 = '-4.13425e-05*hvn_mobility*hvn_mobility+2.83733e-04*hvn_mobility+9.96050e-04'
+ sky130_fd_pr__nfet_g5v0d10v5__u0_diff_13 = '-4.42587e-05*hvn_mobility*hvn_mobility+-4.03625e-05*hvn_mobility+-5.64110e-04'
+ sky130_fd_pr__nfet_g5v0d10v5__u0_diff_14 = '-1.08125e-05*hvn_mobility*hvn_mobility+3.17375e-04*hvn_mobility+1.07100e-03'
+ sky130_fd_pr__nfet_g5v0d10v5__u0_diff_15 = '1.26447e-04*hvn_mobility*hvn_mobility+1.85454e-03*hvn_mobility+4.21570e-03'
+ sky130_fd_pr__nfet_g5v0d10v5__u0_diff_16 = '-1.46031e-05*hvn_mobility*hvn_mobility+3.61638e-04*hvn_mobility+-1.05750e-03'
+ sky130_fd_pr__nfet_g5v0d10v5__u0_diff_17 = '-9.52375e-06*hvn_mobility*hvn_mobility+3.20463e-04*hvn_mobility+-7.02670e-04'
+ sky130_fd_pr__nfet_g5v0d10v5__u0_diff_18 = '-9.49000e-06*hvn_mobility*hvn_mobility+2.19832e-04*hvn_mobility+-9.12430e-04'
+ sky130_fd_pr__nfet_g5v0d10v5__u0_diff_19 = '-1.24641e-05*hvn_mobility*hvn_mobility+8.79613e-05*hvn_mobility+-9.95730e-04'
+ sky130_fd_pr__nfet_g5v0d10v5__u0_diff_2 = '5.92500e-06*hvn_mobility*hvn_mobility+9.91450e-04*hvn_mobility+5.75260e-03'
+ sky130_fd_pr__nfet_g5v0d10v5__u0_diff_20 = '-3.45594e-05*hvn_mobility*hvn_mobility+5.85712e-04*hvn_mobility+2.04650e-03'
+ sky130_fd_pr__nfet_g5v0d10v5__u0_diff_21 = '-3.88516e-05*hvn_mobility*hvn_mobility+1.89781e-04*hvn_mobility+1.23160e-03'
+ sky130_fd_pr__nfet_g5v0d10v5__u0_diff_22 = '-1.19396e-05*hvn_mobility*hvn_mobility+4.28525e-04*hvn_mobility+4.72330e-05'
+ sky130_fd_pr__nfet_g5v0d10v5__u0_diff_23 = '-9.17781e-06*hvn_mobility*hvn_mobility+3.17489e-04*hvn_mobility+-1.66270e-03'
+ sky130_fd_pr__nfet_g5v0d10v5__u0_diff_24 = '-9.35938e-06*hvn_mobility*hvn_mobility+2.08013e-04*hvn_mobility+-2.15460e-03'
+ sky130_fd_pr__nfet_g5v0d10v5__u0_diff_25 = '-1.26000e-05*hvn_mobility*hvn_mobility+3.56750e-05*hvn_mobility+-2.49750e-03'
+ sky130_fd_pr__nfet_g5v0d10v5__u0_diff_26 = '-2.76486e-05*hvn_mobility*hvn_mobility+7.50544e-04*hvn_mobility+3.40790e-03'
+ sky130_fd_pr__nfet_g5v0d10v5__u0_diff_27 = '-3.36691e-05*hvn_mobility*hvn_mobility+2.37101e-04*hvn_mobility+1.79980e-03'
+ sky130_fd_pr__nfet_g5v0d10v5__u0_diff_28 = '-1.17908e-04*hvn_mobility*hvn_mobility+-8.22875e-05*hvn_mobility+1.58670e-04'
+ sky130_fd_pr__nfet_g5v0d10v5__u0_diff_29 = '-1.16491e-05*hvn_mobility*hvn_mobility+4.16404e-04*hvn_mobility+-1.24220e-03'
+ sky130_fd_pr__nfet_g5v0d10v5__u0_diff_3 = '-2.31438e-05*hvn_mobility*hvn_mobility+2.19200e-04*hvn_mobility+-1.89060e-03'
+ sky130_fd_pr__nfet_g5v0d10v5__u0_diff_30 = '-7.79375e-06*hvn_mobility*hvn_mobility+3.19525e-04*hvn_mobility+-2.41470e-03'
+ sky130_fd_pr__nfet_g5v0d10v5__u0_diff_31 = '-9.29375e-06*hvn_mobility*hvn_mobility+1.95600e-04*hvn_mobility+-2.32500e-03'
+ sky130_fd_pr__nfet_g5v0d10v5__u0_diff_32 = '-1.27250e-05*hvn_mobility*hvn_mobility+1.20250e-05*hvn_mobility+-2.89780e-03'
+ sky130_fd_pr__nfet_g5v0d10v5__u0_diff_33 = '-3.05922e-05*hvn_mobility*hvn_mobility+6.93119e-04*hvn_mobility+4.02960e-03'
+ sky130_fd_pr__nfet_g5v0d10v5__u0_diff_34 = '-1.71832e-05*hvn_mobility*hvn_mobility+3.45517e-04*hvn_mobility+-1.14770e-03'
+ sky130_fd_pr__nfet_g5v0d10v5__u0_diff_35 = '-8.34531e-05*hvn_mobility*hvn_mobility+-2.59062e-04*hvn_mobility+-3.15800e-03'
+ sky130_fd_pr__nfet_g5v0d10v5__u0_diff_36 = '-3.90187e-05*hvn_mobility*hvn_mobility+-1.26000e-05*hvn_mobility+-3.20110e-03'
+ sky130_fd_pr__nfet_g5v0d10v5__u0_diff_37 = '-6.98906e-05*hvn_mobility*hvn_mobility+-3.57612e-04*hvn_mobility+-2.98380e-03'
+ sky130_fd_pr__nfet_g5v0d10v5__u0_diff_38 = '-2.93594e-05*hvn_mobility*hvn_mobility+1.86038e-04*hvn_mobility+-2.98950e-03'
+ sky130_fd_pr__nfet_g5v0d10v5__u0_diff_39 = '-2.84500e-05*hvn_mobility*hvn_mobility+1.21850e-04*hvn_mobility+-3.23850e-03'
+ sky130_fd_pr__nfet_g5v0d10v5__u0_diff_4 = '-1.34703e-05*hvn_mobility*hvn_mobility+2.64119e-04*hvn_mobility+-1.30030e-03'
+ sky130_fd_pr__nfet_g5v0d10v5__u0_diff_40 = '-1.27712e-04*hvn_mobility*hvn_mobility+-1.01025e-04*hvn_mobility+-1.08410e-03'
+ sky130_fd_pr__nfet_g5v0d10v5__u0_diff_41 = '-1.51431e-04*hvn_mobility*hvn_mobility+-6.57925e-04*hvn_mobility+-2.79320e-03'
+ sky130_fd_pr__nfet_g5v0d10v5__u0_diff_42 = '-1.29638e-04*hvn_mobility*hvn_mobility+-7.43375e-04*hvn_mobility+-3.05680e-03'
+ sky130_fd_pr__nfet_g5v0d10v5__u0_diff_43 = '-4.69281e-05*hvn_mobility*hvn_mobility+-1.12813e-04*hvn_mobility+-1.20260e-03'
+ sky130_fd_pr__nfet_g5v0d10v5__u0_diff_44 = '-3.64169e-05*hvn_mobility*hvn_mobility+-1.27200e-04*hvn_mobility+-9.53130e-04'
+ sky130_fd_pr__nfet_g5v0d10v5__u0_diff_45 = '-1.26812e-05*hvn_mobility*hvn_mobility+2.27873e-04*hvn_mobility+-9.37710e-04'
+ sky130_fd_pr__nfet_g5v0d10v5__u0_diff_46 = '-7.45319e-05*hvn_mobility*hvn_mobility+4.15575e-05*hvn_mobility+2.01740e-04'
+ sky130_fd_pr__nfet_g5v0d10v5__u0_diff_47 = '-5.95500e-05*hvn_mobility*hvn_mobility+-2.03525e-04*hvn_mobility+-1.01860e-03'
+ sky130_fd_pr__nfet_g5v0d10v5__u0_diff_48 = '-6.66087e-05*hvn_mobility*hvn_mobility+3.55375e-05*hvn_mobility+-5.95410e-04'
+ sky130_fd_pr__nfet_g5v0d10v5__u0_diff_5 = '-1.20960e-05*hvn_mobility*hvn_mobility+1.98846e-04*hvn_mobility+-6.51780e-04'
+ sky130_fd_pr__nfet_g5v0d10v5__u0_diff_6 = '-4.61306e-05*hvn_mobility*hvn_mobility+4.04450e-04*hvn_mobility+5.68390e-04'
+ sky130_fd_pr__nfet_g5v0d10v5__u0_diff_7 = '-1.95196e-05*hvn_mobility*hvn_mobility+9.26537e-05*hvn_mobility+6.46980e-05'
+ sky130_fd_pr__nfet_g5v0d10v5__u0_diff_8 = '-2.48087e-05*hvn_mobility*hvn_mobility+4.47675e-05*hvn_mobility+-2.29840e-04'
+ sky130_fd_pr__nfet_g5v0d10v5__u0_diff_9 = '-9.14038e-06*hvn_mobility*hvn_mobility+2.66504e-04*hvn_mobility+-6.99390e-05'
+ sky130_fd_pr__nfet_g5v0d10v5__ua_diff_0 = '3.08034e-14*hvn_mobility*hvn_mobility+-7.00689e-13*hvn_mobility+-4.02290e-12'
+ sky130_fd_pr__nfet_g5v0d10v5__ua_diff_1 = '1.07072e-13*hvn_mobility*hvn_mobility+1.39237e-13*hvn_mobility+-4.08070e-12'
+ sky130_fd_pr__nfet_g5v0d10v5__ua_diff_10 = '3.56969e-14*hvn_mobility*hvn_mobility+2.05062e-13*hvn_mobility+1.31660e-12'
+ sky130_fd_pr__nfet_g5v0d10v5__ua_diff_11 = '2.69375e-13*hvn_mobility*hvn_mobility+-4.34750e-13*hvn_mobility+1.02950e-11'
+ sky130_fd_pr__nfet_g5v0d10v5__ua_diff_12 = '1.75116e-13*hvn_mobility*hvn_mobility+6.83437e-13*hvn_mobility+5.67640e-12'
+ sky130_fd_pr__nfet_g5v0d10v5__ua_diff_13 = '1.06450e-13*hvn_mobility*hvn_mobility+4.85700e-13*hvn_mobility+5.70160e-12'
+ sky130_fd_pr__nfet_g5v0d10v5__ua_diff_14 = '2.48300e-14*hvn_mobility*hvn_mobility+-2.02645e-13*hvn_mobility+-1.38260e-12'
+ sky130_fd_pr__nfet_g5v0d10v5__ua_diff_15 = '-9.28797e-13*hvn_mobility*hvn_mobility+-2.37851e-12*hvn_mobility+2.14780e-12'
+ sky130_fd_pr__nfet_g5v0d10v5__ua_diff_16 = '6.42416e-14*hvn_mobility*hvn_mobility+-5.33334e-13*hvn_mobility+2.03550e-12'
+ sky130_fd_pr__nfet_g5v0d10v5__ua_diff_17 = '3.74328e-14*hvn_mobility*hvn_mobility+-4.06869e-13*hvn_mobility+1.20120e-12'
+ sky130_fd_pr__nfet_g5v0d10v5__ua_diff_18 = '3.99844e-14*hvn_mobility*hvn_mobility+-2.42625e-14*hvn_mobility+1.88270e-12'
+ sky130_fd_pr__nfet_g5v0d10v5__ua_diff_19 = '2.86406e-14*hvn_mobility*hvn_mobility+-8.25125e-14*hvn_mobility+1.82940e-12'
+ sky130_fd_pr__nfet_g5v0d10v5__ua_diff_2 = '2.92219e-13*hvn_mobility*hvn_mobility+1.84660e-12*hvn_mobility+-3.38710e-12'
+ sky130_fd_pr__nfet_g5v0d10v5__ua_diff_20 = '1.18606e-13*hvn_mobility*hvn_mobility+-4.52450e-13*hvn_mobility+2.98890e-12'
+ sky130_fd_pr__nfet_g5v0d10v5__ua_diff_21 = '9.45531e-14*hvn_mobility*hvn_mobility+-9.03625e-14*hvn_mobility+3.08820e-12'
+ sky130_fd_pr__nfet_g5v0d10v5__ua_diff_22 = '1.91687e-14*hvn_mobility*hvn_mobility+-4.35225e-13*hvn_mobility+-5.02000e-14'
+ sky130_fd_pr__nfet_g5v0d10v5__ua_diff_23 = '3.52531e-14*hvn_mobility*hvn_mobility+-4.77287e-13*hvn_mobility+2.46660e-12'
+ sky130_fd_pr__nfet_g5v0d10v5__ua_diff_24 = '3.50969e-14*hvn_mobility*hvn_mobility+-2.18213e-13*hvn_mobility+2.78140e-12'
+ sky130_fd_pr__nfet_g5v0d10v5__ua_diff_25 = '2.59125e-14*hvn_mobility*hvn_mobility+-1.69350e-13*hvn_mobility+3.09810e-12'
+ sky130_fd_pr__nfet_g5v0d10v5__ua_diff_26 = '1.20585e-13*hvn_mobility*hvn_mobility+-4.14509e-13*hvn_mobility+7.05500e-13'
+ sky130_fd_pr__nfet_g5v0d10v5__ua_diff_27 = '1.10091e-13*hvn_mobility*hvn_mobility+3.48888e-13*hvn_mobility+2.34770e-12'
+ sky130_fd_pr__nfet_g5v0d10v5__ua_diff_28 = '-1.56675e-11*hvn_mobility*hvn_mobility+-6.28976e-11*hvn_mobility+2.27000e-12'
+ sky130_fd_pr__nfet_g5v0d10v5__ua_diff_29 = '6.44584e-14*hvn_mobility*hvn_mobility+-6.00341e-13*hvn_mobility+1.12070e-12'
+ sky130_fd_pr__nfet_g5v0d10v5__ua_diff_3 = '3.19875e-14*hvn_mobility*hvn_mobility+-2.35550e-13*hvn_mobility+2.07000e-12'
+ sky130_fd_pr__nfet_g5v0d10v5__ua_diff_30 = '5.09687e-14*hvn_mobility*hvn_mobility+-2.64275e-13*hvn_mobility+3.37100e-12'
+ sky130_fd_pr__nfet_g5v0d10v5__ua_diff_31 = '3.39000e-14*hvn_mobility*hvn_mobility+-2.17775e-13*hvn_mobility+2.77840e-12'
+ sky130_fd_pr__nfet_g5v0d10v5__ua_diff_32 = '1.94906e-14*hvn_mobility*hvn_mobility+-1.25338e-13*hvn_mobility+3.67290e-12'
+ sky130_fd_pr__nfet_g5v0d10v5__ua_diff_33 = '1.24336e-13*hvn_mobility*hvn_mobility+-2.44977e-13*hvn_mobility+-4.35080e-13'
+ sky130_fd_pr__nfet_g5v0d10v5__ua_diff_34 = '7.73469e-14*hvn_mobility*hvn_mobility+-1.65313e-13*hvn_mobility+1.58570e-12'
+ sky130_fd_pr__nfet_g5v0d10v5__ua_diff_35 = '2.17375e-13*hvn_mobility*hvn_mobility+7.43250e-13*hvn_mobility+1.16200e-11'
+ sky130_fd_pr__nfet_g5v0d10v5__ua_diff_36 = '6.93656e-14*hvn_mobility*hvn_mobility+4.40787e-13*hvn_mobility+7.14500e-12'
+ sky130_fd_pr__nfet_g5v0d10v5__ua_diff_37 = '1.96231e-13*hvn_mobility*hvn_mobility+1.21515e-12*hvn_mobility+8.89170e-12'
+ sky130_fd_pr__nfet_g5v0d10v5__ua_diff_38 = '1.33637e-13*hvn_mobility*hvn_mobility+9.21250e-14*hvn_mobility+8.96230e-12'
+ sky130_fd_pr__nfet_g5v0d10v5__ua_diff_39 = '1.50981e-13*hvn_mobility*hvn_mobility+7.01775e-13*hvn_mobility+8.52320e-12'
+ sky130_fd_pr__nfet_g5v0d10v5__ua_diff_4 = '1.81091e-14*hvn_mobility*hvn_mobility+-2.52514e-13*hvn_mobility+1.38540e-12'
+ sky130_fd_pr__nfet_g5v0d10v5__ua_diff_40 = '2.65928e-13*hvn_mobility*hvn_mobility+7.27012e-13*hvn_mobility+2.38830e-12'
+ sky130_fd_pr__nfet_g5v0d10v5__ua_diff_41 = '1.72400e-13*hvn_mobility*hvn_mobility+7.87250e-13*hvn_mobility+4.30260e-12'
+ sky130_fd_pr__nfet_g5v0d10v5__ua_diff_42 = '4.38437e-14*hvn_mobility*hvn_mobility+5.26150e-13*hvn_mobility+2.70050e-12'
+ sky130_fd_pr__nfet_g5v0d10v5__ua_diff_43 = '1.16775e-13*hvn_mobility*hvn_mobility+5.43025e-13*hvn_mobility+5.97250e-12'
+ sky130_fd_pr__nfet_g5v0d10v5__ua_diff_44 = '8.54156e-14*hvn_mobility*hvn_mobility+5.29613e-13*hvn_mobility+4.46700e-12'
+ sky130_fd_pr__nfet_g5v0d10v5__ua_diff_45 = '1.32266e-13*hvn_mobility*hvn_mobility+8.06362e-13*hvn_mobility+3.72570e-12'
+ sky130_fd_pr__nfet_g5v0d10v5__ua_diff_46 = '2.73187e-13*hvn_mobility*hvn_mobility+9.12750e-13*hvn_mobility+1.22100e-11'
+ sky130_fd_pr__nfet_g5v0d10v5__ua_diff_47 = '1.35281e-13*hvn_mobility*hvn_mobility+8.26400e-13*hvn_mobility+6.09290e-12'
+ sky130_fd_pr__nfet_g5v0d10v5__ua_diff_48 = '1.70203e-13*hvn_mobility*hvn_mobility+2.52012e-13*hvn_mobility+7.17670e-12'
+ sky130_fd_pr__nfet_g5v0d10v5__ua_diff_5 = '4.57406e-14*hvn_mobility*hvn_mobility+5.48125e-14*hvn_mobility+1.57090e-12'
+ sky130_fd_pr__nfet_g5v0d10v5__ua_diff_6 = '1.60738e-13*hvn_mobility*hvn_mobility+-6.40475e-13*hvn_mobility+4.47580e-12'
+ sky130_fd_pr__nfet_g5v0d10v5__ua_diff_7 = '2.82175e-12*hvn_mobility*hvn_mobility+-1.11879e-11*hvn_mobility+7.17340e-13'
+ sky130_fd_pr__nfet_g5v0d10v5__ua_diff_8 = '6.17937e-14*hvn_mobility*hvn_mobility+2.20800e-13*hvn_mobility+2.70320e-12'
+ sky130_fd_pr__nfet_g5v0d10v5__ua_diff_9 = '1.05069e-13*hvn_mobility*hvn_mobility+6.56850e-13*hvn_mobility+2.39370e-12'
+ sky130_fd_pr__nfet_g5v0d10v5__ub_diff_0 = '1.15921e-20*hvn_mobility*hvn_mobility+2.92174e-19*hvn_mobility+8.94030e-19'
+ sky130_fd_pr__nfet_g5v0d10v5__ub_diff_1 = '2.66594e-21*hvn_mobility*hvn_mobility+1.02431e-19*hvn_mobility+-1.91910e-19'
+ sky130_fd_pr__nfet_g5v0d10v5__ub_diff_10 = '-1.33375e-21*hvn_mobility*hvn_mobility+1.20725e-20*hvn_mobility+1.01180e-19'
+ sky130_fd_pr__nfet_g5v0d10v5__ub_diff_11 = '-4.24687e-22*hvn_mobility*hvn_mobility+7.51863e-20*hvn_mobility+9.19250e-19'
+ sky130_fd_pr__nfet_g5v0d10v5__ub_diff_12 = '3.30031e-21*hvn_mobility*hvn_mobility+1.19769e-19*hvn_mobility+6.42020e-19'
+ sky130_fd_pr__nfet_g5v0d10v5__ub_diff_13 = '-8.26562e-22*hvn_mobility*hvn_mobility+4.18387e-20*hvn_mobility+3.38110e-19'
+ sky130_fd_pr__nfet_g5v0d10v5__ub_diff_14 = '3.89375e-21*hvn_mobility*hvn_mobility+1.23202e-19*hvn_mobility+-1.50940e-19'
+ sky130_fd_pr__nfet_g5v0d10v5__ub_diff_15 = '9.36219e-20*hvn_mobility*hvn_mobility+9.59913e-19*hvn_mobility+1.14650e-18'
+ sky130_fd_pr__nfet_g5v0d10v5__ub_diff_16 = '1.57187e-22*hvn_mobility*hvn_mobility+4.73262e-20*hvn_mobility+-7.10500e-20'
+ sky130_fd_pr__nfet_g5v0d10v5__ub_diff_17 = '1.73750e-22*hvn_mobility*hvn_mobility+4.18288e-20*hvn_mobility+-6.53050e-20'
+ sky130_fd_pr__nfet_g5v0d10v5__ub_diff_18 = '3.70750e-22*hvn_mobility*hvn_mobility+4.58463e-20*hvn_mobility+-4.05370e-20'
+ sky130_fd_pr__nfet_g5v0d10v5__ub_diff_19 = '-1.09256e-21*hvn_mobility*hvn_mobility+1.17475e-20*hvn_mobility+-5.11990e-20'
+ sky130_fd_pr__nfet_g5v0d10v5__ub_diff_2 = '1.87434e-20*hvn_mobility*hvn_mobility+3.64904e-19*hvn_mobility+9.49190e-19'
+ sky130_fd_pr__nfet_g5v0d10v5__ub_diff_20 = '3.39687e-22*hvn_mobility*hvn_mobility+1.01271e-19*hvn_mobility+6.92180e-19'
+ sky130_fd_pr__nfet_g5v0d10v5__ub_diff_21 = '-2.19500e-21*hvn_mobility*hvn_mobility+3.66525e-20*hvn_mobility+5.12690e-19'
+ sky130_fd_pr__nfet_g5v0d10v5__ub_diff_22 = '4.09438e-22*hvn_mobility*hvn_mobility+5.29487e-20*hvn_mobility+-3.41860e-20'
+ sky130_fd_pr__nfet_g5v0d10v5__ub_diff_23 = '-6.85938e-23*hvn_mobility*hvn_mobility+3.60306e-20*hvn_mobility+-1.82730e-19'
+ sky130_fd_pr__nfet_g5v0d10v5__ub_diff_24 = '-1.01250e-22*hvn_mobility*hvn_mobility+3.39950e-20*hvn_mobility+-2.65550e-19'
+ sky130_fd_pr__nfet_g5v0d10v5__ub_diff_25 = '-1.36656e-21*hvn_mobility*hvn_mobility+8.46250e-22*hvn_mobility+-2.83300e-19'
+ sky130_fd_pr__nfet_g5v0d10v5__ub_diff_26 = '1.09656e-21*hvn_mobility*hvn_mobility+1.34234e-19*hvn_mobility+7.96520e-19'
+ sky130_fd_pr__nfet_g5v0d10v5__ub_diff_27 = '-1.21875e-22*hvn_mobility*hvn_mobility+7.91650e-20*hvn_mobility+5.73870e-19'
+ sky130_fd_pr__nfet_g5v0d10v5__ub_diff_28 = '1.99306e-20*hvn_mobility*hvn_mobility+1.55958e-19*hvn_mobility+1.96980e-19'
+ sky130_fd_pr__nfet_g5v0d10v5__ub_diff_29 = '4.12594e-22*hvn_mobility*hvn_mobility+5.66779e-20*hvn_mobility+-2.21290e-19'
+ sky130_fd_pr__nfet_g5v0d10v5__ub_diff_3 = '1.85000e-23*hvn_mobility*hvn_mobility+4.33715e-20*hvn_mobility+-1.10470e-19'
+ sky130_fd_pr__nfet_g5v0d10v5__ub_diff_30 = '9.25094e-22*hvn_mobility*hvn_mobility+6.17654e-20*hvn_mobility+-3.03440e-19'
+ sky130_fd_pr__nfet_g5v0d10v5__ub_diff_31 = '-1.77500e-22*hvn_mobility*hvn_mobility+3.38075e-20*hvn_mobility+-3.16760e-19'
+ sky130_fd_pr__nfet_g5v0d10v5__ub_diff_32 = '-1.48625e-21*hvn_mobility*hvn_mobility+-5.42500e-22*hvn_mobility+-3.64590e-19'
+ sky130_fd_pr__nfet_g5v0d10v5__ub_diff_33 = '1.27219e-21*hvn_mobility*hvn_mobility+1.35094e-19*hvn_mobility+8.36370e-19'
+ sky130_fd_pr__nfet_g5v0d10v5__ub_diff_34 = '8.37187e-22*hvn_mobility*hvn_mobility+7.55412e-20*hvn_mobility+-1.47520e-19'
+ sky130_fd_pr__nfet_g5v0d10v5__ub_diff_35 = '-1.65816e-21*hvn_mobility*hvn_mobility+2.87251e-20*hvn_mobility+1.88970e-19'
+ sky130_fd_pr__nfet_g5v0d10v5__ub_diff_36 = '-3.85312e-22*hvn_mobility*hvn_mobility+3.16292e-20*hvn_mobility+-5.09380e-20'
+ sky130_fd_pr__nfet_g5v0d10v5__ub_diff_37 = '-2.53750e-23*hvn_mobility*hvn_mobility+4.21437e-20*hvn_mobility+5.49410e-20'
+ sky130_fd_pr__nfet_g5v0d10v5__ub_diff_38 = '3.32850e-21*hvn_mobility*hvn_mobility+7.56287e-20*hvn_mobility+8.51490e-20'
+ sky130_fd_pr__nfet_g5v0d10v5__ub_diff_39 = '6.35394e-21*hvn_mobility*hvn_mobility+1.07311e-19*hvn_mobility+-3.77180e-20'
+ sky130_fd_pr__nfet_g5v0d10v5__ub_diff_4 = '3.94312e-22*hvn_mobility*hvn_mobility+4.46687e-20*hvn_mobility+-7.73640e-20'
+ sky130_fd_pr__nfet_g5v0d10v5__ub_diff_40 = '1.34156e-21*hvn_mobility*hvn_mobility+1.35964e-19*hvn_mobility+7.42680e-19'
+ sky130_fd_pr__nfet_g5v0d10v5__ub_diff_41 = '-7.83906e-21*hvn_mobility*hvn_mobility+1.66812e-20*hvn_mobility+5.53700e-19'
+ sky130_fd_pr__nfet_g5v0d10v5__ub_diff_42 = '7.30937e-22*hvn_mobility*hvn_mobility+9.59113e-20*hvn_mobility+5.45190e-19'
+ sky130_fd_pr__nfet_g5v0d10v5__ub_diff_43 = '-9.11625e-22*hvn_mobility*hvn_mobility+3.17315e-20*hvn_mobility+2.33840e-19'
+ sky130_fd_pr__nfet_g5v0d10v5__ub_diff_44 = '-7.16750e-22*hvn_mobility*hvn_mobility+2.76720e-20*hvn_mobility+1.36550e-19'
+ sky130_fd_pr__nfet_g5v0d10v5__ub_diff_45 = '6.31719e-21*hvn_mobility*hvn_mobility+1.20509e-19*hvn_mobility+1.50930e-19'
+ sky130_fd_pr__nfet_g5v0d10v5__ub_diff_46 = '2.44750e-21*hvn_mobility*hvn_mobility+1.01710e-19*hvn_mobility+1.00270e-18'
+ sky130_fd_pr__nfet_g5v0d10v5__ub_diff_47 = '-1.37716e-21*hvn_mobility*hvn_mobility+3.99061e-20*hvn_mobility+2.68330e-19'
+ sky130_fd_pr__nfet_g5v0d10v5__ub_diff_48 = '-1.26906e-21*hvn_mobility*hvn_mobility+4.43863e-20*hvn_mobility+4.29170e-19'
+ sky130_fd_pr__nfet_g5v0d10v5__ub_diff_5 = '4.82125e-22*hvn_mobility*hvn_mobility+4.56475e-20*hvn_mobility+1.43960e-20'
+ sky130_fd_pr__nfet_g5v0d10v5__ub_diff_6 = '-1.05406e-21*hvn_mobility*hvn_mobility+6.11812e-20*hvn_mobility+4.79900e-19'
+ sky130_fd_pr__nfet_g5v0d10v5__ub_diff_7 = '-4.96322e-21*hvn_mobility*hvn_mobility+5.01754e-20*hvn_mobility+2.39360e-19'
+ sky130_fd_pr__nfet_g5v0d10v5__ub_diff_8 = '-4.72594e-22*hvn_mobility*hvn_mobility+3.03729e-20*hvn_mobility+1.69050e-19'
+ sky130_fd_pr__nfet_g5v0d10v5__ub_diff_9 = '5.06562e-21*hvn_mobility*hvn_mobility+1.11312e-19*hvn_mobility+2.06970e-19'
+ sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_0 = '7.23906e+01*hvn_saturation*hvn_saturation+2.13531e+03*hvn_saturation+-3.45400e+03'
+ sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_11 = '9.33375e+01*hvn_saturation*hvn_saturation+3.27227e+03*hvn_saturation+-5.02930e+03'
+ sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_12 = '1.37822e+02*hvn_saturation*hvn_saturation+3.34186e+03*hvn_saturation+-5.70370e+03'
+ sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_13 = '1.09897e+02*hvn_saturation*hvn_saturation+3.12029e+03*hvn_saturation+-4.33620e+03'
+ sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_15 = '5.07919e+02*hvn_saturation*hvn_saturation+4.52825e+03*hvn_saturation+-2.32970e+03'
+ sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_2 = '8.07025e+01*hvn_saturation*hvn_saturation+1.98546e+03*hvn_saturation+-2.40090e+02'
+ sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_20 = '4.99500e+01*hvn_saturation*hvn_saturation+2.50510e+03*hvn_saturation+-2.13080e+03'
+ sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_21 = '3.42281e+01*hvn_saturation*hvn_saturation+2.13439e+03*hvn_saturation+-3.42210e+03'
+ sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_26 = '4.06750e+01*hvn_saturation*hvn_saturation+2.00498e+03*hvn_saturation+-3.12090e+03'
+ sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_27 = '3.75469e+01*hvn_saturation*hvn_saturation+2.03714e+03*hvn_saturation+-2.09690e+03'
+ sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_28 = '5.77487e+01*hvn_saturation*hvn_saturation+2.38294e+03*hvn_saturation+-5.46930e+02'
+ sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_33 = '2.92506e+01*hvn_saturation*hvn_saturation+1.93930e+03*hvn_saturation+-7.93310e+02'
+ sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_34 = '4.66125e+01*hvn_saturation*hvn_saturation+2.14698e+03*hvn_saturation+-3.41590e+03'
+ sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_40 = '1.04503e+02*hvn_saturation*hvn_saturation+3.26001e+03*hvn_saturation+-1.26290e+04'
+ sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_41 = '1.14453e+02*hvn_saturation*hvn_saturation+3.32856e+03*hvn_saturation+-1.04990e+04'
+ sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_42 = '2.81169e+02*hvn_saturation*hvn_saturation+4.14200e+03*hvn_saturation+-5.74570e+03'
+ sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_46 = '2.18413e+02*hvn_saturation*hvn_saturation+3.97650e+03*hvn_saturation+-5.37760e+03'
+ sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_47 = '1.29219e+02*hvn_saturation*hvn_saturation+3.28312e+03*hvn_saturation+-6.45600e+03'
+ sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_48 = '1.21291e+02*hvn_saturation*hvn_saturation+3.19459e+03*hvn_saturation+-9.16230e+03'
+ sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_6 = '8.87562e+01*hvn_saturation*hvn_saturation+3.28380e+03*hvn_saturation+-5.80290e+03'
+ sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_0 = '-1.50750e-04*hvn_threshold*hvn_threshold+2.08127e-02*hvn_threshold+-2.96670e-02'
+ sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_1 = '-1.89375e-05*hvn_threshold*hvn_threshold+2.50225e-03*hvn_threshold+-2.74180e-02'
+ sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_10 = '-2.62500e-06*hvn_threshold*hvn_threshold+2.76000e-04*hvn_threshold+-2.53840e-02'
+ sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_11 = '-1.56594e-04*hvn_threshold*hvn_threshold+2.41181e-02*hvn_threshold+-2.99920e-02'
+ sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_12 = '-7.38750e-05*hvn_threshold*hvn_threshold+1.41725e-02*hvn_threshold+-3.88720e-02'
+ sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_13 = '-3.78125e-05*hvn_threshold*hvn_threshold+7.85525e-03*hvn_threshold+-1.83520e-02'
+ sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_14 = '-1.83438e-05*hvn_threshold*hvn_threshold+2.33788e-03*hvn_threshold+-2.38540e-02'
+ sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_15 = '-8.87500e-05*hvn_threshold*hvn_threshold+2.11133e-02*hvn_threshold+-1.81470e-02'
+ sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_16 = '-2.27500e-05*hvn_threshold*hvn_threshold+3.96525e-03*hvn_threshold+-3.01540e-02'
+ sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_17 = '-4.78125e-06*hvn_threshold*hvn_threshold+1.70113e-03*hvn_threshold+-2.98970e-02'
+ sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_18 = '-6.87500e-07*hvn_threshold*hvn_threshold+-5.68000e-04*hvn_threshold+-2.76180e-02'
+ sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_19 = '-4.81250e-06*hvn_threshold*hvn_threshold+-9.20750e-04*hvn_threshold+-3.05590e-02'
+ sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_2 = '-2.89250e-04*hvn_threshold*hvn_threshold+1.98325e-02*hvn_threshold+-1.90020e-02'
+ sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_20 = '-1.63781e-04*hvn_threshold*hvn_threshold+1.98706e-02*hvn_threshold+-2.72770e-02'
+ sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_21 = '-8.61250e-05*hvn_threshold*hvn_threshold+9.63775e-03*hvn_threshold+-1.86990e-02'
+ sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_22 = '-2.27500e-05*hvn_threshold*hvn_threshold+3.31000e-03*hvn_threshold+-3.34990e-02'
+ sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_23 = '-4.56250e-06*hvn_threshold*hvn_threshold+-2.50000e-06*hvn_threshold+-3.27790e-02'
+ sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_24 = '-1.90625e-06*hvn_threshold*hvn_threshold+-1.28687e-03*hvn_threshold+-3.12050e-02'
+ sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_25 = '-6.06250e-06*hvn_threshold*hvn_threshold+-1.23875e-03*hvn_threshold+-2.57730e-02'
+ sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_26 = '-1.63031e-04*hvn_threshold*hvn_threshold+1.71741e-02*hvn_threshold+-3.75350e-02'
+ sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_27 = '-1.46531e-04*hvn_threshold*hvn_threshold+7.56412e-03*hvn_threshold+-1.58760e-02'
+ sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_28 = '-8.76250e-05*hvn_threshold*hvn_threshold+4.41475e-03*hvn_threshold+-3.15400e-02'
+ sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_29 = '-2.29687e-05*hvn_threshold*hvn_threshold+2.12887e-03*hvn_threshold+-3.80360e-02'
+ sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_3 = '-2.51563e-05*hvn_threshold*hvn_threshold+4.95613e-03*hvn_threshold+-4.75280e-02'
+ sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_30 = '-2.37500e-06*hvn_threshold*hvn_threshold+-2.72750e-04*hvn_threshold+-3.46740e-02'
+ sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_31 = '-1.93750e-06*hvn_threshold*hvn_threshold+-9.35750e-04*hvn_threshold+-3.15400e-02'
+ sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_32 = '-5.87500e-06*hvn_threshold*hvn_threshold+-1.09625e-03*hvn_threshold+-2.82100e-02'
+ sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_33 = '-1.64000e-04*hvn_threshold*hvn_threshold+1.83653e-02*hvn_threshold+-3.54850e-02'
+ sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_34 = '-3.44375e-05*hvn_threshold*hvn_threshold+4.08600e-03*hvn_threshold+-2.96060e-02'
+ sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_35 = '1.82813e-05*hvn_threshold*hvn_threshold+1.79899e-02*hvn_threshold+-5.01230e-02'
+ sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_36 = '5.39063e-05*hvn_threshold*hvn_threshold+6.82012e-03*hvn_threshold+-3.22040e-02'
+ sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_37 = '1.38625e-04*hvn_threshold*hvn_threshold+9.64300e-03*hvn_threshold+-2.96180e-02'
+ sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_38 = '6.26562e-05*hvn_threshold*hvn_threshold+9.86612e-03*hvn_threshold+-2.98930e-02'
+ sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_39 = '6.96656e-05*hvn_threshold*hvn_threshold+7.20666e-03*hvn_threshold+-3.64700e-02'
+ sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_4 = '-3.06250e-06*hvn_threshold*hvn_threshold+1.67850e-03*hvn_threshold+-3.61380e-02'
+ sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_40 = '-1.30250e-04*hvn_threshold*hvn_threshold+3.20513e-02*hvn_threshold+-1.78510e-02'
+ sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_41 = '-7.83125e-05*hvn_threshold*hvn_threshold+2.08590e-02*hvn_threshold+-4.45710e-02'
+ sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_42 = '-1.20313e-05*hvn_threshold*hvn_threshold+1.50459e-02*hvn_threshold+-7.28240e-02'
+ sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_43 = '-2.52344e-05*hvn_threshold*hvn_threshold+8.34556e-03*hvn_threshold+-2.32190e-02'
+ sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_44 = '-5.62500e-07*hvn_threshold*hvn_threshold+4.74075e-03*hvn_threshold+-4.36160e-02'
+ sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_45 = '4.62625e-05*hvn_threshold*hvn_threshold+4.49180e-03*hvn_threshold+-2.06840e-02'
+ sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_46 = '-1.94062e-04*hvn_threshold*hvn_threshold+2.41052e-02*hvn_threshold+-2.86840e-02'
+ sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_47 = '-3.50313e-05*hvn_threshold*hvn_threshold+1.02894e-02*hvn_threshold+-2.24510e-02'
+ sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_48 = '-6.53125e-05*hvn_threshold*hvn_threshold+1.57550e-02*hvn_threshold+-3.20320e-02'
+ sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_5 = '1.43750e-06*hvn_threshold*hvn_threshold+3.55250e-04*hvn_threshold+-2.24640e-02'
+ sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_6 = '-1.61813e-04*hvn_threshold*hvn_threshold+2.47148e-02*hvn_threshold+-4.79020e-02'
+ sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_7 = '2.86406e-04*hvn_threshold*hvn_threshold+4.60262e-03*hvn_threshold+-3.71560e-02'
+ sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_8 = '-1.93750e-06*hvn_threshold*hvn_threshold+2.27350e-03*hvn_threshold+-3.10990e-02'
+ sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_9 = '1.74375e-05*hvn_threshold*hvn_threshold+1.55725e-03*hvn_threshold+-2.37280e-02'
+ sky130_fd_pr__nfet_g5v0d10v5__wint_diff = '8.04375e-09*diff_cd'
+ sky130_fd_pr__esd_nfet_g5v0d10v5__a0_diff_5 = '1.21722e-02*hvn_saturation*hvn_saturation+-1.77450e-02*hvn_saturation+-2.13250e-02'
+ sky130_fd_pr__esd_nfet_g5v0d10v5__a0_diff_8 = '9.23726e-03*hvn_saturation*hvn_saturation+-2.88625e-03*hvn_saturation+7.10880e-03'
+ sky130_fd_pr__esd_nfet_g5v0d10v5__ags_diff_5 = '9.07094e-03*hvn_saturation*hvn_saturation+6.95487e-02*hvn_saturation+-2.66940e-01'
+ sky130_fd_pr__esd_nfet_g5v0d10v5__ags_diff_8 = '-5.86561e-03*hvn_saturation*hvn_saturation+7.71338e-02*hvn_saturation+2.45480e-03'
+ sky130_fd_pr__esd_nfet_g5v0d10v5__ajunction_mult = '9.37500e-07*hvn_diode*hvn_diode+4.43837e-02*hvn_diode+9.95050e-01'
+ sky130_fd_pr__esd_nfet_g5v0d10v5__dlc_diff = '-4.33125e-09*poly_cd'
+ sky130_fd_pr__esd_nfet_g5v0d10v5__dwc_diff = '8.04375e-09*diff_cd'
+ sky130_fd_pr__esd_nfet_g5v0d10v5__k2_diff_0 = '-3.84288e-05*hvn_bodyeffect*hvn_bodyeffect+2.56146e-03*hvn_bodyeffect+1.04060e-02'
+ sky130_fd_pr__esd_nfet_g5v0d10v5__k2_diff_1 = '-3.53550e-05*hvn_bodyeffect*hvn_bodyeffect+2.33942e-03*hvn_bodyeffect+1.03270e-02'
+ sky130_fd_pr__esd_nfet_g5v0d10v5__k2_diff_10 = '-2.24406e-05*hvn_bodyeffect*hvn_bodyeffect+1.49279e-03*hvn_bodyeffect+3.17680e-03'
+ sky130_fd_pr__esd_nfet_g5v0d10v5__k2_diff_2 = '-3.61143e-05*hvn_bodyeffect*hvn_bodyeffect+2.42446e-03*hvn_bodyeffect+1.03040e-02'
+ sky130_fd_pr__esd_nfet_g5v0d10v5__k2_diff_3 = '-3.49250e-05*hvn_bodyeffect*hvn_bodyeffect+2.32870e-03*hvn_bodyeffect+1.00340e-02'
+ sky130_fd_pr__esd_nfet_g5v0d10v5__k2_diff_4 = '-4.50438e-05*hvn_bodyeffect*hvn_bodyeffect+2.98052e-03*hvn_bodyeffect+9.97960e-03'
+ sky130_fd_pr__esd_nfet_g5v0d10v5__k2_diff_5 = '5.10000e-05*hvn_bodyeffect*hvn_bodyeffect+-1.45050e-03*hvn_bodyeffect+4.75330e-02'
+ sky130_fd_pr__esd_nfet_g5v0d10v5__k2_diff_6 = '-3.96813e-05*hvn_bodyeffect*hvn_bodyeffect+2.62222e-03*hvn_bodyeffect+1.00190e-02'
+ sky130_fd_pr__esd_nfet_g5v0d10v5__k2_diff_7 = '-4.12750e-05*hvn_bodyeffect*hvn_bodyeffect+2.74135e-03*hvn_bodyeffect+1.02070e-02'
+ sky130_fd_pr__esd_nfet_g5v0d10v5__k2_diff_8 = '3.76875e-05*hvn_bodyeffect*hvn_bodyeffect+-1.03875e-03*hvn_bodyeffect+1.09770e-02'
+ sky130_fd_pr__esd_nfet_g5v0d10v5__k2_diff_9 = '-2.62281e-05*hvn_bodyeffect*hvn_bodyeffect+1.73514e-03*hvn_bodyeffect+1.44880e-03'
+ sky130_fd_pr__esd_nfet_g5v0d10v5__lint_diff = '-4.33125e-09*poly_cd'
+ sky130_fd_pr__esd_nfet_g5v0d10v5__nfactor_diff_0 = '-1.16563e-04*hvn_subvt*hvn_subvt+2.21188e-02*hvn_subvt+2.33620e-01'
+ sky130_fd_pr__esd_nfet_g5v0d10v5__nfactor_diff_1 = '-7.09375e-05*hvn_subvt*hvn_subvt+1.81337e-02*hvn_subvt+2.30140e-01'
+ sky130_fd_pr__esd_nfet_g5v0d10v5__nfactor_diff_10 = '6.03125e-05*hvn_subvt*hvn_subvt+3.73875e-03*hvn_subvt+2.95910e-01'
+ sky130_fd_pr__esd_nfet_g5v0d10v5__nfactor_diff_2 = '-6.06250e-05*hvn_subvt*hvn_subvt+1.65100e-02*hvn_subvt+2.33910e-01'
+ sky130_fd_pr__esd_nfet_g5v0d10v5__nfactor_diff_3 = '-7.93750e-05*hvn_subvt*hvn_subvt+1.88950e-02*hvn_subvt+2.30860e-01'
+ sky130_fd_pr__esd_nfet_g5v0d10v5__nfactor_diff_4 = '-8.00000e-05*hvn_subvt*hvn_subvt+1.98200e-02*hvn_subvt+2.26090e-01'
+ sky130_fd_pr__esd_nfet_g5v0d10v5__nfactor_diff_5 = '-5.07500e-04*hvn_subvt*hvn_subvt+2.27450e-02*hvn_subvt+2.70560e-01'
+ sky130_fd_pr__esd_nfet_g5v0d10v5__nfactor_diff_6 = '-9.40625e-05*hvn_subvt*hvn_subvt+2.09162e-02*hvn_subvt+2.26690e-01'
+ sky130_fd_pr__esd_nfet_g5v0d10v5__nfactor_diff_7 = '-7.46875e-05*hvn_subvt*hvn_subvt+1.86137e-02*hvn_subvt+1.99320e-01'
+ sky130_fd_pr__esd_nfet_g5v0d10v5__nfactor_diff_8 = '-4.22187e-04*hvn_subvt*hvn_subvt+2.04137e-02*hvn_subvt+2.58880e-01'
+ sky130_fd_pr__esd_nfet_g5v0d10v5__nfactor_diff_9 = '-8.62500e-05*hvn_subvt*hvn_subvt+1.96675e-02*hvn_subvt+2.07210e-01'
+ sky130_fd_pr__esd_nfet_g5v0d10v5__overlap_mult = '2.36250e-04*hvtox*hvtox+3.48425e-02*hvtox+8.98050e-01'
+ sky130_fd_pr__esd_nfet_g5v0d10v5__pjunction_mult = '1.87500e-06*hvn_diode*hvn_diode+5.91425e-02*hvn_diode+1.01440e+00'
+ sky130_fd_pr__esd_nfet_g5v0d10v5__toxe_mult = '1.50000e-02*hvtox+1.00000e+00'
+ sky130_fd_pr__esd_nfet_g5v0d10v5__u0_diff_0 = '-3.20281e-05*hvn_mobility*hvn_mobility+4.75612e-04*hvn_mobility+1.24500e-03'
+ sky130_fd_pr__esd_nfet_g5v0d10v5__u0_diff_1 = '-3.30003e-05*hvn_mobility*hvn_mobility+4.71976e-04*hvn_mobility+2.99590e-03'
+ sky130_fd_pr__esd_nfet_g5v0d10v5__u0_diff_10 = '-2.44813e-05*hvn_mobility*hvn_mobility+5.09462e-04*hvn_mobility+-4.50450e-04'
+ sky130_fd_pr__esd_nfet_g5v0d10v5__u0_diff_2 = '-3.33281e-05*hvn_mobility*hvn_mobility+4.49487e-04*hvn_mobility+1.27410e-03'
+ sky130_fd_pr__esd_nfet_g5v0d10v5__u0_diff_3 = '-3.41688e-05*hvn_mobility*hvn_mobility+4.55250e-04*hvn_mobility+1.06280e-03'
+ sky130_fd_pr__esd_nfet_g5v0d10v5__u0_diff_4 = '-3.19456e-05*hvn_mobility*hvn_mobility+4.61832e-04*hvn_mobility+1.39270e-03'
+ sky130_fd_pr__esd_nfet_g5v0d10v5__u0_diff_5 = '-6.00625e-06*hvn_mobility*hvn_mobility+-1.31425e-04*hvn_mobility+-6.39310e-03'
+ sky130_fd_pr__esd_nfet_g5v0d10v5__u0_diff_6 = '-3.14394e-05*hvn_mobility*hvn_mobility+4.70057e-04*hvn_mobility+1.68740e-03'
+ sky130_fd_pr__esd_nfet_g5v0d10v5__u0_diff_7 = '-3.34088e-05*hvn_mobility*hvn_mobility+4.74360e-04*hvn_mobility+1.44680e-03'
+ sky130_fd_pr__esd_nfet_g5v0d10v5__u0_diff_8 = '1.46875e-06*hvn_mobility*hvn_mobility+-6.11250e-05*hvn_mobility+-8.85190e-03'
+ sky130_fd_pr__esd_nfet_g5v0d10v5__u0_diff_9 = '-3.14781e-05*hvn_mobility*hvn_mobility+4.82187e-04*hvn_mobility+3.79850e-03'
+ sky130_fd_pr__esd_nfet_g5v0d10v5__ua_diff_0 = '5.09074e-13*hvn_mobility*hvn_mobility+3.41621e-13*hvn_mobility+-8.83950e-12'
+ sky130_fd_pr__esd_nfet_g5v0d10v5__ua_diff_1 = '5.25375e-13*hvn_mobility*hvn_mobility+7.09250e-13*hvn_mobility+-2.42000e-11'
+ sky130_fd_pr__esd_nfet_g5v0d10v5__ua_diff_10 = '1.67094e-13*hvn_mobility*hvn_mobility+-3.03525e-13*hvn_mobility+2.88030e-12'
+ sky130_fd_pr__esd_nfet_g5v0d10v5__ua_diff_2 = '3.79175e-13*hvn_mobility*hvn_mobility+-6.39625e-13*hvn_mobility+-7.33300e-12'
+ sky130_fd_pr__esd_nfet_g5v0d10v5__ua_diff_3 = '2.58622e-13*hvn_mobility*hvn_mobility+1.02509e-12*hvn_mobility+-1.72010e-12'
+ sky130_fd_pr__esd_nfet_g5v0d10v5__ua_diff_4 = '4.68688e-13*hvn_mobility*hvn_mobility+1.28125e-12*hvn_mobility+-7.65270e-12'
+ sky130_fd_pr__esd_nfet_g5v0d10v5__ua_diff_5 = '7.42594e-13*hvn_mobility*hvn_mobility+-9.06513e-12*hvn_mobility+8.21280e-11'
+ sky130_fd_pr__esd_nfet_g5v0d10v5__ua_diff_6 = '5.02244e-13*hvn_mobility*hvn_mobility+6.89925e-13*hvn_mobility+-7.01280e-12'
+ sky130_fd_pr__esd_nfet_g5v0d10v5__ua_diff_7 = '2.59384e-13*hvn_mobility*hvn_mobility+1.18726e-12*hvn_mobility+3.22280e-12'
+ sky130_fd_pr__esd_nfet_g5v0d10v5__ua_diff_8 = '2.11791e-12*hvn_mobility*hvn_mobility+-7.77887e-12*hvn_mobility+5.53480e-11'
+ sky130_fd_pr__esd_nfet_g5v0d10v5__ua_diff_9 = '4.99034e-13*hvn_mobility*hvn_mobility+1.88939e-12*hvn_mobility+-1.32830e-11'
+ sky130_fd_pr__esd_nfet_g5v0d10v5__ub_diff_0 = '5.92625e-21*hvn_mobility*hvn_mobility+2.93163e-19*hvn_mobility+2.41530e-19'
+ sky130_fd_pr__esd_nfet_g5v0d10v5__ub_diff_1 = '6.03344e-21*hvn_mobility*hvn_mobility+2.96989e-19*hvn_mobility+3.42210e-19'
+ sky130_fd_pr__esd_nfet_g5v0d10v5__ub_diff_10 = '2.85588e-21*hvn_mobility*hvn_mobility+1.73623e-19*hvn_mobility+8.25060e-20'
+ sky130_fd_pr__esd_nfet_g5v0d10v5__ub_diff_2 = '5.99938e-21*hvn_mobility*hvn_mobility+2.95952e-19*hvn_mobility+3.29100e-19'
+ sky130_fd_pr__esd_nfet_g5v0d10v5__ub_diff_3 = '6.22312e-21*hvn_mobility*hvn_mobility+2.94882e-19*hvn_mobility+3.18300e-19'
+ sky130_fd_pr__esd_nfet_g5v0d10v5__ub_diff_4 = '6.13531e-21*hvn_mobility*hvn_mobility+2.98186e-19*hvn_mobility+2.72490e-19'
+ sky130_fd_pr__esd_nfet_g5v0d10v5__ub_diff_5 = '2.72938e-21*hvn_mobility*hvn_mobility+1.12685e-19*hvn_mobility+-6.17830e-19'
+ sky130_fd_pr__esd_nfet_g5v0d10v5__ub_diff_6 = '6.37688e-21*hvn_mobility*hvn_mobility+3.10353e-19*hvn_mobility+6.06660e-19'
+ sky130_fd_pr__esd_nfet_g5v0d10v5__ub_diff_7 = '6.80125e-21*hvn_mobility*hvn_mobility+3.25178e-19*hvn_mobility+9.79770e-19'
+ sky130_fd_pr__esd_nfet_g5v0d10v5__ub_diff_8 = '1.64469e-21*hvn_mobility*hvn_mobility+1.36976e-19*hvn_mobility+-6.76710e-19'
+ sky130_fd_pr__esd_nfet_g5v0d10v5__ub_diff_9 = '6.73650e-21*hvn_mobility*hvn_mobility+3.33554e-19*hvn_mobility+1.30510e-18'
+ sky130_fd_pr__esd_nfet_g5v0d10v5__vsat_diff_0 = '1.94219e+01*hvn_saturation*hvn_saturation+1.43216e+03*hvn_saturation+-1.67220e+03'
+ sky130_fd_pr__esd_nfet_g5v0d10v5__vsat_diff_1 = '2.03500e+01*hvn_saturation*hvn_saturation+1.45195e+03*hvn_saturation+-1.44370e+03'
+ sky130_fd_pr__esd_nfet_g5v0d10v5__vsat_diff_10 = '-9.90625e-01*hvn_saturation*hvn_saturation+1.27424e+03*hvn_saturation+-2.50220e+03'
+ sky130_fd_pr__esd_nfet_g5v0d10v5__vsat_diff_2 = '1.95063e+01*hvn_saturation*hvn_saturation+1.42331e+03*hvn_saturation+-4.34510e+01'
+ sky130_fd_pr__esd_nfet_g5v0d10v5__vsat_diff_3 = '1.97006e+01*hvn_saturation*hvn_saturation+1.41971e+03*hvn_saturation+3.35400e+01'
+ sky130_fd_pr__esd_nfet_g5v0d10v5__vsat_diff_4 = '1.93387e+01*hvn_saturation*hvn_saturation+1.40379e+03*hvn_saturation+-9.07070e+02'
+ sky130_fd_pr__esd_nfet_g5v0d10v5__vsat_diff_6 = '2.31219e+01*hvn_saturation*hvn_saturation+1.48624e+03*hvn_saturation+1.50000e+03'
+ sky130_fd_pr__esd_nfet_g5v0d10v5__vsat_diff_7 = '2.62500e+01*hvn_saturation*hvn_saturation+1.54505e+03*hvn_saturation+3.01920e+03'
+ sky130_fd_pr__esd_nfet_g5v0d10v5__vsat_diff_9 = '2.46125e+01*hvn_saturation*hvn_saturation+1.48247e+03*hvn_saturation+-1.91500e+02'
+ sky130_fd_pr__esd_nfet_g5v0d10v5__vth0_diff_0 = '1.36250e-06*hvn_threshold*hvn_threshold+4.21430e-03*hvn_threshold+1.27690e-02'
+ sky130_fd_pr__esd_nfet_g5v0d10v5__vth0_diff_1 = '1.61875e-06*hvn_threshold*hvn_threshold+4.16602e-03*hvn_threshold+1.40490e-02'
+ sky130_fd_pr__esd_nfet_g5v0d10v5__vth0_diff_10 = '8.78125e-07*hvn_threshold*hvn_threshold+3.82724e-03*hvn_threshold+1.35430e-02'
+ sky130_fd_pr__esd_nfet_g5v0d10v5__vth0_diff_2 = '4.09375e-07*hvn_threshold*hvn_threshold+4.20411e-03*hvn_threshold+1.33260e-02'
+ sky130_fd_pr__esd_nfet_g5v0d10v5__vth0_diff_3 = '1.50312e-06*hvn_threshold*hvn_threshold+3.72349e-03*hvn_threshold+1.31900e-02'
+ sky130_fd_pr__esd_nfet_g5v0d10v5__vth0_diff_4 = '3.39062e-06*hvn_threshold*hvn_threshold+3.96794e-03*hvn_threshold+1.14690e-02'
+ sky130_fd_pr__esd_nfet_g5v0d10v5__vth0_diff_5 = '-1.91996e-04*hvn_threshold*hvn_threshold+1.84923e-03*hvn_threshold+1.04310e-02'
+ sky130_fd_pr__esd_nfet_g5v0d10v5__vth0_diff_6 = '3.31563e-06*hvn_threshold*hvn_threshold+3.81949e-03*hvn_threshold+1.13960e-02'
+ sky130_fd_pr__esd_nfet_g5v0d10v5__vth0_diff_7 = '2.45625e-06*hvn_threshold*hvn_threshold+3.56092e-03*hvn_threshold+1.18990e-02'
+ sky130_fd_pr__esd_nfet_g5v0d10v5__vth0_diff_8 = '-1.47606e-04*hvn_threshold*hvn_threshold+-4.92320e-04*hvn_threshold+-8.01240e-05'
+ sky130_fd_pr__esd_nfet_g5v0d10v5__vth0_diff_9 = '2.53125e-06*hvn_threshold*hvn_threshold+3.37388e-03*hvn_threshold+2.94300e-03'
+ sky130_fd_pr__esd_nfet_g5v0d10v5__wint_diff = '8.04375e-09*diff_cd'
+ sky130_fd_pr__nfet_05v0_nvt__a0_diff_0 = '-5.41731e-04*hvn_saturation*hvn_saturation+2.16290e-02*hvn_saturation+6.43170e-03'
+ sky130_fd_pr__nfet_05v0_nvt__a0_diff_1 = '-2.70961e-04*hvn_saturation*hvn_saturation+1.17641e-02*hvn_saturation+-4.42130e-04'
+ sky130_fd_pr__nfet_05v0_nvt__a0_diff_3 = '-1.55106e-05*hvn_saturation*hvn_saturation+-7.40925e-05*hvn_saturation+1.27670e-03'
+ sky130_fd_pr__nfet_05v0_nvt__a0_diff_4 = '-4.12300e-03*hvn_saturation*hvn_saturation+5.72388e-02*hvn_saturation+-3.56870e-02'
+ sky130_fd_pr__nfet_05v0_nvt__a0_diff_5 = '-8.62875e-04*hvn_saturation*hvn_saturation+2.57815e-02*hvn_saturation+2.76200e-02'
+ sky130_fd_pr__nfet_05v0_nvt__a0_diff_6 = '-3.47939e-04*hvn_saturation*hvn_saturation+1.69583e-02*hvn_saturation+4.37030e-04'
+ sky130_fd_pr__nfet_05v0_nvt__ags_diff_0 = '-8.85550e-05*hvn_saturation*hvn_saturation+1.97016e-03*hvn_saturation+3.40130e-04'
+ sky130_fd_pr__nfet_05v0_nvt__ags_diff_1 = '-4.87700e-05*hvn_saturation*hvn_saturation+1.55635e-03*hvn_saturation+-5.67080e-04'
+ sky130_fd_pr__nfet_05v0_nvt__ags_diff_3 = '-4.15812e-05*hvn_saturation*hvn_saturation+3.52248e-03*hvn_saturation+7.58940e-03'
+ sky130_fd_pr__nfet_05v0_nvt__ags_diff_4 = '-5.52400e-04*hvn_saturation*hvn_saturation+1.27288e-02*hvn_saturation+-8.46860e-03'
+ sky130_fd_pr__nfet_05v0_nvt__ags_diff_5 = '-5.41688e-05*hvn_saturation*hvn_saturation+5.60975e-03*hvn_saturation+5.32370e-03'
+ sky130_fd_pr__nfet_05v0_nvt__ags_diff_6 = '-3.05062e-06*hvn_saturation*hvn_saturation+3.37325e-03*hvn_saturation+-4.17190e-04'
+ sky130_fd_pr__nfet_05v0_nvt__ajunction_mult = '-1.87500e-06*hvn_diode*hvn_diode+1.02953e-01*hvn_diode+9.76020e-01'
+ sky130_fd_pr__nfet_05v0_nvt__b0_diff_8 = '2.71866e-09*hvn_saturation*hvn_saturation+-3.72864e-08*hvn_saturation+8.00960e-08'
+ sky130_fd_pr__nfet_05v0_nvt__b1_diff_8 = '-8.09664e-10*hvn_saturation*hvn_saturation+2.91469e-09*hvn_saturation+1.65140e-09'
+ sky130_fd_pr__nfet_05v0_nvt__dlc_diff = '9.86313e-10*poly_cd*poly_cd+-7.50000e-09*poly_cd+-1.57810e-08'
+ sky130_fd_pr__nfet_05v0_nvt__dwc_diff = '8.04375e-09*diff_cd'
+ sky130_fd_pr__nfet_05v0_nvt__k2_diff_0 = '-1.11344e-06*hvn_bodyeffect*hvn_bodyeffect+1.10706e-04*hvn_bodyeffect+-2.57080e-04'
+ sky130_fd_pr__nfet_05v0_nvt__k2_diff_1 = '-6.42812e-06*hvn_bodyeffect*hvn_bodyeffect+3.87038e-04*hvn_bodyeffect+-3.97190e-03'
+ sky130_fd_pr__nfet_05v0_nvt__k2_diff_10 = '3.12500e-10*hvn_bodyeffect*hvn_bodyeffect+4.14937e-05*hvn_bodyeffect+6.34570e-04'
+ sky130_fd_pr__nfet_05v0_nvt__k2_diff_2 = '-2.03469e-06*hvn_bodyeffect*hvn_bodyeffect+2.35439e-04*hvn_bodyeffect+1.59150e-03'
+ sky130_fd_pr__nfet_05v0_nvt__k2_diff_3 = '-5.44062e-06*hvn_bodyeffect*hvn_bodyeffect+1.77387e-04*hvn_bodyeffect+-4.63050e-03'
+ sky130_fd_pr__nfet_05v0_nvt__k2_diff_4 = '-7.51563e-06*hvn_bodyeffect*hvn_bodyeffect+1.68387e-04*hvn_bodyeffect+-1.68930e-03'
+ sky130_fd_pr__nfet_05v0_nvt__k2_diff_5 = '-6.28969e-06*hvn_bodyeffect*hvn_bodyeffect+2.50559e-04*hvn_bodyeffect+-1.35530e-04'
+ sky130_fd_pr__nfet_05v0_nvt__k2_diff_6 = '-3.71562e-06*hvn_bodyeffect*hvn_bodyeffect+1.37887e-04*hvn_bodyeffect+-2.36150e-03'
+ sky130_fd_pr__nfet_05v0_nvt__k2_diff_7 = '-2.94747e-06*hvn_bodyeffect*hvn_bodyeffect+9.78224e-05*hvn_bodyeffect+3.52320e-04'
+ sky130_fd_pr__nfet_05v0_nvt__k2_diff_8 = '5.23562e-05*hvn_bodyeffect*hvn_bodyeffect+1.74810e-03*hvn_bodyeffect+-4.92830e-03'
+ sky130_fd_pr__nfet_05v0_nvt__k2_diff_9 = '8.21187e-05*hvn_bodyeffect*hvn_bodyeffect+1.66192e-03*hvn_bodyeffect+-3.00360e-03'
+ sky130_fd_pr__nfet_05v0_nvt__lint_diff = '-4.33125e-09*poly_cd'
+ sky130_fd_pr__nfet_05v0_nvt__nfactor_diff_0 = '2.20063e-04*hvn_subvt*hvn_subvt+-1.76015e-02*hvn_subvt+1.03080e-02'
+ sky130_fd_pr__nfet_05v0_nvt__nfactor_diff_1 = '-1.75844e-04*hvn_subvt*hvn_subvt+1.59659e-02*hvn_subvt+2.99520e-02'
+ sky130_fd_pr__nfet_05v0_nvt__nfactor_diff_10 = '5.13875e-04*hvn_subvt*hvn_subvt+-9.62575e-03*hvn_subvt+1.12750e-02'
+ sky130_fd_pr__nfet_05v0_nvt__nfactor_diff_2 = '5.17250e-04*hvn_subvt*hvn_subvt+-4.04375e-02*hvn_subvt+-4.45860e-02'
+ sky130_fd_pr__nfet_05v0_nvt__nfactor_diff_3 = '9.15938e-05*hvn_subvt*hvn_subvt+1.38279e-02*hvn_subvt+6.40230e-02'
+ sky130_fd_pr__nfet_05v0_nvt__nfactor_diff_4 = '-1.02219e-04*hvn_subvt*hvn_subvt+2.56756e-02*hvn_subvt+2.43930e-02'
+ sky130_fd_pr__nfet_05v0_nvt__nfactor_diff_5 = '5.67187e-05*hvn_subvt*hvn_subvt+1.65679e-02*hvn_subvt+5.30810e-02'
+ sky130_fd_pr__nfet_05v0_nvt__nfactor_diff_6 = '-6.23125e-05*hvn_subvt*hvn_subvt+2.42602e-02*hvn_subvt+5.53460e-02'
+ sky130_fd_pr__nfet_05v0_nvt__nfactor_diff_7 = '4.29544e-04*hvn_subvt*hvn_subvt+-1.77286e-02*hvn_subvt+1.62680e-03'
+ sky130_fd_pr__nfet_05v0_nvt__nfactor_diff_8 = '8.34812e-04*hvn_subvt*hvn_subvt+-5.00750e-03*hvn_subvt+1.74670e-02'
+ sky130_fd_pr__nfet_05v0_nvt__nfactor_diff_9 = '6.29125e-04*hvn_subvt*hvn_subvt+3.88913e-02*hvn_subvt+-1.16110e-02'
+ sky130_fd_pr__nfet_05v0_nvt__overlap_mult = '7.40406e-03*hvtox*hvtox+1.20091e-01*hvtox+7.71170e-01'
+ sky130_fd_pr__nfet_05v0_nvt__pjunction_mult = '-3.12500e-07*hvn_diode*hvn_diode+5.06762e-02*hvn_diode+1.04370e+00'
+ sky130_fd_pr__nfet_05v0_nvt__toxe_mult = '1.30000e-02*hvtox+1.00000e+00'
+ sky130_fd_pr__nfet_05v0_nvt__u0_diff_0 = '-6.23125e-06*hvn_mobility*hvn_mobility+5.75375e-04*hvn_mobility+-7.83780e-03'
+ sky130_fd_pr__nfet_05v0_nvt__u0_diff_1 = '-6.85625e-06*hvn_mobility*hvn_mobility+3.84500e-04*hvn_mobility+-7.04340e-03'
+ sky130_fd_pr__nfet_05v0_nvt__u0_diff_10 = '-3.56750e-05*hvn_mobility*hvn_mobility+5.86400e-04*hvn_mobility+-9.64260e-03'
+ sky130_fd_pr__nfet_05v0_nvt__u0_diff_2 = '-8.51250e-06*hvn_mobility*hvn_mobility+6.62950e-04*hvn_mobility+-8.36300e-03'
+ sky130_fd_pr__nfet_05v0_nvt__u0_diff_3 = '-1.51125e-05*hvn_mobility*hvn_mobility+2.88325e-04*hvn_mobility+-6.63220e-03'
+ sky130_fd_pr__nfet_05v0_nvt__u0_diff_4 = '-1.65906e-05*hvn_mobility*hvn_mobility+4.78687e-04*hvn_mobility+-7.84680e-03'
+ sky130_fd_pr__nfet_05v0_nvt__u0_diff_5 = '-2.18625e-05*hvn_mobility*hvn_mobility+2.38325e-04*hvn_mobility+-7.93990e-03'
+ sky130_fd_pr__nfet_05v0_nvt__u0_diff_6 = '-1.49406e-05*hvn_mobility*hvn_mobility+3.24838e-04*hvn_mobility+-6.81880e-03'
+ sky130_fd_pr__nfet_05v0_nvt__u0_diff_7 = '-2.03375e-05*hvn_mobility*hvn_mobility+6.85975e-04*hvn_mobility+-9.49470e-03'
+ sky130_fd_pr__nfet_05v0_nvt__u0_diff_8 = '-5.37406e-05*hvn_mobility*hvn_mobility+6.54963e-04*hvn_mobility+-8.60230e-03'
+ sky130_fd_pr__nfet_05v0_nvt__u0_diff_9 = '-6.21438e-05*hvn_mobility*hvn_mobility+6.55050e-04*hvn_mobility+-8.92250e-03'
+ sky130_fd_pr__nfet_05v0_nvt__ua_diff_0 = '1.16844e-13*hvn_mobility*hvn_mobility+1.35613e-12*hvn_mobility+-2.69100e-11'
+ sky130_fd_pr__nfet_05v0_nvt__ua_diff_1 = '-5.56250e-14*hvn_mobility*hvn_mobility+8.90000e-14*hvn_mobility+-2.43510e-11'
+ sky130_fd_pr__nfet_05v0_nvt__ua_diff_10 = '1.79031e-13*hvn_mobility*hvn_mobility+1.77012e-12*hvn_mobility+-2.50500e-11'
+ sky130_fd_pr__nfet_05v0_nvt__ua_diff_2 = '1.92125e-13*hvn_mobility*hvn_mobility+2.79325e-12*hvn_mobility+-3.34190e-11'
+ sky130_fd_pr__nfet_05v0_nvt__ua_diff_3 = '6.46563e-14*hvn_mobility*hvn_mobility+8.18375e-13*hvn_mobility+-1.69150e-11'
+ sky130_fd_pr__nfet_05v0_nvt__ua_diff_4 = '-1.41250e-14*hvn_mobility*hvn_mobility+-5.57250e-13*hvn_mobility+-2.42900e-11'
+ sky130_fd_pr__nfet_05v0_nvt__ua_diff_5 = '3.88438e-14*hvn_mobility*hvn_mobility+6.15625e-13*hvn_mobility+-2.15010e-11'
+ sky130_fd_pr__nfet_05v0_nvt__ua_diff_6 = '6.12813e-14*hvn_mobility*hvn_mobility+7.13125e-13*hvn_mobility+-1.90140e-11'
+ sky130_fd_pr__nfet_05v0_nvt__ua_diff_7 = '7.74687e-14*hvn_mobility*hvn_mobility+1.22838e-12*hvn_mobility+-2.89800e-11'
+ sky130_fd_pr__nfet_05v0_nvt__ua_diff_8 = '5.67247e-13*hvn_mobility*hvn_mobility+1.87799e-12*hvn_mobility+-2.28730e-11'
+ sky130_fd_pr__nfet_05v0_nvt__ua_diff_9 = '-3.38751e-12*hvn_mobility*hvn_mobility+1.70485e-11*hvn_mobility+-1.37660e-11'
+ sky130_fd_pr__nfet_05v0_nvt__ub_diff_0 = '1.59063e-21*hvn_mobility*hvn_mobility+7.29625e-20*hvn_mobility+-1.36890e-18'
+ sky130_fd_pr__nfet_05v0_nvt__ub_diff_1 = '7.50000e-22*hvn_mobility*hvn_mobility+3.81000e-20*hvn_mobility+-1.24720e-18'
+ sky130_fd_pr__nfet_05v0_nvt__ub_diff_10 = '3.58562e-21*hvn_mobility*hvn_mobility+1.13743e-19*hvn_mobility+-1.31110e-18'
+ sky130_fd_pr__nfet_05v0_nvt__ub_diff_2 = '3.46875e-21*hvn_mobility*hvn_mobility+1.16075e-19*hvn_mobility+-1.52240e-18'
+ sky130_fd_pr__nfet_05v0_nvt__ub_diff_3 = '1.13875e-21*hvn_mobility*hvn_mobility+4.58275e-20*hvn_mobility+-9.68610e-19'
+ sky130_fd_pr__nfet_05v0_nvt__ub_diff_4 = '1.15312e-21*hvn_mobility*hvn_mobility+5.19375e-20*hvn_mobility+-1.28940e-18'
+ sky130_fd_pr__nfet_05v0_nvt__ub_diff_5 = '5.96875e-22*hvn_mobility*hvn_mobility+4.20875e-20*hvn_mobility+-1.20370e-18'
+ sky130_fd_pr__nfet_05v0_nvt__ub_diff_6 = '1.13469e-21*hvn_mobility*hvn_mobility+4.48887e-20*hvn_mobility+-1.05850e-18'
+ sky130_fd_pr__nfet_05v0_nvt__ub_diff_7 = '2.88438e-21*hvn_mobility*hvn_mobility+9.32375e-20*hvn_mobility+-1.42900e-18'
+ sky130_fd_pr__nfet_05v0_nvt__ub_diff_8 = '3.88313e-21*hvn_mobility*hvn_mobility+1.30557e-19*hvn_mobility+-1.22960e-18'
+ sky130_fd_pr__nfet_05v0_nvt__ub_diff_9 = '1.21937e-20*hvn_mobility*hvn_mobility+1.07000e-19*hvn_mobility+-9.12700e-19'
+ sky130_fd_pr__nfet_05v0_nvt__vsat_diff_10 = '2.42281e+01*hvn_saturation*hvn_saturation+1.75294e+03*hvn_saturation+-4.88990e+03'
+ sky130_fd_pr__nfet_05v0_nvt__vsat_diff_2 = '1.93281e+01*hvn_saturation*hvn_saturation+1.35256e+03*hvn_saturation+-2.84850e+03'
+ sky130_fd_pr__nfet_05v0_nvt__vsat_diff_7 = '1.87781e+01*hvn_saturation*hvn_saturation+1.64861e+03*hvn_saturation+-3.14650e+03'
+ sky130_fd_pr__nfet_05v0_nvt__vsat_diff_9 = '8.31875e+00*hvn_saturation*hvn_saturation+1.87810e+03*hvn_saturation+-6.05270e+03'
+ sky130_fd_pr__nfet_05v0_nvt__vth0_diff_0 = '-7.60625e-06*hvn_threshold*hvn_threshold+9.40775e-03*hvn_threshold+-4.60330e-03'
+ sky130_fd_pr__nfet_05v0_nvt__vth0_diff_1 = '-2.86250e-06*hvn_threshold*hvn_threshold+5.74725e-03*hvn_threshold+-2.20020e-03'
+ sky130_fd_pr__nfet_05v0_nvt__vth0_diff_10 = '-4.40000e-05*hvn_threshold*hvn_threshold+9.14950e-03*hvn_threshold+-1.04950e-02'
+ sky130_fd_pr__nfet_05v0_nvt__vth0_diff_2 = '-9.99375e-06*hvn_threshold*hvn_threshold+1.05278e-02*hvn_threshold+-1.19310e-03'
+ sky130_fd_pr__nfet_05v0_nvt__vth0_diff_3 = '-2.01250e-05*hvn_threshold*hvn_threshold+3.86650e-03*hvn_threshold+-1.34460e-02'
+ sky130_fd_pr__nfet_05v0_nvt__vth0_diff_4 = '-4.31250e-07*hvn_threshold*hvn_threshold+5.17538e-03*hvn_threshold+-5.71660e-03'
+ sky130_fd_pr__nfet_05v0_nvt__vth0_diff_5 = '-2.17500e-05*hvn_threshold*hvn_threshold+4.47813e-03*hvn_threshold+-5.05350e-03'
+ sky130_fd_pr__nfet_05v0_nvt__vth0_diff_6 = '-2.10469e-05*hvn_threshold*hvn_threshold+4.52256e-03*hvn_threshold+-1.10780e-02'
+ sky130_fd_pr__nfet_05v0_nvt__vth0_diff_7 = '-2.03750e-05*hvn_threshold*hvn_threshold+8.82050e-03*hvn_threshold+-1.42540e-02'
+ sky130_fd_pr__nfet_05v0_nvt__vth0_diff_8 = '-9.53719e-05*hvn_threshold*hvn_threshold+8.81576e-03*hvn_threshold+-3.15530e-02'
+ sky130_fd_pr__nfet_05v0_nvt__vth0_diff_9 = '-4.05937e-05*hvn_threshold*hvn_threshold+1.15954e-02*hvn_threshold+-1.03330e-02'
+ sky130_fd_pr__nfet_05v0_nvt__wint_diff = '8.04375e-09*diff_cd'
+ sky130_fd_pr__nfet_01v8_lvt__a0_diff_0 = '-1.02478e-03*lvln_saturation*lvln_saturation+7.70888e-03*lvln_saturation+-7.03880e-02'
+ sky130_fd_pr__nfet_01v8_lvt__a0_diff_1 = '-4.91469e-04*lvln_saturation*lvln_saturation+5.74875e-04*lvln_saturation+-6.49450e-02'
+ sky130_fd_pr__nfet_01v8_lvt__a0_diff_14 = '-3.93875e-04*lvln_saturation*lvln_saturation+-8.82750e-04*lvln_saturation+-6.26760e-02'
+ sky130_fd_pr__nfet_01v8_lvt__a0_diff_15 = '-1.38284e-04*lvln_saturation*lvln_saturation+-2.07531e-03*lvln_saturation+-5.02620e-03'
+ sky130_fd_pr__nfet_01v8_lvt__a0_diff_16 = '3.86375e-05*lvln_saturation*lvln_saturation+8.65625e-04*lvln_saturation+7.77730e-03'
+ sky130_fd_pr__nfet_01v8_lvt__a0_diff_2 = '2.62281e-05*lvln_saturation*lvln_saturation+-1.31721e-03*lvln_saturation+7.11550e-03'
+ sky130_fd_pr__nfet_01v8_lvt__a0_diff_21 = '-3.12337e-04*lvln_saturation*lvln_saturation+-7.56100e-03*lvln_saturation+-6.29860e-03'
+ sky130_fd_pr__nfet_01v8_lvt__a0_diff_22 = '-1.37497e-04*lvln_saturation*lvln_saturation+-4.34501e-03*lvln_saturation+-2.48090e-02'
+ sky130_fd_pr__nfet_01v8_lvt__a0_diff_23 = '2.61344e-05*lvln_saturation*lvln_saturation+7.48413e-04*lvln_saturation+3.44490e-03'
+ sky130_fd_pr__nfet_01v8_lvt__a0_diff_7 = '-5.68281e-04*lvln_saturation*lvln_saturation+-1.29937e-03*lvln_saturation+-5.85100e-02'
+ sky130_fd_pr__nfet_01v8_lvt__a0_diff_8 = '-2.96531e-04*lvln_saturation*lvln_saturation+-4.13812e-03*lvln_saturation+-5.19000e-02'
+ sky130_fd_pr__nfet_01v8_lvt__a0_diff_9 = '3.87094e-05*lvln_saturation*lvln_saturation+-9.32625e-05*lvln_saturation+7.85690e-03'
+ sky130_fd_pr__nfet_01v8_lvt__ags_diff_0 = '-1.67312e-03*lvln_saturation*lvln_saturation+1.22500e-02*lvln_saturation+-1.24230e-01'
+ sky130_fd_pr__nfet_01v8_lvt__ags_diff_1 = '-9.88125e-04*lvln_saturation*lvln_saturation+8.77500e-04*lvln_saturation+-1.41890e-01'
+ sky130_fd_pr__nfet_01v8_lvt__ags_diff_14 = '-5.44625e-04*lvln_saturation*lvln_saturation+-1.48875e-03*lvln_saturation+-9.09510e-02'
+ sky130_fd_pr__nfet_01v8_lvt__ags_diff_15 = '-3.75328e-04*lvln_saturation*lvln_saturation+-6.27344e-03*lvln_saturation+-2.83510e-02'
+ sky130_fd_pr__nfet_01v8_lvt__ags_diff_16 = '-2.32500e-04*lvln_saturation*lvln_saturation+-3.98000e-03*lvln_saturation+-4.80530e-02'
+ sky130_fd_pr__nfet_01v8_lvt__ags_diff_2 = '-3.14438e-04*lvln_saturation*lvln_saturation+1.10003e-02*lvln_saturation+2.20060e-02'
+ sky130_fd_pr__nfet_01v8_lvt__ags_diff_21 = '-3.99500e-04*lvln_saturation*lvln_saturation+-9.25325e-03*lvln_saturation+-1.41080e-02'
+ sky130_fd_pr__nfet_01v8_lvt__ags_diff_22 = '-3.85281e-04*lvln_saturation*lvln_saturation+-1.05526e-02*lvln_saturation+-6.54450e-02'
+ sky130_fd_pr__nfet_01v8_lvt__ags_diff_23 = '-1.99359e-04*lvln_saturation*lvln_saturation+-3.43179e-03*lvln_saturation+9.13260e-03'
+ sky130_fd_pr__nfet_01v8_lvt__ags_diff_7 = '-6.61031e-04*lvln_saturation*lvln_saturation+-1.73888e-03*lvln_saturation+-7.46270e-02'
+ sky130_fd_pr__nfet_01v8_lvt__ags_diff_8 = '-4.48906e-04*lvln_saturation*lvln_saturation+-6.35113e-03*lvln_saturation+-8.01930e-02'
+ sky130_fd_pr__nfet_01v8_lvt__ags_diff_9 = '-2.60744e-04*lvln_saturation*lvln_saturation+1.86352e-03*lvln_saturation+-1.17090e-02'
+ sky130_fd_pr__nfet_01v8_lvt__ajunction_mult = '-2.59375e-05*lvn_diode*lvn_diode+4.38787e-02*lvn_diode+1.00040e+00'
+ sky130_fd_pr__nfet_01v8_lvt__b0_diff_28 = '2.69131e-09*lvln_saturation*lvln_saturation+-1.69675e-08*lvln_saturation+8.06090e-08'
+ sky130_fd_pr__nfet_01v8_lvt__b1_diff_28 = '4.11456e-10*lvln_saturation*lvln_saturation+1.72440e-09*lvln_saturation+2.22210e-09'
+ sky130_fd_pr__nfet_01v8_lvt__dlc_diff = '-4.91625e-11*poly_cd*poly_cd+-3.37112e-09*poly_cd+-1.36190e-09'
+ sky130_fd_pr__nfet_01v8_lvt__dwc_diff = '8.04375e-09*diff_cd'
+ sky130_fd_pr__nfet_01v8_lvt__k2_diff_0 = '1.29219e-05*lvln_bodyeffect*lvln_bodyeffect+4.47375e-05*lvln_bodyeffect+8.15680e-03'
+ sky130_fd_pr__nfet_01v8_lvt__k2_diff_1 = '9.51875e-06*lvln_bodyeffect*lvln_bodyeffect+-1.41525e-04*lvln_bodyeffect+7.33230e-03'
+ sky130_fd_pr__nfet_01v8_lvt__k2_diff_10 = '8.12781e-04*lvln_bodyeffect*lvln_bodyeffect+-9.65787e-03*lvln_bodyeffect+3.07900e-03'
+ sky130_fd_pr__nfet_01v8_lvt__k2_diff_11 = '3.89181e-04*lvln_bodyeffect*lvln_bodyeffect+-6.54650e-03*lvln_bodyeffect+4.21110e-03'
+ sky130_fd_pr__nfet_01v8_lvt__k2_diff_12 = '1.38847e-04*lvln_bodyeffect*lvln_bodyeffect+-1.98154e-03*lvln_bodyeffect+7.72530e-03'
+ sky130_fd_pr__nfet_01v8_lvt__k2_diff_13 = '7.43750e-06*lvln_bodyeffect*lvln_bodyeffect+-3.20750e-04*lvln_bodyeffect+1.11500e-02'
+ sky130_fd_pr__nfet_01v8_lvt__k2_diff_14 = '-3.31250e-07*lvln_bodyeffect*lvln_bodyeffect+1.04000e-04*lvln_bodyeffect+3.23330e-03'
+ sky130_fd_pr__nfet_01v8_lvt__k2_diff_15 = '5.31250e-07*lvln_bodyeffect*lvln_bodyeffect+6.29250e-05*lvln_bodyeffect+-5.88460e-03'
+ sky130_fd_pr__nfet_01v8_lvt__k2_diff_16 = '-2.26562e-06*lvln_bodyeffect*lvln_bodyeffect+3.58562e-04*lvln_bodyeffect+9.61400e-03'
+ sky130_fd_pr__nfet_01v8_lvt__k2_diff_17 = '8.61656e-04*lvln_bodyeffect*lvln_bodyeffect+-1.05986e-02*lvln_bodyeffect+2.83200e-03'
+ sky130_fd_pr__nfet_01v8_lvt__k2_diff_18 = '3.84850e-04*lvln_bodyeffect*lvln_bodyeffect+-6.49788e-03*lvln_bodyeffect+4.96990e-03'
+ sky130_fd_pr__nfet_01v8_lvt__k2_diff_19 = '1.11193e-04*lvln_bodyeffect*lvln_bodyeffect+-1.86765e-03*lvln_bodyeffect+5.43530e-03'
+ sky130_fd_pr__nfet_01v8_lvt__k2_diff_2 = '9.06875e-06*lvln_bodyeffect*lvln_bodyeffect+-7.32500e-05*lvln_bodyeffect+9.75390e-03'
+ sky130_fd_pr__nfet_01v8_lvt__k2_diff_20 = '-4.34375e-07*lvln_bodyeffect*lvln_bodyeffect+3.76487e-04*lvln_bodyeffect+3.04780e-03'
+ sky130_fd_pr__nfet_01v8_lvt__k2_diff_21 = '-7.63750e-06*lvln_bodyeffect*lvln_bodyeffect+3.93125e-04*lvln_bodyeffect+-3.59820e-03'
+ sky130_fd_pr__nfet_01v8_lvt__k2_diff_22 = '-3.68750e-06*lvln_bodyeffect*lvln_bodyeffect+3.08425e-04*lvln_bodyeffect+8.57370e-03'
+ sky130_fd_pr__nfet_01v8_lvt__k2_diff_23 = '-2.90625e-07*lvln_bodyeffect*lvln_bodyeffect+2.78188e-04*lvln_bodyeffect+7.57100e-03'
+ sky130_fd_pr__nfet_01v8_lvt__k2_diff_24 = '7.68256e-04*lvln_bodyeffect*lvln_bodyeffect+-9.34400e-03*lvln_bodyeffect+8.56890e-03'
+ sky130_fd_pr__nfet_01v8_lvt__k2_diff_25 = '3.60403e-04*lvln_bodyeffect*lvln_bodyeffect+-5.08014e-03*lvln_bodyeffect+6.58600e-03'
+ sky130_fd_pr__nfet_01v8_lvt__k2_diff_26 = '1.06734e-04*lvln_bodyeffect*lvln_bodyeffect+-1.78299e-03*lvln_bodyeffect+6.75130e-03'
+ sky130_fd_pr__nfet_01v8_lvt__k2_diff_27 = '2.84688e-06*lvln_bodyeffect*lvln_bodyeffect+6.56375e-05*lvln_bodyeffect+3.92910e-03'
+ sky130_fd_pr__nfet_01v8_lvt__k2_diff_28 = '1.32722e-04*lvln_bodyeffect*lvln_bodyeffect+-4.41488e-04*lvln_bodyeffect+2.71000e-03'
+ sky130_fd_pr__nfet_01v8_lvt__k2_diff_29 = '8.47700e-04*lvln_bodyeffect*lvln_bodyeffect+-8.66187e-03*lvln_bodyeffect+1.00930e-03'
+ sky130_fd_pr__nfet_01v8_lvt__k2_diff_3 = '8.27400e-04*lvln_bodyeffect*lvln_bodyeffect+-8.65362e-03*lvln_bodyeffect+2.54710e-03'
+ sky130_fd_pr__nfet_01v8_lvt__k2_diff_30 = '4.03418e-04*lvln_bodyeffect*lvln_bodyeffect+-3.90980e-03*lvln_bodyeffect+-8.08890e-04'
+ sky130_fd_pr__nfet_01v8_lvt__k2_diff_31 = '7.72275e-04*lvln_bodyeffect*lvln_bodyeffect+-5.87550e-03*lvln_bodyeffect+-3.12040e-03'
+ sky130_fd_pr__nfet_01v8_lvt__k2_diff_32 = '7.72819e-04*lvln_bodyeffect*lvln_bodyeffect+-6.20550e-03*lvln_bodyeffect+-4.04610e-03'
+ sky130_fd_pr__nfet_01v8_lvt__k2_diff_33 = '7.81106e-04*lvln_bodyeffect*lvln_bodyeffect+-6.15838e-03*lvln_bodyeffect+-4.96220e-03'
+ sky130_fd_pr__nfet_01v8_lvt__k2_diff_34 = '7.52500e-04*lvln_bodyeffect*lvln_bodyeffect+-8.31525e-03*lvln_bodyeffect+4.71900e-03'
+ sky130_fd_pr__nfet_01v8_lvt__k2_diff_35 = '7.82919e-04*lvln_bodyeffect*lvln_bodyeffect+-9.51225e-03*lvln_bodyeffect+2.23630e-03'
+ sky130_fd_pr__nfet_01v8_lvt__k2_diff_36 = '8.64638e-04*lvln_bodyeffect*lvln_bodyeffect+-1.05616e-02*lvln_bodyeffect+3.15830e-03'
+ sky130_fd_pr__nfet_01v8_lvt__k2_diff_37 = '1.03573e-04*lvln_bodyeffect*lvln_bodyeffect+-1.86916e-03*lvln_bodyeffect+5.17620e-03'
+ sky130_fd_pr__nfet_01v8_lvt__k2_diff_4 = '3.85494e-04*lvln_bodyeffect*lvln_bodyeffect+-5.62800e-03*lvln_bodyeffect+1.98710e-03'
+ sky130_fd_pr__nfet_01v8_lvt__k2_diff_5 = '2.52759e-04*lvln_bodyeffect*lvln_bodyeffect+-6.58137e-04*lvln_bodyeffect+5.45730e-03'
+ sky130_fd_pr__nfet_01v8_lvt__k2_diff_6 = '2.42156e-05*lvln_bodyeffect*lvln_bodyeffect+6.79638e-04*lvln_bodyeffect+1.20100e-03'
+ sky130_fd_pr__nfet_01v8_lvt__k2_diff_7 = '-2.92500e-06*lvln_bodyeffect*lvln_bodyeffect+3.72600e-04*lvln_bodyeffect+4.86510e-03'
+ sky130_fd_pr__nfet_01v8_lvt__k2_diff_8 = '-3.30375e-06*lvln_bodyeffect*lvln_bodyeffect+5.57840e-04*lvln_bodyeffect+2.93230e-03'
+ sky130_fd_pr__nfet_01v8_lvt__k2_diff_9 = '-2.43750e-07*lvln_bodyeffect*lvln_bodyeffect+2.00325e-04*lvln_bodyeffect+6.42030e-03'
+ sky130_fd_pr__nfet_01v8_lvt__lint_diff = '-4.33125e-09*poly_cd'
+ sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_0 = '-1.33094e-03*lvn_subvt*lvn_subvt+4.33588e-02*lvn_subvt+8.91660e-01'
+ sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_1 = '-2.87500e-05*lvn_subvt*lvn_subvt+-8.84750e-03*lvn_subvt+4.31950e-01'
+ sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_10 = '7.80000e-03*lvn_subvt*lvn_subvt+8.37500e-03*lvn_subvt+1.36320e+00'
+ sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_11 = '-2.00000e-04*lvn_subvt*lvn_subvt+5.19250e-02*lvn_subvt+1.37830e+00'
+ sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_12 = '-2.88438e-03*lvn_subvt*lvn_subvt+1.39375e-02*lvn_subvt+1.06580e+00'
+ sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_13 = '2.37500e-04*lvn_subvt*lvn_subvt+-5.00000e-05*lvn_subvt+1.24980e+00'
+ sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_14 = '-3.86562e-04*lvn_subvt*lvn_subvt+1.41712e-02*lvn_subvt+6.91020e-01'
+ sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_15 = '-6.21562e-04*lvn_subvt*lvn_subvt+3.38113e-02*lvn_subvt+6.31960e-01'
+ sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_16 = '-5.67812e-04*lvn_subvt*lvn_subvt+1.00862e-02*lvn_subvt+1.51080e-01'
+ sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_17 = '1.06250e-04*lvn_subvt*lvn_subvt+2.38500e-02*lvn_subvt+1.44370e+00'
+ sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_18 = '3.50000e-04*lvn_subvt*lvn_subvt+7.80000e-03*lvn_subvt+1.32020e+00'
+ sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_19 = '2.91250e-04*lvn_subvt*lvn_subvt+7.12350e-02*lvn_subvt+1.01290e+00'
+ sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_2 = '1.64375e-04*lvn_subvt*lvn_subvt+3.35750e-02*lvn_subvt+8.71670e-01'
+ sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_20 = '2.10000e-04*lvn_subvt*lvn_subvt+-4.46100e-02*lvn_subvt+1.04000e+00'
+ sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_21 = '6.65625e-05*lvn_subvt*lvn_subvt+-2.53125e-03*lvn_subvt+7.56520e-01'
+ sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_22 = '-2.19687e-04*lvn_subvt*lvn_subvt+9.51625e-03*lvn_subvt+4.99700e-01'
+ sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_23 = '-8.57812e-04*lvn_subvt*lvn_subvt+1.63212e-02*lvn_subvt+3.92360e-01'
+ sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_24 = '1.65625e-04*lvn_subvt*lvn_subvt+3.06375e-02*lvn_subvt+1.45750e+00'
+ sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_25 = '3.34375e-04*lvn_subvt*lvn_subvt+1.26875e-02*lvn_subvt+1.30490e+00'
+ sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_26 = '7.73750e-04*lvn_subvt*lvn_subvt+8.33550e-02*lvn_subvt+1.01830e+00'
+ sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_27 = '-2.99375e-04*lvn_subvt*lvn_subvt+2.64975e-02*lvn_subvt+1.08420e+00'
+ sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_28 = '-1.32592e-02*lvn_subvt*lvn_subvt+9.60744e-02*lvn_subvt+6.11740e-01'
+ sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_29 = '6.03125e-04*lvn_subvt*lvn_subvt+-5.33750e-03*lvn_subvt+1.64280e+00'
+ sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_3 = '9.71875e-04*lvn_subvt*lvn_subvt+2.34875e-02*lvn_subvt+1.58130e+00'
+ sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_30 = '1.06250e-04*lvn_subvt*lvn_subvt+-2.92000e-02*lvn_subvt+1.51060e+00'
+ sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_31 = '3.66250e-03*lvn_subvt*lvn_subvt+-6.83250e-02*lvn_subvt+1.98940e+00'
+ sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_32 = '-4.06250e-04*lvn_subvt*lvn_subvt+-2.35750e-02*lvn_subvt+2.15590e+00'
+ sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_33 = '1.29063e-03*lvn_subvt*lvn_subvt+4.61250e-03*lvn_subvt+1.96860e+00'
+ sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_34 = '1.41875e-03*lvn_subvt*lvn_subvt+-8.09000e-02*lvn_subvt+1.45480e+00'
+ sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_35 = '4.03125e-04*lvn_subvt*lvn_subvt+3.80875e-02*lvn_subvt+1.41390e+00'
+ sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_36 = '1.56250e-04*lvn_subvt*lvn_subvt+3.24500e-02*lvn_subvt+1.56910e+00'
+ sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_37 = '9.44062e-04*lvn_subvt*lvn_subvt+7.01987e-02*lvn_subvt+1.13410e+00'
+ sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_4 = '4.90625e-04*lvn_subvt*lvn_subvt+2.17625e-02*lvn_subvt+1.61480e+00'
+ sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_5 = '-2.30487e-02*lvn_subvt*lvn_subvt+-1.74875e-02*lvn_subvt+1.24440e+00'
+ sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_6 = '-4.55625e-03*lvn_subvt*lvn_subvt+-6.65500e-02*lvn_subvt+1.24350e+00'
+ sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_7 = '-5.62187e-04*lvn_subvt*lvn_subvt+1.75462e-02*lvn_subvt+8.58750e-01'
+ sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_8 = '-4.74687e-04*lvn_subvt*lvn_subvt+4.50625e-03*lvn_subvt+4.02580e-01'
+ sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_9 = '-5.33750e-04*lvn_subvt*lvn_subvt+2.14575e-02*lvn_subvt+5.10990e-01'
+ sky130_fd_pr__nfet_01v8_lvt__overlap_mult = '-2.39062e-04*lvtox*lvtox+1.49487e-02*lvtox+9.24290e-01'
+ sky130_fd_pr__nfet_01v8_lvt__pjunction_mult = '4.43125e-04*lvn_diode*lvn_diode+3.72125e-02*lvn_diode+8.91760e-01'
+ sky130_fd_pr__rf_nfet_01v8_lvt__aw_cap_mult = '3.75000e-02*nfet_01v8_lvt+1.00000e+00'
+ sky130_fd_pr__rf_nfet_01v8_lvt__aw_cap_mult_p42 = '3.75000e-02*nfet_01v8_lvt+1.00000e+00'
+ sky130_fd_pr__rf_nfet_01v8_lvt__aw_rgate_dist_mult = '3.12500e-03*nfet_01v8_lvt*nfet_01v8_lvt+7.50000e-02*nfet_01v8_lvt+1.00000e+00'
+ sky130_fd_pr__rf_nfet_01v8_lvt__aw_rgate_dist_mult_p42 = '8.75000e-02*nfet_01v8_lvt+1.00000e+00'
+ sky130_fd_pr__rf_nfet_01v8_lvt__aw_rgate_stub_mult = '3.12500e-03*lvln_mobility*lvln_mobility+7.50000e-02*lvln_mobility+1.00000e+00'
+ sky130_fd_pr__rf_nfet_01v8_lvt__aw_rgate_stub_mult_p42 = '8.75000e-02*lvln_mobility+1.00000e+00'
+ sky130_fd_pr__rf_nfet_01v8_lvt_b__ajunction_mult = '-2.59375e-05*lvn_diode*lvn_diode+4.38787e-02*lvn_diode+1.00040e+00'
+ sky130_fd_pr__rf_nfet_01v8_lvt_b__dlc_diff = '-4.91625e-11*poly_cd*poly_cd+-3.37112e-09*poly_cd+-1.36190e-09'
+ sky130_fd_pr__rf_nfet_01v8_lvt_b__lint_diff = '-4.33125e-09*poly_cd'
+ sky130_fd_pr__rf_nfet_01v8_lvt_b__overlap_mult = '-2.39062e-04*lvtox*lvtox+1.49487e-02*lvtox+9.24290e-01'
+ sky130_fd_pr__rf_nfet_01v8_lvt_b__pjunction_mult = '4.43125e-04*lvn_diode*lvn_diode+3.72125e-02*lvn_diode+8.91760e-01'
+ sky130_fd_pr__rf_nfet_01v8_lvt_b__rbpb_mult = '5.00000e-02*lvln_bodyeffect+1.00000e+00'
+ sky130_fd_pr__rf_nfet_01v8_lvt_b__rshg_diff = '1.75000e+00*ic_res'
+ sky130_fd_pr__rf_nfet_01v8_lvt_b__toxe_mult = '1.30000e-02*lvtox+1.00000e+00'
+ sky130_fd_pr__rf_nfet_01v8_lvt_b__wint_diff = '8.04375e-09*diff_cd'
+ sky130_fd_pr__rf_nfet_01v8_lvt_b__xgw_diff = '1.60625e-08*diff_cd'
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__k2_diff_0 = '2.16537e-04*lvln_bodyeffect*lvln_bodyeffect+-2.62240e-03*lvln_bodyeffect+-1.78380e-02'
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__k2_diff_1 = '1.35078e-04*lvln_bodyeffect*lvln_bodyeffect+-2.77109e-03*lvln_bodyeffect+-8.88490e-03'
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__k2_diff_2 = '2.44556e-05*lvln_bodyeffect*lvln_bodyeffect+4.77047e-04*lvln_bodyeffect+-1.89470e-03'
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__k2_diff_3 = '3.99562e-04*lvln_bodyeffect*lvln_bodyeffect+-5.82675e-03*lvln_bodyeffect+-1.30740e-02'
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__k2_diff_4 = '1.72656e-04*lvln_bodyeffect*lvln_bodyeffect+-4.12787e-03*lvln_bodyeffect+-8.65900e-03'
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__k2_diff_5 = '5.23656e-05*lvln_bodyeffect*lvln_bodyeffect+-1.42609e-03*lvln_bodyeffect+-1.49170e-03'
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__k2_diff_6 = '2.87944e-04*lvln_bodyeffect*lvln_bodyeffect+-4.77777e-03*lvln_bodyeffect+-2.04570e-02'
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__k2_diff_7 = '1.70841e-04*lvln_bodyeffect*lvln_bodyeffect+-3.84876e-03*lvln_bodyeffect+-9.14240e-03'
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__k2_diff_8 = '4.93312e-05*lvln_bodyeffect*lvln_bodyeffect+-1.29807e-03*lvln_bodyeffect+-1.35180e-03'
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__u0_diff_0 = '-1.27475e-05*lvln_mobility*lvln_mobility+-3.77012e-04*lvln_mobility+-2.59890e-04'
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__u0_diff_1 = '-3.12666e-05*lvln_mobility*lvln_mobility+-1.65496e-04*lvln_mobility+6.88700e-04'
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__u0_diff_2 = '-3.05450e-05*lvln_mobility*lvln_mobility+-3.54088e-04*lvln_mobility+7.01070e-04'
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__u0_diff_3 = '-2.20438e-05*lvln_mobility*lvln_mobility+-1.72850e-04*lvln_mobility+-4.13870e-03'
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__u0_diff_4 = '-2.53094e-05*lvln_mobility*lvln_mobility+2.66612e-04*lvln_mobility+-2.15790e-03'
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__u0_diff_5 = '-2.68078e-05*lvln_mobility*lvln_mobility+-3.03044e-04*lvln_mobility+-1.04250e-03'
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__u0_diff_6 = '-2.88062e-05*lvln_mobility*lvln_mobility+1.33150e-04*lvln_mobility+-8.36300e-03'
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__u0_diff_7 = '-2.50531e-05*lvln_mobility*lvln_mobility+1.44313e-04*lvln_mobility+-4.23970e-03'
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__u0_diff_8 = '-2.64838e-05*lvln_mobility*lvln_mobility+-4.36215e-04*lvln_mobility+-1.91930e-03'
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__vsat_diff_0 = '7.32625e+01*lvln_saturation*lvln_saturation+7.38425e+03*lvln_saturation+-4.14020e+03'
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__vsat_diff_1 = '2.23044e+02*lvln_saturation*lvln_saturation+7.08838e+03*lvln_saturation+-1.70920e+03'
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__vsat_diff_2 = '1.66750e+02*lvln_saturation*lvln_saturation+4.82325e+03*lvln_saturation+-3.89100e+03'
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__vsat_diff_3 = '1.01919e+02*lvln_saturation*lvln_saturation+8.30375e+03*lvln_saturation+-6.08870e+03'
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__vsat_diff_4 = '7.99125e+01*lvln_saturation*lvln_saturation+6.43850e+03*lvln_saturation+-1.51960e+03'
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__vsat_diff_5 = '2.15024e+02*lvln_saturation*lvln_saturation+5.42662e+03*lvln_saturation+-4.15880e+02'
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__vsat_diff_6 = '-5.46875e+00*lvln_saturation*lvln_saturation+6.40075e+03*lvln_saturation+-5.55550e+03'
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__vsat_diff_7 = '8.60469e+01*lvln_saturation*lvln_saturation+5.73812e+03*lvln_saturation+-7.90250e+02'
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__vsat_diff_8 = '3.04746e+02*lvln_saturation*lvln_saturation+5.30988e+03*lvln_saturation+-1.05440e+02'
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__vth0_diff_0 = '-2.61075e-04*lvln_threshold*lvln_threshold+1.48638e-02*lvln_threshold+-1.90980e-03'
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__vth0_diff_1 = '-1.89812e-04*lvln_threshold*lvln_threshold+1.33500e-02*lvln_threshold+-2.59700e-03'
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__vth0_diff_2 = '-8.61250e-05*lvln_threshold*lvln_threshold+7.26675e-03*lvln_threshold+-1.23440e-02'
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__vth0_diff_3 = '-4.21469e-04*lvln_threshold*lvln_threshold+1.39709e-02*lvln_threshold+-1.12620e-02'
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__vth0_diff_4 = '-2.22750e-04*lvln_threshold*lvln_threshold+1.09125e-02*lvln_threshold+-2.00030e-02'
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__vth0_diff_5 = '-9.39187e-05*lvln_threshold*lvln_threshold+5.23312e-03*lvln_threshold+-7.42980e-03'
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__vth0_diff_6 = '-3.57906e-04*lvln_threshold*lvln_threshold+1.21069e-02*lvln_threshold+-1.02570e-02'
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__vth0_diff_7 = '-2.25563e-04*lvln_threshold*lvln_threshold+9.05225e-03*lvln_threshold+-1.70600e-02'
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__vth0_diff_8 = '-9.28219e-05*lvln_threshold*lvln_threshold+4.10981e-03*lvln_threshold+-6.94560e-03'
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__k2_diff_0 = '2.12059e-04*lvln_bodyeffect*lvln_bodyeffect+-2.43399e-03*lvln_bodyeffect+-1.75260e-02'
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__k2_diff_1 = '1.29553e-04*lvln_bodyeffect*lvln_bodyeffect+-2.65451e-03*lvln_bodyeffect+-9.39780e-03'
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__k2_diff_2 = '4.61625e-05*lvln_bodyeffect*lvln_bodyeffect+-1.24362e-03*lvln_bodyeffect+-2.33740e-03'
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__k2_diff_3 = '3.91781e-04*lvln_bodyeffect*lvln_bodyeffect+-5.71988e-03*lvln_bodyeffect+-1.42820e-02'
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__k2_diff_4 = '1.47672e-04*lvln_bodyeffect*lvln_bodyeffect+-3.83104e-03*lvln_bodyeffect+-9.64160e-03'
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__k2_diff_5 = '4.74750e-05*lvln_bodyeffect*lvln_bodyeffect+-1.34908e-03*lvln_bodyeffect+-2.71180e-03'
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__k2_diff_6 = '3.32397e-04*lvln_bodyeffect*lvln_bodyeffect+-5.34884e-03*lvln_bodyeffect+-1.91600e-02'
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__k2_diff_7 = '1.37456e-04*lvln_bodyeffect*lvln_bodyeffect+-3.47033e-03*lvln_bodyeffect+-1.14380e-02'
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__k2_diff_8 = '4.66500e-05*lvln_bodyeffect*lvln_bodyeffect+-1.20602e-03*lvln_bodyeffect+-2.83740e-03'
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__u0_diff_0 = '-1.76219e-05*lvln_mobility*lvln_mobility+-2.84613e-04*lvln_mobility+-6.03480e-03'
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__u0_diff_1 = '-3.21063e-05*lvln_mobility*lvln_mobility+-6.38750e-05*lvln_mobility+-2.81360e-03'
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__u0_diff_2 = '-2.79550e-05*lvln_mobility*lvln_mobility+-3.72130e-04*lvln_mobility+-1.72530e-03'
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__u0_diff_3 = '-2.89937e-05*lvln_mobility*lvln_mobility+-9.04500e-05*lvln_mobility+-4.67570e-03'
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__u0_diff_4 = '-2.23969e-05*lvln_mobility*lvln_mobility+2.08213e-04*lvln_mobility+-6.94280e-03'
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__u0_diff_5 = '-2.35313e-05*lvln_mobility*lvln_mobility+-2.96250e-04*lvln_mobility+-4.24740e-03'
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__u0_diff_6 = '-3.00687e-05*lvln_mobility*lvln_mobility+1.03425e-04*lvln_mobility+-6.15790e-03'
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__u0_diff_7 = '-2.47250e-05*lvln_mobility*lvln_mobility+5.17000e-05*lvln_mobility+-8.45140e-03'
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__u0_diff_8 = '-2.26906e-05*lvln_mobility*lvln_mobility+-4.28638e-04*lvln_mobility+-6.56350e-03'
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__vsat_diff_0 = '1.74569e+02*lvln_saturation*lvln_saturation+7.96162e+03*lvln_saturation+1.45400e+02'
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__vsat_diff_1 = '2.40744e+02*lvln_saturation*lvln_saturation+7.13262e+03*lvln_saturation+-1.62240e+03'
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__vsat_diff_2 = '1.56794e+02*lvln_saturation*lvln_saturation+5.01475e+03*lvln_saturation+2.32830e+03'
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__vsat_diff_3 = '1.09244e+02*lvln_saturation*lvln_saturation+8.25900e+03*lvln_saturation+-6.71990e+03'
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__vsat_diff_4 = '1.60491e+02*lvln_saturation*lvln_saturation+6.83362e+03*lvln_saturation+3.27640e+02'
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__vsat_diff_5 = '3.10119e+02*lvln_saturation*lvln_saturation+5.98098e+03*lvln_saturation+9.08320e+03'
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__vsat_diff_6 = '6.03562e+01*lvln_saturation*lvln_saturation+7.56138e+03*lvln_saturation+-6.43120e+03'
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__vsat_diff_7 = '1.54125e+02*lvln_saturation*lvln_saturation+6.14912e+03*lvln_saturation+-2.62550e+03'
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__vsat_diff_8 = '5.30047e+02*lvln_saturation*lvln_saturation+7.52931e+03*lvln_saturation+1.41900e+04'
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__vth0_diff_0 = '-2.69669e-04*lvln_threshold*lvln_threshold+1.48915e-02*lvln_threshold+-5.11330e-03'
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__vth0_diff_1 = '-1.94688e-04*lvln_threshold*lvln_threshold+1.34505e-02*lvln_threshold+-1.00420e-02'
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__vth0_diff_2 = '-8.10625e-05*lvln_threshold*lvln_threshold+7.25900e-03*lvln_threshold+-1.77560e-02'
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__vth0_diff_3 = '-4.34213e-04*lvln_threshold*lvln_threshold+1.42046e-02*lvln_threshold+-8.51510e-03'
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__vth0_diff_4 = '-1.97313e-04*lvln_threshold*lvln_threshold+1.04557e-02*lvln_threshold+-1.70880e-02'
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__vth0_diff_5 = '-8.34781e-05*lvln_threshold*lvln_threshold+4.97284e-03*lvln_threshold+-1.99910e-02'
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__vth0_diff_6 = '-3.76781e-04*lvln_threshold*lvln_threshold+1.26681e-02*lvln_threshold+-1.30210e-02'
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__vth0_diff_7 = '-1.85438e-04*lvln_threshold*lvln_threshold+8.48675e-03*lvln_threshold+-1.86740e-02'
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__vth0_diff_8 = '-8.59000e-05*lvln_threshold*lvln_threshold+3.90465e-03*lvln_threshold+-2.40190e-02'
+ sky130_fd_pr__nfet_01v8_lvt__toxe_mult = '1.30000e-02*lvtox+1.00000e+00'
+ sky130_fd_pr__nfet_01v8_lvt__u0_diff_0 = '-3.86092e-05*lvln_mobility*lvln_mobility+-4.16513e-04*lvln_mobility+7.37980e-05'
+ sky130_fd_pr__nfet_01v8_lvt__u0_diff_1 = '-3.57631e-05*lvln_mobility*lvln_mobility+-3.84433e-04*lvln_mobility+-9.77360e-04'
+ sky130_fd_pr__nfet_01v8_lvt__u0_diff_10 = '-2.15503e-05*lvln_mobility*lvln_mobility+4.08574e-04*lvln_mobility+-1.91150e-03'
+ sky130_fd_pr__nfet_01v8_lvt__u0_diff_11 = '-2.95187e-05*lvln_mobility*lvln_mobility+3.32838e-04*lvln_mobility+3.56250e-04'
+ sky130_fd_pr__nfet_01v8_lvt__u0_diff_12 = '-1.37567e-04*lvln_mobility*lvln_mobility+-6.57826e-04*lvln_mobility+-2.18920e-04'
+ sky130_fd_pr__nfet_01v8_lvt__u0_diff_13 = '-1.86809e-05*lvln_mobility*lvln_mobility+2.57876e-04*lvln_mobility+4.82990e-04'
+ sky130_fd_pr__nfet_01v8_lvt__u0_diff_14 = '-1.40191e-05*lvln_mobility*lvln_mobility+1.27701e-04*lvln_mobility+9.56300e-04'
+ sky130_fd_pr__nfet_01v8_lvt__u0_diff_15 = '-1.27256e-05*lvln_mobility*lvln_mobility+5.49375e-05*lvln_mobility+6.92510e-04'
+ sky130_fd_pr__nfet_01v8_lvt__u0_diff_16 = '-1.13497e-05*lvln_mobility*lvln_mobility+7.42537e-05*lvln_mobility+3.78290e-04'
+ sky130_fd_pr__nfet_01v8_lvt__u0_diff_17 = '-2.43906e-05*lvln_mobility*lvln_mobility+5.07813e-04*lvln_mobility+4.62100e-04'
+ sky130_fd_pr__nfet_01v8_lvt__u0_diff_18 = '-2.28106e-05*lvln_mobility*lvln_mobility+3.66405e-04*lvln_mobility+-3.94910e-04'
+ sky130_fd_pr__nfet_01v8_lvt__u0_diff_19 = '-1.00201e-04*lvln_mobility*lvln_mobility+-6.48670e-04*lvln_mobility+-1.74080e-03'
+ sky130_fd_pr__nfet_01v8_lvt__u0_diff_2 = '-3.00291e-05*lvln_mobility*lvln_mobility+-3.85434e-04*lvln_mobility+-1.29460e-03'
+ sky130_fd_pr__nfet_01v8_lvt__u0_diff_20 = '-1.40184e-05*lvln_mobility*lvln_mobility+3.95024e-04*lvln_mobility+1.57340e-03'
+ sky130_fd_pr__nfet_01v8_lvt__u0_diff_21 = '-1.47719e-05*lvln_mobility*lvln_mobility+1.08937e-04*lvln_mobility+1.28280e-03'
+ sky130_fd_pr__nfet_01v8_lvt__u0_diff_22 = '-1.21544e-05*lvln_mobility*lvln_mobility+9.58801e-05*lvln_mobility+6.29700e-04'
+ sky130_fd_pr__nfet_01v8_lvt__u0_diff_23 = '-1.01947e-05*lvln_mobility*lvln_mobility+6.50313e-05*lvln_mobility+8.78370e-04'
+ sky130_fd_pr__nfet_01v8_lvt__u0_diff_24 = '-3.74313e-05*lvln_mobility*lvln_mobility+5.48800e-04*lvln_mobility+-3.23000e-03'
+ sky130_fd_pr__nfet_01v8_lvt__u0_diff_25 = '-1.25669e-05*lvln_mobility*lvln_mobility+7.07800e-04*lvln_mobility+-4.96930e-04'
+ sky130_fd_pr__nfet_01v8_lvt__u0_diff_26 = '-6.45937e-05*lvln_mobility*lvln_mobility+-4.27510e-04*lvln_mobility+-4.89460e-04'
+ sky130_fd_pr__nfet_01v8_lvt__u0_diff_27 = '-1.40362e-05*lvln_mobility*lvln_mobility+3.05595e-04*lvln_mobility+1.19390e-03'
+ sky130_fd_pr__nfet_01v8_lvt__u0_diff_28 = '-1.41781e-04*lvln_mobility*lvln_mobility+-1.39063e-03*lvln_mobility+-2.06260e-03'
+ sky130_fd_pr__nfet_01v8_lvt__u0_diff_29 = '-7.21519e-05*lvln_mobility*lvln_mobility+3.20915e-04*lvln_mobility+-7.93510e-04'
+ sky130_fd_pr__nfet_01v8_lvt__u0_diff_3 = '-4.21187e-06*lvln_mobility*lvln_mobility+7.52375e-04*lvln_mobility+1.62590e-04'
+ sky130_fd_pr__nfet_01v8_lvt__u0_diff_30 = '-7.39863e-05*lvln_mobility*lvln_mobility+4.83988e-04*lvln_mobility+5.02030e-04'
+ sky130_fd_pr__nfet_01v8_lvt__u0_diff_31 = '-1.23581e-05*lvln_mobility*lvln_mobility+3.96567e-04*lvln_mobility+-1.94520e-03'
+ sky130_fd_pr__nfet_01v8_lvt__u0_diff_32 = '-2.41344e-05*lvln_mobility*lvln_mobility+-6.31625e-05*lvln_mobility+-1.33080e-03'
+ sky130_fd_pr__nfet_01v8_lvt__u0_diff_33 = '-3.64437e-05*lvln_mobility*lvln_mobility+1.67300e-04*lvln_mobility+-1.39320e-03'
+ sky130_fd_pr__nfet_01v8_lvt__u0_diff_34 = '-3.54500e-05*lvln_mobility*lvln_mobility+4.06725e-04*lvln_mobility+-2.34620e-03'
+ sky130_fd_pr__nfet_01v8_lvt__u0_diff_35 = '-3.06662e-05*lvln_mobility*lvln_mobility+4.54335e-04*lvln_mobility+-1.86530e-03'
+ sky130_fd_pr__nfet_01v8_lvt__u0_diff_36 = '-3.16563e-05*lvln_mobility*lvln_mobility+5.75500e-04*lvln_mobility+5.08000e-04'
+ sky130_fd_pr__nfet_01v8_lvt__u0_diff_37 = '-6.58597e-05*lvln_mobility*lvln_mobility+-5.49211e-04*lvln_mobility+-1.74940e-03'
+ sky130_fd_pr__nfet_01v8_lvt__u0_diff_4 = '-3.29316e-05*lvln_mobility*lvln_mobility+3.32549e-04*lvln_mobility+-1.46780e-03'
+ sky130_fd_pr__nfet_01v8_lvt__u0_diff_5 = '-1.01594e-04*lvln_mobility*lvln_mobility+-9.45900e-04*lvln_mobility+-7.97300e-04'
+ sky130_fd_pr__nfet_01v8_lvt__u0_diff_6 = '-4.56734e-05*lvln_mobility*lvln_mobility+-1.80359e-04*lvln_mobility+-4.91890e-04'
+ sky130_fd_pr__nfet_01v8_lvt__u0_diff_7 = '-1.95638e-05*lvln_mobility*lvln_mobility+-6.41828e-05*lvln_mobility+6.47410e-04'
+ sky130_fd_pr__nfet_01v8_lvt__u0_diff_8 = '-1.34928e-05*lvln_mobility*lvln_mobility+7.41785e-05*lvln_mobility+4.88970e-04'
+ sky130_fd_pr__nfet_01v8_lvt__u0_diff_9 = '-1.30312e-05*lvln_mobility*lvln_mobility+6.65250e-06*lvln_mobility+-1.53310e-04'
+ sky130_fd_pr__nfet_01v8_lvt__ua_diff_0 = '3.23531e-14*lvln_mobility*lvln_mobility+-3.90095e-13*lvln_mobility+6.43770e-13'
+ sky130_fd_pr__nfet_01v8_lvt__ua_diff_1 = '3.90156e-14*lvln_mobility*lvln_mobility+3.34863e-13*lvln_mobility+3.55080e-12'
+ sky130_fd_pr__nfet_01v8_lvt__ua_diff_10 = '2.48473e-12*lvln_mobility*lvln_mobility+-1.20772e-11*lvln_mobility+3.92450e-12'
+ sky130_fd_pr__nfet_01v8_lvt__ua_diff_11 = '7.85019e-13*lvln_mobility*lvln_mobility+-6.68875e-12*lvln_mobility+1.11470e-12'
+ sky130_fd_pr__nfet_01v8_lvt__ua_diff_12 = '-8.65970e-12*lvln_mobility*lvln_mobility+-1.59774e-11*lvln_mobility+1.64680e-13'
+ sky130_fd_pr__nfet_01v8_lvt__ua_diff_13 = '5.81250e-15*lvln_mobility*lvln_mobility+-7.20700e-13*lvln_mobility+-1.21300e-12'
+ sky130_fd_pr__nfet_01v8_lvt__ua_diff_14 = '2.11500e-14*lvln_mobility*lvln_mobility+-3.26040e-13*lvln_mobility+-6.88440e-13'
+ sky130_fd_pr__nfet_01v8_lvt__ua_diff_15 = '5.05062e-15*lvln_mobility*lvln_mobility+-2.11202e-13*lvln_mobility+-1.49760e-12'
+ sky130_fd_pr__nfet_01v8_lvt__ua_diff_16 = '1.24178e-14*lvln_mobility*lvln_mobility+-1.99791e-13*lvln_mobility+1.86750e-13'
+ sky130_fd_pr__nfet_01v8_lvt__ua_diff_17 = '1.13526e-12*lvln_mobility*lvln_mobility+-9.67137e-12*lvln_mobility+-1.00560e-12'
+ sky130_fd_pr__nfet_01v8_lvt__ua_diff_18 = '1.06420e-12*lvln_mobility*lvln_mobility+-7.09760e-12*lvln_mobility+1.65140e-12'
+ sky130_fd_pr__nfet_01v8_lvt__ua_diff_19 = '-3.09654e-12*lvln_mobility*lvln_mobility+-5.29575e-12*lvln_mobility+3.47870e-12'
+ sky130_fd_pr__nfet_01v8_lvt__ua_diff_2 = '2.05775e-14*lvln_mobility*lvln_mobility+2.79925e-14*lvln_mobility+-6.24430e-13'
+ sky130_fd_pr__nfet_01v8_lvt__ua_diff_20 = '-8.85938e-16*lvln_mobility*lvln_mobility+-7.44656e-13*lvln_mobility+-3.35610e-12'
+ sky130_fd_pr__nfet_01v8_lvt__ua_diff_21 = '5.94688e-15*lvln_mobility*lvln_mobility+-2.73875e-14*lvln_mobility+-2.73720e-12'
+ sky130_fd_pr__nfet_01v8_lvt__ua_diff_22 = '1.48947e-14*lvln_mobility*lvln_mobility+-1.17019e-13*lvln_mobility+-7.01450e-13'
+ sky130_fd_pr__nfet_01v8_lvt__ua_diff_23 = '1.44750e-14*lvln_mobility*lvln_mobility+-1.55275e-13*lvln_mobility+-2.36020e-12'
+ sky130_fd_pr__nfet_01v8_lvt__ua_diff_24 = '-3.85717e-13*lvln_mobility*lvln_mobility+-7.01892e-14*lvln_mobility+6.39210e-12'
+ sky130_fd_pr__nfet_01v8_lvt__ua_diff_25 = '1.76484e-13*lvln_mobility*lvln_mobility+-1.72011e-12*lvln_mobility+2.77980e-12'
+ sky130_fd_pr__nfet_01v8_lvt__ua_diff_26 = '3.49188e-14*lvln_mobility*lvln_mobility+-3.50000e-15*lvln_mobility+1.79840e-12'
+ sky130_fd_pr__nfet_01v8_lvt__ua_diff_27 = '1.90781e-14*lvln_mobility*lvln_mobility+-5.86737e-13*lvln_mobility+-3.95450e-12'
+ sky130_fd_pr__nfet_01v8_lvt__ua_diff_28 = '-2.99312e-14*lvln_mobility*lvln_mobility+6.01250e-14*lvln_mobility+2.82320e-12'
+ sky130_fd_pr__nfet_01v8_lvt__ua_diff_29 = '-3.38898e-12*lvln_mobility*lvln_mobility+-6.19243e-12*lvln_mobility+7.15050e-11'
+ sky130_fd_pr__nfet_01v8_lvt__ua_diff_3 = '3.35049e-12*lvln_mobility*lvln_mobility+5.89087e-12*lvln_mobility+-1.44380e-13'
+ sky130_fd_pr__nfet_01v8_lvt__ua_diff_30 = '5.00950e-13*lvln_mobility*lvln_mobility+-6.26525e-12*lvln_mobility+4.44580e-12'
+ sky130_fd_pr__nfet_01v8_lvt__ua_diff_31 = '1.92415e-12*lvln_mobility*lvln_mobility+-1.20252e-11*lvln_mobility+1.57360e-11'
+ sky130_fd_pr__nfet_01v8_lvt__ua_diff_32 = '6.27485e-12*lvln_mobility*lvln_mobility+-2.96279e-11*lvln_mobility+1.28110e-11'
+ sky130_fd_pr__nfet_01v8_lvt__ua_diff_33 = '1.93873e-12*lvln_mobility*lvln_mobility+-1.06509e-11*lvln_mobility+8.20570e-12'
+ sky130_fd_pr__nfet_01v8_lvt__ua_diff_34 = '3.68572e-14*lvln_mobility*lvln_mobility+1.56125e-15*lvln_mobility+2.80470e-13'
+ sky130_fd_pr__nfet_01v8_lvt__ua_diff_35 = '1.57366e-14*lvln_mobility*lvln_mobility+-1.30449e-13*lvln_mobility+2.41120e-13'
+ sky130_fd_pr__nfet_01v8_lvt__ua_diff_36 = '8.28031e-15*lvln_mobility*lvln_mobility+-1.67366e-13*lvln_mobility+-2.87570e-13'
+ sky130_fd_pr__nfet_01v8_lvt__ua_diff_37 = '8.88580e-13*lvln_mobility*lvln_mobility+3.56654e-12*lvln_mobility+2.21560e-13'
+ sky130_fd_pr__nfet_01v8_lvt__ua_diff_4 = '1.21394e-13*lvln_mobility*lvln_mobility+-2.57740e-12*lvln_mobility+2.72310e-12'
+ sky130_fd_pr__nfet_01v8_lvt__ua_diff_5 = '-8.18859e-13*lvln_mobility*lvln_mobility+-3.90956e-12*lvln_mobility+-1.44400e-12'
+ sky130_fd_pr__nfet_01v8_lvt__ua_diff_6 = '-1.40188e-13*lvln_mobility*lvln_mobility+-1.57715e-12*lvln_mobility+-5.51540e-12'
+ sky130_fd_pr__nfet_01v8_lvt__ua_diff_7 = '1.73319e-14*lvln_mobility*lvln_mobility+-1.79228e-13*lvln_mobility+-1.29770e-12'
+ sky130_fd_pr__nfet_01v8_lvt__ua_diff_8 = '1.40134e-14*lvln_mobility*lvln_mobility+-7.46137e-14*lvln_mobility+4.24790e-13'
+ sky130_fd_pr__nfet_01v8_lvt__ua_diff_9 = '9.35781e-15*lvln_mobility*lvln_mobility+-1.44094e-13*lvln_mobility+-9.09750e-13'
+ sky130_fd_pr__nfet_01v8_lvt__ub_diff_0 = '-3.88122e-21*lvln_mobility*lvln_mobility+-5.34299e-20*lvln_mobility+2.32690e-19'
+ sky130_fd_pr__nfet_01v8_lvt__ub_diff_1 = '-3.42228e-21*lvln_mobility*lvln_mobility+-3.52966e-20*lvln_mobility+1.82120e-19'
+ sky130_fd_pr__nfet_01v8_lvt__ub_diff_10 = '-2.99487e-21*lvln_mobility*lvln_mobility+1.95815e-20*lvln_mobility+-3.28860e-20'
+ sky130_fd_pr__nfet_01v8_lvt__ub_diff_11 = '-1.72731e-21*lvln_mobility*lvln_mobility+-1.02493e-20*lvln_mobility+1.60970e-19'
+ sky130_fd_pr__nfet_01v8_lvt__ub_diff_12 = '3.20400e-21*lvln_mobility*lvln_mobility+-5.06315e-20*lvln_mobility+2.45170e-19'
+ sky130_fd_pr__nfet_01v8_lvt__ub_diff_13 = '-1.62394e-21*lvln_mobility*lvln_mobility+-1.65433e-20*lvln_mobility+1.82520e-19'
+ sky130_fd_pr__nfet_01v8_lvt__ub_diff_14 = '-1.68000e-21*lvln_mobility*lvln_mobility+-1.18825e-20*lvln_mobility+1.78320e-19'
+ sky130_fd_pr__nfet_01v8_lvt__ub_diff_15 = '-1.68428e-21*lvln_mobility*lvln_mobility+-1.58096e-20*lvln_mobility+1.81050e-19'
+ sky130_fd_pr__nfet_01v8_lvt__ub_diff_16 = '-1.47297e-21*lvln_mobility*lvln_mobility+-5.71937e-21*lvln_mobility+1.42120e-19'
+ sky130_fd_pr__nfet_01v8_lvt__ub_diff_17 = '-1.20375e-21*lvln_mobility*lvln_mobility+1.66275e-20*lvln_mobility+1.93080e-19'
+ sky130_fd_pr__nfet_01v8_lvt__ub_diff_18 = '-1.87809e-21*lvln_mobility*lvln_mobility+5.47238e-21*lvln_mobility+1.20880e-19'
+ sky130_fd_pr__nfet_01v8_lvt__ub_diff_19 = '-2.06375e-21*lvln_mobility*lvln_mobility+-6.02625e-20*lvln_mobility+1.60910e-19'
+ sky130_fd_pr__nfet_01v8_lvt__ub_diff_2 = '-2.86156e-21*lvln_mobility*lvln_mobility+-3.10087e-20*lvln_mobility+1.68790e-19'
+ sky130_fd_pr__nfet_01v8_lvt__ub_diff_20 = '-1.41781e-21*lvln_mobility*lvln_mobility+-2.31125e-21*lvln_mobility+2.44270e-19'
+ sky130_fd_pr__nfet_01v8_lvt__ub_diff_21 = '-1.77562e-21*lvln_mobility*lvln_mobility+-1.27100e-20*lvln_mobility+2.04760e-19'
+ sky130_fd_pr__nfet_01v8_lvt__ub_diff_22 = '-1.60084e-21*lvln_mobility*lvln_mobility+-9.44087e-21*lvln_mobility+1.58750e-19'
+ sky130_fd_pr__nfet_01v8_lvt__ub_diff_23 = '-1.32469e-21*lvln_mobility*lvln_mobility+-2.59625e-21*lvln_mobility+2.01510e-19'
+ sky130_fd_pr__nfet_01v8_lvt__ub_diff_24 = '-1.15000e-22*lvln_mobility*lvln_mobility+-9.85000e-22*lvln_mobility+-1.36800e-19'
+ sky130_fd_pr__nfet_01v8_lvt__ub_diff_25 = '-3.87187e-23*lvln_mobility*lvln_mobility+3.39449e-20*lvln_mobility+1.08890e-19'
+ sky130_fd_pr__nfet_01v8_lvt__ub_diff_26 = '-4.07472e-21*lvln_mobility*lvln_mobility+-3.54914e-20*lvln_mobility+2.69840e-19'
+ sky130_fd_pr__nfet_01v8_lvt__ub_diff_27 = '-1.35000e-21*lvln_mobility*lvln_mobility+-1.14750e-21*lvln_mobility+2.11620e-19'
+ sky130_fd_pr__nfet_01v8_lvt__ub_diff_28 = '-1.23722e-20*lvln_mobility*lvln_mobility+-1.17416e-19*lvln_mobility+2.52160e-19'
+ sky130_fd_pr__nfet_01v8_lvt__ub_diff_29 = '2.59725e-21*lvln_mobility*lvln_mobility+-6.67525e-20*lvln_mobility+-3.59960e-20'
+ sky130_fd_pr__nfet_01v8_lvt__ub_diff_3 = '-3.21397e-21*lvln_mobility*lvln_mobility+-2.02784e-20*lvln_mobility+1.67480e-19'
+ sky130_fd_pr__nfet_01v8_lvt__ub_diff_30 = '-4.12284e-21*lvln_mobility*lvln_mobility+-9.60664e-20*lvln_mobility+4.64070e-19'
+ sky130_fd_pr__nfet_01v8_lvt__ub_diff_31 = '1.11187e-21*lvln_mobility*lvln_mobility+1.90450e-20*lvln_mobility+-2.58500e-19'
+ sky130_fd_pr__nfet_01v8_lvt__ub_diff_32 = '-6.02016e-21*lvln_mobility*lvln_mobility+-5.02894e-20*lvln_mobility+-1.46930e-19'
+ sky130_fd_pr__nfet_01v8_lvt__ub_diff_33 = '-1.99953e-21*lvln_mobility*lvln_mobility+-3.53194e-20*lvln_mobility+-1.39090e-19'
+ sky130_fd_pr__nfet_01v8_lvt__ub_diff_34 = '-5.29281e-22*lvln_mobility*lvln_mobility+-7.69688e-21*lvln_mobility+-9.14840e-20'
+ sky130_fd_pr__nfet_01v8_lvt__ub_diff_35 = '-2.14125e-22*lvln_mobility*lvln_mobility+4.22550e-21*lvln_mobility+-3.18000e-20'
+ sky130_fd_pr__nfet_01v8_lvt__ub_diff_36 = '-3.12500e-22*lvln_mobility*lvln_mobility+7.23250e-21*lvln_mobility+2.22680e-19'
+ sky130_fd_pr__nfet_01v8_lvt__ub_diff_37 = '-5.40187e-21*lvln_mobility*lvln_mobility+-6.66650e-20*lvln_mobility+1.56820e-19'
+ sky130_fd_pr__nfet_01v8_lvt__ub_diff_4 = '-1.11956e-21*lvln_mobility*lvln_mobility+-2.72841e-20*lvln_mobility+4.49480e-22'
+ sky130_fd_pr__nfet_01v8_lvt__ub_diff_5 = '-5.92469e-21*lvln_mobility*lvln_mobility+-1.00884e-19*lvln_mobility+1.83830e-19'
+ sky130_fd_pr__nfet_01v8_lvt__ub_diff_6 = '-3.76375e-21*lvln_mobility*lvln_mobility+-5.08225e-20*lvln_mobility+1.27320e-19'
+ sky130_fd_pr__nfet_01v8_lvt__ub_diff_7 = '-2.26207e-21*lvln_mobility*lvln_mobility+-2.68083e-20*lvln_mobility+1.52660e-19'
+ sky130_fd_pr__nfet_01v8_lvt__ub_diff_8 = '-1.60281e-21*lvln_mobility*lvln_mobility+-6.88875e-21*lvln_mobility+1.73150e-19'
+ sky130_fd_pr__nfet_01v8_lvt__ub_diff_9 = '-1.58569e-21*lvln_mobility*lvln_mobility+-9.60525e-21*lvln_mobility+1.06710e-19'
+ sky130_fd_pr__nfet_01v8_lvt__vsat_diff_10 = '-1.00031e+02*lvln_saturation*lvln_saturation+7.57588e+03*lvln_saturation+-7.78010e+02'
+ sky130_fd_pr__nfet_01v8_lvt__vsat_diff_11 = '-2.39563e+00*lvln_saturation*lvln_saturation+5.61650e+03*lvln_saturation+2.21330e+02'
+ sky130_fd_pr__nfet_01v8_lvt__vsat_diff_12 = '1.41525e+02*lvln_saturation*lvln_saturation+4.65038e+03*lvln_saturation+1.20610e+03'
+ sky130_fd_pr__nfet_01v8_lvt__vsat_diff_13 = '8.17563e+01*lvln_saturation*lvln_saturation+4.39412e+03*lvln_saturation+3.58740e+03'
+ sky130_fd_pr__nfet_01v8_lvt__vsat_diff_17 = '-1.23756e+02*lvln_saturation*lvln_saturation+7.07712e+03*lvln_saturation+3.79360e+03'
+ sky130_fd_pr__nfet_01v8_lvt__vsat_diff_18 = '-3.68438e+01*lvln_saturation*lvln_saturation+5.08038e+03*lvln_saturation+-4.51000e+03'
+ sky130_fd_pr__nfet_01v8_lvt__vsat_diff_19 = '1.53488e+02*lvln_saturation*lvln_saturation+4.14275e+03*lvln_saturation+-5.63980e+03'
+ sky130_fd_pr__nfet_01v8_lvt__vsat_diff_20 = '-2.67500e+00*lvln_saturation*lvln_saturation+3.77390e+03*lvln_saturation+5.86820e+03'
+ sky130_fd_pr__nfet_01v8_lvt__vsat_diff_24 = '-2.36017e+02*lvln_saturation*lvln_saturation+6.04750e+03*lvln_saturation+6.93270e+02'
+ sky130_fd_pr__nfet_01v8_lvt__vsat_diff_25 = '2.65625e+01*lvln_saturation*lvln_saturation+5.86838e+03*lvln_saturation+-1.05850e+03'
+ sky130_fd_pr__nfet_01v8_lvt__vsat_diff_26 = '3.59644e+02*lvln_saturation*lvln_saturation+6.03150e+03*lvln_saturation+8.18690e+02'
+ sky130_fd_pr__nfet_01v8_lvt__vsat_diff_27 = '-3.56750e+01*lvln_saturation*lvln_saturation+9.62700e+02*lvln_saturation+-1.09760e+03'
+ sky130_fd_pr__nfet_01v8_lvt__vsat_diff_29 = '4.80025e+02*lvln_saturation*lvln_saturation+1.28522e+04*lvln_saturation+6.64600e+02'
+ sky130_fd_pr__nfet_01v8_lvt__vsat_diff_3 = '3.27812e+01*lvln_saturation*lvln_saturation+8.89738e+03*lvln_saturation+-4.93500e+03'
+ sky130_fd_pr__nfet_01v8_lvt__vsat_diff_30 = '1.00850e+02*lvln_saturation*lvln_saturation+9.04762e+03*lvln_saturation+-3.70710e+03'
+ sky130_fd_pr__nfet_01v8_lvt__vsat_diff_31 = '8.63281e+02*lvln_saturation*lvln_saturation+1.35634e+04*lvln_saturation+-1.00410e+04'
+ sky130_fd_pr__nfet_01v8_lvt__vsat_diff_32 = '-2.10962e+02*lvln_saturation*lvln_saturation+7.99738e+03*lvln_saturation+-1.23210e+03'
+ sky130_fd_pr__nfet_01v8_lvt__vsat_diff_33 = '-1.11363e+02*lvln_saturation*lvln_saturation+6.81800e+03*lvln_saturation+-1.36020e+03'
+ sky130_fd_pr__nfet_01v8_lvt__vsat_diff_34 = '-1.23716e+02*lvln_saturation*lvln_saturation+7.56725e+03*lvln_saturation+2.52460e+02'
+ sky130_fd_pr__nfet_01v8_lvt__vsat_diff_35 = '-1.06119e+02*lvln_saturation*lvln_saturation+7.27888e+03*lvln_saturation+-3.45160e+03'
+ sky130_fd_pr__nfet_01v8_lvt__vsat_diff_36 = '-1.28244e+02*lvln_saturation*lvln_saturation+7.13175e+03*lvln_saturation+3.91490e+03'
+ sky130_fd_pr__nfet_01v8_lvt__vsat_diff_37 = '1.71325e+02*lvln_saturation*lvln_saturation+4.31712e+03*lvln_saturation+-4.16070e+03'
+ sky130_fd_pr__nfet_01v8_lvt__vsat_diff_4 = '5.09125e+01*lvln_saturation*lvln_saturation+6.80012e+03*lvln_saturation+-6.62310e+03'
+ sky130_fd_pr__nfet_01v8_lvt__vsat_diff_5 = '-5.33875e+01*lvln_saturation*lvln_saturation+2.63403e+03*lvln_saturation+-8.60970e+03'
+ sky130_fd_pr__nfet_01v8_lvt__vsat_diff_6 = '1.42425e+02*lvln_saturation*lvln_saturation+6.02062e+03*lvln_saturation+2.48870e+03'
+ sky130_fd_pr__nfet_01v8_lvt__vth0_diff_0 = '-7.12581e-05*lvln_threshold*lvln_threshold+1.16099e-03*lvln_threshold+-4.27890e-03'
+ sky130_fd_pr__nfet_01v8_lvt__vth0_diff_1 = '-4.29156e-05*lvln_threshold*lvln_threshold+9.84113e-04*lvln_threshold+-5.08880e-03'
+ sky130_fd_pr__nfet_01v8_lvt__vth0_diff_10 = '-4.56781e-04*lvln_threshold*lvln_threshold+1.61439e-02*lvln_threshold+-3.94960e-02'
+ sky130_fd_pr__nfet_01v8_lvt__vth0_diff_11 = '-3.74719e-04*lvln_threshold*lvln_threshold+1.30024e-02*lvln_threshold+-2.47600e-02'
+ sky130_fd_pr__nfet_01v8_lvt__vth0_diff_12 = '-3.19275e-04*lvln_threshold*lvln_threshold+5.20225e-03*lvln_threshold+-3.99160e-03'
+ sky130_fd_pr__nfet_01v8_lvt__vth0_diff_13 = '-2.47844e-05*lvln_threshold*lvln_threshold+1.46319e-03*lvln_threshold+-3.86670e-03'
+ sky130_fd_pr__nfet_01v8_lvt__vth0_diff_14 = '-1.44500e-05*lvln_threshold*lvln_threshold+5.80750e-04*lvln_threshold+-6.75860e-03'
+ sky130_fd_pr__nfet_01v8_lvt__vth0_diff_15 = '-1.30125e-05*lvln_threshold*lvln_threshold+-3.71287e-04*lvln_threshold+-2.64250e-04'
+ sky130_fd_pr__nfet_01v8_lvt__vth0_diff_16 = '-1.59250e-05*lvln_threshold*lvln_threshold+7.47000e-04*lvln_threshold+-8.16220e-03'
+ sky130_fd_pr__nfet_01v8_lvt__vth0_diff_17 = '-4.03969e-04*lvln_threshold*lvln_threshold+1.57459e-02*lvln_threshold+-2.74230e-02'
+ sky130_fd_pr__nfet_01v8_lvt__vth0_diff_18 = '-3.69219e-04*lvln_threshold*lvln_threshold+1.21114e-02*lvln_threshold+-1.12530e-02'
+ sky130_fd_pr__nfet_01v8_lvt__vth0_diff_19 = '-2.38881e-04*lvln_threshold*lvln_threshold+4.18448e-03*lvln_threshold+-1.54580e-02'
+ sky130_fd_pr__nfet_01v8_lvt__vth0_diff_2 = '-3.97187e-05*lvln_threshold*lvln_threshold+-1.92825e-04*lvln_threshold+-5.06750e-03'
+ sky130_fd_pr__nfet_01v8_lvt__vth0_diff_20 = '-2.76094e-05*lvln_threshold*lvln_threshold+9.04612e-04*lvln_threshold+-8.77380e-03'
+ sky130_fd_pr__nfet_01v8_lvt__vth0_diff_21 = '-1.05902e-05*lvln_threshold*lvln_threshold+1.07378e-04*lvln_threshold+5.54920e-04'
+ sky130_fd_pr__nfet_01v8_lvt__vth0_diff_22 = '-9.80625e-06*lvln_threshold*lvln_threshold+2.71650e-04*lvln_threshold+-4.72750e-03'
+ sky130_fd_pr__nfet_01v8_lvt__vth0_diff_23 = '-1.79844e-05*lvln_threshold*lvln_threshold+1.22763e-04*lvln_threshold+-3.91200e-03'
+ sky130_fd_pr__nfet_01v8_lvt__vth0_diff_24 = '-2.90531e-04*lvln_threshold*lvln_threshold+1.53124e-02*lvln_threshold+-4.51820e-02'
+ sky130_fd_pr__nfet_01v8_lvt__vth0_diff_25 = '-3.66353e-04*lvln_threshold*lvln_threshold+7.85734e-03*lvln_threshold+-2.25100e-02'
+ sky130_fd_pr__nfet_01v8_lvt__vth0_diff_26 = '-2.06312e-04*lvln_threshold*lvln_threshold+2.19175e-03*lvln_threshold+-1.21990e-02'
+ sky130_fd_pr__nfet_01v8_lvt__vth0_diff_27 = '-2.39075e-05*lvln_threshold*lvln_threshold+7.17170e-04*lvln_threshold+-3.00640e-03'
+ sky130_fd_pr__nfet_01v8_lvt__vth0_diff_28 = '-4.56762e-04*lvln_threshold*lvln_threshold+2.40400e-03*lvln_threshold+-9.03780e-03'
+ sky130_fd_pr__nfet_01v8_lvt__vth0_diff_29 = '-6.38187e-04*lvln_threshold*lvln_threshold+3.10375e-02*lvln_threshold+-2.64690e-02'
+ sky130_fd_pr__nfet_01v8_lvt__vth0_diff_3 = '-3.83128e-04*lvln_threshold*lvln_threshold+1.97771e-02*lvln_threshold+-2.43460e-04'
+ sky130_fd_pr__nfet_01v8_lvt__vth0_diff_30 = '-4.63062e-04*lvln_threshold*lvln_threshold+2.07850e-02*lvln_threshold+-4.47810e-02'
+ sky130_fd_pr__nfet_01v8_lvt__vth0_diff_31 = '-5.34375e-04*lvln_threshold*lvln_threshold+3.65425e-02*lvln_threshold+-2.85300e-02'
+ sky130_fd_pr__nfet_01v8_lvt__vth0_diff_32 = '-5.15531e-04*lvln_threshold*lvln_threshold+3.42974e-02*lvln_threshold+-3.53320e-02'
+ sky130_fd_pr__nfet_01v8_lvt__vth0_diff_33 = '-5.55250e-04*lvln_threshold*lvln_threshold+3.38413e-02*lvln_threshold+-2.74810e-02'
+ sky130_fd_pr__nfet_01v8_lvt__vth0_diff_34 = '-3.44563e-04*lvln_threshold*lvln_threshold+2.10698e-02*lvln_threshold+-2.65980e-02'
+ sky130_fd_pr__nfet_01v8_lvt__vth0_diff_35 = '-3.37188e-04*lvln_threshold*lvln_threshold+1.56512e-02*lvln_threshold+-3.72500e-02'
+ sky130_fd_pr__nfet_01v8_lvt__vth0_diff_36 = '-4.17688e-04*lvln_threshold*lvln_threshold+1.56768e-02*lvln_threshold+-2.51020e-02'
+ sky130_fd_pr__nfet_01v8_lvt__vth0_diff_37 = '-2.14734e-04*lvln_threshold*lvln_threshold+4.24656e-03*lvln_threshold+-1.08830e-02'
+ sky130_fd_pr__nfet_01v8_lvt__vth0_diff_4 = '-4.36313e-04*lvln_threshold*lvln_threshold+1.66855e-02*lvln_threshold+-3.33570e-02'
+ sky130_fd_pr__nfet_01v8_lvt__vth0_diff_5 = '-6.77606e-04*lvln_threshold*lvln_threshold+4.28337e-03*lvln_threshold+5.83420e-03'
+ sky130_fd_pr__nfet_01v8_lvt__vth0_diff_6 = '-1.42826e-04*lvln_threshold*lvln_threshold+1.81757e-03*lvln_threshold+-5.20750e-03'
+ sky130_fd_pr__nfet_01v8_lvt__vth0_diff_7 = '-2.34403e-05*lvln_threshold*lvln_threshold+1.21741e-04*lvln_threshold+3.58670e-04'
+ sky130_fd_pr__nfet_01v8_lvt__vth0_diff_8 = '-1.60750e-05*lvln_threshold*lvln_threshold+-3.93750e-05*lvln_threshold+-5.90520e-03'
+ sky130_fd_pr__nfet_01v8_lvt__vth0_diff_9 = '-1.65250e-05*lvln_threshold*lvln_threshold+-7.14025e-04*lvln_threshold+-2.43500e-03'
+ sky130_fd_pr__nfet_01v8_lvt__wint_diff = '8.04375e-09*diff_cd'
+ sky130_fd_pr__special_nfet_pass_lvt__ajunction_mult = '-2.59375e-05*lvn_diode*lvn_diode+4.38787e-02*lvn_diode+1.00040e+00'
+ sky130_fd_pr__special_nfet_pass_lvt__dlc_diff = '-4.91625e-11*poly_cd*poly_cd+3.37112e-09*poly_cd+-1.36190e-09'
+ sky130_fd_pr__special_nfet_pass_lvt__dwc_diff = '8.04375e-09*diff_cd'
+ sky130_fd_pr__special_nfet_pass_lvt__lint_diff = '4.33125e-09*poly_cd'
+ sky130_fd_pr__special_nfet_pass_lvt__nfactor_diff_0 = '-2.46134e-02*lvn_subvt*lvn_subvt+1.00321e-01*lvn_subvt+3.97550e-01'
+ sky130_fd_pr__special_nfet_pass_lvt__overlap_mult = '-2.39062e-04*lvtox*lvtox+1.49487e-02*lvtox+9.24290e-01'
+ sky130_fd_pr__special_nfet_pass_lvt__pjunction_mult = '4.43125e-04*lvn_diode*lvn_diode+3.72125e-02*lvn_diode+8.91760e-01'
+ sky130_fd_pr__special_nfet_pass_lvt__rshn_mult = '5.00000e-02*special_nfet_pass_lvt+1.00000e+00'
+ sky130_fd_pr__special_nfet_pass_lvt__toxe_mult = '1.30000e-02*lvtox+1.00000e+00'
+ sky130_fd_pr__special_nfet_pass_lvt__u0_diff_0 = '-3.63906e-05*lvln_mobility*lvln_mobility+3.15216e-03*lvln_mobility+-6.97310e-03'
+ sky130_fd_pr__special_nfet_pass_lvt__vsat_diff_0 = '6.84562e+01*lvln_saturation*lvln_saturation+1.18361e+04*lvln_saturation+8.11120e+03'
+ sky130_fd_pr__special_nfet_pass_lvt__vth0_diff_0 = '5.66969e-04*lvln_threshold*lvln_threshold+3.27404e-02*lvln_threshold+2.47670e-02'
+ sky130_fd_pr__special_nfet_pass_lvt__wint_diff = '8.04375e-09*diff_cd'
+ sky130_fd_pr__special_nfet_pass__ajunction_mult = '9.37500e-07*lvn_diode*lvn_diode+3.87638e-02*lvn_diode+9.95430e-01'
+ sky130_fd_pr__special_nfet_pass__dlc_diff = '-3.03188e-09*poly_cd'
+ sky130_fd_pr__special_nfet_pass__dwc_diff = '5.63000e-09*diff_cd'
+ sky130_fd_pr__special_nfet_pass__lint_diff = '-3.03188e-09*poly_cd'
+ sky130_fd_pr__special_nfet_pass__overlap_mult = '-1.27188e-04*lvtox*lvtox+8.00875e-03*lvtox+9.84200e-01'
+ sky130_fd_pr__special_nfet_pass__pjunction_mult = '-9.37500e-07*lvn_diode*lvn_diode+3.97287e-02*lvn_diode+1.02040e+00'
+ sky130_fd_pr__special_nfet_pass__tox_mult = '9.12500e-03*lvtox+1.00000e+00'
+ sky130_fd_pr__special_nfet_pass__u0_diff_0 = '3.55678e-04*lvn_mobility*lvn_mobility+3.05794e-03*lvn_mobility+-2.92260e-03'
+ sky130_fd_pr__special_nfet_pass__vth0_diff_0 = '-2.68250e-04*lvn_threshold*lvn_threshold+4.27650e-02*lvn_threshold+2.75220e-02'
+ sky130_fd_pr__special_nfet_pass__wint_diff = '5.63000e-09*diff_cd'
+ sky130_fd_pr__special_nfet_latch__ajunction_mult = '9.37500e-07*lvn_diode*lvn_diode+3.87638e-02*lvn_diode+9.95430e-01'
+ sky130_fd_pr__special_nfet_latch__dlc_diff = '-3.03188e-09*poly_cd'
+ sky130_fd_pr__special_nfet_latch__dwc_diff = '5.63000e-09*diff_cd'
+ sky130_fd_pr__special_nfet_latch__lint_diff = '-3.03188e-09*poly_cd'
+ sky130_fd_pr__special_nfet_latch__overlap_mult = '-1.27188e-04*lvtox*lvtox+8.00875e-03*lvtox+9.84200e-01'
+ sky130_fd_pr__special_nfet_latch__pjunction_mult = '-9.37500e-07*lvn_diode*lvn_diode+3.97287e-02*lvn_diode+1.02040e+00'
+ sky130_fd_pr__special_nfet_latch__tox_mult = '9.12500e-03*lvtox+1.00000e+00'
+ sky130_fd_pr__special_nfet_latch__u0_diff_0 = '6.25750e-06*lvn_mobility*lvn_mobility+2.32240e-03*lvn_mobility+3.03680e-04'
+ sky130_fd_pr__special_nfet_latch__vth0_diff_0 = '-9.35625e-05*lvn_threshold*lvn_threshold+3.22038e-02*lvn_threshold+2.09520e-02'
+ sky130_fd_pr__special_nfet_latch__wint_diff = '5.63000e-09*diff_cd'
+ sky130_fd_pr__nfet_01v8__a0_diff_11 = '3.67969e-04*lvn_saturation*lvn_saturation+-8.67875e-04*lvn_saturation+1.64720e-02'
+ sky130_fd_pr__nfet_01v8__a0_diff_12 = '6.65219e-04*lvn_saturation*lvn_saturation+5.39312e-03*lvn_saturation+4.47690e-02'
+ sky130_fd_pr__nfet_01v8__a0_diff_13 = '3.04491e-03*lvn_saturation*lvn_saturation+1.40759e-02*lvn_saturation+2.16880e-02'
+ sky130_fd_pr__nfet_01v8__a0_diff_14 = '5.19531e-04*lvn_saturation*lvn_saturation+3.75538e-03*lvn_saturation+4.22500e-02'
+ sky130_fd_pr__nfet_01v8__a0_diff_19 = '-8.78438e-05*lvn_saturation*lvn_saturation+-2.64375e-04*lvn_saturation+1.37280e-02'
+ sky130_fd_pr__nfet_01v8__a0_diff_2 = '3.24813e-04*lvn_saturation*lvn_saturation+-4.01708e-02*lvn_saturation+2.34120e-01'
+ sky130_fd_pr__nfet_01v8__a0_diff_20 = '8.89375e-04*lvn_saturation*lvn_saturation+5.34350e-03*lvn_saturation+3.90450e-02'
+ sky130_fd_pr__nfet_01v8__a0_diff_21 = '5.39094e-04*lvn_saturation*lvn_saturation+6.08238e-03*lvn_saturation+6.58450e-02'
+ sky130_fd_pr__nfet_01v8__a0_diff_22 = '5.14556e-04*lvn_saturation*lvn_saturation+3.49980e-03*lvn_saturation+8.66190e-03'
+ sky130_fd_pr__nfet_01v8__a0_diff_27 = '9.21281e-04*lvn_saturation*lvn_saturation+-9.08375e-04*lvn_saturation+6.61330e-02'
+ sky130_fd_pr__nfet_01v8__a0_diff_28 = '7.51656e-04*lvn_saturation*lvn_saturation+1.18891e-02*lvn_saturation+4.06470e-02'
+ sky130_fd_pr__nfet_01v8__a0_diff_29 = '5.38228e-04*lvn_saturation*lvn_saturation+4.58516e-03*lvn_saturation+-2.12760e-02'
+ sky130_fd_pr__nfet_01v8__a0_diff_3 = '9.32625e-04*lvn_saturation*lvn_saturation+-2.31588e-02*lvn_saturation+3.06930e-02'
+ sky130_fd_pr__nfet_01v8__a0_diff_30 = '4.59594e-04*lvn_saturation*lvn_saturation+6.86962e-03*lvn_saturation+1.46190e-02'
+ sky130_fd_pr__nfet_01v8__a0_diff_4 = '9.22750e-04*lvn_saturation*lvn_saturation+-2.91350e-03*lvn_saturation+3.43960e-02'
+ sky130_fd_pr__nfet_01v8__a0_diff_5 = '6.45531e-04*lvn_saturation*lvn_saturation+-1.23063e-03*lvn_saturation+4.38220e-02'
+ sky130_fd_pr__nfet_01v8__ags_diff_11 = '-1.73869e-03*lvn_saturation*lvn_saturation+2.58087e-02*lvn_saturation+-2.90260e-02'
+ sky130_fd_pr__nfet_01v8__ags_diff_12 = '-4.93875e-04*lvn_saturation*lvn_saturation+-5.54525e-03*lvn_saturation+-3.79560e-02'
+ sky130_fd_pr__nfet_01v8__ags_diff_13 = '4.31968e-04*lvn_saturation*lvn_saturation+-1.53185e-03*lvn_saturation+-1.74090e-03'
+ sky130_fd_pr__nfet_01v8__ags_diff_14 = '-2.70097e-04*lvn_saturation*lvn_saturation+-4.36786e-03*lvn_saturation+-2.27340e-02'
+ sky130_fd_pr__nfet_01v8__ags_diff_19 = '-1.04715e-03*lvn_saturation*lvn_saturation+-2.27879e-03*lvn_saturation+4.47060e-03'
+ sky130_fd_pr__nfet_01v8__ags_diff_2 = '-2.98569e-03*lvn_saturation*lvn_saturation+2.21567e-02*lvn_saturation+-5.28720e-02'
+ sky130_fd_pr__nfet_01v8__ags_diff_20 = '-3.99281e-04*lvn_saturation*lvn_saturation+-2.94388e-03*lvn_saturation+-1.69250e-02'
+ sky130_fd_pr__nfet_01v8__ags_diff_21 = '-2.76750e-04*lvn_saturation*lvn_saturation+-4.47300e-03*lvn_saturation+-4.74760e-02'
+ sky130_fd_pr__nfet_01v8__ags_diff_22 = '-2.42650e-04*lvn_saturation*lvn_saturation+-3.64775e-03*lvn_saturation+6.58540e-03'
+ sky130_fd_pr__nfet_01v8__ags_diff_27 = '-8.62656e-04*lvn_saturation*lvn_saturation+1.41487e-03*lvn_saturation+-5.63720e-02'
+ sky130_fd_pr__nfet_01v8__ags_diff_28 = '-3.73075e-04*lvn_saturation*lvn_saturation+-9.30645e-03*lvn_saturation+-2.43290e-02'
+ sky130_fd_pr__nfet_01v8__ags_diff_29 = '-2.43719e-04*lvn_saturation*lvn_saturation+-2.97937e-03*lvn_saturation+2.29170e-02'
+ sky130_fd_pr__nfet_01v8__ags_diff_3 = '-5.90388e-04*lvn_saturation*lvn_saturation+1.30913e-02*lvn_saturation+-8.64580e-03'
+ sky130_fd_pr__nfet_01v8__ags_diff_30 = '-2.11113e-04*lvn_saturation*lvn_saturation+-5.44163e-03*lvn_saturation+-1.80700e-04'
+ sky130_fd_pr__nfet_01v8__ags_diff_4 = '-4.42016e-04*lvn_saturation*lvn_saturation+2.45219e-03*lvn_saturation+-1.13910e-02'
+ sky130_fd_pr__nfet_01v8__ags_diff_5 = '-3.79438e-04*lvn_saturation*lvn_saturation+2.40125e-03*lvn_saturation+-1.83730e-02'
+ sky130_fd_pr__nfet_01v8__ajunction_mult = '-1.87500e-06*lvn_diode*lvn_diode+5.53750e-02*lvn_diode+9.95430e-01'
+ sky130_fd_pr__nfet_01v8__b0_diff_35 = '1.49206e-09*lvn_saturation*lvn_saturation+-3.40957e-08*lvn_saturation+-1.41470e-07'
+ sky130_fd_pr__nfet_01v8__b0_diff_36 = '9.53875e-10*lvn_saturation*lvn_saturation+-1.32235e-08*lvn_saturation+2.33280e-08'
+ sky130_fd_pr__nfet_01v8__b0_diff_37 = '1.66556e-09*lvn_saturation*lvn_saturation+-2.90920e-08*lvn_saturation+4.25530e-08'
+ sky130_fd_pr__nfet_01v8__b0_diff_38 = '1.17094e-09*lvn_saturation*lvn_saturation+-1.90767e-08*lvn_saturation+4.05090e-09'
+ sky130_fd_pr__nfet_01v8__b0_diff_39 = '1.01979e-09*lvn_saturation*lvn_saturation+-1.39236e-08*lvn_saturation+3.94090e-08'
+ sky130_fd_pr__nfet_01v8__b0_diff_40 = '-2.14281e-08*lvn_saturation*lvn_saturation+-2.32050e-08*lvn_saturation'
+ sky130_fd_pr__nfet_01v8__b0_diff_41 = '3.12511e-08*lvn_saturation*lvn_saturation+-1.42596e-07*lvn_saturation'
+ sky130_fd_pr__nfet_01v8__b0_diff_42 = '6.36281e-09*lvn_saturation*lvn_saturation+-6.14762e-08*lvn_saturation'
+ sky130_fd_pr__nfet_01v8__b0_diff_43 = '2.70466e-09*lvn_saturation*lvn_saturation+-3.48314e-08*lvn_saturation+1.14180e-07'
+ sky130_fd_pr__nfet_01v8__b0_diff_44 = '1.58822e-09*lvn_saturation*lvn_saturation+-2.76301e-08*lvn_saturation+6.61280e-08'
+ sky130_fd_pr__nfet_01v8__b0_diff_45 = '1.22031e-09*lvn_saturation*lvn_saturation+-2.18563e-08*lvn_saturation+3.31900e-08'
+ sky130_fd_pr__nfet_01v8__b0_diff_46 = '1.02753e-09*lvn_saturation*lvn_saturation+-1.41096e-08*lvn_saturation+2.19740e-08'
+ sky130_fd_pr__nfet_01v8__b0_diff_47 = '-1.30375e-09*lvn_saturation*lvn_saturation+-1.19735e-07*lvn_saturation'
+ sky130_fd_pr__nfet_01v8__b0_diff_50 = '1.06494e-08*lvn_saturation*lvn_saturation+-1.00063e-07*lvn_saturation'
+ sky130_fd_pr__nfet_01v8__b0_diff_51 = '5.92856e-09*lvn_saturation*lvn_saturation+-5.69935e-08*lvn_saturation'
+ sky130_fd_pr__nfet_01v8__b0_diff_52 = '-3.51168e-08*lvn_saturation*lvn_saturation+4.45300e-08*lvn_saturation'
+ sky130_fd_pr__nfet_01v8__b0_diff_53 = '-2.77995e-08*lvn_saturation*lvn_saturation+8.08000e-09*lvn_saturation'
+ sky130_fd_pr__nfet_01v8__b0_diff_54 = '-5.11553e-09*lvn_saturation*lvn_saturation+-1.01686e-07*lvn_saturation'
+ sky130_fd_pr__nfet_01v8__b0_diff_55 = '-2.53025e-09*lvn_saturation*lvn_saturation+-1.13938e-07*lvn_saturation'
+ sky130_fd_pr__nfet_01v8__b0_diff_56 = '-6.83937e-10*lvn_saturation*lvn_saturation+-7.52690e-08*lvn_saturation'
+ sky130_fd_pr__nfet_01v8__b0_diff_57 = '-3.86469e-10*lvn_saturation*lvn_saturation+-4.83431e-08*lvn_saturation'
+ sky130_fd_pr__nfet_01v8__b0_diff_58 = '-2.66219e-10*lvn_saturation*lvn_saturation+-3.56064e-08*lvn_saturation'
+ sky130_fd_pr__nfet_01v8__b0_diff_59 = '6.59159e-10*lvn_saturation*lvn_saturation+-6.51724e-09*lvn_saturation'
+ sky130_fd_pr__nfet_01v8__b0_diff_60 = '6.59159e-10*lvn_saturation*lvn_saturation+-6.51724e-09*lvn_saturation'
+ sky130_fd_pr__nfet_01v8__b0_diff_62 = '1.06126e-18*lvn_saturation*lvn_saturation+-9.39251e-18*lvn_saturation'
+ sky130_fd_pr__nfet_01v8__b1_diff_35 = '6.83684e-10*lvn_saturation*lvn_saturation+1.54376e-09*lvn_saturation+4.95200e-09'
+ sky130_fd_pr__nfet_01v8__b1_diff_36 = '1.92562e-10*lvn_saturation*lvn_saturation+1.34565e-09*lvn_saturation+3.91140e-09'
+ sky130_fd_pr__nfet_01v8__b1_diff_37 = '4.09550e-10*lvn_saturation*lvn_saturation+-2.03750e-10*lvn_saturation+8.16020e-09'
+ sky130_fd_pr__nfet_01v8__b1_diff_38 = '-1.52253e-10*lvn_saturation*lvn_saturation+4.96212e-10*lvn_saturation+5.78290e-09'
+ sky130_fd_pr__nfet_01v8__b1_diff_39 = '-3.17594e-11*lvn_saturation*lvn_saturation+3.49738e-10*lvn_saturation+3.43480e-09'
+ sky130_fd_pr__nfet_01v8__b1_diff_40 = '1.13437e-08*lvn_saturation*lvn_saturation+3.96652e-08*lvn_saturation'
+ sky130_fd_pr__nfet_01v8__b1_diff_41 = '-8.04969e-10*lvn_saturation*lvn_saturation+-7.31413e-09*lvn_saturation'
+ sky130_fd_pr__nfet_01v8__b1_diff_42 = '5.73969e-10*lvn_saturation*lvn_saturation+9.35375e-10*lvn_saturation'
+ sky130_fd_pr__nfet_01v8__b1_diff_43 = '1.04818e-09*lvn_saturation*lvn_saturation+2.92948e-09*lvn_saturation+2.20320e-09'
+ sky130_fd_pr__nfet_01v8__b1_diff_44 = '1.55447e-10*lvn_saturation*lvn_saturation+1.20824e-09*lvn_saturation+8.04990e-09'
+ sky130_fd_pr__nfet_01v8__b1_diff_45 = '2.67438e-11*lvn_saturation*lvn_saturation+1.36925e-10*lvn_saturation+3.34370e-09'
+ sky130_fd_pr__nfet_01v8__b1_diff_46 = '6.36900e-11*lvn_saturation*lvn_saturation+5.54465e-10*lvn_saturation+1.96690e-09'
+ sky130_fd_pr__nfet_01v8__b1_diff_47 = '3.60744e-09*lvn_saturation*lvn_saturation+1.02280e-08*lvn_saturation'
+ sky130_fd_pr__nfet_01v8__b1_diff_50 = '4.89452e-09*lvn_saturation*lvn_saturation+1.97819e-08*lvn_saturation'
+ sky130_fd_pr__nfet_01v8__b1_diff_51 = '2.83486e-09*lvn_saturation*lvn_saturation+1.14548e-08*lvn_saturation'
+ sky130_fd_pr__nfet_01v8__b1_diff_52 = '1.75849e-08*lvn_saturation*lvn_saturation+6.35869e-08*lvn_saturation'
+ sky130_fd_pr__nfet_01v8__b1_diff_53 = '1.41344e-08*lvn_saturation*lvn_saturation+5.03446e-08*lvn_saturation'
+ sky130_fd_pr__nfet_01v8__b1_diff_54 = '4.96185e-09*lvn_saturation*lvn_saturation+1.53621e-08*lvn_saturation'
+ sky130_fd_pr__nfet_01v8__b1_diff_55 = '4.03811e-09*lvn_saturation*lvn_saturation+1.18596e-08*lvn_saturation'
+ sky130_fd_pr__nfet_01v8__b1_diff_56 = '2.25685e-09*lvn_saturation*lvn_saturation+6.36614e-09*lvn_saturation'
+ sky130_fd_pr__nfet_01v8__b1_diff_57 = '1.44527e-09*lvn_saturation*lvn_saturation+4.06406e-09*lvn_saturation'
+ sky130_fd_pr__nfet_01v8__b1_diff_58 = '1.06301e-09*lvn_saturation*lvn_saturation+2.98470e-09*lvn_saturation'
+ sky130_fd_pr__nfet_01v8__b1_diff_59 = '3.30612e-10*lvn_saturation*lvn_saturation+1.33553e-09*lvn_saturation'
+ sky130_fd_pr__nfet_01v8__b1_diff_60 = '3.30612e-10*lvn_saturation*lvn_saturation+1.33553e-09*lvn_saturation'
+ sky130_fd_pr__nfet_01v8__b1_diff_62 = '-4.38675e-19*lvn_saturation*lvn_saturation+-1.20933e-18*lvn_saturation'
+ sky130_fd_pr__nfet_01v8__dlc_diff = '-1.06849e-10*poly_cd*poly_cd+-3.77438e-09*poly_cd+-6.14920e-10'
+ sky130_fd_pr__nfet_01v8__dwc_diff = '8.04375e-09*diff_cd'
+ sky130_fd_pr__nfet_01v8__eta0_diff_51 = '-4.71629e-18*lvn_threshold*lvn_threshold+-6.72209e-18*lvn_threshold'
+ sky130_fd_pr__nfet_01v8__eta0_diff_52 = '1.01678e-06*lvn_threshold*lvn_threshold+-4.06712e-06*lvn_threshold'
+ sky130_fd_pr__nfet_01v8__eta0_diff_53 = '3.62462e-07*lvn_threshold*lvn_threshold+-1.44985e-06*lvn_threshold'
+ sky130_fd_pr__nfet_01v8__eta0_diff_54 = '3.90850e-08*lvn_threshold*lvn_threshold+1.15713e-06*lvn_threshold'
+ sky130_fd_pr__nfet_01v8__eta0_diff_55 = '1.37988e-08*lvn_threshold*lvn_threshold+4.25668e-07*lvn_threshold'
+ sky130_fd_pr__nfet_01v8__eta0_diff_56 = '-2.36359e-08*lvn_threshold*lvn_threshold+-7.87924e-07*lvn_threshold'
+ sky130_fd_pr__nfet_01v8__eta0_diff_57 = '-2.35059e-08*lvn_threshold*lvn_threshold+-8.12811e-07*lvn_threshold'
+ sky130_fd_pr__nfet_01v8__eta0_diff_58 = '-2.00447e-08*lvn_threshold*lvn_threshold+-7.05589e-07*lvn_threshold'
+ sky130_fd_pr__nfet_01v8__eta0_diff_59 = '-2.26278e-19*lvn_threshold*lvn_threshold+1.12122e-17*lvn_threshold'
+ sky130_fd_pr__nfet_01v8__eta0_diff_60 = '3.18769e-13*lvn_threshold*lvn_threshold+7.26373e-12*lvn_threshold'
+ sky130_fd_pr__nfet_01v8__k2_diff_0 = '3.05637e-04*lvn_bodyeffect*lvn_bodyeffect+-8.07963e-03*lvn_bodyeffect+3.18430e-03'
+ sky130_fd_pr__nfet_01v8__k2_diff_1 = '3.03088e-04*lvn_bodyeffect*lvn_bodyeffect+-7.01887e-03*lvn_bodyeffect+4.71710e-03'
+ sky130_fd_pr__nfet_01v8__k2_diff_10 = '3.04575e-04*lvn_bodyeffect*lvn_bodyeffect+-8.26013e-03*lvn_bodyeffect+3.60330e-03'
+ sky130_fd_pr__nfet_01v8__k2_diff_11 = '6.91875e-06*lvn_bodyeffect*lvn_bodyeffect+-4.54975e-04*lvn_bodyeffect+-3.17990e-03'
+ sky130_fd_pr__nfet_01v8__k2_diff_12 = '-2.86250e-06*lvn_bodyeffect*lvn_bodyeffect+5.47500e-05*lvn_bodyeffect+3.25700e-03'
+ sky130_fd_pr__nfet_01v8__k2_diff_13 = '1.76625e-05*lvn_bodyeffect*lvn_bodyeffect+-4.17825e-04*lvn_bodyeffect+3.33930e-03'
+ sky130_fd_pr__nfet_01v8__k2_diff_14 = '7.40000e-06*lvn_bodyeffect*lvn_bodyeffect+-4.53275e-04*lvn_bodyeffect+4.55990e-03'
+ sky130_fd_pr__nfet_01v8__k2_diff_15 = '2.85375e-04*lvn_bodyeffect*lvn_bodyeffect+-8.07800e-03*lvn_bodyeffect+1.04640e-02'
+ sky130_fd_pr__nfet_01v8__k2_diff_16 = '7.51063e-05*lvn_bodyeffect*lvn_bodyeffect+-5.72575e-03*lvn_bodyeffect+9.84030e-03'
+ sky130_fd_pr__nfet_01v8__k2_diff_17 = '-4.65625e-07*lvn_bodyeffect*lvn_bodyeffect+-2.22731e-03*lvn_bodyeffect+7.23320e-03'
+ sky130_fd_pr__nfet_01v8__k2_diff_18 = '-5.45000e-06*lvn_bodyeffect*lvn_bodyeffect+-3.39450e-04*lvn_bodyeffect+3.25310e-03'
+ sky130_fd_pr__nfet_01v8__k2_diff_19 = '-2.41875e-06*lvn_bodyeffect*lvn_bodyeffect+5.49000e-05*lvn_bodyeffect+5.13730e-03'
+ sky130_fd_pr__nfet_01v8__k2_diff_2 = '1.46875e-05*lvn_bodyeffect*lvn_bodyeffect+-4.69625e-04*lvn_bodyeffect+-6.62380e-03'
+ sky130_fd_pr__nfet_01v8__k2_diff_20 = '-2.14375e-06*lvn_bodyeffect*lvn_bodyeffect+1.44750e-04*lvn_bodyeffect+3.58390e-03'
+ sky130_fd_pr__nfet_01v8__k2_diff_21 = '-2.48750e-06*lvn_bodyeffect*lvn_bodyeffect+1.84250e-04*lvn_bodyeffect+3.18590e-03'
+ sky130_fd_pr__nfet_01v8__k2_diff_22 = '7.01250e-06*lvn_bodyeffect*lvn_bodyeffect+-4.18850e-04*lvn_bodyeffect+5.08360e-03'
+ sky130_fd_pr__nfet_01v8__k2_diff_23 = '2.68019e-04*lvn_bodyeffect*lvn_bodyeffect+-7.72088e-03*lvn_bodyeffect+3.42220e-03'
+ sky130_fd_pr__nfet_01v8__k2_diff_24 = '6.38563e-05*lvn_bodyeffect*lvn_bodyeffect+-5.46987e-03*lvn_bodyeffect+8.84780e-03'
+ sky130_fd_pr__nfet_01v8__k2_diff_25 = '3.01250e-06*lvn_bodyeffect*lvn_bodyeffect+-2.25387e-03*lvn_bodyeffect+5.63730e-03'
+ sky130_fd_pr__nfet_01v8__k2_diff_26 = '-8.35000e-06*lvn_bodyeffect*lvn_bodyeffect+-1.67500e-05*lvn_bodyeffect+2.32370e-03'
+ sky130_fd_pr__nfet_01v8__k2_diff_27 = '1.26562e-06*lvn_bodyeffect*lvn_bodyeffect+-1.31663e-04*lvn_bodyeffect+3.16510e-03'
+ sky130_fd_pr__nfet_01v8__k2_diff_28 = '4.65625e-07*lvn_bodyeffect*lvn_bodyeffect+-9.56250e-06*lvn_bodyeffect+4.32460e-03'
+ sky130_fd_pr__nfet_01v8__k2_diff_29 = '-2.27187e-06*lvn_bodyeffect*lvn_bodyeffect+1.20212e-04*lvn_bodyeffect+2.66230e-03'
+ sky130_fd_pr__nfet_01v8__k2_diff_3 = '7.65625e-06*lvn_bodyeffect*lvn_bodyeffect+-2.78600e-04*lvn_bodyeffect+-5.27070e-03'
+ sky130_fd_pr__nfet_01v8__k2_diff_30 = '4.81250e-07*lvn_bodyeffect*lvn_bodyeffect+2.15000e-06*lvn_bodyeffect+4.30650e-03'
+ sky130_fd_pr__nfet_01v8__k2_diff_31 = '2.71919e-04*lvn_bodyeffect*lvn_bodyeffect+-7.55225e-03*lvn_bodyeffect+-2.14770e-03'
+ sky130_fd_pr__nfet_01v8__k2_diff_32 = '6.77812e-05*lvn_bodyeffect*lvn_bodyeffect+-5.48500e-03*lvn_bodyeffect+7.18450e-03'
+ sky130_fd_pr__nfet_01v8__k2_diff_33 = '6.84375e-06*lvn_bodyeffect*lvn_bodyeffect+-2.44152e-03*lvn_bodyeffect+6.04440e-03'
+ sky130_fd_pr__nfet_01v8__k2_diff_34 = '-7.08437e-06*lvn_bodyeffect*lvn_bodyeffect+-1.52787e-04*lvn_bodyeffect+1.85090e-03'
+ sky130_fd_pr__nfet_01v8__k2_diff_35 = '1.95441e-05*lvn_bodyeffect*lvn_bodyeffect+-3.38149e-04*lvn_bodyeffect+1.71410e-03'
+ sky130_fd_pr__nfet_01v8__k2_diff_36 = '1.32156e-05*lvn_bodyeffect*lvn_bodyeffect+1.08181e-03*lvn_bodyeffect+5.11590e-03'
+ sky130_fd_pr__nfet_01v8__k2_diff_37 = '8.02500e-06*lvn_bodyeffect*lvn_bodyeffect+-1.86775e-04*lvn_bodyeffect+4.02200e-03'
+ sky130_fd_pr__nfet_01v8__k2_diff_38 = '1.29781e-05*lvn_bodyeffect*lvn_bodyeffect+-3.09963e-04*lvn_bodyeffect+8.42700e-03'
+ sky130_fd_pr__nfet_01v8__k2_diff_39 = '1.37837e-05*lvn_bodyeffect*lvn_bodyeffect+4.40600e-04*lvn_bodyeffect+-1.82840e-04'
+ sky130_fd_pr__nfet_01v8__k2_diff_4 = '2.96875e-07*lvn_bodyeffect*lvn_bodyeffect+6.65375e-05*lvn_bodyeffect+4.48600e-03'
+ sky130_fd_pr__nfet_01v8__k2_diff_40 = '1.65694e-04*lvn_bodyeffect*lvn_bodyeffect+-7.11450e-03*lvn_bodyeffect+1.97590e-03'
+ sky130_fd_pr__nfet_01v8__k2_diff_41 = '1.95556e-04*lvn_bodyeffect*lvn_bodyeffect+-4.06788e-03*lvn_bodyeffect+-3.36840e-03'
+ sky130_fd_pr__nfet_01v8__k2_diff_42 = '1.36094e-05*lvn_bodyeffect*lvn_bodyeffect+2.59312e-04*lvn_bodyeffect+1.02510e-02'
+ sky130_fd_pr__nfet_01v8__k2_diff_43 = '4.60375e-05*lvn_bodyeffect*lvn_bodyeffect+-1.13343e-03*lvn_bodyeffect+6.31570e-03'
+ sky130_fd_pr__nfet_01v8__k2_diff_44 = '-2.63750e-06*lvn_bodyeffect*lvn_bodyeffect+3.96975e-04*lvn_bodyeffect+5.59830e-03'
+ sky130_fd_pr__nfet_01v8__k2_diff_45 = '1.18781e-05*lvn_bodyeffect*lvn_bodyeffect+-5.47962e-04*lvn_bodyeffect+3.07880e-03'
+ sky130_fd_pr__nfet_01v8__k2_diff_46 = '8.15625e-06*lvn_bodyeffect*lvn_bodyeffect+4.51100e-04*lvn_bodyeffect+3.76140e-03'
+ sky130_fd_pr__nfet_01v8__k2_diff_47 = '2.36362e-04*lvn_bodyeffect*lvn_bodyeffect+-7.45412e-03*lvn_bodyeffect+1.50070e-03'
+ sky130_fd_pr__nfet_01v8__k2_diff_48 = '2.92844e-05*lvn_bodyeffect*lvn_bodyeffect+1.85812e-04*lvn_bodyeffect+2.27280e-03'
+ sky130_fd_pr__nfet_01v8__k2_diff_49 = '3.01706e-04*lvn_bodyeffect*lvn_bodyeffect+-7.72088e-03*lvn_bodyeffect+4.09920e-03'
+ sky130_fd_pr__nfet_01v8__k2_diff_5 = '1.08125e-06*lvn_bodyeffect*lvn_bodyeffect+2.45075e-04*lvn_bodyeffect+6.64350e-03'
+ sky130_fd_pr__nfet_01v8__k2_diff_50 = '2.98110e-04*lvn_bodyeffect*lvn_bodyeffect+-7.44412e-03*lvn_bodyeffect+7.61740e-04'
+ sky130_fd_pr__nfet_01v8__k2_diff_51 = '3.00294e-04*lvn_bodyeffect*lvn_bodyeffect+-7.55461e-03*lvn_bodyeffect'
+ sky130_fd_pr__nfet_01v8__k2_diff_52 = '1.21750e-05*lvn_bodyeffect*lvn_bodyeffect+-2.12830e-03*lvn_bodyeffect+1.16330e-02'
+ sky130_fd_pr__nfet_01v8__k2_diff_53 = '7.49312e-05*lvn_bodyeffect*lvn_bodyeffect+-3.00255e-03*lvn_bodyeffect+9.06490e-03'
+ sky130_fd_pr__nfet_01v8__k2_diff_54 = '2.15938e-04*lvn_bodyeffect*lvn_bodyeffect+-6.63250e-03*lvn_bodyeffect'
+ sky130_fd_pr__nfet_01v8__k2_diff_55 = '2.21906e-04*lvn_bodyeffect*lvn_bodyeffect+-6.90613e-03*lvn_bodyeffect'
+ sky130_fd_pr__nfet_01v8__k2_diff_56 = '2.50844e-04*lvn_bodyeffect*lvn_bodyeffect+-6.66188e-03*lvn_bodyeffect'
+ sky130_fd_pr__nfet_01v8__k2_diff_57 = '2.63563e-04*lvn_bodyeffect*lvn_bodyeffect+-6.56725e-03*lvn_bodyeffect'
+ sky130_fd_pr__nfet_01v8__k2_diff_58 = '2.72563e-04*lvn_bodyeffect*lvn_bodyeffect+-6.50475e-03*lvn_bodyeffect'
+ sky130_fd_pr__nfet_01v8__k2_diff_59 = '2.88500e-04*lvn_bodyeffect*lvn_bodyeffect+-6.32100e-03*lvn_bodyeffect'
+ sky130_fd_pr__nfet_01v8__k2_diff_6 = '3.11900e-04*lvn_bodyeffect*lvn_bodyeffect+-8.15963e-03*lvn_bodyeffect+1.04010e-03'
+ sky130_fd_pr__nfet_01v8__k2_diff_60 = '6.64688e-05*lvn_bodyeffect*lvn_bodyeffect+-2.87088e-03*lvn_bodyeffect'
+ sky130_fd_pr__nfet_01v8__k2_diff_61 = '-8.13750e-06*lvn_bodyeffect*lvn_bodyeffect+-1.49147e-03*lvn_bodyeffect'
+ sky130_fd_pr__nfet_01v8__k2_diff_62 = '3.66125e-05*lvn_bodyeffect*lvn_bodyeffect+7.42975e-04*lvn_bodyeffect'
+ sky130_fd_pr__nfet_01v8__k2_diff_7 = '6.06563e-05*lvn_bodyeffect*lvn_bodyeffect+-4.50700e-03*lvn_bodyeffect+2.66650e-03'
+ sky130_fd_pr__nfet_01v8__k2_diff_8 = '-8.96000e-06*lvn_bodyeffect*lvn_bodyeffect+-1.83821e-03*lvn_bodyeffect+3.31910e-04'
+ sky130_fd_pr__nfet_01v8__k2_diff_9 = '-3.37188e-06*lvn_bodyeffect*lvn_bodyeffect+-2.74862e-04*lvn_bodyeffect+4.85380e-03'
+ sky130_fd_pr__nfet_01v8__keta_diff_52 = '-4.89387e-05*lvn_bodyeffect*lvn_bodyeffect+-9.62142e-04*lvn_bodyeffect'
+ sky130_fd_pr__nfet_01v8__keta_diff_53 = '-1.55894e-05*lvn_bodyeffect*lvn_bodyeffect+-3.35558e-04*lvn_bodyeffect'
+ sky130_fd_pr__nfet_01v8__keta_diff_54 = '3.68250e-06*lvn_bodyeffect*lvn_bodyeffect+1.09023e-04*lvn_bodyeffect'
+ sky130_fd_pr__nfet_01v8__keta_diff_55 = '1.30031e-06*lvn_bodyeffect*lvn_bodyeffect+4.01063e-05*lvn_bodyeffect'
+ sky130_fd_pr__nfet_01v8__kt1_diff_51 = '-3.86647e-07*lvn_subvt*lvn_subvt+-1.67345e-05*lvn_subvt'
+ sky130_fd_pr__nfet_01v8__kt1_diff_56 = '3.40509e-07*lvn_subvt*lvn_subvt+1.13509e-05*lvn_subvt'
+ sky130_fd_pr__nfet_01v8__kt1_diff_57 = '3.38634e-07*lvn_subvt*lvn_subvt+1.17095e-05*lvn_subvt'
+ sky130_fd_pr__nfet_01v8__kt1_diff_58 = '2.88769e-07*lvn_subvt*lvn_subvt+1.01648e-05*lvn_subvt'
+ sky130_fd_pr__nfet_01v8__lint_diff = '-1.62422e-10*poly_cd*poly_cd+-3.68156e-09*poly_cd'
+ sky130_fd_pr__nfet_01v8__nfactor_diff_0 = '-2.45906e-03*lvn_subvt*lvn_subvt+-1.63649e-01*lvn_subvt+3.76680e-01'
+ sky130_fd_pr__nfet_01v8__nfactor_diff_1 = '-4.44781e-03*lvn_subvt*lvn_subvt+-1.98201e-01*lvn_subvt+3.19360e-01'
+ sky130_fd_pr__nfet_01v8__nfactor_diff_10 = '-2.57119e-03*lvn_subvt*lvn_subvt+-1.28687e-01*lvn_subvt+5.84990e-01'
+ sky130_fd_pr__nfet_01v8__nfactor_diff_11 = '-7.04687e-04*lvn_subvt*lvn_subvt+1.08712e-02*lvn_subvt+9.63200e-01'
+ sky130_fd_pr__nfet_01v8__nfactor_diff_12 = '1.40937e-04*lvn_subvt*lvn_subvt+-1.29613e-02*lvn_subvt+1.01730e+00'
+ sky130_fd_pr__nfet_01v8__nfactor_diff_13 = '-9.31250e-05*lvn_subvt*lvn_subvt+-1.22530e-01*lvn_subvt+9.81670e-01'
+ sky130_fd_pr__nfet_01v8__nfactor_diff_14 = '3.54688e-04*lvn_subvt*lvn_subvt+-6.97438e-02*lvn_subvt+9.14250e-01'
+ sky130_fd_pr__nfet_01v8__nfactor_diff_15 = '-1.24063e-04*lvn_subvt*lvn_subvt+-4.28463e-02*lvn_subvt+1.02340e+00'
+ sky130_fd_pr__nfet_01v8__nfactor_diff_16 = '5.62187e-04*lvn_subvt*lvn_subvt+2.32337e-02*lvn_subvt+6.32660e-01'
+ sky130_fd_pr__nfet_01v8__nfactor_diff_17 = '3.15625e-04*lvn_subvt*lvn_subvt+2.84375e-02*lvn_subvt+1.35870e+00'
+ sky130_fd_pr__nfet_01v8__nfactor_diff_18 = '-1.99375e-04*lvn_subvt*lvn_subvt+1.16325e-02*lvn_subvt+9.86560e-01'
+ sky130_fd_pr__nfet_01v8__nfactor_diff_19 = '-1.42500e-04*lvn_subvt*lvn_subvt+1.25625e-02*lvn_subvt+9.15550e-01'
+ sky130_fd_pr__nfet_01v8__nfactor_diff_2 = '-1.02375e-03*lvn_subvt*lvn_subvt+-3.21200e-02*lvn_subvt+1.11000e+00'
+ sky130_fd_pr__nfet_01v8__nfactor_diff_20 = '1.53437e-04*lvn_subvt*lvn_subvt+-7.10125e-03*lvn_subvt+9.87040e-01'
+ sky130_fd_pr__nfet_01v8__nfactor_diff_21 = '-1.69063e-04*lvn_subvt*lvn_subvt+1.31213e-02*lvn_subvt+8.74210e-01'
+ sky130_fd_pr__nfet_01v8__nfactor_diff_22 = '4.17500e-04*lvn_subvt*lvn_subvt+-6.35875e-02*lvn_subvt+9.12570e-01'
+ sky130_fd_pr__nfet_01v8__nfactor_diff_23 = '-1.10937e-03*lvn_subvt*lvn_subvt+-5.84625e-02*lvn_subvt+1.37570e+00'
+ sky130_fd_pr__nfet_01v8__nfactor_diff_24 = '4.12500e-04*lvn_subvt*lvn_subvt+9.70000e-03*lvn_subvt+1.60870e+00'
+ sky130_fd_pr__nfet_01v8__nfactor_diff_25 = '5.66562e-04*lvn_subvt*lvn_subvt+5.15838e-02*lvn_subvt+1.19140e+00'
+ sky130_fd_pr__nfet_01v8__nfactor_diff_26 = '-3.75000e-05*lvn_subvt*lvn_subvt+6.30000e-03*lvn_subvt+1.13970e+00'
+ sky130_fd_pr__nfet_01v8__nfactor_diff_27 = '-1.56562e-04*lvn_subvt*lvn_subvt+4.14375e-03*lvn_subvt+9.76110e-01'
+ sky130_fd_pr__nfet_01v8__nfactor_diff_28 = '-4.40625e-05*lvn_subvt*lvn_subvt+3.97125e-03*lvn_subvt+9.55690e-01'
+ sky130_fd_pr__nfet_01v8__nfactor_diff_29 = '-6.21875e-05*lvn_subvt*lvn_subvt+7.81125e-03*lvn_subvt+8.74530e-01'
+ sky130_fd_pr__nfet_01v8__nfactor_diff_3 = '-4.42500e-04*lvn_subvt*lvn_subvt+-2.55175e-02*lvn_subvt+8.12720e-01'
+ sky130_fd_pr__nfet_01v8__nfactor_diff_30 = '-1.15312e-04*lvn_subvt*lvn_subvt+1.32663e-02*lvn_subvt+8.33310e-01'
+ sky130_fd_pr__nfet_01v8__nfactor_diff_31 = '3.47578e-03*lvn_subvt*lvn_subvt+-1.07061e-01*lvn_subvt+-5.42090e-01'
+ sky130_fd_pr__nfet_01v8__nfactor_diff_32 = '3.78125e-04*lvn_subvt*lvn_subvt+1.43375e-02*lvn_subvt+1.51010e+00'
+ sky130_fd_pr__nfet_01v8__nfactor_diff_33 = '4.65312e-04*lvn_subvt*lvn_subvt+8.35387e-02*lvn_subvt+1.01770e+00'
+ sky130_fd_pr__nfet_01v8__nfactor_diff_34 = '-1.37500e-04*lvn_subvt*lvn_subvt+1.32000e-02*lvn_subvt+1.08620e+00'
+ sky130_fd_pr__nfet_01v8__nfactor_diff_35 = '2.37500e-04*lvn_subvt*lvn_subvt+-1.86450e-01*lvn_subvt+1.76540e+00'
+ sky130_fd_pr__nfet_01v8__nfactor_diff_36 = '3.75625e-04*lvn_subvt*lvn_subvt+1.42722e-01*lvn_subvt+1.54530e+00'
+ sky130_fd_pr__nfet_01v8__nfactor_diff_37 = '2.91250e-03*lvn_subvt*lvn_subvt+-9.84000e-02*lvn_subvt+1.42710e+00'
+ sky130_fd_pr__nfet_01v8__nfactor_diff_38 = '2.17813e-03*lvn_subvt*lvn_subvt+-4.01375e-02*lvn_subvt+1.21190e+00'
+ sky130_fd_pr__nfet_01v8__nfactor_diff_39 = '8.00000e-04*lvn_subvt*lvn_subvt+9.06000e-02*lvn_subvt+1.29570e+00'
+ sky130_fd_pr__nfet_01v8__nfactor_diff_4 = '3.40625e-04*lvn_subvt*lvn_subvt+4.51250e-03*lvn_subvt+1.09140e+00'
+ sky130_fd_pr__nfet_01v8__nfactor_diff_40 = '8.06094e-03*lvn_subvt*lvn_subvt+-1.03019e-01*lvn_subvt+7.29050e-01'
+ sky130_fd_pr__nfet_01v8__nfactor_diff_41 = '-3.72563e-03*lvn_subvt*lvn_subvt+-1.41125e-01*lvn_subvt+1.92300e-01'
+ sky130_fd_pr__nfet_01v8__nfactor_diff_42 = '-5.79469e-02*lvn_subvt*lvn_subvt+-2.21912e-01*lvn_subvt+1.76350e+00'
+ sky130_fd_pr__nfet_01v8__nfactor_diff_43 = '-3.28875e-03*lvn_subvt*lvn_subvt+-1.51980e-01*lvn_subvt+1.48220e+00'
+ sky130_fd_pr__nfet_01v8__nfactor_diff_44 = '1.89375e-03*lvn_subvt*lvn_subvt+-1.44750e-02*lvn_subvt+1.44430e+00'
+ sky130_fd_pr__nfet_01v8__nfactor_diff_45 = '9.57500e-04*lvn_subvt*lvn_subvt+-8.96700e-02*lvn_subvt+1.11600e+00'
+ sky130_fd_pr__nfet_01v8__nfactor_diff_46 = '-1.97812e-04*lvn_subvt*lvn_subvt+1.02516e-01*lvn_subvt+1.06300e+00'
+ sky130_fd_pr__nfet_01v8__nfactor_diff_47 = '5.59281e-03*lvn_subvt*lvn_subvt+-9.91587e-02*lvn_subvt+6.35380e-01'
+ sky130_fd_pr__nfet_01v8__nfactor_diff_48 = '-4.40312e-03*lvn_subvt*lvn_subvt+-2.55375e-02*lvn_subvt+1.65690e+00'
+ sky130_fd_pr__nfet_01v8__nfactor_diff_49 = '-3.15312e-03*lvn_subvt*lvn_subvt+-1.30705e-01*lvn_subvt+4.69740e-01'
+ sky130_fd_pr__nfet_01v8__nfactor_diff_5 = '-5.63437e-04*lvn_subvt*lvn_subvt+7.01037e-02*lvn_subvt+1.12050e+00'
+ sky130_fd_pr__nfet_01v8__nfactor_diff_50 = '1.18344e-04*lvn_subvt*lvn_subvt+-6.29541e-02*lvn_subvt+3.17290e-01'
+ sky130_fd_pr__nfet_01v8__nfactor_diff_51 = '-1.17296e-03*lvn_subvt*lvn_subvt+-9.20900e-02*lvn_subvt'
+ sky130_fd_pr__nfet_01v8__nfactor_diff_52 = '9.62568e-03*lvn_subvt*lvn_subvt+-1.09887e-01*lvn_subvt'
+ sky130_fd_pr__nfet_01v8__nfactor_diff_53 = '8.80955e-03*lvn_subvt*lvn_subvt+-1.05720e-01*lvn_subvt'
+ sky130_fd_pr__nfet_01v8__nfactor_diff_54 = '6.06442e-03*lvn_subvt*lvn_subvt+-9.94092e-02*lvn_subvt'
+ sky130_fd_pr__nfet_01v8__nfactor_diff_55 = '5.74449e-03*lvn_subvt*lvn_subvt+-9.92172e-02*lvn_subvt'
+ sky130_fd_pr__nfet_01v8__nfactor_diff_56 = '2.30512e-03*lvn_subvt*lvn_subvt+-1.11215e-01*lvn_subvt'
+ sky130_fd_pr__nfet_01v8__nfactor_diff_57 = '3.37291e-04*lvn_subvt*lvn_subvt+-1.18320e-01*lvn_subvt'
+ sky130_fd_pr__nfet_01v8__nfactor_diff_58 = '-5.87593e-04*lvn_subvt*lvn_subvt+-1.21629e-01*lvn_subvt'
+ sky130_fd_pr__nfet_01v8__nfactor_diff_59 = '-2.91092e-03*lvn_subvt*lvn_subvt+-1.26286e-01*lvn_subvt'
+ sky130_fd_pr__nfet_01v8__nfactor_diff_6 = '-5.87278e-03*lvn_subvt*lvn_subvt+-1.83076e-01*lvn_subvt+8.53660e-01'
+ sky130_fd_pr__nfet_01v8__nfactor_diff_60 = '-2.91092e-03*lvn_subvt*lvn_subvt+-1.26286e-01*lvn_subvt'
+ sky130_fd_pr__nfet_01v8__nfactor_diff_61 = '-1.10881e-02*lvn_subvt*lvn_subvt+-1.60178e-01*lvn_subvt'
+ sky130_fd_pr__nfet_01v8__nfactor_diff_62 = '-4.40312e-03*lvn_subvt*lvn_subvt+-2.55375e-02*lvn_subvt'
+ sky130_fd_pr__nfet_01v8__nfactor_diff_7 = '1.82700e-03*lvn_subvt*lvn_subvt+-1.88567e-01*lvn_subvt+6.39180e-02'
+ sky130_fd_pr__nfet_01v8__nfactor_diff_8 = '-1.10881e-02*lvn_subvt*lvn_subvt+-1.60178e-01*lvn_subvt+1.10530e+00'
+ sky130_fd_pr__nfet_01v8__nfactor_diff_9 = '-1.59375e-04*lvn_subvt*lvn_subvt+-3.71125e-02*lvn_subvt+1.41730e+00'
+ sky130_fd_pr__nfet_01v8__overlap_mult = '-6.32500e-04*lvtox*lvtox+1.48000e-03*lvtox+9.64200e-01'
+ sky130_fd_pr__nfet_01v8__pclm_diff_51 = '-2.12219e-06*lvn_saturation*lvn_saturation+-9.18562e-05*lvn_saturation'
+ sky130_fd_pr__nfet_01v8__pclm_diff_52 = '-1.46666e-05*lvn_saturation*lvn_saturation+-2.88349e-04*lvn_saturation'
+ sky130_fd_pr__nfet_01v8__pclm_diff_53 = '-4.67188e-06*lvn_saturation*lvn_saturation+-1.00565e-04*lvn_saturation'
+ sky130_fd_pr__nfet_01v8__pclm_diff_54 = '1.10344e-06*lvn_saturation*lvn_saturation+3.26738e-05*lvn_saturation'
+ sky130_fd_pr__nfet_01v8__pclm_diff_55 = '3.89634e-07*lvn_saturation*lvn_saturation+1.20196e-05*lvn_saturation'
+ sky130_fd_pr__nfet_01v8__pclm_diff_56 = '6.67394e-07*lvn_saturation*lvn_saturation+2.22478e-05*lvn_saturation'
+ sky130_fd_pr__nfet_01v8__pclm_diff_57 = '6.63669e-07*lvn_saturation*lvn_saturation+2.29503e-05*lvn_saturation'
+ sky130_fd_pr__nfet_01v8__pclm_diff_58 = '5.65991e-07*lvn_saturation*lvn_saturation+1.99230e-05*lvn_saturation'
+ sky130_fd_pr__nfet_01v8__pclm_diff_59 = '-6.12516e-07*lvn_saturation*lvn_saturation+-2.30824e-05*lvn_saturation'
+ sky130_fd_pr__nfet_01v8__pclm_diff_60 = '-6.12528e-07*lvn_saturation*lvn_saturation+-2.30824e-05*lvn_saturation'
+ sky130_fd_pr__nfet_01v8__pjunction_mult = '-1.25000e-06*lvn_diode*lvn_diode+5.67550e-02*lvn_diode+1.02040e+00'
+ sky130_fd_pr__rf_nfet_01v8_b__ajunction_mult = '-1.87500e-06*lvn_diode*lvn_diode+5.53750e-02*lvn_diode+9.95430e-01'
+ sky130_fd_pr__rf_nfet_01v8_b__dlc_diff = '-1.06849e-10*poly_cd*poly_cd+-3.77438e-09*poly_cd+-6.14920e-10'
+ sky130_fd_pr__rf_nfet_01v8_b__lint_diff = '-4.33125e-09*poly_cd'
+ sky130_fd_pr__rf_nfet_01v8_b__overlap_mult = '-6.32500e-04*lvtox*lvtox+1.48000e-03*lvtox+9.64200e-01'
+ sky130_fd_pr__rf_nfet_01v8_b__pjunction_mult = '-1.25000e-06*lvn_diode*lvn_diode+5.67550e-02*lvn_diode+1.02040e+00'
+ sky130_fd_pr__rf_nfet_01v8_b__rbpb_mult = '5.00000e-02*lvn_bodyeffect+1.00000e+00'
+ sky130_fd_pr__rf_nfet_01v8_b__rshg_diff = '1.75000e+00*ic_res'
+ sky130_fd_pr__rf_nfet_01v8_b__toxe_mult = '1.30000e-02*lvtox+1.00000e+00'
+ sky130_fd_pr__rf_nfet_01v8_b__wint_diff = '8.04375e-09*diff_cd'
+ sky130_fd_pr__rf_nfet_01v8_b__xgw_diff = '1.60625e-08*diff_cd'
+ sky130_fd_pr__rf_nfet_01v8_bM02__k2_diff_0 = '9.86813e-05*lvn_bodyeffect*lvn_bodyeffect+-2.16475e-04*lvn_bodyeffect+7.64020e-03'
+ sky130_fd_pr__rf_nfet_01v8_bM02__k2_diff_1 = '3.98437e-05*lvn_bodyeffect*lvn_bodyeffect+-8.01375e-04*lvn_bodyeffect+1.68400e-02'
+ sky130_fd_pr__rf_nfet_01v8_bM02__k2_diff_2 = '2.04688e-05*lvn_bodyeffect*lvn_bodyeffect+-7.86125e-04*lvn_bodyeffect+3.45610e-02'
+ sky130_fd_pr__rf_nfet_01v8_bM02__k2_diff_3 = '1.15172e-04*lvn_bodyeffect*lvn_bodyeffect+-1.04921e-03*lvn_bodyeffect+4.58640e-03'
+ sky130_fd_pr__rf_nfet_01v8_bM02__k2_diff_4 = '8.01562e-05*lvn_bodyeffect*lvn_bodyeffect+-2.15937e-03*lvn_bodyeffect+2.04550e-02'
+ sky130_fd_pr__rf_nfet_01v8_bM02__k2_diff_5 = '3.81250e-05*lvn_bodyeffect*lvn_bodyeffect+-1.28100e-03*lvn_bodyeffect+3.72450e-02'
+ sky130_fd_pr__rf_nfet_01v8_bM02__k2_diff_6 = '1.12641e-04*lvn_bodyeffect*lvn_bodyeffect+-6.86062e-04*lvn_bodyeffect+1.94870e-03'
+ sky130_fd_pr__rf_nfet_01v8_bM02__k2_diff_7 = '7.50000e-05*lvn_bodyeffect*lvn_bodyeffect+-1.86975e-03*lvn_bodyeffect+1.77710e-02'
+ sky130_fd_pr__rf_nfet_01v8_bM02__k2_diff_8 = '3.85937e-05*lvn_bodyeffect*lvn_bodyeffect+-1.41812e-03*lvn_bodyeffect+3.54600e-02'
+ sky130_fd_pr__rf_nfet_01v8_bM02__u0_diff_0 = '-2.03169e-05*lvn_mobility*lvn_mobility+-7.14350e-05*lvn_mobility+7.86820e-04'
+ sky130_fd_pr__rf_nfet_01v8_bM02__u0_diff_1 = '-2.40125e-05*lvn_mobility*lvn_mobility+-2.04582e-04*lvn_mobility+6.95070e-04'
+ sky130_fd_pr__rf_nfet_01v8_bM02__u0_diff_2 = '-2.55544e-05*lvn_mobility*lvn_mobility+-3.10587e-04*lvn_mobility+-1.86680e-04'
+ sky130_fd_pr__rf_nfet_01v8_bM02__u0_diff_3 = '-1.55000e-05*lvn_mobility*lvn_mobility+-4.14350e-04*lvn_mobility+-5.08880e-03'
+ sky130_fd_pr__rf_nfet_01v8_bM02__u0_diff_4 = '-2.01469e-05*lvn_mobility*lvn_mobility+-9.54875e-05*lvn_mobility+-3.38250e-03'
+ sky130_fd_pr__rf_nfet_01v8_bM02__u0_diff_5 = '-2.12863e-05*lvn_mobility*lvn_mobility+-3.87613e-04*lvn_mobility+-1.08370e-04'
+ sky130_fd_pr__rf_nfet_01v8_bM02__u0_diff_6 = '-1.66125e-05*lvn_mobility*lvn_mobility+-1.83325e-04*lvn_mobility+-3.81310e-03'
+ sky130_fd_pr__rf_nfet_01v8_bM02__u0_diff_7 = '-1.86562e-05*lvn_mobility*lvn_mobility+-7.10500e-05*lvn_mobility+-3.65260e-03'
+ sky130_fd_pr__rf_nfet_01v8_bM02__u0_diff_8 = '-2.01562e-05*lvn_mobility*lvn_mobility+-3.97775e-04*lvn_mobility+-2.32590e-03'
+ sky130_fd_pr__rf_nfet_01v8_bM02__vsat_diff_0 = '-1.15489e+02*lvn_saturation*lvn_saturation+5.36138e+03*lvn_saturation+8.76330e+02'
+ sky130_fd_pr__rf_nfet_01v8_bM02__vsat_diff_1 = '4.23912e+01*lvn_saturation*lvn_saturation+5.05100e+03*lvn_saturation+2.92740e+02'
+ sky130_fd_pr__rf_nfet_01v8_bM02__vsat_diff_2 = '2.37344e+02*lvn_saturation*lvn_saturation+6.14662e+03*lvn_saturation+4.00800e+03'
+ sky130_fd_pr__rf_nfet_01v8_bM02__vsat_diff_3 = '-1.44812e+01*lvn_saturation*lvn_saturation+5.13850e+03*lvn_saturation+-7.67730e+03'
+ sky130_fd_pr__rf_nfet_01v8_bM02__vsat_diff_4 = '1.45662e+02*lvn_saturation*lvn_saturation+6.06888e+03*lvn_saturation+-3.22610e+03'
+ sky130_fd_pr__rf_nfet_01v8_bM02__vsat_diff_5 = '2.18925e+02*lvn_saturation*lvn_saturation+5.16400e+03*lvn_saturation+-3.10380e+03'
+ sky130_fd_pr__rf_nfet_01v8_bM02__vsat_diff_6 = '-1.10087e+02*lvn_saturation*lvn_saturation+4.09440e+03*lvn_saturation+-1.05210e+04'
+ sky130_fd_pr__rf_nfet_01v8_bM02__vsat_diff_7 = '1.07662e+02*lvn_saturation*lvn_saturation+5.22625e+03*lvn_saturation+-3.85660e+03'
+ sky130_fd_pr__rf_nfet_01v8_bM02__vsat_diff_8 = '1.96437e+02*lvn_saturation*lvn_saturation+4.60912e+03*lvn_saturation+-7.49490e+02'
+ sky130_fd_pr__rf_nfet_01v8_bM02__vth0_diff_0 = '-1.62094e-04*lvn_threshold*lvn_threshold+1.35881e-02*lvn_threshold+-1.90450e-02'
+ sky130_fd_pr__rf_nfet_01v8_bM02__vth0_diff_1 = '-7.34188e-05*lvn_threshold*lvn_threshold+8.96013e-03*lvn_threshold+-2.47180e-03'
+ sky130_fd_pr__rf_nfet_01v8_bM02__vth0_diff_2 = '-4.36562e-05*lvn_threshold*lvn_threshold+7.71487e-03*lvn_threshold+-1.14640e-02'
+ sky130_fd_pr__rf_nfet_01v8_bM02__vth0_diff_3 = '-1.64381e-04*lvn_threshold*lvn_threshold+8.90112e-03*lvn_threshold+3.12960e-03'
+ sky130_fd_pr__rf_nfet_01v8_bM02__vth0_diff_4 = '-1.15569e-04*lvn_threshold*lvn_threshold+7.71322e-03*lvn_threshold+-1.91180e-02'
+ sky130_fd_pr__rf_nfet_01v8_bM02__vth0_diff_5 = '-5.94469e-05*lvn_threshold*lvn_threshold+5.11071e-03*lvn_threshold+-1.09280e-02'
+ sky130_fd_pr__rf_nfet_01v8_bM02__vth0_diff_6 = '-1.75688e-04*lvn_threshold*lvn_threshold+7.06775e-03*lvn_threshold+-1.03570e-02'
+ sky130_fd_pr__rf_nfet_01v8_bM02__vth0_diff_7 = '-1.04675e-04*lvn_threshold*lvn_threshold+6.36330e-03*lvn_threshold+-1.86330e-02'
+ sky130_fd_pr__rf_nfet_01v8_bM02__vth0_diff_8 = '-5.97938e-05*lvn_threshold*lvn_threshold+4.31957e-03*lvn_threshold+-1.47380e-02'
+ sky130_fd_pr__rf_nfet_01v8_bM04__k2_diff_0 = '1.01206e-04*lvn_bodyeffect*lvn_bodyeffect+-2.39325e-04*lvn_bodyeffect+6.60760e-03'
+ sky130_fd_pr__rf_nfet_01v8_bM04__k2_diff_1 = '7.19375e-05*lvn_bodyeffect*lvn_bodyeffect+-1.34700e-03*lvn_bodyeffect+2.24380e-02'
+ sky130_fd_pr__rf_nfet_01v8_bM04__k2_diff_2 = '3.36875e-05*lvn_bodyeffect*lvn_bodyeffect+-1.03250e-03*lvn_bodyeffect+3.75000e-02'
+ sky130_fd_pr__rf_nfet_01v8_bM04__k2_diff_3 = '1.50000e-04*lvn_bodyeffect*lvn_bodyeffect+-1.47690e-03*lvn_bodyeffect+5.54840e-03'
+ sky130_fd_pr__rf_nfet_01v8_bM04__k2_diff_4 = '9.85312e-05*lvn_bodyeffect*lvn_bodyeffect+-2.44437e-03*lvn_bodyeffect+2.36230e-02'
+ sky130_fd_pr__rf_nfet_01v8_bM04__k2_diff_5 = '4.27812e-05*lvn_bodyeffect*lvn_bodyeffect+-1.40612e-03*lvn_bodyeffect+3.90920e-02'
+ sky130_fd_pr__rf_nfet_01v8_bM04__k2_diff_6 = '1.46059e-04*lvn_bodyeffect*lvn_bodyeffect+-1.06724e-03*lvn_bodyeffect+2.99510e-03'
+ sky130_fd_pr__rf_nfet_01v8_bM04__k2_diff_7 = '9.85000e-05*lvn_bodyeffect*lvn_bodyeffect+-2.19400e-03*lvn_bodyeffect+2.15790e-02'
+ sky130_fd_pr__rf_nfet_01v8_bM04__k2_diff_8 = '4.26875e-05*lvn_bodyeffect*lvn_bodyeffect+-1.52550e-03*lvn_bodyeffect+3.73290e-02'
+ sky130_fd_pr__rf_nfet_01v8_bM04__u0_diff_0 = '-2.36125e-05*lvn_mobility*lvn_mobility+-9.13050e-05*lvn_mobility+-6.96680e-04'
+ sky130_fd_pr__rf_nfet_01v8_bM04__u0_diff_1 = '-2.69156e-05*lvn_mobility*lvn_mobility+-1.03337e-04*lvn_mobility+-1.34750e-03'
+ sky130_fd_pr__rf_nfet_01v8_bM04__u0_diff_2 = '-2.58159e-05*lvn_mobility*lvn_mobility+-2.66011e-04*lvn_mobility+-1.00130e-03'
+ sky130_fd_pr__rf_nfet_01v8_bM04__u0_diff_3 = '-1.96437e-05*lvn_mobility*lvn_mobility+-3.09800e-04*lvn_mobility+-5.73800e-03'
+ sky130_fd_pr__rf_nfet_01v8_bM04__u0_diff_4 = '-2.20062e-05*lvn_mobility*lvn_mobility+1.62250e-05*lvn_mobility+-6.72530e-03'
+ sky130_fd_pr__rf_nfet_01v8_bM04__u0_diff_5 = '-2.11250e-05*lvn_mobility*lvn_mobility+-2.42950e-04*lvn_mobility+-4.97740e-03'
+ sky130_fd_pr__rf_nfet_01v8_bM04__u0_diff_6 = '-1.91562e-05*lvn_mobility*lvn_mobility+-1.70875e-04*lvn_mobility+-3.71750e-03'
+ sky130_fd_pr__rf_nfet_01v8_bM04__u0_diff_7 = '-2.06969e-05*lvn_mobility*lvn_mobility+4.18625e-05*lvn_mobility+-5.53610e-03'
+ sky130_fd_pr__rf_nfet_01v8_bM04__u0_diff_8 = '-2.02562e-05*lvn_mobility*lvn_mobility+-3.29650e-04*lvn_mobility+-4.09270e-03'
+ sky130_fd_pr__rf_nfet_01v8_bM04__vsat_diff_0 = '-6.86938e+01*lvn_saturation*lvn_saturation+5.32662e+03*lvn_saturation+-9.57840e+03'
+ sky130_fd_pr__rf_nfet_01v8_bM04__vsat_diff_1 = '1.42819e+02*lvn_saturation*lvn_saturation+5.97550e+03*lvn_saturation+-1.94710e+03'
+ sky130_fd_pr__rf_nfet_01v8_bM04__vsat_diff_2 = '4.07231e+02*lvn_saturation*lvn_saturation+7.37000e+03*lvn_saturation+3.93430e+03'
+ sky130_fd_pr__rf_nfet_01v8_bM04__vsat_diff_3 = '-1.55125e+01*lvn_saturation*lvn_saturation+5.34838e+03*lvn_saturation+-9.28630e+03'
+ sky130_fd_pr__rf_nfet_01v8_bM04__vsat_diff_4 = '2.14356e+02*lvn_saturation*lvn_saturation+6.49375e+03*lvn_saturation+-2.37570e+03'
+ sky130_fd_pr__rf_nfet_01v8_bM04__vsat_diff_5 = '5.62681e+02*lvn_saturation*lvn_saturation+7.95552e+03*lvn_saturation+1.42910e+04'
+ sky130_fd_pr__rf_nfet_01v8_bM04__vsat_diff_6 = '-1.00753e+02*lvn_saturation*lvn_saturation+4.25624e+03*lvn_saturation+-1.13210e+04'
+ sky130_fd_pr__rf_nfet_01v8_bM04__vsat_diff_7 = '7.49312e+01*lvn_saturation*lvn_saturation+4.89662e+03*lvn_saturation+-8.60840e+03'
+ sky130_fd_pr__rf_nfet_01v8_bM04__vsat_diff_8 = '5.51006e+02*lvn_saturation*lvn_saturation+7.46000e+03*lvn_saturation+9.12790e+03'
+ sky130_fd_pr__rf_nfet_01v8_bM04__vth0_diff_0 = '-1.63794e-04*lvn_threshold*lvn_threshold+1.35991e-02*lvn_threshold+5.51620e-03'
+ sky130_fd_pr__rf_nfet_01v8_bM04__vth0_diff_1 = '-1.14875e-04*lvn_threshold*lvn_threshold+9.79050e-03*lvn_threshold+-1.71250e-02'
+ sky130_fd_pr__rf_nfet_01v8_bM04__vth0_diff_2 = '-6.13437e-05*lvn_threshold*lvn_threshold+8.03163e-03*lvn_threshold+-1.35250e-02'
+ sky130_fd_pr__rf_nfet_01v8_bM04__vth0_diff_3 = '-2.02750e-04*lvn_threshold*lvn_threshold+9.64162e-03*lvn_threshold+-5.00650e-03'
+ sky130_fd_pr__rf_nfet_01v8_bM04__vth0_diff_4 = '-1.44725e-04*lvn_threshold*lvn_threshold+8.33085e-03*lvn_threshold+-2.55090e-02'
+ sky130_fd_pr__rf_nfet_01v8_bM04__vth0_diff_5 = '-6.63719e-05*lvn_threshold*lvn_threshold+5.42226e-03*lvn_threshold+-1.84290e-02'
+ sky130_fd_pr__rf_nfet_01v8_bM04__vth0_diff_6 = '-2.01062e-04*lvn_threshold*lvn_threshold+7.62525e-03*lvn_threshold+-1.13020e-02'
+ sky130_fd_pr__rf_nfet_01v8_bM04__vth0_diff_7 = '-1.45200e-04*lvn_threshold*lvn_threshold+7.05445e-03*lvn_threshold+-2.98950e-02'
+ sky130_fd_pr__rf_nfet_01v8_bM04__vth0_diff_8 = '-6.84031e-05*lvn_threshold*lvn_threshold+4.64789e-03*lvn_threshold+-1.92140e-02'
+ sky130_fd_pr__nfet_01v8__toxe_mult = '1.30000e-02*lvtox+1.00000e+00'
+ sky130_fd_pr__nfet_01v8__u0_diff_0 = '1.58094e-06*lvn_mobility*lvn_mobility+6.34224e-04*lvn_mobility+-3.48940e-03'
+ sky130_fd_pr__nfet_01v8__u0_diff_1 = '-1.75356e-05*lvn_mobility*lvn_mobility+5.36507e-04*lvn_mobility+-2.69800e-03'
+ sky130_fd_pr__nfet_01v8__u0_diff_10 = '-5.42531e-06*lvn_mobility*lvn_mobility+6.60349e-04*lvn_mobility+-1.78280e-03'
+ sky130_fd_pr__nfet_01v8__u0_diff_11 = '-9.25413e-06*lvn_mobility*lvn_mobility+-9.35910e-05*lvn_mobility+-3.07710e-04'
+ sky130_fd_pr__nfet_01v8__u0_diff_12 = '-9.53750e-06*lvn_mobility*lvn_mobility+-1.23000e-04*lvn_mobility+-3.16130e-03'
+ sky130_fd_pr__nfet_01v8__u0_diff_13 = '-1.51469e-05*lvn_mobility*lvn_mobility+1.62563e-04*lvn_mobility+-3.17090e-03'
+ sky130_fd_pr__nfet_01v8__u0_diff_14 = '-9.50000e-06*lvn_mobility*lvn_mobility+8.99000e-05*lvn_mobility+-2.42050e-03'
+ sky130_fd_pr__nfet_01v8__u0_diff_15 = '5.20375e-06*lvn_mobility*lvn_mobility+8.82115e-04*lvn_mobility+-3.87010e-03'
+ sky130_fd_pr__nfet_01v8__u0_diff_16 = '-1.43656e-05*lvn_mobility*lvn_mobility+2.35788e-04*lvn_mobility+-1.96160e-03'
+ sky130_fd_pr__nfet_01v8__u0_diff_17 = '-2.14863e-05*lvn_mobility*lvn_mobility+-3.03005e-04*lvn_mobility+-1.34480e-03'
+ sky130_fd_pr__nfet_01v8__u0_diff_18 = '-2.58437e-06*lvn_mobility*lvn_mobility+6.68875e-05*lvn_mobility+-1.05560e-03'
+ sky130_fd_pr__nfet_01v8__u0_diff_19 = '-5.64406e-06*lvn_mobility*lvn_mobility+1.04125e-06*lvn_mobility+-3.54510e-04'
+ sky130_fd_pr__nfet_01v8__u0_diff_2 = '-2.55651e-05*lvn_mobility*lvn_mobility+-3.54116e-04*lvn_mobility+-9.22930e-05'
+ sky130_fd_pr__nfet_01v8__u0_diff_20 = '-7.00937e-06*lvn_mobility*lvn_mobility+-8.97875e-05*lvn_mobility+-4.28810e-03'
+ sky130_fd_pr__nfet_01v8__u0_diff_21 = '-8.37500e-06*lvn_mobility*lvn_mobility+-8.75250e-05*lvn_mobility+-2.87590e-03'
+ sky130_fd_pr__nfet_01v8__u0_diff_22 = '-8.98438e-06*lvn_mobility*lvn_mobility+7.16625e-05*lvn_mobility+-1.69540e-03'
+ sky130_fd_pr__nfet_01v8__u0_diff_23 = '1.41739e-05*lvn_mobility*lvn_mobility+6.90413e-04*lvn_mobility+3.96780e-06'
+ sky130_fd_pr__nfet_01v8__u0_diff_24 = '1.43281e-05*lvn_mobility*lvn_mobility+6.82738e-04*lvn_mobility+-7.32880e-03'
+ sky130_fd_pr__nfet_01v8__u0_diff_25 = '-1.65922e-05*lvn_mobility*lvn_mobility+-2.46006e-04*lvn_mobility+-1.07820e-03'
+ sky130_fd_pr__nfet_01v8__u0_diff_26 = '1.39062e-06*lvn_mobility*lvn_mobility+1.75765e-04*lvn_mobility+-3.54490e-04'
+ sky130_fd_pr__nfet_01v8__u0_diff_27 = '-4.52500e-06*lvn_mobility*lvn_mobility+-1.25000e-07*lvn_mobility+-1.49210e-03'
+ sky130_fd_pr__nfet_01v8__u0_diff_28 = '-7.25000e-06*lvn_mobility*lvn_mobility+-8.80750e-05*lvn_mobility+-1.76470e-03'
+ sky130_fd_pr__nfet_01v8__u0_diff_29 = '-9.00938e-06*lvn_mobility*lvn_mobility+-1.14887e-04*lvn_mobility+-1.45690e-03'
+ sky130_fd_pr__nfet_01v8__u0_diff_3 = '-2.27147e-05*lvn_mobility*lvn_mobility+-2.37156e-04*lvn_mobility+-4.33940e-04'
+ sky130_fd_pr__nfet_01v8__u0_diff_30 = '-8.44375e-06*lvn_mobility*lvn_mobility+-6.60500e-05*lvn_mobility+-1.21260e-03'
+ sky130_fd_pr__nfet_01v8__u0_diff_31 = '2.42316e-05*lvn_mobility*lvn_mobility+5.29099e-04*lvn_mobility+2.04660e-03'
+ sky130_fd_pr__nfet_01v8__u0_diff_32 = '8.95937e-06*lvn_mobility*lvn_mobility+6.43862e-04*lvn_mobility+-5.79780e-03'
+ sky130_fd_pr__nfet_01v8__u0_diff_33 = '-1.52313e-05*lvn_mobility*lvn_mobility+-2.55550e-04*lvn_mobility+-1.24650e-03'
+ sky130_fd_pr__nfet_01v8__u0_diff_34 = '1.86719e-06*lvn_mobility*lvn_mobility+1.72144e-04*lvn_mobility+-3.72100e-04'
+ sky130_fd_pr__nfet_01v8__u0_diff_35 = '-7.57813e-05*lvn_mobility*lvn_mobility+-6.24100e-04*lvn_mobility+-5.11790e-03'
+ sky130_fd_pr__nfet_01v8__u0_diff_36 = '-3.09031e-05*lvn_mobility*lvn_mobility+-4.65837e-04*lvn_mobility+-3.60190e-03'
+ sky130_fd_pr__nfet_01v8__u0_diff_37 = '-5.99438e-05*lvn_mobility*lvn_mobility+-4.96325e-04*lvn_mobility+-6.13530e-03'
+ sky130_fd_pr__nfet_01v8__u0_diff_38 = '-3.79875e-05*lvn_mobility*lvn_mobility+-2.39400e-04*lvn_mobility+-3.95830e-03'
+ sky130_fd_pr__nfet_01v8__u0_diff_39 = '-3.60906e-05*lvn_mobility*lvn_mobility+-4.02112e-04*lvn_mobility+-3.76550e-03'
+ sky130_fd_pr__nfet_01v8__u0_diff_4 = '-1.44688e-05*lvn_mobility*lvn_mobility+-9.78750e-05*lvn_mobility+-1.75270e-03'
+ sky130_fd_pr__nfet_01v8__u0_diff_40 = '-9.37781e-05*lvn_mobility*lvn_mobility+3.60888e-04*lvn_mobility+1.92950e-03'
+ sky130_fd_pr__nfet_01v8__u0_diff_41 = '-8.78937e-05*lvn_mobility*lvn_mobility+-4.84000e-04*lvn_mobility+-6.66270e-03'
+ sky130_fd_pr__nfet_01v8__u0_diff_42 = '-6.41875e-05*lvn_mobility*lvn_mobility+-6.92550e-04*lvn_mobility+-5.08400e-03'
+ sky130_fd_pr__nfet_01v8__u0_diff_43 = '-6.43153e-05*lvn_mobility*lvn_mobility+-6.40239e-04*lvn_mobility+-2.37280e-03'
+ sky130_fd_pr__nfet_01v8__u0_diff_44 = '-3.69937e-05*lvn_mobility*lvn_mobility+-4.40425e-04*lvn_mobility+-7.55660e-03'
+ sky130_fd_pr__nfet_01v8__u0_diff_45 = '-3.51063e-05*lvn_mobility*lvn_mobility+-2.25300e-04*lvn_mobility+-4.32120e-03'
+ sky130_fd_pr__nfet_01v8__u0_diff_46 = '-2.58094e-05*lvn_mobility*lvn_mobility+-3.28387e-04*lvn_mobility+-2.64090e-03'
+ sky130_fd_pr__nfet_01v8__u0_diff_47 = '1.51094e-05*lvn_mobility*lvn_mobility+5.11687e-04*lvn_mobility+-4.10870e-03'
+ sky130_fd_pr__nfet_01v8__u0_diff_48 = '-8.01200e-05*lvn_mobility*lvn_mobility+-6.72770e-04*lvn_mobility+-2.10610e-03'
+ sky130_fd_pr__nfet_01v8__u0_diff_49 = '-5.47625e-05*lvn_mobility*lvn_mobility+5.70000e-05*lvn_mobility+-2.91030e-03'
+ sky130_fd_pr__nfet_01v8__u0_diff_5 = '-1.33437e-05*lvn_mobility*lvn_mobility+-1.65925e-04*lvn_mobility+-2.13500e-03'
+ sky130_fd_pr__nfet_01v8__u0_diff_50 = '-1.06641e-05*lvn_mobility*lvn_mobility+6.09869e-04*lvn_mobility+-2.71830e-03'
+ sky130_fd_pr__nfet_01v8__u0_diff_51 = '-2.86319e-05*lvn_mobility*lvn_mobility+3.73023e-04*lvn_mobility'
+ sky130_fd_pr__nfet_01v8__u0_diff_52 = '-2.37247e-04*lvn_mobility*lvn_mobility+3.55538e-04*lvn_mobility+-3.13230e-03'
+ sky130_fd_pr__nfet_01v8__u0_diff_53 = '-1.61281e-04*lvn_mobility*lvn_mobility+4.51625e-04*lvn_mobility+-2.90360e-03'
+ sky130_fd_pr__nfet_01v8__u0_diff_54 = '-4.65912e-05*lvn_mobility*lvn_mobility+-6.57850e-05*lvn_mobility'
+ sky130_fd_pr__nfet_01v8__u0_diff_55 = '-1.27769e-05*lvn_mobility*lvn_mobility+1.89463e-04*lvn_mobility'
+ sky130_fd_pr__nfet_01v8__u0_diff_56 = '-4.04112e-05*lvn_mobility*lvn_mobility+-3.25105e-04*lvn_mobility'
+ sky130_fd_pr__nfet_01v8__u0_diff_57 = '-5.57719e-05*lvn_mobility*lvn_mobility+-6.17837e-04*lvn_mobility'
+ sky130_fd_pr__nfet_01v8__u0_diff_58 = '-6.01281e-05*lvn_mobility*lvn_mobility+-6.57087e-04*lvn_mobility'
+ sky130_fd_pr__nfet_01v8__u0_diff_59 = '-1.07150e-04*lvn_mobility*lvn_mobility+-8.53200e-04*lvn_mobility'
+ sky130_fd_pr__nfet_01v8__u0_diff_6 = '-2.60656e-05*lvn_mobility*lvn_mobility+4.59038e-04*lvn_mobility+-3.90890e-03'
+ sky130_fd_pr__nfet_01v8__u0_diff_60 = '-7.39672e-05*lvn_mobility*lvn_mobility+-4.91106e-04*lvn_mobility'
+ sky130_fd_pr__nfet_01v8__u0_diff_61 = '-1.01219e-04*lvn_mobility*lvn_mobility+-1.16565e-03*lvn_mobility'
+ sky130_fd_pr__nfet_01v8__u0_diff_62 = '-9.16531e-05*lvn_mobility*lvn_mobility+-7.28088e-04*lvn_mobility'
+ sky130_fd_pr__nfet_01v8__u0_diff_7 = '-1.01750e-05*lvn_mobility*lvn_mobility+-1.08775e-04*lvn_mobility+-3.73740e-03'
+ sky130_fd_pr__nfet_01v8__u0_diff_8 = '-7.90406e-05*lvn_mobility*lvn_mobility+-1.27304e-03*lvn_mobility+-5.20520e-03'
+ sky130_fd_pr__nfet_01v8__u0_diff_9 = '-1.45781e-05*lvn_mobility*lvn_mobility+-6.47375e-05*lvn_mobility+-2.59860e-03'
+ sky130_fd_pr__nfet_01v8__ua_diff_0 = '3.84213e-12*lvn_mobility*lvn_mobility+5.58350e-12*lvn_mobility+1.39350e-11'
+ sky130_fd_pr__nfet_01v8__ua_diff_1 = '2.95259e-12*lvn_mobility*lvn_mobility+6.55412e-12*lvn_mobility+1.03810e-11'
+ sky130_fd_pr__nfet_01v8__ua_diff_10 = '2.25768e-12*lvn_mobility*lvn_mobility+3.68863e-12*lvn_mobility+6.53870e-12'
+ sky130_fd_pr__nfet_01v8__ua_diff_11 = '9.80418e-14*lvn_mobility*lvn_mobility+-4.24396e-13*lvn_mobility+3.59480e-14'
+ sky130_fd_pr__nfet_01v8__ua_diff_12 = '1.38266e-13*lvn_mobility*lvn_mobility+-3.75637e-13*lvn_mobility+8.17920e-12'
+ sky130_fd_pr__nfet_01v8__ua_diff_13 = '-8.13550e-13*lvn_mobility*lvn_mobility+-5.20162e-12*lvn_mobility+8.16830e-12'
+ sky130_fd_pr__nfet_01v8__ua_diff_14 = '1.33734e-13*lvn_mobility*lvn_mobility+-7.84762e-13*lvn_mobility+5.86820e-12'
+ sky130_fd_pr__nfet_01v8__ua_diff_15 = '5.54809e-13*lvn_mobility*lvn_mobility+-4.36126e-12*lvn_mobility+1.38180e-11'
+ sky130_fd_pr__nfet_01v8__ua_diff_16 = '3.10531e-13*lvn_mobility*lvn_mobility+-1.82330e-12*lvn_mobility+7.43030e-12'
+ sky130_fd_pr__nfet_01v8__ua_diff_17 = '1.59625e-13*lvn_mobility*lvn_mobility+7.18225e-13*lvn_mobility+3.33770e-12'
+ sky130_fd_pr__nfet_01v8__ua_diff_18 = '7.31184e-14*lvn_mobility*lvn_mobility+-6.40726e-13*lvn_mobility+2.26840e-12'
+ sky130_fd_pr__nfet_01v8__ua_diff_19 = '3.09737e-14*lvn_mobility*lvn_mobility+-2.89325e-14*lvn_mobility+4.42090e-13'
+ sky130_fd_pr__nfet_01v8__ua_diff_2 = '1.87183e-13*lvn_mobility*lvn_mobility+3.19863e-13*lvn_mobility+4.54620e-13'
+ sky130_fd_pr__nfet_01v8__ua_diff_20 = '2.01125e-13*lvn_mobility*lvn_mobility+-6.51750e-13*lvn_mobility+1.20210e-11'
+ sky130_fd_pr__nfet_01v8__ua_diff_21 = '1.30144e-13*lvn_mobility*lvn_mobility+-3.86875e-13*lvn_mobility+7.49520e-12'
+ sky130_fd_pr__nfet_01v8__ua_diff_22 = '1.04291e-13*lvn_mobility*lvn_mobility+-5.78837e-13*lvn_mobility+4.08040e-12'
+ sky130_fd_pr__nfet_01v8__ua_diff_23 = '-2.54063e-13*lvn_mobility*lvn_mobility+-4.48000e-12*lvn_mobility+-6.85990e-13'
+ sky130_fd_pr__nfet_01v8__ua_diff_24 = '1.00712e-12*lvn_mobility*lvn_mobility+-3.00550e-12*lvn_mobility+2.52290e-11'
+ sky130_fd_pr__nfet_01v8__ua_diff_25 = '2.13497e-13*lvn_mobility*lvn_mobility+9.64737e-13*lvn_mobility+2.72610e-12'
+ sky130_fd_pr__nfet_01v8__ua_diff_26 = '2.36606e-14*lvn_mobility*lvn_mobility+-8.37175e-13*lvn_mobility+-1.47270e-13'
+ sky130_fd_pr__nfet_01v8__ua_diff_27 = '1.00531e-13*lvn_mobility*lvn_mobility+-3.64475e-13*lvn_mobility+4.67450e-12'
+ sky130_fd_pr__nfet_01v8__ua_diff_28 = '8.25500e-14*lvn_mobility*lvn_mobility+-1.21175e-13*lvn_mobility+4.78560e-12'
+ sky130_fd_pr__nfet_01v8__ua_diff_29 = '6.84781e-14*lvn_mobility*lvn_mobility+-1.62375e-14*lvn_mobility+3.79530e-12'
+ sky130_fd_pr__nfet_01v8__ua_diff_3 = '6.63819e-14*lvn_mobility*lvn_mobility+4.79432e-13*lvn_mobility+5.22860e-13'
+ sky130_fd_pr__nfet_01v8__ua_diff_30 = '5.78000e-14*lvn_mobility*lvn_mobility+-5.50750e-14*lvn_mobility+2.90640e-12'
+ sky130_fd_pr__nfet_01v8__ua_diff_31 = '2.12782e-12*lvn_mobility*lvn_mobility+6.54126e-12*lvn_mobility+-6.15620e-12'
+ sky130_fd_pr__nfet_01v8__ua_diff_32 = '8.45000e-13*lvn_mobility*lvn_mobility+-3.16750e-12*lvn_mobility+2.04070e-11'
+ sky130_fd_pr__nfet_01v8__ua_diff_33 = '2.56778e-13*lvn_mobility*lvn_mobility+1.12251e-12*lvn_mobility+3.60450e-12'
+ sky130_fd_pr__nfet_01v8__ua_diff_34 = '2.59168e-14*lvn_mobility*lvn_mobility+-8.25575e-13*lvn_mobility+3.63060e-15'
+ sky130_fd_pr__nfet_01v8__ua_diff_35 = '5.74406e-13*lvn_mobility*lvn_mobility+2.10463e-12*lvn_mobility+1.42920e-11'
+ sky130_fd_pr__nfet_01v8__ua_diff_36 = '1.73394e-13*lvn_mobility*lvn_mobility+4.74775e-13*lvn_mobility+7.43060e-12'
+ sky130_fd_pr__nfet_01v8__ua_diff_37 = '4.01250e-13*lvn_mobility*lvn_mobility+1.01000e-13*lvn_mobility+1.73340e-11'
+ sky130_fd_pr__nfet_01v8__ua_diff_38 = '2.25969e-13*lvn_mobility*lvn_mobility+-2.24375e-13*lvn_mobility+1.03350e-11'
+ sky130_fd_pr__nfet_01v8__ua_diff_39 = '-9.60188e-14*lvn_mobility*lvn_mobility+-9.00875e-13*lvn_mobility+8.76080e-12'
+ sky130_fd_pr__nfet_01v8__ua_diff_4 = '9.36156e-14*lvn_mobility*lvn_mobility+-2.56437e-13*lvn_mobility+4.18970e-12'
+ sky130_fd_pr__nfet_01v8__ua_diff_40 = '1.23310e-12*lvn_mobility*lvn_mobility+-1.48421e-12*lvn_mobility+-6.38250e-12'
+ sky130_fd_pr__nfet_01v8__ua_diff_41 = '2.54181e-12*lvn_mobility*lvn_mobility+5.95750e-12*lvn_mobility+2.75640e-11'
+ sky130_fd_pr__nfet_01v8__ua_diff_42 = '1.63156e-13*lvn_mobility*lvn_mobility+7.32875e-13*lvn_mobility+1.54710e-11'
+ sky130_fd_pr__nfet_01v8__ua_diff_43 = '2.00634e-13*lvn_mobility*lvn_mobility+1.66984e-12*lvn_mobility+5.50550e-12'
+ sky130_fd_pr__nfet_01v8__ua_diff_44 = '3.68250e-13*lvn_mobility*lvn_mobility+-2.89750e-13*lvn_mobility+2.00250e-11'
+ sky130_fd_pr__nfet_01v8__ua_diff_45 = '2.51437e-13*lvn_mobility*lvn_mobility+-2.11750e-13*lvn_mobility+1.14580e-11'
+ sky130_fd_pr__nfet_01v8__ua_diff_46 = '1.55753e-13*lvn_mobility*lvn_mobility+2.90013e-13*lvn_mobility+6.46290e-12'
+ sky130_fd_pr__nfet_01v8__ua_diff_47 = '4.27953e-12*lvn_mobility*lvn_mobility+-1.34981e-11*lvn_mobility+1.63150e-11'
+ sky130_fd_pr__nfet_01v8__ua_diff_48 = '-4.32666e-12*lvn_mobility*lvn_mobility+-1.80467e-11*lvn_mobility+3.93320e-12'
+ sky130_fd_pr__nfet_01v8__ua_diff_49 = '3.58147e-12*lvn_mobility*lvn_mobility+9.16987e-12*lvn_mobility+1.14870e-11'
+ sky130_fd_pr__nfet_01v8__ua_diff_5 = '1.07928e-13*lvn_mobility*lvn_mobility+-8.50875e-14*lvn_mobility+5.03360e-12'
+ sky130_fd_pr__nfet_01v8__ua_diff_50 = '1.21353e-12*lvn_mobility*lvn_mobility+-1.87363e-12*lvn_mobility+1.06290e-11'
+ sky130_fd_pr__nfet_01v8__ua_diff_51 = '2.20748e-12*lvn_mobility*lvn_mobility+2.78343e-12*lvn_mobility'
+ sky130_fd_pr__nfet_01v8__ua_diff_52 = '-8.94306e-13*lvn_mobility*lvn_mobility+6.48447e-12*lvn_mobility'
+ sky130_fd_pr__nfet_01v8__ua_diff_53 = '2.49861e-13*lvn_mobility*lvn_mobility+2.24851e-12*lvn_mobility'
+ sky130_fd_pr__nfet_01v8__ua_diff_54 = '3.70812e-12*lvn_mobility*lvn_mobility+-1.11995e-11*lvn_mobility'
+ sky130_fd_pr__nfet_01v8__ua_diff_55 = '4.09590e-12*lvn_mobility*lvn_mobility+-1.27574e-11*lvn_mobility'
+ sky130_fd_pr__nfet_01v8__ua_diff_56 = '4.04600e-12*lvn_mobility*lvn_mobility+-5.10256e-12*lvn_mobility'
+ sky130_fd_pr__nfet_01v8__ua_diff_57 = '3.88983e-12*lvn_mobility*lvn_mobility+-5.71250e-15*lvn_mobility'
+ sky130_fd_pr__nfet_01v8__ua_diff_58 = '3.81208e-12*lvn_mobility*lvn_mobility+2.40867e-12*lvn_mobility'
+ sky130_fd_pr__nfet_01v8__ua_diff_59 = '3.42089e-12*lvn_mobility*lvn_mobility+8.42639e-12*lvn_mobility'
+ sky130_fd_pr__nfet_01v8__ua_diff_6 = '3.44894e-12*lvn_mobility*lvn_mobility+6.18550e-12*lvn_mobility+1.49190e-11'
+ sky130_fd_pr__nfet_01v8__ua_diff_60 = '3.42089e-12*lvn_mobility*lvn_mobility+8.42639e-12*lvn_mobility'
+ sky130_fd_pr__nfet_01v8__ua_diff_61 = '1.83287e-12*lvn_mobility*lvn_mobility+9.60850e-12*lvn_mobility'
+ sky130_fd_pr__nfet_01v8__ua_diff_62 = '-4.32665e-12*lvn_mobility*lvn_mobility+-1.80467e-11*lvn_mobility'
+ sky130_fd_pr__nfet_01v8__ua_diff_7 = '3.95350e-12*lvn_mobility*lvn_mobility+1.40183e-11*lvn_mobility+1.47410e-11'
+ sky130_fd_pr__nfet_01v8__ua_diff_8 = '1.83287e-12*lvn_mobility*lvn_mobility+9.60850e-12*lvn_mobility+1.93880e-11'
+ sky130_fd_pr__nfet_01v8__ua_diff_9 = '1.49697e-13*lvn_mobility*lvn_mobility+-5.33363e-13*lvn_mobility+6.05940e-12'
+ sky130_fd_pr__nfet_01v8__ub_diff_0 = '-6.72156e-21*lvn_mobility*lvn_mobility+-2.70112e-20*lvn_mobility+-1.16750e-19'
+ sky130_fd_pr__nfet_01v8__ub_diff_1 = '-7.35572e-21*lvn_mobility*lvn_mobility+-5.75321e-20*lvn_mobility+-1.69790e-19'
+ sky130_fd_pr__nfet_01v8__ub_diff_10 = '-5.95000e-21*lvn_mobility*lvn_mobility+-4.71550e-20*lvn_mobility+-1.67730e-19'
+ sky130_fd_pr__nfet_01v8__ub_diff_11 = '-2.00672e-21*lvn_mobility*lvn_mobility+-2.68984e-20*lvn_mobility+6.11940e-20'
+ sky130_fd_pr__nfet_01v8__ub_diff_12 = '-2.07200e-21*lvn_mobility*lvn_mobility+-4.34595e-20*lvn_mobility+-2.26030e-19'
+ sky130_fd_pr__nfet_01v8__ub_diff_13 = '-4.07500e-22*lvn_mobility*lvn_mobility+-5.54250e-21*lvn_mobility+-2.10770e-19'
+ sky130_fd_pr__nfet_01v8__ub_diff_14 = '-1.54156e-21*lvn_mobility*lvn_mobility+-1.59313e-20*lvn_mobility+-1.72380e-19'
+ sky130_fd_pr__nfet_01v8__ub_diff_15 = '-2.17719e-21*lvn_mobility*lvn_mobility+2.40162e-20*lvn_mobility+-3.65250e-19'
+ sky130_fd_pr__nfet_01v8__ub_diff_16 = '-3.37581e-21*lvn_mobility*lvn_mobility+-3.46362e-20*lvn_mobility+-3.93420e-20'
+ sky130_fd_pr__nfet_01v8__ub_diff_17 = '-3.01675e-21*lvn_mobility*lvn_mobility+-3.58263e-20*lvn_mobility+8.18030e-20'
+ sky130_fd_pr__nfet_01v8__ub_diff_18 = '-1.55100e-21*lvn_mobility*lvn_mobility+-1.87215e-20*lvn_mobility+5.98900e-20'
+ sky130_fd_pr__nfet_01v8__ub_diff_19 = '-1.54099e-21*lvn_mobility*lvn_mobility+-1.57402e-20*lvn_mobility+8.08050e-20'
+ sky130_fd_pr__nfet_01v8__ub_diff_2 = '-2.98222e-21*lvn_mobility*lvn_mobility+-4.00739e-20*lvn_mobility+1.65480e-19'
+ sky130_fd_pr__nfet_01v8__ub_diff_20 = '-1.77781e-21*lvn_mobility*lvn_mobility+-3.18888e-20*lvn_mobility+-3.41490e-19'
+ sky130_fd_pr__nfet_01v8__ub_diff_21 = '-1.64281e-21*lvn_mobility*lvn_mobility+-2.92913e-20*lvn_mobility+-2.42570e-19'
+ sky130_fd_pr__nfet_01v8__ub_diff_22 = '-1.37744e-21*lvn_mobility*lvn_mobility+-1.25327e-20*lvn_mobility+-8.90700e-20'
+ sky130_fd_pr__nfet_01v8__ub_diff_23 = '-5.92500e-23*lvn_mobility*lvn_mobility+3.42235e-20*lvn_mobility+5.44640e-20'
+ sky130_fd_pr__nfet_01v8__ub_diff_24 = '-2.56969e-21*lvn_mobility*lvn_mobility+2.38750e-22*lvn_mobility+-4.48400e-19'
+ sky130_fd_pr__nfet_01v8__ub_diff_25 = '-2.65135e-21*lvn_mobility*lvn_mobility+-2.51654e-20*lvn_mobility+1.36750e-19'
+ sky130_fd_pr__nfet_01v8__ub_diff_26 = '-1.15075e-21*lvn_mobility*lvn_mobility+-4.96749e-21*lvn_mobility+3.15990e-20'
+ sky130_fd_pr__nfet_01v8__ub_diff_27 = '-1.56503e-21*lvn_mobility*lvn_mobility+-1.65546e-20*lvn_mobility+-1.00310e-20'
+ sky130_fd_pr__nfet_01v8__ub_diff_28 = '-1.65556e-21*lvn_mobility*lvn_mobility+-2.86882e-20*lvn_mobility+-7.35480e-20'
+ sky130_fd_pr__nfet_01v8__ub_diff_29 = '-1.64519e-21*lvn_mobility*lvn_mobility+-3.13983e-20*lvn_mobility+-4.18640e-20'
+ sky130_fd_pr__nfet_01v8__ub_diff_3 = '-2.77500e-21*lvn_mobility*lvn_mobility+-4.91287e-20*lvn_mobility+9.83550e-20'
+ sky130_fd_pr__nfet_01v8__ub_diff_30 = '-1.34403e-21*lvn_mobility*lvn_mobility+-2.05494e-20*lvn_mobility+-6.35080e-20'
+ sky130_fd_pr__nfet_01v8__ub_diff_31 = '-2.59562e-21*lvn_mobility*lvn_mobility+8.32000e-21*lvn_mobility+2.64240e-19'
+ sky130_fd_pr__nfet_01v8__ub_diff_32 = '-2.71406e-21*lvn_mobility*lvn_mobility+5.15375e-21*lvn_mobility+-3.05350e-19'
+ sky130_fd_pr__nfet_01v8__ub_diff_33 = '-2.61844e-21*lvn_mobility*lvn_mobility+-2.13215e-20*lvn_mobility+9.67890e-20'
+ sky130_fd_pr__nfet_01v8__ub_diff_34 = '-1.18216e-21*lvn_mobility*lvn_mobility+-6.78937e-21*lvn_mobility+2.10290e-20'
+ sky130_fd_pr__nfet_01v8__ub_diff_35 = '-6.78178e-21*lvn_mobility*lvn_mobility+-7.64729e-20*lvn_mobility+-1.06700e-19'
+ sky130_fd_pr__nfet_01v8__ub_diff_36 = '-3.53281e-21*lvn_mobility*lvn_mobility+-7.29562e-20*lvn_mobility+-1.17200e-19'
+ sky130_fd_pr__nfet_01v8__ub_diff_37 = '-5.48241e-21*lvn_mobility*lvn_mobility+-7.66854e-20*lvn_mobility+-2.48860e-19'
+ sky130_fd_pr__nfet_01v8__ub_diff_38 = '-4.22094e-21*lvn_mobility*lvn_mobility+-6.92388e-20*lvn_mobility+-1.01550e-19'
+ sky130_fd_pr__nfet_01v8__ub_diff_39 = '-3.53016e-21*lvn_mobility*lvn_mobility+-7.24944e-20*lvn_mobility+-1.63340e-19'
+ sky130_fd_pr__nfet_01v8__ub_diff_4 = '-2.04331e-21*lvn_mobility*lvn_mobility+-4.11950e-20*lvn_mobility+-1.62470e-20'
+ sky130_fd_pr__nfet_01v8__ub_diff_40 = '-9.09125e-21*lvn_mobility*lvn_mobility+-8.78650e-20*lvn_mobility+6.55000e-19'
+ sky130_fd_pr__nfet_01v8__ub_diff_41 = '-8.46875e-21*lvn_mobility*lvn_mobility+-1.57645e-19*lvn_mobility+-2.27360e-19'
+ sky130_fd_pr__nfet_01v8__ub_diff_42 = '-5.18469e-21*lvn_mobility*lvn_mobility+-9.76962e-20*lvn_mobility+-1.30380e-19'
+ sky130_fd_pr__nfet_01v8__ub_diff_43 = '-6.00806e-21*lvn_mobility*lvn_mobility+-8.11263e-20*lvn_mobility+5.32840e-20'
+ sky130_fd_pr__nfet_01v8__ub_diff_44 = '-4.08469e-21*lvn_mobility*lvn_mobility+-7.68262e-20*lvn_mobility+-4.82090e-19'
+ sky130_fd_pr__nfet_01v8__ub_diff_45 = '-3.86963e-21*lvn_mobility*lvn_mobility+-5.59690e-20*lvn_mobility+-1.95090e-19'
+ sky130_fd_pr__nfet_01v8__ub_diff_46 = '-2.93187e-21*lvn_mobility*lvn_mobility+-5.86612e-20*lvn_mobility+-7.45030e-22'
+ sky130_fd_pr__nfet_01v8__ub_diff_47 = '-1.73026e-21*lvn_mobility*lvn_mobility+2.56802e-20*lvn_mobility+-6.69850e-20'
+ sky130_fd_pr__nfet_01v8__ub_diff_48 = '-3.99387e-22*lvn_mobility*lvn_mobility+-6.44525e-20*lvn_mobility+-3.75980e-21'
+ sky130_fd_pr__nfet_01v8__ub_diff_49 = '-8.91219e-21*lvn_mobility*lvn_mobility+-1.19659e-19*lvn_mobility+-1.30930e-19'
+ sky130_fd_pr__nfet_01v8__ub_diff_5 = '-1.88538e-21*lvn_mobility*lvn_mobility+-4.24613e-20*lvn_mobility+-2.19790e-20'
+ sky130_fd_pr__nfet_01v8__ub_diff_50 = '-2.76611e-21*lvn_mobility*lvn_mobility+-2.02952e-20*lvn_mobility+-4.81130e-21'
+ sky130_fd_pr__nfet_01v8__ub_diff_51 = '-5.22284e-21*lvn_mobility*lvn_mobility+-6.24046e-20*lvn_mobility'
+ sky130_fd_pr__nfet_01v8__ub_diff_52 = '-1.59262e-20*lvn_mobility*lvn_mobility+-1.67728e-19*lvn_mobility'
+ sky130_fd_pr__nfet_01v8__ub_diff_53 = '-1.20702e-20*lvn_mobility*lvn_mobility+-1.24730e-19*lvn_mobility'
+ sky130_fd_pr__nfet_01v8__ub_diff_54 = '-2.90361e-21*lvn_mobility*lvn_mobility+4.47132e-21*lvn_mobility'
+ sky130_fd_pr__nfet_01v8__ub_diff_55 = '-2.09722e-21*lvn_mobility*lvn_mobility+1.88696e-20*lvn_mobility'
+ sky130_fd_pr__nfet_01v8__ub_diff_56 = '-4.56945e-21*lvn_mobility*lvn_mobility+-2.86792e-20*lvn_mobility'
+ sky130_fd_pr__nfet_01v8__ub_diff_57 = '-6.18966e-21*lvn_mobility*lvn_mobility+-6.13751e-20*lvn_mobility'
+ sky130_fd_pr__nfet_01v8__ub_diff_58 = '-6.93009e-21*lvn_mobility*lvn_mobility+-7.67831e-20*lvn_mobility'
+ sky130_fd_pr__nfet_01v8__ub_diff_59 = '-8.46431e-21*lvn_mobility*lvn_mobility+-1.13021e-19*lvn_mobility'
+ sky130_fd_pr__nfet_01v8__ub_diff_6 = '-8.39844e-21*lvn_mobility*lvn_mobility+-7.75813e-20*lvn_mobility+-3.44300e-19'
+ sky130_fd_pr__nfet_01v8__ub_diff_60 = '-8.46431e-21*lvn_mobility*lvn_mobility+-1.13021e-19*lvn_mobility'
+ sky130_fd_pr__nfet_01v8__ub_diff_61 = '-1.01141e-20*lvn_mobility*lvn_mobility+-1.55569e-19*lvn_mobility'
+ sky130_fd_pr__nfet_01v8__ub_diff_62 = '-3.99375e-22*lvn_mobility*lvn_mobility+-6.44525e-20*lvn_mobility'
+ sky130_fd_pr__nfet_01v8__ub_diff_7 = '-7.19787e-21*lvn_mobility*lvn_mobility+-1.10406e-19*lvn_mobility+-2.51130e-19'
+ sky130_fd_pr__nfet_01v8__ub_diff_8 = '-1.01141e-20*lvn_mobility*lvn_mobility+-1.55569e-19*lvn_mobility+-7.59090e-20'
+ sky130_fd_pr__nfet_01v8__ub_diff_9 = '-2.38741e-21*lvn_mobility*lvn_mobility+-3.57479e-20*lvn_mobility+-1.18010e-19'
+ sky130_fd_pr__nfet_01v8__voff_diff_42 = '-1.25000e-03*lvn_subvt*lvn_subvt+-5.00000e-03*lvn_subvt'
+ sky130_fd_pr__nfet_01v8__vsat_diff_0 = '7.09474e+02*lvn_saturation*lvn_saturation+1.17592e+04*lvn_saturation+5.94410e+02'
+ sky130_fd_pr__nfet_01v8__vsat_diff_1 = '1.52729e+02*lvn_saturation*lvn_saturation+7.53112e+03*lvn_saturation+2.49830e+02'
+ sky130_fd_pr__nfet_01v8__vsat_diff_10 = '2.23662e+02*lvn_saturation*lvn_saturation+7.94875e+03*lvn_saturation+-3.16260e+03'
+ sky130_fd_pr__nfet_01v8__vsat_diff_15 = '2.69429e+02*lvn_saturation*lvn_saturation+7.55350e+03*lvn_saturation+-6.47870e+02'
+ sky130_fd_pr__nfet_01v8__vsat_diff_16 = '3.62381e+02*lvn_saturation*lvn_saturation+7.10150e+03*lvn_saturation+-1.58610e+03'
+ sky130_fd_pr__nfet_01v8__vsat_diff_17 = '6.09281e+02*lvn_saturation*lvn_saturation+7.54788e+03*lvn_saturation+-3.38400e+03'
+ sky130_fd_pr__nfet_01v8__vsat_diff_18 = '7.61531e+01*lvn_saturation*lvn_saturation+3.23781e+03*lvn_saturation+2.23030e+03'
+ sky130_fd_pr__nfet_01v8__vsat_diff_23 = '1.70319e+02*lvn_saturation*lvn_saturation+6.72600e+03*lvn_saturation+4.44490e+03'
+ sky130_fd_pr__nfet_01v8__vsat_diff_24 = '1.98919e+02*lvn_saturation*lvn_saturation+5.05962e+03*lvn_saturation+-1.45120e+03'
+ sky130_fd_pr__nfet_01v8__vsat_diff_25 = '4.32406e+02*lvn_saturation*lvn_saturation+5.77375e+03*lvn_saturation+-3.53350e+03'
+ sky130_fd_pr__nfet_01v8__vsat_diff_26 = '2.45594e+01*lvn_saturation*lvn_saturation+2.18921e+03*lvn_saturation+-3.04310e+03'
+ sky130_fd_pr__nfet_01v8__vsat_diff_31 = '8.80187e+01*lvn_saturation*lvn_saturation+5.45425e+03*lvn_saturation+5.59670e+03'
+ sky130_fd_pr__nfet_01v8__vsat_diff_32 = '2.03096e+02*lvn_saturation*lvn_saturation+5.19212e+03*lvn_saturation+-3.60040e+02'
+ sky130_fd_pr__nfet_01v8__vsat_diff_33 = '4.97444e+02*lvn_saturation*lvn_saturation+6.21538e+03*lvn_saturation+-3.88360e+03'
+ sky130_fd_pr__nfet_01v8__vsat_diff_34 = '1.90437e+01*lvn_saturation*lvn_saturation+1.92215e+03*lvn_saturation+-1.50430e+03'
+ sky130_fd_pr__nfet_01v8__vsat_diff_40 = '3.89909e+02*lvn_saturation*lvn_saturation+1.59162e+04*lvn_saturation+-1.05370e+01'
+ sky130_fd_pr__nfet_01v8__vsat_diff_41 = '2.30675e+03*lvn_saturation*lvn_saturation+7.95950e+03*lvn_saturation+-1.45440e+04'
+ sky130_fd_pr__nfet_01v8__vsat_diff_42 = '1.21966e+03*lvn_saturation*lvn_saturation+-4.14300e+02*lvn_saturation+-1.48840e+04'
+ sky130_fd_pr__nfet_01v8__vsat_diff_47 = '7.42744e+02*lvn_saturation*lvn_saturation+1.45985e+04*lvn_saturation+-1.43690e+03'
+ sky130_fd_pr__nfet_01v8__vsat_diff_48 = '1.90759e+03*lvn_saturation*lvn_saturation+1.78664e+04*lvn_saturation+-1.23460e+04'
+ sky130_fd_pr__nfet_01v8__vsat_diff_49 = '8.13200e+02*lvn_saturation*lvn_saturation+1.31471e+04*lvn_saturation+2.64330e+03'
+ sky130_fd_pr__nfet_01v8__vsat_diff_50 = '9.90925e+02*lvn_saturation*lvn_saturation+1.32719e+04*lvn_saturation+5.76370e+03'
+ sky130_fd_pr__nfet_01v8__vsat_diff_51 = '9.15613e+02*lvn_saturation*lvn_saturation+1.32436e+04*lvn_saturation'
+ sky130_fd_pr__nfet_01v8__vsat_diff_52 = '4.11062e+01*lvn_saturation*lvn_saturation+1.57946e+04*lvn_saturation+-2.54620e+03'
+ sky130_fd_pr__nfet_01v8__vsat_diff_53 = '3.84625e+01*lvn_saturation*lvn_saturation+1.44640e+04*lvn_saturation+-1.95040e+03'
+ sky130_fd_pr__nfet_01v8__vsat_diff_54 = '1.59831e+03*lvn_saturation*lvn_saturation+1.86568e+04*lvn_saturation'
+ sky130_fd_pr__nfet_01v8__vsat_diff_55 = '1.24697e+03*lvn_saturation*lvn_saturation+1.69561e+04*lvn_saturation'
+ sky130_fd_pr__nfet_01v8__vsat_diff_56 = '2.37288e+03*lvn_saturation*lvn_saturation+2.15210e+04*lvn_saturation'
+ sky130_fd_pr__nfet_01v8__vsat_diff_57 = '3.81800e+03*lvn_saturation*lvn_saturation+2.75955e+04*lvn_saturation'
+ sky130_fd_pr__nfet_01v8__vsat_diff_58 = '3.85119e+03*lvn_saturation*lvn_saturation+2.78478e+04*lvn_saturation'
+ sky130_fd_pr__nfet_01v8__vsat_diff_59 = '2.71669e+03*lvn_saturation*lvn_saturation+2.14882e+04*lvn_saturation'
+ sky130_fd_pr__nfet_01v8__vsat_diff_6 = '3.62862e+02*lvn_saturation*lvn_saturation+1.00955e+04*lvn_saturation+-2.39180e+03'
+ sky130_fd_pr__nfet_01v8__vsat_diff_60 = '1.95016e+03*lvn_saturation*lvn_saturation+1.81569e+04*lvn_saturation'
+ sky130_fd_pr__nfet_01v8__vsat_diff_61 = '1.78216e+03*lvn_saturation*lvn_saturation+1.65241e+04*lvn_saturation'
+ sky130_fd_pr__nfet_01v8__vsat_diff_62 = '4.67028e+03*lvn_saturation*lvn_saturation+3.10614e+04*lvn_saturation'
+ sky130_fd_pr__nfet_01v8__vsat_diff_7 = '5.76819e+02*lvn_saturation*lvn_saturation+9.95512e+03*lvn_saturation+-5.17260e+03'
+ sky130_fd_pr__nfet_01v8__vsat_diff_8 = '5.61125e+02*lvn_saturation*lvn_saturation+8.09275e+03*lvn_saturation+-1.36730e+04'
+ sky130_fd_pr__nfet_01v8__vsat_diff_9 = '2.13875e+02*lvn_saturation*lvn_saturation+5.02938e+03*lvn_saturation+-6.75850e+03'
+ sky130_fd_pr__nfet_01v8__vth0_diff_0 = '-3.20594e-04*lvn_threshold*lvn_threshold+1.97749e-02*lvn_threshold+-2.44410e-02'
+ sky130_fd_pr__nfet_01v8__vth0_diff_1 = '-3.51837e-04*lvn_threshold*lvn_threshold+1.97401e-02*lvn_threshold+6.49090e-03'
+ sky130_fd_pr__nfet_01v8__vth0_diff_10 = '-2.98250e-04*lvn_threshold*lvn_threshold+1.75417e-02*lvn_threshold+4.97300e-03'
+ sky130_fd_pr__nfet_01v8__vth0_diff_11 = '-2.43031e-05*lvn_threshold*lvn_threshold+1.06164e-03*lvn_threshold+5.85760e-03'
+ sky130_fd_pr__nfet_01v8__vth0_diff_12 = '-1.93437e-05*lvn_threshold*lvn_threshold+3.73750e-05*lvn_threshold+-1.08730e-02'
+ sky130_fd_pr__nfet_01v8__vth0_diff_13 = '-5.60500e-05*lvn_threshold*lvn_threshold+1.53207e-03*lvn_threshold+-7.49090e-03'
+ sky130_fd_pr__nfet_01v8__vth0_diff_14 = '-2.18437e-05*lvn_threshold*lvn_threshold+2.98850e-04*lvn_threshold+-7.39820e-03'
+ sky130_fd_pr__nfet_01v8__vth0_diff_15 = '-2.50094e-04*lvn_threshold*lvn_threshold+1.69979e-02*lvn_threshold+-1.80990e-02'
+ sky130_fd_pr__nfet_01v8__vth0_diff_16 = '-4.64187e-05*lvn_threshold*lvn_threshold+1.00962e-02*lvn_threshold+-3.91930e-03'
+ sky130_fd_pr__nfet_01v8__vth0_diff_17 = '-2.00281e-05*lvn_threshold*lvn_threshold+4.29489e-03*lvn_threshold+-1.84420e-02'
+ sky130_fd_pr__nfet_01v8__vth0_diff_18 = '1.85944e-06*lvn_threshold*lvn_threshold+2.14489e-03*lvn_threshold+-8.57020e-03'
+ sky130_fd_pr__nfet_01v8__vth0_diff_19 = '-7.74375e-06*lvn_threshold*lvn_threshold+-1.66075e-04*lvn_threshold+2.22920e-03'
+ sky130_fd_pr__nfet_01v8__vth0_diff_2 = '-6.27813e-05*lvn_threshold*lvn_threshold+3.11655e-03*lvn_threshold+6.56330e-03'
+ sky130_fd_pr__nfet_01v8__vth0_diff_20 = '-1.73750e-05*lvn_threshold*lvn_threshold+5.15750e-04*lvn_threshold+-1.36280e-02'
+ sky130_fd_pr__nfet_01v8__vth0_diff_21 = '-1.62188e-05*lvn_threshold*lvn_threshold+-1.63875e-04*lvn_threshold+-1.10820e-02'
+ sky130_fd_pr__nfet_01v8__vth0_diff_22 = '-1.90687e-05*lvn_threshold*lvn_threshold+5.52200e-04*lvn_threshold+-4.04530e-03'
+ sky130_fd_pr__nfet_01v8__vth0_diff_23 = '-2.53350e-04*lvn_threshold*lvn_threshold+1.58884e-02*lvn_threshold+-3.87790e-03'
+ sky130_fd_pr__nfet_01v8__vth0_diff_24 = '-3.57188e-05*lvn_threshold*lvn_threshold+9.77562e-03*lvn_threshold+-2.17450e-02'
+ sky130_fd_pr__nfet_01v8__vth0_diff_25 = '-4.26250e-06*lvn_threshold*lvn_threshold+3.52237e-03*lvn_threshold+-3.52730e-03'
+ sky130_fd_pr__nfet_01v8__vth0_diff_26 = '5.64062e-06*lvn_threshold*lvn_threshold+2.45611e-03*lvn_threshold+-3.43180e-03'
+ sky130_fd_pr__nfet_01v8__vth0_diff_27 = '-1.39687e-05*lvn_threshold*lvn_threshold+-8.86250e-05*lvn_threshold+-1.33240e-02'
+ sky130_fd_pr__nfet_01v8__vth0_diff_28 = '-1.74875e-05*lvn_threshold*lvn_threshold+-3.11675e-04*lvn_threshold+-6.87920e-03'
+ sky130_fd_pr__nfet_01v8__vth0_diff_29 = '-1.54813e-05*lvn_threshold*lvn_threshold+-1.93775e-04*lvn_threshold+-9.51120e-03'
+ sky130_fd_pr__nfet_01v8__vth0_diff_3 = '-5.18188e-05*lvn_threshold*lvn_threshold+2.67343e-03*lvn_threshold+-1.63620e-03'
+ sky130_fd_pr__nfet_01v8__vth0_diff_30 = '-1.36670e-05*lvn_threshold*lvn_threshold+-6.75932e-04*lvn_threshold+-2.39070e-03'
+ sky130_fd_pr__nfet_01v8__vth0_diff_31 = '-1.93244e-04*lvn_threshold*lvn_threshold+1.21945e-02*lvn_threshold+3.66890e-03'
+ sky130_fd_pr__nfet_01v8__vth0_diff_32 = '-3.78750e-05*lvn_threshold*lvn_threshold+7.79850e-03*lvn_threshold+-1.95640e-02'
+ sky130_fd_pr__nfet_01v8__vth0_diff_33 = '-4.21563e-06*lvn_threshold*lvn_threshold+2.61654e-03*lvn_threshold+-6.04640e-03'
+ sky130_fd_pr__nfet_01v8__vth0_diff_34 = '6.61875e-06*lvn_threshold*lvn_threshold+2.28225e-03*lvn_threshold+-6.02990e-03'
+ sky130_fd_pr__nfet_01v8__vth0_diff_35 = '-2.03437e-04*lvn_threshold*lvn_threshold+8.41625e-03*lvn_threshold+-1.08410e-02'
+ sky130_fd_pr__nfet_01v8__vth0_diff_36 = '-1.64084e-04*lvn_threshold*lvn_threshold+-1.27574e-03*lvn_threshold+-8.21770e-03'
+ sky130_fd_pr__nfet_01v8__vth0_diff_37 = '-1.36531e-04*lvn_threshold*lvn_threshold+6.07687e-03*lvn_threshold+-3.96450e-02'
+ sky130_fd_pr__nfet_01v8__vth0_diff_38 = '-1.11625e-04*lvn_threshold*lvn_threshold+3.41975e-03*lvn_threshold+-2.60400e-02'
+ sky130_fd_pr__nfet_01v8__vth0_diff_39 = '-1.45347e-04*lvn_threshold*lvn_threshold+3.67962e-04*lvn_threshold+-4.46610e-03'
+ sky130_fd_pr__nfet_01v8__vth0_diff_4 = '-3.26469e-05*lvn_threshold*lvn_threshold+1.56989e-03*lvn_threshold+-8.28310e-03'
+ sky130_fd_pr__nfet_01v8__vth0_diff_40 = '-5.71250e-05*lvn_threshold*lvn_threshold+3.17300e-02*lvn_threshold+-2.11360e-02'
+ sky130_fd_pr__nfet_01v8__vth0_diff_41 = '-5.90031e-04*lvn_threshold*lvn_threshold+2.06576e-02*lvn_threshold+-3.93390e-02'
+ sky130_fd_pr__nfet_01v8__vth0_diff_42 = '7.19375e-05*lvn_threshold*lvn_threshold+8.78950e-03*lvn_threshold+-1.16110e-02'
+ sky130_fd_pr__nfet_01v8__vth0_diff_43 = '-1.98212e-04*lvn_threshold*lvn_threshold+6.19263e-03*lvn_threshold+2.76090e-03'
+ sky130_fd_pr__nfet_01v8__vth0_diff_44 = '-8.29563e-05*lvn_threshold*lvn_threshold+3.98818e-03*lvn_threshold+-2.21110e-02'
+ sky130_fd_pr__nfet_01v8__vth0_diff_45 = '-8.25781e-05*lvn_threshold*lvn_threshold+3.02966e-03*lvn_threshold+-9.38710e-03'
+ sky130_fd_pr__nfet_01v8__vth0_diff_46 = '-9.13812e-05*lvn_threshold*lvn_threshold+6.20825e-04*lvn_threshold+-2.40930e-03'
+ sky130_fd_pr__nfet_01v8__vth0_diff_47 = '2.87500e-04*lvn_threshold*lvn_threshold+3.40500e-02*lvn_threshold+-2.21800e-02'
+ sky130_fd_pr__nfet_01v8__vth0_diff_48 = '-2.00906e-04*lvn_threshold*lvn_threshold+6.99988e-03*lvn_threshold+-1.02260e-02'
+ sky130_fd_pr__nfet_01v8__vth0_diff_49 = '-3.88375e-04*lvn_threshold*lvn_threshold+2.47857e-02*lvn_threshold+1.13610e-02'
+ sky130_fd_pr__nfet_01v8__vth0_diff_5 = '-3.73719e-05*lvn_threshold*lvn_threshold+2.20138e-04*lvn_threshold+-9.42950e-03'
+ sky130_fd_pr__nfet_01v8__vth0_diff_50 = '-3.35500e-04*lvn_threshold*lvn_threshold+2.48002e-02*lvn_threshold+-1.74810e-02'
+ sky130_fd_pr__nfet_01v8__vth0_diff_51 = '-3.58060e-04*lvn_threshold*lvn_threshold+2.47965e-02*lvn_threshold'
+ sky130_fd_pr__nfet_01v8__vth0_diff_52 = '-1.23063e-04*lvn_threshold*lvn_threshold+4.05688e-02*lvn_threshold+4.20040e-02'
+ sky130_fd_pr__nfet_01v8__vth0_diff_53 = '-7.83750e-05*lvn_threshold*lvn_threshold+4.00962e-02*lvn_threshold+3.21090e-02'
+ sky130_fd_pr__nfet_01v8__vth0_diff_54 = '-1.35625e-04*lvn_threshold*lvn_threshold+3.79525e-02*lvn_threshold'
+ sky130_fd_pr__nfet_01v8__vth0_diff_55 = '-1.38437e-04*lvn_threshold*lvn_threshold+3.68438e-02*lvn_threshold'
+ sky130_fd_pr__nfet_01v8__vth0_diff_56 = '-2.30625e-04*lvn_threshold*lvn_threshold+3.55175e-02*lvn_threshold'
+ sky130_fd_pr__nfet_01v8__vth0_diff_57 = '-2.83438e-04*lvn_threshold*lvn_threshold+3.42262e-02*lvn_threshold'
+ sky130_fd_pr__nfet_01v8__vth0_diff_58 = '-3.18750e-04*lvn_threshold*lvn_threshold+3.37650e-02*lvn_threshold'
+ sky130_fd_pr__nfet_01v8__vth0_diff_59 = '-4.11250e-04*lvn_threshold*lvn_threshold+3.29000e-02*lvn_threshold'
+ sky130_fd_pr__nfet_01v8__vth0_diff_6 = '-3.94069e-04*lvn_threshold*lvn_threshold+2.09175e-02*lvn_threshold+-1.51290e-03'
+ sky130_fd_pr__nfet_01v8__vth0_diff_60 = '-1.75344e-04*lvn_threshold*lvn_threshold+2.32764e-02*lvn_threshold'
+ sky130_fd_pr__nfet_01v8__vth0_diff_61 = '-2.67469e-04*lvn_threshold*lvn_threshold+1.07809e-02*lvn_threshold'
+ sky130_fd_pr__nfet_01v8__vth0_diff_62 = '-2.28219e-04*lvn_threshold*lvn_threshold+8.48662e-03*lvn_threshold'
+ sky130_fd_pr__nfet_01v8__vth0_diff_7 = '-1.00156e-04*lvn_threshold*lvn_threshold+1.35479e-02*lvn_threshold+-1.22030e-02'
+ sky130_fd_pr__nfet_01v8__vth0_diff_8 = '-2.57312e-04*lvn_threshold*lvn_threshold+7.41500e-03*lvn_threshold+-1.00360e-02'
+ sky130_fd_pr__nfet_01v8__vth0_diff_9 = '-3.24062e-05*lvn_threshold*lvn_threshold+3.24788e-03*lvn_threshold+1.98500e-03'
+ sky130_fd_pr__nfet_01v8__wint_diff = '8.04375e-09*diff_cd'
+ sky130_fd_pr__esd_nfet_01v8__ajunction_mult = '-6.25000e-07*lvn_diode*lvn_diode+5.53700e-02*lvn_diode+9.95430e-01'
+ sky130_fd_pr__esd_nfet_01v8__dlc_diff = '-5.05994e-11*poly_cd*poly_cd+-3.24937e-09*poly_cd+-6.14910e-10'
+ sky130_fd_pr__esd_nfet_01v8__dwc_diff = '8.04375e-09*diff_cd'
+ sky130_fd_pr__esd_nfet_01v8__k2_diff_0 = '4.43913e-04*lvn_bodyeffect*lvn_bodyeffect+-5.74310e-03*lvn_bodyeffect+1.76280e-02'
+ sky130_fd_pr__esd_nfet_01v8__k2_diff_1 = '3.98588e-04*lvn_bodyeffect*lvn_bodyeffect+-5.11850e-03*lvn_bodyeffect+-3.04040e-03'
+ sky130_fd_pr__esd_nfet_01v8__k2_diff_2 = '2.59872e-04*lvn_bodyeffect*lvn_bodyeffect+-3.80556e-03*lvn_bodyeffect+3.28980e-03'
+ sky130_fd_pr__esd_nfet_01v8__lint_diff = '-4.33125e-09*poly_cd'
+ sky130_fd_pr__esd_nfet_01v8__nfactor_diff_0 = '6.32993e-03*lvn_subvt*lvn_subvt+5.56838e-02*lvn_subvt+4.38610e-03'
+ sky130_fd_pr__esd_nfet_01v8__nfactor_diff_1 = '9.06125e-03*lvn_subvt*lvn_subvt+2.91225e-02*lvn_subvt+-5.31690e-01'
+ sky130_fd_pr__esd_nfet_01v8__nfactor_diff_2 = '8.35813e-03*lvn_subvt*lvn_subvt+2.15100e-02*lvn_subvt+-6.67760e-01'
+ sky130_fd_pr__esd_nfet_01v8__overlap_mult = '-2.66875e-04*lvtox*lvtox+1.14425e-02*lvtox+9.84200e-01'
+ sky130_fd_pr__esd_nfet_01v8__pjunction_mult = '-1.25000e-06*lvn_diode*lvn_diode+5.67550e-02*lvn_diode+1.02040e+00'
+ sky130_fd_pr__esd_nfet_01v8__toxe_mult = '1.30000e-02*lvtox+1.00000e+00'
+ sky130_fd_pr__esd_nfet_01v8__u0_diff_0 = '2.78625e-05*lvn_mobility*lvn_mobility+1.45907e-03*lvn_mobility+-3.81750e-03'
+ sky130_fd_pr__esd_nfet_01v8__u0_diff_1 = '3.35781e-05*lvn_mobility*lvn_mobility+1.58924e-03*lvn_mobility+-3.14350e-03'
+ sky130_fd_pr__esd_nfet_01v8__u0_diff_2 = '3.55094e-05*lvn_mobility*lvn_mobility+1.39709e-03*lvn_mobility+-4.34170e-03'
+ sky130_fd_pr__esd_nfet_01v8__ua_diff_0 = '5.15581e-12*lvn_mobility*lvn_mobility+5.24075e-12*lvn_mobility+3.48540e-11'
+ sky130_fd_pr__esd_nfet_01v8__ua_diff_1 = '3.91206e-12*lvn_mobility*lvn_mobility+6.70925e-12*lvn_mobility+2.33900e-11'
+ sky130_fd_pr__esd_nfet_01v8__ua_diff_2 = '4.07072e-12*lvn_mobility*lvn_mobility+8.74338e-12*lvn_mobility+2.87150e-11'
+ sky130_fd_pr__esd_nfet_01v8__ub_diff_0 = '-4.68234e-21*lvn_mobility*lvn_mobility+8.93806e-20*lvn_mobility+-3.61550e-19'
+ sky130_fd_pr__esd_nfet_01v8__ub_diff_1 = '-2.14625e-21*lvn_mobility*lvn_mobility+9.83550e-20*lvn_mobility+-1.24960e-19'
+ sky130_fd_pr__esd_nfet_01v8__ub_diff_2 = '-2.79437e-21*lvn_mobility*lvn_mobility+6.78800e-20*lvn_mobility+-4.87630e-19'
+ sky130_fd_pr__esd_nfet_01v8__vsat_diff_0 = '2.28506e+02*lvn_saturation*lvn_saturation+7.65712e+03*lvn_saturation+-4.45260e+03'
+ sky130_fd_pr__esd_nfet_01v8__vsat_diff_1 = '-7.08011e+01*lvn_saturation*lvn_saturation+4.23062e+03*lvn_saturation+-9.36830e+01'
+ sky130_fd_pr__esd_nfet_01v8__vsat_diff_2 = '1.40144e+02*lvn_saturation*lvn_saturation+5.82562e+03*lvn_saturation+1.06020e+03'
+ sky130_fd_pr__esd_nfet_01v8__vth0_diff_0 = '-5.42006e-04*lvn_threshold*lvn_threshold+1.97986e-02*lvn_threshold+-8.44540e-03'
+ sky130_fd_pr__esd_nfet_01v8__vth0_diff_1 = '-4.66000e-04*lvn_threshold*lvn_threshold+1.88445e-02*lvn_threshold+-1.26510e-02'
+ sky130_fd_pr__esd_nfet_01v8__vth0_diff_2 = '-3.14781e-04*lvn_threshold*lvn_threshold+1.91984e-02*lvn_threshold+-1.55380e-02'
+ sky130_fd_pr__esd_nfet_01v8__wint_diff = '8.04375e-09*diff_cd'
+ sky130_fd_pr__nfet_03v3_nvt__ajunction_mult = '-1.87500e-06*hvn_diode*hvn_diode+1.02953e-01*hvn_diode+9.76020e-01'
+ sky130_fd_pr__nfet_03v3_nvt__dlc_diff = '9.86313e-10*poly_cd*poly_cd+-7.50000e-09*poly_cd+-1.57810e-08'
+ sky130_fd_pr__nfet_03v3_nvt__dwc_diff = '8.04375e-09*diff_cd'
+ sky130_fd_pr__nfet_03v3_nvt__k2_diff_0 = '-1.53563e-04*hvn_bodyeffect*hvn_bodyeffect+6.48713e-03*hvn_bodyeffect+1.91350e-03'
+ sky130_fd_pr__nfet_03v3_nvt__k2_diff_1 = '-9.16781e-05*hvn_bodyeffect*hvn_bodyeffect+3.45939e-03*hvn_bodyeffect+9.67430e-03'
+ sky130_fd_pr__nfet_03v3_nvt__k2_diff_2 = '-2.04419e-05*hvn_bodyeffect*hvn_bodyeffect+1.56259e-03*hvn_bodyeffect+5.77670e-03'
+ sky130_fd_pr__nfet_03v3_nvt__k2_diff_3 = '-1.63819e-04*hvn_bodyeffect*hvn_bodyeffect+6.07375e-03*hvn_bodyeffect+3.27210e-03'
+ sky130_fd_pr__nfet_03v3_nvt__k2_diff_4 = '-1.20169e-04*hvn_bodyeffect*hvn_bodyeffect+2.84050e-04*hvn_bodyeffect+1.00040e-02'
+ sky130_fd_pr__nfet_03v3_nvt__k2_diff_5 = '-2.98969e-05*hvn_bodyeffect*hvn_bodyeffect+2.32684e-03*hvn_bodyeffect+1.27150e-02'
+ sky130_fd_pr__nfet_03v3_nvt__k2_diff_6 = '-3.09000e-05*hvn_bodyeffect*hvn_bodyeffect+2.13685e-03*hvn_bodyeffect+1.20660e-02'
+ sky130_fd_pr__nfet_03v3_nvt__k2_diff_7 = '-1.13381e-04*hvn_bodyeffect*hvn_bodyeffect+3.09352e-03*hvn_bodyeffect+1.11170e-02'
+ sky130_fd_pr__nfet_03v3_nvt__k2_diff_8 = '-3.59781e-05*hvn_bodyeffect*hvn_bodyeffect+1.49849e-03*hvn_bodyeffect+8.47970e-03'
+ sky130_fd_pr__nfet_03v3_nvt__lint_diff = '-4.33125e-09*poly_cd'
+ sky130_fd_pr__nfet_03v3_nvt__nfactor_diff_0 = '-2.07188e-03*hvn_subvt*hvn_subvt+-9.57625e-02*hvn_subvt+-1.38380e+00'
+ sky130_fd_pr__nfet_03v3_nvt__nfactor_diff_1 = '-1.39031e-02*hvn_subvt*hvn_subvt+2.21875e-02*hvn_subvt+-1.39580e+00'
+ sky130_fd_pr__nfet_03v3_nvt__nfactor_diff_2 = '4.80625e-04*hvn_subvt*hvn_subvt+5.11000e-03*hvn_subvt+-4.65030e-01'
+ sky130_fd_pr__nfet_03v3_nvt__nfactor_diff_3 = '-2.09125e-03*hvn_subvt*hvn_subvt+-1.10060e-01*hvn_subvt+-1.36210e+00'
+ sky130_fd_pr__nfet_03v3_nvt__nfactor_diff_4 = '-6.67812e-03*hvn_subvt*hvn_subvt+6.17125e-02*hvn_subvt+-1.34040e+00'
+ sky130_fd_pr__nfet_03v3_nvt__nfactor_diff_5 = '1.92500e-03*hvn_subvt*hvn_subvt+-9.12500e-03*hvn_subvt+-1.64340e+00'
+ sky130_fd_pr__nfet_03v3_nvt__nfactor_diff_6 = '1.63438e-03*hvn_subvt*hvn_subvt+4.66500e-03*hvn_subvt+-7.46000e-01'
+ sky130_fd_pr__nfet_03v3_nvt__nfactor_diff_7 = '-1.02438e-02*hvn_subvt*hvn_subvt+8.05000e-03*hvn_subvt+-1.34360e+00'
+ sky130_fd_pr__nfet_03v3_nvt__nfactor_diff_8 = '6.08125e-04*hvn_subvt*hvn_subvt+2.39550e-02*hvn_subvt+-4.37240e-01'
+ sky130_fd_pr__nfet_03v3_nvt__overlap_mult = '7.40406e-03*hvtox*hvtox+1.20091e-01*hvtox+7.71170e-01'
+ sky130_fd_pr__nfet_03v3_nvt__pjunction_mult = '-3.12500e-07*hvn_diode*hvn_diode+5.06762e-02*hvn_diode+1.04370e+00'
+ sky130_fd_pr__nfet_03v3_nvt__toxe_mult = '1.30000e-02*hvtox+1.00000e+00'
+ sky130_fd_pr__nfet_03v3_nvt__u0_diff_0 = '-6.24522e-05*hvn_mobility*hvn_mobility+-4.56099e-04*hvn_mobility+-6.56970e-04'
+ sky130_fd_pr__nfet_03v3_nvt__u0_diff_1 = '-9.07750e-05*hvn_mobility*hvn_mobility+6.29500e-05*hvn_mobility+-1.15940e-03'
+ sky130_fd_pr__nfet_03v3_nvt__u0_diff_2 = '-5.09822e-05*hvn_mobility*hvn_mobility+1.47733e-03*hvn_mobility+6.32540e-03'
+ sky130_fd_pr__nfet_03v3_nvt__u0_diff_3 = '-9.15600e-05*hvn_mobility*hvn_mobility+-6.82875e-04*hvn_mobility+-1.10740e-04'
+ sky130_fd_pr__nfet_03v3_nvt__u0_diff_4 = '1.25828e-04*hvn_mobility*hvn_mobility+3.20487e-04*hvn_mobility+-1.88560e-03'
+ sky130_fd_pr__nfet_03v3_nvt__u0_diff_5 = '-2.02756e-04*hvn_mobility*hvn_mobility+-2.46625e-04*hvn_mobility+1.12410e-02'
+ sky130_fd_pr__nfet_03v3_nvt__u0_diff_6 = '-1.29997e-04*hvn_mobility*hvn_mobility+-2.02963e-04*hvn_mobility+7.88100e-03'
+ sky130_fd_pr__nfet_03v3_nvt__u0_diff_7 = '-7.02625e-05*hvn_mobility*hvn_mobility+-6.15275e-04*hvn_mobility+-1.76890e-03'
+ sky130_fd_pr__nfet_03v3_nvt__u0_diff_8 = '-9.27019e-05*hvn_mobility*hvn_mobility+9.01008e-04*hvn_mobility+5.95200e-03'
+ sky130_fd_pr__nfet_03v3_nvt__ua_diff_0 = '3.50625e-14*hvn_mobility*hvn_mobility+-5.93600e-12*hvn_mobility+3.49770e-11'
+ sky130_fd_pr__nfet_03v3_nvt__ua_diff_1 = '1.53853e-12*hvn_mobility*hvn_mobility+-1.28913e-12*hvn_mobility+5.34070e-11'
+ sky130_fd_pr__nfet_03v3_nvt__ua_diff_2 = '4.12563e-13*hvn_mobility*hvn_mobility+5.89600e-12*hvn_mobility+5.82040e-11'
+ sky130_fd_pr__nfet_03v3_nvt__ua_diff_3 = '2.43597e-12*hvn_mobility*hvn_mobility+4.61762e-12*hvn_mobility+3.73970e-11'
+ sky130_fd_pr__nfet_03v3_nvt__ua_diff_4 = '1.63500e-13*hvn_mobility*hvn_mobility+-3.64850e-12*hvn_mobility+2.22680e-11'
+ sky130_fd_pr__nfet_03v3_nvt__ua_diff_5 = '1.87872e-12*hvn_mobility*hvn_mobility+1.52754e-11*hvn_mobility+7.29690e-11'
+ sky130_fd_pr__nfet_03v3_nvt__ua_diff_6 = '4.43409e-12*hvn_mobility*hvn_mobility+2.19319e-11*hvn_mobility+8.57370e-11'
+ sky130_fd_pr__nfet_03v3_nvt__ua_diff_7 = '-1.15409e-12*hvn_mobility*hvn_mobility+-1.19221e-11*hvn_mobility+4.00610e-11'
+ sky130_fd_pr__nfet_03v3_nvt__ua_diff_8 = '-2.06165e-12*hvn_mobility*hvn_mobility+-5.70359e-12*hvn_mobility+5.55250e-11'
+ sky130_fd_pr__nfet_03v3_nvt__ub_diff_0 = '-9.28844e-21*hvn_mobility*hvn_mobility+-1.77516e-19*hvn_mobility+-1.41320e-19'
+ sky130_fd_pr__nfet_03v3_nvt__ub_diff_1 = '-1.73537e-20*hvn_mobility*hvn_mobility+-1.50575e-19*hvn_mobility+1.04290e-19'
+ sky130_fd_pr__nfet_03v3_nvt__ub_diff_2 = '5.45000e-21*hvn_mobility*hvn_mobility+4.09100e-19*hvn_mobility+2.60950e-18'
+ sky130_fd_pr__nfet_03v3_nvt__ub_diff_3 = '-3.28819e-20*hvn_mobility*hvn_mobility+-4.14170e-19*hvn_mobility+-3.33610e-19'
+ sky130_fd_pr__nfet_03v3_nvt__ub_diff_4 = '1.15728e-19*hvn_mobility*hvn_mobility+5.13355e-19*hvn_mobility+3.72240e-19'
+ sky130_fd_pr__nfet_03v3_nvt__ub_diff_5 = '-6.25937e-21*hvn_mobility*hvn_mobility+3.11513e-19*hvn_mobility+3.05970e-18'
+ sky130_fd_pr__nfet_03v3_nvt__ub_diff_6 = '-1.16094e-20*hvn_mobility*hvn_mobility+1.68012e-19*hvn_mobility+2.39730e-18'
+ sky130_fd_pr__nfet_03v3_nvt__ub_diff_7 = '7.50312e-21*hvn_mobility*hvn_mobility+-2.11445e-19*hvn_mobility+2.65470e-19'
+ sky130_fd_pr__nfet_03v3_nvt__ub_diff_8 = '2.65625e-22*hvn_mobility*hvn_mobility+2.90237e-19*hvn_mobility+2.46450e-18'
+ sky130_fd_pr__nfet_03v3_nvt__voff_diff_0 = '-2.48287e-04*hvn_subvt*hvn_subvt+8.88265e-03*hvn_subvt+3.84490e-02'
+ sky130_fd_pr__nfet_03v3_nvt__voff_diff_1 = '-8.10188e-04*hvn_subvt*hvn_subvt+1.02485e-02*hvn_subvt+3.30820e-02'
+ sky130_fd_pr__nfet_03v3_nvt__voff_diff_3 = '-2.09394e-04*hvn_subvt*hvn_subvt+9.99958e-03*hvn_subvt+4.06730e-02'
+ sky130_fd_pr__nfet_03v3_nvt__voff_diff_4 = '-1.26547e-03*hvn_subvt*hvn_subvt+-1.94287e-03*hvn_subvt+4.54530e-02'
+ sky130_fd_pr__nfet_03v3_nvt__voff_diff_7 = '-6.99647e-04*hvn_subvt*hvn_subvt+9.64659e-03*hvn_subvt+4.19300e-02'
+ sky130_fd_pr__nfet_03v3_nvt__vsat_diff_0 = '-3.11031e+01*hvn_saturation*hvn_saturation+-9.64125e+01*hvn_saturation+-3.83720e+03'
+ sky130_fd_pr__nfet_03v3_nvt__vsat_diff_1 = '1.41694e+01*hvn_saturation*hvn_saturation+1.86873e+03*hvn_saturation+-6.76380e+03'
+ sky130_fd_pr__nfet_03v3_nvt__vsat_diff_2 = '4.09813e+01*hvn_saturation*hvn_saturation+2.25872e+03*hvn_saturation+-4.05680e+03'
+ sky130_fd_pr__nfet_03v3_nvt__vsat_diff_3 = '-2.83000e+01*hvn_saturation*hvn_saturation+3.24725e+02*hvn_saturation+-4.39620e+03'
+ sky130_fd_pr__nfet_03v3_nvt__vsat_diff_4 = '-2.70219e+01*hvn_saturation*hvn_saturation+9.54388e+02*hvn_saturation+-8.37610e+03'
+ sky130_fd_pr__nfet_03v3_nvt__vsat_diff_5 = '-5.53031e+01*hvn_saturation*hvn_saturation+9.38238e+02*hvn_saturation+-6.84320e+03'
+ sky130_fd_pr__nfet_03v3_nvt__vsat_diff_6 = '-5.74375e+00*hvn_saturation*hvn_saturation+1.44970e+03*hvn_saturation+-3.53490e+03'
+ sky130_fd_pr__nfet_03v3_nvt__vsat_diff_7 = '4.76875e+00*hvn_saturation*hvn_saturation+1.60227e+03*hvn_saturation+-7.89320e+03'
+ sky130_fd_pr__nfet_03v3_nvt__vsat_diff_8 = '9.51750e+01*hvn_saturation*hvn_saturation+2.19348e+03*hvn_saturation+-5.52890e+03'
+ sky130_fd_pr__nfet_03v3_nvt__vth0_diff_0 = '9.58750e-05*hvn_threshold*hvn_threshold+8.24050e-03*hvn_threshold+-1.58360e-02'
+ sky130_fd_pr__nfet_03v3_nvt__vth0_diff_1 = '1.10000e-05*hvn_threshold*hvn_threshold+1.14372e-02*hvn_threshold+-1.53240e-02'
+ sky130_fd_pr__nfet_03v3_nvt__vth0_diff_2 = '7.45000e-06*hvn_threshold*hvn_threshold+1.34726e-02*hvn_threshold+3.23230e-03'
+ sky130_fd_pr__nfet_03v3_nvt__vth0_diff_3 = '4.54062e-05*hvn_threshold*hvn_threshold+7.61013e-03*hvn_threshold+-1.87500e-02'
+ sky130_fd_pr__nfet_03v3_nvt__vth0_diff_4 = '9.10906e-04*hvn_threshold*hvn_threshold+1.99769e-02*hvn_threshold+-1.83380e-02'
+ sky130_fd_pr__nfet_03v3_nvt__vth0_diff_5 = '2.38438e-06*hvn_threshold*hvn_threshold+1.33790e-02*hvn_threshold+5.18760e-02'
+ sky130_fd_pr__nfet_03v3_nvt__vth0_diff_6 = '1.35000e-05*hvn_threshold*hvn_threshold+9.29750e-03*hvn_threshold+2.20080e-02'
+ sky130_fd_pr__nfet_03v3_nvt__vth0_diff_7 = '1.10437e-04*hvn_threshold*hvn_threshold+1.03045e-02*hvn_threshold+-1.41540e-02'
+ sky130_fd_pr__nfet_03v3_nvt__vth0_diff_8 = '1.19375e-06*hvn_threshold*hvn_threshold+1.33917e-02*hvn_threshold+-3.47710e-03'
+ sky130_fd_pr__nfet_03v3_nvt__wint_diff = '8.04375e-09*diff_cd'
+ sky130_fd_pr__nfet_g5v0d16v0__ajunction_mult = '9.37500e-07*hvn_diode*hvn_diode+4.43837e-02*hvn_diode+9.95050e-01'
+ sky130_fd_pr__nfet_g5v0d16v0__cf_mult = '-6.25000e-02*nfet_g5v0d16v0*nfet_g5v0d16v0+1.00000e+00'
+ sky130_fd_pr__nfet_g5v0d16v0__cgdl_mult = '-6.25000e-02*nfet_g5v0d16v0*nfet_g5v0d16v0+1.00000e+00'
+ sky130_fd_pr__nfet_g5v0d16v0__cgdo_mult = '-6.25000e-02*nfet_g5v0d16v0*nfet_g5v0d16v0+1.00000e+00'
+ sky130_fd_pr__nfet_g5v0d16v0__cgsl_mult = '-6.25000e-02*nfet_g5v0d16v0*nfet_g5v0d16v0+1.00000e+00'
+ sky130_fd_pr__nfet_g5v0d16v0__cgso_mult = '-6.25000e-02*nfet_g5v0d16v0*nfet_g5v0d16v0+1.00000e+00'
+ sky130_fd_pr__nfet_g5v0d16v0__cjs_mult = '-6.25000e-02*nfet_g5v0d16v0*nfet_g5v0d16v0+1.00000e+00'
+ sky130_fd_pr__nfet_g5v0d16v0__cjswgs_mult = '-6.25000e-02*nfet_g5v0d16v0*nfet_g5v0d16v0+1.00000e+00'
+ sky130_fd_pr__nfet_g5v0d16v0__cjsws_mult = '-6.25000e-02*nfet_g5v0d16v0*nfet_g5v0d16v0+1.00000e+00'
+ sky130_fd_pr__nfet_g5v0d16v0__dlc_diff = '-4.33125e-09*poly_cd'
+ sky130_fd_pr__nfet_g5v0d16v0__dwc_diff = '8.04375e-09*diff_cd'
+ sky130_fd_pr__nfet_g5v0d16v0__lint_diff = '-4.33125e-09*poly_cd'
+ sky130_fd_pr__nfet_g5v0d16v0__overlap_mult = '1.14375e-04*hvtox*hvtox+2.24843e-01*hvtox+1.00000e+00'
+ sky130_fd_pr__nfet_g5v0d16v0__pjunction_mult = '1.87500e-06*hvn_diode*hvn_diode+5.91425e-02*hvn_diode+1.01440e+00'
+ sky130_fd_pr__nfet_g5v0d16v0__rdiff_mult = '1.33031e-02*nfet_g5v0d16v0*nfet_g5v0d16v0+1.57087e-01*nfet_g5v0d16v0+1.05880e+00'
+ sky130_fd_pr__nfet_g5v0d16v0__toxe_mult = '1.50000e-02*hvtox+1.00000e+00'
+ sky130_fd_pr__nfet_g5v0d16v0__toxp_mult = '-3.12500e-02*hvtox*hvtox+-1.25000e-01*hvtox+1.00000e+00'
+ sky130_fd_pr__nfet_g5v0d16v0__u0_diff_0 = '2.71181e-04*hvn_mobility*hvn_mobility+-4.83587e-03*hvn_mobility+-1.49140e-03'
+ sky130_fd_pr__nfet_g5v0d16v0__u0_diff_1 = '2.69350e-04*hvn_mobility*hvn_mobility+-4.08888e-03*hvn_mobility+-5.09310e-03'
+ sky130_fd_pr__nfet_g5v0d16v0__u0_diff_2 = '1.58044e-04*hvn_mobility*hvn_mobility+-3.99450e-03*hvn_mobility+-1.90570e-03'
+ sky130_fd_pr__nfet_g5v0d16v0__u0_diff_3 = '-5.32094e-05*hvn_mobility*hvn_mobility+-1.61681e-03*hvn_mobility+-1.38990e-03'
+ sky130_fd_pr__nfet_g5v0d16v0__u0_diff_4 = '-5.91031e-05*hvn_mobility*hvn_mobility+-1.50351e-03*hvn_mobility+-2.98810e-03'
+ sky130_fd_pr__nfet_g5v0d16v0__vth0_diff_0 = '-9.43750e-06*hvn_threshold*hvn_threshold+3.61550e-02*hvn_threshold+1.05210e-02'
+ sky130_fd_pr__nfet_g5v0d16v0__vth0_diff_1 = '-2.29756e-05*hvn_threshold*hvn_threshold+3.52888e-02*hvn_threshold+9.82610e-04'
+ sky130_fd_pr__nfet_g5v0d16v0__vth0_diff_2 = '-1.95625e-05*hvn_threshold*hvn_threshold+3.63600e-02*hvn_threshold+8.61300e-03'
+ sky130_fd_pr__nfet_g5v0d16v0__vth0_diff_3 = '2.59375e-05*hvn_threshold*hvn_threshold+2.71480e-02*hvn_threshold+1.08530e-02'
+ sky130_fd_pr__nfet_g5v0d16v0__vth0_diff_4 = '1.59375e-05*hvn_threshold*hvn_threshold+2.71535e-02*hvn_threshold+1.74610e-02'
+ sky130_fd_pr__nfet_g5v0d16v0__wint_diff = '8.04375e-09*diff_cd'
+ sky130_fd_pr__model__parasitic__diode_ps2nw__ajunction_mult = '6.93889e-18*well_diode*well_diode+4.81850e-02*well_diode+9.82860e-01'
+ sky130_fd_pr__model__parasitic__diode_ps2nw__pjunction_mult = '6.93889e-18*well_diode*well_diode+1.80650e-02*well_diode+9.89540e-01'
+ sky130_fd_pr__pfet_20v0__ajunction_mult = '3.10000e-04*hvp_diode*hvp_diode+1.81850e-02*hvp_diode+1.00000e+00'
+ sky130_fd_pr__pfet_20v0__dlc_diff = '2.17734e-09*poly_cd*poly_cd+-1.30406e-08*poly_cd'
+ sky130_fd_pr__pfet_20v0__dwc_diff = '8.04375e-09*pdiff_cd'
+ sky130_fd_pr__pfet_20v0__lint_diff = '-4.33125e-09*poly_cd'
+ sky130_fd_pr__pfet_20v0__overlap_mult = '1.85000e-02*hvtox*hvtox+2.99000e-01*hvtox+1.00000e+00'
+ sky130_fd_pr__pfet_20v0__pjunction_mult = '5.61250e-04*hvp_diode*hvp_diode+1.61550e-02*hvp_diode+1.00000e+00'
+ sky130_fd_pr__pfet_20v0__rdrift_mult = '6.55156e-03*pfet_20v0*pfet_20v0+6.84013e-02*pfet_20v0+9.17770e-01'
+ sky130_fd_pr__pfet_20v0__toxe_mult = '2.50000e-04*hvtox*hvtox+1.40000e-02*hvtox+1.00000e+00'
+ sky130_fd_pr__pfet_20v0__u0_diff = '1.20212e-04*hvp_mobility*hvp_mobility+-2.71625e-03*hvp_mobility+-1.24040e-03'
+ sky130_fd_pr__pfet_20v0__vth0_diff = '-2.11250e-05*hvp_threshold*hvp_threshold+-3.65555e-02*hvp_threshold+8.31760e-02'
+ sky130_fd_pr__pfet_20v0__wint_diff = '8.04375e-09*pdiff_cd'
+ sky130_fd_pr__pfet_01v8_hvt__a0_diff_10 = '2.52306e-04*lvhp_saturation*lvhp_saturation+-9.42350e-04*lvhp_saturation+1.92370e-03'
+ sky130_fd_pr__pfet_01v8_hvt__a0_diff_11 = '-2.81234e-04*lvhp_saturation*lvhp_saturation+2.32376e-03*lvhp_saturation+3.66080e-03'
+ sky130_fd_pr__pfet_01v8_hvt__a0_diff_12 = '-1.78934e-03*lvhp_saturation*lvhp_saturation+4.56022e-03*lvhp_saturation+4.63140e-03'
+ sky130_fd_pr__pfet_01v8_hvt__a0_diff_13 = '-1.05071e-03*lvhp_saturation*lvhp_saturation+1.48690e-03*lvhp_saturation+1.58990e-03'
+ sky130_fd_pr__pfet_01v8_hvt__a0_diff_18 = '3.04378e-03*lvhp_saturation*lvhp_saturation+-7.07263e-03*lvhp_saturation+-6.52630e-02'
+ sky130_fd_pr__pfet_01v8_hvt__a0_diff_19 = '4.19245e-03*lvhp_saturation*lvhp_saturation+4.37479e-03*lvhp_saturation+-8.90780e-02'
+ sky130_fd_pr__pfet_01v8_hvt__a0_diff_2 = '-3.27375e-04*lvhp_saturation*lvhp_saturation+-6.24113e-02*lvhp_saturation+-1.74370e-02'
+ sky130_fd_pr__pfet_01v8_hvt__a0_diff_20 = '2.88148e-03*lvhp_saturation*lvhp_saturation+1.50743e-03*lvhp_saturation+-5.58890e-02'
+ sky130_fd_pr__pfet_01v8_hvt__a0_diff_21 = '-2.00503e-03*lvhp_saturation*lvhp_saturation+1.04381e-02*lvhp_saturation+2.96450e-02'
+ sky130_fd_pr__pfet_01v8_hvt__a0_diff_26 = '5.44393e-03*lvhp_saturation*lvhp_saturation+2.30349e-03*lvhp_saturation+-9.96070e-02'
+ sky130_fd_pr__pfet_01v8_hvt__a0_diff_27 = '4.57466e-03*lvhp_saturation*lvhp_saturation+1.03346e-02*lvhp_saturation+-8.02170e-02'
+ sky130_fd_pr__pfet_01v8_hvt__a0_diff_28 = '7.44362e-04*lvhp_saturation*lvhp_saturation+-7.00150e-04*lvhp_saturation+-9.10920e-03'
+ sky130_fd_pr__pfet_01v8_hvt__a0_diff_29 = '2.17591e-04*lvhp_saturation*lvhp_saturation+-2.17712e-04*lvhp_saturation+-2.61060e-03'
+ sky130_fd_pr__pfet_01v8_hvt__a0_diff_3 = '1.06489e-03*lvhp_saturation*lvhp_saturation+-2.82903e-02*lvhp_saturation+-2.89930e-03'
+ sky130_fd_pr__pfet_01v8_hvt__a0_diff_33 = '-9.37500e-03*lvhp_saturation*lvhp_saturation+-3.75000e-02*lvhp_saturation'
+ sky130_fd_pr__pfet_01v8_hvt__a0_diff_4 = '1.16825e-03*lvhp_saturation*lvhp_saturation+-3.12605e-02*lvhp_saturation+4.14160e-02'
+ sky130_fd_pr__pfet_01v8_hvt__a0_diff_5 = '4.07437e-04*lvhp_saturation*lvhp_saturation+-2.07017e-02*lvhp_saturation+-3.75420e-02'
+ sky130_fd_pr__pfet_01v8_hvt__a0_diff_59 = '8.88562e-06*lvhp_saturation*lvhp_saturation+3.76285e-04*lvhp_saturation'
+ sky130_fd_pr__pfet_01v8_hvt__a0_diff_60 = '8.45750e-06*lvhp_saturation*lvhp_saturation+3.84450e-04*lvhp_saturation'
+ sky130_fd_pr__pfet_01v8_hvt__a0_diff_61 = '5.45688e-06*lvhp_saturation*lvhp_saturation+2.61618e-04*lvhp_saturation'
+ sky130_fd_pr__pfet_01v8_hvt__a0_diff_62 = '2.33469e-06*lvhp_saturation*lvhp_saturation+1.16289e-04*lvhp_saturation'
+ sky130_fd_pr__pfet_01v8_hvt__a0_diff_63 = '2.33469e-06*lvhp_saturation*lvhp_saturation+1.16289e-04*lvhp_saturation'
+ sky130_fd_pr__pfet_01v8_hvt__a0_diff_64 = '-2.58875e-06*lvhp_saturation*lvhp_saturation+-1.28937e-04*lvhp_saturation'
+ sky130_fd_pr__pfet_01v8_hvt__a0_diff_66 = '-1.65656e-06*lvhp_saturation*lvhp_saturation+-8.66237e-05*lvhp_saturation'
+ sky130_fd_pr__pfet_01v8_hvt__a0_diff_67 = '-2.70031e-06*lvhp_saturation*lvhp_saturation+-1.54634e-04*lvhp_saturation'
+ sky130_fd_pr__pfet_01v8_hvt__agidl_diff_59 = '-2.79584e-14*lvp_subvt*lvp_subvt+-1.18398e-12*lvp_subvt'
+ sky130_fd_pr__pfet_01v8_hvt__agidl_diff_60 = '-2.66119e-14*lvp_subvt*lvp_subvt+-1.20968e-12*lvp_subvt'
+ sky130_fd_pr__pfet_01v8_hvt__agidl_diff_61 = '-1.71700e-14*lvp_subvt*lvp_subvt+-8.23180e-13*lvp_subvt'
+ sky130_fd_pr__pfet_01v8_hvt__agidl_diff_62 = '-7.34625e-15*lvp_subvt*lvp_subvt+-3.65905e-13*lvp_subvt'
+ sky130_fd_pr__pfet_01v8_hvt__agidl_diff_63 = '-7.34625e-15*lvp_subvt*lvp_subvt+-3.65905e-13*lvp_subvt'
+ sky130_fd_pr__pfet_01v8_hvt__agidl_diff_64 = '-8.52500e-15*lvp_subvt*lvp_subvt+-4.24600e-13*lvp_subvt'
+ sky130_fd_pr__pfet_01v8_hvt__agidl_diff_66 = '2.34919e-15*lvp_subvt*lvp_subvt+1.22871e-13*lvp_subvt'
+ sky130_fd_pr__pfet_01v8_hvt__agidl_diff_67 = '3.82972e-15*lvp_subvt*lvp_subvt+2.19338e-13*lvp_subvt'
+ sky130_fd_pr__pfet_01v8_hvt__ags_diff_10 = '-9.80531e-05*lvhp_saturation*lvhp_saturation+4.01545e-04*lvhp_saturation+-5.31770e-04'
+ sky130_fd_pr__pfet_01v8_hvt__ags_diff_11 = '8.02281e-04*lvhp_saturation*lvhp_saturation+-3.56410e-03*lvhp_saturation+-1.27090e-03'
+ sky130_fd_pr__pfet_01v8_hvt__ags_diff_12 = '2.85175e-03*lvhp_saturation*lvhp_saturation+-7.03875e-03*lvhp_saturation+-6.18600e-03'
+ sky130_fd_pr__pfet_01v8_hvt__ags_diff_13 = '1.72285e-03*lvhp_saturation*lvhp_saturation+-3.30387e-03*lvhp_saturation+-2.93710e-03'
+ sky130_fd_pr__pfet_01v8_hvt__ags_diff_18 = '-2.29741e-03*lvhp_saturation*lvhp_saturation+5.15688e-03*lvhp_saturation+4.84340e-02'
+ sky130_fd_pr__pfet_01v8_hvt__ags_diff_19 = '-3.74273e-03*lvhp_saturation*lvhp_saturation+-4.42540e-03*lvhp_saturation+8.11240e-02'
+ sky130_fd_pr__pfet_01v8_hvt__ags_diff_2 = '-6.64813e-04*lvhp_saturation*lvhp_saturation+4.24788e-02*lvhp_saturation+1.31320e-02'
+ sky130_fd_pr__pfet_01v8_hvt__ags_diff_20 = '-2.56912e-03*lvhp_saturation*lvhp_saturation+-1.68822e-03*lvhp_saturation+5.06340e-02'
+ sky130_fd_pr__pfet_01v8_hvt__ags_diff_21 = '-4.43981e-03*lvhp_saturation*lvhp_saturation+-3.20900e-03*lvhp_saturation+1.99940e-02'
+ sky130_fd_pr__pfet_01v8_hvt__ags_diff_26 = '-4.06706e-03*lvhp_saturation*lvhp_saturation+-1.87225e-03*lvhp_saturation+7.50880e-02'
+ sky130_fd_pr__pfet_01v8_hvt__ags_diff_27 = '-3.98172e-03*lvhp_saturation*lvhp_saturation+-9.53713e-03*lvhp_saturation+7.13000e-02'
+ sky130_fd_pr__pfet_01v8_hvt__ags_diff_28 = '-1.27549e-03*lvhp_saturation*lvhp_saturation+1.03473e-03*lvhp_saturation+1.62690e-02'
+ sky130_fd_pr__pfet_01v8_hvt__ags_diff_29 = '-2.26715e-04*lvhp_saturation*lvhp_saturation+8.37612e-05*lvhp_saturation+3.29240e-03'
+ sky130_fd_pr__pfet_01v8_hvt__ags_diff_3 = '-1.29131e-03*lvhp_saturation*lvhp_saturation+2.50560e-02*lvhp_saturation+3.29500e-03'
+ sky130_fd_pr__pfet_01v8_hvt__ags_diff_4 = '-7.10469e-04*lvhp_saturation*lvhp_saturation+1.41151e-02*lvhp_saturation+-1.75890e-02'
+ sky130_fd_pr__pfet_01v8_hvt__ags_diff_5 = '-6.80375e-04*lvhp_saturation*lvhp_saturation+2.03152e-02*lvhp_saturation+3.96750e-02'
+ sky130_fd_pr__pfet_01v8_hvt__ags_diff_64 = '2.53000e-06*lvhp_saturation*lvhp_saturation+1.26018e-04*lvhp_saturation'
+ sky130_fd_pr__pfet_01v8_hvt__ajunction_mult = '-6.25000e-07*lvp_diode*lvp_diode+2.33625e-02*lvp_diode+9.83660e-01'
+ sky130_fd_pr__pfet_01v8_hvt__b0_diff_34 = '1.62434e-09*lvhp_saturation*lvhp_saturation+-2.75431e-08*lvhp_saturation+-6.40670e-08'
+ sky130_fd_pr__pfet_01v8_hvt__b0_diff_35 = '2.44183e-09*lvhp_saturation*lvhp_saturation+1.35698e-08*lvhp_saturation+-8.76200e-08'
+ sky130_fd_pr__pfet_01v8_hvt__b0_diff_36 = '-2.25081e-09*lvhp_saturation*lvhp_saturation+-1.80975e-08*lvhp_saturation+2.03010e-08'
+ sky130_fd_pr__pfet_01v8_hvt__b0_diff_37 = '1.02841e-09*lvhp_saturation*lvhp_saturation+-3.25456e-08*lvhp_saturation+-5.14020e-08'
+ sky130_fd_pr__pfet_01v8_hvt__b0_diff_38 = '-4.83363e-09*lvhp_saturation*lvhp_saturation+-3.04500e-08*lvhp_saturation+-2.53620e-08'
+ sky130_fd_pr__pfet_01v8_hvt__b0_diff_41 = '-2.36922e-09*lvhp_saturation*lvhp_saturation+-9.47687e-09*lvhp_saturation'
+ sky130_fd_pr__pfet_01v8_hvt__b0_diff_42 = '2.03513e-09*lvhp_saturation*lvhp_saturation+-4.19788e-08*lvhp_saturation+-9.38270e-08'
+ sky130_fd_pr__pfet_01v8_hvt__b0_diff_43 = '1.83800e-09*lvhp_saturation*lvhp_saturation+-3.12012e-08*lvhp_saturation+-3.97830e-08'
+ sky130_fd_pr__pfet_01v8_hvt__b0_diff_44 = '1.79172e-09*lvhp_saturation*lvhp_saturation+-3.40334e-08*lvhp_saturation+-6.99140e-08'
+ sky130_fd_pr__pfet_01v8_hvt__b0_diff_45 = '-3.54791e-09*lvhp_saturation*lvhp_saturation+-2.79161e-08*lvhp_saturation+2.24710e-08'
+ sky130_fd_pr__pfet_01v8_hvt__b0_diff_47 = '-2.55800e-09*lvhp_saturation*lvhp_saturation+-1.02320e-08*lvhp_saturation'
+ sky130_fd_pr__pfet_01v8_hvt__b0_diff_49 = '-1.82959e-09*lvhp_saturation*lvhp_saturation+-7.31838e-09*lvhp_saturation'
+ sky130_fd_pr__pfet_01v8_hvt__b0_diff_50 = '4.49422e-16*lvhp_saturation*lvhp_saturation+1.79769e-15*lvhp_saturation'
+ sky130_fd_pr__pfet_01v8_hvt__b0_diff_54 = '-1.82959e-09*lvhp_saturation*lvhp_saturation+-7.31838e-09*lvhp_saturation'
+ sky130_fd_pr__pfet_01v8_hvt__b0_diff_57 = '-4.54938e-09*lvhp_saturation*lvhp_saturation+-1.81975e-08*lvhp_saturation'
+ sky130_fd_pr__pfet_01v8_hvt__b0_diff_58 = '-2.84809e-09*lvhp_saturation*lvhp_saturation+-1.13924e-08*lvhp_saturation'
+ sky130_fd_pr__pfet_01v8_hvt__b0_diff_59 = '-3.37438e-09*lvhp_saturation*lvhp_saturation+-1.34975e-08*lvhp_saturation'
+ sky130_fd_pr__pfet_01v8_hvt__b0_diff_60 = '-4.13594e-09*lvhp_saturation*lvhp_saturation+-1.65437e-08*lvhp_saturation'
+ sky130_fd_pr__pfet_01v8_hvt__b0_diff_61 = '-5.23187e-09*lvhp_saturation*lvhp_saturation+-2.09275e-08*lvhp_saturation'
+ sky130_fd_pr__pfet_01v8_hvt__b0_diff_62 = '-5.51187e-09*lvhp_saturation*lvhp_saturation+-2.20475e-08*lvhp_saturation'
+ sky130_fd_pr__pfet_01v8_hvt__b0_diff_63 = '-4.62625e-09*lvhp_saturation*lvhp_saturation+-1.85050e-08*lvhp_saturation'
+ sky130_fd_pr__pfet_01v8_hvt__b0_diff_64 = '3.71862e-17*lvhp_saturation*lvhp_saturation+1.48745e-16*lvhp_saturation'
+ sky130_fd_pr__pfet_01v8_hvt__b0_diff_66 = '-5.45344e-09*lvhp_saturation*lvhp_saturation+-2.18137e-08*lvhp_saturation'
+ sky130_fd_pr__pfet_01v8_hvt__b0_diff_67 = '-5.54781e-09*lvhp_saturation*lvhp_saturation+-2.21913e-08*lvhp_saturation'
+ sky130_fd_pr__pfet_01v8_hvt__b1_diff_34 = '1.73324e-09*lvhp_saturation*lvhp_saturation+-5.71710e-09*lvhp_saturation+1.78730e-10'
+ sky130_fd_pr__pfet_01v8_hvt__b1_diff_35 = '1.60997e-09*lvhp_saturation*lvhp_saturation+4.16953e-09*lvhp_saturation+-6.76360e-09'
+ sky130_fd_pr__pfet_01v8_hvt__b1_diff_36 = '3.86362e-10*lvhp_saturation*lvhp_saturation+-2.21441e-09*lvhp_saturation+1.25570e-11'
+ sky130_fd_pr__pfet_01v8_hvt__b1_diff_37 = '4.13213e-10*lvhp_saturation*lvhp_saturation+1.36585e-09*lvhp_saturation+-2.17530e-09'
+ sky130_fd_pr__pfet_01v8_hvt__b1_diff_38 = '-3.80871e-09*lvhp_saturation*lvhp_saturation+5.02788e-08*lvhp_saturation+-5.65820e-12'
+ sky130_fd_pr__pfet_01v8_hvt__b1_diff_41 = '8.02875e-11*lvhp_saturation*lvhp_saturation+3.21150e-10*lvhp_saturation'
+ sky130_fd_pr__pfet_01v8_hvt__b1_diff_42 = '3.07022e-10*lvhp_saturation*lvhp_saturation+-1.16456e-09*lvhp_saturation+-1.24720e-10'
+ sky130_fd_pr__pfet_01v8_hvt__b1_diff_43 = '3.52550e-11*lvhp_saturation*lvhp_saturation+1.57595e-10*lvhp_saturation+-1.56320e-09'
+ sky130_fd_pr__pfet_01v8_hvt__b1_diff_44 = '2.87047e-11*lvhp_saturation*lvhp_saturation+-4.12724e-10*lvhp_saturation+2.03530e-10'
+ sky130_fd_pr__pfet_01v8_hvt__b1_diff_45 = '1.45038e-10*lvhp_saturation*lvhp_saturation+4.11874e-10*lvhp_saturation+2.92040e-11'
+ sky130_fd_pr__pfet_01v8_hvt__b1_diff_47 = '-9.21750e-11*lvhp_saturation*lvhp_saturation+-3.68700e-10*lvhp_saturation'
+ sky130_fd_pr__pfet_01v8_hvt__b1_diff_49 = '1.53400e-16*lvhp_saturation*lvhp_saturation+6.13600e-16*lvhp_saturation'
+ sky130_fd_pr__pfet_01v8_hvt__b1_diff_50 = '1.46945e-23*lvhp_saturation*lvhp_saturation+5.87780e-23*lvhp_saturation'
+ sky130_fd_pr__pfet_01v8_hvt__b1_diff_54 = '1.53400e-16*lvhp_saturation*lvhp_saturation+6.13600e-16*lvhp_saturation'
+ sky130_fd_pr__pfet_01v8_hvt__b1_diff_56 = '2.73263e-31*lvhp_saturation*lvhp_saturation+1.09305e-30*lvhp_saturation'
+ sky130_fd_pr__pfet_01v8_hvt__b1_diff_57 = '2.10686e-31*lvhp_saturation*lvhp_saturation+8.42744e-31*lvhp_saturation'
+ sky130_fd_pr__pfet_01v8_hvt__b1_diff_58 = '5.20578e-33*lvhp_saturation*lvhp_saturation+2.08231e-32*lvhp_saturation'
+ sky130_fd_pr__pfet_01v8_hvt__b1_diff_59 = '5.64634e-17*lvhp_saturation*lvhp_saturation+2.25854e-16*lvhp_saturation'
+ sky130_fd_pr__pfet_01v8_hvt__b1_diff_60 = '9.57556e-17*lvhp_saturation*lvhp_saturation+3.83023e-16*lvhp_saturation'
+ sky130_fd_pr__pfet_01v8_hvt__b1_diff_61 = '1.23187e-16*lvhp_saturation*lvhp_saturation+4.92750e-16*lvhp_saturation'
+ sky130_fd_pr__pfet_01v8_hvt__b1_diff_62 = '1.41807e-16*lvhp_saturation*lvhp_saturation+5.67228e-16*lvhp_saturation'
+ sky130_fd_pr__pfet_01v8_hvt__b1_diff_63 = '1.41807e-16*lvhp_saturation*lvhp_saturation+5.67228e-16*lvhp_saturation'
+ sky130_fd_pr__pfet_01v8_hvt__b1_diff_64 = '-9.78869e-20*lvhp_saturation*lvhp_saturation+-3.91548e-19*lvhp_saturation'
+ sky130_fd_pr__pfet_01v8_hvt__b1_diff_66 = '1.30770e-16*lvhp_saturation*lvhp_saturation+5.23079e-16*lvhp_saturation'
+ sky130_fd_pr__pfet_01v8_hvt__b1_diff_67 = '5.08119e-17*lvhp_saturation*lvhp_saturation+2.03248e-16*lvhp_saturation'
+ sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_64 = '2.37304e+03*lvp_subvt*lvp_subvt+1.18195e+05*lvp_subvt'
+ sky130_fd_pr__pfet_01v8_hvt__dlc_diff = '-4.33125e-09*poly_cd'
+ sky130_fd_pr__pfet_01v8_hvt__dwc_diff = '8.04375e-09*diff_cd'
+ sky130_fd_pr__pfet_01v8_hvt__eta0_diff_59 = '-9.38312e-06*lvhp_threshold*lvhp_threshold+-3.97363e-04*lvhp_threshold'
+ sky130_fd_pr__pfet_01v8_hvt__eta0_diff_60 = '-8.93125e-06*lvhp_threshold*lvhp_threshold+-4.05985e-04*lvhp_threshold'
+ sky130_fd_pr__pfet_01v8_hvt__eta0_diff_61 = '-5.76281e-06*lvhp_threshold*lvhp_threshold+-2.76271e-04*lvhp_threshold'
+ sky130_fd_pr__pfet_01v8_hvt__eta0_diff_62 = '-2.46562e-06*lvhp_threshold*lvhp_threshold+-1.22802e-04*lvhp_threshold'
+ sky130_fd_pr__pfet_01v8_hvt__eta0_diff_63 = '-2.46562e-06*lvhp_threshold*lvhp_threshold+-1.22802e-04*lvhp_threshold'
+ sky130_fd_pr__pfet_01v8_hvt__eta0_diff_66 = '-1.34800e-07*lvhp_threshold*lvhp_threshold+-7.03908e-06*lvhp_threshold'
+ sky130_fd_pr__pfet_01v8_hvt__eta0_diff_67 = '-2.19600e-07*lvhp_threshold*lvhp_threshold+-1.25650e-05*lvhp_threshold'
+ sky130_fd_pr__pfet_01v8_hvt__k2_diff_0 = '3.65916e-04*lvhp_bodyeffect*lvhp_bodyeffect+-8.85140e-04*lvhp_bodyeffect+-8.42000e-03'
+ sky130_fd_pr__pfet_01v8_hvt__k2_diff_1 = '4.38053e-04*lvhp_bodyeffect*lvhp_bodyeffect+-6.01213e-04*lvhp_bodyeffect+-1.62920e-02'
+ sky130_fd_pr__pfet_01v8_hvt__k2_diff_10 = '2.89966e-04*lvhp_bodyeffect*lvhp_bodyeffect+3.77363e-04*lvhp_bodyeffect+-1.32420e-02'
+ sky130_fd_pr__pfet_01v8_hvt__k2_diff_11 = '2.48925e-04*lvhp_bodyeffect*lvhp_bodyeffect+3.16700e-04*lvhp_bodyeffect+-1.44670e-02'
+ sky130_fd_pr__pfet_01v8_hvt__k2_diff_12 = '-3.02281e-05*lvhp_bodyeffect*lvhp_bodyeffect+1.67959e-03*lvhp_bodyeffect+-3.50300e-03'
+ sky130_fd_pr__pfet_01v8_hvt__k2_diff_13 = '1.19191e-04*lvhp_bodyeffect*lvhp_bodyeffect+1.23751e-03*lvhp_bodyeffect+-5.38700e-03'
+ sky130_fd_pr__pfet_01v8_hvt__k2_diff_14 = '3.19247e-04*lvhp_bodyeffect*lvhp_bodyeffect+-4.81987e-04*lvhp_bodyeffect+-1.12400e-02'
+ sky130_fd_pr__pfet_01v8_hvt__k2_diff_15 = '2.42638e-04*lvhp_bodyeffect*lvhp_bodyeffect+-2.35730e-03*lvhp_bodyeffect+-1.33930e-02'
+ sky130_fd_pr__pfet_01v8_hvt__k2_diff_16 = '-2.71381e-04*lvhp_bodyeffect*lvhp_bodyeffect+-1.76525e-04*lvhp_bodyeffect+6.46190e-03'
+ sky130_fd_pr__pfet_01v8_hvt__k2_diff_17 = '-2.00766e-04*lvhp_bodyeffect*lvhp_bodyeffect+1.41238e-04*lvhp_bodyeffect+-3.10580e-03'
+ sky130_fd_pr__pfet_01v8_hvt__k2_diff_18 = '2.19063e-05*lvhp_bodyeffect*lvhp_bodyeffect+1.31625e-04*lvhp_bodyeffect+-1.17230e-02'
+ sky130_fd_pr__pfet_01v8_hvt__k2_diff_19 = '2.24019e-04*lvhp_bodyeffect*lvhp_bodyeffect+9.98178e-04*lvhp_bodyeffect+-7.79110e-03'
+ sky130_fd_pr__pfet_01v8_hvt__k2_diff_2 = '-5.82719e-05*lvhp_bodyeffect*lvhp_bodyeffect+-8.95213e-04*lvhp_bodyeffect+-5.70080e-03'
+ sky130_fd_pr__pfet_01v8_hvt__k2_diff_20 = '2.34578e-04*lvhp_bodyeffect*lvhp_bodyeffect+1.09586e-03*lvhp_bodyeffect+-7.10710e-03'
+ sky130_fd_pr__pfet_01v8_hvt__k2_diff_21 = '1.69347e-04*lvhp_bodyeffect*lvhp_bodyeffect+1.23609e-03*lvhp_bodyeffect+-4.46030e-03'
+ sky130_fd_pr__pfet_01v8_hvt__k2_diff_22 = '3.38917e-04*lvhp_bodyeffect*lvhp_bodyeffect+-1.66342e-03*lvhp_bodyeffect+-1.16240e-02'
+ sky130_fd_pr__pfet_01v8_hvt__k2_diff_23 = '3.67694e-04*lvhp_bodyeffect*lvhp_bodyeffect+-2.27965e-03*lvhp_bodyeffect+-7.38350e-03'
+ sky130_fd_pr__pfet_01v8_hvt__k2_diff_24 = '1.00869e-04*lvhp_bodyeffect*lvhp_bodyeffect+-1.18198e-03*lvhp_bodyeffect+-4.53080e-03'
+ sky130_fd_pr__pfet_01v8_hvt__k2_diff_25 = '7.57969e-05*lvhp_bodyeffect*lvhp_bodyeffect+-1.66375e-05*lvhp_bodyeffect+-9.90050e-03'
+ sky130_fd_pr__pfet_01v8_hvt__k2_diff_26 = '1.35334e-04*lvhp_bodyeffect*lvhp_bodyeffect+5.71537e-04*lvhp_bodyeffect+-9.50460e-03'
+ sky130_fd_pr__pfet_01v8_hvt__k2_diff_27 = '2.77000e-04*lvhp_bodyeffect*lvhp_bodyeffect+1.80950e-03*lvhp_bodyeffect+-7.63600e-03'
+ sky130_fd_pr__pfet_01v8_hvt__k2_diff_28 = '2.48450e-04*lvhp_bodyeffect*lvhp_bodyeffect+1.31272e-03*lvhp_bodyeffect+-5.36360e-03'
+ sky130_fd_pr__pfet_01v8_hvt__k2_diff_29 = '1.14552e-04*lvhp_bodyeffect*lvhp_bodyeffect+9.96835e-04*lvhp_bodyeffect+-8.85950e-03'
+ sky130_fd_pr__pfet_01v8_hvt__k2_diff_3 = '3.61563e-06*lvhp_bodyeffect*lvhp_bodyeffect+-5.52113e-04*lvhp_bodyeffect+-8.56140e-03'
+ sky130_fd_pr__pfet_01v8_hvt__k2_diff_30 = '4.08031e-04*lvhp_bodyeffect*lvhp_bodyeffect+-9.80625e-04*lvhp_bodyeffect+-2.97490e-02'
+ sky130_fd_pr__pfet_01v8_hvt__k2_diff_31 = '2.67191e-04*lvhp_bodyeffect*lvhp_bodyeffect+-2.14026e-03*lvhp_bodyeffect+-1.12810e-02'
+ sky130_fd_pr__pfet_01v8_hvt__k2_diff_32 = '1.88350e-04*lvhp_bodyeffect*lvhp_bodyeffect+2.98711e-05*lvhp_bodyeffect+-2.81170e-03'
+ sky130_fd_pr__pfet_01v8_hvt__k2_diff_33 = '9.97125e-05*lvhp_bodyeffect*lvhp_bodyeffect+1.47575e-04*lvhp_bodyeffect+-1.01710e-02'
+ sky130_fd_pr__pfet_01v8_hvt__k2_diff_34 = '4.71356e-04*lvhp_bodyeffect*lvhp_bodyeffect+4.04487e-03*lvhp_bodyeffect+-3.13120e-03'
+ sky130_fd_pr__pfet_01v8_hvt__k2_diff_35 = '3.64844e-04*lvhp_bodyeffect*lvhp_bodyeffect+3.39238e-03*lvhp_bodyeffect+-9.36100e-03'
+ sky130_fd_pr__pfet_01v8_hvt__k2_diff_36 = '-5.62906e-04*lvhp_bodyeffect*lvhp_bodyeffect+4.05725e-03*lvhp_bodyeffect+6.93850e-03'
+ sky130_fd_pr__pfet_01v8_hvt__k2_diff_37 = '-3.74588e-05*lvhp_bodyeffect*lvhp_bodyeffect+1.46861e-03*lvhp_bodyeffect+-5.57420e-03'
+ sky130_fd_pr__pfet_01v8_hvt__k2_diff_38 = '-5.46688e-04*lvhp_bodyeffect*lvhp_bodyeffect+1.43933e-03*lvhp_bodyeffect+-1.96470e-03'
+ sky130_fd_pr__pfet_01v8_hvt__k2_diff_39 = '8.61444e-04*lvhp_bodyeffect*lvhp_bodyeffect+2.29383e-03*lvhp_bodyeffect+-6.40940e-03'
+ sky130_fd_pr__pfet_01v8_hvt__k2_diff_4 = '-6.44375e-06*lvhp_bodyeffect*lvhp_bodyeffect+-2.80425e-04*lvhp_bodyeffect+-9.81320e-03'
+ sky130_fd_pr__pfet_01v8_hvt__k2_diff_40 = '1.59434e-04*lvhp_bodyeffect*lvhp_bodyeffect+8.99188e-04*lvhp_bodyeffect+-7.55350e-03'
+ sky130_fd_pr__pfet_01v8_hvt__k2_diff_41 = '-1.31250e-05*lvhp_bodyeffect*lvhp_bodyeffect+3.12950e-03*lvhp_bodyeffect+-1.09910e-02'
+ sky130_fd_pr__pfet_01v8_hvt__k2_diff_42 = '-1.18281e-04*lvhp_bodyeffect*lvhp_bodyeffect+5.77625e-04*lvhp_bodyeffect+-1.06030e-02'
+ sky130_fd_pr__pfet_01v8_hvt__k2_diff_43 = '-7.93813e-05*lvhp_bodyeffect*lvhp_bodyeffect+5.20400e-04*lvhp_bodyeffect+-2.83990e-03'
+ sky130_fd_pr__pfet_01v8_hvt__k2_diff_44 = '-3.09469e-05*lvhp_bodyeffect*lvhp_bodyeffect+6.34287e-04*lvhp_bodyeffect+-4.82610e-03'
+ sky130_fd_pr__pfet_01v8_hvt__k2_diff_45 = '-5.22070e-04*lvhp_bodyeffect*lvhp_bodyeffect+2.52737e-04*lvhp_bodyeffect+5.31470e-04'
+ sky130_fd_pr__pfet_01v8_hvt__k2_diff_46 = '1.85447e-03*lvhp_bodyeffect*lvhp_bodyeffect+4.65087e-03*lvhp_bodyeffect+-2.75100e-02'
+ sky130_fd_pr__pfet_01v8_hvt__k2_diff_47 = '-7.33750e-06*lvhp_bodyeffect*lvhp_bodyeffect+1.33058e-03*lvhp_bodyeffect+-2.65490e-03'
+ sky130_fd_pr__pfet_01v8_hvt__k2_diff_48 = '6.36075e-04*lvhp_bodyeffect*lvhp_bodyeffect+2.27887e-03*lvhp_bodyeffect+-8.41570e-03'
+ sky130_fd_pr__pfet_01v8_hvt__k2_diff_49 = '-1.69538e-04*lvhp_bodyeffect*lvhp_bodyeffect+-1.50460e-03*lvhp_bodyeffect+-1.01900e-02'
+ sky130_fd_pr__pfet_01v8_hvt__k2_diff_5 = '-2.60625e-05*lvhp_bodyeffect*lvhp_bodyeffect+-2.32500e-04*lvhp_bodyeffect+-1.08150e-02'
+ sky130_fd_pr__pfet_01v8_hvt__k2_diff_50 = '6.36075e-04*lvhp_bodyeffect*lvhp_bodyeffect+2.27888e-03*lvhp_bodyeffect'
+ sky130_fd_pr__pfet_01v8_hvt__k2_diff_51 = '3.19246e-04*lvhp_bodyeffect*lvhp_bodyeffect+-4.81988e-04*lvhp_bodyeffect'
+ sky130_fd_pr__pfet_01v8_hvt__k2_diff_52 = '4.94343e-04*lvhp_bodyeffect*lvhp_bodyeffect+-1.12813e-03*lvhp_bodyeffect'
+ sky130_fd_pr__pfet_01v8_hvt__k2_diff_53 = '4.38052e-04*lvhp_bodyeffect*lvhp_bodyeffect+-6.01211e-04*lvhp_bodyeffect'
+ sky130_fd_pr__pfet_01v8_hvt__k2_diff_54 = '-1.69536e-04*lvhp_bodyeffect*lvhp_bodyeffect+-1.50460e-03*lvhp_bodyeffect'
+ sky130_fd_pr__pfet_01v8_hvt__k2_diff_55 = '2.42638e-04*lvhp_bodyeffect*lvhp_bodyeffect+-2.35730e-03*lvhp_bodyeffect'
+ sky130_fd_pr__pfet_01v8_hvt__k2_diff_56 = '2.11381e-04*lvhp_bodyeffect*lvhp_bodyeffect+-2.72927e-03*lvhp_bodyeffect+-2.09340e-02'
+ sky130_fd_pr__pfet_01v8_hvt__k2_diff_57 = '3.10831e-04*lvhp_bodyeffect*lvhp_bodyeffect+-3.70433e-03*lvhp_bodyeffect+-1.43480e-02'
+ sky130_fd_pr__pfet_01v8_hvt__k2_diff_58 = '3.68653e-04*lvhp_bodyeffect*lvhp_bodyeffect+-3.76611e-03*lvhp_bodyeffect+-1.58010e-02'
+ sky130_fd_pr__pfet_01v8_hvt__k2_diff_59 = '-8.37813e-05*lvhp_bodyeffect*lvhp_bodyeffect+-2.53462e-03*lvhp_bodyeffect+-1.44450e-02'
+ sky130_fd_pr__pfet_01v8_hvt__k2_diff_6 = '4.94344e-04*lvhp_bodyeffect*lvhp_bodyeffect+-1.12812e-03*lvhp_bodyeffect+-2.54630e-02'
+ sky130_fd_pr__pfet_01v8_hvt__k2_diff_60 = '-1.55828e-04*lvhp_bodyeffect*lvhp_bodyeffect+-2.87994e-03*lvhp_bodyeffect+-1.37850e-02'
+ sky130_fd_pr__pfet_01v8_hvt__k2_diff_61 = '-1.72534e-04*lvhp_bodyeffect*lvhp_bodyeffect+-2.89261e-03*lvhp_bodyeffect+-1.33080e-02'
+ sky130_fd_pr__pfet_01v8_hvt__k2_diff_62 = '-1.84084e-04*lvhp_bodyeffect*lvhp_bodyeffect+-2.99191e-03*lvhp_bodyeffect+-1.19490e-02'
+ sky130_fd_pr__pfet_01v8_hvt__k2_diff_63 = '-3.03994e-04*lvhp_bodyeffect*lvhp_bodyeffect+-2.20625e-04*lvhp_bodyeffect+-9.89160e-03'
+ sky130_fd_pr__pfet_01v8_hvt__k2_diff_64 = '-4.51906e-05*lvhp_bodyeffect*lvhp_bodyeffect+-3.14531e-03*lvhp_bodyeffect+-6.88970e-03'
+ sky130_fd_pr__pfet_01v8_hvt__k2_diff_65 = '1.60712e-04*lvhp_bodyeffect*lvhp_bodyeffect+-7.81975e-04*lvhp_bodyeffect+-7.30460e-03'
+ sky130_fd_pr__pfet_01v8_hvt__k2_diff_66 = '-9.93313e-05*lvhp_bodyeffect*lvhp_bodyeffect+-2.92992e-03*lvhp_bodyeffect+-1.25630e-02'
+ sky130_fd_pr__pfet_01v8_hvt__k2_diff_67 = '1.85362e-04*lvhp_bodyeffect*lvhp_bodyeffect+-2.14045e-03*lvhp_bodyeffect+-1.27900e-02'
+ sky130_fd_pr__pfet_01v8_hvt__k2_diff_7 = '4.31653e-04*lvhp_bodyeffect*lvhp_bodyeffect+-2.29881e-03*lvhp_bodyeffect+-2.91970e-03'
+ sky130_fd_pr__pfet_01v8_hvt__k2_diff_8 = '5.64844e-05*lvhp_bodyeffect*lvhp_bodyeffect+-2.72324e-03*lvhp_bodyeffect+-5.28680e-03'
+ sky130_fd_pr__pfet_01v8_hvt__k2_diff_9 = '3.47809e-04*lvhp_bodyeffect*lvhp_bodyeffect+2.05949e-03*lvhp_bodyeffect+-9.60400e-03'
+ sky130_fd_pr__pfet_01v8_hvt__keta_diff_52 = '4.61422e-09*lvhp_bodyeffect*lvhp_bodyeffect+3.76186e-08*lvhp_bodyeffect'
+ sky130_fd_pr__pfet_01v8_hvt__keta_diff_59 = '4.62369e-07*lvhp_bodyeffect*lvhp_bodyeffect+1.95804e-05*lvhp_bodyeffect'
+ sky130_fd_pr__pfet_01v8_hvt__keta_diff_60 = '4.40106e-07*lvhp_bodyeffect*lvhp_bodyeffect+2.00053e-05*lvhp_bodyeffect'
+ sky130_fd_pr__pfet_01v8_hvt__keta_diff_61 = '2.83956e-07*lvhp_bodyeffect*lvhp_bodyeffect+1.36136e-05*lvhp_bodyeffect'
+ sky130_fd_pr__pfet_01v8_hvt__keta_diff_62 = '1.21494e-07*lvhp_bodyeffect*lvhp_bodyeffect+6.05125e-06*lvhp_bodyeffect'
+ sky130_fd_pr__pfet_01v8_hvt__keta_diff_63 = '1.21478e-07*lvhp_bodyeffect*lvhp_bodyeffect+6.05124e-06*lvhp_bodyeffect'
+ sky130_fd_pr__pfet_01v8_hvt__keta_diff_64 = '-1.89178e-07*lvhp_bodyeffect*lvhp_bodyeffect+-9.42226e-06*lvhp_bodyeffect'
+ sky130_fd_pr__pfet_01v8_hvt__keta_diff_66 = '-9.84500e-09*lvhp_bodyeffect*lvhp_bodyeffect+-5.18847e-07*lvhp_bodyeffect'
+ sky130_fd_pr__pfet_01v8_hvt__keta_diff_67 = '-1.61016e-08*lvhp_bodyeffect*lvhp_bodyeffect+-9.26179e-07*lvhp_bodyeffect'
+ sky130_fd_pr__pfet_01v8_hvt__kt1_diff_59 = '1.74906e-06*lvp_subvt*lvp_subvt+7.40612e-05*lvp_subvt'
+ sky130_fd_pr__pfet_01v8_hvt__kt1_diff_60 = '1.66469e-06*lvp_subvt*lvp_subvt+7.56687e-05*lvp_subvt'
+ sky130_fd_pr__pfet_01v8_hvt__kt1_diff_61 = '1.07406e-06*lvp_subvt*lvp_subvt+5.14913e-05*lvp_subvt'
+ sky130_fd_pr__pfet_01v8_hvt__kt1_diff_62 = '4.59538e-07*lvp_subvt*lvp_subvt+2.28883e-05*lvp_subvt'
+ sky130_fd_pr__pfet_01v8_hvt__kt1_diff_63 = '4.59541e-07*lvp_subvt*lvp_subvt+2.28883e-05*lvp_subvt'
+ sky130_fd_pr__pfet_01v8_hvt__kt1_diff_64 = '6.31562e-07*lvp_subvt*lvp_subvt+3.14512e-05*lvp_subvt'
+ sky130_fd_pr__pfet_01v8_hvt__kt1_diff_67 = '-3.74159e-07*lvp_subvt*lvp_subvt+-2.14284e-05*lvp_subvt'
+ sky130_fd_pr__pfet_01v8_hvt__lint_diff = '-4.33125e-09*poly_cd'
+ sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_0 = '2.60594e-03*lvp_subvt*lvp_subvt+-3.22204e-01*lvp_subvt+3.39690e-01'
+ sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_1 = '1.02134e-02*lvp_subvt*lvp_subvt+-2.37229e-01*lvp_subvt+6.08570e-01'
+ sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_10 = '-1.45492e-03*lvp_subvt*lvp_subvt+-3.09847e-02*lvp_subvt+1.49740e-01'
+ sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_11 = '-1.80097e-02*lvp_subvt*lvp_subvt+2.67764e-02*lvp_subvt+2.17550e-01'
+ sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_12 = '-3.50584e-02*lvp_subvt*lvp_subvt+9.16337e-02*lvp_subvt+1.19940e+00'
+ sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_13 = '-6.58228e-02*lvp_subvt*lvp_subvt+-2.25763e-02*lvp_subvt+1.23430e+00'
+ sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_14 = '1.50991e-02*lvp_subvt*lvp_subvt+-1.81374e-01*lvp_subvt+2.87420e-01'
+ sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_15 = '2.43281e-02*lvp_subvt*lvp_subvt+-3.65175e-02*lvp_subvt+1.26140e-01'
+ sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_16 = '1.73452e-02*lvp_subvt*lvp_subvt+-7.62594e-02*lvp_subvt+1.24570e-01'
+ sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_17 = '-7.65722e-02*lvp_subvt*lvp_subvt+-1.17771e-01*lvp_subvt+1.28230e+00'
+ sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_18 = '5.70878e-03*lvp_subvt*lvp_subvt+-3.11466e-02*lvp_subvt+6.65630e-02'
+ sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_19 = '-6.58649e-03*lvp_subvt*lvp_subvt+-1.70085e-02*lvp_subvt+1.64730e-01'
+ sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_2 = '1.13113e-02*lvp_subvt*lvp_subvt+-1.25043e-01*lvp_subvt+2.08020e-01'
+ sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_20 = '-6.35269e-03*lvp_subvt*lvp_subvt+-3.84983e-02*lvp_subvt+2.15100e-01'
+ sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_21 = '3.75222e-02*lvp_subvt*lvp_subvt+-3.20987e-02*lvp_subvt+-3.63210e-01'
+ sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_22 = '7.40656e-03*lvp_subvt*lvp_subvt+-1.82554e-01*lvp_subvt+2.33980e-01'
+ sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_23 = '-2.13056e-02*lvp_subvt*lvp_subvt+-1.17538e-01*lvp_subvt+5.86980e-01'
+ sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_24 = '3.09694e-03*lvp_subvt*lvp_subvt+-4.70227e-02*lvp_subvt+7.76780e-02'
+ sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_25 = '5.07625e-03*lvp_subvt*lvp_subvt+-1.34547e-01*lvp_subvt+-3.30530e-01'
+ sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_26 = '4.04004e-03*lvp_subvt*lvp_subvt+-1.26998e-02*lvp_subvt+-3.29570e-04'
+ sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_27 = '-8.99309e-03*lvp_subvt*lvp_subvt+-7.33487e-03*lvp_subvt+8.90970e-02'
+ sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_28 = '-8.75597e-02*lvp_subvt*lvp_subvt+-1.37994e-01*lvp_subvt+1.21660e+00'
+ sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_29 = '-3.40856e-02*lvp_subvt*lvp_subvt+-7.56125e-02*lvp_subvt+1.21870e+00'
+ sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_3 = '-7.93688e-04*lvp_subvt*lvp_subvt+-7.26897e-02*lvp_subvt+2.87260e-01'
+ sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_30 = '9.91969e-04*lvp_subvt*lvp_subvt+-1.36027e-01*lvp_subvt+6.14820e-01'
+ sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_31 = '4.66881e-03*lvp_subvt*lvp_subvt+-6.25797e-02*lvp_subvt+1.00050e-01'
+ sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_32 = '2.03109e-03*lvp_subvt*lvp_subvt+-5.03581e-02*lvp_subvt+1.23660e-01'
+ sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_33 = '-9.39834e-02*lvp_subvt*lvp_subvt+-2.96341e-01*lvp_subvt+1.28910e+00'
+ sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_34 = '-8.68375e-02*lvp_subvt*lvp_subvt+-2.74275e-01*lvp_subvt+1.38700e+00'
+ sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_35 = '-1.10131e-03*lvp_subvt*lvp_subvt+-7.18003e-02*lvp_subvt+2.29530e-01'
+ sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_36 = '-4.53853e-02*lvp_subvt*lvp_subvt+-4.60262e-02*lvp_subvt+1.23810e+00'
+ sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_37 = '1.54769e-02*lvp_subvt*lvp_subvt+-6.82175e-02*lvp_subvt+2.29120e-01'
+ sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_38 = '-5.30781e-02*lvp_subvt*lvp_subvt+-3.60375e-02*lvp_subvt+1.24230e+00'
+ sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_39 = '4.10688e-03*lvp_subvt*lvp_subvt+-3.36020e-01*lvp_subvt+8.68910e-01'
+ sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_4 = '7.64000e-04*lvp_subvt*lvp_subvt+-3.60790e-02*lvp_subvt+2.13960e-01'
+ sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_40 = '8.91687e-02*lvp_subvt*lvp_subvt+-1.19711e-01*lvp_subvt+4.65560e-02'
+ sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_41 = '-7.28094e-02*lvp_subvt*lvp_subvt+-3.49638e-01*lvp_subvt+1.41090e+00'
+ sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_42 = '2.68237e-02*lvp_subvt*lvp_subvt+-1.47690e-01*lvp_subvt+2.97460e-01'
+ sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_43 = '1.27791e-02*lvp_subvt*lvp_subvt+-6.44337e-02*lvp_subvt+2.71930e-01'
+ sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_44 = '4.91750e-03*lvp_subvt*lvp_subvt+-2.99775e-02*lvp_subvt+2.93010e-01'
+ sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_45 = '8.87159e-03*lvp_subvt*lvp_subvt+-3.28019e-02*lvp_subvt+8.89470e-02'
+ sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_46 = '2.35089e-02*lvp_subvt*lvp_subvt+-2.60637e-01*lvp_subvt+6.70210e-01'
+ sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_47 = '-1.38500e-02*lvp_subvt*lvp_subvt+-6.27650e-01*lvp_subvt+1.39920e+00'
+ sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_48 = '1.30237e-02*lvp_subvt*lvp_subvt+-3.77937e-01*lvp_subvt+8.06070e-01'
+ sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_49 = '-3.12539e-02*lvp_subvt*lvp_subvt+-2.24216e-01*lvp_subvt+1.41450e+00'
+ sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_5 = '4.52047e-03*lvp_subvt*lvp_subvt+-6.38931e-02*lvp_subvt+2.61110e-01'
+ sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_50 = '1.30238e-02*lvp_subvt*lvp_subvt+-3.77938e-01*lvp_subvt'
+ sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_51 = '1.50991e-02*lvp_subvt*lvp_subvt+-1.81374e-01*lvp_subvt'
+ sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_52 = '2.17517e-03*lvp_subvt*lvp_subvt+-2.95474e-01*lvp_subvt'
+ sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_53 = '1.02134e-02*lvp_subvt*lvp_subvt+-2.37229e-01*lvp_subvt'
+ sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_54 = '-3.12539e-02*lvp_subvt*lvp_subvt+-2.24216e-01*lvp_subvt'
+ sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_55 = '2.43281e-02*lvp_subvt*lvp_subvt+-3.65175e-02*lvp_subvt'
+ sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_59 = '-2.75228e-03*lvp_subvt*lvp_subvt+-3.21786e-01*lvp_subvt'
+ sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_6 = '2.17522e-03*lvp_subvt*lvp_subvt+-2.95474e-01*lvp_subvt+1.13110e+00'
+ sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_60 = '-1.40848e-02*lvp_subvt*lvp_subvt+-2.82421e-01*lvp_subvt'
+ sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_61 = '-2.21735e-02*lvp_subvt*lvp_subvt+-2.54791e-01*lvp_subvt'
+ sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_62 = '-2.77481e-02*lvp_subvt*lvp_subvt+-2.35966e-01*lvp_subvt'
+ sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_63 = '-2.77481e-02*lvp_subvt*lvp_subvt+-2.35966e-01*lvp_subvt'
+ sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_64 = '-7.29347e-03*lvp_subvt*lvp_subvt+-2.31757e-01*lvp_subvt'
+ sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_66 = '-2.64125e-02*lvp_subvt*lvp_subvt+-2.34828e-01*lvp_subvt'
+ sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_67 = '-9.05755e-03*lvp_subvt*lvp_subvt+-2.72049e-01*lvp_subvt'
+ sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_7 = '4.33035e-02*lvp_subvt*lvp_subvt+-1.26533e-01*lvp_subvt+-1.32090e-01'
+ sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_8 = '-9.07781e-03*lvp_subvt*lvp_subvt+-2.19426e-01*lvp_subvt+5.65240e-01'
+ sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_9 = '-4.07313e-03*lvp_subvt*lvp_subvt+-3.57825e-01*lvp_subvt+1.12170e-01'
+ sky130_fd_pr__pfet_01v8_hvt__overlap_mult = '4.16563e-03*lvtox*lvtox+3.61700e-02*lvtox+9.88670e-01'
+ sky130_fd_pr__pfet_01v8_hvt__pjunction_mult = '-6.25000e-07*lvp_diode*lvp_diode+2.44275e-02*lvp_diode+1.02860e+00'
+ sky130_fd_pr__pfet_01v8_hvt__toxe_mult = '1.30000e-02*lvtox+1.00000e+00'
+ sky130_fd_pr__pfet_01v8_hvt__u0_diff_0 = '3.31306e-06*lvhp_mobility*lvhp_mobility+-1.12818e-04*lvhp_mobility+3.60800e-04'
+ sky130_fd_pr__pfet_01v8_hvt__u0_diff_1 = '-1.89697e-05*lvhp_mobility*lvhp_mobility+5.39563e-05*lvhp_mobility+1.06740e-03'
+ sky130_fd_pr__pfet_01v8_hvt__u0_diff_10 = '1.89670e-05*lvhp_mobility*lvhp_mobility+-2.87502e-04*lvhp_mobility+8.78420e-04'
+ sky130_fd_pr__pfet_01v8_hvt__u0_diff_11 = '8.76474e-05*lvhp_mobility*lvhp_mobility+-4.49975e-04*lvhp_mobility+2.99040e-04'
+ sky130_fd_pr__pfet_01v8_hvt__u0_diff_12 = '1.26353e-04*lvhp_mobility*lvhp_mobility+-4.74234e-04*lvhp_mobility+2.54520e-04'
+ sky130_fd_pr__pfet_01v8_hvt__u0_diff_13 = '1.50375e-04*lvhp_mobility*lvhp_mobility+-5.76068e-04*lvhp_mobility+1.22430e-04'
+ sky130_fd_pr__pfet_01v8_hvt__u0_diff_14 = '1.26931e-05*lvhp_mobility*lvhp_mobility+4.31200e-05*lvhp_mobility+3.87300e-04'
+ sky130_fd_pr__pfet_01v8_hvt__u0_diff_15 = '2.64753e-05*lvhp_mobility*lvhp_mobility+1.55888e-05*lvhp_mobility+5.32540e-04'
+ sky130_fd_pr__pfet_01v8_hvt__u0_diff_16 = '2.29216e-05*lvhp_mobility*lvhp_mobility+-1.27579e-04*lvhp_mobility+3.48540e-04'
+ sky130_fd_pr__pfet_01v8_hvt__u0_diff_17 = '5.67106e-05*lvhp_mobility*lvhp_mobility+-3.89200e-04*lvhp_mobility+1.55630e-04'
+ sky130_fd_pr__pfet_01v8_hvt__u0_diff_18 = '-1.32021e-05*lvhp_mobility*lvhp_mobility+-2.90758e-04*lvhp_mobility+1.36610e-03'
+ sky130_fd_pr__pfet_01v8_hvt__u0_diff_19 = '1.12822e-05*lvhp_mobility*lvhp_mobility+-4.29821e-04*lvhp_mobility+1.21890e-03'
+ sky130_fd_pr__pfet_01v8_hvt__u0_diff_2 = '7.85844e-05*lvhp_mobility*lvhp_mobility+1.54413e-04*lvhp_mobility+1.53290e-03'
+ sky130_fd_pr__pfet_01v8_hvt__u0_diff_20 = '2.51739e-05*lvhp_mobility*lvhp_mobility+-5.80154e-04*lvhp_mobility+1.91420e-03'
+ sky130_fd_pr__pfet_01v8_hvt__u0_diff_21 = '1.64298e-04*lvhp_mobility*lvhp_mobility+-6.11334e-04*lvhp_mobility+-1.08380e-03'
+ sky130_fd_pr__pfet_01v8_hvt__u0_diff_22 = '1.61613e-05*lvhp_mobility*lvhp_mobility+4.41725e-05*lvhp_mobility+3.45800e-04'
+ sky130_fd_pr__pfet_01v8_hvt__u0_diff_23 = '-2.56553e-05*lvhp_mobility*lvhp_mobility+1.71250e-07*lvhp_mobility+1.07310e-03'
+ sky130_fd_pr__pfet_01v8_hvt__u0_diff_24 = '5.93125e-07*lvhp_mobility*lvhp_mobility+-1.26395e-04*lvhp_mobility+3.33250e-04'
+ sky130_fd_pr__pfet_01v8_hvt__u0_diff_25 = '-5.51231e-05*lvhp_mobility*lvhp_mobility+-3.07889e-04*lvhp_mobility+-1.58760e-05'
+ sky130_fd_pr__pfet_01v8_hvt__u0_diff_26 = '-2.61072e-05*lvhp_mobility*lvhp_mobility+-4.71204e-04*lvhp_mobility+1.84710e-03'
+ sky130_fd_pr__pfet_01v8_hvt__u0_diff_27 = '1.55484e-05*lvhp_mobility*lvhp_mobility+-6.10406e-04*lvhp_mobility+1.82160e-03'
+ sky130_fd_pr__pfet_01v8_hvt__u0_diff_28 = '4.99387e-05*lvhp_mobility*lvhp_mobility+-6.85795e-04*lvhp_mobility+1.43520e-03'
+ sky130_fd_pr__pfet_01v8_hvt__u0_diff_29 = '1.94228e-04*lvhp_mobility*lvhp_mobility+-1.09454e-03*lvhp_mobility+1.74190e-03'
+ sky130_fd_pr__pfet_01v8_hvt__u0_diff_3 = '4.72187e-06*lvhp_mobility*lvhp_mobility+-1.22313e-04*lvhp_mobility+1.45490e-03'
+ sky130_fd_pr__pfet_01v8_hvt__u0_diff_30 = '-4.43344e-06*lvhp_mobility*lvhp_mobility+7.99837e-05*lvhp_mobility+1.22990e-03'
+ sky130_fd_pr__pfet_01v8_hvt__u0_diff_31 = '1.09972e-05*lvhp_mobility*lvhp_mobility+1.61788e-05*lvhp_mobility+1.35140e-04'
+ sky130_fd_pr__pfet_01v8_hvt__u0_diff_32 = '1.23973e-05*lvhp_mobility*lvhp_mobility+-8.00756e-05*lvhp_mobility+1.67790e-04'
+ sky130_fd_pr__pfet_01v8_hvt__u0_diff_33 = '-2.50956e-05*lvhp_mobility*lvhp_mobility+-3.65983e-04*lvhp_mobility+1.08990e-03'
+ sky130_fd_pr__pfet_01v8_hvt__u0_diff_34 = '7.90934e-05*lvhp_mobility*lvhp_mobility+-5.60176e-04*lvhp_mobility+1.49660e-03'
+ sky130_fd_pr__pfet_01v8_hvt__u0_diff_35 = '1.27188e-07*lvhp_mobility*lvhp_mobility+-3.29566e-04*lvhp_mobility+2.13070e-03'
+ sky130_fd_pr__pfet_01v8_hvt__u0_diff_36 = '2.47470e-04*lvhp_mobility*lvhp_mobility+-6.16917e-04*lvhp_mobility+-2.13990e-04'
+ sky130_fd_pr__pfet_01v8_hvt__u0_diff_37 = '1.15325e-04*lvhp_mobility*lvhp_mobility+1.80550e-04*lvhp_mobility+2.02120e-03'
+ sky130_fd_pr__pfet_01v8_hvt__u0_diff_38 = '2.74406e-04*lvhp_mobility*lvhp_mobility+-2.24962e-04*lvhp_mobility+7.52060e-04'
+ sky130_fd_pr__pfet_01v8_hvt__u0_diff_39 = '5.08148e-05*lvhp_mobility*lvhp_mobility+-3.16581e-04*lvhp_mobility+4.65540e-04'
+ sky130_fd_pr__pfet_01v8_hvt__u0_diff_4 = '1.12281e-05*lvhp_mobility*lvhp_mobility+-5.51625e-05*lvhp_mobility+1.22350e-03'
+ sky130_fd_pr__pfet_01v8_hvt__u0_diff_40 = '8.55806e-05*lvhp_mobility*lvhp_mobility+-4.48575e-04*lvhp_mobility+-9.82290e-04'
+ sky130_fd_pr__pfet_01v8_hvt__u0_diff_41 = '1.30416e-04*lvhp_mobility*lvhp_mobility+-7.12706e-04*lvhp_mobility+7.74820e-04'
+ sky130_fd_pr__pfet_01v8_hvt__u0_diff_42 = '8.86281e-05*lvhp_mobility*lvhp_mobility+-2.92513e-04*lvhp_mobility+2.11190e-03'
+ sky130_fd_pr__pfet_01v8_hvt__u0_diff_43 = '8.82438e-05*lvhp_mobility*lvhp_mobility+-1.43925e-04*lvhp_mobility+1.30840e-03'
+ sky130_fd_pr__pfet_01v8_hvt__u0_diff_44 = '3.22781e-05*lvhp_mobility*lvhp_mobility+-1.95625e-05*lvhp_mobility+1.86790e-03'
+ sky130_fd_pr__pfet_01v8_hvt__u0_diff_45 = '1.24147e-04*lvhp_mobility*lvhp_mobility+2.26250e-05*lvhp_mobility+5.58520e-05'
+ sky130_fd_pr__pfet_01v8_hvt__u0_diff_46 = '-2.81225e-05*lvhp_mobility*lvhp_mobility+-1.76157e-04*lvhp_mobility+7.12120e-04'
+ sky130_fd_pr__pfet_01v8_hvt__u0_diff_47 = '4.17675e-04*lvhp_mobility*lvhp_mobility+-2.00504e-03*lvhp_mobility+9.28030e-04'
+ sky130_fd_pr__pfet_01v8_hvt__u0_diff_48 = '5.37374e-05*lvhp_mobility*lvhp_mobility+-9.74113e-05*lvhp_mobility+-3.19430e-05'
+ sky130_fd_pr__pfet_01v8_hvt__u0_diff_49 = '1.57980e-04*lvhp_mobility*lvhp_mobility+2.31375e-04*lvhp_mobility+1.92820e-04'
+ sky130_fd_pr__pfet_01v8_hvt__u0_diff_5 = '2.70688e-05*lvhp_mobility*lvhp_mobility+-2.94250e-05*lvhp_mobility+1.55300e-03'
+ sky130_fd_pr__pfet_01v8_hvt__u0_diff_50 = '5.37372e-05*lvhp_mobility*lvhp_mobility+-9.74112e-05*lvhp_mobility'
+ sky130_fd_pr__pfet_01v8_hvt__u0_diff_51 = '1.26931e-05*lvhp_mobility*lvhp_mobility+4.31200e-05*lvhp_mobility'
+ sky130_fd_pr__pfet_01v8_hvt__u0_diff_52 = '-1.43562e-05*lvhp_mobility*lvhp_mobility+-1.39475e-04*lvhp_mobility'
+ sky130_fd_pr__pfet_01v8_hvt__u0_diff_53 = '-1.89697e-05*lvhp_mobility*lvhp_mobility+5.39563e-05*lvhp_mobility'
+ sky130_fd_pr__pfet_01v8_hvt__u0_diff_54 = '1.57980e-04*lvhp_mobility*lvhp_mobility+2.31375e-04*lvhp_mobility'
+ sky130_fd_pr__pfet_01v8_hvt__u0_diff_55 = '2.64753e-05*lvhp_mobility*lvhp_mobility+1.55887e-05*lvhp_mobility'
+ sky130_fd_pr__pfet_01v8_hvt__u0_diff_56 = '-9.59688e-07*lvhp_mobility*lvhp_mobility+2.08456e-04*lvhp_mobility+-1.75820e-04'
+ sky130_fd_pr__pfet_01v8_hvt__u0_diff_57 = '-8.28725e-06*lvhp_mobility*lvhp_mobility+6.39085e-05*lvhp_mobility+-1.76180e-04'
+ sky130_fd_pr__pfet_01v8_hvt__u0_diff_58 = '-5.31313e-06*lvhp_mobility*lvhp_mobility+5.99425e-05*lvhp_mobility+-2.01890e-04'
+ sky130_fd_pr__pfet_01v8_hvt__u0_diff_59 = '8.58569e-05*lvhp_mobility*lvhp_mobility+-2.60625e-05*lvhp_mobility+-1.63460e-04'
+ sky130_fd_pr__pfet_01v8_hvt__u0_diff_6 = '-1.43562e-05*lvhp_mobility*lvhp_mobility+-1.39475e-04*lvhp_mobility+1.20820e-03'
+ sky130_fd_pr__pfet_01v8_hvt__u0_diff_60 = '1.08603e-04*lvhp_mobility*lvhp_mobility+6.67875e-05*lvhp_mobility+-1.81900e-04'
+ sky130_fd_pr__pfet_01v8_hvt__u0_diff_61 = '1.23424e-04*lvhp_mobility*lvhp_mobility+1.05550e-04*lvhp_mobility+-2.19980e-04'
+ sky130_fd_pr__pfet_01v8_hvt__u0_diff_62 = '1.34194e-04*lvhp_mobility*lvhp_mobility+1.38263e-04*lvhp_mobility+-2.21450e-04'
+ sky130_fd_pr__pfet_01v8_hvt__u0_diff_63 = '1.36827e-04*lvhp_mobility*lvhp_mobility+1.29025e-04*lvhp_mobility+-1.56030e-04'
+ sky130_fd_pr__pfet_01v8_hvt__u0_diff_64 = '6.43731e-05*lvhp_mobility*lvhp_mobility+-3.26512e-04*lvhp_mobility+-1.17220e-04'
+ sky130_fd_pr__pfet_01v8_hvt__u0_diff_65 = '-1.30872e-05*lvhp_mobility*lvhp_mobility+1.65162e-05*lvhp_mobility+-3.14530e-04'
+ sky130_fd_pr__pfet_01v8_hvt__u0_diff_66 = '1.19247e-04*lvhp_mobility*lvhp_mobility+1.05813e-04*lvhp_mobility+-2.41200e-04'
+ sky130_fd_pr__pfet_01v8_hvt__u0_diff_67 = '3.88975e-05*lvhp_mobility*lvhp_mobility+-5.17525e-05*lvhp_mobility+-2.95950e-04'
+ sky130_fd_pr__pfet_01v8_hvt__u0_diff_7 = '4.63056e-05*lvhp_mobility*lvhp_mobility+-2.64050e-04*lvhp_mobility+-7.21490e-04'
+ sky130_fd_pr__pfet_01v8_hvt__u0_diff_8 = '6.11519e-05*lvhp_mobility*lvhp_mobility+-3.35215e-04*lvhp_mobility+-1.85390e-04'
+ sky130_fd_pr__pfet_01v8_hvt__u0_diff_9 = '-3.60937e-06*lvhp_mobility*lvhp_mobility+-7.91962e-04*lvhp_mobility+1.42060e-03'
+ sky130_fd_pr__pfet_01v8_hvt__ua_diff_0 = '3.29139e-12*lvhp_mobility*lvhp_mobility+-2.30284e-11*lvhp_mobility+3.73740e-11'
+ sky130_fd_pr__pfet_01v8_hvt__ua_diff_1 = '-4.94687e-12*lvhp_mobility*lvhp_mobility+1.91250e-11*lvhp_mobility+3.45860e-10'
+ sky130_fd_pr__pfet_01v8_hvt__ua_diff_10 = '-1.02742e-12*lvhp_mobility*lvhp_mobility+1.72948e-11*lvhp_mobility+-5.80820e-11'
+ sky130_fd_pr__pfet_01v8_hvt__ua_diff_11 = '-2.36751e-12*lvhp_mobility*lvhp_mobility+1.69550e-11*lvhp_mobility+-3.41100e-11'
+ sky130_fd_pr__pfet_01v8_hvt__ua_diff_12 = '-4.69559e-12*lvhp_mobility*lvhp_mobility+2.13106e-11*lvhp_mobility+-1.14080e-11'
+ sky130_fd_pr__pfet_01v8_hvt__ua_diff_13 = '-1.03067e-11*lvhp_mobility*lvhp_mobility+4.05101e-11*lvhp_mobility+-1.12320e-11'
+ sky130_fd_pr__pfet_01v8_hvt__ua_diff_14 = '4.87622e-12*lvhp_mobility*lvhp_mobility+5.27563e-12*lvhp_mobility+3.78280e-11'
+ sky130_fd_pr__pfet_01v8_hvt__ua_diff_15 = '1.00166e-11*lvhp_mobility*lvhp_mobility+-4.33750e-12*lvhp_mobility+-1.45650e-11'
+ sky130_fd_pr__pfet_01v8_hvt__ua_diff_16 = '4.20839e-12*lvhp_mobility*lvhp_mobility+-1.42874e-11*lvhp_mobility+5.63620e-12'
+ sky130_fd_pr__pfet_01v8_hvt__ua_diff_17 = '7.40494e-12*lvhp_mobility*lvhp_mobility+-7.92500e-13*lvhp_mobility+-1.10890e-11'
+ sky130_fd_pr__pfet_01v8_hvt__ua_diff_18 = '1.38469e-13*lvhp_mobility*lvhp_mobility+1.72519e-11*lvhp_mobility+-9.67780e-11'
+ sky130_fd_pr__pfet_01v8_hvt__ua_diff_19 = '5.14778e-12*lvhp_mobility*lvhp_mobility+3.37161e-11*lvhp_mobility+-2.01910e-10'
+ sky130_fd_pr__pfet_01v8_hvt__ua_diff_2 = '8.40762e-12*lvhp_mobility*lvhp_mobility+-2.90260e-11*lvhp_mobility+-4.63760e-11'
+ sky130_fd_pr__pfet_01v8_hvt__ua_diff_20 = '1.54639e-12*lvhp_mobility*lvhp_mobility+4.22356e-11*lvhp_mobility+-1.92090e-10'
+ sky130_fd_pr__pfet_01v8_hvt__ua_diff_21 = '2.88022e-11*lvhp_mobility*lvhp_mobility+6.57238e-11*lvhp_mobility+-6.12710e-10'
+ sky130_fd_pr__pfet_01v8_hvt__ua_diff_22 = '5.78644e-12*lvhp_mobility*lvhp_mobility+2.90000e-13*lvhp_mobility+4.09770e-11'
+ sky130_fd_pr__pfet_01v8_hvt__ua_diff_23 = '-5.50786e-12*lvhp_mobility*lvhp_mobility+-1.91489e-11*lvhp_mobility+1.62270e-10'
+ sky130_fd_pr__pfet_01v8_hvt__ua_diff_24 = '2.49187e-12*lvhp_mobility*lvhp_mobility+-2.99122e-12*lvhp_mobility+-5.21200e-11'
+ sky130_fd_pr__pfet_01v8_hvt__ua_diff_25 = '-1.58720e-11*lvhp_mobility*lvhp_mobility+-9.99246e-11*lvhp_mobility+-1.58780e-10'
+ sky130_fd_pr__pfet_01v8_hvt__ua_diff_26 = '6.92000e-13*lvhp_mobility*lvhp_mobility+3.83030e-11*lvhp_mobility+-1.49360e-10'
+ sky130_fd_pr__pfet_01v8_hvt__ua_diff_27 = '1.35156e-12*lvhp_mobility*lvhp_mobility+5.57213e-11*lvhp_mobility+-1.76670e-10'
+ sky130_fd_pr__pfet_01v8_hvt__ua_diff_28 = '-5.60487e-12*lvhp_mobility*lvhp_mobility+7.74625e-11*lvhp_mobility+-1.36720e-11'
+ sky130_fd_pr__pfet_01v8_hvt__ua_diff_29 = '8.77272e-12*lvhp_mobility*lvhp_mobility+4.46921e-11*lvhp_mobility+-1.48520e-11'
+ sky130_fd_pr__pfet_01v8_hvt__ua_diff_3 = '-2.80322e-12*lvhp_mobility*lvhp_mobility+-2.18088e-12*lvhp_mobility+-1.96580e-11'
+ sky130_fd_pr__pfet_01v8_hvt__ua_diff_30 = '-1.34656e-12*lvhp_mobility*lvhp_mobility+2.64625e-12*lvhp_mobility+3.18130e-10'
+ sky130_fd_pr__pfet_01v8_hvt__ua_diff_31 = '3.92984e-12*lvhp_mobility*lvhp_mobility+-1.56194e-11*lvhp_mobility+-1.42250e-10'
+ sky130_fd_pr__pfet_01v8_hvt__ua_diff_32 = '3.06959e-12*lvhp_mobility*lvhp_mobility+8.60625e-13*lvhp_mobility+-1.72430e-11'
+ sky130_fd_pr__pfet_01v8_hvt__ua_diff_33 = '-4.95281e-12*lvhp_mobility*lvhp_mobility+-7.39675e-11*lvhp_mobility+-2.48850e-11'
+ sky130_fd_pr__pfet_01v8_hvt__ua_diff_34 = '5.89781e-12*lvhp_mobility*lvhp_mobility+4.44662e-11*lvhp_mobility+-2.37100e-11'
+ sky130_fd_pr__pfet_01v8_hvt__ua_diff_35 = '-1.45906e-12*lvhp_mobility*lvhp_mobility+7.41875e-12*lvhp_mobility+-1.44560e-10'
+ sky130_fd_pr__pfet_01v8_hvt__ua_diff_36 = '9.11124e-12*lvhp_mobility*lvhp_mobility+1.89052e-11*lvhp_mobility+-9.00080e-12'
+ sky130_fd_pr__pfet_01v8_hvt__ua_diff_37 = '-5.07844e-12*lvhp_mobility*lvhp_mobility+-8.03212e-11*lvhp_mobility+-1.36290e-10'
+ sky130_fd_pr__pfet_01v8_hvt__ua_diff_38 = '1.74837e-11*lvhp_mobility*lvhp_mobility+-1.29782e-10*lvhp_mobility+-2.52700e-11'
+ sky130_fd_pr__pfet_01v8_hvt__ua_diff_39 = '3.25996e-11*lvhp_mobility*lvhp_mobility+1.34875e-12*lvhp_mobility+7.71020e-11'
+ sky130_fd_pr__pfet_01v8_hvt__ua_diff_4 = '-1.15875e-12*lvhp_mobility*lvhp_mobility+-7.55600e-12*lvhp_mobility+-7.28960e-11'
+ sky130_fd_pr__pfet_01v8_hvt__ua_diff_40 = '3.66619e-11*lvhp_mobility*lvhp_mobility+-1.13940e-10*lvhp_mobility+-4.85380e-10'
+ sky130_fd_pr__pfet_01v8_hvt__ua_diff_41 = '2.22794e-11*lvhp_mobility*lvhp_mobility+-2.49113e-11*lvhp_mobility+-2.54850e-11'
+ sky130_fd_pr__pfet_01v8_hvt__ua_diff_42 = '1.20141e-11*lvhp_mobility*lvhp_mobility+-1.05901e-10*lvhp_mobility+1.11790e-10'
+ sky130_fd_pr__pfet_01v8_hvt__ua_diff_43 = '8.18737e-12*lvhp_mobility*lvhp_mobility+-5.25875e-11*lvhp_mobility+-5.50280e-11'
+ sky130_fd_pr__pfet_01v8_hvt__ua_diff_44 = '-2.32738e-12*lvhp_mobility*lvhp_mobility+-1.95260e-11*lvhp_mobility+-8.73180e-11'
+ sky130_fd_pr__pfet_01v8_hvt__ua_diff_45 = '-1.27791e-11*lvhp_mobility*lvhp_mobility+-1.55087e-11*lvhp_mobility+-4.96980e-12'
+ sky130_fd_pr__pfet_01v8_hvt__ua_diff_46 = '-1.03297e-11*lvhp_mobility*lvhp_mobility+-5.72313e-11*lvhp_mobility+1.54490e-10'
+ sky130_fd_pr__pfet_01v8_hvt__ua_diff_47 = '7.07464e-11*lvhp_mobility*lvhp_mobility+-2.16721e-10*lvhp_mobility+1.17270e-12'
+ sky130_fd_pr__pfet_01v8_hvt__ua_diff_48 = '3.43469e-11*lvhp_mobility*lvhp_mobility+5.07125e-11*lvhp_mobility+-8.67210e-11'
+ sky130_fd_pr__pfet_01v8_hvt__ua_diff_49 = '6.11944e-11*lvhp_mobility*lvhp_mobility+1.12381e-10*lvhp_mobility+-7.93530e-12'
+ sky130_fd_pr__pfet_01v8_hvt__ua_diff_5 = '2.23878e-12*lvhp_mobility*lvhp_mobility+-8.49662e-12*lvhp_mobility+-3.48930e-11'
+ sky130_fd_pr__pfet_01v8_hvt__ua_diff_50 = '3.43469e-11*lvhp_mobility*lvhp_mobility+5.07125e-11*lvhp_mobility'
+ sky130_fd_pr__pfet_01v8_hvt__ua_diff_51 = '4.87622e-12*lvhp_mobility*lvhp_mobility+5.27564e-12*lvhp_mobility'
+ sky130_fd_pr__pfet_01v8_hvt__ua_diff_52 = '-2.02407e-12*lvhp_mobility*lvhp_mobility+-2.41712e-11*lvhp_mobility'
+ sky130_fd_pr__pfet_01v8_hvt__ua_diff_53 = '-4.94688e-12*lvhp_mobility*lvhp_mobility+1.91250e-11*lvhp_mobility'
+ sky130_fd_pr__pfet_01v8_hvt__ua_diff_54 = '6.11942e-11*lvhp_mobility*lvhp_mobility+1.12381e-10*lvhp_mobility'
+ sky130_fd_pr__pfet_01v8_hvt__ua_diff_55 = '1.00166e-11*lvhp_mobility*lvhp_mobility+-4.33750e-12*lvhp_mobility'
+ sky130_fd_pr__pfet_01v8_hvt__ua_diff_59 = '4.41631e-11*lvhp_mobility*lvhp_mobility+7.37328e-11*lvhp_mobility'
+ sky130_fd_pr__pfet_01v8_hvt__ua_diff_6 = '-2.02406e-12*lvhp_mobility*lvhp_mobility+-2.41713e-11*lvhp_mobility+3.46900e-10'
+ sky130_fd_pr__pfet_01v8_hvt__ua_diff_60 = '5.10381e-11*lvhp_mobility*lvhp_mobility+8.95350e-11*lvhp_mobility'
+ sky130_fd_pr__pfet_01v8_hvt__ua_diff_61 = '5.58609e-11*lvhp_mobility*lvhp_mobility+1.00459e-10*lvhp_mobility'
+ sky130_fd_pr__pfet_01v8_hvt__ua_diff_62 = '5.91450e-11*lvhp_mobility*lvhp_mobility+1.07820e-10*lvhp_mobility'
+ sky130_fd_pr__pfet_01v8_hvt__ua_diff_63 = '5.91447e-11*lvhp_mobility*lvhp_mobility+1.07819e-10*lvhp_mobility'
+ sky130_fd_pr__pfet_01v8_hvt__ua_diff_64 = '3.11262e-11*lvhp_mobility*lvhp_mobility+5.90796e-11*lvhp_mobility'
+ sky130_fd_pr__pfet_01v8_hvt__ua_diff_66 = '5.19170e-11*lvhp_mobility*lvhp_mobility+9.21769e-11*lvhp_mobility'
+ sky130_fd_pr__pfet_01v8_hvt__ua_diff_67 = '1.90034e-11*lvhp_mobility*lvhp_mobility+2.09540e-11*lvhp_mobility'
+ sky130_fd_pr__pfet_01v8_hvt__ua_diff_7 = '2.41375e-11*lvhp_mobility*lvhp_mobility+-4.13650e-11*lvhp_mobility+-4.50140e-10'
+ sky130_fd_pr__pfet_01v8_hvt__ua_diff_8 = '3.08406e-11*lvhp_mobility*lvhp_mobility+5.92500e-11*lvhp_mobility+1.60040e-10'
+ sky130_fd_pr__pfet_01v8_hvt__ua_diff_9 = '5.04919e-12*lvhp_mobility*lvhp_mobility+-1.59655e-10*lvhp_mobility+5.78330e-11'
+ sky130_fd_pr__pfet_01v8_hvt__ub_diff_0 = '-1.59750e-21*lvhp_mobility*lvhp_mobility+-7.15500e-22*lvhp_mobility+9.17100e-20'
+ sky130_fd_pr__pfet_01v8_hvt__ub_diff_1 = '4.37419e-21*lvhp_mobility*lvhp_mobility+-3.30443e-20*lvhp_mobility+-2.29020e-19'
+ sky130_fd_pr__pfet_01v8_hvt__ub_diff_10 = '6.74816e-21*lvhp_mobility*lvhp_mobility+-9.33349e-20*lvhp_mobility+2.45750e-19'
+ sky130_fd_pr__pfet_01v8_hvt__ub_diff_11 = '2.42146e-20*lvhp_mobility*lvhp_mobility+-1.23923e-19*lvhp_mobility+6.20770e-20'
+ sky130_fd_pr__pfet_01v8_hvt__ub_diff_12 = '3.38680e-20*lvhp_mobility*lvhp_mobility+-1.29661e-19*lvhp_mobility+1.84700e-20'
+ sky130_fd_pr__pfet_01v8_hvt__ub_diff_13 = '4.72352e-20*lvhp_mobility*lvhp_mobility+-1.78104e-19*lvhp_mobility+-2.08020e-21'
+ sky130_fd_pr__pfet_01v8_hvt__ub_diff_14 = '-2.74809e-21*lvhp_mobility*lvhp_mobility+-3.63763e-21*lvhp_mobility+7.06590e-20'
+ sky130_fd_pr__pfet_01v8_hvt__ub_diff_15 = '-6.86944e-21*lvhp_mobility*lvhp_mobility+-8.52750e-22*lvhp_mobility+2.08020e-19'
+ sky130_fd_pr__pfet_01v8_hvt__ub_diff_16 = '1.68281e-21*lvhp_mobility*lvhp_mobility+-1.27488e-20*lvhp_mobility+1.75980e-19'
+ sky130_fd_pr__pfet_01v8_hvt__ub_diff_17 = '4.59606e-21*lvhp_mobility*lvhp_mobility+-9.80350e-20*lvhp_mobility+4.25830e-20'
+ sky130_fd_pr__pfet_01v8_hvt__ub_diff_18 = '-3.02222e-21*lvhp_mobility*lvhp_mobility+-9.32439e-20*lvhp_mobility+4.41020e-19'
+ sky130_fd_pr__pfet_01v8_hvt__ub_diff_19 = '-4.71719e-21*lvhp_mobility*lvhp_mobility+-1.39831e-19*lvhp_mobility+5.22250e-19'
+ sky130_fd_pr__pfet_01v8_hvt__ub_diff_2 = '8.88437e-21*lvhp_mobility*lvhp_mobility+8.76475e-20*lvhp_mobility+3.87060e-19'
+ sky130_fd_pr__pfet_01v8_hvt__ub_diff_20 = '3.34313e-21*lvhp_mobility*lvhp_mobility+-1.78160e-19*lvhp_mobility+6.36170e-19'
+ sky130_fd_pr__pfet_01v8_hvt__ub_diff_21 = '-6.72219e-21*lvhp_mobility*lvhp_mobility+-2.13789e-19*lvhp_mobility+6.06700e-19'
+ sky130_fd_pr__pfet_01v8_hvt__ub_diff_22 = '-3.56972e-21*lvhp_mobility*lvhp_mobility+3.99362e-21*lvhp_mobility+2.71140e-20'
+ sky130_fd_pr__pfet_01v8_hvt__ub_diff_23 = '4.58250e-21*lvhp_mobility*lvhp_mobility+1.83585e-20*lvhp_mobility+7.60560e-20'
+ sky130_fd_pr__pfet_01v8_hvt__ub_diff_24 = '-2.10187e-21*lvhp_mobility*lvhp_mobility+-2.93725e-20*lvhp_mobility+2.66330e-19'
+ sky130_fd_pr__pfet_01v8_hvt__ub_diff_25 = '1.22391e-20*lvhp_mobility*lvhp_mobility+7.20937e-20*lvhp_mobility+2.63360e-19'
+ sky130_fd_pr__pfet_01v8_hvt__ub_diff_26 = '-6.50688e-21*lvhp_mobility*lvhp_mobility+-1.56975e-19*lvhp_mobility+5.62210e-19'
+ sky130_fd_pr__pfet_01v8_hvt__ub_diff_27 = '1.48437e-21*lvhp_mobility*lvhp_mobility+-2.00495e-19*lvhp_mobility+5.88070e-19'
+ sky130_fd_pr__pfet_01v8_hvt__ub_diff_28 = '1.79338e-20*lvhp_mobility*lvhp_mobility+-2.43848e-19*lvhp_mobility+2.98470e-19'
+ sky130_fd_pr__pfet_01v8_hvt__ub_diff_29 = '2.58419e-20*lvhp_mobility*lvhp_mobility+-2.76780e-19*lvhp_mobility+3.36710e-19'
+ sky130_fd_pr__pfet_01v8_hvt__ub_diff_3 = '6.69594e-21*lvhp_mobility*lvhp_mobility+-2.05687e-20*lvhp_mobility+3.29240e-19'
+ sky130_fd_pr__pfet_01v8_hvt__ub_diff_30 = '2.96844e-21*lvhp_mobility*lvhp_mobility+8.57375e-21*lvhp_mobility+-1.87160e-19'
+ sky130_fd_pr__pfet_01v8_hvt__ub_diff_31 = '-1.97781e-21*lvhp_mobility*lvhp_mobility+2.20462e-20*lvhp_mobility+3.08330e-19'
+ sky130_fd_pr__pfet_01v8_hvt__ub_diff_32 = '5.58906e-22*lvhp_mobility*lvhp_mobility+-1.97319e-20*lvhp_mobility+1.64510e-19'
+ sky130_fd_pr__pfet_01v8_hvt__ub_diff_33 = '2.43094e-21*lvhp_mobility*lvhp_mobility+2.82838e-20*lvhp_mobility+2.54240e-19'
+ sky130_fd_pr__pfet_01v8_hvt__ub_diff_34 = '1.27341e-20*lvhp_mobility*lvhp_mobility+-1.97249e-19*lvhp_mobility+3.43760e-19'
+ sky130_fd_pr__pfet_01v8_hvt__ub_diff_35 = '4.53844e-21*lvhp_mobility*lvhp_mobility+-9.73587e-20*lvhp_mobility+5.20050e-19'
+ sky130_fd_pr__pfet_01v8_hvt__ub_diff_36 = '3.76741e-20*lvhp_mobility*lvhp_mobility+-1.69749e-19*lvhp_mobility+-2.42810e-20'
+ sky130_fd_pr__pfet_01v8_hvt__ub_diff_37 = '3.60194e-20*lvhp_mobility*lvhp_mobility+1.62625e-19*lvhp_mobility+5.31590e-19'
+ sky130_fd_pr__pfet_01v8_hvt__ub_diff_38 = '3.19092e-20*lvhp_mobility*lvhp_mobility+1.43365e-19*lvhp_mobility+9.77920e-20'
+ sky130_fd_pr__pfet_01v8_hvt__ub_diff_39 = '-2.75590e-20*lvhp_mobility*lvhp_mobility+-1.47170e-19*lvhp_mobility+8.15540e-20'
+ sky130_fd_pr__pfet_01v8_hvt__ub_diff_4 = '5.38469e-21*lvhp_mobility*lvhp_mobility+-2.00625e-21*lvhp_mobility+3.56870e-19'
+ sky130_fd_pr__pfet_01v8_hvt__ub_diff_40 = '-2.53422e-20*lvhp_mobility*lvhp_mobility+6.67862e-21*lvhp_mobility+4.95610e-19'
+ sky130_fd_pr__pfet_01v8_hvt__ub_diff_41 = '8.17188e-22*lvhp_mobility*lvhp_mobility+-1.54674e-19*lvhp_mobility+2.19970e-19'
+ sky130_fd_pr__pfet_01v8_hvt__ub_diff_42 = '4.61309e-21*lvhp_mobility*lvhp_mobility+9.67026e-20*lvhp_mobility+2.69040e-19'
+ sky130_fd_pr__pfet_01v8_hvt__ub_diff_43 = '1.03094e-20*lvhp_mobility*lvhp_mobility+6.61975e-20*lvhp_mobility+3.84820e-19'
+ sky130_fd_pr__pfet_01v8_hvt__ub_diff_44 = '1.28866e-20*lvhp_mobility*lvhp_mobility+2.85563e-20*lvhp_mobility+4.68000e-19'
+ sky130_fd_pr__pfet_01v8_hvt__ub_diff_45 = '4.53268e-20*lvhp_mobility*lvhp_mobility+2.83750e-20*lvhp_mobility+-3.45390e-20'
+ sky130_fd_pr__pfet_01v8_hvt__ub_diff_46 = '6.20703e-21*lvhp_mobility*lvhp_mobility+-2.20709e-20*lvhp_mobility+-2.83760e-20'
+ sky130_fd_pr__pfet_01v8_hvt__ub_diff_47 = '1.49531e-21*lvhp_mobility*lvhp_mobility+-2.08989e-19*lvhp_mobility+2.76820e-19'
+ sky130_fd_pr__pfet_01v8_hvt__ub_diff_48 = '-3.47972e-20*lvhp_mobility*lvhp_mobility+-1.42679e-19*lvhp_mobility+1.59470e-19'
+ sky130_fd_pr__pfet_01v8_hvt__ub_diff_49 = '-5.00816e-20*lvhp_mobility*lvhp_mobility+-1.49984e-19*lvhp_mobility+7.60400e-20'
+ sky130_fd_pr__pfet_01v8_hvt__ub_diff_5 = '3.85625e-21*lvhp_mobility*lvhp_mobility+5.59250e-21*lvhp_mobility+3.63070e-19'
+ sky130_fd_pr__pfet_01v8_hvt__ub_diff_50 = '-3.47972e-20*lvhp_mobility*lvhp_mobility+-1.42679e-19*lvhp_mobility'
+ sky130_fd_pr__pfet_01v8_hvt__ub_diff_51 = '-2.74809e-21*lvhp_mobility*lvhp_mobility+-3.63762e-21*lvhp_mobility'
+ sky130_fd_pr__pfet_01v8_hvt__ub_diff_52 = '2.14317e-21*lvhp_mobility*lvhp_mobility+-1.73326e-20*lvhp_mobility'
+ sky130_fd_pr__pfet_01v8_hvt__ub_diff_53 = '4.37419e-21*lvhp_mobility*lvhp_mobility+-3.30443e-20*lvhp_mobility'
+ sky130_fd_pr__pfet_01v8_hvt__ub_diff_54 = '-5.00816e-20*lvhp_mobility*lvhp_mobility+-1.49984e-19*lvhp_mobility'
+ sky130_fd_pr__pfet_01v8_hvt__ub_diff_55 = '-6.86944e-21*lvhp_mobility*lvhp_mobility+-8.52750e-22*lvhp_mobility'
+ sky130_fd_pr__pfet_01v8_hvt__ub_diff_59 = '-4.03444e-20*lvhp_mobility*lvhp_mobility+-1.45695e-19*lvhp_mobility'
+ sky130_fd_pr__pfet_01v8_hvt__ub_diff_6 = '2.14313e-21*lvhp_mobility*lvhp_mobility+-1.73325e-20*lvhp_mobility+-2.42240e-19'
+ sky130_fd_pr__pfet_01v8_hvt__ub_diff_60 = '-4.42575e-20*lvhp_mobility*lvhp_mobility+-1.47573e-19*lvhp_mobility'
+ sky130_fd_pr__pfet_01v8_hvt__ub_diff_61 = '-4.70164e-20*lvhp_mobility*lvhp_mobility+-1.48772e-19*lvhp_mobility'
+ sky130_fd_pr__pfet_01v8_hvt__ub_diff_62 = '-4.89020e-20*lvhp_mobility*lvhp_mobility+-1.49532e-19*lvhp_mobility'
+ sky130_fd_pr__pfet_01v8_hvt__ub_diff_63 = '-4.89020e-20*lvhp_mobility*lvhp_mobility+-1.49532e-19*lvhp_mobility'
+ sky130_fd_pr__pfet_01v8_hvt__ub_diff_64 = '-2.57202e-20*lvhp_mobility*lvhp_mobility+-2.00142e-19*lvhp_mobility'
+ sky130_fd_pr__pfet_01v8_hvt__ub_diff_66 = '-4.24099e-20*lvhp_mobility*lvhp_mobility+-1.30415e-19*lvhp_mobility'
+ sky130_fd_pr__pfet_01v8_hvt__ub_diff_67 = '-1.52140e-20*lvhp_mobility*lvhp_mobility+-6.12742e-20*lvhp_mobility'
+ sky130_fd_pr__pfet_01v8_hvt__ub_diff_7 = '-2.05929e-20*lvhp_mobility*lvhp_mobility+-4.01990e-20*lvhp_mobility+5.06610e-19'
+ sky130_fd_pr__pfet_01v8_hvt__ub_diff_8 = '-2.49204e-20*lvhp_mobility*lvhp_mobility+-2.04647e-19*lvhp_mobility+-7.40840e-20'
+ sky130_fd_pr__pfet_01v8_hvt__ub_diff_9 = '-5.90225e-21*lvhp_mobility*lvhp_mobility+3.00315e-20*lvhp_mobility+2.56470e-19'
+ sky130_fd_pr__pfet_01v8_hvt__voff_diff_0 = '4.86250e-05*lvp_subvt*lvp_subvt+1.79668e-02*lvp_subvt+-2.69220e-02'
+ sky130_fd_pr__pfet_01v8_hvt__voff_diff_1 = '-2.52531e-04*lvp_subvt*lvp_subvt+2.26864e-02*lvp_subvt+-3.22440e-02'
+ sky130_fd_pr__pfet_01v8_hvt__voff_diff_10 = '9.43406e-05*lvp_subvt*lvp_subvt+8.51136e-03*lvp_subvt+-3.85630e-02'
+ sky130_fd_pr__pfet_01v8_hvt__voff_diff_11 = '-5.69625e-04*lvp_subvt*lvp_subvt+1.15847e-02*lvp_subvt+-4.72570e-02'
+ sky130_fd_pr__pfet_01v8_hvt__voff_diff_12 = '-1.20240e-03*lvp_subvt*lvp_subvt+1.20790e-02*lvp_subvt+1.79410e-04'
+ sky130_fd_pr__pfet_01v8_hvt__voff_diff_13 = '-1.29145e-03*lvp_subvt*lvp_subvt+9.42404e-03*lvp_subvt+-7.97770e-03'
+ sky130_fd_pr__pfet_01v8_hvt__voff_diff_14 = '-2.24219e-04*lvp_subvt*lvp_subvt+1.97096e-02*lvp_subvt+-4.13240e-02'
+ sky130_fd_pr__pfet_01v8_hvt__voff_diff_15 = '3.46406e-04*lvp_subvt*lvp_subvt+1.04041e-02*lvp_subvt+-5.76800e-02'
+ sky130_fd_pr__pfet_01v8_hvt__voff_diff_16 = '4.12300e-04*lvp_subvt*lvp_subvt+5.32395e-03*lvp_subvt+-2.99910e-02'
+ sky130_fd_pr__pfet_01v8_hvt__voff_diff_17 = '-8.33047e-04*lvp_subvt*lvp_subvt+9.70706e-03*lvp_subvt+-2.11290e-02'
+ sky130_fd_pr__pfet_01v8_hvt__voff_diff_18 = '1.67813e-04*lvp_subvt*lvp_subvt+6.87600e-03*lvp_subvt+-4.02010e-02'
+ sky130_fd_pr__pfet_01v8_hvt__voff_diff_19 = '4.57481e-04*lvp_subvt*lvp_subvt+9.91218e-03*lvp_subvt+-4.47170e-02'
+ sky130_fd_pr__pfet_01v8_hvt__voff_diff_2 = '-6.75625e-05*lvp_subvt*lvp_subvt+3.40200e-03*lvp_subvt+-3.85210e-02'
+ sky130_fd_pr__pfet_01v8_hvt__voff_diff_20 = '5.27806e-04*lvp_subvt*lvp_subvt+9.35373e-03*lvp_subvt+-3.70850e-02'
+ sky130_fd_pr__pfet_01v8_hvt__voff_diff_21 = '2.09194e-03*lvp_subvt*lvp_subvt+9.06525e-03*lvp_subvt+-4.09900e-02'
+ sky130_fd_pr__pfet_01v8_hvt__voff_diff_22 = '-1.43719e-04*lvp_subvt*lvp_subvt+1.53789e-02*lvp_subvt+-2.07790e-02'
+ sky130_fd_pr__pfet_01v8_hvt__voff_diff_23 = '-5.64450e-04*lvp_subvt*lvp_subvt+7.05170e-03*lvp_subvt+-1.09740e-02'
+ sky130_fd_pr__pfet_01v8_hvt__voff_diff_24 = '7.09281e-05*lvp_subvt*lvp_subvt+5.22071e-03*lvp_subvt+-3.09090e-02'
+ sky130_fd_pr__pfet_01v8_hvt__voff_diff_25 = '1.36862e-04*lvp_subvt*lvp_subvt+6.06045e-03*lvp_subvt+-3.41500e-02'
+ sky130_fd_pr__pfet_01v8_hvt__voff_diff_26 = '5.88491e-04*lvp_subvt*lvp_subvt+7.80546e-03*lvp_subvt+-4.47410e-02'
+ sky130_fd_pr__pfet_01v8_hvt__voff_diff_27 = '6.60063e-04*lvp_subvt*lvp_subvt+9.55275e-03*lvp_subvt+-3.04870e-02'
+ sky130_fd_pr__pfet_01v8_hvt__voff_diff_28 = '-9.54478e-04*lvp_subvt*lvp_subvt+6.06299e-03*lvp_subvt+-5.90340e-03'
+ sky130_fd_pr__pfet_01v8_hvt__voff_diff_29 = '5.20437e-05*lvp_subvt*lvp_subvt+6.90763e-03*lvp_subvt+-7.82520e-03'
+ sky130_fd_pr__pfet_01v8_hvt__voff_diff_3 = '-1.16500e-04*lvp_subvt*lvp_subvt+3.09325e-03*lvp_subvt+-2.60130e-02'
+ sky130_fd_pr__pfet_01v8_hvt__voff_diff_30 = '-3.18000e-04*lvp_subvt*lvp_subvt+1.35643e-02*lvp_subvt+-2.88430e-02'
+ sky130_fd_pr__pfet_01v8_hvt__voff_diff_31 = '-1.30312e-04*lvp_subvt*lvp_subvt+9.28725e-03*lvp_subvt+-4.74650e-02'
+ sky130_fd_pr__pfet_01v8_hvt__voff_diff_32 = '1.93341e-04*lvp_subvt*lvp_subvt+9.34436e-03*lvp_subvt+-3.26360e-02'
+ sky130_fd_pr__pfet_01v8_hvt__voff_diff_33 = '-1.37116e-03*lvp_subvt*lvp_subvt+3.10638e-03*lvp_subvt+-1.29800e-02'
+ sky130_fd_pr__pfet_01v8_hvt__voff_diff_34 = '-5.81344e-04*lvp_subvt*lvp_subvt+1.60289e-02*lvp_subvt+-5.41930e-02'
+ sky130_fd_pr__pfet_01v8_hvt__voff_diff_35 = '7.44541e-04*lvp_subvt*lvp_subvt+1.28379e-02*lvp_subvt+-5.54370e-02'
+ sky130_fd_pr__pfet_01v8_hvt__voff_diff_36 = '-1.94313e-03*lvp_subvt*lvp_subvt+1.42368e-02*lvp_subvt+-1.18200e-02'
+ sky130_fd_pr__pfet_01v8_hvt__voff_diff_37 = '6.46875e-06*lvp_subvt*lvp_subvt+6.58388e-03*lvp_subvt+-5.01470e-02'
+ sky130_fd_pr__pfet_01v8_hvt__voff_diff_38 = '-2.84900e-03*lvp_subvt*lvp_subvt+6.47500e-03*lvp_subvt+-1.57280e-02'
+ sky130_fd_pr__pfet_01v8_hvt__voff_diff_39 = '1.58594e-03*lvp_subvt*lvp_subvt+3.73340e-02*lvp_subvt+-7.57190e-02'
+ sky130_fd_pr__pfet_01v8_hvt__voff_diff_4 = '-1.47813e-04*lvp_subvt*lvp_subvt+5.17900e-03*lvp_subvt+-4.04910e-02'
+ sky130_fd_pr__pfet_01v8_hvt__voff_diff_40 = '1.52678e-03*lvp_subvt*lvp_subvt+3.66794e-02*lvp_subvt+-7.44510e-02'
+ sky130_fd_pr__pfet_01v8_hvt__voff_diff_41 = '-8.88125e-05*lvp_subvt*lvp_subvt+1.28568e-02*lvp_subvt+-4.01660e-02'
+ sky130_fd_pr__pfet_01v8_hvt__voff_diff_42 = '9.24375e-05*lvp_subvt*lvp_subvt+5.78475e-03*lvp_subvt+-6.67700e-02'
+ sky130_fd_pr__pfet_01v8_hvt__voff_diff_43 = '-1.55969e-04*lvp_subvt*lvp_subvt+4.29838e-03*lvp_subvt+-4.21590e-02'
+ sky130_fd_pr__pfet_01v8_hvt__voff_diff_44 = '-1.91719e-04*lvp_subvt*lvp_subvt+4.93563e-03*lvp_subvt+-4.65460e-02'
+ sky130_fd_pr__pfet_01v8_hvt__voff_diff_45 = '-1.96322e-03*lvp_subvt*lvp_subvt+4.73913e-03*lvp_subvt+-1.72830e-02'
+ sky130_fd_pr__pfet_01v8_hvt__voff_diff_46 = '3.89831e-03*lvp_subvt*lvp_subvt+3.83875e-02*lvp_subvt+-4.71330e-02'
+ sky130_fd_pr__pfet_01v8_hvt__voff_diff_47 = '6.37813e-05*lvp_subvt*lvp_subvt+1.04361e-02*lvp_subvt+-3.49900e-02'
+ sky130_fd_pr__pfet_01v8_hvt__voff_diff_48 = '2.24866e-03*lvp_subvt*lvp_subvt+3.48319e-02*lvp_subvt+-9.22610e-02'
+ sky130_fd_pr__pfet_01v8_hvt__voff_diff_49 = '-1.91982e-03*lvp_subvt*lvp_subvt+1.97850e-02*lvp_subvt+-4.90030e-02'
+ sky130_fd_pr__pfet_01v8_hvt__voff_diff_5 = '-7.64688e-05*lvp_subvt*lvp_subvt+4.97413e-03*lvp_subvt+-4.22550e-02'
+ sky130_fd_pr__pfet_01v8_hvt__voff_diff_50 = '2.24866e-03*lvp_subvt*lvp_subvt+3.48319e-02*lvp_subvt'
+ sky130_fd_pr__pfet_01v8_hvt__voff_diff_51 = '-2.24219e-04*lvp_subvt*lvp_subvt+1.97096e-02*lvp_subvt'
+ sky130_fd_pr__pfet_01v8_hvt__voff_diff_52 = '4.02291e-04*lvp_subvt*lvp_subvt+1.96197e-02*lvp_subvt'
+ sky130_fd_pr__pfet_01v8_hvt__voff_diff_53 = '-2.52532e-04*lvp_subvt*lvp_subvt+2.26864e-02*lvp_subvt'
+ sky130_fd_pr__pfet_01v8_hvt__voff_diff_54 = '-1.91982e-03*lvp_subvt*lvp_subvt+1.97850e-02*lvp_subvt'
+ sky130_fd_pr__pfet_01v8_hvt__voff_diff_55 = '3.46406e-04*lvp_subvt*lvp_subvt+1.04041e-02*lvp_subvt'
+ sky130_fd_pr__pfet_01v8_hvt__voff_diff_59 = '7.18244e-04*lvp_subvt*lvp_subvt+2.93487e-02*lvp_subvt'
+ sky130_fd_pr__pfet_01v8_hvt__voff_diff_6 = '4.02291e-04*lvp_subvt*lvp_subvt+1.96197e-02*lvp_subvt+-8.08380e-02'
+ sky130_fd_pr__pfet_01v8_hvt__voff_diff_60 = '-3.49498e-04*lvp_subvt*lvp_subvt+2.54957e-02*lvp_subvt'
+ sky130_fd_pr__pfet_01v8_hvt__voff_diff_61 = '-1.09622e-03*lvp_subvt*lvp_subvt+2.27869e-02*lvp_subvt'
+ sky130_fd_pr__pfet_01v8_hvt__voff_diff_62 = '-1.60365e-03*lvp_subvt*lvp_subvt+2.09392e-02*lvp_subvt'
+ sky130_fd_pr__pfet_01v8_hvt__voff_diff_63 = '-1.60365e-03*lvp_subvt*lvp_subvt+2.09392e-02*lvp_subvt'
+ sky130_fd_pr__pfet_01v8_hvt__voff_diff_64 = '7.27984e-04*lvp_subvt*lvp_subvt+9.05166e-03*lvp_subvt'
+ sky130_fd_pr__pfet_01v8_hvt__voff_diff_66 = '-1.58140e-03*lvp_subvt*lvp_subvt+1.97567e-02*lvp_subvt'
+ sky130_fd_pr__pfet_01v8_hvt__voff_diff_67 = '-3.74228e-04*lvp_subvt*lvp_subvt+1.96674e-02*lvp_subvt'
+ sky130_fd_pr__pfet_01v8_hvt__voff_diff_7 = '1.56884e-03*lvp_subvt*lvp_subvt+2.51996e-02*lvp_subvt+-3.74530e-02'
+ sky130_fd_pr__pfet_01v8_hvt__voff_diff_8 = '6.13419e-04*lvp_subvt*lvp_subvt+6.86367e-03*lvp_subvt+-2.76990e-02'
+ sky130_fd_pr__pfet_01v8_hvt__voff_diff_9 = '3.86750e-04*lvp_subvt*lvp_subvt+9.16700e-03*lvp_subvt+-4.28560e-02'
+ sky130_fd_pr__pfet_01v8_hvt__vsat_diff_0 = '1.64331e+02*lvhp_saturation*lvhp_saturation+6.22162e+03*lvhp_saturation+-7.41680e+03'
+ sky130_fd_pr__pfet_01v8_hvt__vsat_diff_1 = '-9.78231e+02*lvhp_saturation*lvhp_saturation+1.40625e+02*lvhp_saturation+-7.42680e+03'
+ sky130_fd_pr__pfet_01v8_hvt__vsat_diff_14 = '-6.06156e+02*lvhp_saturation*lvhp_saturation+1.12288e+03*lvhp_saturation+-1.02540e+04'
+ sky130_fd_pr__pfet_01v8_hvt__vsat_diff_15 = '-1.07521e+03*lvhp_saturation*lvhp_saturation+5.55657e+03*lvhp_saturation+3.29240e+04'
+ sky130_fd_pr__pfet_01v8_hvt__vsat_diff_16 = '5.39688e+01*lvhp_saturation*lvhp_saturation+6.91325e+03*lvhp_saturation+-1.97250e+03'
+ sky130_fd_pr__pfet_01v8_hvt__vsat_diff_17 = '6.87227e+02*lvhp_saturation*lvhp_saturation+-6.74562e+02*lvhp_saturation+1.65110e+02'
+ sky130_fd_pr__pfet_01v8_hvt__vsat_diff_22 = '-5.92656e+02*lvhp_saturation*lvhp_saturation+1.05638e+03*lvhp_saturation+-1.30870e+04'
+ sky130_fd_pr__pfet_01v8_hvt__vsat_diff_23 = '-8.09312e+02*lvhp_saturation*lvhp_saturation+6.60575e+03*lvhp_saturation+1.87530e+04'
+ sky130_fd_pr__pfet_01v8_hvt__vsat_diff_24 = '-5.81913e+02*lvhp_saturation*lvhp_saturation+2.90275e+03*lvhp_saturation+9.90560e+03'
+ sky130_fd_pr__pfet_01v8_hvt__vsat_diff_25 = '9.05003e+02*lvhp_saturation*lvhp_saturation+1.53600e+04*lvhp_saturation+4.40800e+04'
+ sky130_fd_pr__pfet_01v8_hvt__vsat_diff_30 = '-6.31100e+02*lvhp_saturation*lvhp_saturation+5.64000e+02*lvhp_saturation+-6.54340e+03'
+ sky130_fd_pr__pfet_01v8_hvt__vsat_diff_31 = '-6.80000e+02*lvhp_saturation*lvhp_saturation+4.32300e+03*lvhp_saturation+2.39240e+04'
+ sky130_fd_pr__pfet_01v8_hvt__vsat_diff_32 = '-4.31146e+02*lvhp_saturation*lvhp_saturation+1.46679e+03*lvhp_saturation+1.01050e+03'
+ sky130_fd_pr__pfet_01v8_hvt__vsat_diff_33 = '-7.86906e+02*lvhp_saturation*lvhp_saturation+1.28389e+04*lvhp_saturation+3.12350e+04'
+ sky130_fd_pr__pfet_01v8_hvt__vsat_diff_34 = '5.44125e+00*lvhp_saturation*lvhp_saturation+2.17650e+01*lvhp_saturation'
+ sky130_fd_pr__pfet_01v8_hvt__vsat_diff_36 = '-1.23431e+00*lvhp_saturation*lvhp_saturation+-4.93725e+00*lvhp_saturation'
+ sky130_fd_pr__pfet_01v8_hvt__vsat_diff_39 = '-1.70516e+03*lvhp_saturation*lvhp_saturation+6.23900e+03*lvhp_saturation+2.23850e+03'
+ sky130_fd_pr__pfet_01v8_hvt__vsat_diff_40 = '-1.32234e+03*lvhp_saturation*lvhp_saturation+1.42086e+04*lvhp_saturation+3.28430e+04'
+ sky130_fd_pr__pfet_01v8_hvt__vsat_diff_41 = '-2.37009e+03*lvhp_saturation*lvhp_saturation+6.00715e+03*lvhp_saturation+2.30610e+04'
+ sky130_fd_pr__pfet_01v8_hvt__vsat_diff_46 = '-2.82200e+02*lvhp_saturation*lvhp_saturation+1.12629e+04*lvhp_saturation+8.98470e+03'
+ sky130_fd_pr__pfet_01v8_hvt__vsat_diff_47 = '-1.06888e+03*lvhp_saturation*lvhp_saturation+4.93250e+03*lvhp_saturation+-1.31680e+04'
+ sky130_fd_pr__pfet_01v8_hvt__vsat_diff_48 = '-1.27238e+03*lvhp_saturation*lvhp_saturation+2.38386e+03*lvhp_saturation+5.42160e+03'
+ sky130_fd_pr__pfet_01v8_hvt__vsat_diff_49 = '-5.78133e+02*lvhp_saturation*lvhp_saturation+3.83962e+03*lvhp_saturation+-6.14640e+03'
+ sky130_fd_pr__pfet_01v8_hvt__vsat_diff_50 = '-1.27238e+03*lvhp_saturation*lvhp_saturation+2.38386e+03*lvhp_saturation'
+ sky130_fd_pr__pfet_01v8_hvt__vsat_diff_51 = '-6.06158e+02*lvhp_saturation*lvhp_saturation+1.12287e+03*lvhp_saturation'
+ sky130_fd_pr__pfet_01v8_hvt__vsat_diff_52 = '-2.06312e+02*lvhp_saturation*lvhp_saturation+5.82725e+03*lvhp_saturation'
+ sky130_fd_pr__pfet_01v8_hvt__vsat_diff_53 = '-9.78231e+02*lvhp_saturation*lvhp_saturation+1.40624e+02*lvhp_saturation'
+ sky130_fd_pr__pfet_01v8_hvt__vsat_diff_54 = '-5.78130e+02*lvhp_saturation*lvhp_saturation+3.83962e+03*lvhp_saturation'
+ sky130_fd_pr__pfet_01v8_hvt__vsat_diff_55 = '-1.07521e+03*lvhp_saturation*lvhp_saturation+5.55658e+03*lvhp_saturation'
+ sky130_fd_pr__pfet_01v8_hvt__vsat_diff_56 = '-4.50444e+03*lvhp_saturation*lvhp_saturation+1.00225e+04*lvhp_saturation+8.19810e+04'
+ sky130_fd_pr__pfet_01v8_hvt__vsat_diff_57 = '7.65094e+02*lvhp_saturation*lvhp_saturation+3.20841e+04*lvhp_saturation+7.83720e+04'
+ sky130_fd_pr__pfet_01v8_hvt__vsat_diff_58 = '2.16531e+03*lvhp_saturation*lvhp_saturation+2.53708e+04*lvhp_saturation+3.62020e+04'
+ sky130_fd_pr__pfet_01v8_hvt__vsat_diff_59 = '4.37484e+03*lvhp_saturation*lvhp_saturation+3.07001e+04*lvhp_saturation+2.56020e+04'
+ sky130_fd_pr__pfet_01v8_hvt__vsat_diff_6 = '-2.06312e+02*lvhp_saturation*lvhp_saturation+5.82725e+03*lvhp_saturation+-1.06000e+03'
+ sky130_fd_pr__pfet_01v8_hvt__vsat_diff_60 = '5.74216e+03*lvhp_saturation*lvhp_saturation+3.56804e+04*lvhp_saturation+2.54540e+04'
+ sky130_fd_pr__pfet_01v8_hvt__vsat_diff_61 = '6.66816e+03*lvhp_saturation*lvhp_saturation+4.16316e+04*lvhp_saturation+3.60530e+04'
+ sky130_fd_pr__pfet_01v8_hvt__vsat_diff_62 = '6.69912e+03*lvhp_saturation*lvhp_saturation+4.17638e+04*lvhp_saturation+3.79690e+04'
+ sky130_fd_pr__pfet_01v8_hvt__vsat_diff_63 = '5.68928e+03*lvhp_saturation*lvhp_saturation+3.55581e+04*lvhp_saturation+2.76690e+04'
+ sky130_fd_pr__pfet_01v8_hvt__vsat_diff_64 = '-1.88616e+03*lvhp_saturation*lvhp_saturation+1.19129e+04*lvhp_saturation+5.86070e+04'
+ sky130_fd_pr__pfet_01v8_hvt__vsat_diff_65 = '-2.09984e+03*lvhp_saturation*lvhp_saturation+8.14838e+03*lvhp_saturation+5.10040e+04'
+ sky130_fd_pr__pfet_01v8_hvt__vsat_diff_66 = '5.38934e+03*lvhp_saturation*lvhp_saturation+3.95031e+04*lvhp_saturation+5.28180e+04'
+ sky130_fd_pr__pfet_01v8_hvt__vsat_diff_67 = '5.06166e+03*lvhp_saturation*lvhp_saturation+4.08251e+04*lvhp_saturation+6.46030e+04'
+ sky130_fd_pr__pfet_01v8_hvt__vsat_diff_7 = '-2.72381e+03*lvhp_saturation*lvhp_saturation+6.54775e+03*lvhp_saturation+5.37820e+04'
+ sky130_fd_pr__pfet_01v8_hvt__vsat_diff_8 = '-2.06085e+03*lvhp_saturation*lvhp_saturation+-1.28762e+03*lvhp_saturation+-2.12090e+03'
+ sky130_fd_pr__pfet_01v8_hvt__vsat_diff_9 = '9.47016e+03*lvhp_saturation*lvhp_saturation+5.13171e+04*lvhp_saturation+4.32090e+04'
+ sky130_fd_pr__pfet_01v8_hvt__vth0_diff_0 = '-1.37425e-03*lvhp_threshold*lvhp_threshold+8.90425e-03*lvhp_threshold+2.72530e-02'
+ sky130_fd_pr__pfet_01v8_hvt__vth0_diff_1 = '-1.21278e-03*lvhp_threshold*lvhp_threshold+1.29531e-02*lvhp_threshold+1.19210e-02'
+ sky130_fd_pr__pfet_01v8_hvt__vth0_diff_10 = '1.65700e-04*lvhp_threshold*lvhp_threshold+-3.98325e-03*lvhp_threshold+1.56780e-03'
+ sky130_fd_pr__pfet_01v8_hvt__vth0_diff_11 = '2.15707e-04*lvhp_threshold*lvhp_threshold+-2.77416e-03*lvhp_threshold+-9.26960e-04'
+ sky130_fd_pr__pfet_01v8_hvt__vth0_diff_12 = '-5.77237e-04*lvhp_threshold*lvhp_threshold+1.80947e-03*lvhp_threshold+-8.99310e-04'
+ sky130_fd_pr__pfet_01v8_hvt__vth0_diff_13 = '-3.88134e-04*lvhp_threshold*lvhp_threshold+5.71712e-04*lvhp_threshold+1.07670e-02'
+ sky130_fd_pr__pfet_01v8_hvt__vth0_diff_14 = '-1.46084e-03*lvhp_threshold*lvhp_threshold+1.30116e-02*lvhp_threshold+2.55280e-02'
+ sky130_fd_pr__pfet_01v8_hvt__vth0_diff_15 = '-1.14877e-03*lvhp_threshold*lvhp_threshold+1.09909e-02*lvhp_threshold+-8.91020e-03'
+ sky130_fd_pr__pfet_01v8_hvt__vth0_diff_16 = '-3.02344e-04*lvhp_threshold*lvhp_threshold+-4.37037e-03*lvhp_threshold+-1.43260e-02'
+ sky130_fd_pr__pfet_01v8_hvt__vth0_diff_17 = '1.70794e-04*lvhp_threshold*lvhp_threshold+-2.44167e-03*lvhp_threshold+4.05460e-03'
+ sky130_fd_pr__pfet_01v8_hvt__vth0_diff_18 = '1.53830e-04*lvhp_threshold*lvhp_threshold+-3.65675e-03*lvhp_threshold+-9.67280e-04'
+ sky130_fd_pr__pfet_01v8_hvt__vth0_diff_19 = '6.83278e-04*lvhp_threshold*lvhp_threshold+3.74887e-04*lvhp_threshold+-6.52710e-03'
+ sky130_fd_pr__pfet_01v8_hvt__vth0_diff_2 = '-2.83625e-04*lvhp_threshold*lvhp_threshold+-1.06702e-02*lvhp_threshold+-1.16230e-02'
+ sky130_fd_pr__pfet_01v8_hvt__vth0_diff_20 = '6.29834e-04*lvhp_threshold*lvhp_threshold+3.84738e-04*lvhp_threshold+-7.06010e-03'
+ sky130_fd_pr__pfet_01v8_hvt__vth0_diff_21 = '5.08844e-04*lvhp_threshold*lvhp_threshold+8.13625e-04*lvhp_threshold+1.21930e-02'
+ sky130_fd_pr__pfet_01v8_hvt__vth0_diff_22 = '-1.45443e-03*lvhp_threshold*lvhp_threshold+1.44575e-02*lvhp_threshold+9.52590e-03'
+ sky130_fd_pr__pfet_01v8_hvt__vth0_diff_23 = '-8.30800e-04*lvhp_threshold*lvhp_threshold+1.11301e-02*lvhp_threshold+7.53730e-03'
+ sky130_fd_pr__pfet_01v8_hvt__vth0_diff_24 = '-2.22569e-04*lvhp_threshold*lvhp_threshold+-2.52973e-03*lvhp_threshold+-1.42740e-02'
+ sky130_fd_pr__pfet_01v8_hvt__vth0_diff_25 = '1.90750e-05*lvhp_threshold*lvhp_threshold+-5.39650e-03*lvhp_threshold+6.63580e-03'
+ sky130_fd_pr__pfet_01v8_hvt__vth0_diff_26 = '5.89734e-04*lvhp_threshold*lvhp_threshold+-1.06999e-03*lvhp_threshold+-7.12890e-03'
+ sky130_fd_pr__pfet_01v8_hvt__vth0_diff_27 = '8.46712e-04*lvhp_threshold*lvhp_threshold+1.72790e-03*lvhp_threshold+-3.64800e-03'
+ sky130_fd_pr__pfet_01v8_hvt__vth0_diff_28 = '4.25681e-04*lvhp_threshold*lvhp_threshold+-4.49625e-04*lvhp_threshold+9.13660e-03'
+ sky130_fd_pr__pfet_01v8_hvt__vth0_diff_29 = '1.08875e-04*lvhp_threshold*lvhp_threshold+-8.57125e-04*lvhp_threshold+3.59050e-03'
+ sky130_fd_pr__pfet_01v8_hvt__vth0_diff_3 = '-9.69750e-05*lvhp_threshold*lvhp_threshold+-8.72137e-03*lvhp_threshold+3.56510e-03'
+ sky130_fd_pr__pfet_01v8_hvt__vth0_diff_30 = '-1.30456e-03*lvhp_threshold*lvhp_threshold+1.38431e-02*lvhp_threshold+2.51740e-03'
+ sky130_fd_pr__pfet_01v8_hvt__vth0_diff_31 = '-1.07006e-03*lvhp_threshold*lvhp_threshold+1.20820e-02*lvhp_threshold+-1.98520e-02'
+ sky130_fd_pr__pfet_01v8_hvt__vth0_diff_32 = '-6.65969e-05*lvhp_threshold*lvhp_threshold+-5.44037e-04*lvhp_threshold+-4.67620e-03'
+ sky130_fd_pr__pfet_01v8_hvt__vth0_diff_33 = '1.08456e-04*lvhp_threshold*lvhp_threshold+-4.25412e-03*lvhp_threshold+-5.31080e-03'
+ sky130_fd_pr__pfet_01v8_hvt__vth0_diff_34 = '3.34219e-04*lvhp_threshold*lvhp_threshold+-1.33746e-02*lvhp_threshold+-1.26190e-02'
+ sky130_fd_pr__pfet_01v8_hvt__vth0_diff_35 = '5.64709e-04*lvhp_threshold*lvhp_threshold+-6.58159e-03*lvhp_threshold+-4.41120e-02'
+ sky130_fd_pr__pfet_01v8_hvt__vth0_diff_36 = '-2.15413e-03*lvhp_threshold*lvhp_threshold+-1.07874e-02*lvhp_threshold+5.18360e-03'
+ sky130_fd_pr__pfet_01v8_hvt__vth0_diff_37 = '-6.18188e-04*lvhp_threshold*lvhp_threshold+-1.63155e-02*lvhp_threshold+-2.15150e-02'
+ sky130_fd_pr__pfet_01v8_hvt__vth0_diff_38 = '-2.14915e-03*lvhp_threshold*lvhp_threshold+-1.45129e-02*lvhp_threshold+-2.02020e-02'
+ sky130_fd_pr__pfet_01v8_hvt__vth0_diff_39 = '6.56156e-04*lvhp_threshold*lvhp_threshold+2.66363e-03*lvhp_threshold+4.02580e-02'
+ sky130_fd_pr__pfet_01v8_hvt__vth0_diff_4 = '-1.07527e-04*lvhp_threshold*lvhp_threshold+-8.00875e-03*lvhp_threshold+-8.89570e-04'
+ sky130_fd_pr__pfet_01v8_hvt__vth0_diff_40 = '-6.03719e-04*lvhp_threshold*lvhp_threshold+3.12212e-03*lvhp_threshold+2.71580e-02'
+ sky130_fd_pr__pfet_01v8_hvt__vth0_diff_41 = '2.30375e-04*lvhp_threshold*lvhp_threshold+-1.45493e-02*lvhp_threshold+2.95960e-02'
+ sky130_fd_pr__pfet_01v8_hvt__vth0_diff_42 = '-5.29906e-04*lvhp_threshold*lvhp_threshold+-1.57471e-02*lvhp_threshold+-1.98440e-02'
+ sky130_fd_pr__pfet_01v8_hvt__vth0_diff_43 = '-4.59306e-04*lvhp_threshold*lvhp_threshold+-1.32059e-02*lvhp_threshold+-3.78860e-03'
+ sky130_fd_pr__pfet_01v8_hvt__vth0_diff_44 = '-3.40094e-04*lvhp_threshold*lvhp_threshold+-1.23694e-02*lvhp_threshold+-1.12460e-02'
+ sky130_fd_pr__pfet_01v8_hvt__vth0_diff_45 = '-2.01334e-03*lvhp_threshold*lvhp_threshold+-1.13054e-02*lvhp_threshold+1.32750e-02'
+ sky130_fd_pr__pfet_01v8_hvt__vth0_diff_46 = '2.24391e-03*lvhp_threshold*lvhp_threshold+1.58096e-02*lvhp_threshold+-1.21260e-02'
+ sky130_fd_pr__pfet_01v8_hvt__vth0_diff_47 = '-1.77250e-04*lvhp_threshold*lvhp_threshold+-1.49235e-02*lvhp_threshold+1.78500e-02'
+ sky130_fd_pr__pfet_01v8_hvt__vth0_diff_48 = '-2.81250e-06*lvhp_threshold*lvhp_threshold+1.03083e-02*lvhp_threshold+1.80440e-02'
+ sky130_fd_pr__pfet_01v8_hvt__vth0_diff_49 = '-2.27750e-03*lvhp_threshold*lvhp_threshold+6.03500e-03*lvhp_threshold+4.81610e-02'
+ sky130_fd_pr__pfet_01v8_hvt__vth0_diff_5 = '-1.51988e-04*lvhp_threshold*lvhp_threshold+-7.21588e-03*lvhp_threshold+-1.28270e-03'
+ sky130_fd_pr__pfet_01v8_hvt__vth0_diff_50 = '-2.81094e-06*lvhp_threshold*lvhp_threshold+1.03083e-02*lvhp_threshold'
+ sky130_fd_pr__pfet_01v8_hvt__vth0_diff_51 = '-1.46084e-03*lvhp_threshold*lvhp_threshold+1.30116e-02*lvhp_threshold'
+ sky130_fd_pr__pfet_01v8_hvt__vth0_diff_52 = '-1.06863e-03*lvhp_threshold*lvhp_threshold+9.01263e-03*lvhp_threshold'
+ sky130_fd_pr__pfet_01v8_hvt__vth0_diff_53 = '-1.21278e-03*lvhp_threshold*lvhp_threshold+1.29531e-02*lvhp_threshold'
+ sky130_fd_pr__pfet_01v8_hvt__vth0_diff_54 = '-2.27750e-03*lvhp_threshold*lvhp_threshold+6.03500e-03*lvhp_threshold'
+ sky130_fd_pr__pfet_01v8_hvt__vth0_diff_55 = '-1.14877e-03*lvhp_threshold*lvhp_threshold+1.09909e-02*lvhp_threshold'
+ sky130_fd_pr__pfet_01v8_hvt__vth0_diff_56 = '-9.18812e-04*lvhp_threshold*lvhp_threshold+-1.93938e-02*lvhp_threshold+2.05860e-02'
+ sky130_fd_pr__pfet_01v8_hvt__vth0_diff_57 = '-1.34041e-03*lvhp_threshold*lvhp_threshold+-6.53501e-03*lvhp_threshold+3.92560e-03'
+ sky130_fd_pr__pfet_01v8_hvt__vth0_diff_58 = '-1.25868e-03*lvhp_threshold*lvhp_threshold+-3.03244e-03*lvhp_threshold+7.57570e-03'
+ sky130_fd_pr__pfet_01v8_hvt__vth0_diff_59 = '-1.99181e-03*lvhp_threshold*lvhp_threshold+4.06675e-03*lvhp_threshold+3.40290e-03'
+ sky130_fd_pr__pfet_01v8_hvt__vth0_diff_6 = '-1.06863e-03*lvhp_threshold*lvhp_threshold+9.01262e-03*lvhp_threshold+-2.02380e-04'
+ sky130_fd_pr__pfet_01v8_hvt__vth0_diff_60 = '-2.27551e-03*lvhp_threshold*lvhp_threshold+4.08075e-03*lvhp_threshold+2.65110e-03'
+ sky130_fd_pr__pfet_01v8_hvt__vth0_diff_61 = '-2.36310e-03*lvhp_threshold*lvhp_threshold+4.18575e-03*lvhp_threshold+1.98360e-03'
+ sky130_fd_pr__pfet_01v8_hvt__vth0_diff_62 = '-2.40726e-03*lvhp_threshold*lvhp_threshold+4.93288e-03*lvhp_threshold+3.62560e-03'
+ sky130_fd_pr__pfet_01v8_hvt__vth0_diff_63 = '-1.97434e-03*lvhp_threshold*lvhp_threshold+2.45750e-03*lvhp_threshold+6.64540e-03'
+ sky130_fd_pr__pfet_01v8_hvt__vth0_diff_64 = '3.74875e-05*lvhp_threshold*lvhp_threshold+-5.75063e-03*lvhp_threshold+-4.39430e-03'
+ sky130_fd_pr__pfet_01v8_hvt__vth0_diff_65 = '2.64581e-04*lvhp_threshold*lvhp_threshold+-1.01461e-02*lvhp_threshold+2.11120e-03'
+ sky130_fd_pr__pfet_01v8_hvt__vth0_diff_66 = '-2.26757e-03*lvhp_threshold*lvhp_threshold+6.00560e-03*lvhp_threshold+3.53550e-03'
+ sky130_fd_pr__pfet_01v8_hvt__vth0_diff_67 = '-1.70992e-03*lvhp_threshold*lvhp_threshold+6.76985e-03*lvhp_threshold+7.20120e-03'
+ sky130_fd_pr__pfet_01v8_hvt__vth0_diff_7 = '-4.19437e-04*lvhp_threshold*lvhp_threshold+8.85450e-03*lvhp_threshold+-1.73090e-02'
+ sky130_fd_pr__pfet_01v8_hvt__vth0_diff_8 = '3.76600e-04*lvhp_threshold*lvhp_threshold+-9.03463e-03*lvhp_threshold+-4.82210e-03'
+ sky130_fd_pr__pfet_01v8_hvt__vth0_diff_9 = '5.18775e-04*lvhp_threshold*lvhp_threshold+-9.03750e-03*lvhp_threshold+8.16600e-04'
+ sky130_fd_pr__pfet_01v8_hvt__wint_diff = '8.04375e-09*diff_cd'
+ sky130_fd_pr__pfet_g5v0d10v5__a0_diff_1 = '5.78513e-04*hvp_saturation*hvp_saturation+2.05655e-03*hvp_saturation+-2.26790e-02'
+ sky130_fd_pr__pfet_g5v0d10v5__a0_diff_10 = '4.09738e-04*hvp_saturation*hvp_saturation+1.26371e-03*hvp_saturation+7.75350e-04'
+ sky130_fd_pr__pfet_g5v0d10v5__a0_diff_14 = '4.81500e-04*hvp_saturation*hvp_saturation+4.85000e-04*hvp_saturation+-2.24290e-02'
+ sky130_fd_pr__pfet_g5v0d10v5__a0_diff_16 = '5.24506e-04*hvp_saturation*hvp_saturation+4.02562e-03*hvp_saturation+-8.79260e-03'
+ sky130_fd_pr__pfet_g5v0d10v5__a0_diff_17 = '8.21006e-04*hvp_saturation*hvp_saturation+3.95717e-03*hvp_saturation+4.21820e-03'
+ sky130_fd_pr__pfet_g5v0d10v5__a0_diff_18 = '3.56503e-04*hvp_saturation*hvp_saturation+1.74664e-03*hvp_saturation+3.12640e-03'
+ sky130_fd_pr__pfet_g5v0d10v5__a0_diff_19 = '-1.47333e-02*hvp_saturation*hvp_saturation+1.85613e-03*hvp_saturation+2.43820e-01'
+ sky130_fd_pr__pfet_g5v0d10v5__a0_diff_22 = '8.44394e-03*hvp_saturation*hvp_saturation+2.98640e-02*hvp_saturation+-2.62690e-02'
+ sky130_fd_pr__pfet_g5v0d10v5__a0_diff_23 = '3.95966e-05*hvp_saturation*hvp_saturation+1.81021e-04*hvp_saturation+3.00570e-04'
+ sky130_fd_pr__pfet_g5v0d10v5__a0_diff_24 = '4.36234e-04*hvp_saturation*hvp_saturation+2.30521e-03*hvp_saturation+3.33540e-03'
+ sky130_fd_pr__pfet_g5v0d10v5__a0_diff_25 = '4.88250e-04*hvp_saturation*hvp_saturation+2.52785e-03*hvp_saturation+1.44360e-03'
+ sky130_fd_pr__pfet_g5v0d10v5__a0_diff_29 = '4.26750e-04*hvp_saturation*hvp_saturation+1.62525e-03*hvp_saturation+-3.05130e-02'
+ sky130_fd_pr__pfet_g5v0d10v5__a0_diff_3 = '1.05056e-03*hvp_saturation*hvp_saturation+-2.35819e-03*hvp_saturation+1.99280e-04'
+ sky130_fd_pr__pfet_g5v0d10v5__a0_diff_30 = '6.09223e-04*hvp_saturation*hvp_saturation+4.14651e-03*hvp_saturation+5.98040e-03'
+ sky130_fd_pr__pfet_g5v0d10v5__a0_diff_31 = '3.15544e-04*hvp_saturation*hvp_saturation+1.91990e-03*hvp_saturation+1.57770e-03'
+ sky130_fd_pr__pfet_g5v0d10v5__a0_diff_32 = '3.73541e-04*hvp_saturation*hvp_saturation+2.14771e-03*hvp_saturation+1.21950e-03'
+ sky130_fd_pr__pfet_g5v0d10v5__a0_diff_4 = '8.29675e-04*hvp_saturation*hvp_saturation+2.03030e-03*hvp_saturation+1.75300e-03'
+ sky130_fd_pr__pfet_g5v0d10v5__a0_diff_5 = '4.73362e-04*hvp_saturation*hvp_saturation+1.67323e-03*hvp_saturation+-1.17170e-03'
+ sky130_fd_pr__pfet_g5v0d10v5__a0_diff_7 = '8.10078e-04*hvp_saturation*hvp_saturation+9.34475e-03*hvp_saturation+5.86760e-04'
+ sky130_fd_pr__pfet_g5v0d10v5__a0_diff_8 = '4.74038e-04*hvp_saturation*hvp_saturation+4.31740e-03*hvp_saturation+-2.27090e-02'
+ sky130_fd_pr__pfet_g5v0d10v5__a0_diff_9 = '8.80753e-04*hvp_saturation*hvp_saturation+2.72849e-03*hvp_saturation+1.55500e-03'
+ sky130_fd_pr__pfet_g5v0d10v5__ags_diff_1 = '-3.03594e-04*hvp_saturation*hvp_saturation+-2.99037e-03*hvp_saturation+-4.20280e-02'
+ sky130_fd_pr__pfet_g5v0d10v5__ags_diff_10 = '-6.48438e-05*hvp_saturation*hvp_saturation+4.89462e-03*hvp_saturation+4.76400e-03'
+ sky130_fd_pr__pfet_g5v0d10v5__ags_diff_14 = '-6.54187e-04*hvp_saturation*hvp_saturation+-6.73500e-03*hvp_saturation+-4.34710e-02'
+ sky130_fd_pr__pfet_g5v0d10v5__ags_diff_16 = '-7.11812e-04*hvp_saturation*hvp_saturation+5.90000e-05*hvp_saturation+-1.91380e-02'
+ sky130_fd_pr__pfet_g5v0d10v5__ags_diff_17 = '-1.09068e-04*hvp_saturation*hvp_saturation+2.94213e-03*hvp_saturation+3.02590e-04'
+ sky130_fd_pr__pfet_g5v0d10v5__ags_diff_18 = '-1.05012e-04*hvp_saturation*hvp_saturation+2.80050e-04*hvp_saturation+-6.78520e-03'
+ sky130_fd_pr__pfet_g5v0d10v5__ags_diff_19 = '-1.80150e-03*hvp_saturation*hvp_saturation+9.38025e-04*hvp_saturation+2.75640e-02'
+ sky130_fd_pr__pfet_g5v0d10v5__ags_diff_22 = '-2.27850e-03*hvp_saturation*hvp_saturation+-1.65165e-02*hvp_saturation+-4.67880e-02'
+ sky130_fd_pr__pfet_g5v0d10v5__ags_diff_23 = '-2.02259e-04*hvp_saturation*hvp_saturation+9.37563e-04*hvp_saturation+3.18860e-03'
+ sky130_fd_pr__pfet_g5v0d10v5__ags_diff_24 = '-6.36094e-05*hvp_saturation*hvp_saturation+-7.71788e-04*hvp_saturation+-5.51890e-03'
+ sky130_fd_pr__pfet_g5v0d10v5__ags_diff_25 = '-8.68219e-05*hvp_saturation*hvp_saturation+-9.84938e-04*hvp_saturation+1.72630e-03'
+ sky130_fd_pr__pfet_g5v0d10v5__ags_diff_29 = '-6.50969e-04*hvp_saturation*hvp_saturation+-3.68637e-03*hvp_saturation+-5.36940e-02'
+ sky130_fd_pr__pfet_g5v0d10v5__ags_diff_3 = '-1.12594e-04*hvp_saturation*hvp_saturation+1.73526e-02*hvp_saturation+1.69100e-03'
+ sky130_fd_pr__pfet_g5v0d10v5__ags_diff_30 = '-1.24188e-04*hvp_saturation*hvp_saturation+9.35200e-04*hvp_saturation+9.21620e-03'
+ sky130_fd_pr__pfet_g5v0d10v5__ags_diff_31 = '-1.06362e-04*hvp_saturation*hvp_saturation+-1.78722e-03*hvp_saturation+2.53720e-03'
+ sky130_fd_pr__pfet_g5v0d10v5__ags_diff_32 = '-8.52219e-05*hvp_saturation*hvp_saturation+-1.44499e-03*hvp_saturation+2.47340e-03'
+ sky130_fd_pr__pfet_g5v0d10v5__ags_diff_4 = '-5.51139e-05*hvp_saturation*hvp_saturation+7.56100e-03*hvp_saturation+5.38230e-05'
+ sky130_fd_pr__pfet_g5v0d10v5__ags_diff_5 = '-9.71131e-05*hvp_saturation*hvp_saturation+3.04770e-03*hvp_saturation+1.39070e-02'
+ sky130_fd_pr__pfet_g5v0d10v5__ags_diff_7 = '-1.18200e-03*hvp_saturation*hvp_saturation+7.06005e-03*hvp_saturation+-3.17570e-05'
+ sky130_fd_pr__pfet_g5v0d10v5__ags_diff_8 = '-6.87656e-04*hvp_saturation*hvp_saturation+7.57375e-04*hvp_saturation+-3.95060e-02'
+ sky130_fd_pr__pfet_g5v0d10v5__ags_diff_9 = '-1.37375e-05*hvp_saturation*hvp_saturation+6.61250e-03*hvp_saturation+1.34780e-03'
+ sky130_fd_pr__pfet_g5v0d10v5__ajunction_mult = '-2.50000e-06*hvp_diode*hvp_diode+1.81850e-02*hvp_diode+1.00500e+00'
+ sky130_fd_pr__pfet_g5v0d10v5__b0_diff_35 = '-1.24613e-08*hvp_saturation*hvp_saturation+-7.01645e-08*hvp_saturation+-1.99310e-08'
+ sky130_fd_pr__pfet_g5v0d10v5__b0_diff_36 = '-1.27834e-09*hvp_saturation*hvp_saturation+-1.53426e-08*hvp_saturation+-1.72900e-08'
+ sky130_fd_pr__pfet_g5v0d10v5__b0_diff_37 = '4.14719e-10*hvp_saturation*hvp_saturation+-1.78901e-08*hvp_saturation+-1.06550e-08'
+ sky130_fd_pr__pfet_g5v0d10v5__b0_diff_38 = '-2.95000e-10*hvp_saturation*hvp_saturation+-1.45738e-08*hvp_saturation+1.30150e-08'
+ sky130_fd_pr__pfet_g5v0d10v5__b0_diff_39 = '2.67594e-10*hvp_saturation*hvp_saturation+-1.33869e-08*hvp_saturation+6.02300e-09'
+ sky130_fd_pr__pfet_g5v0d10v5__b0_diff_43 = '1.71694e-09*hvp_saturation*hvp_saturation+-3.01300e-08*hvp_saturation+8.99490e-08'
+ sky130_fd_pr__pfet_g5v0d10v5__b0_diff_44 = '1.22287e-09*hvp_saturation*hvp_saturation+-1.62662e-08*hvp_saturation+6.67090e-08'
+ sky130_fd_pr__pfet_g5v0d10v5__b0_diff_45 = '-2.12413e-10*hvp_saturation*hvp_saturation+-2.35773e-08*hvp_saturation+2.85760e-09'
+ sky130_fd_pr__pfet_g5v0d10v5__b1_diff_35 = '1.01576e-07*hvp_saturation*hvp_saturation+4.19222e-07*hvp_saturation+5.29010e-08'
+ sky130_fd_pr__pfet_g5v0d10v5__b1_diff_36 = '1.55838e-08*hvp_saturation*hvp_saturation+6.23693e-08*hvp_saturation+1.18150e-09'
+ sky130_fd_pr__pfet_g5v0d10v5__b1_diff_37 = '2.79198e-09*hvp_saturation*hvp_saturation+-3.15975e-09*hvp_saturation+6.84530e-09'
+ sky130_fd_pr__pfet_g5v0d10v5__b1_diff_38 = '1.79298e-08*hvp_saturation*hvp_saturation+7.16693e-08*hvp_saturation+6.67620e-09'
+ sky130_fd_pr__pfet_g5v0d10v5__b1_diff_39 = '1.16331e-08*hvp_saturation*hvp_saturation+2.80474e-08*hvp_saturation+4.50410e-10'
+ sky130_fd_pr__pfet_g5v0d10v5__b1_diff_43 = '-1.55723e-08*hvp_saturation*hvp_saturation+-6.21021e-08*hvp_saturation+1.03500e-09'
+ sky130_fd_pr__pfet_g5v0d10v5__b1_diff_44 = '7.82657e-09*hvp_saturation*hvp_saturation+3.13162e-08*hvp_saturation+3.90100e-10'
+ sky130_fd_pr__pfet_g5v0d10v5__b1_diff_45 = '1.03807e-08*hvp_saturation*hvp_saturation+4.14538e-08*hvp_saturation+3.29820e-11'
+ sky130_fd_pr__pfet_g5v0d10v5__dlc_diff = '-4.33125e-09*poly_cd'
+ sky130_fd_pr__pfet_g5v0d10v5__dwc_diff = '8.04375e-09*diff_cd'
+ sky130_fd_pr__pfet_g5v0d10v5__k2_diff_0 = '6.33750e-05*hvp_bodyeffect*hvp_bodyeffect+-8.87000e-04*hvp_bodyeffect+1.47030e-02'
+ sky130_fd_pr__pfet_g5v0d10v5__k2_diff_1 = '-3.51219e-05*hvp_bodyeffect*hvp_bodyeffect+1.12199e-03*hvp_bodyeffect+1.30830e-02'
+ sky130_fd_pr__pfet_g5v0d10v5__k2_diff_10 = '1.51250e-06*hvp_bodyeffect*hvp_bodyeffect+3.67575e-04*hvp_bodyeffect+4.75430e-03'
+ sky130_fd_pr__pfet_g5v0d10v5__k2_diff_11 = '8.53312e-05*hvp_bodyeffect*hvp_bodyeffect+-1.97417e-03*hvp_bodyeffect+1.00500e-02'
+ sky130_fd_pr__pfet_g5v0d10v5__k2_diff_12 = '3.28969e-05*hvp_bodyeffect*hvp_bodyeffect+-1.24881e-03*hvp_bodyeffect+6.41540e-03'
+ sky130_fd_pr__pfet_g5v0d10v5__k2_diff_13 = '1.02781e-05*hvp_bodyeffect*hvp_bodyeffect+-4.23388e-04*hvp_bodyeffect+1.07680e-02'
+ sky130_fd_pr__pfet_g5v0d10v5__k2_diff_14 = '-1.20000e-05*hvp_bodyeffect*hvp_bodyeffect+1.06050e-03*hvp_bodyeffect+1.29450e-02'
+ sky130_fd_pr__pfet_g5v0d10v5__k2_diff_15 = '6.46875e-05*hvp_bodyeffect*hvp_bodyeffect+-7.73250e-04*hvp_bodyeffect+1.42500e-02'
+ sky130_fd_pr__pfet_g5v0d10v5__k2_diff_16 = '-2.78125e-06*hvp_bodyeffect*hvp_bodyeffect+7.32875e-04*hvp_bodyeffect+1.17840e-02'
+ sky130_fd_pr__pfet_g5v0d10v5__k2_diff_17 = '-3.59844e-05*hvp_bodyeffect*hvp_bodyeffect+8.13563e-04*hvp_bodyeffect+5.43680e-03'
+ sky130_fd_pr__pfet_g5v0d10v5__k2_diff_18 = '-1.09000e-05*hvp_bodyeffect*hvp_bodyeffect+7.91200e-04*hvp_bodyeffect+6.33700e-03'
+ sky130_fd_pr__pfet_g5v0d10v5__k2_diff_19 = '-3.53544e-05*hvp_bodyeffect*hvp_bodyeffect+9.49092e-04*hvp_bodyeffect+5.02710e-03'
+ sky130_fd_pr__pfet_g5v0d10v5__k2_diff_2 = '7.31875e-05*hvp_bodyeffect*hvp_bodyeffect+-1.36875e-03*hvp_bodyeffect+1.41510e-02'
+ sky130_fd_pr__pfet_g5v0d10v5__k2_diff_20 = '8.37812e-05*hvp_bodyeffect*hvp_bodyeffect+-1.24787e-03*hvp_bodyeffect+1.41840e-02'
+ sky130_fd_pr__pfet_g5v0d10v5__k2_diff_21 = '1.15937e-05*hvp_bodyeffect*hvp_bodyeffect+-1.93125e-04*hvp_bodyeffect+1.45130e-02'
+ sky130_fd_pr__pfet_g5v0d10v5__k2_diff_22 = '-2.60156e-05*hvp_bodyeffect*hvp_bodyeffect+1.53956e-03*hvp_bodyeffect+1.05890e-02'
+ sky130_fd_pr__pfet_g5v0d10v5__k2_diff_23 = '-2.15025e-05*hvp_bodyeffect*hvp_bodyeffect+1.21979e-03*hvp_bodyeffect+5.53490e-03'
+ sky130_fd_pr__pfet_g5v0d10v5__k2_diff_24 = '-1.84687e-06*hvp_bodyeffect*hvp_bodyeffect+8.45737e-04*hvp_bodyeffect+7.01160e-03'
+ sky130_fd_pr__pfet_g5v0d10v5__k2_diff_25 = '-1.42853e-05*hvp_bodyeffect*hvp_bodyeffect+1.10767e-03*hvp_bodyeffect+5.18560e-03'
+ sky130_fd_pr__pfet_g5v0d10v5__k2_diff_26 = '5.01875e-05*hvp_bodyeffect*hvp_bodyeffect+-6.96250e-04*hvp_bodyeffect+1.22900e-02'
+ sky130_fd_pr__pfet_g5v0d10v5__k2_diff_27 = '2.20000e-05*hvp_bodyeffect*hvp_bodyeffect+-1.98000e-04*hvp_bodyeffect+1.42390e-02'
+ sky130_fd_pr__pfet_g5v0d10v5__k2_diff_28 = '-7.35000e-06*hvp_bodyeffect*hvp_bodyeffect+6.94400e-04*hvp_bodyeffect+1.03000e-02'
+ sky130_fd_pr__pfet_g5v0d10v5__k2_diff_29 = '-1.17187e-05*hvp_bodyeffect*hvp_bodyeffect+9.81625e-04*hvp_bodyeffect+1.27370e-02'
+ sky130_fd_pr__pfet_g5v0d10v5__k2_diff_3 = '1.21875e-06*hvp_bodyeffect*hvp_bodyeffect+6.34400e-04*hvp_bodyeffect+5.73650e-03'
+ sky130_fd_pr__pfet_g5v0d10v5__k2_diff_30 = '-2.09441e-05*hvp_bodyeffect*hvp_bodyeffect+1.21325e-03*hvp_bodyeffect+5.96010e-03'
+ sky130_fd_pr__pfet_g5v0d10v5__k2_diff_31 = '-2.03063e-05*hvp_bodyeffect*hvp_bodyeffect+1.01465e-03*hvp_bodyeffect+7.34130e-03'
+ sky130_fd_pr__pfet_g5v0d10v5__k2_diff_32 = '-2.27006e-05*hvp_bodyeffect*hvp_bodyeffect+1.13043e-03*hvp_bodyeffect+5.35340e-03'
+ sky130_fd_pr__pfet_g5v0d10v5__k2_diff_33 = '5.46250e-05*hvp_bodyeffect*hvp_bodyeffect+-9.52250e-04*hvp_bodyeffect+1.48030e-02'
+ sky130_fd_pr__pfet_g5v0d10v5__k2_diff_34 = '-1.30062e-05*hvp_bodyeffect*hvp_bodyeffect+6.05275e-04*hvp_bodyeffect+1.06530e-02'
+ sky130_fd_pr__pfet_g5v0d10v5__k2_diff_35 = '1.31284e-04*hvp_bodyeffect*hvp_bodyeffect+4.95288e-04*hvp_bodyeffect+3.44010e-03'
+ sky130_fd_pr__pfet_g5v0d10v5__k2_diff_36 = '-4.35184e-05*hvp_bodyeffect*hvp_bodyeffect+7.99899e-04*hvp_bodyeffect+3.63810e-03'
+ sky130_fd_pr__pfet_g5v0d10v5__k2_diff_37 = '-2.13219e-05*hvp_bodyeffect*hvp_bodyeffect+1.36300e-04*hvp_bodyeffect+-4.59550e-04'
+ sky130_fd_pr__pfet_g5v0d10v5__k2_diff_38 = '-1.31797e-05*hvp_bodyeffect*hvp_bodyeffect+4.99269e-04*hvp_bodyeffect+2.23250e-03'
+ sky130_fd_pr__pfet_g5v0d10v5__k2_diff_39 = '-4.22500e-06*hvp_bodyeffect*hvp_bodyeffect+4.32450e-04*hvp_bodyeffect+3.54350e-03'
+ sky130_fd_pr__pfet_g5v0d10v5__k2_diff_4 = '-2.97812e-06*hvp_bodyeffect*hvp_bodyeffect+4.71712e-04*hvp_bodyeffect+4.60610e-03'
+ sky130_fd_pr__pfet_g5v0d10v5__k2_diff_40 = '6.11406e-05*hvp_bodyeffect*hvp_bodyeffect+-4.57494e-03*hvp_bodyeffect+1.20330e-02'
+ sky130_fd_pr__pfet_g5v0d10v5__k2_diff_41 = '8.07813e-06*hvp_bodyeffect*hvp_bodyeffect+-2.39114e-03*hvp_bodyeffect+3.89520e-03'
+ sky130_fd_pr__pfet_g5v0d10v5__k2_diff_42 = '3.91250e-06*hvp_bodyeffect*hvp_bodyeffect+-1.29688e-03*hvp_bodyeffect+8.06790e-03'
+ sky130_fd_pr__pfet_g5v0d10v5__k2_diff_43 = '-3.84375e-07*hvp_bodyeffect*hvp_bodyeffect+2.20062e-04*hvp_bodyeffect+8.81360e-03'
+ sky130_fd_pr__pfet_g5v0d10v5__k2_diff_44 = '2.81250e-07*hvp_bodyeffect*hvp_bodyeffect+-1.30400e-04*hvp_bodyeffect+8.38500e-03'
+ sky130_fd_pr__pfet_g5v0d10v5__k2_diff_45 = '3.12500e-06*hvp_bodyeffect*hvp_bodyeffect+-1.04500e-05*hvp_bodyeffect+5.25730e-03'
+ sky130_fd_pr__pfet_g5v0d10v5__k2_diff_46 = '8.35938e-05*hvp_bodyeffect*hvp_bodyeffect+-2.67263e-03*hvp_bodyeffect+1.14890e-02'
+ sky130_fd_pr__pfet_g5v0d10v5__k2_diff_47 = '3.65625e-06*hvp_bodyeffect*hvp_bodyeffect+5.28750e-05*hvp_bodyeffect+1.15670e-02'
+ sky130_fd_pr__pfet_g5v0d10v5__k2_diff_48 = '2.11062e-05*hvp_bodyeffect*hvp_bodyeffect+-8.54225e-04*hvp_bodyeffect+7.47340e-03'
+ sky130_fd_pr__pfet_g5v0d10v5__k2_diff_5 = '-5.60312e-06*hvp_bodyeffect*hvp_bodyeffect+4.84438e-04*hvp_bodyeffect+6.73600e-03'
+ sky130_fd_pr__pfet_g5v0d10v5__k2_diff_6 = '7.83125e-05*hvp_bodyeffect*hvp_bodyeffect+-1.64875e-03*hvp_bodyeffect+1.11930e-02'
+ sky130_fd_pr__pfet_g5v0d10v5__k2_diff_7 = '8.68125e-06*hvp_bodyeffect*hvp_bodyeffect+1.46475e-04*hvp_bodyeffect+8.91590e-03'
+ sky130_fd_pr__pfet_g5v0d10v5__k2_diff_8 = '1.60312e-06*hvp_bodyeffect*hvp_bodyeffect+1.07938e-04*hvp_bodyeffect+7.16650e-03'
+ sky130_fd_pr__pfet_g5v0d10v5__k2_diff_9 = '-2.30937e-06*hvp_bodyeffect*hvp_bodyeffect+2.54538e-04*hvp_bodyeffect+3.59520e-03'
+ sky130_fd_pr__pfet_g5v0d10v5__lint_diff = '-4.33125e-09*poly_cd'
+ sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_0 = '7.10000e-04*hvp_subvt*hvp_subvt+-8.33875e-02*hvp_subvt+5.77880e-01'
+ sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_1 = '2.82938e-03*hvp_subvt*hvp_subvt+-6.85500e-03*hvp_subvt+2.83000e-01'
+ sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_10 = '1.13188e-03*hvp_subvt*hvp_subvt+-2.45700e-02*hvp_subvt+6.50790e-01'
+ sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_11 = '9.07187e-05*hvp_subvt*hvp_subvt+-1.12317e-01*hvp_subvt+3.59520e-01'
+ sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_12 = '1.21334e-03*hvp_subvt*hvp_subvt+-4.81591e-02*hvp_subvt+2.14700e-01'
+ sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_13 = '1.24900e-03*hvp_subvt*hvp_subvt+-6.13338e-02*hvp_subvt+8.42510e-02'
+ sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_14 = '1.17187e-04*hvp_subvt*hvp_subvt+-8.89375e-03*hvp_subvt+2.53290e-01'
+ sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_15 = '2.03063e-04*hvp_subvt*hvp_subvt+-9.54003e-02*hvp_subvt+4.68090e-01'
+ sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_16 = '9.17500e-04*hvp_subvt*hvp_subvt+-2.96900e-02*hvp_subvt+3.63090e-01'
+ sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_17 = '5.83053e-03*hvp_subvt*hvp_subvt+-2.37339e-02*hvp_subvt+-3.55140e-02'
+ sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_18 = '6.57500e-04*hvp_subvt*hvp_subvt+-1.66600e-02*hvp_subvt+9.45840e-01'
+ sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_19 = '1.31750e-03*hvp_subvt*hvp_subvt+-1.33900e-02*hvp_subvt+6.54750e-01'
+ sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_2 = '7.60625e-04*hvp_subvt*hvp_subvt+1.84475e-02*hvp_subvt+5.01840e-01'
+ sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_20 = '-1.04219e-03*hvp_subvt*hvp_subvt+-1.32849e-01*hvp_subvt+4.09960e-01'
+ sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_21 = '1.01769e-03*hvp_subvt*hvp_subvt+-6.14568e-02*hvp_subvt+2.69400e-01'
+ sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_22 = '1.56531e-03*hvp_subvt*hvp_subvt+7.97875e-03*hvp_subvt+2.60220e-01'
+ sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_24 = '-1.24687e-04*hvp_subvt*hvp_subvt+-2.46588e-02*hvp_subvt+9.57160e-01'
+ sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_25 = '2.68438e-04*hvp_subvt*hvp_subvt+-9.88875e-03*hvp_subvt+6.81510e-01'
+ sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_27 = '8.93562e-04*hvp_subvt*hvp_subvt+-7.16583e-02*hvp_subvt+2.10740e-01'
+ sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_28 = '7.97750e-04*hvp_subvt*hvp_subvt+-2.93015e-02*hvp_subvt+1.93250e-01'
+ sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_29 = '3.39687e-04*hvp_subvt*hvp_subvt+-2.60037e-02*hvp_subvt+3.59730e-01'
+ sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_3 = '6.85312e-04*hvp_subvt*hvp_subvt+-2.99537e-02*hvp_subvt+3.88500e-01'
+ sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_30 = '1.07116e-03*hvp_subvt*hvp_subvt+-9.58662e-03*hvp_subvt+7.27250e-02'
+ sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_31 = '3.78125e-04*hvp_subvt*hvp_subvt+-1.59825e-02*hvp_subvt+9.24650e-01'
+ sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_32 = '5.88437e-04*hvp_subvt*hvp_subvt+-1.24587e-02*hvp_subvt+6.55190e-01'
+ sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_33 = '9.24063e-04*hvp_subvt*hvp_subvt+-7.08488e-02*hvp_subvt+5.75900e-01'
+ sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_34 = '8.73875e-04*hvp_subvt*hvp_subvt+-4.34520e-02*hvp_subvt+1.77380e-01'
+ sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_35 = '-1.43688e-03*hvp_subvt*hvp_subvt+1.71150e-02*hvp_subvt+3.32760e-01'
+ sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_36 = '2.76875e-03*hvp_subvt*hvp_subvt+1.01250e-02*hvp_subvt+1.00310e+00'
+ sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_37 = '-1.54406e-03*hvp_subvt*hvp_subvt+-5.67125e-03*hvp_subvt+2.94850e-01'
+ sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_38 = '5.23000e-03*hvp_subvt*hvp_subvt+2.48175e-02*hvp_subvt+2.56100e-01'
+ sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_39 = '2.51875e-03*hvp_subvt*hvp_subvt+-6.81250e-03*hvp_subvt+5.71760e-01'
+ sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_4 = '4.26562e-04*hvp_subvt*hvp_subvt+-1.66287e-02*hvp_subvt+4.65990e-01'
+ sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_40 = '2.57813e-03*hvp_subvt*hvp_subvt+-1.18835e-01*hvp_subvt+1.99470e-01'
+ sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_42 = '1.02844e-03*hvp_subvt*hvp_subvt+-1.29444e-01*hvp_subvt+2.96520e-01'
+ sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_43 = '1.49618e-03*hvp_subvt*hvp_subvt+-5.29453e-02*hvp_subvt+1.94480e-01'
+ sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_44 = '1.20844e-03*hvp_subvt*hvp_subvt+-3.21862e-02*hvp_subvt+3.16280e-01'
+ sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_45 = '1.07469e-03*hvp_subvt*hvp_subvt+-4.16737e-02*hvp_subvt+5.92520e-01'
+ sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_46 = '3.78312e-04*hvp_subvt*hvp_subvt+-1.44914e-01*hvp_subvt+7.36020e-02'
+ sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_47 = '1.47816e-03*hvp_subvt*hvp_subvt+-5.79799e-02*hvp_subvt+1.90950e-01'
+ sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_5 = '5.94687e-04*hvp_subvt*hvp_subvt+-1.90637e-02*hvp_subvt+5.43860e-01'
+ sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_6 = '8.94594e-04*hvp_subvt*hvp_subvt+-8.16266e-02*hvp_subvt+2.87440e-01'
+ sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_7 = '8.10625e-04*hvp_subvt*hvp_subvt+-4.47600e-02*hvp_subvt+3.34010e-01'
+ sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_8 = '9.49375e-04*hvp_subvt*hvp_subvt+-3.01950e-02*hvp_subvt+3.90000e-01'
+ sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_9 = '1.19969e-03*hvp_subvt*hvp_subvt+-2.33363e-02*hvp_subvt+6.67710e-01'
+ sky130_fd_pr__pfet_g5v0d10v5__overlap_mult = '8.68750e-04*hvtox*hvtox+7.40000e-02*hvtox+9.82100e-01'
+ sky130_fd_pr__pfet_g5v0d10v5__pjunction_mult = '-1.25000e-06*hvp_diode*hvp_diode+1.61550e-02*hvp_diode+1.00900e+00'
+ sky130_fd_pr__pfet_g5v0d10v5__toxe_mult = '1.50000e-02*hvtox+1.00000e+00'
+ sky130_fd_pr__pfet_g5v0d10v5__u0_diff_0 = '-1.59434e-05*hvp_mobility*hvp_mobility+1.97826e-04*hvp_mobility+-1.41240e-03'
+ sky130_fd_pr__pfet_g5v0d10v5__u0_diff_1 = '-1.78206e-05*hvp_mobility*hvp_mobility+-1.92167e-04*hvp_mobility+-1.40110e-03'
+ sky130_fd_pr__pfet_g5v0d10v5__u0_diff_10 = '-8.11000e-06*hvp_mobility*hvp_mobility+8.70125e-05*hvp_mobility+-5.87390e-04'
+ sky130_fd_pr__pfet_g5v0d10v5__u0_diff_11 = '-1.18994e-05*hvp_mobility*hvp_mobility+3.29575e-04*hvp_mobility+-3.97810e-04'
+ sky130_fd_pr__pfet_g5v0d10v5__u0_diff_12 = '1.76747e-05*hvp_mobility*hvp_mobility+3.56299e-04*hvp_mobility+-1.96720e-03'
+ sky130_fd_pr__pfet_g5v0d10v5__u0_diff_13 = '-9.20938e-06*hvp_mobility*hvp_mobility+2.15863e-04*hvp_mobility+-1.04820e-03'
+ sky130_fd_pr__pfet_g5v0d10v5__u0_diff_14 = '-5.31562e-06*hvp_mobility*hvp_mobility+6.61875e-05*hvp_mobility+-1.21490e-03'
+ sky130_fd_pr__pfet_g5v0d10v5__u0_diff_15 = '-1.56434e-05*hvp_mobility*hvp_mobility+2.37151e-04*hvp_mobility+-1.59630e-03'
+ sky130_fd_pr__pfet_g5v0d10v5__u0_diff_16 = '-8.38750e-06*hvp_mobility*hvp_mobility+9.33250e-05*hvp_mobility+-2.04100e-03'
+ sky130_fd_pr__pfet_g5v0d10v5__u0_diff_17 = '-9.12656e-06*hvp_mobility*hvp_mobility+4.10937e-05*hvp_mobility+-3.78080e-04'
+ sky130_fd_pr__pfet_g5v0d10v5__u0_diff_18 = '-1.02031e-05*hvp_mobility*hvp_mobility+-9.66250e-06*hvp_mobility+-2.00890e-03'
+ sky130_fd_pr__pfet_g5v0d10v5__u0_diff_19 = '-3.20938e-06*hvp_mobility*hvp_mobility+-1.68625e-05*hvp_mobility+-1.46800e-03'
+ sky130_fd_pr__pfet_g5v0d10v5__u0_diff_2 = '-1.72594e-05*hvp_mobility*hvp_mobility+8.46625e-05*hvp_mobility+-1.57910e-03'
+ sky130_fd_pr__pfet_g5v0d10v5__u0_diff_20 = '-1.90228e-05*hvp_mobility*hvp_mobility+3.07901e-04*hvp_mobility+-5.76630e-04'
+ sky130_fd_pr__pfet_g5v0d10v5__u0_diff_21 = '-1.17188e-05*hvp_mobility*hvp_mobility+1.94300e-04*hvp_mobility+-2.24180e-03'
+ sky130_fd_pr__pfet_g5v0d10v5__u0_diff_22 = '-1.82347e-05*hvp_mobility*hvp_mobility+-1.45786e-04*hvp_mobility+-4.01900e-04'
+ sky130_fd_pr__pfet_g5v0d10v5__u0_diff_23 = '-1.05431e-05*hvp_mobility*hvp_mobility+-1.68750e-06*hvp_mobility+-9.95960e-04'
+ sky130_fd_pr__pfet_g5v0d10v5__u0_diff_24 = '-6.62812e-06*hvp_mobility*hvp_mobility+4.27625e-05*hvp_mobility+-2.23220e-03'
+ sky130_fd_pr__pfet_g5v0d10v5__u0_diff_25 = '-6.88750e-06*hvp_mobility*hvp_mobility+-9.50000e-06*hvp_mobility+-1.98880e-03'
+ sky130_fd_pr__pfet_g5v0d10v5__u0_diff_26 = '-1.70244e-05*hvp_mobility*hvp_mobility+1.97652e-04*hvp_mobility+-1.23390e-03'
+ sky130_fd_pr__pfet_g5v0d10v5__u0_diff_27 = '-1.90406e-05*hvp_mobility*hvp_mobility+2.39862e-04*hvp_mobility+-3.53360e-03'
+ sky130_fd_pr__pfet_g5v0d10v5__u0_diff_28 = '-9.33750e-06*hvp_mobility*hvp_mobility+1.14275e-04*hvp_mobility+-2.68450e-03'
+ sky130_fd_pr__pfet_g5v0d10v5__u0_diff_29 = '-5.73125e-06*hvp_mobility*hvp_mobility+1.04825e-04*hvp_mobility+-1.46420e-03'
+ sky130_fd_pr__pfet_g5v0d10v5__u0_diff_3 = '-1.25606e-05*hvp_mobility*hvp_mobility+7.71575e-05*hvp_mobility+-7.05500e-04'
+ sky130_fd_pr__pfet_g5v0d10v5__u0_diff_30 = '-7.65312e-06*hvp_mobility*hvp_mobility+-5.46250e-06*hvp_mobility+-1.02120e-03'
+ sky130_fd_pr__pfet_g5v0d10v5__u0_diff_31 = '-7.79687e-06*hvp_mobility*hvp_mobility+5.96250e-06*hvp_mobility+-2.29940e-03'
+ sky130_fd_pr__pfet_g5v0d10v5__u0_diff_32 = '-6.84063e-06*hvp_mobility*hvp_mobility+-1.91875e-05*hvp_mobility+-1.91440e-03'
+ sky130_fd_pr__pfet_g5v0d10v5__u0_diff_33 = '-1.43656e-05*hvp_mobility*hvp_mobility+2.51562e-04*hvp_mobility+-1.80920e-03'
+ sky130_fd_pr__pfet_g5v0d10v5__u0_diff_34 = '-7.60937e-06*hvp_mobility*hvp_mobility+1.70913e-04*hvp_mobility+-2.82760e-03'
+ sky130_fd_pr__pfet_g5v0d10v5__u0_diff_35 = '-6.11103e-05*hvp_mobility*hvp_mobility+-5.49819e-04*hvp_mobility+-3.82760e-04'
+ sky130_fd_pr__pfet_g5v0d10v5__u0_diff_36 = '-2.51965e-05*hvp_mobility*hvp_mobility+-1.28891e-04*hvp_mobility+-1.67690e-04'
+ sky130_fd_pr__pfet_g5v0d10v5__u0_diff_37 = '-3.66013e-05*hvp_mobility*hvp_mobility+-2.53900e-04*hvp_mobility+5.61320e-04'
+ sky130_fd_pr__pfet_g5v0d10v5__u0_diff_38 = '-2.90391e-05*hvp_mobility*hvp_mobility+-1.04189e-04*hvp_mobility+7.08030e-04'
+ sky130_fd_pr__pfet_g5v0d10v5__u0_diff_39 = '-2.38741e-05*hvp_mobility*hvp_mobility+-5.48112e-05*hvp_mobility+-2.40140e-04'
+ sky130_fd_pr__pfet_g5v0d10v5__u0_diff_4 = '-8.11281e-06*hvp_mobility*hvp_mobility+7.12463e-05*hvp_mobility+-5.49120e-04'
+ sky130_fd_pr__pfet_g5v0d10v5__u0_diff_40 = '-5.35219e-05*hvp_mobility*hvp_mobility+2.90125e-05*hvp_mobility+-3.31020e-03'
+ sky130_fd_pr__pfet_g5v0d10v5__u0_diff_41 = '-4.55813e-05*hvp_mobility*hvp_mobility+-8.62475e-05*hvp_mobility+5.42130e-04'
+ sky130_fd_pr__pfet_g5v0d10v5__u0_diff_42 = '-4.59456e-05*hvp_mobility*hvp_mobility+-1.91125e-05*hvp_mobility+-7.49220e-04'
+ sky130_fd_pr__pfet_g5v0d10v5__u0_diff_43 = '-1.98313e-05*hvp_mobility*hvp_mobility+2.50250e-05*hvp_mobility+-1.64690e-03'
+ sky130_fd_pr__pfet_g5v0d10v5__u0_diff_44 = '-1.40594e-05*hvp_mobility*hvp_mobility+-9.12500e-07*hvp_mobility+-2.18650e-03'
+ sky130_fd_pr__pfet_g5v0d10v5__u0_diff_45 = '-5.70719e-06*hvp_mobility*hvp_mobility+5.42262e-05*hvp_mobility+-9.62880e-04'
+ sky130_fd_pr__pfet_g5v0d10v5__u0_diff_46 = '-1.67122e-05*hvp_mobility*hvp_mobility+3.38401e-04*hvp_mobility+-1.78270e-03'
+ sky130_fd_pr__pfet_g5v0d10v5__u0_diff_47 = '-1.85938e-05*hvp_mobility*hvp_mobility+9.23250e-05*hvp_mobility+-2.42490e-03'
+ sky130_fd_pr__pfet_g5v0d10v5__u0_diff_48 = '-2.12809e-05*hvp_mobility*hvp_mobility+1.05744e-04*hvp_mobility+3.59190e-04'
+ sky130_fd_pr__pfet_g5v0d10v5__u0_diff_5 = '-7.41875e-06*hvp_mobility*hvp_mobility+6.32250e-05*hvp_mobility+-1.50510e-03'
+ sky130_fd_pr__pfet_g5v0d10v5__u0_diff_6 = '-8.64500e-06*hvp_mobility*hvp_mobility+3.42245e-04*hvp_mobility+-1.94100e-03'
+ sky130_fd_pr__pfet_g5v0d10v5__u0_diff_7 = '-8.63375e-06*hvp_mobility*hvp_mobility+1.05445e-04*hvp_mobility+-8.12580e-04'
+ sky130_fd_pr__pfet_g5v0d10v5__u0_diff_8 = '-1.02312e-05*hvp_mobility*hvp_mobility+5.20750e-05*hvp_mobility+-1.08730e-03'
+ sky130_fd_pr__pfet_g5v0d10v5__u0_diff_9 = '-7.61906e-06*hvp_mobility*hvp_mobility+7.68212e-05*hvp_mobility+-6.45410e-04'
+ sky130_fd_pr__pfet_g5v0d10v5__ua_diff_0 = '2.06314e-12*hvp_mobility*hvp_mobility+8.38543e-12*hvp_mobility+-5.80220e-14'
+ sky130_fd_pr__pfet_g5v0d10v5__ua_diff_1 = '1.89620e-12*hvp_mobility*hvp_mobility+7.42031e-12*hvp_mobility+6.76490e-13'
+ sky130_fd_pr__pfet_g5v0d10v5__ua_diff_10 = '6.61409e-13*hvp_mobility*hvp_mobility+2.48603e-12*hvp_mobility+-2.62680e-13'
+ sky130_fd_pr__pfet_g5v0d10v5__ua_diff_11 = '2.31099e-12*hvp_mobility*hvp_mobility+1.30790e-11*hvp_mobility+1.61980e-11'
+ sky130_fd_pr__pfet_g5v0d10v5__ua_diff_12 = '1.56844e-11*hvp_mobility*hvp_mobility+6.26056e-11*hvp_mobility+-1.37290e-12'
+ sky130_fd_pr__pfet_g5v0d10v5__ua_diff_13 = '1.84419e-12*hvp_mobility*hvp_mobility+9.74039e-12*hvp_mobility+8.10740e-12'
+ sky130_fd_pr__pfet_g5v0d10v5__ua_diff_14 = '1.94659e-12*hvp_mobility*hvp_mobility+7.98322e-12*hvp_mobility+1.44570e-12'
+ sky130_fd_pr__pfet_g5v0d10v5__ua_diff_15 = '1.83013e-12*hvp_mobility*hvp_mobility+7.47352e-12*hvp_mobility+1.00890e-12'
+ sky130_fd_pr__pfet_g5v0d10v5__ua_diff_16 = '1.85194e-12*hvp_mobility*hvp_mobility+7.10433e-12*hvp_mobility+-7.48320e-13'
+ sky130_fd_pr__pfet_g5v0d10v5__ua_diff_17 = '1.85177e-12*hvp_mobility*hvp_mobility+7.56409e-12*hvp_mobility+2.06640e-12'
+ sky130_fd_pr__pfet_g5v0d10v5__ua_diff_18 = '2.78012e-13*hvp_mobility*hvp_mobility+7.87659e-13*hvp_mobility+-8.48230e-13'
+ sky130_fd_pr__pfet_g5v0d10v5__ua_diff_19 = '4.52236e-12*hvp_mobility*hvp_mobility+3.63107e-12*hvp_mobility+-5.72190e-11'
+ sky130_fd_pr__pfet_g5v0d10v5__ua_diff_2 = '1.88557e-12*hvp_mobility*hvp_mobility+7.56018e-12*hvp_mobility+3.27190e-13'
+ sky130_fd_pr__pfet_g5v0d10v5__ua_diff_20 = '2.01225e-12*hvp_mobility*hvp_mobility+9.77611e-12*hvp_mobility+8.36560e-12'
+ sky130_fd_pr__pfet_g5v0d10v5__ua_diff_21 = '1.80428e-12*hvp_mobility*hvp_mobility+6.83710e-12*hvp_mobility+-2.07690e-12'
+ sky130_fd_pr__pfet_g5v0d10v5__ua_diff_22 = '3.98790e-13*hvp_mobility*hvp_mobility+1.15686e-12*hvp_mobility+5.68910e-13'
+ sky130_fd_pr__pfet_g5v0d10v5__ua_diff_23 = '3.30000e-16*hvp_mobility*hvp_mobility+-2.96037e-13*hvp_mobility+1.09270e-13'
+ sky130_fd_pr__pfet_g5v0d10v5__ua_diff_24 = '3.80460e-13*hvp_mobility*hvp_mobility+1.20029e-12*hvp_mobility+-3.96520e-13'
+ sky130_fd_pr__pfet_g5v0d10v5__ua_diff_25 = '4.25585e-13*hvp_mobility*hvp_mobility+1.42399e-12*hvp_mobility+-3.06310e-13'
+ sky130_fd_pr__pfet_g5v0d10v5__ua_diff_26 = '4.64431e-14*hvp_mobility*hvp_mobility+-2.86875e-13*hvp_mobility+8.18810e-13'
+ sky130_fd_pr__pfet_g5v0d10v5__ua_diff_27 = '1.09521e-12*hvp_mobility*hvp_mobility+5.21640e-12*hvp_mobility+4.58110e-12'
+ sky130_fd_pr__pfet_g5v0d10v5__ua_diff_28 = '1.43774e-12*hvp_mobility*hvp_mobility+7.31546e-12*hvp_mobility+5.74930e-12'
+ sky130_fd_pr__pfet_g5v0d10v5__ua_diff_29 = '1.86734e-12*hvp_mobility*hvp_mobility+7.19696e-12*hvp_mobility+-3.32360e-15'
+ sky130_fd_pr__pfet_g5v0d10v5__ua_diff_3 = '1.59026e-12*hvp_mobility*hvp_mobility+6.11891e-12*hvp_mobility+-6.97850e-13'
+ sky130_fd_pr__pfet_g5v0d10v5__ua_diff_30 = '1.73848e-12*hvp_mobility*hvp_mobility+7.63179e-12*hvp_mobility+3.76610e-12'
+ sky130_fd_pr__pfet_g5v0d10v5__ua_diff_31 = '4.39826e-13*hvp_mobility*hvp_mobility+1.34487e-12*hvp_mobility+-1.94710e-13'
+ sky130_fd_pr__pfet_g5v0d10v5__ua_diff_32 = '9.72440e-13*hvp_mobility*hvp_mobility+3.62433e-12*hvp_mobility+-2.33480e-14'
+ sky130_fd_pr__pfet_g5v0d10v5__ua_diff_33 = '1.65074e-12*hvp_mobility*hvp_mobility+6.80998e-12*hvp_mobility+1.11620e-12'
+ sky130_fd_pr__pfet_g5v0d10v5__ua_diff_34 = '1.70476e-12*hvp_mobility*hvp_mobility+7.01491e-12*hvp_mobility+1.17220e-12'
+ sky130_fd_pr__pfet_g5v0d10v5__ua_diff_35 = '3.17154e-12*hvp_mobility*hvp_mobility+1.18834e-11*hvp_mobility+-2.61220e-12'
+ sky130_fd_pr__pfet_g5v0d10v5__ua_diff_36 = '1.45641e-13*hvp_mobility*hvp_mobility+3.27515e-13*hvp_mobility+-5.47820e-13'
+ sky130_fd_pr__pfet_g5v0d10v5__ua_diff_37 = '-3.90922e-14*hvp_mobility*hvp_mobility+-1.94016e-13*hvp_mobility+-2.77760e-13'
+ sky130_fd_pr__pfet_g5v0d10v5__ua_diff_38 = '8.31056e-14*hvp_mobility*hvp_mobility+4.45905e-13*hvp_mobility+8.47790e-13'
+ sky130_fd_pr__pfet_g5v0d10v5__ua_diff_39 = '1.59322e-13*hvp_mobility*hvp_mobility+5.65896e-13*hvp_mobility+-6.32300e-14'
+ sky130_fd_pr__pfet_g5v0d10v5__ua_diff_4 = '1.70222e-12*hvp_mobility*hvp_mobility+6.55469e-12*hvp_mobility+-1.21530e-12'
+ sky130_fd_pr__pfet_g5v0d10v5__ua_diff_40 = '1.74526e-12*hvp_mobility*hvp_mobility+6.65447e-12*hvp_mobility+-6.39800e-12'
+ sky130_fd_pr__pfet_g5v0d10v5__ua_diff_41 = '-2.66875e-14*hvp_mobility*hvp_mobility+-7.62100e-13*hvp_mobility+-2.88840e-12'
+ sky130_fd_pr__pfet_g5v0d10v5__ua_diff_42 = '3.57898e-12*hvp_mobility*hvp_mobility+1.38684e-11*hvp_mobility+7.32690e-13'
+ sky130_fd_pr__pfet_g5v0d10v5__ua_diff_43 = '1.96807e-12*hvp_mobility*hvp_mobility+7.75675e-12*hvp_mobility+-2.96510e-12'
+ sky130_fd_pr__pfet_g5v0d10v5__ua_diff_44 = '1.94521e-12*hvp_mobility*hvp_mobility+7.64160e-12*hvp_mobility+-2.82570e-12'
+ sky130_fd_pr__pfet_g5v0d10v5__ua_diff_45 = '5.10664e-12*hvp_mobility*hvp_mobility+2.03476e-11*hvp_mobility+-3.96820e-13'
+ sky130_fd_pr__pfet_g5v0d10v5__ua_diff_46 = '2.19922e-12*hvp_mobility*hvp_mobility+8.79411e-12*hvp_mobility+-3.67190e-12'
+ sky130_fd_pr__pfet_g5v0d10v5__ua_diff_47 = '2.09181e-12*hvp_mobility*hvp_mobility+8.53110e-12*hvp_mobility+-1.09830e-12'
+ sky130_fd_pr__pfet_g5v0d10v5__ua_diff_48 = '1.73623e-13*hvp_mobility*hvp_mobility+-3.26794e-13*hvp_mobility+-4.11470e-12'
+ sky130_fd_pr__pfet_g5v0d10v5__ua_diff_5 = '1.10617e-12*hvp_mobility*hvp_mobility+4.17061e-12*hvp_mobility+-8.92110e-13'
+ sky130_fd_pr__pfet_g5v0d10v5__ua_diff_6 = '1.64766e-12*hvp_mobility*hvp_mobility+6.32755e-12*hvp_mobility+-3.23770e-12'
+ sky130_fd_pr__pfet_g5v0d10v5__ua_diff_7 = '2.47501e-12*hvp_mobility*hvp_mobility+9.80362e-12*hvp_mobility+-7.36630e-13'
+ sky130_fd_pr__pfet_g5v0d10v5__ua_diff_8 = '1.64924e-12*hvp_mobility*hvp_mobility+6.50413e-12*hvp_mobility+-9.57280e-13'
+ sky130_fd_pr__pfet_g5v0d10v5__ua_diff_9 = '1.82103e-12*hvp_mobility*hvp_mobility+7.18883e-12*hvp_mobility+-4.10750e-13'
+ sky130_fd_pr__pfet_g5v0d10v5__ub_diff_0 = '-2.78950e-21*hvp_mobility*hvp_mobility+1.02867e-19*hvp_mobility+-3.54580e-19'
+ sky130_fd_pr__pfet_g5v0d10v5__ub_diff_1 = '-1.03816e-20*hvp_mobility*hvp_mobility+-9.21912e-20*hvp_mobility+-3.03520e-19'
+ sky130_fd_pr__pfet_g5v0d10v5__ub_diff_10 = '-2.15738e-21*hvp_mobility*hvp_mobility+1.75112e-20*hvp_mobility+-9.31970e-20'
+ sky130_fd_pr__pfet_g5v0d10v5__ub_diff_11 = '-4.37031e-21*hvp_mobility*hvp_mobility+6.74987e-20*hvp_mobility+-7.89000e-20'
+ sky130_fd_pr__pfet_g5v0d10v5__ub_diff_12 = '-1.85347e-20*hvp_mobility*hvp_mobility+-1.46987e-20*hvp_mobility+-6.09720e-19'
+ sky130_fd_pr__pfet_g5v0d10v5__ub_diff_13 = '-3.46000e-21*hvp_mobility*hvp_mobility+4.29825e-20*hvp_mobility+-4.70240e-19'
+ sky130_fd_pr__pfet_g5v0d10v5__ub_diff_14 = '-3.59844e-21*hvp_mobility*hvp_mobility+1.78963e-20*hvp_mobility+-2.72780e-19'
+ sky130_fd_pr__pfet_g5v0d10v5__ub_diff_15 = '-3.45328e-21*hvp_mobility*hvp_mobility+8.96794e-20*hvp_mobility+-3.75040e-19'
+ sky130_fd_pr__pfet_g5v0d10v5__ub_diff_16 = '-5.74000e-21*hvp_mobility*hvp_mobility+-1.84250e-20*hvp_mobility+-6.45970e-19'
+ sky130_fd_pr__pfet_g5v0d10v5__ub_diff_17 = '-7.56744e-21*hvp_mobility*hvp_mobility+-3.93150e-20*hvp_mobility+-2.04810e-20'
+ sky130_fd_pr__pfet_g5v0d10v5__ub_diff_18 = '-4.40156e-21*hvp_mobility*hvp_mobility+-5.21037e-20*hvp_mobility+-6.99740e-19'
+ sky130_fd_pr__pfet_g5v0d10v5__ub_diff_19 = '-1.05372e-20*hvp_mobility*hvp_mobility+-4.88813e-20*hvp_mobility+-3.42630e-19'
+ sky130_fd_pr__pfet_g5v0d10v5__ub_diff_2 = '-4.05344e-21*hvp_mobility*hvp_mobility+5.22562e-20*hvp_mobility+-3.67290e-19'
+ sky130_fd_pr__pfet_g5v0d10v5__ub_diff_20 = '-7.36747e-21*hvp_mobility*hvp_mobility+4.54426e-20*hvp_mobility+-1.57650e-19'
+ sky130_fd_pr__pfet_g5v0d10v5__ub_diff_21 = '-6.03000e-21*hvp_mobility*hvp_mobility+-9.49000e-21*hvp_mobility+-8.34280e-19'
+ sky130_fd_pr__pfet_g5v0d10v5__ub_diff_22 = '-6.39706e-21*hvp_mobility*hvp_mobility+-9.56513e-20*hvp_mobility+-3.74720e-20'
+ sky130_fd_pr__pfet_g5v0d10v5__ub_diff_23 = '-3.46000e-21*hvp_mobility*hvp_mobility+-2.57825e-20*hvp_mobility+-2.83850e-19'
+ sky130_fd_pr__pfet_g5v0d10v5__ub_diff_24 = '-2.99469e-21*hvp_mobility*hvp_mobility+-3.56188e-20*hvp_mobility+-7.27610e-19'
+ sky130_fd_pr__pfet_g5v0d10v5__ub_diff_25 = '-3.63469e-21*hvp_mobility*hvp_mobility+-4.45612e-20*hvp_mobility+-6.24500e-19'
+ sky130_fd_pr__pfet_g5v0d10v5__ub_diff_26 = '-1.31281e-21*hvp_mobility*hvp_mobility+2.59988e-20*hvp_mobility+-2.60250e-19'
+ sky130_fd_pr__pfet_g5v0d10v5__ub_diff_27 = '-6.14375e-21*hvp_mobility*hvp_mobility+1.96500e-20*hvp_mobility+-1.22540e-18'
+ sky130_fd_pr__pfet_g5v0d10v5__ub_diff_28 = '-3.76625e-21*hvp_mobility*hvp_mobility+1.88750e-21*hvp_mobility+-9.59190e-19'
+ sky130_fd_pr__pfet_g5v0d10v5__ub_diff_29 = '-4.63375e-21*hvp_mobility*hvp_mobility+-8.46500e-21*hvp_mobility+-4.07000e-19'
+ sky130_fd_pr__pfet_g5v0d10v5__ub_diff_3 = '-4.89344e-21*hvp_mobility*hvp_mobility+-2.27125e-21*hvp_mobility+-2.66150e-19'
+ sky130_fd_pr__pfet_g5v0d10v5__ub_diff_30 = '-5.83969e-21*hvp_mobility*hvp_mobility+-3.57763e-20*hvp_mobility+-2.77390e-19'
+ sky130_fd_pr__pfet_g5v0d10v5__ub_diff_31 = '-3.65906e-21*hvp_mobility*hvp_mobility+-4.67637e-20*hvp_mobility+-6.69520e-19'
+ sky130_fd_pr__pfet_g5v0d10v5__ub_diff_32 = '-4.53594e-21*hvp_mobility*hvp_mobility+-4.90613e-20*hvp_mobility+-5.69030e-19'
+ sky130_fd_pr__pfet_g5v0d10v5__ub_diff_33 = '-4.42938e-21*hvp_mobility*hvp_mobility+5.32875e-20*hvp_mobility+-5.36590e-19'
+ sky130_fd_pr__pfet_g5v0d10v5__ub_diff_34 = '-4.58750e-21*hvp_mobility*hvp_mobility+6.75000e-21*hvp_mobility+-9.18000e-19'
+ sky130_fd_pr__pfet_g5v0d10v5__ub_diff_35 = '-1.42341e-20*hvp_mobility*hvp_mobility+-2.01131e-19*hvp_mobility+-3.25830e-19'
+ sky130_fd_pr__pfet_g5v0d10v5__ub_diff_36 = '-5.94803e-21*hvp_mobility*hvp_mobility+-2.32516e-20*hvp_mobility+8.96610e-20'
+ sky130_fd_pr__pfet_g5v0d10v5__ub_diff_37 = '-5.16625e-21*hvp_mobility*hvp_mobility+-4.68500e-20*hvp_mobility+1.43530e-19'
+ sky130_fd_pr__pfet_g5v0d10v5__ub_diff_38 = '-4.78281e-21*hvp_mobility*hvp_mobility+-5.28750e-22*hvp_mobility+2.95830e-19'
+ sky130_fd_pr__pfet_g5v0d10v5__ub_diff_39 = '-3.91106e-21*hvp_mobility*hvp_mobility+3.35250e-21*hvp_mobility+1.28700e-20'
+ sky130_fd_pr__pfet_g5v0d10v5__ub_diff_4 = '-4.77750e-21*hvp_mobility*hvp_mobility+-1.54075e-20*hvp_mobility+-2.88840e-19'
+ sky130_fd_pr__pfet_g5v0d10v5__ub_diff_40 = '-1.37469e-20*hvp_mobility*hvp_mobility+-7.62500e-22*hvp_mobility+-1.61270e-18'
+ sky130_fd_pr__pfet_g5v0d10v5__ub_diff_41 = '-1.22027e-20*hvp_mobility*hvp_mobility+-7.07868e-20*hvp_mobility+-1.71850e-19'
+ sky130_fd_pr__pfet_g5v0d10v5__ub_diff_42 = '-1.82180e-20*hvp_mobility*hvp_mobility+-5.65000e-20*hvp_mobility+-5.07720e-20'
+ sky130_fd_pr__pfet_g5v0d10v5__ub_diff_43 = '-7.39531e-21*hvp_mobility*hvp_mobility+-1.48062e-20*hvp_mobility+-8.08530e-19'
+ sky130_fd_pr__pfet_g5v0d10v5__ub_diff_44 = '-5.46125e-21*hvp_mobility*hvp_mobility+-9.62500e-21*hvp_mobility+-9.02120e-19'
+ sky130_fd_pr__pfet_g5v0d10v5__ub_diff_45 = '-8.34000e-21*hvp_mobility*hvp_mobility+-1.11150e-20*hvp_mobility+-2.45170e-19'
+ sky130_fd_pr__pfet_g5v0d10v5__ub_diff_46 = '-4.37500e-21*hvp_mobility*hvp_mobility+8.60950e-20*hvp_mobility+-9.11020e-19'
+ sky130_fd_pr__pfet_g5v0d10v5__ub_diff_47 = '-5.41344e-21*hvp_mobility*hvp_mobility+2.49613e-20*hvp_mobility+-8.30740e-19'
+ sky130_fd_pr__pfet_g5v0d10v5__ub_diff_48 = '-4.63437e-21*hvp_mobility*hvp_mobility+-6.01875e-21*hvp_mobility+-7.92450e-20'
+ sky130_fd_pr__pfet_g5v0d10v5__ub_diff_5 = '-4.05250e-21*hvp_mobility*hvp_mobility+-1.65975e-20*hvp_mobility+-5.06050e-19'
+ sky130_fd_pr__pfet_g5v0d10v5__ub_diff_6 = '-3.60438e-21*hvp_mobility*hvp_mobility+4.77500e-20*hvp_mobility+-9.20030e-19'
+ sky130_fd_pr__pfet_g5v0d10v5__ub_diff_7 = '-4.74875e-21*hvp_mobility*hvp_mobility+2.19100e-20*hvp_mobility+-2.59750e-19'
+ sky130_fd_pr__pfet_g5v0d10v5__ub_diff_8 = '-4.11594e-21*hvp_mobility*hvp_mobility+1.24412e-20*hvp_mobility+-3.92510e-19'
+ sky130_fd_pr__pfet_g5v0d10v5__ub_diff_9 = '-4.09906e-21*hvp_mobility*hvp_mobility+9.64875e-21*hvp_mobility+-1.55970e-19'
+ sky130_fd_pr__pfet_g5v0d10v5__voff_diff_22 = '7.57187e-05*hvp_subvt*hvp_subvt+3.82337e-03*hvp_subvt+-1.65050e-02'
+ sky130_fd_pr__pfet_g5v0d10v5__voff_diff_35 = '1.34170e-03*hvp_subvt*hvp_subvt+1.13463e-02*hvp_subvt+-8.80620e-03'
+ sky130_fd_pr__pfet_g5v0d10v5__voff_diff_37 = '-2.26531e-04*hvp_subvt*hvp_subvt+5.09875e-04*hvp_subvt+-3.88520e-02'
+ sky130_fd_pr__pfet_g5v0d10v5__voff_diff_38 = '1.23781e-04*hvp_subvt*hvp_subvt+1.58062e-03*hvp_subvt+-3.65400e-02'
+ sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_0 = '-3.31937e+01*hvp_saturation*hvp_saturation+6.19750e+01*hvp_saturation+-3.18610e+03'
+ sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_11 = '2.98375e+02*hvp_saturation*hvp_saturation+5.76075e+03*hvp_saturation+-2.66900e+03'
+ sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_12 = '3.51125e+01*hvp_saturation*hvp_saturation+1.80067e+03*hvp_saturation+-2.87640e+03'
+ sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_13 = '-1.16500e+01*hvp_saturation*hvp_saturation+7.84600e+02*hvp_saturation+-1.10210e+03'
+ sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_15 = '-3.99562e+01*hvp_saturation*hvp_saturation+-1.97025e+02*hvp_saturation+-4.03310e+03'
+ sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_2 = '-4.29469e+01*hvp_saturation*hvp_saturation+-2.92312e+02*hvp_saturation+-3.56980e+03'
+ sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_20 = '1.92456e+02*hvp_saturation*hvp_saturation+4.94512e+03*hvp_saturation+-7.26080e+03'
+ sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_21 = '-2.68250e+01*hvp_saturation*hvp_saturation+6.78150e+02*hvp_saturation+-4.65850e+03'
+ sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_26 = '-3.71813e+01*hvp_saturation*hvp_saturation+-3.74250e+01*hvp_saturation+-4.33720e+03'
+ sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_27 = '-2.60875e+01*hvp_saturation*hvp_saturation+-4.81500e+01*hvp_saturation+-2.67600e+03'
+ sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_28 = '-2.51844e+01*hvp_saturation*hvp_saturation+8.70375e+01*hvp_saturation+-2.38100e+03'
+ sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_33 = '-3.82156e+01*hvp_saturation*hvp_saturation+-8.80625e+01*hvp_saturation+-4.05180e+03'
+ sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_34 = '-2.93219e+01*hvp_saturation*hvp_saturation+2.46375e+01*hvp_saturation+-2.16630e+03'
+ sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_40 = '6.16375e+01*hvp_saturation*hvp_saturation+2.71443e+03*hvp_saturation+-8.18450e+03'
+ sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_41 = '1.61500e+01*hvp_saturation*hvp_saturation+2.28962e+03*hvp_saturation+-2.86290e+03'
+ sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_42 = '5.47806e+01*hvp_saturation*hvp_saturation+2.23829e+03*hvp_saturation+-7.58340e+02'
+ sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_46 = '1.32625e+01*hvp_saturation*hvp_saturation+1.86915e+03*hvp_saturation+-3.56460e+03'
+ sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_47 = '9.99125e+01*hvp_saturation*hvp_saturation+2.42845e+03*hvp_saturation+-3.10380e+03'
+ sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_48 = '5.60312e+00*hvp_saturation*hvp_saturation+1.34291e+03*hvp_saturation+-3.50820e+03'
+ sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_6 = '-9.06562e+00*hvp_saturation*hvp_saturation+1.44669e+03*hvp_saturation+-4.01460e+03'
+ sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_0 = '-3.69375e-05*hvp_threshold*hvp_threshold+-1.47107e-02*hvp_threshold+-2.83710e-02'
+ sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_1 = '-1.81250e-05*hvp_threshold*hvp_threshold+-1.16695e-02*hvp_threshold+-2.18830e-02'
+ sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_10 = '3.28125e-06*hvp_threshold*hvp_threshold+-1.22281e-02*hvp_threshold+-1.15090e-02'
+ sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_11 = '-7.59375e-06*hvp_threshold*hvp_threshold+-2.11184e-02*hvp_threshold+-5.29850e-02'
+ sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_12 = '-1.82437e-05*hvp_threshold*hvp_threshold+-1.77556e-02*hvp_threshold+-5.68060e-03'
+ sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_13 = '1.50312e-05*hvp_threshold*hvp_threshold+-1.96836e-02*hvp_threshold+-3.67360e-02'
+ sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_14 = '2.68438e-05*hvp_threshold*hvp_threshold+-1.24334e-02*hvp_threshold+-2.57480e-02'
+ sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_15 = '-2.00938e-05*hvp_threshold*hvp_threshold+-1.44011e-02*hvp_threshold+-3.08980e-02'
+ sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_16 = '2.33750e-05*hvp_threshold*hvp_threshold+-1.34247e-02*hvp_threshold+-1.32800e-02'
+ sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_17 = '-1.29375e-04*hvp_threshold*hvp_threshold+-1.22735e-02*hvp_threshold+-2.41500e-02'
+ sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_18 = '1.56375e-05*hvp_threshold*hvp_threshold+-1.17236e-02*hvp_threshold+-5.30670e-03'
+ sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_19 = '-1.85381e-04*hvp_threshold*hvp_threshold+-1.17102e-02*hvp_threshold+-8.44390e-03'
+ sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_2 = '-6.27188e-05*hvp_threshold*hvp_threshold+-1.75204e-02*hvp_threshold+-2.73320e-02'
+ sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_20 = '4.30312e-05*hvp_threshold*hvp_threshold+-1.72169e-02*hvp_threshold+-4.49610e-02'
+ sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_21 = '-7.12500e-06*hvp_threshold*hvp_threshold+-1.78290e-02*hvp_threshold+-1.39050e-02'
+ sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_22 = '-7.62278e-04*hvp_threshold*hvp_threshold+-1.34176e-02*hvp_threshold+-3.90110e-02'
+ sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_23 = '1.94687e-05*hvp_threshold*hvp_threshold+-1.22009e-02*hvp_threshold+-3.08610e-02'
+ sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_24 = '2.93437e-05*hvp_threshold*hvp_threshold+-1.17679e-02*hvp_threshold+-1.02160e-02'
+ sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_25 = '1.93438e-05*hvp_threshold*hvp_threshold+-1.13241e-02*hvp_threshold+-1.13580e-02'
+ sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_26 = '-5.50938e-05*hvp_threshold*hvp_threshold+-1.41464e-02*hvp_threshold+-3.53710e-02'
+ sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_27 = '9.09375e-06*hvp_threshold*hvp_threshold+-1.45484e-02*hvp_threshold+-3.03830e-02'
+ sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_28 = '1.22188e-05*hvp_threshold*hvp_threshold+-1.41714e-02*hvp_threshold+-3.20780e-02'
+ sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_29 = '2.30938e-05*hvp_threshold*hvp_threshold+-1.34341e-02*hvp_threshold+-1.82110e-02'
+ sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_3 = '3.22000e-05*hvp_threshold*hvp_threshold+-1.45950e-02*hvp_threshold+-9.89020e-03'
+ sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_30 = '-4.75000e-06*hvp_threshold*hvp_threshold+-1.17795e-02*hvp_threshold+-3.10000e-02'
+ sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_31 = '1.30938e-05*hvp_threshold*hvp_threshold+-1.18634e-02*hvp_threshold+-1.09980e-02'
+ sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_32 = '1.14687e-05*hvp_threshold*hvp_threshold+-1.15724e-02*hvp_threshold+-1.10280e-02'
+ sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_33 = '-5.51562e-05*hvp_threshold*hvp_threshold+-1.46231e-02*hvp_threshold+-3.57980e-02'
+ sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_34 = '1.09375e-05*hvp_threshold*hvp_threshold+-1.40602e-02*hvp_threshold+-2.40290e-02'
+ sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_35 = '1.72250e-03*hvp_threshold*hvp_threshold+-9.76100e-03*hvp_threshold+-3.83990e-02'
+ sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_36 = '-7.08750e-05*hvp_threshold*hvp_threshold+-1.07607e-02*hvp_threshold+-2.02940e-02'
+ sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_37 = '-1.64594e-04*hvp_threshold*hvp_threshold+-1.47446e-02*hvp_threshold+-1.94380e-02'
+ sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_38 = '-5.93125e-05*hvp_threshold*hvp_threshold+-1.29327e-02*hvp_threshold+-1.96540e-02'
+ sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_39 = '-8.39250e-05*hvp_threshold*hvp_threshold+-1.25435e-02*hvp_threshold+-6.04220e-03'
+ sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_4 = '2.78750e-05*hvp_threshold*hvp_threshold+-1.33815e-02*hvp_threshold+-2.03600e-02'
+ sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_40 = '4.18125e-05*hvp_threshold*hvp_threshold+-2.88485e-02*hvp_threshold+2.65970e-02'
+ sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_41 = '-3.14688e-05*hvp_threshold*hvp_threshold+-2.55204e-02*hvp_threshold+-4.03650e-02'
+ sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_42 = '4.50625e-05*hvp_threshold*hvp_threshold+-2.66540e-02*hvp_threshold+-1.68850e-02'
+ sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_43 = '2.40313e-05*hvp_threshold*hvp_threshold+-1.82301e-02*hvp_threshold+-2.19180e-02'
+ sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_44 = '2.50000e-05*hvp_threshold*hvp_threshold+-1.42752e-02*hvp_threshold+-1.60430e-02'
+ sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_45 = '8.50000e-06*hvp_threshold*hvp_threshold+-1.39445e-02*hvp_threshold+-1.40800e-02'
+ sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_46 = '-9.71875e-06*hvp_threshold*hvp_threshold+-2.51645e-02*hvp_threshold+-7.89650e-03'
+ sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_47 = '2.03125e-05*hvp_threshold*hvp_threshold+-1.77300e-02*hvp_threshold+-2.01350e-02'
+ sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_48 = '-4.14687e-05*hvp_threshold*hvp_threshold+-2.43451e-02*hvp_threshold+-6.32560e-02'
+ sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_5 = '1.40625e-05*hvp_threshold*hvp_threshold+-1.18798e-02*hvp_threshold+-1.26520e-02'
+ sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_6 = '-5.08000e-05*hvp_threshold*hvp_threshold+-1.80235e-02*hvp_threshold+-1.89820e-03'
+ sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_7 = '3.11250e-05*hvp_threshold*hvp_threshold+-1.52023e-02*hvp_threshold+-1.17440e-02'
+ sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_8 = '1.94812e-05*hvp_threshold*hvp_threshold+-1.40639e-02*hvp_threshold+-8.11420e-03'
+ sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_9 = '1.24375e-05*hvp_threshold*hvp_threshold+-1.29505e-02*hvp_threshold+-2.01470e-02'
+ sky130_fd_pr__pfet_g5v0d10v5__wint_diff = '8.04375e-09*diff_cd'
+ sky130_fd_pr__esd_pfet_g5v0d10v5__ajunction_mult = '-2.50000e-06*hvp_diode*hvp_diode+1.81850e-02*hvp_diode+1.00500e+00'
+ sky130_fd_pr__esd_pfet_g5v0d10v5__dlc_diff = '-4.33125e-09*poly_cd'
+ sky130_fd_pr__esd_pfet_g5v0d10v5__dwc_diff = '8.04375e-09*diff_cd'
+ sky130_fd_pr__esd_pfet_g5v0d10v5__k2_diff_0 = '-2.10781e-05*hvp_bodyeffect*hvp_bodyeffect+1.52921e-03*hvp_bodyeffect+2.59040e-03'
+ sky130_fd_pr__esd_pfet_g5v0d10v5__k2_diff_1 = '2.11122e-04*hvp_bodyeffect*hvp_bodyeffect+2.48336e-03*hvp_bodyeffect+2.52960e-03'
+ sky130_fd_pr__esd_pfet_g5v0d10v5__k2_diff_2 = '1.54622e-04*hvp_bodyeffect*hvp_bodyeffect+1.79881e-03*hvp_bodyeffect+1.17380e-03'
+ sky130_fd_pr__esd_pfet_g5v0d10v5__k2_diff_3 = '4.56875e-06*hvp_bodyeffect*hvp_bodyeffect+1.63363e-03*hvp_bodyeffect+2.50330e-03'
+ sky130_fd_pr__esd_pfet_g5v0d10v5__k2_diff_4 = '-3.78437e-06*hvp_bodyeffect*hvp_bodyeffect+1.55779e-03*hvp_bodyeffect+2.72320e-03'
+ sky130_fd_pr__esd_pfet_g5v0d10v5__k2_diff_5 = '2.21903e-04*hvp_bodyeffect*hvp_bodyeffect+2.59791e-03*hvp_bodyeffect+2.60990e-03'
+ sky130_fd_pr__esd_pfet_g5v0d10v5__k2_diff_6 = '2.05675e-04*hvp_bodyeffect*hvp_bodyeffect+2.49152e-03*hvp_bodyeffect+2.81810e-03'
+ sky130_fd_pr__esd_pfet_g5v0d10v5__k2_diff_7 = '2.38472e-04*hvp_bodyeffect*hvp_bodyeffect+2.56914e-03*hvp_bodyeffect+2.43090e-03'
+ sky130_fd_pr__esd_pfet_g5v0d10v5__lint_diff = '-4.33125e-09*poly_cd'
+ sky130_fd_pr__esd_pfet_g5v0d10v5__nfactor_diff_0 = '-1.27274e-02*hvp_subvt*hvp_subvt+-3.96912e-02*hvp_subvt+-6.31470e-02'
+ sky130_fd_pr__esd_pfet_g5v0d10v5__nfactor_diff_1 = '1.98816e-02*hvp_subvt*hvp_subvt+6.77894e-02*hvp_subvt+-7.47430e-02'
+ sky130_fd_pr__esd_pfet_g5v0d10v5__nfactor_diff_2 = '2.11058e-02*hvp_subvt*hvp_subvt+5.53791e-02*hvp_subvt+-1.83720e-01'
+ sky130_fd_pr__esd_pfet_g5v0d10v5__nfactor_diff_3 = '6.86153e-03*hvp_subvt*hvp_subvt+2.68401e-02*hvp_subvt+-8.88150e-02'
+ sky130_fd_pr__esd_pfet_g5v0d10v5__nfactor_diff_4 = '-3.06744e-03*hvp_subvt*hvp_subvt+-1.25690e-02*hvp_subvt+-6.78450e-02'
+ sky130_fd_pr__esd_pfet_g5v0d10v5__nfactor_diff_5 = '1.84450e-02*hvp_subvt*hvp_subvt+8.36988e-02*hvp_subvt+-6.07250e-02'
+ sky130_fd_pr__esd_pfet_g5v0d10v5__nfactor_diff_6 = '1.63519e-02*hvp_subvt*hvp_subvt+6.95986e-02*hvp_subvt+-6.75050e-02'
+ sky130_fd_pr__esd_pfet_g5v0d10v5__nfactor_diff_7 = '1.76127e-02*hvp_subvt*hvp_subvt+8.56312e-02*hvp_subvt+-5.34990e-02'
+ sky130_fd_pr__esd_pfet_g5v0d10v5__overlap_mult = '8.68750e-04*hvtox*hvtox+7.40000e-02*hvtox+9.82100e-01'
+ sky130_fd_pr__esd_pfet_g5v0d10v5__pjunction_mult = '-1.25000e-06*hvp_diode*hvp_diode+1.61550e-02*hvp_diode+1.00900e+00'
+ sky130_fd_pr__esd_pfet_g5v0d10v5__toxe_mult = '1.50000e-02*hvtox+1.00000e+00'
+ sky130_fd_pr__esd_pfet_g5v0d10v5__u0_diff_0 = '5.65938e-06*hvp_mobility*hvp_mobility+3.15263e-04*hvp_mobility+1.32160e-03'
+ sky130_fd_pr__esd_pfet_g5v0d10v5__u0_diff_1 = '-2.87138e-04*hvp_mobility*hvp_mobility+-8.66623e-04*hvp_mobility+1.39910e-03'
+ sky130_fd_pr__esd_pfet_g5v0d10v5__u0_diff_2 = '-5.23449e-05*hvp_mobility*hvp_mobility+3.43595e-05*hvp_mobility+9.45920e-04'
+ sky130_fd_pr__esd_pfet_g5v0d10v5__u0_diff_3 = '-2.04478e-05*hvp_mobility*hvp_mobility+2.05116e-04*hvp_mobility+1.52690e-03'
+ sky130_fd_pr__esd_pfet_g5v0d10v5__u0_diff_4 = '-5.65434e-06*hvp_mobility*hvp_mobility+2.72167e-04*hvp_mobility+1.08030e-03'
+ sky130_fd_pr__esd_pfet_g5v0d10v5__u0_diff_5 = '-3.07647e-04*hvp_mobility*hvp_mobility+-9.55186e-04*hvp_mobility+1.36540e-03'
+ sky130_fd_pr__esd_pfet_g5v0d10v5__u0_diff_6 = '-3.20093e-04*hvp_mobility*hvp_mobility+-9.21868e-04*hvp_mobility+1.18510e-03'
+ sky130_fd_pr__esd_pfet_g5v0d10v5__u0_diff_7 = '-2.78399e-04*hvp_mobility*hvp_mobility+-8.08280e-04*hvp_mobility+1.39250e-03'
+ sky130_fd_pr__esd_pfet_g5v0d10v5__ua_diff_0 = '5.20158e-12*hvp_mobility*hvp_mobility+2.34789e-11*hvp_mobility+1.32290e-11'
+ sky130_fd_pr__esd_pfet_g5v0d10v5__ua_diff_1 = '-2.59361e-12*hvp_mobility*hvp_mobility+-6.92929e-12*hvp_mobility+1.40790e-11'
+ sky130_fd_pr__esd_pfet_g5v0d10v5__ua_diff_2 = '2.41118e-12*hvp_mobility*hvp_mobility+3.73976e-12*hvp_mobility+-1.68180e-11'
+ sky130_fd_pr__esd_pfet_g5v0d10v5__ua_diff_3 = '1.59362e-12*hvp_mobility*hvp_mobility+8.06351e-12*hvp_mobility+1.43170e-11'
+ sky130_fd_pr__esd_pfet_g5v0d10v5__ua_diff_4 = '1.04375e-12*hvp_mobility*hvp_mobility+7.83376e-12*hvp_mobility+1.10800e-11'
+ sky130_fd_pr__esd_pfet_g5v0d10v5__ua_diff_5 = '-2.40611e-12*hvp_mobility*hvp_mobility+-6.97082e-12*hvp_mobility+1.37110e-11'
+ sky130_fd_pr__esd_pfet_g5v0d10v5__ua_diff_6 = '-2.20597e-12*hvp_mobility*hvp_mobility+-5.40387e-12*hvp_mobility+1.63660e-11'
+ sky130_fd_pr__esd_pfet_g5v0d10v5__ua_diff_7 = '-8.73837e-13*hvp_mobility*hvp_mobility+3.15810e-12*hvp_mobility+1.81600e-11'
+ sky130_fd_pr__esd_pfet_g5v0d10v5__ub_diff_0 = '1.44281e-21*hvp_mobility*hvp_mobility+1.79234e-19*hvp_mobility+3.17180e-19'
+ sky130_fd_pr__esd_pfet_g5v0d10v5__ub_diff_1 = '-1.25421e-19*hvp_mobility*hvp_mobility+-3.36819e-19*hvp_mobility+3.16310e-19'
+ sky130_fd_pr__esd_pfet_g5v0d10v5__ub_diff_2 = '-2.15400e-20*hvp_mobility*hvp_mobility+6.46875e-20*hvp_mobility+2.83220e-19'
+ sky130_fd_pr__esd_pfet_g5v0d10v5__ub_diff_3 = '-4.89781e-21*hvp_mobility*hvp_mobility+1.36454e-19*hvp_mobility+2.96490e-19'
+ sky130_fd_pr__esd_pfet_g5v0d10v5__ub_diff_4 = '7.80313e-22*hvp_mobility*hvp_mobility+1.71104e-19*hvp_mobility+2.86280e-19'
+ sky130_fd_pr__esd_pfet_g5v0d10v5__ub_diff_5 = '-1.35431e-19*hvp_mobility*hvp_mobility+-3.89545e-19*hvp_mobility+3.62470e-19'
+ sky130_fd_pr__esd_pfet_g5v0d10v5__ub_diff_6 = '-1.55654e-19*hvp_mobility*hvp_mobility+-4.54207e-19*hvp_mobility+3.71300e-19'
+ sky130_fd_pr__esd_pfet_g5v0d10v5__ub_diff_7 = '-1.24436e-19*hvp_mobility*hvp_mobility+-3.02338e-19*hvp_mobility+4.24420e-19'
+ sky130_fd_pr__esd_pfet_g5v0d10v5__voff_diff_0 = '-6.25416e-04*hvp_subvt*hvp_subvt+-2.64591e-03*hvp_subvt+1.94320e-02'
+ sky130_fd_pr__esd_pfet_g5v0d10v5__voff_diff_1 = '3.93169e-03*hvp_subvt*hvp_subvt+1.78005e-02*hvp_subvt+1.89810e-02'
+ sky130_fd_pr__esd_pfet_g5v0d10v5__voff_diff_2 = '1.15994e-03*hvp_subvt*hvp_subvt+4.76000e-03*hvp_subvt+1.64930e-02'
+ sky130_fd_pr__esd_pfet_g5v0d10v5__voff_diff_3 = '3.41375e-04*hvp_subvt*hvp_subvt+1.85075e-03*hvp_subvt+2.01980e-02'
+ sky130_fd_pr__esd_pfet_g5v0d10v5__voff_diff_4 = '-1.33625e-04*hvp_subvt*hvp_subvt+8.00000e-04*hvp_subvt+2.17230e-02'
+ sky130_fd_pr__esd_pfet_g5v0d10v5__voff_diff_5 = '4.28875e-03*hvp_subvt*hvp_subvt+1.78815e-02*hvp_subvt+2.23340e-02'
+ sky130_fd_pr__esd_pfet_g5v0d10v5__voff_diff_6 = '4.94750e-03*hvp_subvt*hvp_subvt+2.10115e-02*hvp_subvt+2.29640e-02'
+ sky130_fd_pr__esd_pfet_g5v0d10v5__voff_diff_7 = '3.76809e-03*hvp_subvt*hvp_subvt+1.54001e-02*hvp_subvt+2.25300e-02'
+ sky130_fd_pr__esd_pfet_g5v0d10v5__vsat_diff_0 = '2.10246e+03*hvp_saturation*hvp_saturation+1.67444e+04*hvp_saturation+-5.98380e+03'
+ sky130_fd_pr__esd_pfet_g5v0d10v5__vsat_diff_1 = '1.17156e+02*hvp_saturation*hvp_saturation+7.30638e+03*hvp_saturation+-9.02000e+03'
+ sky130_fd_pr__esd_pfet_g5v0d10v5__vsat_diff_2 = '9.62440e+02*hvp_saturation*hvp_saturation+1.25120e+04*hvp_saturation+-8.40040e+02'
+ sky130_fd_pr__esd_pfet_g5v0d10v5__vsat_diff_3 = '9.42719e+02*hvp_saturation*hvp_saturation+1.05574e+04*hvp_saturation+-1.41430e+04'
+ sky130_fd_pr__esd_pfet_g5v0d10v5__vsat_diff_4 = '6.18219e+02*hvp_saturation*hvp_saturation+1.00669e+04*hvp_saturation+-2.26100e+03'
+ sky130_fd_pr__esd_pfet_g5v0d10v5__vsat_diff_5 = '6.99437e+01*hvp_saturation*hvp_saturation+7.46788e+03*hvp_saturation+-2.37860e+03'
+ sky130_fd_pr__esd_pfet_g5v0d10v5__vsat_diff_6 = '2.48053e+02*hvp_saturation*hvp_saturation+9.17688e+03*hvp_saturation+-2.32340e+02'
+ sky130_fd_pr__esd_pfet_g5v0d10v5__vsat_diff_7 = '-1.70669e+02*hvp_saturation*hvp_saturation+6.31912e+03*hvp_saturation+-1.15780e+03'
+ sky130_fd_pr__esd_pfet_g5v0d10v5__vth0_diff_0 = '-5.75750e-05*hvp_threshold*hvp_threshold+-1.47074e-02*hvp_threshold+1.19570e-03'
+ sky130_fd_pr__esd_pfet_g5v0d10v5__vth0_diff_1 = '3.84315e-03*hvp_threshold*hvp_threshold+5.33625e-04*hvp_threshold+7.28410e-03'
+ sky130_fd_pr__esd_pfet_g5v0d10v5__vth0_diff_2 = '4.81844e-04*hvp_threshold*hvp_threshold+-1.22659e-02*hvp_threshold+1.16330e-02'
+ sky130_fd_pr__esd_pfet_g5v0d10v5__vth0_diff_3 = '1.15800e-04*hvp_threshold*hvp_threshold+-1.44595e-02*hvp_threshold+3.01220e-03'
+ sky130_fd_pr__esd_pfet_g5v0d10v5__vth0_diff_4 = '-1.67846e-04*hvp_threshold*hvp_threshold+-1.56219e-02*hvp_threshold+-6.96650e-06'
+ sky130_fd_pr__esd_pfet_g5v0d10v5__vth0_diff_5 = '4.32071e-03*hvp_threshold*hvp_threshold+2.16613e-03*hvp_threshold+1.14220e-03'
+ sky130_fd_pr__esd_pfet_g5v0d10v5__vth0_diff_6 = '5.19909e-03*hvp_threshold*hvp_threshold+5.96600e-03*hvp_threshold+3.74060e-03'
+ sky130_fd_pr__esd_pfet_g5v0d10v5__vth0_diff_7 = '3.70357e-03*hvp_threshold*hvp_threshold+-4.89250e-04*hvp_threshold+2.31290e-03'
+ sky130_fd_pr__esd_pfet_g5v0d10v5__wint_diff = '8.04375e-09*diff_cd'
+ sky130_fd_pr__pfet_01v8_lvt__a0_diff_0 = '-1.31375e-03*lvlp_saturation*lvlp_saturation+-3.00382e-02*lvlp_saturation+6.05170e-02'
+ sky130_fd_pr__pfet_01v8_lvt__a0_diff_1 = '-1.06844e-04*lvlp_saturation*lvlp_saturation+-1.22319e-02*lvlp_saturation+8.91620e-02'
+ sky130_fd_pr__pfet_01v8_lvt__a0_diff_10 = '-1.04312e-04*lvlp_saturation*lvlp_saturation+-2.07575e-03*lvlp_saturation+9.41760e-02'
+ sky130_fd_pr__pfet_01v8_lvt__a0_diff_12 = '-1.41875e-05*lvlp_saturation*lvlp_saturation+-4.49000e-03*lvlp_saturation+7.73390e-02'
+ sky130_fd_pr__pfet_01v8_lvt__a0_diff_13 = '9.52313e-03*lvlp_saturation*lvlp_saturation+3.61900e-02*lvlp_saturation+1.02870e-01'
+ sky130_fd_pr__pfet_01v8_lvt__a0_diff_14 = '-6.02719e-04*lvlp_saturation*lvlp_saturation+-1.19209e-02*lvlp_saturation+1.08600e-01'
+ sky130_fd_pr__pfet_01v8_lvt__a0_diff_15 = '-5.64656e-04*lvlp_saturation*lvlp_saturation+-6.79113e-03*lvlp_saturation+1.04690e-01'
+ sky130_fd_pr__pfet_01v8_lvt__a0_diff_16 = '-7.53125e-05*lvlp_saturation*lvlp_saturation+-8.62500e-05*lvlp_saturation+1.06920e-01'
+ sky130_fd_pr__pfet_01v8_lvt__a0_diff_17 = '-5.00000e-05*lvlp_saturation*lvlp_saturation+-4.60000e-04*lvlp_saturation+1.02670e-01'
+ sky130_fd_pr__pfet_01v8_lvt__a0_diff_19 = '-3.49609e-05*lvlp_saturation*lvlp_saturation+-1.41871e-02*lvlp_saturation+5.81010e-02'
+ sky130_fd_pr__pfet_01v8_lvt__a0_diff_2 = '-6.72531e-04*lvlp_saturation*lvlp_saturation+-1.32376e-02*lvlp_saturation+1.14640e-01'
+ sky130_fd_pr__pfet_01v8_lvt__a0_diff_20 = '-1.29100e-03*lvlp_saturation*lvlp_saturation+-2.92113e-02*lvlp_saturation+4.75510e-02'
+ sky130_fd_pr__pfet_01v8_lvt__a0_diff_21 = '-1.30634e-03*lvlp_saturation*lvlp_saturation+-1.82431e-02*lvlp_saturation+7.30490e-02'
+ sky130_fd_pr__pfet_01v8_lvt__a0_diff_22 = '-7.04357e-04*lvlp_saturation*lvlp_saturation+-1.23797e-02*lvlp_saturation+6.08440e-02'
+ sky130_fd_pr__pfet_01v8_lvt__a0_diff_23 = '-7.75000e-05*lvlp_saturation*lvlp_saturation+-8.05000e-04*lvlp_saturation+1.16730e-01'
+ sky130_fd_pr__pfet_01v8_lvt__a0_diff_24 = '-1.36875e-04*lvlp_saturation*lvlp_saturation+-1.86750e-03*lvlp_saturation+1.13390e-01'
+ sky130_fd_pr__pfet_01v8_lvt__a0_diff_26 = '-7.97719e-04*lvlp_saturation*lvlp_saturation+-1.02771e-02*lvlp_saturation+6.77150e-02'
+ sky130_fd_pr__pfet_01v8_lvt__a0_diff_3 = '-9.41094e-04*lvlp_saturation*lvlp_saturation+-1.58579e-02*lvlp_saturation+9.31460e-02'
+ sky130_fd_pr__pfet_01v8_lvt__a0_diff_6 = '-4.18781e-04*lvlp_saturation*lvlp_saturation+-1.61636e-02*lvlp_saturation+1.78800e-02'
+ sky130_fd_pr__pfet_01v8_lvt__a0_diff_7 = '-5.78194e-04*lvlp_saturation*lvlp_saturation+-1.24393e-02*lvlp_saturation+6.49640e-02'
+ sky130_fd_pr__pfet_01v8_lvt__a0_diff_8 = '-3.56519e-04*lvlp_saturation*lvlp_saturation+-1.03186e-02*lvlp_saturation+5.33830e-02'
+ sky130_fd_pr__pfet_01v8_lvt__a0_diff_9 = '-2.81656e-04*lvlp_saturation*lvlp_saturation+-5.69188e-03*lvlp_saturation+7.30880e-02'
+ sky130_fd_pr__pfet_01v8_lvt__ags_diff_0 = '1.41275e-03*lvlp_saturation*lvlp_saturation+5.62615e-02*lvlp_saturation+1.74640e-01'
+ sky130_fd_pr__pfet_01v8_lvt__ags_diff_1 = '-2.77812e-04*lvlp_saturation*lvlp_saturation+3.50738e-02*lvlp_saturation+1.29380e-01'
+ sky130_fd_pr__pfet_01v8_lvt__ags_diff_10 = '1.79937e-04*lvlp_saturation*lvlp_saturation+2.49228e-02*lvlp_saturation+1.19260e-01'
+ sky130_fd_pr__pfet_01v8_lvt__ags_diff_13 = '1.78416e-03*lvlp_saturation*lvlp_saturation+5.11221e-02*lvlp_saturation+8.51250e-02'
+ sky130_fd_pr__pfet_01v8_lvt__ags_diff_14 = '4.30875e-04*lvlp_saturation*lvlp_saturation+4.75062e-02*lvlp_saturation+7.88110e-02'
+ sky130_fd_pr__pfet_01v8_lvt__ags_diff_15 = '1.57984e-03*lvlp_saturation*lvlp_saturation+4.85781e-02*lvlp_saturation+1.01360e-01'
+ sky130_fd_pr__pfet_01v8_lvt__ags_diff_16 = '2.39406e-04*lvlp_saturation*lvlp_saturation+2.60261e-02*lvlp_saturation+8.36850e-02'
+ sky130_fd_pr__pfet_01v8_lvt__ags_diff_17 = '8.39125e-05*lvlp_saturation*lvlp_saturation+2.32446e-02*lvlp_saturation+9.49890e-02'
+ sky130_fd_pr__pfet_01v8_lvt__ags_diff_2 = '1.45200e-03*lvlp_saturation*lvlp_saturation+4.78838e-02*lvlp_saturation+6.75030e-02'
+ sky130_fd_pr__pfet_01v8_lvt__ags_diff_20 = '5.39187e-04*lvlp_saturation*lvlp_saturation+4.35557e-02*lvlp_saturation+1.81470e-01'
+ sky130_fd_pr__pfet_01v8_lvt__ags_diff_21 = '2.25400e-03*lvlp_saturation*lvlp_saturation+6.95915e-02*lvlp_saturation+2.13090e-01'
+ sky130_fd_pr__pfet_01v8_lvt__ags_diff_22 = '1.00750e-03*lvlp_saturation*lvlp_saturation+3.65400e-02*lvlp_saturation+2.19510e-01'
+ sky130_fd_pr__pfet_01v8_lvt__ags_diff_23 = '2.10219e-04*lvlp_saturation*lvlp_saturation+2.70881e-02*lvlp_saturation+4.99240e-02'
+ sky130_fd_pr__pfet_01v8_lvt__ags_diff_24 = '2.45969e-04*lvlp_saturation*lvlp_saturation+2.63671e-02*lvlp_saturation+6.83560e-02'
+ sky130_fd_pr__pfet_01v8_lvt__ags_diff_3 = '2.37463e-03*lvlp_saturation*lvlp_saturation+5.29615e-02*lvlp_saturation+1.15910e-01'
+ sky130_fd_pr__pfet_01v8_lvt__ags_diff_6 = '3.99063e-04*lvlp_saturation*lvlp_saturation+3.83063e-02*lvlp_saturation+2.64260e-01'
+ sky130_fd_pr__pfet_01v8_lvt__ags_diff_7 = '8.63562e-04*lvlp_saturation*lvlp_saturation+4.47207e-02*lvlp_saturation+2.30410e-01'
+ sky130_fd_pr__pfet_01v8_lvt__ags_diff_8 = '4.91250e-04*lvlp_saturation*lvlp_saturation+3.47925e-02*lvlp_saturation+2.03510e-01'
+ sky130_fd_pr__pfet_01v8_lvt__ags_diff_9 = '4.49250e-04*lvlp_saturation*lvlp_saturation+2.97730e-02*lvlp_saturation+1.88030e-01'
+ sky130_fd_pr__pfet_01v8_lvt__ajunction_mult = '-3.12500e-07*lvp_diode*lvp_diode+2.36612e-02*lvp_diode+9.96260e-01'
+ sky130_fd_pr__pfet_01v8_lvt__b0_diff_12 = '-4.54063e-10*lvlp_saturation*lvlp_saturation+-2.23634e-07*lvlp_saturation+-1.09850e-06'
+ sky130_fd_pr__pfet_01v8_lvt__b0_diff_19 = '1.51469e-09*lvlp_saturation*lvlp_saturation+-4.14259e-07*lvlp_saturation+-1.24070e-06'
+ sky130_fd_pr__pfet_01v8_lvt__b0_diff_26 = '-1.58431e-08*lvlp_saturation*lvlp_saturation+-2.28520e-07*lvlp_saturation+-7.38830e-07'
+ sky130_fd_pr__pfet_01v8_lvt__b0_diff_27 = '-8.30000e-10*lvlp_saturation*lvlp_saturation+-9.04525e-08*lvlp_saturation+-1.60460e-07'
+ sky130_fd_pr__pfet_01v8_lvt__b0_diff_28 = '2.57816e-09*lvlp_saturation*lvlp_saturation+-2.62976e-08*lvlp_saturation+-1.30140e-07'
+ sky130_fd_pr__pfet_01v8_lvt__b0_diff_29 = '2.89312e-09*lvlp_saturation*lvlp_saturation+-4.48850e-08*lvlp_saturation+-1.10830e-07'
+ sky130_fd_pr__pfet_01v8_lvt__b0_diff_30 = '2.64194e-09*lvlp_saturation*lvlp_saturation+-3.62802e-08*lvlp_saturation+-1.22600e-07'
+ sky130_fd_pr__pfet_01v8_lvt__b0_diff_31 = '1.74688e-09*lvlp_saturation*lvlp_saturation+-4.30550e-08*lvlp_saturation+-5.34000e-08'
+ sky130_fd_pr__pfet_01v8_lvt__b0_diff_33 = '2.10687e-09*lvlp_saturation*lvlp_saturation+-7.58525e-08*lvlp_saturation+-1.89610e-07'
+ sky130_fd_pr__pfet_01v8_lvt__b0_diff_34 = '1.44625e-09*lvlp_saturation*lvlp_saturation+-9.36075e-08*lvlp_saturation+-7.52000e-08'
+ sky130_fd_pr__pfet_01v8_lvt__b0_diff_35 = '2.51906e-09*lvlp_saturation*lvlp_saturation+-6.28063e-08*lvlp_saturation+-1.05030e-07'
+ sky130_fd_pr__pfet_01v8_lvt__b0_diff_36 = '1.39438e-09*lvlp_saturation*lvlp_saturation+-8.79625e-08*lvlp_saturation+-1.48220e-07'
+ sky130_fd_pr__pfet_01v8_lvt__b0_diff_37 = '2.11537e-09*lvlp_saturation*lvlp_saturation+-5.60125e-08*lvlp_saturation+-8.38960e-08'
+ sky130_fd_pr__pfet_01v8_lvt__b0_diff_39 = '9.30438e-09*lvlp_saturation*lvlp_saturation+-6.72900e-08*lvlp_saturation+-1.79310e-07'
+ sky130_fd_pr__pfet_01v8_lvt__b0_diff_4 = '-3.56156e-10*lvlp_saturation*lvlp_saturation+-5.61004e-08*lvlp_saturation+-1.75460e-07'
+ sky130_fd_pr__pfet_01v8_lvt__b0_diff_5 = '-2.94813e-09*lvlp_saturation*lvlp_saturation+-1.48538e-07*lvlp_saturation+-1.10200e-07'
+ sky130_fd_pr__pfet_01v8_lvt__b1_diff_27 = '2.18125e-09*lvlp_saturation*lvlp_saturation+6.11250e-09*lvlp_saturation+4.40490e-07'
+ sky130_fd_pr__pfet_01v8_lvt__b1_diff_28 = '1.81250e-11*lvlp_saturation*lvlp_saturation+-7.27250e-09*lvlp_saturation+2.28950e-07'
+ sky130_fd_pr__pfet_01v8_lvt__b1_diff_29 = '-1.24500e-09*lvlp_saturation*lvlp_saturation+-2.70750e-09*lvlp_saturation+2.27840e-07'
+ sky130_fd_pr__pfet_01v8_lvt__b1_diff_30 = '-2.72594e-09*lvlp_saturation*lvlp_saturation+-4.95375e-09*lvlp_saturation+2.48210e-07'
+ sky130_fd_pr__pfet_01v8_lvt__b1_diff_31 = '-1.93312e-09*lvlp_saturation*lvlp_saturation+2.91250e-09*lvlp_saturation+2.26990e-07'
+ sky130_fd_pr__pfet_01v8_lvt__b1_diff_33 = '-1.25000e-12*lvlp_saturation*lvlp_saturation+4.17500e-10*lvlp_saturation+2.11680e-07'
+ sky130_fd_pr__pfet_01v8_lvt__b1_diff_34 = '9.78125e-09*lvlp_saturation*lvlp_saturation+-6.61744e-24*lvlp_saturation+3.43500e-07'
+ sky130_fd_pr__pfet_01v8_lvt__b1_diff_35 = '-4.44687e-10*lvlp_saturation*lvlp_saturation+-3.55375e-09*lvlp_saturation+2.02970e-07'
+ sky130_fd_pr__pfet_01v8_lvt__b1_diff_36 = '-8.00625e-10*lvlp_saturation*lvlp_saturation+-3.45250e-09*lvlp_saturation+2.02280e-07'
+ sky130_fd_pr__pfet_01v8_lvt__b1_diff_37 = '-1.43750e-11*lvlp_saturation*lvlp_saturation+-2.05750e-09*lvlp_saturation+2.04180e-07'
+ sky130_fd_pr__pfet_01v8_lvt__b1_diff_39 = '-1.07792e-08*lvlp_saturation*lvlp_saturation+-3.59516e-08*lvlp_saturation+4.11800e-07'
+ sky130_fd_pr__pfet_01v8_lvt__b1_diff_4 = '-1.39625e-09*lvlp_saturation*lvlp_saturation+-4.93250e-09*lvlp_saturation+2.05850e-07'
+ sky130_fd_pr__pfet_01v8_lvt__b1_diff_5 = '2.32575e-08*lvlp_saturation*lvlp_saturation+4.55000e-10*lvlp_saturation+1.11810e-07'
+ sky130_fd_pr__pfet_01v8_lvt__dlc_diff = '-5.03437e-11*poly_cd*poly_cd+-1.17439e-08*poly_cd+-1.20000e-08'
+ sky130_fd_pr__pfet_01v8_lvt__dwc_diff = '8.04375e-09*diff_cd'
+ sky130_fd_pr__pfet_01v8_lvt__k2_diff_0 = '3.76031e-04*lvlp_bodyeffect*lvlp_bodyeffect+-1.58067e-02*lvlp_bodyeffect+7.10150e-03'
+ sky130_fd_pr__pfet_01v8_lvt__k2_diff_1 = '2.65721e-04*lvlp_bodyeffect*lvlp_bodyeffect+-1.09444e-02*lvlp_bodyeffect+-3.04030e-04'
+ sky130_fd_pr__pfet_01v8_lvt__k2_diff_10 = '2.66913e-04*lvlp_bodyeffect*lvlp_bodyeffect+-1.02802e-02*lvlp_bodyeffect+1.45140e-03'
+ sky130_fd_pr__pfet_01v8_lvt__k2_diff_11 = '3.41338e-04*lvlp_bodyeffect*lvlp_bodyeffect+-1.21610e-02*lvlp_bodyeffect+7.86360e-03'
+ sky130_fd_pr__pfet_01v8_lvt__k2_diff_12 = '1.90619e-04*lvlp_bodyeffect*lvlp_bodyeffect+-8.40800e-03*lvlp_bodyeffect+-4.61910e-04'
+ sky130_fd_pr__pfet_01v8_lvt__k2_diff_13 = '3.87894e-04*lvlp_bodyeffect*lvlp_bodyeffect+-1.17699e-02*lvlp_bodyeffect+-2.22800e-04'
+ sky130_fd_pr__pfet_01v8_lvt__k2_diff_14 = '2.61592e-04*lvlp_bodyeffect*lvlp_bodyeffect+-1.10719e-02*lvlp_bodyeffect+2.11020e-04'
+ sky130_fd_pr__pfet_01v8_lvt__k2_diff_15 = '4.36175e-04*lvlp_bodyeffect*lvlp_bodyeffect+-1.35081e-02*lvlp_bodyeffect+1.21370e-03'
+ sky130_fd_pr__pfet_01v8_lvt__k2_diff_16 = '3.72731e-04*lvlp_bodyeffect*lvlp_bodyeffect+-1.35305e-02*lvlp_bodyeffect+1.96730e-03'
+ sky130_fd_pr__pfet_01v8_lvt__k2_diff_17 = '3.07275e-04*lvlp_bodyeffect*lvlp_bodyeffect+-1.10043e-02*lvlp_bodyeffect+2.51260e-03'
+ sky130_fd_pr__pfet_01v8_lvt__k2_diff_18 = '2.89144e-04*lvlp_bodyeffect*lvlp_bodyeffect+-1.11160e-02*lvlp_bodyeffect+3.58570e-03'
+ sky130_fd_pr__pfet_01v8_lvt__k2_diff_19 = '2.13750e-04*lvlp_bodyeffect*lvlp_bodyeffect+-8.96537e-03*lvlp_bodyeffect+-3.68750e-03'
+ sky130_fd_pr__pfet_01v8_lvt__k2_diff_2 = '2.67806e-04*lvlp_bodyeffect*lvlp_bodyeffect+-1.06950e-02*lvlp_bodyeffect+4.50810e-03'
+ sky130_fd_pr__pfet_01v8_lvt__k2_diff_20 = '2.58637e-04*lvlp_bodyeffect*lvlp_bodyeffect+-1.06519e-02*lvlp_bodyeffect+-7.49970e-03'
+ sky130_fd_pr__pfet_01v8_lvt__k2_diff_21 = '3.21569e-04*lvlp_bodyeffect*lvlp_bodyeffect+-1.53447e-02*lvlp_bodyeffect+-3.30810e-03'
+ sky130_fd_pr__pfet_01v8_lvt__k2_diff_22 = '3.62225e-04*lvlp_bodyeffect*lvlp_bodyeffect+-1.72476e-02*lvlp_bodyeffect+-5.41510e-03'
+ sky130_fd_pr__pfet_01v8_lvt__k2_diff_23 = '3.15937e-04*lvlp_bodyeffect*lvlp_bodyeffect+-1.15916e-02*lvlp_bodyeffect+1.62950e-03'
+ sky130_fd_pr__pfet_01v8_lvt__k2_diff_24 = '3.25196e-04*lvlp_bodyeffect*lvlp_bodyeffect+-1.12300e-02*lvlp_bodyeffect+5.13870e-04'
+ sky130_fd_pr__pfet_01v8_lvt__k2_diff_25 = '2.81900e-04*lvlp_bodyeffect*lvlp_bodyeffect+-1.08309e-02*lvlp_bodyeffect+1.42710e-03'
+ sky130_fd_pr__pfet_01v8_lvt__k2_diff_26 = '2.01863e-04*lvlp_bodyeffect*lvlp_bodyeffect+-9.78863e-03*lvlp_bodyeffect+-4.43630e-03'
+ sky130_fd_pr__pfet_01v8_lvt__k2_diff_27 = '4.33319e-04*lvlp_bodyeffect*lvlp_bodyeffect+-1.85039e-02*lvlp_bodyeffect+-7.96860e-03'
+ sky130_fd_pr__pfet_01v8_lvt__k2_diff_28 = '2.29763e-04*lvlp_bodyeffect*lvlp_bodyeffect+-7.19775e-03*lvlp_bodyeffect+-6.20320e-03'
+ sky130_fd_pr__pfet_01v8_lvt__k2_diff_29 = '3.33919e-04*lvlp_bodyeffect*lvlp_bodyeffect+-1.11314e-02*lvlp_bodyeffect+-7.16320e-03'
+ sky130_fd_pr__pfet_01v8_lvt__k2_diff_3 = '3.00675e-04*lvlp_bodyeffect*lvlp_bodyeffect+-1.24371e-02*lvlp_bodyeffect+-1.24030e-03'
+ sky130_fd_pr__pfet_01v8_lvt__k2_diff_30 = '3.27956e-04*lvlp_bodyeffect*lvlp_bodyeffect+-1.15346e-02*lvlp_bodyeffect+-5.55780e-03'
+ sky130_fd_pr__pfet_01v8_lvt__k2_diff_31 = '3.37419e-04*lvlp_bodyeffect*lvlp_bodyeffect+-1.18815e-02*lvlp_bodyeffect+-3.79770e-03'
+ sky130_fd_pr__pfet_01v8_lvt__k2_diff_32 = '4.26356e-04*lvlp_bodyeffect*lvlp_bodyeffect+-1.38191e-02*lvlp_bodyeffect+8.04180e-03'
+ sky130_fd_pr__pfet_01v8_lvt__k2_diff_33 = '4.05219e-04*lvlp_bodyeffect*lvlp_bodyeffect+-1.42134e-02*lvlp_bodyeffect+-1.27860e-02'
+ sky130_fd_pr__pfet_01v8_lvt__k2_diff_34 = '3.87669e-04*lvlp_bodyeffect*lvlp_bodyeffect+-1.67144e-02*lvlp_bodyeffect+1.65480e-03'
+ sky130_fd_pr__pfet_01v8_lvt__k2_diff_35 = '3.97344e-04*lvlp_bodyeffect*lvlp_bodyeffect+-1.17296e-02*lvlp_bodyeffect+1.17720e-02'
+ sky130_fd_pr__pfet_01v8_lvt__k2_diff_36 = '3.62375e-04*lvlp_bodyeffect*lvlp_bodyeffect+-1.30607e-02*lvlp_bodyeffect+1.18670e-02'
+ sky130_fd_pr__pfet_01v8_lvt__k2_diff_37 = '2.68981e-04*lvlp_bodyeffect*lvlp_bodyeffect+-9.54663e-03*lvlp_bodyeffect+9.06380e-03'
+ sky130_fd_pr__pfet_01v8_lvt__k2_diff_38 = '3.81869e-04*lvlp_bodyeffect*lvlp_bodyeffect+-1.38899e-02*lvlp_bodyeffect+-5.54940e-03'
+ sky130_fd_pr__pfet_01v8_lvt__k2_diff_39 = '4.18594e-04*lvlp_bodyeffect*lvlp_bodyeffect+-1.46381e-02*lvlp_bodyeffect+-1.91370e-02'
+ sky130_fd_pr__pfet_01v8_lvt__k2_diff_4 = '5.61625e-04*lvlp_bodyeffect*lvlp_bodyeffect+-1.79358e-02*lvlp_bodyeffect+-1.16570e-02'
+ sky130_fd_pr__pfet_01v8_lvt__k2_diff_5 = '4.23131e-04*lvlp_bodyeffect*lvlp_bodyeffect+-1.50295e-02*lvlp_bodyeffect+-4.46210e-03'
+ sky130_fd_pr__pfet_01v8_lvt__k2_diff_6 = '2.65663e-04*lvlp_bodyeffect*lvlp_bodyeffect+-1.07644e-02*lvlp_bodyeffect+-1.99410e-03'
+ sky130_fd_pr__pfet_01v8_lvt__k2_diff_7 = '3.26912e-04*lvlp_bodyeffect*lvlp_bodyeffect+-1.65866e-02*lvlp_bodyeffect+1.10690e-03'
+ sky130_fd_pr__pfet_01v8_lvt__k2_diff_8 = '3.19563e-04*lvlp_bodyeffect*lvlp_bodyeffect+-1.20547e-02*lvlp_bodyeffect+1.51100e-03'
+ sky130_fd_pr__pfet_01v8_lvt__k2_diff_9 = '3.07606e-04*lvlp_bodyeffect*lvlp_bodyeffect+-1.16611e-02*lvlp_bodyeffect+5.48580e-03'
+ sky130_fd_pr__pfet_01v8_lvt__keta_diff_27 = '-2.50000e-04*lvlp_bodyeffect*lvlp_bodyeffect+1.00000e-03*lvlp_bodyeffect'
+ sky130_fd_pr__pfet_01v8_lvt__lint_diff = '-4.33125e-09*poly_cd'
+ sky130_fd_pr__pfet_01v8_lvt__overlap_mult = '-6.25000e-03*lvtox*lvtox+2.00000e-01'
+ sky130_fd_pr__pfet_01v8_lvt__pjunction_mult = '-1.57187e-04*lvp_diode*lvp_diode+2.31288e-02*lvp_diode+1.00090e+00'
+ sky130_fd_pr__pfet_01v8_lvt__toxe_mult = '1.30000e-02*lvtox+1.00000e+00'
+ sky130_fd_pr__pfet_01v8_lvt__u0_diff_0 = '-2.91850e-06*lvlp_mobility*lvlp_mobility+3.91413e-05*lvlp_mobility+2.14510e-05'
+ sky130_fd_pr__pfet_01v8_lvt__u0_diff_1 = '-3.48622e-06*lvlp_mobility*lvlp_mobility+1.99174e-05*lvlp_mobility+2.09090e-05'
+ sky130_fd_pr__pfet_01v8_lvt__u0_diff_10 = '3.79687e-07*lvlp_mobility*lvlp_mobility+7.00862e-05*lvlp_mobility+-1.58050e-04'
+ sky130_fd_pr__pfet_01v8_lvt__u0_diff_11 = '-2.21250e-07*lvlp_mobility*lvlp_mobility+1.07562e-04*lvlp_mobility+-1.93990e-04'
+ sky130_fd_pr__pfet_01v8_lvt__u0_diff_12 = '-1.27216e-06*lvlp_mobility*lvlp_mobility+7.40139e-05*lvlp_mobility+-2.37000e-04'
+ sky130_fd_pr__pfet_01v8_lvt__u0_diff_13 = '-9.19813e-07*lvlp_mobility*lvlp_mobility+6.83350e-05*lvlp_mobility+-8.10630e-05'
+ sky130_fd_pr__pfet_01v8_lvt__u0_diff_14 = '-3.62762e-07*lvlp_mobility*lvlp_mobility+6.78938e-05*lvlp_mobility+9.42920e-06'
+ sky130_fd_pr__pfet_01v8_lvt__u0_diff_15 = '2.06831e-06*lvlp_mobility*lvlp_mobility+1.00615e-04*lvlp_mobility+-6.66930e-05'
+ sky130_fd_pr__pfet_01v8_lvt__u0_diff_16 = '7.49563e-07*lvlp_mobility*lvlp_mobility+7.17137e-05*lvlp_mobility+-7.49380e-05'
+ sky130_fd_pr__pfet_01v8_lvt__u0_diff_17 = '5.43000e-07*lvlp_mobility*lvlp_mobility+6.69038e-05*lvlp_mobility+-9.60030e-05'
+ sky130_fd_pr__pfet_01v8_lvt__u0_diff_18 = '-2.01500e-06*lvlp_mobility*lvlp_mobility+7.45837e-05*lvlp_mobility+-7.13750e-05'
+ sky130_fd_pr__pfet_01v8_lvt__u0_diff_19 = '-3.97750e-07*lvlp_mobility*lvlp_mobility+9.28112e-05*lvlp_mobility+-2.10010e-05'
+ sky130_fd_pr__pfet_01v8_lvt__u0_diff_2 = '-3.40103e-06*lvlp_mobility*lvlp_mobility+1.68986e-05*lvlp_mobility+-7.56190e-05'
+ sky130_fd_pr__pfet_01v8_lvt__u0_diff_20 = '3.19313e-07*lvlp_mobility*lvlp_mobility+7.43850e-05*lvlp_mobility+-2.38890e-05'
+ sky130_fd_pr__pfet_01v8_lvt__u0_diff_21 = '1.91250e-08*lvlp_mobility*lvlp_mobility+8.09300e-05*lvlp_mobility+-2.31860e-05'
+ sky130_fd_pr__pfet_01v8_lvt__u0_diff_22 = '3.96525e-07*lvlp_mobility*lvlp_mobility+7.00050e-05*lvlp_mobility+7.33560e-06'
+ sky130_fd_pr__pfet_01v8_lvt__u0_diff_23 = '7.75125e-07*lvlp_mobility*lvlp_mobility+7.33875e-05*lvlp_mobility+-1.81220e-05'
+ sky130_fd_pr__pfet_01v8_lvt__u0_diff_24 = '6.91631e-07*lvlp_mobility*lvlp_mobility+7.22350e-05*lvlp_mobility+8.28390e-06'
+ sky130_fd_pr__pfet_01v8_lvt__u0_diff_25 = '-1.64006e-06*lvlp_mobility*lvlp_mobility+9.23962e-05*lvlp_mobility+1.33360e-05'
+ sky130_fd_pr__pfet_01v8_lvt__u0_diff_26 = '-8.71312e-07*lvlp_mobility*lvlp_mobility+7.67550e-05*lvlp_mobility+-4.05590e-05'
+ sky130_fd_pr__pfet_01v8_lvt__u0_diff_27 = '-3.90041e-06*lvlp_mobility*lvlp_mobility+8.82041e-05*lvlp_mobility+4.86410e-04'
+ sky130_fd_pr__pfet_01v8_lvt__u0_diff_28 = '-1.96422e-06*lvlp_mobility*lvlp_mobility+4.34731e-05*lvlp_mobility+-7.10100e-05'
+ sky130_fd_pr__pfet_01v8_lvt__u0_diff_29 = '-2.95938e-06*lvlp_mobility*lvlp_mobility+5.69550e-05*lvlp_mobility+1.22300e-05'
+ sky130_fd_pr__pfet_01v8_lvt__u0_diff_3 = '-3.18813e-06*lvlp_mobility*lvlp_mobility+1.98580e-05*lvlp_mobility+1.71820e-05'
+ sky130_fd_pr__pfet_01v8_lvt__u0_diff_30 = '-6.73813e-07*lvlp_mobility*lvlp_mobility+7.65950e-05*lvlp_mobility+6.23910e-05'
+ sky130_fd_pr__pfet_01v8_lvt__u0_diff_31 = '-7.25938e-07*lvlp_mobility*lvlp_mobility+6.91713e-05*lvlp_mobility+-3.48900e-05'
+ sky130_fd_pr__pfet_01v8_lvt__u0_diff_32 = '-6.08225e-06*lvlp_mobility*lvlp_mobility+5.02625e-05*lvlp_mobility+2.76960e-05'
+ sky130_fd_pr__pfet_01v8_lvt__u0_diff_33 = '-2.85212e-06*lvlp_mobility*lvlp_mobility+9.85213e-05*lvlp_mobility+4.02890e-05'
+ sky130_fd_pr__pfet_01v8_lvt__u0_diff_34 = '-2.94862e-06*lvlp_mobility*lvlp_mobility+6.23637e-05*lvlp_mobility+3.36030e-05'
+ sky130_fd_pr__pfet_01v8_lvt__u0_diff_35 = '-2.58381e-06*lvlp_mobility*lvlp_mobility+4.77437e-05*lvlp_mobility+3.58460e-05'
+ sky130_fd_pr__pfet_01v8_lvt__u0_diff_36 = '-1.70012e-06*lvlp_mobility*lvlp_mobility+4.85238e-05*lvlp_mobility+1.62690e-06'
+ sky130_fd_pr__pfet_01v8_lvt__u0_diff_37 = '-8.28500e-07*lvlp_mobility*lvlp_mobility+5.92450e-05*lvlp_mobility+-6.57400e-06'
+ sky130_fd_pr__pfet_01v8_lvt__u0_diff_38 = '-4.14438e-06*lvlp_mobility*lvlp_mobility+5.87075e-05*lvlp_mobility+1.08120e-04'
+ sky130_fd_pr__pfet_01v8_lvt__u0_diff_39 = '-3.90312e-07*lvlp_mobility*lvlp_mobility+1.15444e-04*lvlp_mobility+3.52710e-04'
+ sky130_fd_pr__pfet_01v8_lvt__u0_diff_4 = '-3.21587e-06*lvlp_mobility*lvlp_mobility+8.12250e-05*lvlp_mobility+-7.07160e-05'
+ sky130_fd_pr__pfet_01v8_lvt__u0_diff_5 = '-3.00375e-07*lvlp_mobility*lvlp_mobility+8.43112e-05*lvlp_mobility+-2.48290e-05'
+ sky130_fd_pr__pfet_01v8_lvt__u0_diff_6 = '-2.14875e-07*lvlp_mobility*lvlp_mobility+5.99780e-05*lvlp_mobility+-1.69570e-04'
+ sky130_fd_pr__pfet_01v8_lvt__u0_diff_7 = '-9.55375e-07*lvlp_mobility*lvlp_mobility+6.85100e-05*lvlp_mobility+-1.44440e-05'
+ sky130_fd_pr__pfet_01v8_lvt__u0_diff_8 = '3.59531e-07*lvlp_mobility*lvlp_mobility+6.86356e-05*lvlp_mobility+-1.97920e-04'
+ sky130_fd_pr__pfet_01v8_lvt__u0_diff_9 = '2.11437e-07*lvlp_mobility*lvlp_mobility+6.37832e-05*lvlp_mobility+-1.93050e-04'
+ sky130_fd_pr__pfet_01v8_lvt__uc_diff_21 = '-2.25000e-12*lvlp_mobility'
+ sky130_fd_pr__pfet_01v8_lvt__uc_diff_22 = '1.25000e-13*lvlp_mobility*lvlp_mobility+-2.75000e-12*lvlp_mobility'
+ sky130_fd_pr__pfet_01v8_lvt__uc_diff_7 = '3.12500e-14*lvlp_mobility*lvlp_mobility+-2.37500e-12*lvlp_mobility'
+ sky130_fd_pr__pfet_01v8_lvt__vsat_diff_11 = '3.41459e+02*lvlp_saturation*lvlp_saturation+8.40266e+03*lvlp_saturation+1.89160e+04'
+ sky130_fd_pr__pfet_01v8_lvt__vsat_diff_12 = '-1.57203e+02*lvlp_saturation*lvlp_saturation+2.88109e+03*lvlp_saturation+-6.36840e+03'
+ sky130_fd_pr__pfet_01v8_lvt__vsat_diff_18 = '1.36739e+03*lvlp_saturation*lvlp_saturation+1.24566e+04*lvlp_saturation+8.29520e+03'
+ sky130_fd_pr__pfet_01v8_lvt__vsat_diff_19 = '-8.69000e+01*lvlp_saturation*lvlp_saturation+3.29415e+03*lvlp_saturation+-9.99700e+03'
+ sky130_fd_pr__pfet_01v8_lvt__vsat_diff_25 = '2.25753e+02*lvlp_saturation*lvlp_saturation+5.51474e+03*lvlp_saturation+1.07040e+04'
+ sky130_fd_pr__pfet_01v8_lvt__vsat_diff_26 = '2.25750e+02*lvlp_saturation*lvlp_saturation+8.90975e+03*lvlp_saturation+1.21240e+04'
+ sky130_fd_pr__pfet_01v8_lvt__vsat_diff_32 = '8.00250e+02*lvlp_saturation*lvlp_saturation+1.23778e+04*lvlp_saturation+1.50690e+04'
+ sky130_fd_pr__pfet_01v8_lvt__vsat_diff_33 = '-1.09156e+02*lvlp_saturation*lvlp_saturation+7.18625e+02*lvlp_saturation+-1.71610e+04'
+ sky130_fd_pr__pfet_01v8_lvt__vsat_diff_38 = '1.08434e+03*lvlp_saturation*lvlp_saturation+1.13641e+04*lvlp_saturation+1.71940e+04'
+ sky130_fd_pr__pfet_01v8_lvt__vsat_diff_39 = '5.85906e+02*lvlp_saturation*lvlp_saturation+5.33788e+03*lvlp_saturation+-1.56260e+04'
+ sky130_fd_pr__pfet_01v8_lvt__vsat_diff_4 = '8.70812e+02*lvlp_saturation*lvlp_saturation+1.00090e+04*lvlp_saturation+1.60310e+04'
+ sky130_fd_pr__pfet_01v8_lvt__vsat_diff_5 = '-2.37781e+02*lvlp_saturation*lvlp_saturation+1.95288e+03*lvlp_saturation+-1.91870e+04'
+ sky130_fd_pr__pfet_01v8_lvt__vth0_diff_0 = '5.17875e-04*lvlp_threshold*lvlp_threshold+-3.56763e-02*lvlp_threshold+-4.54710e-02'
+ sky130_fd_pr__pfet_01v8_lvt__vth0_diff_1 = '4.52875e-04*lvlp_threshold*lvlp_threshold+-2.92138e-02*lvlp_threshold+-1.32210e-02'
+ sky130_fd_pr__pfet_01v8_lvt__vth0_diff_10 = '3.46263e-04*lvlp_threshold*lvlp_threshold+-3.32750e-02*lvlp_threshold+-9.77020e-03'
+ sky130_fd_pr__pfet_01v8_lvt__vth0_diff_11 = '2.43062e-04*lvlp_threshold*lvlp_threshold+-3.44678e-02*lvlp_threshold+-4.75880e-02'
+ sky130_fd_pr__pfet_01v8_lvt__vth0_diff_12 = '2.93875e-04*lvlp_threshold*lvlp_threshold+-3.15875e-02*lvlp_threshold+-2.94720e-02'
+ sky130_fd_pr__pfet_01v8_lvt__vth0_diff_13 = '6.26688e-04*lvlp_threshold*lvlp_threshold+-3.38725e-02*lvlp_threshold+-2.45370e-02'
+ sky130_fd_pr__pfet_01v8_lvt__vth0_diff_14 = '2.91219e-04*lvlp_threshold*lvlp_threshold+-2.90014e-02*lvlp_threshold+-3.27340e-02'
+ sky130_fd_pr__pfet_01v8_lvt__vth0_diff_15 = '6.33687e-04*lvlp_threshold*lvlp_threshold+-4.28763e-02*lvlp_threshold+-2.80440e-02'
+ sky130_fd_pr__pfet_01v8_lvt__vth0_diff_16 = '4.42437e-04*lvlp_threshold*lvlp_threshold+-3.63513e-02*lvlp_threshold+-2.02940e-02'
+ sky130_fd_pr__pfet_01v8_lvt__vth0_diff_17 = '4.06250e-04*lvlp_threshold*lvlp_threshold+-3.43325e-02*lvlp_threshold+-1.38600e-02'
+ sky130_fd_pr__pfet_01v8_lvt__vth0_diff_18 = '1.58031e-04*lvlp_threshold*lvlp_threshold+-3.37189e-02*lvlp_threshold+-6.63030e-02'
+ sky130_fd_pr__pfet_01v8_lvt__vth0_diff_19 = '3.19406e-04*lvlp_threshold*lvlp_threshold+-3.41991e-02*lvlp_threshold+-5.77840e-02'
+ sky130_fd_pr__pfet_01v8_lvt__vth0_diff_2 = '4.71788e-04*lvlp_threshold*lvlp_threshold+-3.02800e-02*lvlp_threshold+-9.60860e-03'
+ sky130_fd_pr__pfet_01v8_lvt__vth0_diff_20 = '3.03813e-04*lvlp_threshold*lvlp_threshold+-3.18275e-02*lvlp_threshold+-4.30410e-02'
+ sky130_fd_pr__pfet_01v8_lvt__vth0_diff_21 = '2.54625e-04*lvlp_threshold*lvlp_threshold+-3.09997e-02*lvlp_threshold+-4.43650e-02'
+ sky130_fd_pr__pfet_01v8_lvt__vth0_diff_22 = '2.67281e-04*lvlp_threshold*lvlp_threshold+-3.18586e-02*lvlp_threshold+-4.52420e-02'
+ sky130_fd_pr__pfet_01v8_lvt__vth0_diff_23 = '3.97438e-04*lvlp_threshold*lvlp_threshold+-3.48975e-02*lvlp_threshold+-2.30690e-02'
+ sky130_fd_pr__pfet_01v8_lvt__vth0_diff_24 = '4.46187e-04*lvlp_threshold*lvlp_threshold+-3.59675e-02*lvlp_threshold+-3.25090e-02'
+ sky130_fd_pr__pfet_01v8_lvt__vth0_diff_25 = '1.19656e-04*lvlp_threshold*lvlp_threshold+-2.96494e-02*lvlp_threshold+-7.99170e-02'
+ sky130_fd_pr__pfet_01v8_lvt__vth0_diff_26 = '1.84531e-04*lvlp_threshold*lvlp_threshold+-2.89846e-02*lvlp_threshold+-4.51240e-02'
+ sky130_fd_pr__pfet_01v8_lvt__vth0_diff_27 = '7.55500e-04*lvlp_threshold*lvlp_threshold+-4.16640e-02*lvlp_threshold+-9.49120e-02'
+ sky130_fd_pr__pfet_01v8_lvt__vth0_diff_28 = '5.75644e-04*lvlp_threshold*lvlp_threshold+-2.05389e-02*lvlp_threshold+-2.79480e-03'
+ sky130_fd_pr__pfet_01v8_lvt__vth0_diff_29 = '7.73375e-04*lvlp_threshold*lvlp_threshold+-3.41075e-02*lvlp_threshold+-1.32340e-02'
+ sky130_fd_pr__pfet_01v8_lvt__vth0_diff_3 = '4.68875e-04*lvlp_threshold*lvlp_threshold+-3.24088e-02*lvlp_threshold+-2.39870e-02'
+ sky130_fd_pr__pfet_01v8_lvt__vth0_diff_30 = '6.33188e-04*lvlp_threshold*lvlp_threshold+-3.15025e-02*lvlp_threshold+-3.23110e-02'
+ sky130_fd_pr__pfet_01v8_lvt__vth0_diff_31 = '6.64781e-04*lvlp_threshold*lvlp_threshold+-3.45937e-02*lvlp_threshold+-1.48150e-03'
+ sky130_fd_pr__pfet_01v8_lvt__vth0_diff_32 = '7.74437e-04*lvlp_threshold*lvlp_threshold+-3.45092e-02*lvlp_threshold+2.95120e-02'
+ sky130_fd_pr__pfet_01v8_lvt__vth0_diff_33 = '9.04500e-04*lvlp_threshold*lvlp_threshold+-4.53725e-02*lvlp_threshold+-5.83420e-02'
+ sky130_fd_pr__pfet_01v8_lvt__vth0_diff_34 = '6.28200e-04*lvlp_threshold*lvlp_threshold+-3.77863e-02*lvlp_threshold+-8.76620e-03'
+ sky130_fd_pr__pfet_01v8_lvt__vth0_diff_35 = '8.36563e-04*lvlp_threshold*lvlp_threshold+-3.49337e-02*lvlp_threshold+-2.36500e-02'
+ sky130_fd_pr__pfet_01v8_lvt__vth0_diff_36 = '6.75000e-04*lvlp_threshold*lvlp_threshold+-3.60162e-02*lvlp_threshold+-2.64150e-02'
+ sky130_fd_pr__pfet_01v8_lvt__vth0_diff_37 = '5.20500e-04*lvlp_threshold*lvlp_threshold+-2.94825e-02*lvlp_threshold+-1.80880e-02'
+ sky130_fd_pr__pfet_01v8_lvt__vth0_diff_38 = '5.05906e-04*lvlp_threshold*lvlp_threshold+-3.75561e-02*lvlp_threshold+-1.05690e-01'
+ sky130_fd_pr__pfet_01v8_lvt__vth0_diff_39 = '7.66844e-04*lvlp_threshold*lvlp_threshold+-4.71574e-02*lvlp_threshold+-1.23640e-01'
+ sky130_fd_pr__pfet_01v8_lvt__vth0_diff_4 = '7.30562e-04*lvlp_threshold*lvlp_threshold+-4.94613e-02*lvlp_threshold+-9.38440e-02'
+ sky130_fd_pr__pfet_01v8_lvt__vth0_diff_5 = '7.42000e-04*lvlp_threshold*lvlp_threshold+-5.12263e-02*lvlp_threshold+-2.35270e-02'
+ sky130_fd_pr__pfet_01v8_lvt__vth0_diff_6 = '3.31250e-04*lvlp_threshold*lvlp_threshold+-3.16625e-02*lvlp_threshold+-4.31300e-02'
+ sky130_fd_pr__pfet_01v8_lvt__vth0_diff_7 = '2.51219e-04*lvlp_threshold*lvlp_threshold+-2.83526e-02*lvlp_threshold+-4.12290e-02'
+ sky130_fd_pr__pfet_01v8_lvt__vth0_diff_8 = '4.04938e-04*lvlp_threshold*lvlp_threshold+-3.55987e-02*lvlp_threshold+-1.48840e-02'
+ sky130_fd_pr__pfet_01v8_lvt__vth0_diff_9 = '3.94250e-04*lvlp_threshold*lvlp_threshold+-3.51837e-02*lvlp_threshold+-2.13030e-02'
+ sky130_fd_pr__pfet_01v8_lvt__wint_diff = '8.04375e-09*diff_cd'
+ sky130_fd_pr__pfet_01v8_mvt__ajunction_mult = '-3.12500e-07*lvp_diode*lvp_diode+2.36612e-02*lvp_diode+9.96260e-01'
+ sky130_fd_pr__pfet_01v8_mvt__dlc_diff = '-4.33125e-09*poly_cd'
+ sky130_fd_pr__pfet_01v8_mvt__dwc_diff = '8.04375e-09*diff_cd'
+ sky130_fd_pr__pfet_01v8_mvt__k2_diff_0 = '-9.21756e-03*lvp_bodyeffect*lvp_bodyeffect+4.31298e-02*lvp_bodyeffect'
+ sky130_fd_pr__pfet_01v8_mvt__k2_diff_1 = '-7.88292e-03*lvp_bodyeffect*lvp_bodyeffect+3.35458e-02*lvp_bodyeffect'
+ sky130_fd_pr__pfet_01v8_mvt__lint_diff = '-4.33125e-09*poly_cd'
+ sky130_fd_pr__pfet_01v8_mvt__overlap_mult = '7.47062e-03*lvtox*lvtox+2.98800e-02*lvtox+9.54350e-01'
+ sky130_fd_pr__pfet_01v8_mvt__pjunction_mult = '2.18750e-06*lvp_diode*lvp_diode+2.37662e-02*lvp_diode+1.00090e+00'
+ sky130_fd_pr__rf_pfet_01v8_mvt__aw_cap_mult = '3.75000e-02*pfet_01v8_mvt+1.00000e+00'
+ sky130_fd_pr__rf_pfet_01v8_mvt__aw_rgate_dist_mult = '6.25000e-03*pfet_01v8_mvt*pfet_01v8_mvt+8.75000e-02*pfet_01v8_mvt+1.00000e+00'
+ sky130_fd_pr__rf_pfet_01v8_mvt__aw_rgate_dist_mult_2 = '3.12500e-03*pfet_01v8_mvt*pfet_01v8_mvt+1.00000e-01*pfet_01v8_mvt+1.00000e+00'
+ sky130_fd_pr__rf_pfet_01v8_mvt__aw_rgate_stub_mult = '6.25000e-03*lvp_mobility*lvp_mobility+8.75000e-02*lvp_mobility+1.00000e+00'
+ sky130_fd_pr__rf_pfet_01v8_mvt__aw_rgate_stub_mult_2 = '3.12500e-03*lvp_mobility*lvp_mobility+1.00000e-01*lvp_mobility+1.00000e+00'
+ sky130_fd_pr__pfet_01v8_mvt__toxe_mult = '1.30000e-02*lvtox+1.00000e+00'
+ sky130_fd_pr__pfet_01v8_mvt__u0_diff_0 = '-9.56406e-06*lvp_mobility*lvp_mobility+-2.17375e-06*lvp_mobility'
+ sky130_fd_pr__pfet_01v8_mvt__u0_diff_1 = '-1.31759e-05*lvp_mobility*lvp_mobility+-7.05625e-06*lvp_mobility'
+ sky130_fd_pr__pfet_01v8_mvt__vsat_diff_0 = '1.90562e+02*lvp_saturation*lvp_saturation+4.51050e+03*lvp_saturation'
+ sky130_fd_pr__pfet_01v8_mvt__vsat_diff_1 = '1.04844e+02*lvp_saturation*lvp_saturation+3.88288e+03*lvp_saturation'
+ sky130_fd_pr__pfet_01v8_mvt__vth0_diff_0 = '-1.50000e-05*lvp_threshold*lvp_threshold+-2.82625e-02*lvp_threshold'
+ sky130_fd_pr__pfet_01v8_mvt__vth0_diff_1 = '2.57469e-03*lvp_threshold*lvp_threshold+-4.77988e-02*lvp_threshold'
+ sky130_fd_pr__pfet_01v8_mvt__wint_diff = '8.04375e-09*diff_cd'
+ sky130_fd_pr__special_pfet_pass__ajunction_mult = '2.33750e-04*lvp_diode*lvp_diode+-1.38778e-17*lvp_diode+9.96260e-01'
+ sky130_fd_pr__special_pfet_pass__overlap_mult = '2.85312e-03*lvtox*lvtox+9.54350e-01'
+ sky130_fd_pr__special_pfet_pass__pjunction_mult = '-5.62500e-05*lvp_diode*lvp_diode+1.00090e+00'
+ sky130_fd_pr__special_pfet_pass__u0_diff_0 = '-9.11563e-07*lvp_mobility*lvp_mobility+-2.98259e-04*lvp_mobility+-4.44680e-04'
+ sky130_fd_pr__special_pfet_pass__vth0_diff_0 = '8.09813e-05*lvp_threshold*lvp_threshold+-4.19525e-02*lvp_threshold+8.19430e-03'
+ sky130_fd_pr__pfet_01v8__a0_diff_11 = '3.15701e-03*lvp_saturation*lvp_saturation+1.06738e-02*lvp_saturation+-8.73550e-02'
+ sky130_fd_pr__pfet_01v8__a0_diff_12 = '2.62199e-03*lvp_saturation*lvp_saturation+7.72522e-03*lvp_saturation+-7.20230e-02'
+ sky130_fd_pr__pfet_01v8__a0_diff_13 = '1.62044e-03*lvp_saturation*lvp_saturation+1.99900e-03*lvp_saturation+-4.10370e-02'
+ sky130_fd_pr__pfet_01v8__a0_diff_14 = '1.77066e-03*lvp_saturation*lvp_saturation+4.73438e-03*lvp_saturation+-2.02150e-02'
+ sky130_fd_pr__pfet_01v8__a0_diff_19 = '3.01987e-04*lvp_saturation*lvp_saturation+1.11857e-02*lvp_saturation+-4.50260e-02'
+ sky130_fd_pr__pfet_01v8__a0_diff_2 = '7.36063e-03*lvp_saturation*lvp_saturation+8.85324e-03*lvp_saturation+-8.02300e-02'
+ sky130_fd_pr__pfet_01v8__a0_diff_20 = '1.67681e-03*lvp_saturation*lvp_saturation+-2.69000e-04*lvp_saturation+-3.97820e-02'
+ sky130_fd_pr__pfet_01v8__a0_diff_21 = '1.63154e-03*lvp_saturation*lvp_saturation+5.36284e-03*lvp_saturation+-1.28540e-02'
+ sky130_fd_pr__pfet_01v8__a0_diff_22 = '1.52681e-03*lvp_saturation*lvp_saturation+6.05850e-03*lvp_saturation+-1.15030e-02'
+ sky130_fd_pr__pfet_01v8__a0_diff_27 = '2.72275e-03*lvp_saturation*lvp_saturation+6.97350e-03*lvp_saturation+-1.34710e-01'
+ sky130_fd_pr__pfet_01v8__a0_diff_28 = '1.91247e-03*lvp_saturation*lvp_saturation+6.34238e-03*lvp_saturation+-6.67330e-02'
+ sky130_fd_pr__pfet_01v8__a0_diff_29 = '1.59591e-03*lvp_saturation*lvp_saturation+6.02988e-03*lvp_saturation+-1.91740e-02'
+ sky130_fd_pr__pfet_01v8__a0_diff_3 = '4.56485e-03*lvp_saturation*lvp_saturation+-3.42888e-04*lvp_saturation+-7.03840e-02'
+ sky130_fd_pr__pfet_01v8__a0_diff_30 = '1.81791e-03*lvp_saturation*lvp_saturation+1.69709e-02*lvp_saturation+1.68200e-02'
+ sky130_fd_pr__pfet_01v8__a0_diff_4 = '3.88384e-03*lvp_saturation*lvp_saturation+5.60190e-03*lvp_saturation+-4.43630e-02'
+ sky130_fd_pr__pfet_01v8__a0_diff_5 = '3.24284e-03*lvp_saturation*lvp_saturation+3.93888e-03*lvp_saturation+-8.15850e-02'
+ sky130_fd_pr__pfet_01v8__ags_diff_11 = '-2.29793e-03*lvp_saturation*lvp_saturation+-8.43549e-03*lvp_saturation+6.71700e-02'
+ sky130_fd_pr__pfet_01v8__ags_diff_12 = '-2.06099e-03*lvp_saturation*lvp_saturation+-6.76197e-03*lvp_saturation+6.02380e-02'
+ sky130_fd_pr__pfet_01v8__ags_diff_13 = '-1.34241e-03*lvp_saturation*lvp_saturation+-1.80038e-03*lvp_saturation+3.48810e-02'
+ sky130_fd_pr__pfet_01v8__ags_diff_14 = '-1.32793e-03*lvp_saturation*lvp_saturation+-3.59304e-03*lvp_saturation+1.57870e-02'
+ sky130_fd_pr__pfet_01v8__ags_diff_19 = '-1.05813e-05*lvp_saturation*lvp_saturation+-1.09251e-02*lvp_saturation+4.05640e-02'
+ sky130_fd_pr__pfet_01v8__ags_diff_2 = '-7.29072e-03*lvp_saturation*lvp_saturation+-8.15537e-03*lvp_saturation+8.19170e-02'
+ sky130_fd_pr__pfet_01v8__ags_diff_20 = '-1.43191e-03*lvp_saturation*lvp_saturation+1.34125e-04*lvp_saturation+3.42610e-02'
+ sky130_fd_pr__pfet_01v8__ags_diff_21 = '-1.32829e-03*lvp_saturation*lvp_saturation+-4.39635e-03*lvp_saturation+1.10090e-02'
+ sky130_fd_pr__pfet_01v8__ags_diff_22 = '-1.22639e-03*lvp_saturation*lvp_saturation+-4.99725e-03*lvp_saturation+9.94820e-03'
+ sky130_fd_pr__pfet_01v8__ags_diff_27 = '-1.76269e-03*lvp_saturation*lvp_saturation+-5.34150e-03*lvp_saturation+9.03960e-02'
+ sky130_fd_pr__pfet_01v8__ags_diff_28 = '-1.55645e-03*lvp_saturation*lvp_saturation+-5.85080e-03*lvp_saturation+5.73440e-02'
+ sky130_fd_pr__pfet_01v8__ags_diff_29 = '-1.25981e-03*lvp_saturation*lvp_saturation+-4.69175e-03*lvp_saturation+1.57690e-02'
+ sky130_fd_pr__pfet_01v8__ags_diff_3 = '-3.99271e-03*lvp_saturation*lvp_saturation+3.15875e-04*lvp_saturation+6.15440e-02'
+ sky130_fd_pr__pfet_01v8__ags_diff_30 = '-1.37472e-03*lvp_saturation*lvp_saturation+-1.41679e-02*lvp_saturation+-1.42480e-02'
+ sky130_fd_pr__pfet_01v8__ags_diff_4 = '-3.67510e-03*lvp_saturation*lvp_saturation+-5.25410e-03*lvp_saturation+4.29790e-02'
+ sky130_fd_pr__pfet_01v8__ags_diff_5 = '-3.36803e-03*lvp_saturation*lvp_saturation+-4.42138e-03*lvp_saturation+8.56250e-02'
+ sky130_fd_pr__pfet_01v8__ajunction_mult = '-3.12500e-07*lvp_diode*lvp_diode+2.36612e-02*lvp_diode+9.96260e-01'
+ sky130_fd_pr__pfet_01v8__b0_diff_35 = '3.58916e-09*lvp_saturation*lvp_saturation+1.14113e-09*lvp_saturation+-3.96030e-08'
+ sky130_fd_pr__pfet_01v8__b0_diff_36 = '2.04428e-09*lvp_saturation*lvp_saturation+-7.78339e-09*lvp_saturation+-7.36180e-08'
+ sky130_fd_pr__pfet_01v8__b0_diff_37 = '-2.05056e-09*lvp_saturation*lvp_saturation+-2.38137e-09*lvp_saturation+-7.14480e-10'
+ sky130_fd_pr__pfet_01v8__b0_diff_38 = '-1.76159e-09*lvp_saturation*lvp_saturation+6.94125e-10*lvp_saturation+-1.99090e-08'
+ sky130_fd_pr__pfet_01v8__b0_diff_39 = '2.20819e-09*lvp_saturation*lvp_saturation+-1.77613e-08*lvp_saturation+3.62140e-08'
+ sky130_fd_pr__pfet_01v8__b0_diff_40 = '9.46581e-09*lvp_saturation*lvp_saturation+-5.52987e-08*lvp_saturation+-5.06080e-08'
+ sky130_fd_pr__pfet_01v8__b0_diff_41 = '3.20806e-09*lvp_saturation*lvp_saturation+-6.03925e-09*lvp_saturation+-7.59860e-08'
+ sky130_fd_pr__pfet_01v8__b0_diff_42 = '4.56753e-09*lvp_saturation*lvp_saturation+-1.82788e-09*lvp_saturation+-4.35830e-08'
+ sky130_fd_pr__pfet_01v8__b0_diff_43 = '8.25928e-09*lvp_saturation*lvp_saturation+-7.63212e-09*lvp_saturation+-3.90870e-08'
+ sky130_fd_pr__pfet_01v8__b0_diff_44 = '4.05193e-09*lvp_saturation*lvp_saturation+2.41098e-09*lvp_saturation+-7.46750e-08'
+ sky130_fd_pr__pfet_01v8__b0_diff_45 = '9.15062e-10*lvp_saturation*lvp_saturation+-1.52822e-08*lvp_saturation+1.69120e-08'
+ sky130_fd_pr__pfet_01v8__b0_diff_46 = '3.01391e-09*lvp_saturation*lvp_saturation+-1.42113e-09*lvp_saturation+-7.52160e-08'
+ sky130_fd_pr__pfet_01v8__b0_diff_47 = '1.47652e-08*lvp_saturation*lvp_saturation+-1.04270e-07*lvp_saturation+2.69470e-08'
+ sky130_fd_pr__pfet_01v8__b0_diff_48 = '5.02447e-09*lvp_saturation*lvp_saturation+-3.05513e-09*lvp_saturation+-6.82210e-08'
+ sky130_fd_pr__pfet_01v8__b0_diff_49 = '1.53625e-08*lvp_saturation*lvp_saturation+-1.21745e-07*lvp_saturation+1.36730e-07'
+ sky130_fd_pr__pfet_01v8__b1_diff_35 = '1.83845e-09*lvp_saturation*lvp_saturation+5.01975e-09*lvp_saturation+9.65870e-10'
+ sky130_fd_pr__pfet_01v8__b1_diff_36 = '2.61900e-10*lvp_saturation*lvp_saturation+8.95750e-10*lvp_saturation+1.87010e-09'
+ sky130_fd_pr__pfet_01v8__b1_diff_37 = '5.42668e-10*lvp_saturation*lvp_saturation+6.72862e-10*lvp_saturation+7.96860e-10'
+ sky130_fd_pr__pfet_01v8__b1_diff_38 = '1.52752e-10*lvp_saturation*lvp_saturation+3.65238e-10*lvp_saturation+1.73020e-10'
+ sky130_fd_pr__pfet_01v8__b1_diff_39 = '-2.93809e-10*lvp_saturation*lvp_saturation+4.19690e-10*lvp_saturation+3.37030e-09'
+ sky130_fd_pr__pfet_01v8__b1_diff_40 = '8.40006e-10*lvp_saturation*lvp_saturation+-1.12613e-09*lvp_saturation+2.64140e-09'
+ sky130_fd_pr__pfet_01v8__b1_diff_41 = '-6.49602e-10*lvp_saturation*lvp_saturation+-8.10442e-10*lvp_saturation+7.22730e-09'
+ sky130_fd_pr__pfet_01v8__b1_diff_42 = '-3.27580e-10*lvp_saturation*lvp_saturation+3.73956e-10*lvp_saturation+4.45920e-09'
+ sky130_fd_pr__pfet_01v8__b1_diff_43 = '-7.83652e-11*lvp_saturation*lvp_saturation+2.03770e-10*lvp_saturation+-5.01760e-11'
+ sky130_fd_pr__pfet_01v8__b1_diff_44 = '-6.41406e-13*lvp_saturation*lvp_saturation+-3.50906e-11*lvp_saturation+2.28950e-10'
+ sky130_fd_pr__pfet_01v8__b1_diff_45 = '-1.39303e-11*lvp_saturation*lvp_saturation+5.85963e-11*lvp_saturation+1.53340e-10'
+ sky130_fd_pr__pfet_01v8__b1_diff_46 = '1.30647e-10*lvp_saturation*lvp_saturation+-4.25750e-11*lvp_saturation+-1.29500e-11'
+ sky130_fd_pr__pfet_01v8__b1_diff_47 = '5.15772e-10*lvp_saturation*lvp_saturation+-3.13734e-09*lvp_saturation+2.52230e-09'
+ sky130_fd_pr__pfet_01v8__b1_diff_48 = '2.39769e-10*lvp_saturation*lvp_saturation+-3.08657e-09*lvp_saturation+3.31390e-10'
+ sky130_fd_pr__pfet_01v8__b1_diff_49 = '1.09084e-09*lvp_saturation*lvp_saturation+2.05499e-09*lvp_saturation+6.49550e-10'
+ sky130_fd_pr__pfet_01v8__dlc_diff = '-4.33125e-09*poly_cd'
+ sky130_fd_pr__pfet_01v8__dwc_diff = '8.04375e-09*diff_cd'
+ sky130_fd_pr__pfet_01v8__k2_diff_0 = '7.05787e-04*lvp_bodyeffect*lvp_bodyeffect+-3.18165e-03*lvp_bodyeffect+-1.94680e-02'
+ sky130_fd_pr__pfet_01v8__k2_diff_1 = '6.67959e-04*lvp_bodyeffect*lvp_bodyeffect+-3.15859e-03*lvp_bodyeffect+-2.32770e-02'
+ sky130_fd_pr__pfet_01v8__k2_diff_10 = '1.53956e-03*lvp_bodyeffect*lvp_bodyeffect+-8.34925e-03*lvp_bodyeffect+-1.82590e-02'
+ sky130_fd_pr__pfet_01v8__k2_diff_11 = '3.26563e-05*lvp_bodyeffect*lvp_bodyeffect+-4.03750e-05*lvp_bodyeffect+-1.52750e-02'
+ sky130_fd_pr__pfet_01v8__k2_diff_12 = '2.43156e-05*lvp_bodyeffect*lvp_bodyeffect+-4.81513e-04*lvp_bodyeffect+-1.04560e-02'
+ sky130_fd_pr__pfet_01v8__k2_diff_13 = '1.94375e-05*lvp_bodyeffect*lvp_bodyeffect+-5.02800e-04*lvp_bodyeffect+-8.56880e-03'
+ sky130_fd_pr__pfet_01v8__k2_diff_14 = '3.02156e-05*lvp_bodyeffect*lvp_bodyeffect+-3.10537e-04*lvp_bodyeffect+-8.11600e-03'
+ sky130_fd_pr__pfet_01v8__k2_diff_15 = '5.71901e-04*lvp_bodyeffect*lvp_bodyeffect+-2.67810e-03*lvp_bodyeffect+-1.90650e-02'
+ sky130_fd_pr__pfet_01v8__k2_diff_16 = '3.83431e-04*lvp_bodyeffect*lvp_bodyeffect+-3.10823e-03*lvp_bodyeffect+-1.55610e-02'
+ sky130_fd_pr__pfet_01v8__k2_diff_17 = '8.59125e-05*lvp_bodyeffect*lvp_bodyeffect+-1.98038e-03*lvp_bodyeffect+-7.32510e-03'
+ sky130_fd_pr__pfet_01v8__k2_diff_18 = '1.72500e-05*lvp_bodyeffect*lvp_bodyeffect+-6.70250e-04*lvp_bodyeffect+-1.54950e-02'
+ sky130_fd_pr__pfet_01v8__k2_diff_19 = '-3.88438e-05*lvp_bodyeffect*lvp_bodyeffect+-1.24625e-04*lvp_bodyeffect+-9.61600e-03'
+ sky130_fd_pr__pfet_01v8__k2_diff_2 = '8.15844e-05*lvp_bodyeffect*lvp_bodyeffect+-2.97962e-04*lvp_bodyeffect+-1.00760e-02'
+ sky130_fd_pr__pfet_01v8__k2_diff_20 = '1.59281e-05*lvp_bodyeffect*lvp_bodyeffect+-6.40713e-04*lvp_bodyeffect+-1.19310e-02'
+ sky130_fd_pr__pfet_01v8__k2_diff_21 = '1.81312e-05*lvp_bodyeffect*lvp_bodyeffect+-4.84525e-04*lvp_bodyeffect+-1.18870e-02'
+ sky130_fd_pr__pfet_01v8__k2_diff_22 = '2.18438e-05*lvp_bodyeffect*lvp_bodyeffect+-4.94375e-04*lvp_bodyeffect+-1.21090e-02'
+ sky130_fd_pr__pfet_01v8__k2_diff_23 = '1.68828e-03*lvp_bodyeffect*lvp_bodyeffect+-7.02262e-03*lvp_bodyeffect+-1.47580e-02'
+ sky130_fd_pr__pfet_01v8__k2_diff_24 = '3.57697e-04*lvp_bodyeffect*lvp_bodyeffect+-2.70029e-03*lvp_bodyeffect+-1.12360e-02'
+ sky130_fd_pr__pfet_01v8__k2_diff_25 = '1.03217e-04*lvp_bodyeffect*lvp_bodyeffect+-1.58204e-03*lvp_bodyeffect+-8.15730e-03'
+ sky130_fd_pr__pfet_01v8__k2_diff_26 = '1.38750e-05*lvp_bodyeffect*lvp_bodyeffect+-8.28250e-04*lvp_bodyeffect+-1.52440e-02'
+ sky130_fd_pr__pfet_01v8__k2_diff_27 = '1.81187e-05*lvp_bodyeffect*lvp_bodyeffect+-3.88475e-04*lvp_bodyeffect+-1.01500e-02'
+ sky130_fd_pr__pfet_01v8__k2_diff_28 = '1.56875e-05*lvp_bodyeffect*lvp_bodyeffect+-4.61250e-04*lvp_bodyeffect+-1.28930e-02'
+ sky130_fd_pr__pfet_01v8__k2_diff_29 = '1.43750e-05*lvp_bodyeffect*lvp_bodyeffect+-4.39000e-04*lvp_bodyeffect+-1.23670e-02'
+ sky130_fd_pr__pfet_01v8__k2_diff_3 = '3.11966e-04*lvp_bodyeffect*lvp_bodyeffect+9.17112e-04*lvp_bodyeffect+-1.35080e-02'
+ sky130_fd_pr__pfet_01v8__k2_diff_30 = '1.91562e-05*lvp_bodyeffect*lvp_bodyeffect+-5.18875e-04*lvp_bodyeffect+-1.32100e-02'
+ sky130_fd_pr__pfet_01v8__k2_diff_31 = '6.62528e-04*lvp_bodyeffect*lvp_bodyeffect+-2.47711e-03*lvp_bodyeffect+-1.71210e-02'
+ sky130_fd_pr__pfet_01v8__k2_diff_32 = '3.56166e-04*lvp_bodyeffect*lvp_bodyeffect+-2.49491e-03*lvp_bodyeffect+-1.44440e-02'
+ sky130_fd_pr__pfet_01v8__k2_diff_33 = '9.02437e-05*lvp_bodyeffect*lvp_bodyeffect+-1.54297e-03*lvp_bodyeffect+-1.08220e-02'
+ sky130_fd_pr__pfet_01v8__k2_diff_34 = '-8.58437e-05*lvp_bodyeffect*lvp_bodyeffect+-6.84625e-04*lvp_bodyeffect+-1.60000e-02'
+ sky130_fd_pr__pfet_01v8__k2_diff_35 = '4.86212e-04*lvp_bodyeffect*lvp_bodyeffect+2.42957e-03*lvp_bodyeffect+-6.68970e-03'
+ sky130_fd_pr__pfet_01v8__k2_diff_36 = '1.82681e-04*lvp_bodyeffect*lvp_bodyeffect+2.89478e-03*lvp_bodyeffect+6.48600e-03'
+ sky130_fd_pr__pfet_01v8__k2_diff_37 = '-1.23409e-04*lvp_bodyeffect*lvp_bodyeffect+2.01944e-03*lvp_bodyeffect+3.16150e-03'
+ sky130_fd_pr__pfet_01v8__k2_diff_38 = '-1.49109e-04*lvp_bodyeffect*lvp_bodyeffect+2.07381e-03*lvp_bodyeffect+-1.69800e-03'
+ sky130_fd_pr__pfet_01v8__k2_diff_39 = '1.54059e-04*lvp_bodyeffect*lvp_bodyeffect+-1.31559e-03*lvp_bodyeffect+1.66750e-03'
+ sky130_fd_pr__pfet_01v8__k2_diff_4 = '1.91416e-04*lvp_bodyeffect*lvp_bodyeffect+5.44663e-04*lvp_bodyeffect+-1.41490e-02'
+ sky130_fd_pr__pfet_01v8__k2_diff_40 = '7.42069e-04*lvp_bodyeffect*lvp_bodyeffect+-2.86202e-03*lvp_bodyeffect+-3.01160e-02'
+ sky130_fd_pr__pfet_01v8__k2_diff_41 = '8.42053e-04*lvp_bodyeffect*lvp_bodyeffect+3.88621e-03*lvp_bodyeffect+-2.31780e-02'
+ sky130_fd_pr__pfet_01v8__k2_diff_42 = '6.75963e-04*lvp_bodyeffect*lvp_bodyeffect+2.84285e-03*lvp_bodyeffect+-6.54280e-03'
+ sky130_fd_pr__pfet_01v8__k2_diff_43 = '6.59938e-04*lvp_bodyeffect*lvp_bodyeffect+3.68475e-03*lvp_bodyeffect+-1.13200e-02'
+ sky130_fd_pr__pfet_01v8__k2_diff_44 = '1.70816e-04*lvp_bodyeffect*lvp_bodyeffect+8.59162e-04*lvp_bodyeffect+-8.36270e-03'
+ sky130_fd_pr__pfet_01v8__k2_diff_45 = '5.24504e-04*lvp_bodyeffect*lvp_bodyeffect+-3.17550e-04*lvp_bodyeffect+7.87730e-04'
+ sky130_fd_pr__pfet_01v8__k2_diff_46 = '4.67903e-04*lvp_bodyeffect*lvp_bodyeffect+2.37036e-03*lvp_bodyeffect+-1.13710e-02'
+ sky130_fd_pr__pfet_01v8__k2_diff_47 = '1.52205e-03*lvp_bodyeffect*lvp_bodyeffect+-2.37570e-03*lvp_bodyeffect+-2.48650e-02'
+ sky130_fd_pr__pfet_01v8__k2_diff_48 = '1.36559e-03*lvp_bodyeffect*lvp_bodyeffect+4.82488e-03*lvp_bodyeffect+-1.88860e-02'
+ sky130_fd_pr__pfet_01v8__k2_diff_49 = '5.92188e-04*lvp_bodyeffect*lvp_bodyeffect+-4.47850e-03*lvp_bodyeffect+-1.31150e-02'
+ sky130_fd_pr__pfet_01v8__k2_diff_5 = '4.09531e-04*lvp_bodyeffect*lvp_bodyeffect+1.58388e-03*lvp_bodyeffect+-1.52900e-02'
+ sky130_fd_pr__pfet_01v8__k2_diff_50 = '4.37750e-04*lvp_bodyeffect*lvp_bodyeffect+-2.14875e-03*lvp_bodyeffect+-4.02950e-02'
+ sky130_fd_pr__pfet_01v8__k2_diff_51 = '6.78900e-04*lvp_bodyeffect*lvp_bodyeffect+-3.83635e-03*lvp_bodyeffect+-3.07030e-02'
+ sky130_fd_pr__pfet_01v8__k2_diff_6 = '1.46225e-03*lvp_bodyeffect*lvp_bodyeffect+-6.89475e-03*lvp_bodyeffect+-2.58480e-02'
+ sky130_fd_pr__pfet_01v8__k2_diff_7 = '6.12393e-04*lvp_bodyeffect*lvp_bodyeffect+-1.98232e-03*lvp_bodyeffect+-1.84930e-02'
+ sky130_fd_pr__pfet_01v8__k2_diff_8 = '1.11597e-04*lvp_bodyeffect*lvp_bodyeffect+-1.31224e-03*lvp_bodyeffect+-9.23160e-03'
+ sky130_fd_pr__pfet_01v8__k2_diff_9 = '4.79875e-05*lvp_bodyeffect*lvp_bodyeffect+-2.82700e-04*lvp_bodyeffect+-1.06500e-02'
+ sky130_fd_pr__pfet_01v8__lint_diff = '-4.33125e-09*poly_cd'
+ sky130_fd_pr__pfet_01v8__nfactor_diff_0 = '3.84303e-02*lvp_subvt*lvp_subvt+-3.57384e-01*lvp_subvt+6.60780e-01'
+ sky130_fd_pr__pfet_01v8__nfactor_diff_1 = '2.73244e-02*lvp_subvt*lvp_subvt+-3.60525e-01*lvp_subvt+7.98710e-01'
+ sky130_fd_pr__pfet_01v8__nfactor_diff_10 = '-2.73984e-02*lvp_subvt*lvp_subvt+-1.90661e-01*lvp_subvt+8.83130e-01'
+ sky130_fd_pr__pfet_01v8__nfactor_diff_11 = '7.69385e-03*lvp_subvt*lvp_subvt+-2.64316e-02*lvp_subvt+-2.51980e-02'
+ sky130_fd_pr__pfet_01v8__nfactor_diff_12 = '5.15490e-03*lvp_subvt*lvp_subvt+-2.31182e-02*lvp_subvt+1.13690e-02'
+ sky130_fd_pr__pfet_01v8__nfactor_diff_13 = '3.09959e-03*lvp_subvt*lvp_subvt+-2.10771e-02*lvp_subvt+4.65280e-02'
+ sky130_fd_pr__pfet_01v8__nfactor_diff_14 = '3.91160e-03*lvp_subvt*lvp_subvt+-2.60876e-02*lvp_subvt+3.87940e-02'
+ sky130_fd_pr__pfet_01v8__nfactor_diff_15 = '1.76816e-02*lvp_subvt*lvp_subvt+-3.66229e-01*lvp_subvt+8.44480e-01'
+ sky130_fd_pr__pfet_01v8__nfactor_diff_16 = '2.63777e-02*lvp_subvt*lvp_subvt+-1.89422e-01*lvp_subvt+3.30970e-01'
+ sky130_fd_pr__pfet_01v8__nfactor_diff_17 = '3.13750e-02*lvp_subvt*lvp_subvt+-9.87356e-02*lvp_subvt+-5.70730e-02'
+ sky130_fd_pr__pfet_01v8__nfactor_diff_18 = '1.15203e-02*lvp_subvt*lvp_subvt+-4.99837e-02*lvp_subvt+1.34850e-01'
+ sky130_fd_pr__pfet_01v8__nfactor_diff_19 = '1.34827e-03*lvp_subvt*lvp_subvt+6.08759e-03*lvp_subvt+-3.90410e-02'
+ sky130_fd_pr__pfet_01v8__nfactor_diff_2 = '1.12942e-02*lvp_subvt*lvp_subvt+-1.25319e-02*lvp_subvt+-7.99440e-02'
+ sky130_fd_pr__pfet_01v8__nfactor_diff_20 = '3.08258e-03*lvp_subvt*lvp_subvt+-2.37317e-02*lvp_subvt+4.81120e-02'
+ sky130_fd_pr__pfet_01v8__nfactor_diff_21 = '2.06494e-03*lvp_subvt*lvp_subvt+-1.49210e-02*lvp_subvt+5.66070e-02'
+ sky130_fd_pr__pfet_01v8__nfactor_diff_22 = '3.48603e-03*lvp_subvt*lvp_subvt+-2.43421e-02*lvp_subvt+6.08450e-02'
+ sky130_fd_pr__pfet_01v8__nfactor_diff_23 = '6.84062e-04*lvp_subvt*lvp_subvt+-1.81874e-01*lvp_subvt+5.92860e-01'
+ sky130_fd_pr__pfet_01v8__nfactor_diff_24 = '2.99061e-02*lvp_subvt*lvp_subvt+-1.97116e-01*lvp_subvt+2.84140e-01'
+ sky130_fd_pr__pfet_01v8__nfactor_diff_25 = '1.43391e-02*lvp_subvt*lvp_subvt+-5.52662e-02*lvp_subvt+1.10820e-01'
+ sky130_fd_pr__pfet_01v8__nfactor_diff_26 = '4.93313e-03*lvp_subvt*lvp_subvt+-3.41275e-02*lvp_subvt+1.75260e-01'
+ sky130_fd_pr__pfet_01v8__nfactor_diff_27 = '4.86519e-03*lvp_subvt*lvp_subvt+-9.81925e-03*lvp_subvt+-7.78750e-02'
+ sky130_fd_pr__pfet_01v8__nfactor_diff_28 = '2.74741e-03*lvp_subvt*lvp_subvt+-1.51735e-02*lvp_subvt+3.76740e-03'
+ sky130_fd_pr__pfet_01v8__nfactor_diff_29 = '2.92334e-03*lvp_subvt*lvp_subvt+-1.96666e-02*lvp_subvt+6.06700e-02'
+ sky130_fd_pr__pfet_01v8__nfactor_diff_3 = '1.41390e-03*lvp_subvt*lvp_subvt+-2.20167e-02*lvp_subvt+7.40910e-02'
+ sky130_fd_pr__pfet_01v8__nfactor_diff_30 = '4.43869e-03*lvp_subvt*lvp_subvt+-3.01965e-02*lvp_subvt+9.34650e-02'
+ sky130_fd_pr__pfet_01v8__nfactor_diff_31 = '1.46009e-02*lvp_subvt*lvp_subvt+-2.28531e-01*lvp_subvt+5.70960e-01'
+ sky130_fd_pr__pfet_01v8__nfactor_diff_32 = '1.37156e-02*lvp_subvt*lvp_subvt+-1.36392e-01*lvp_subvt+2.11590e-01'
+ sky130_fd_pr__pfet_01v8__nfactor_diff_33 = '1.60181e-02*lvp_subvt*lvp_subvt+9.41750e-03*lvp_subvt+1.04370e-01'
+ sky130_fd_pr__pfet_01v8__nfactor_diff_34 = '-2.31187e-03*lvp_subvt*lvp_subvt+-1.24500e-03*lvp_subvt+2.79190e-01'
+ sky130_fd_pr__pfet_01v8__nfactor_diff_35 = '1.09280e-02*lvp_subvt*lvp_subvt+-1.24823e-01*lvp_subvt+2.34410e-01'
+ sky130_fd_pr__pfet_01v8__nfactor_diff_36 = '1.20758e-02*lvp_subvt*lvp_subvt+-9.32187e-02*lvp_subvt+2.92220e-02'
+ sky130_fd_pr__pfet_01v8__nfactor_diff_37 = '8.82813e-03*lvp_subvt*lvp_subvt+-5.76705e-02*lvp_subvt+5.12680e-02'
+ sky130_fd_pr__pfet_01v8__nfactor_diff_38 = '9.08134e-03*lvp_subvt*lvp_subvt+-6.97446e-02*lvp_subvt+4.43100e-02'
+ sky130_fd_pr__pfet_01v8__nfactor_diff_39 = '3.71031e-04*lvp_subvt*lvp_subvt+-4.14913e-03*lvp_subvt+1.06600e-02'
+ sky130_fd_pr__pfet_01v8__nfactor_diff_4 = '2.31746e-02*lvp_subvt*lvp_subvt+6.33700e-02*lvp_subvt+6.52360e-02'
+ sky130_fd_pr__pfet_01v8__nfactor_diff_40 = '1.82406e-02*lvp_subvt*lvp_subvt+-6.49987e-01*lvp_subvt+1.10810e+00'
+ sky130_fd_pr__pfet_01v8__nfactor_diff_41 = '8.59884e-02*lvp_subvt*lvp_subvt+-6.66546e-01*lvp_subvt+1.14840e+00'
+ sky130_fd_pr__pfet_01v8__nfactor_diff_42 = '5.63731e-02*lvp_subvt*lvp_subvt+1.43300e-02*lvp_subvt+1.41810e-01'
+ sky130_fd_pr__pfet_01v8__nfactor_diff_43 = '1.47086e-01*lvp_subvt*lvp_subvt+-2.13438e-01*lvp_subvt+1.40770e-01'
+ sky130_fd_pr__pfet_01v8__nfactor_diff_44 = '1.85312e-02*lvp_subvt*lvp_subvt+2.00625e-02*lvp_subvt+1.00720e-01'
+ sky130_fd_pr__pfet_01v8__nfactor_diff_45 = '-9.06087e-03*lvp_subvt*lvp_subvt+2.54895e-02*lvp_subvt+2.93620e-02'
+ sky130_fd_pr__pfet_01v8__nfactor_diff_46 = '4.69084e-03*lvp_subvt*lvp_subvt+-8.52991e-02*lvp_subvt+1.83700e-01'
+ sky130_fd_pr__pfet_01v8__nfactor_diff_47 = '5.56556e-02*lvp_subvt*lvp_subvt+-5.21253e-01*lvp_subvt+1.00260e+00'
+ sky130_fd_pr__pfet_01v8__nfactor_diff_48 = '1.04121e-02*lvp_subvt*lvp_subvt+-5.31566e-02*lvp_subvt+1.03760e-01'
+ sky130_fd_pr__pfet_01v8__nfactor_diff_49 = '8.31250e-04*lvp_subvt*lvp_subvt+-7.25000e-01*lvp_subvt+1.08670e+00'
+ sky130_fd_pr__pfet_01v8__nfactor_diff_5 = '3.61128e-03*lvp_subvt*lvp_subvt+-3.88401e-02*lvp_subvt+8.67190e-02'
+ sky130_fd_pr__pfet_01v8__nfactor_diff_50 = '1.26725e-02*lvp_subvt*lvp_subvt+-5.88025e-01*lvp_subvt+9.49340e-01'
+ sky130_fd_pr__pfet_01v8__nfactor_diff_51 = '4.52959e-02*lvp_subvt*lvp_subvt+-4.05256e-01*lvp_subvt+5.24740e-01'
+ sky130_fd_pr__pfet_01v8__nfactor_diff_6 = '3.14344e-03*lvp_subvt*lvp_subvt+-3.20794e-01*lvp_subvt+8.42530e-01'
+ sky130_fd_pr__pfet_01v8__nfactor_diff_7 = '-1.39813e-03*lvp_subvt*lvp_subvt+-3.98800e-01*lvp_subvt+4.17570e-01'
+ sky130_fd_pr__pfet_01v8__nfactor_diff_8 = '3.48203e-02*lvp_subvt*lvp_subvt+-1.48192e-01*lvp_subvt+-2.74920e-02'
+ sky130_fd_pr__pfet_01v8__nfactor_diff_9 = '8.81575e-03*lvp_subvt*lvp_subvt+-3.46595e-02*lvp_subvt+-1.54010e-03'
+ sky130_fd_pr__pfet_01v8__overlap_mult = '7.47062e-03*lvtox*lvtox+2.98800e-02*lvtox+9.54350e-01'
+ sky130_fd_pr__pfet_01v8__pjunction_mult = '2.18750e-06*lvp_diode*lvp_diode+2.37662e-02*lvp_diode+1.00090e+00'
+ sky130_fd_pr__rf_pfet_01v8__aw_cap_mult = '3.75000e-02*pfet_01v8+1.00000e+00'
+ sky130_fd_pr__rf_pfet_01v8__aw_cap_mult_2 = '3.75000e-02*pfet_01v8+1.00000e+00'
+ sky130_fd_pr__rf_pfet_01v8__aw_rgate_dist_mult = '6.87500e-03*pfet_01v8*pfet_01v8+8.50000e-02*pfet_01v8+1.00000e+00'
+ sky130_fd_pr__rf_pfet_01v8__aw_rgate_dist_mult_2 = '3.12500e-03*pfet_01v8*pfet_01v8+6.25000e-02*pfet_01v8+1.00000e+00'
+ sky130_fd_pr__rf_pfet_01v8__aw_rgate_stub_mult = '6.87500e-03*lvp_mobility*lvp_mobility+8.50000e-02*lvp_mobility+1.00000e+00'
+ sky130_fd_pr__rf_pfet_01v8__aw_rgate_stub_mult_2 = '3.12500e-03*lvp_mobility*lvp_mobility+6.25000e-02*lvp_mobility+1.00000e+00'
+ sky130_fd_pr__rf_pfet_01v8_b__ajunction_mult = '-3.12500e-07*lvp_diode*lvp_diode+2.36612e-02*lvp_diode+9.96260e-01'
+ sky130_fd_pr__rf_pfet_01v8_b__dlc_diff = '-4.33125e-09*poly_cd'
+ sky130_fd_pr__rf_pfet_01v8_b__lint_diff = '-4.33125e-09*poly_cd'
+ sky130_fd_pr__rf_pfet_01v8_b__overlap_mult = '7.47062e-03*lvtox*lvtox+2.98800e-02*lvtox+9.54350e-01'
+ sky130_fd_pr__rf_pfet_01v8_b__pjunction_mult = '2.18750e-06*lvp_diode*lvp_diode+2.37662e-02*lvp_diode+1.00090e+00'
+ sky130_fd_pr__rf_pfet_01v8_b__rbpb_mult = '5.00000e-02*lvp_bodyeffect+1.00000e+00'
+ sky130_fd_pr__rf_pfet_01v8_b__rshg_diff = '1.75000e+00*ic_res'
+ sky130_fd_pr__rf_pfet_01v8_b__toxe_mult = '1.30000e-02*lvtox+1.00000e+00'
+ sky130_fd_pr__rf_pfet_01v8_b__wint_diff = '8.04375e-09*diff_cd'
+ sky130_fd_pr__rf_pfet_01v8_b__xgw_diff = '1.60625e-08*diff_cd'
+ sky130_fd_pr__rf_pfet_01v8_bM02__k2_diff_0 = '7.88925e-04*lvp_bodyeffect*lvp_bodyeffect+-3.74695e-03*lvp_bodyeffect+-2.39530e-02'
+ sky130_fd_pr__rf_pfet_01v8_bM02__k2_diff_1 = '4.12838e-04*lvp_bodyeffect*lvp_bodyeffect+-7.85000e-05*lvp_bodyeffect+-1.46000e-02'
+ sky130_fd_pr__rf_pfet_01v8_bM02__k2_diff_2 = '8.07491e-05*lvp_bodyeffect*lvp_bodyeffect+4.28325e-03*lvp_bodyeffect+-1.75040e-02'
+ sky130_fd_pr__rf_pfet_01v8_bM02__k2_diff_3 = '8.30297e-04*lvp_bodyeffect*lvp_bodyeffect+-2.77369e-03*lvp_bodyeffect+-2.56720e-02'
+ sky130_fd_pr__rf_pfet_01v8_bM02__k2_diff_4 = '4.43511e-04*lvp_bodyeffect*lvp_bodyeffect+-2.39504e-03*lvp_bodyeffect+-1.64290e-02'
+ sky130_fd_pr__rf_pfet_01v8_bM02__k2_diff_5 = '1.27375e-04*lvp_bodyeffect*lvp_bodyeffect+1.05000e-05*lvp_bodyeffect+-1.85780e-02'
+ sky130_fd_pr__rf_pfet_01v8_bM02__k2_diff_6 = '8.48497e-04*lvp_bodyeffect*lvp_bodyeffect+-2.83474e-03*lvp_bodyeffect+-2.63870e-02'
+ sky130_fd_pr__rf_pfet_01v8_bM02__k2_diff_7 = '4.38997e-04*lvp_bodyeffect*lvp_bodyeffect+-1.75149e-03*lvp_bodyeffect+-1.36950e-02'
+ sky130_fd_pr__rf_pfet_01v8_bM02__k2_diff_8 = '1.16562e-04*lvp_bodyeffect*lvp_bodyeffect+8.99500e-04*lvp_bodyeffect+-1.78310e-02'
+ sky130_fd_pr__rf_pfet_01v8_bM02__u0_diff_0 = '-2.95281e-06*lvp_mobility*lvp_mobility+1.07038e-05*lvp_mobility+-2.56080e-04'
+ sky130_fd_pr__rf_pfet_01v8_bM02__u0_diff_1 = '-3.17469e-06*lvp_mobility*lvp_mobility+-7.32625e-06*lvp_mobility+-1.75340e-04'
+ sky130_fd_pr__rf_pfet_01v8_bM02__u0_diff_2 = '-5.07816e-06*lvp_mobility*lvp_mobility+-4.14349e-05*lvp_mobility+-1.15280e-04'
+ sky130_fd_pr__rf_pfet_01v8_bM02__u0_diff_3 = '-1.61219e-06*lvp_mobility*lvp_mobility+-4.63037e-05*lvp_mobility+-4.39530e-04'
+ sky130_fd_pr__rf_pfet_01v8_bM02__u0_diff_4 = '-2.81625e-06*lvp_mobility*lvp_mobility+-8.32000e-06*lvp_mobility+-4.02980e-04'
+ sky130_fd_pr__rf_pfet_01v8_bM02__u0_diff_5 = '-3.43469e-06*lvp_mobility*lvp_mobility+-2.94162e-05*lvp_mobility+-2.29660e-04'
+ sky130_fd_pr__rf_pfet_01v8_bM02__u0_diff_6 = '-1.04187e-06*lvp_mobility*lvp_mobility+-6.76675e-05*lvp_mobility+-7.89060e-04'
+ sky130_fd_pr__rf_pfet_01v8_bM02__u0_diff_7 = '-3.19031e-06*lvp_mobility*lvp_mobility+-2.56063e-05*lvp_mobility+-3.06110e-04'
+ sky130_fd_pr__rf_pfet_01v8_bM02__u0_diff_8 = '-2.76312e-06*lvp_mobility*lvp_mobility+-4.04825e-05*lvp_mobility+-3.26940e-04'
+ sky130_fd_pr__rf_pfet_01v8_bM02__vsat_diff_0 = '-2.19959e+02*lvp_saturation*lvp_saturation+3.58099e+03*lvp_saturation+-1.79270e+03'
+ sky130_fd_pr__rf_pfet_01v8_bM02__vsat_diff_1 = '-6.67469e+02*lvp_saturation*lvp_saturation+2.31875e+02*lvp_saturation+-3.93900e+03'
+ sky130_fd_pr__rf_pfet_01v8_bM02__vsat_diff_2 = '-3.74053e+02*lvp_saturation*lvp_saturation+-8.13988e+02*lvp_saturation+-3.70520e+03'
+ sky130_fd_pr__rf_pfet_01v8_bM02__vsat_diff_3 = '-4.49481e+02*lvp_saturation*lvp_saturation+9.72500e+02*lvp_saturation+-7.60430e+03'
+ sky130_fd_pr__rf_pfet_01v8_bM02__vsat_diff_4 = '-5.17684e+02*lvp_saturation*lvp_saturation+8.18238e+02*lvp_saturation+2.22900e+02'
+ sky130_fd_pr__rf_pfet_01v8_bM02__vsat_diff_5 = '-1.04765e+03*lvp_saturation*lvp_saturation+-8.24300e+02*lvp_saturation+1.23580e+04'
+ sky130_fd_pr__rf_pfet_01v8_bM02__vsat_diff_6 = '-5.68250e+02*lvp_saturation*lvp_saturation+8.48900e+02*lvp_saturation+-3.99640e+03'
+ sky130_fd_pr__rf_pfet_01v8_bM02__vsat_diff_7 = '-6.26394e+02*lvp_saturation*lvp_saturation+6.40750e+02*lvp_saturation+-5.40770e+03'
+ sky130_fd_pr__rf_pfet_01v8_bM02__vsat_diff_8 = '-8.45866e+02*lvp_saturation*lvp_saturation+-1.39554e+03*lvp_saturation+2.23200e+03'
+ sky130_fd_pr__rf_pfet_01v8_bM02__vth0_diff_0 = '-2.08957e-03*lvp_threshold*lvp_threshold+1.60973e-02*lvp_threshold+5.41510e-03'
+ sky130_fd_pr__rf_pfet_01v8_bM02__vth0_diff_1 = '-1.03035e-03*lvp_threshold*lvp_threshold+1.53896e-02*lvp_threshold+-1.32890e-03'
+ sky130_fd_pr__rf_pfet_01v8_bM02__vth0_diff_2 = '-2.39119e-04*lvp_threshold*lvp_threshold+6.98988e-03*lvp_threshold+1.68740e-03'
+ sky130_fd_pr__rf_pfet_01v8_bM02__vth0_diff_3 = '-2.17209e-03*lvp_threshold*lvp_threshold+2.30241e-02*lvp_threshold+5.54000e-03'
+ sky130_fd_pr__rf_pfet_01v8_bM02__vth0_diff_4 = '-1.09537e-03*lvp_threshold*lvp_threshold+1.57754e-02*lvp_threshold+9.01640e-03'
+ sky130_fd_pr__rf_pfet_01v8_bM02__vth0_diff_5 = '-2.77719e-04*lvp_threshold*lvp_threshold+6.42650e-03*lvp_threshold+4.31850e-03'
+ sky130_fd_pr__rf_pfet_01v8_bM02__vth0_diff_6 = '-2.17009e-03*lvp_threshold*lvp_threshold+2.74224e-02*lvp_threshold+1.32910e-02'
+ sky130_fd_pr__rf_pfet_01v8_bM02__vth0_diff_7 = '-1.05824e-03*lvp_threshold*lvp_threshold+1.65510e-02*lvp_threshold+5.46190e-03'
+ sky130_fd_pr__rf_pfet_01v8_bM02__vth0_diff_8 = '-2.81481e-04*lvp_threshold*lvp_threshold+8.40712e-03*lvp_threshold+3.05520e-03'
+ sky130_fd_pr__rf_pfet_01v8_bM04__k2_diff_0 = '8.11859e-04*lvp_bodyeffect*lvp_bodyeffect+-3.96794e-03*lvp_bodyeffect+-2.22710e-02'
+ sky130_fd_pr__rf_pfet_01v8_bM04__k2_diff_1 = '4.22813e-04*lvp_bodyeffect*lvp_bodyeffect+-2.25700e-04*lvp_bodyeffect+-1.40490e-02'
+ sky130_fd_pr__rf_pfet_01v8_bM04__k2_diff_2 = '7.11859e-05*lvp_bodyeffect*lvp_bodyeffect+4.23974e-03*lvp_bodyeffect+-1.85950e-02'
+ sky130_fd_pr__rf_pfet_01v8_bM04__k2_diff_3 = '8.25749e-04*lvp_bodyeffect*lvp_bodyeffect+-2.75950e-03*lvp_bodyeffect+-2.34610e-02'
+ sky130_fd_pr__rf_pfet_01v8_bM04__k2_diff_4 = '4.42350e-04*lvp_bodyeffect*lvp_bodyeffect+-2.42190e-03*lvp_bodyeffect+-1.27890e-02'
+ sky130_fd_pr__rf_pfet_01v8_bM04__k2_diff_5 = '1.26969e-04*lvp_bodyeffect*lvp_bodyeffect+-2.36250e-05*lvp_bodyeffect+-1.85990e-02'
+ sky130_fd_pr__rf_pfet_01v8_bM04__k2_diff_6 = '8.47931e-04*lvp_bodyeffect*lvp_bodyeffect+-2.95897e-03*lvp_bodyeffect+-2.51000e-02'
+ sky130_fd_pr__rf_pfet_01v8_bM04__k2_diff_7 = '4.38387e-04*lvp_bodyeffect*lvp_bodyeffect+-1.69255e-03*lvp_bodyeffect+-1.09530e-02'
+ sky130_fd_pr__rf_pfet_01v8_bM04__k2_diff_8 = '1.15937e-04*lvp_bodyeffect*lvp_bodyeffect+8.62750e-04*lvp_bodyeffect+-1.66060e-02'
+ sky130_fd_pr__rf_pfet_01v8_bM04__u0_diff_0 = '-3.02500e-06*lvp_mobility*lvp_mobility+6.14500e-06*lvp_mobility+-4.34040e-04'
+ sky130_fd_pr__rf_pfet_01v8_bM04__u0_diff_1 = '-3.78563e-06*lvp_mobility*lvp_mobility+-1.01825e-05*lvp_mobility+-2.53300e-04'
+ sky130_fd_pr__rf_pfet_01v8_bM04__u0_diff_2 = '-3.14672e-06*lvp_mobility*lvp_mobility+-4.08281e-05*lvp_mobility+-1.85700e-04'
+ sky130_fd_pr__rf_pfet_01v8_bM04__u0_diff_3 = '-5.81562e-07*lvp_mobility*lvp_mobility+-4.06338e-05*lvp_mobility+-5.35030e-04'
+ sky130_fd_pr__rf_pfet_01v8_bM04__u0_diff_4 = '-2.25750e-06*lvp_mobility*lvp_mobility+-1.96525e-05*lvp_mobility+-6.24650e-04'
+ sky130_fd_pr__rf_pfet_01v8_bM04__u0_diff_5 = '-3.40312e-06*lvp_mobility*lvp_mobility+-3.32025e-05*lvp_mobility+-3.34450e-04'
+ sky130_fd_pr__rf_pfet_01v8_bM04__u0_diff_6 = '-7.05625e-07*lvp_mobility*lvp_mobility+-7.59700e-05*lvp_mobility+-6.46020e-04'
+ sky130_fd_pr__rf_pfet_01v8_bM04__u0_diff_7 = '-3.02000e-06*lvp_mobility*lvp_mobility+-2.82000e-05*lvp_mobility+-5.75480e-04'
+ sky130_fd_pr__rf_pfet_01v8_bM04__u0_diff_8 = '-2.91781e-06*lvp_mobility*lvp_mobility+-4.52087e-05*lvp_mobility+-4.40410e-04'
+ sky130_fd_pr__rf_pfet_01v8_bM04__vsat_diff_0 = '-3.93106e+02*lvp_saturation*lvp_saturation+3.06255e+03*lvp_saturation+-1.65610e+03'
+ sky130_fd_pr__rf_pfet_01v8_bM04__vsat_diff_1 = '-4.90413e+02*lvp_saturation*lvp_saturation+1.33069e+03*lvp_saturation+8.76350e+02'
+ sky130_fd_pr__rf_pfet_01v8_bM04__vsat_diff_2 = '-1.32498e+03*lvp_saturation*lvp_saturation+-1.38783e+03*lvp_saturation+1.59210e+04'
+ sky130_fd_pr__rf_pfet_01v8_bM04__vsat_diff_3 = '-6.36825e+02*lvp_saturation*lvp_saturation+7.42250e+02*lvp_saturation+-2.98080e+03'
+ sky130_fd_pr__rf_pfet_01v8_bM04__vsat_diff_4 = '-6.15031e+02*lvp_saturation*lvp_saturation+1.22375e+02*lvp_saturation+-1.15500e+03'
+ sky130_fd_pr__rf_pfet_01v8_bM04__vsat_diff_5 = '-1.24004e+03*lvp_saturation*lvp_saturation+-8.54950e+02*lvp_saturation+9.11750e+03'
+ sky130_fd_pr__rf_pfet_01v8_bM04__vsat_diff_6 = '-5.66359e+02*lvp_saturation*lvp_saturation+1.15776e+03*lvp_saturation+-2.85020e+03'
+ sky130_fd_pr__rf_pfet_01v8_bM04__vsat_diff_7 = '-6.28938e+02*lvp_saturation*lvp_saturation+3.11750e+02*lvp_saturation+-3.91400e+03'
+ sky130_fd_pr__rf_pfet_01v8_bM04__vsat_diff_8 = '-1.01133e+03*lvp_saturation*lvp_saturation+-2.22694e+03*lvp_saturation+1.14100e+04'
+ sky130_fd_pr__rf_pfet_01v8_bM04__vth0_diff_0 = '-2.10059e-03*lvp_threshold*lvp_threshold+1.63614e-02*lvp_threshold+1.80470e-02'
+ sky130_fd_pr__rf_pfet_01v8_bM04__vth0_diff_1 = '-1.01603e-03*lvp_threshold*lvp_threshold+1.54661e-02*lvp_threshold+1.24260e-02'
+ sky130_fd_pr__rf_pfet_01v8_bM04__vth0_diff_2 = '-2.85394e-04*lvp_threshold*lvp_threshold+6.92225e-03*lvp_threshold+9.47730e-03'
+ sky130_fd_pr__rf_pfet_01v8_bM04__vth0_diff_3 = '-2.19548e-03*lvp_threshold*lvp_threshold+2.26099e-02*lvp_threshold+6.48720e-03'
+ sky130_fd_pr__rf_pfet_01v8_bM04__vth0_diff_4 = '-1.11394e-03*lvp_threshold*lvp_threshold+1.57338e-02*lvp_threshold+2.23420e-02'
+ sky130_fd_pr__rf_pfet_01v8_bM04__vth0_diff_5 = '-2.83188e-04*lvp_threshold*lvp_threshold+6.39900e-03*lvp_threshold+1.20970e-02'
+ sky130_fd_pr__rf_pfet_01v8_bM04__vth0_diff_6 = '-2.17306e-03*lvp_threshold*lvp_threshold+2.71660e-02*lvp_threshold+1.77530e-02'
+ sky130_fd_pr__rf_pfet_01v8_bM04__vth0_diff_7 = '-1.05896e-03*lvp_threshold*lvp_threshold+1.65740e-02*lvp_threshold+9.71640e-03'
+ sky130_fd_pr__rf_pfet_01v8_bM04__vth0_diff_8 = '-2.80031e-04*lvp_threshold*lvp_threshold+8.37688e-03*lvp_threshold+1.54910e-02'
+ sky130_fd_pr__pfet_01v8__toxe_mult = '1.30000e-02*lvtox+1.00000e+00'
+ sky130_fd_pr__pfet_01v8__u0_diff_0 = '-1.77547e-06*lvp_mobility*lvp_mobility+-7.12994e-05*lvp_mobility+3.89970e-04'
+ sky130_fd_pr__pfet_01v8__u0_diff_1 = '1.51812e-06*lvp_mobility*lvp_mobility+5.09500e-06*lvp_mobility+3.45790e-04'
+ sky130_fd_pr__pfet_01v8__u0_diff_10 = '-1.95455e-05*lvp_mobility*lvp_mobility+1.70299e-04*lvp_mobility+4.29110e-04'
+ sky130_fd_pr__pfet_01v8__u0_diff_11 = '-4.77000e-06*lvp_mobility*lvp_mobility+-1.25705e-04*lvp_mobility+1.39280e-03'
+ sky130_fd_pr__pfet_01v8__u0_diff_12 = '-3.81875e-06*lvp_mobility*lvp_mobility+-1.68125e-04*lvp_mobility+1.81130e-03'
+ sky130_fd_pr__pfet_01v8__u0_diff_13 = '-4.82344e-06*lvp_mobility*lvp_mobility+-2.11894e-04*lvp_mobility+1.79860e-03'
+ sky130_fd_pr__pfet_01v8__u0_diff_14 = '-9.49187e-06*lvp_mobility*lvp_mobility+-3.15118e-04*lvp_mobility+1.95090e-03'
+ sky130_fd_pr__pfet_01v8__u0_diff_15 = '2.67088e-05*lvp_mobility*lvp_mobility+-5.86375e-05*lvp_mobility+4.47610e-04'
+ sky130_fd_pr__pfet_01v8__u0_diff_16 = '-8.12500e-07*lvp_mobility*lvp_mobility+2.79800e-05*lvp_mobility+5.52440e-04'
+ sky130_fd_pr__pfet_01v8__u0_diff_17 = '8.39625e-06*lvp_mobility*lvp_mobility+1.62425e-05*lvp_mobility+2.05890e-04'
+ sky130_fd_pr__pfet_01v8__u0_diff_18 = '-2.67313e-06*lvp_mobility*lvp_mobility+-1.22902e-04*lvp_mobility+9.34260e-04'
+ sky130_fd_pr__pfet_01v8__u0_diff_19 = '3.27875e-06*lvp_mobility*lvp_mobility+-7.87600e-05*lvp_mobility+1.09650e-03'
+ sky130_fd_pr__pfet_01v8__u0_diff_2 = '-1.03053e-05*lvp_mobility*lvp_mobility+-2.71646e-04*lvp_mobility+1.42180e-03'
+ sky130_fd_pr__pfet_01v8__u0_diff_20 = '-1.56750e-06*lvp_mobility*lvp_mobility+-1.04745e-04*lvp_mobility+1.25940e-03'
+ sky130_fd_pr__pfet_01v8__u0_diff_21 = '-4.92656e-06*lvp_mobility*lvp_mobility+-1.75956e-04*lvp_mobility+1.62980e-03'
+ sky130_fd_pr__pfet_01v8__u0_diff_22 = '-4.80969e-06*lvp_mobility*lvp_mobility+-1.88214e-04*lvp_mobility+1.79410e-03'
+ sky130_fd_pr__pfet_01v8__u0_diff_23 = '-2.95686e-05*lvp_mobility*lvp_mobility+1.48595e-04*lvp_mobility+4.40060e-04'
+ sky130_fd_pr__pfet_01v8__u0_diff_24 = '1.86856e-06*lvp_mobility*lvp_mobility+6.39183e-05*lvp_mobility+3.24490e-04'
+ sky130_fd_pr__pfet_01v8__u0_diff_25 = '1.87688e-06*lvp_mobility*lvp_mobility+5.03650e-05*lvp_mobility+6.08760e-04'
+ sky130_fd_pr__pfet_01v8__u0_diff_26 = '4.52187e-07*lvp_mobility*lvp_mobility+-6.82413e-05*lvp_mobility+1.24720e-03'
+ sky130_fd_pr__pfet_01v8__u0_diff_27 = '-1.11781e-06*lvp_mobility*lvp_mobility+-1.29171e-04*lvp_mobility+1.21780e-03'
+ sky130_fd_pr__pfet_01v8__u0_diff_28 = '-2.11656e-06*lvp_mobility*lvp_mobility+-1.11366e-04*lvp_mobility+1.41190e-03'
+ sky130_fd_pr__pfet_01v8__u0_diff_29 = '-4.56563e-06*lvp_mobility*lvp_mobility+-1.75762e-04*lvp_mobility+1.88770e-03'
+ sky130_fd_pr__pfet_01v8__u0_diff_3 = '-1.60131e-05*lvp_mobility*lvp_mobility+-3.85027e-04*lvp_mobility+1.57820e-03'
+ sky130_fd_pr__pfet_01v8__u0_diff_30 = '-3.24687e-06*lvp_mobility*lvp_mobility+-1.62337e-04*lvp_mobility+2.03670e-03'
+ sky130_fd_pr__pfet_01v8__u0_diff_31 = '2.87559e-06*lvp_mobility*lvp_mobility+9.28626e-05*lvp_mobility+3.62570e-04'
+ sky130_fd_pr__pfet_01v8__u0_diff_32 = '3.55281e-06*lvp_mobility*lvp_mobility+9.35313e-05*lvp_mobility+5.09260e-04'
+ sky130_fd_pr__pfet_01v8__u0_diff_33 = '6.01406e-06*lvp_mobility*lvp_mobility+8.31137e-05*lvp_mobility+6.10720e-04'
+ sky130_fd_pr__pfet_01v8__u0_diff_34 = '-1.02813e-06*lvp_mobility*lvp_mobility+-5.09125e-05*lvp_mobility+1.36990e-03'
+ sky130_fd_pr__pfet_01v8__u0_diff_35 = '-2.60708e-05*lvp_mobility*lvp_mobility+-3.48258e-04*lvp_mobility+1.71710e-03'
+ sky130_fd_pr__pfet_01v8__u0_diff_36 = '-1.79204e-05*lvp_mobility*lvp_mobility+3.16784e-05*lvp_mobility+1.28950e-04'
+ sky130_fd_pr__pfet_01v8__u0_diff_37 = '1.19033e-04*lvp_mobility*lvp_mobility+-4.20024e-04*lvp_mobility+-3.73230e-04'
+ sky130_fd_pr__pfet_01v8__u0_diff_38 = '9.08794e-05*lvp_mobility*lvp_mobility+-2.66160e-04*lvp_mobility+4.43390e-04'
+ sky130_fd_pr__pfet_01v8__u0_diff_39 = '-1.12425e-05*lvp_mobility*lvp_mobility+1.14943e-04*lvp_mobility+2.93840e-04'
+ sky130_fd_pr__pfet_01v8__u0_diff_4 = '4.99375e-07*lvp_mobility*lvp_mobility+-3.38252e-04*lvp_mobility+1.55430e-03'
+ sky130_fd_pr__pfet_01v8__u0_diff_40 = '-1.03638e-06*lvp_mobility*lvp_mobility+-6.58655e-05*lvp_mobility+3.41390e-04'
+ sky130_fd_pr__pfet_01v8__u0_diff_41 = '9.09303e-05*lvp_mobility*lvp_mobility+-5.84764e-04*lvp_mobility+4.97860e-04'
+ sky130_fd_pr__pfet_01v8__u0_diff_42 = '-2.28819e-05*lvp_mobility*lvp_mobility+-2.69527e-04*lvp_mobility+1.17030e-03'
+ sky130_fd_pr__pfet_01v8__u0_diff_43 = '5.55044e-05*lvp_mobility*lvp_mobility+-5.84407e-04*lvp_mobility+1.17850e-03'
+ sky130_fd_pr__pfet_01v8__u0_diff_44 = '-7.59406e-06*lvp_mobility*lvp_mobility+-3.68926e-04*lvp_mobility+1.72200e-03'
+ sky130_fd_pr__pfet_01v8__u0_diff_45 = '-1.77012e-05*lvp_mobility*lvp_mobility+9.43037e-05*lvp_mobility+9.60150e-05'
+ sky130_fd_pr__pfet_01v8__u0_diff_46 = '1.77969e-06*lvp_mobility*lvp_mobility+-4.51056e-04*lvp_mobility+1.65710e-03'
+ sky130_fd_pr__pfet_01v8__u0_diff_47 = '-1.45387e-05*lvp_mobility*lvp_mobility+-1.62590e-04*lvp_mobility+2.65240e-04'
+ sky130_fd_pr__pfet_01v8__u0_diff_48 = '-4.97366e-05*lvp_mobility*lvp_mobility+-2.22479e-04*lvp_mobility+1.15640e-03'
+ sky130_fd_pr__pfet_01v8__u0_diff_49 = '3.48724e-05*lvp_mobility*lvp_mobility+1.00802e-04*lvp_mobility+3.27510e-05'
+ sky130_fd_pr__pfet_01v8__u0_diff_5 = '-1.05437e-05*lvp_mobility*lvp_mobility+-2.93775e-04*lvp_mobility+1.41130e-03'
+ sky130_fd_pr__pfet_01v8__u0_diff_50 = '1.53825e-05*lvp_mobility*lvp_mobility+1.36867e-04*lvp_mobility+5.77710e-04'
+ sky130_fd_pr__pfet_01v8__u0_diff_51 = '9.25000e-08*lvp_mobility*lvp_mobility+4.89625e-05*lvp_mobility+5.62200e-04'
+ sky130_fd_pr__pfet_01v8__u0_diff_6 = '-3.30975e-05*lvp_mobility*lvp_mobility+5.26266e-05*lvp_mobility+4.44360e-04'
+ sky130_fd_pr__pfet_01v8__u0_diff_7 = '-7.62719e-06*lvp_mobility*lvp_mobility+-1.63999e-04*lvp_mobility+2.00570e-04'
+ sky130_fd_pr__pfet_01v8__u0_diff_8 = '-8.27187e-07*lvp_mobility*lvp_mobility+-1.49521e-04*lvp_mobility+-5.41380e-04'
+ sky130_fd_pr__pfet_01v8__u0_diff_9 = '-1.09897e-05*lvp_mobility*lvp_mobility+-1.38181e-04*lvp_mobility+7.93810e-04'
+ sky130_fd_pr__pfet_01v8__ua_diff_0 = '1.39598e-12*lvp_mobility*lvp_mobility+3.58983e-12*lvp_mobility+-1.03090e-11'
+ sky130_fd_pr__pfet_01v8__ua_diff_1 = '1.63084e-12*lvp_mobility*lvp_mobility+8.69413e-12*lvp_mobility+-2.95280e-11'
+ sky130_fd_pr__pfet_01v8__ua_diff_10 = '-1.50005e-11*lvp_mobility*lvp_mobility+7.48250e-12*lvp_mobility+-2.67420e-11'
+ sky130_fd_pr__pfet_01v8__ua_diff_11 = '5.96125e-13*lvp_mobility*lvp_mobility+2.61325e-12*lvp_mobility+-3.80000e-11'
+ sky130_fd_pr__pfet_01v8__ua_diff_12 = '2.93866e-13*lvp_mobility*lvp_mobility+5.48314e-13*lvp_mobility+-7.06670e-12'
+ sky130_fd_pr__pfet_01v8__ua_diff_13 = '2.72563e-14*lvp_mobility*lvp_mobility+2.25475e-13*lvp_mobility+-2.91210e-12'
+ sky130_fd_pr__pfet_01v8__ua_diff_14 = '1.59947e-13*lvp_mobility*lvp_mobility+3.97713e-13*lvp_mobility+-4.05910e-12'
+ sky130_fd_pr__pfet_01v8__ua_diff_15 = '1.00850e-11*lvp_mobility*lvp_mobility+-3.29194e-11*lvp_mobility+5.23250e-13'
+ sky130_fd_pr__pfet_01v8__ua_diff_16 = '7.75881e-13*lvp_mobility*lvp_mobility+-1.60745e-12*lvp_mobility+2.00710e-12'
+ sky130_fd_pr__pfet_01v8__ua_diff_17 = '3.04803e-12*lvp_mobility*lvp_mobility+3.97988e-12*lvp_mobility+-5.08890e-11'
+ sky130_fd_pr__pfet_01v8__ua_diff_18 = '8.69691e-13*lvp_mobility*lvp_mobility+1.26500e-13*lvp_mobility+9.29940e-13'
+ sky130_fd_pr__pfet_01v8__ua_diff_19 = '3.24125e-13*lvp_mobility*lvp_mobility+1.27930e-12*lvp_mobility+-9.32660e-12'
+ sky130_fd_pr__pfet_01v8__ua_diff_2 = '1.81608e-12*lvp_mobility*lvp_mobility+1.63769e-12*lvp_mobility+-1.89990e-11'
+ sky130_fd_pr__pfet_01v8__ua_diff_20 = '7.94094e-14*lvp_mobility*lvp_mobility+7.86250e-15*lvp_mobility+-3.62600e-12'
+ sky130_fd_pr__pfet_01v8__ua_diff_21 = '2.46844e-15*lvp_mobility*lvp_mobility+4.37749e-13*lvp_mobility+-2.45080e-12'
+ sky130_fd_pr__pfet_01v8__ua_diff_22 = '1.59675e-13*lvp_mobility*lvp_mobility+4.45625e-13*lvp_mobility+-2.97960e-12'
+ sky130_fd_pr__pfet_01v8__ua_diff_23 = '-1.33174e-11*lvp_mobility*lvp_mobility+5.98127e-11*lvp_mobility+-1.52050e-12'
+ sky130_fd_pr__pfet_01v8__ua_diff_24 = '8.07106e-13*lvp_mobility*lvp_mobility+2.53037e-12*lvp_mobility+-8.57920e-12'
+ sky130_fd_pr__pfet_01v8__ua_diff_25 = '7.69986e-13*lvp_mobility*lvp_mobility+2.54635e-12*lvp_mobility+-5.39170e-13'
+ sky130_fd_pr__pfet_01v8__ua_diff_26 = '8.82388e-13*lvp_mobility*lvp_mobility+-1.04812e-12*lvp_mobility+5.74530e-12'
+ sky130_fd_pr__pfet_01v8__ua_diff_27 = '7.30109e-13*lvp_mobility*lvp_mobility+-1.38786e-12*lvp_mobility+-1.08290e-11'
+ sky130_fd_pr__pfet_01v8__ua_diff_28 = '2.38756e-13*lvp_mobility*lvp_mobility+7.99500e-14*lvp_mobility+-7.24650e-12'
+ sky130_fd_pr__pfet_01v8__ua_diff_29 = '1.86983e-13*lvp_mobility*lvp_mobility+3.30655e-13*lvp_mobility+-3.57330e-12'
+ sky130_fd_pr__pfet_01v8__ua_diff_3 = '4.29044e-13*lvp_mobility*lvp_mobility+2.89276e-13*lvp_mobility+-8.11280e-12'
+ sky130_fd_pr__pfet_01v8__ua_diff_30 = '1.33970e-13*lvp_mobility*lvp_mobility+6.43256e-13*lvp_mobility+-5.09770e-12'
+ sky130_fd_pr__pfet_01v8__ua_diff_31 = '3.01250e-14*lvp_mobility*lvp_mobility+5.42512e-12*lvp_mobility+-3.58050e-12'
+ sky130_fd_pr__pfet_01v8__ua_diff_32 = '8.44256e-13*lvp_mobility*lvp_mobility+-1.12375e-13*lvp_mobility+4.83440e-12'
+ sky130_fd_pr__pfet_01v8__ua_diff_33 = '1.66363e-12*lvp_mobility*lvp_mobility+7.90240e-12*lvp_mobility+8.17830e-12'
+ sky130_fd_pr__pfet_01v8__ua_diff_34 = '-9.71031e-14*lvp_mobility*lvp_mobility+1.83141e-12*lvp_mobility+1.21520e-11'
+ sky130_fd_pr__pfet_01v8__ua_diff_35 = '3.31294e-13*lvp_mobility*lvp_mobility+-1.22340e-12*lvp_mobility+-8.81770e-12'
+ sky130_fd_pr__pfet_01v8__ua_diff_36 = '-4.85634e-13*lvp_mobility*lvp_mobility+4.81159e-12*lvp_mobility+-4.99550e-12'
+ sky130_fd_pr__pfet_01v8__ua_diff_37 = '-7.60250e-14*lvp_mobility*lvp_mobility+2.48825e-13*lvp_mobility+-4.99600e-12'
+ sky130_fd_pr__pfet_01v8__ua_diff_38 = '3.59099e-13*lvp_mobility*lvp_mobility+3.00629e-13*lvp_mobility+-4.92820e-12'
+ sky130_fd_pr__pfet_01v8__ua_diff_39 = '4.99450e-13*lvp_mobility*lvp_mobility+3.00137e-12*lvp_mobility+-7.19070e-12'
+ sky130_fd_pr__pfet_01v8__ua_diff_4 = '2.40729e-12*lvp_mobility*lvp_mobility+7.58530e-12*lvp_mobility+-7.82480e-12'
+ sky130_fd_pr__pfet_01v8__ua_diff_40 = '7.31444e-12*lvp_mobility*lvp_mobility+4.17952e-11*lvp_mobility+-2.75120e-11'
+ sky130_fd_pr__pfet_01v8__ua_diff_41 = '3.12103e-11*lvp_mobility*lvp_mobility+-1.03879e-10*lvp_mobility+-2.73200e-11'
+ sky130_fd_pr__pfet_01v8__ua_diff_42 = '1.94538e-12*lvp_mobility*lvp_mobility+6.55725e-12*lvp_mobility+-1.50500e-11'
+ sky130_fd_pr__pfet_01v8__ua_diff_43 = '2.17847e-11*lvp_mobility*lvp_mobility+-8.00853e-11*lvp_mobility+-3.00870e-11'
+ sky130_fd_pr__pfet_01v8__ua_diff_44 = '3.47296e-12*lvp_mobility*lvp_mobility+1.10758e-11*lvp_mobility+-1.74260e-12'
+ sky130_fd_pr__pfet_01v8__ua_diff_45 = '-3.12863e-13*lvp_mobility*lvp_mobility+-1.39225e-13*lvp_mobility+-4.87430e-12'
+ sky130_fd_pr__pfet_01v8__ua_diff_46 = '5.57509e-13*lvp_mobility*lvp_mobility+9.52538e-13*lvp_mobility+-7.58750e-12'
+ sky130_fd_pr__pfet_01v8__ua_diff_47 = '1.49469e-12*lvp_mobility*lvp_mobility+1.07060e-11*lvp_mobility+-2.31280e-11'
+ sky130_fd_pr__pfet_01v8__ua_diff_48 = '-1.35364e-11*lvp_mobility*lvp_mobility+-5.60621e-11*lvp_mobility+-1.26290e-11'
+ sky130_fd_pr__pfet_01v8__ua_diff_49 = '2.30003e-11*lvp_mobility*lvp_mobility+1.13194e-10*lvp_mobility+-1.20780e-10'
+ sky130_fd_pr__pfet_01v8__ua_diff_5 = '1.25657e-12*lvp_mobility*lvp_mobility+6.95723e-13*lvp_mobility+-2.35720e-11'
+ sky130_fd_pr__pfet_01v8__ua_diff_50 = '9.61925e-12*lvp_mobility*lvp_mobility+9.26525e-11*lvp_mobility+-2.45180e-11'
+ sky130_fd_pr__pfet_01v8__ua_diff_51 = '7.47000e-14*lvp_mobility*lvp_mobility+5.81750e-12*lvp_mobility+-6.74720e-12'
+ sky130_fd_pr__pfet_01v8__ua_diff_6 = '-1.33523e-11*lvp_mobility*lvp_mobility+6.48500e-11*lvp_mobility+-2.69630e-11'
+ sky130_fd_pr__pfet_01v8__ua_diff_7 = '3.06062e-13*lvp_mobility*lvp_mobility+-3.82350e-11*lvp_mobility+-2.92670e-11'
+ sky130_fd_pr__pfet_01v8__ua_diff_8 = '2.21090e-12*lvp_mobility*lvp_mobility+-3.33489e-12*lvp_mobility+-2.12980e-11'
+ sky130_fd_pr__pfet_01v8__ua_diff_9 = '4.02456e-13*lvp_mobility*lvp_mobility+-4.18225e-13*lvp_mobility+-7.01500e-12'
+ sky130_fd_pr__pfet_01v8__ub_diff_0 = '-2.45750e-22*lvp_mobility*lvp_mobility+-4.53130e-20*lvp_mobility+2.37660e-19'
+ sky130_fd_pr__pfet_01v8__ub_diff_1 = '-5.85531e-22*lvp_mobility*lvp_mobility+-2.88346e-20*lvp_mobility+1.99280e-19'
+ sky130_fd_pr__pfet_01v8__ub_diff_10 = '2.26338e-20*lvp_mobility*lvp_mobility+5.90050e-20*lvp_mobility+2.04700e-19'
+ sky130_fd_pr__pfet_01v8__ub_diff_11 = '-1.73125e-21*lvp_mobility*lvp_mobility+-3.78850e-20*lvp_mobility+3.73350e-19'
+ sky130_fd_pr__pfet_01v8__ub_diff_12 = '-1.06906e-21*lvp_mobility*lvp_mobility+-4.00637e-20*lvp_mobility+3.97540e-19'
+ sky130_fd_pr__pfet_01v8__ub_diff_13 = '-1.03125e-21*lvp_mobility*lvp_mobility+-4.99125e-20*lvp_mobility+3.83000e-19'
+ sky130_fd_pr__pfet_01v8__ub_diff_14 = '-2.52156e-21*lvp_mobility*lvp_mobility+-7.23637e-20*lvp_mobility+4.10370e-19'
+ sky130_fd_pr__pfet_01v8__ub_diff_15 = '-7.01431e-21*lvp_mobility*lvp_mobility+2.69348e-20*lvp_mobility+1.64150e-19'
+ sky130_fd_pr__pfet_01v8__ub_diff_16 = '-4.87500e-23*lvp_mobility*lvp_mobility+-2.12500e-22*lvp_mobility+1.94530e-19'
+ sky130_fd_pr__pfet_01v8__ub_diff_17 = '-1.01250e-21*lvp_mobility*lvp_mobility+-5.20000e-22*lvp_mobility+2.66120e-19'
+ sky130_fd_pr__pfet_01v8__ub_diff_18 = '-1.46891e-21*lvp_mobility*lvp_mobility+-3.86931e-20*lvp_mobility+2.23880e-19'
+ sky130_fd_pr__pfet_01v8__ub_diff_19 = '7.40000e-22*lvp_mobility*lvp_mobility+-2.21575e-20*lvp_mobility+2.63490e-19'
+ sky130_fd_pr__pfet_01v8__ub_diff_2 = '-4.21062e-21*lvp_mobility*lvp_mobility+-7.60800e-20*lvp_mobility+3.09750e-19'
+ sky130_fd_pr__pfet_01v8__ub_diff_20 = '-2.39375e-22*lvp_mobility*lvp_mobility+-2.25450e-20*lvp_mobility+2.73530e-19'
+ sky130_fd_pr__pfet_01v8__ub_diff_21 = '-1.04219e-21*lvp_mobility*lvp_mobility+-4.20688e-20*lvp_mobility+3.18490e-19'
+ sky130_fd_pr__pfet_01v8__ub_diff_22 = '-1.36000e-21*lvp_mobility*lvp_mobility+-4.28550e-20*lvp_mobility+3.54560e-19'
+ sky130_fd_pr__pfet_01v8__ub_diff_23 = '1.14247e-20*lvp_mobility*lvp_mobility+-3.12763e-20*lvp_mobility+1.67110e-19'
+ sky130_fd_pr__pfet_01v8__ub_diff_24 = '6.53125e-22*lvp_mobility*lvp_mobility+8.77000e-21*lvp_mobility+1.67680e-19'
+ sky130_fd_pr__pfet_01v8__ub_diff_25 = '9.62188e-22*lvp_mobility*lvp_mobility+1.44888e-20*lvp_mobility+2.43810e-19'
+ sky130_fd_pr__pfet_01v8__ub_diff_26 = '-4.67500e-22*lvp_mobility*lvp_mobility+-1.43550e-20*lvp_mobility+2.80550e-19'
+ sky130_fd_pr__pfet_01v8__ub_diff_27 = '-9.99375e-22*lvp_mobility*lvp_mobility+-2.88675e-20*lvp_mobility+2.90280e-19'
+ sky130_fd_pr__pfet_01v8__ub_diff_28 = '-6.75312e-22*lvp_mobility*lvp_mobility+-2.65387e-20*lvp_mobility+2.95800e-19'
+ sky130_fd_pr__pfet_01v8__ub_diff_29 = '-1.29688e-21*lvp_mobility*lvp_mobility+-3.97525e-20*lvp_mobility+3.65940e-19'
+ sky130_fd_pr__pfet_01v8__ub_diff_3 = '-3.04972e-21*lvp_mobility*lvp_mobility+-8.35614e-20*lvp_mobility+3.49610e-19'
+ sky130_fd_pr__pfet_01v8__ub_diff_30 = '-9.80312e-22*lvp_mobility*lvp_mobility+-3.61513e-20*lvp_mobility+3.94610e-19'
+ sky130_fd_pr__pfet_01v8__ub_diff_31 = '2.45250e-21*lvp_mobility*lvp_mobility+1.62150e-20*lvp_mobility+1.46850e-19'
+ sky130_fd_pr__pfet_01v8__ub_diff_32 = '1.47938e-21*lvp_mobility*lvp_mobility+2.62225e-20*lvp_mobility+1.88500e-19'
+ sky130_fd_pr__pfet_01v8__ub_diff_33 = '6.38125e-22*lvp_mobility*lvp_mobility+1.43300e-20*lvp_mobility+2.20260e-19'
+ sky130_fd_pr__pfet_01v8__ub_diff_34 = '5.38125e-22*lvp_mobility*lvp_mobility+-2.67425e-20*lvp_mobility+2.80170e-19'
+ sky130_fd_pr__pfet_01v8__ub_diff_35 = '-3.38584e-21*lvp_mobility*lvp_mobility+-8.04409e-20*lvp_mobility+3.34940e-19'
+ sky130_fd_pr__pfet_01v8__ub_diff_36 = '-1.94125e-23*lvp_mobility*lvp_mobility+-3.32123e-21*lvp_mobility+7.67070e-21'
+ sky130_fd_pr__pfet_01v8__ub_diff_37 = '2.68218e-20*lvp_mobility*lvp_mobility+-9.30260e-20*lvp_mobility+-7.04530e-20'
+ sky130_fd_pr__pfet_01v8__ub_diff_38 = '1.92390e-20*lvp_mobility*lvp_mobility+-7.01464e-20*lvp_mobility+1.42800e-20'
+ sky130_fd_pr__pfet_01v8__ub_diff_39 = '-1.06338e-21*lvp_mobility*lvp_mobility+6.14650e-21*lvp_mobility+1.42670e-20'
+ sky130_fd_pr__pfet_01v8__ub_diff_4 = '-2.36631e-21*lvp_mobility*lvp_mobility+-8.29527e-20*lvp_mobility+3.23880e-19'
+ sky130_fd_pr__pfet_01v8__ub_diff_40 = '-7.24563e-21*lvp_mobility*lvp_mobility+-1.29312e-19*lvp_mobility+2.11950e-19'
+ sky130_fd_pr__pfet_01v8__ub_diff_41 = '-1.32003e-20*lvp_mobility*lvp_mobility+-6.14963e-20*lvp_mobility+2.70270e-19'
+ sky130_fd_pr__pfet_01v8__ub_diff_42 = '-5.05437e-21*lvp_mobility*lvp_mobility+-9.14975e-20*lvp_mobility+2.78140e-19'
+ sky130_fd_pr__pfet_01v8__ub_diff_43 = '-1.90819e-20*lvp_mobility*lvp_mobility+-8.36700e-21*lvp_mobility+2.77970e-19'
+ sky130_fd_pr__pfet_01v8__ub_diff_44 = '-5.42375e-21*lvp_mobility*lvp_mobility+-1.02715e-19*lvp_mobility+3.44670e-19'
+ sky130_fd_pr__pfet_01v8__ub_diff_45 = '-4.20003e-22*lvp_mobility*lvp_mobility+4.68574e-21*lvp_mobility+-1.30620e-20'
+ sky130_fd_pr__pfet_01v8__ub_diff_46 = '2.07432e-21*lvp_mobility*lvp_mobility+-8.64852e-20*lvp_mobility+3.13090e-19'
+ sky130_fd_pr__pfet_01v8__ub_diff_47 = '-2.48625e-21*lvp_mobility*lvp_mobility+-9.55700e-20*lvp_mobility+2.36700e-19'
+ sky130_fd_pr__pfet_01v8__ub_diff_48 = '6.91375e-21*lvp_mobility*lvp_mobility+-2.11275e-20*lvp_mobility+2.93910e-19'
+ sky130_fd_pr__pfet_01v8__ub_diff_49 = '-2.43809e-20*lvp_mobility*lvp_mobility+-1.96676e-19*lvp_mobility+2.26380e-19'
+ sky130_fd_pr__pfet_01v8__ub_diff_5 = '-3.35581e-21*lvp_mobility*lvp_mobility+-6.23933e-20*lvp_mobility+3.21810e-19'
+ sky130_fd_pr__pfet_01v8__ub_diff_50 = '-9.89031e-21*lvp_mobility*lvp_mobility+-1.32886e-19*lvp_mobility+2.71210e-19'
+ sky130_fd_pr__pfet_01v8__ub_diff_51 = '1.41875e-21*lvp_mobility*lvp_mobility+-1.52300e-20*lvp_mobility+2.31630e-19'
+ sky130_fd_pr__pfet_01v8__ub_diff_6 = '1.23578e-20*lvp_mobility*lvp_mobility+-9.23737e-20*lvp_mobility+2.15280e-19'
+ sky130_fd_pr__pfet_01v8__ub_diff_7 = '8.75000e-23*lvp_mobility*lvp_mobility+-7.86500e-21*lvp_mobility+1.89970e-19'
+ sky130_fd_pr__pfet_01v8__ub_diff_8 = '-8.50313e-22*lvp_mobility*lvp_mobility+-3.86562e-20*lvp_mobility+1.50690e-19'
+ sky130_fd_pr__pfet_01v8__ub_diff_9 = '-2.45056e-21*lvp_mobility*lvp_mobility+-6.06973e-20*lvp_mobility+2.42470e-19'
+ sky130_fd_pr__pfet_01v8__voff_diff_0 = '1.84528e-03*lvp_subvt*lvp_subvt+3.70986e-02*lvp_subvt+-1.15980e-01'
+ sky130_fd_pr__pfet_01v8__voff_diff_1 = '1.99084e-03*lvp_subvt*lvp_subvt+3.30734e-02*lvp_subvt+-1.09520e-01'
+ sky130_fd_pr__pfet_01v8__voff_diff_10 = '3.75750e-03*lvp_subvt*lvp_subvt+7.23000e-03*lvp_subvt+-1.32330e-01'
+ sky130_fd_pr__pfet_01v8__voff_diff_11 = '-2.02359e-04*lvp_subvt*lvp_subvt+1.27293e-02*lvp_subvt+-5.58550e-02'
+ sky130_fd_pr__pfet_01v8__voff_diff_12 = '-2.57484e-04*lvp_subvt*lvp_subvt+1.18046e-02*lvp_subvt+-5.17620e-02'
+ sky130_fd_pr__pfet_01v8__voff_diff_13 = '-2.11594e-04*lvp_subvt*lvp_subvt+1.00219e-02*lvp_subvt+-4.83430e-02'
+ sky130_fd_pr__pfet_01v8__voff_diff_14 = '-1.12209e-04*lvp_subvt*lvp_subvt+1.07142e-02*lvp_subvt+-3.84210e-02'
+ sky130_fd_pr__pfet_01v8__voff_diff_15 = '1.98247e-03*lvp_subvt*lvp_subvt+2.69369e-02*lvp_subvt+-9.71020e-02'
+ sky130_fd_pr__pfet_01v8__voff_diff_16 = '-6.98944e-04*lvp_subvt*lvp_subvt+3.49017e-02*lvp_subvt+-1.21180e-01'
+ sky130_fd_pr__pfet_01v8__voff_diff_17 = '-8.34244e-04*lvp_subvt*lvp_subvt+2.72888e-02*lvp_subvt+-8.99170e-02'
+ sky130_fd_pr__pfet_01v8__voff_diff_18 = '-6.85831e-04*lvp_subvt*lvp_subvt+1.79934e-02*lvp_subvt+-5.89230e-02'
+ sky130_fd_pr__pfet_01v8__voff_diff_19 = '-5.52453e-04*lvp_subvt*lvp_subvt+1.10612e-02*lvp_subvt+-3.84210e-02'
+ sky130_fd_pr__pfet_01v8__voff_diff_2 = '3.72250e-04*lvp_subvt*lvp_subvt+9.47375e-03*lvp_subvt+-6.57390e-02'
+ sky130_fd_pr__pfet_01v8__voff_diff_20 = '-2.52866e-04*lvp_subvt*lvp_subvt+9.65054e-03*lvp_subvt+-4.32210e-02'
+ sky130_fd_pr__pfet_01v8__voff_diff_21 = '-1.92219e-04*lvp_subvt*lvp_subvt+8.77013e-03*lvp_subvt+-4.30220e-02'
+ sky130_fd_pr__pfet_01v8__voff_diff_22 = '-9.67000e-05*lvp_subvt*lvp_subvt+9.02170e-03*lvp_subvt+-4.10620e-02'
+ sky130_fd_pr__pfet_01v8__voff_diff_23 = '3.60316e-03*lvp_subvt*lvp_subvt+2.49651e-02*lvp_subvt+-1.26280e-01'
+ sky130_fd_pr__pfet_01v8__voff_diff_24 = '-9.67656e-04*lvp_subvt*lvp_subvt+3.49559e-02*lvp_subvt+-9.93240e-02'
+ sky130_fd_pr__pfet_01v8__voff_diff_25 = '-2.01074e-03*lvp_subvt*lvp_subvt+2.59323e-02*lvp_subvt+-6.79690e-02'
+ sky130_fd_pr__pfet_01v8__voff_diff_26 = '-3.49784e-04*lvp_subvt*lvp_subvt+1.27294e-02*lvp_subvt+-4.19180e-02'
+ sky130_fd_pr__pfet_01v8__voff_diff_27 = '-1.27947e-04*lvp_subvt*lvp_subvt+9.80471e-03*lvp_subvt+-3.15860e-02'
+ sky130_fd_pr__pfet_01v8__voff_diff_28 = '-1.25031e-04*lvp_subvt*lvp_subvt+8.16862e-03*lvp_subvt+-4.34360e-02'
+ sky130_fd_pr__pfet_01v8__voff_diff_29 = '-1.02844e-04*lvp_subvt*lvp_subvt+8.33937e-03*lvp_subvt+-4.52970e-02'
+ sky130_fd_pr__pfet_01v8__voff_diff_3 = '7.44519e-04*lvp_subvt*lvp_subvt+1.22363e-02*lvp_subvt+-6.84270e-02'
+ sky130_fd_pr__pfet_01v8__voff_diff_30 = '-5.80625e-05*lvp_subvt*lvp_subvt+9.13775e-03*lvp_subvt+-5.09260e-02'
+ sky130_fd_pr__pfet_01v8__voff_diff_31 = '1.85189e-03*lvp_subvt*lvp_subvt+2.32900e-02*lvp_subvt+-1.27230e-01'
+ sky130_fd_pr__pfet_01v8__voff_diff_32 = '-9.65156e-04*lvp_subvt*lvp_subvt+2.46389e-02*lvp_subvt+-4.72620e-02'
+ sky130_fd_pr__pfet_01v8__voff_diff_33 = '-1.13853e-03*lvp_subvt*lvp_subvt+1.92991e-02*lvp_subvt+-4.15270e-02'
+ sky130_fd_pr__pfet_01v8__voff_diff_34 = '-7.08188e-04*lvp_subvt*lvp_subvt+1.02575e-02*lvp_subvt+-5.75790e-02'
+ sky130_fd_pr__pfet_01v8__voff_diff_35 = '9.48656e-04*lvp_subvt*lvp_subvt+2.62259e-02*lvp_subvt+-9.57050e-02'
+ sky130_fd_pr__pfet_01v8__voff_diff_36 = '-1.12500e-05*lvp_subvt*lvp_subvt+1.98460e-02*lvp_subvt+-3.04560e-02'
+ sky130_fd_pr__pfet_01v8__voff_diff_37 = '-1.69800e-03*lvp_subvt*lvp_subvt+2.03583e-02*lvp_subvt+-3.71790e-02'
+ sky130_fd_pr__pfet_01v8__voff_diff_38 = '-1.45206e-03*lvp_subvt*lvp_subvt+1.83082e-02*lvp_subvt+-3.69940e-02'
+ sky130_fd_pr__pfet_01v8__voff_diff_39 = '2.48666e-04*lvp_subvt*lvp_subvt+8.18616e-03*lvp_subvt+-3.03520e-02'
+ sky130_fd_pr__pfet_01v8__voff_diff_4 = '7.61209e-04*lvp_subvt*lvp_subvt+1.29526e-02*lvp_subvt+-6.63590e-02'
+ sky130_fd_pr__pfet_01v8__voff_diff_40 = '2.58219e-03*lvp_subvt*lvp_subvt+4.03663e-02*lvp_subvt+-1.02780e-01'
+ sky130_fd_pr__pfet_01v8__voff_diff_41 = '7.39406e-03*lvp_subvt*lvp_subvt+4.39937e-02*lvp_subvt+-1.94280e-01'
+ sky130_fd_pr__pfet_01v8__voff_diff_42 = '9.60594e-04*lvp_subvt*lvp_subvt+3.44449e-02*lvp_subvt+-8.90000e-02'
+ sky130_fd_pr__pfet_01v8__voff_diff_43 = '4.70069e-03*lvp_subvt*lvp_subvt+1.69063e-02*lvp_subvt+-8.38040e-02'
+ sky130_fd_pr__pfet_01v8__voff_diff_44 = '7.34741e-04*lvp_subvt*lvp_subvt+1.43547e-02*lvp_subvt+-7.13070e-02'
+ sky130_fd_pr__pfet_01v8__voff_diff_45 = '7.43625e-04*lvp_subvt*lvp_subvt+8.94400e-03*lvp_subvt+-3.54230e-02'
+ sky130_fd_pr__pfet_01v8__voff_diff_46 = '1.17166e-03*lvp_subvt*lvp_subvt+1.97399e-02*lvp_subvt+-8.25670e-02'
+ sky130_fd_pr__pfet_01v8__voff_diff_47 = '6.00375e-03*lvp_subvt*lvp_subvt+4.02600e-02*lvp_subvt+-1.57100e-01'
+ sky130_fd_pr__pfet_01v8__voff_diff_48 = '1.82313e-03*lvp_subvt*lvp_subvt+3.08162e-02*lvp_subvt+-8.00250e-02'
+ sky130_fd_pr__pfet_01v8__voff_diff_49 = '-5.07002e-03*lvp_subvt*lvp_subvt+2.27464e-02*lvp_subvt+-5.27400e-03'
+ sky130_fd_pr__pfet_01v8__voff_diff_5 = '9.26172e-04*lvp_subvt*lvp_subvt+1.54829e-02*lvp_subvt+-7.34970e-02'
+ sky130_fd_pr__pfet_01v8__voff_diff_50 = '1.29687e-03*lvp_subvt*lvp_subvt+3.22650e-02*lvp_subvt+-4.98100e-02'
+ sky130_fd_pr__pfet_01v8__voff_diff_51 = '1.40006e-03*lvp_subvt*lvp_subvt+3.97462e-02*lvp_subvt+-8.13860e-02'
+ sky130_fd_pr__pfet_01v8__voff_diff_6 = '3.78162e-03*lvp_subvt*lvp_subvt+2.92865e-02*lvp_subvt+-1.05450e-01'
+ sky130_fd_pr__pfet_01v8__voff_diff_7 = '4.88406e-04*lvp_subvt*lvp_subvt+3.63611e-02*lvp_subvt+-1.24520e-01'
+ sky130_fd_pr__pfet_01v8__voff_diff_8 = '-8.45187e-04*lvp_subvt*lvp_subvt+3.08185e-02*lvp_subvt+-7.05630e-02'
+ sky130_fd_pr__pfet_01v8__voff_diff_9 = '-1.06575e-04*lvp_subvt*lvp_subvt+1.42927e-02*lvp_subvt+-5.69140e-02'
+ sky130_fd_pr__pfet_01v8__vsat_diff_0 = '-1.04972e+03*lvp_saturation*lvp_saturation+3.16912e+03*lvp_saturation+1.64310e+04'
+ sky130_fd_pr__pfet_01v8__vsat_diff_1 = '-5.65789e+02*lvp_saturation*lvp_saturation+1.64989e+03*lvp_saturation+-3.75820e+02'
+ sky130_fd_pr__pfet_01v8__vsat_diff_10 = '2.21887e+03*lvp_saturation*lvp_saturation+1.50000e+04*lvp_saturation+4.49810e+03'
+ sky130_fd_pr__pfet_01v8__vsat_diff_11 = '-2.03906e+02*lvp_saturation*lvp_saturation+-9.35625e+02*lvp_saturation+2.67140e+04'
+ sky130_fd_pr__pfet_01v8__vsat_diff_15 = '-3.95987e+02*lvp_saturation*lvp_saturation+1.60130e+03*lvp_saturation+-7.25900e+03'
+ sky130_fd_pr__pfet_01v8__vsat_diff_16 = '-6.56250e+02*lvp_saturation*lvp_saturation+3.71388e+03*lvp_saturation+8.56750e+03'
+ sky130_fd_pr__pfet_01v8__vsat_diff_17 = '-2.32690e+03*lvp_saturation*lvp_saturation+-2.80435e+03*lvp_saturation+5.67930e+04'
+ sky130_fd_pr__pfet_01v8__vsat_diff_18 = '-1.00800e+03*lvp_saturation*lvp_saturation+-3.82500e+03*lvp_saturation+1.59860e+04'
+ sky130_fd_pr__pfet_01v8__vsat_diff_23 = '-4.98528e+02*lvp_saturation*lvp_saturation+2.25904e+03*lvp_saturation+-2.98740e+03'
+ sky130_fd_pr__pfet_01v8__vsat_diff_24 = '-8.23337e+02*lvp_saturation*lvp_saturation+1.42022e+03*lvp_saturation+1.51650e+04'
+ sky130_fd_pr__pfet_01v8__vsat_diff_25 = '-9.00925e+02*lvp_saturation*lvp_saturation+-2.77528e+03*lvp_saturation+7.60290e+03'
+ sky130_fd_pr__pfet_01v8__vsat_diff_26 = '-5.66150e+02*lvp_saturation*lvp_saturation+1.46932e+03*lvp_saturation+7.61280e+03'
+ sky130_fd_pr__pfet_01v8__vsat_diff_31 = '-4.64388e+02*lvp_saturation*lvp_saturation+1.16383e+03*lvp_saturation+-4.71650e+03'
+ sky130_fd_pr__pfet_01v8__vsat_diff_32 = '-6.97209e+02*lvp_saturation*lvp_saturation+1.58389e+03*lvp_saturation+8.57060e+03'
+ sky130_fd_pr__pfet_01v8__vsat_diff_33 = '-1.10430e+03*lvp_saturation*lvp_saturation+-3.52305e+03*lvp_saturation+1.17610e+04'
+ sky130_fd_pr__pfet_01v8__vsat_diff_34 = '4.13299e+02*lvp_saturation*lvp_saturation+-2.24948e+03*lvp_saturation+2.99830e+03'
+ sky130_fd_pr__pfet_01v8__vsat_diff_36 = '-1.25000e-01*lvp_saturation*lvp_saturation+-1.00000e+00*lvp_saturation+2.00040e+04'
+ sky130_fd_pr__pfet_01v8__vsat_diff_39 = '-1.25119e+03*lvp_saturation*lvp_saturation+2.00190e+04'
+ sky130_fd_pr__pfet_01v8__vsat_diff_40 = '-6.97500e+01*lvp_saturation*lvp_saturation+9.47500e+01*lvp_saturation+1.96870e+04'
+ sky130_fd_pr__pfet_01v8__vsat_diff_41 = '2.83438e+01*lvp_saturation*lvp_saturation+-2.12125e+02*lvp_saturation+1.96600e+04'
+ sky130_fd_pr__pfet_01v8__vsat_diff_42 = '-4.95938e+01*lvp_saturation*lvp_saturation+-4.11250e+01*lvp_saturation+2.04660e+04'
+ sky130_fd_pr__pfet_01v8__vsat_diff_43 = '3.10531e+03*lvp_saturation*lvp_saturation+-1.25052e+04*lvp_saturation+2.02240e+04'
+ sky130_fd_pr__pfet_01v8__vsat_diff_45 = '-6.26938e+02*lvp_saturation*lvp_saturation+2.50300e+03*lvp_saturation+2.00430e+04'
+ sky130_fd_pr__pfet_01v8__vsat_diff_47 = '2.50000e+01*lvp_saturation*lvp_saturation+-2.82250e+02*lvp_saturation+2.00300e+04'
+ sky130_fd_pr__pfet_01v8__vsat_diff_48 = '-6.44625e+02*lvp_saturation*lvp_saturation+-2.47625e+03*lvp_saturation+2.02190e+04'
+ sky130_fd_pr__pfet_01v8__vsat_diff_49 = '1.00000e+01*lvp_saturation*lvp_saturation+-6.23250e+02*lvp_saturation+2.15780e+04'
+ sky130_fd_pr__pfet_01v8__vsat_diff_50 = '1.55882e+02*lvp_saturation*lvp_saturation+5.61700e+03*lvp_saturation+-2.61090e+01'
+ sky130_fd_pr__pfet_01v8__vsat_diff_51 = '-1.99375e+02*lvp_saturation*lvp_saturation+3.99288e+03*lvp_saturation+2.38750e+03'
+ sky130_fd_pr__pfet_01v8__vsat_diff_6 = '4.56256e+01*lvp_saturation*lvp_saturation+5.51688e+03*lvp_saturation+1.10490e+02'
+ sky130_fd_pr__pfet_01v8__vsat_diff_7 = '1.23150e+03*lvp_saturation*lvp_saturation+1.50000e+04*lvp_saturation+2.02960e+04'
+ sky130_fd_pr__pfet_01v8__vsat_diff_8 = '-3.01847e+03*lvp_saturation*lvp_saturation+3.96362e+03*lvp_saturation+5.24970e+04'
+ sky130_fd_pr__pfet_01v8__vsat_diff_9 = '-1.04415e+03*lvp_saturation*lvp_saturation+5.63587e+02*lvp_saturation+1.59280e+04'
+ sky130_fd_pr__pfet_01v8__vth0_diff_0 = '-2.08684e-03*lvp_threshold*lvp_threshold+1.43804e-02*lvp_threshold+3.59530e-02'
+ sky130_fd_pr__pfet_01v8__vth0_diff_1 = '-2.18450e-03*lvp_threshold*lvp_threshold+1.86855e-02*lvp_threshold+-1.70060e-02'
+ sky130_fd_pr__pfet_01v8__vth0_diff_10 = '3.41116e-04*lvp_threshold*lvp_threshold+9.77596e-03*lvp_threshold+-5.27390e-02'
+ sky130_fd_pr__pfet_01v8__vth0_diff_11 = '1.11475e-04*lvp_threshold*lvp_threshold+-3.98390e-03*lvp_threshold+-1.41310e-02'
+ sky130_fd_pr__pfet_01v8__vth0_diff_12 = '7.41031e-05*lvp_threshold*lvp_threshold+-3.18791e-03*lvp_threshold+-1.01810e-02'
+ sky130_fd_pr__pfet_01v8__vth0_diff_13 = '5.95556e-05*lvp_threshold*lvp_threshold+-3.14138e-03*lvp_threshold+-3.58390e-04'
+ sky130_fd_pr__pfet_01v8__vth0_diff_14 = '1.27941e-04*lvp_threshold*lvp_threshold+-2.80311e-03*lvp_threshold+2.42350e-03'
+ sky130_fd_pr__pfet_01v8__vth0_diff_15 = '-2.50291e-03*lvp_threshold*lvp_threshold+2.43549e-02*lvp_threshold+-2.74840e-02'
+ sky130_fd_pr__pfet_01v8__vth0_diff_16 = '-1.10076e-03*lvp_threshold*lvp_threshold+1.32889e-02*lvp_threshold+-5.72430e-03'
+ sky130_fd_pr__pfet_01v8__vth0_diff_17 = '-4.20500e-04*lvp_threshold*lvp_threshold+1.79825e-03*lvp_threshold+-1.77960e-02'
+ sky130_fd_pr__pfet_01v8__vth0_diff_18 = '1.85375e-05*lvp_threshold*lvp_threshold+-4.11875e-03*lvp_threshold+1.87840e-03'
+ sky130_fd_pr__pfet_01v8__vth0_diff_19 = '-1.03563e-04*lvp_threshold*lvp_threshold+-4.03500e-03*lvp_threshold+6.90000e-03'
+ sky130_fd_pr__pfet_01v8__vth0_diff_2 = '2.80531e-04*lvp_threshold*lvp_threshold+-4.37875e-03*lvp_threshold+-5.80450e-03'
+ sky130_fd_pr__pfet_01v8__vth0_diff_20 = '2.83000e-05*lvp_threshold*lvp_threshold+-3.69687e-03*lvp_threshold+1.37770e-03'
+ sky130_fd_pr__pfet_01v8__vth0_diff_21 = '5.72031e-05*lvp_threshold*lvp_threshold+-3.54736e-03*lvp_threshold+4.80830e-03'
+ sky130_fd_pr__pfet_01v8__vth0_diff_22 = '6.97088e-05*lvp_threshold*lvp_threshold+-2.94661e-03*lvp_threshold+8.64210e-04'
+ sky130_fd_pr__pfet_01v8__vth0_diff_23 = '5.58125e-05*lvp_threshold*lvp_threshold+1.76405e-02*lvp_threshold+-2.58130e-02'
+ sky130_fd_pr__pfet_01v8__vth0_diff_24 = '-1.14266e-03*lvp_threshold*lvp_threshold+1.39094e-02*lvp_threshold+-1.62910e-02'
+ sky130_fd_pr__pfet_01v8__vth0_diff_25 = '-3.45563e-04*lvp_threshold*lvp_threshold+3.75525e-03*lvp_threshold+-2.57500e-02'
+ sky130_fd_pr__pfet_01v8__vth0_diff_26 = '-1.40875e-05*lvp_threshold*lvp_threshold+-3.71487e-03*lvp_threshold+-3.39410e-03'
+ sky130_fd_pr__pfet_01v8__vth0_diff_27 = '5.33875e-05*lvp_threshold*lvp_threshold+-2.76775e-03*lvp_threshold+-1.09620e-03'
+ sky130_fd_pr__pfet_01v8__vth0_diff_28 = '4.12969e-05*lvp_threshold*lvp_threshold+-3.48354e-03*lvp_threshold+3.54110e-03'
+ sky130_fd_pr__pfet_01v8__vth0_diff_29 = '5.64244e-05*lvp_threshold*lvp_threshold+-2.99850e-03*lvp_threshold+8.05210e-04'
+ sky130_fd_pr__pfet_01v8__vth0_diff_3 = '3.39756e-04*lvp_threshold*lvp_threshold+-4.19197e-03*lvp_threshold+-7.22990e-04'
+ sky130_fd_pr__pfet_01v8__vth0_diff_30 = '5.53444e-05*lvp_threshold*lvp_threshold+-2.67850e-03*lvp_threshold+-2.53510e-04'
+ sky130_fd_pr__pfet_01v8__vth0_diff_31 = '-2.13447e-03*lvp_threshold*lvp_threshold+2.40561e-02*lvp_threshold+-2.75140e-02'
+ sky130_fd_pr__pfet_01v8__vth0_diff_32 = '-1.10959e-03*lvp_threshold*lvp_threshold+1.47369e-02*lvp_threshold+-1.47030e-02'
+ sky130_fd_pr__pfet_01v8__vth0_diff_33 = '-3.71031e-04*lvp_threshold*lvp_threshold+3.37838e-03*lvp_threshold+-2.38520e-02'
+ sky130_fd_pr__pfet_01v8__vth0_diff_34 = '-1.23709e-04*lvp_threshold*lvp_threshold+-7.22787e-04*lvp_threshold+-2.01030e-03'
+ sky130_fd_pr__pfet_01v8__vth0_diff_35 = '9.01219e-04*lvp_threshold*lvp_threshold+-7.80088e-03*lvp_threshold+-3.19990e-02'
+ sky130_fd_pr__pfet_01v8__vth0_diff_36 = '3.34719e-04*lvp_threshold*lvp_threshold+-7.15737e-03*lvp_threshold+2.14700e-03'
+ sky130_fd_pr__pfet_01v8__vth0_diff_37 = '-1.20413e-03*lvp_threshold*lvp_threshold+-7.40525e-03*lvp_threshold+2.20990e-02'
+ sky130_fd_pr__pfet_01v8__vth0_diff_38 = '-1.09569e-03*lvp_threshold*lvp_threshold+-4.34177e-03*lvp_threshold+5.68120e-04'
+ sky130_fd_pr__pfet_01v8__vth0_diff_39 = '1.44000e-04*lvp_threshold*lvp_threshold+-1.45429e-02*lvp_threshold+4.82750e-03'
+ sky130_fd_pr__pfet_01v8__vth0_diff_4 = '5.83066e-04*lvp_threshold*lvp_threshold+-2.59851e-03*lvp_threshold+-1.30350e-02'
+ sky130_fd_pr__pfet_01v8__vth0_diff_40 = '-1.11549e-03*lvp_threshold*lvp_threshold+-1.81496e-03*lvp_threshold+2.15870e-02'
+ sky130_fd_pr__pfet_01v8__vth0_diff_41 = '2.51312e-04*lvp_threshold*lvp_threshold+1.10105e-02*lvp_threshold+3.90210e-02'
+ sky130_fd_pr__pfet_01v8__vth0_diff_42 = '1.44487e-03*lvp_threshold*lvp_threshold+-8.07650e-03*lvp_threshold+-1.75650e-02'
+ sky130_fd_pr__pfet_01v8__vth0_diff_43 = '6.08687e-04*lvp_threshold*lvp_threshold+-4.49600e-03*lvp_threshold+-3.88930e-02'
+ sky130_fd_pr__pfet_01v8__vth0_diff_44 = '5.36649e-04*lvp_threshold*lvp_threshold+-4.47631e-03*lvp_threshold+5.95360e-04'
+ sky130_fd_pr__pfet_01v8__vth0_diff_45 = '1.48512e-03*lvp_threshold*lvp_threshold+-9.65164e-03*lvp_threshold+5.55750e-03'
+ sky130_fd_pr__pfet_01v8__vth0_diff_46 = '9.08213e-04*lvp_threshold*lvp_threshold+-2.63010e-03*lvp_threshold+-2.10940e-02'
+ sky130_fd_pr__pfet_01v8__vth0_diff_47 = '1.80969e-04*lvp_threshold*lvp_threshold+1.14771e-02*lvp_threshold+2.96470e-02'
+ sky130_fd_pr__pfet_01v8__vth0_diff_48 = '1.96826e-03*lvp_threshold*lvp_threshold+-2.37650e-03*lvp_threshold+-2.09920e-03'
+ sky130_fd_pr__pfet_01v8__vth0_diff_49 = '-1.76091e-03*lvp_threshold*lvp_threshold+7.26912e-03*lvp_threshold+-4.54090e-02'
+ sky130_fd_pr__pfet_01v8__vth0_diff_5 = '9.72916e-04*lvp_threshold*lvp_threshold+2.91087e-04*lvp_threshold+-2.36870e-02'
+ sky130_fd_pr__pfet_01v8__vth0_diff_50 = '-2.23153e-03*lvp_threshold*lvp_threshold+1.15259e-02*lvp_threshold+-4.26620e-02'
+ sky130_fd_pr__pfet_01v8__vth0_diff_51 = '-2.18039e-03*lvp_threshold*lvp_threshold+1.88592e-02*lvp_threshold+1.26330e-03'
+ sky130_fd_pr__pfet_01v8__vth0_diff_6 = '-9.48156e-05*lvp_threshold*lvp_threshold+1.22615e-02*lvp_threshold+-5.21570e-02'
+ sky130_fd_pr__pfet_01v8__vth0_diff_7 = '-5.59606e-04*lvp_threshold*lvp_threshold+1.02758e-02*lvp_threshold+-3.64650e-02'
+ sky130_fd_pr__pfet_01v8__vth0_diff_8 = '-3.90721e-04*lvp_threshold*lvp_threshold+-3.64288e-03*lvp_threshold+2.05320e-02'
+ sky130_fd_pr__pfet_01v8__vth0_diff_9 = '1.22221e-04*lvp_threshold*lvp_threshold+-5.50987e-03*lvp_threshold+2.07330e-02'
+ sky130_fd_pr__pfet_01v8__wint_diff = '8.04375e-09*diff_cd'
+ sky130_fd_pr__pfet_g5v0d16v0__ajunction_mult = '-2.50000e-06*hvp_diode*hvp_diode+1.81850e-02*hvp_diode+1.00500e+00'
+ sky130_fd_pr__pfet_g5v0d16v0__dlc_diff = '-4.33125e-09*poly_cd'
+ sky130_fd_pr__pfet_g5v0d16v0__doverlap_mult = '3.12500e-03*hvtox*hvtox+2.25000e-01*hvtox+1.00000e+00'
+ sky130_fd_pr__pfet_g5v0d16v0__dwc_diff = '8.04375e-09*diff_cd'
+ sky130_fd_pr__pfet_g5v0d16v0__lint_diff = '-4.33125e-09*poly_cd'
+ sky130_fd_pr__pfet_g5v0d16v0__pjunction_mult = '-1.25000e-06*hvp_diode*hvp_diode+1.61550e-02*hvp_diode+1.00900e+00'
+ sky130_fd_pr__pfet_g5v0d16v0__rdiff_mult = '1.31656e-02*pfet_g5v0d16v0*pfet_g5v0d16v0+1.62338e-01*pfet_g5v0d16v0+1.04110e+00'
+ sky130_fd_pr__pfet_g5v0d16v0__soverlap_mult = '3.12500e-03*hvtox*hvtox+2.25000e-01*hvtox+1.00000e+00'
+ sky130_fd_pr__pfet_g5v0d16v0__toxe_mult = '1.30000e-02*hvtox+1.00000e+00'
+ sky130_fd_pr__pfet_g5v0d16v0__u0_diff_0 = '-1.39312e-05*hvp_mobility*hvp_mobility+-1.39642e-03*hvp_mobility+-2.68140e-03'
+ sky130_fd_pr__pfet_g5v0d16v0__u0_diff_1 = '-4.75450e-05*hvp_mobility*hvp_mobility+-1.27673e-03*hvp_mobility+-9.22380e-04'
+ sky130_fd_pr__pfet_g5v0d16v0__vth0_diff_0 = '-3.50000e-05*hvp_threshold*hvp_threshold+-2.57500e-02*hvp_threshold+-3.14400e-02'
+ sky130_fd_pr__pfet_g5v0d16v0__vth0_diff_1 = '-7.37500e-06*hvp_threshold*hvp_threshold+-2.50735e-02*hvp_threshold+-5.85880e-02'
+ sky130_fd_pr__pfet_g5v0d16v0__wint_diff = '8.04375e-09*diff_cd'
+ rcl1 = '1.75000e-01*ic_res*ic_res+2.62500e+00*ic_res+9.30000e+00'
+ rcn = '1.59375e+00*ic_res_ndiff*ic_res_ndiff+3.43750e+01*ic_res_ndiff+1.82000e+02'
+ rcp = '6.75000e+01*ic_res_pdiff+6.00000e+02'
+ rcp1 = '-6.87500e-01*ic_res_poly*ic_res_poly+2.72500e+01*ic_res_poly+1.45280e+02'
+ rcrdlcon = '2.18750e-05*ic_res*ic_res+3.87500e-04*ic_res+5.80000e-03'
+ rcvia = '2.50000e-01*ic_res*ic_res+1.62500e+00*ic_res+4.50000e+00'
+ rcvia2 = '5.25000e-02*ic_res*ic_res+9.37500e-01*ic_res+3.41000e+00'
+ rcvia3 = '5.25000e-02*ic_res*ic_res+9.37500e-01*ic_res+3.41000e+00'
+ rcvia4 = '4.46875e-03*ic_res*ic_res+1.09875e-01*ic_res+3.80000e-01'
+ rdn = '3.00000e+00*ic_res_ndiff+1.20000e+02'
+ rdn_hv = '3.00000e+00*ic_res_ndiff+1.14000e+02'
+ rdp = '7.75000e+00*ic_res_pdiff+1.97000e+02'
+ rdp_hv = '7.75000e+00*ic_res_pdiff+1.91000e+02'
+ rl1 = '-3.12500e-03*ic_res*ic_res+6.62500e-01*ic_res+1.22000e+01'
+ rm1 = '5.00000e-03*ic_res+1.25000e-01'
+ rm2 = '5.00000e-03*ic_res+1.25000e-01'
+ rm3 = '2.25000e-03*ic_res+4.70000e-02'
+ rm4 = '2.25000e-03*ic_res+4.70000e-02'
+ rm5 = '-2.16840e-19*ic_res*ic_res+1.82500e-03*ic_res+2.85000e-02'
+ rnw = '1.15000e+02*ic_res+1.70000e+03'
+ rp1 = '5.00000e-02*ic_res_poly*ic_res_poly+1.70000e+00*ic_res_poly+4.82000e+01'
+ rrdl = '2.18750e-05*ic_res*ic_res+3.37500e-04*ic_res+5.00000e-03'
+ rspwres = '2.53250e+02*ic_res_pwell+3.81600e+03'
+ tol_li = '-5.00000e-09*ic_res'
+ tol_m1 = '-6.25000e-09*ic_res'
+ tol_m2 = '-6.25000e-09*ic_res'
+ tol_m3 = '-1.62500e-08*ic_res'
+ tol_m4 = '-1.62500e-08*ic_res'
+ tol_m5 = '-4.25000e-08*ic_res'
+ tol_nfom = '-1.72500e-08*ic_res'
+ tol_nw = '-1.72500e-08*ic_res'
+ tol_pfom = '-1.50000e-08*ic_res'
+ tol_poly = '-1.02500e-08*ic_res'
+ tol_rdl = '-2.50000e-07*ic_res'
+ sky130_fd_pr__cap_vpp_11p5x11p7_l1m1m2_noshield__cor = '3.30000e-02*ic_cap+1.00000e+00'
+ sky130_fd_pr__cap_vpp_11p5x11p7_m1m2m3m4_shieldl1m5__cor = '3.60000e-02*ic_cap+1.00000e+00'
+ sky130_fd_pr__cap_vpp_11p5x11p7_m1m2_shieldl1__cor = '3.30000e-02*ic_cap+1.00000e+00'
+ sky130_fd_pr__cap_vpp_11p5x11p7_m1m2m3_shieldl1__cor = '3.62500e-02*ic_cap+1.00000e+00'
+ sky130_fd_pr__cap_vpp_11p5x11p7_l1m1m2_shieldpom3__cor = '2.87500e-02*ic_cap+1.00000e+00'
+ sky130_fd_pr__cap_vpp_11p5x11p7_l1m1m2m3_shieldm4__cor = '5.00000e-02*ic_cap+1.00000e+00'
+ sky130_fd_pr__cap_vpp_11p5x11p7_l1m1m2m3m4_shieldm5__cor = '3.60000e-02*ic_cap+1.00000e+00'
+ sky130_fd_pr__cap_vpp_11p5x11p7_l1m1m2m3m4_shieldpom5__cor = '3.60000e-02*ic_cap+1.00000e+00'
+ sky130_fd_pr__cap_vpp_01p8x01p8_m1m2_noshield__cor = '5.35000e-02*ic_cap+1.00000e+00'
+ sky130_fd_pr__cap_vpp_03p9x03p9_m1m2_shieldl1_floatm3__cor = '-4.37500e-04*ic_cap*ic_cap+3.25000e-02*ic_cap+1.00000e+00'
+ sky130_fd_pr__cap_vpp_04p4x04p6_l1m1m2_noshield__cor = '5.10000e-02*ic_cap+1.00000e+00'
+ sky130_fd_pr__cap_vpp_04p4x04p6_m1m2_shieldl1__cor = '5.10000e-02*ic_cap+1.00000e+00'
+ sky130_fd_pr__cap_vpp_04p4x04p6_m1m2m3_shieldl1__cor = '5.62500e-02*ic_cap+1.00000e+00'
+ sky130_fd_pr__cap_vpp_04p4x04p6_l1m1m2_shieldpo_floatm3__cor = '4.60000e-02*ic_cap+1.00000e+00'
+ sky130_fd_pr__cap_vpp_06p8x06p1_l1m1m2_noshield__cor = '5.00000e-02*ic_cap+1.00000e+00'
+ sky130_fd_pr__cap_vpp_08p6x07p8_l1m1m2_noshield__cor = '4.32500e-02*ic_cap+1.00000e+00'
+ sky130_fd_pr__cap_vpp_08p6x07p8_m1m2_shieldl1__cor = '4.32500e-02*ic_cap+1.00000e+00'
+ sky130_fd_pr__cap_vpp_08p6x07p8_m1m2m3_shieldl1m5_floatm4__cor = '5.20000e-02*ic_cap+1.00000e+00'
+ sky130_fd_pr__cap_vpp_08p6x07p8_m1m2m3_shieldl1__cor = '4.75000e-02*ic_cap+1.00000e+00'
+ sky130_fd_pr__cap_vpp_08p6x07p8_l1m1m2_shieldpo_floatm3__cor = '3.85000e-02*ic_cap+1.00000e+00'
+ sky130_fd_pr__model__cap_vpp_finger__cor = '5.00000e-02*ic_cap+1.00000e+00'
+ sky130_fd_pr__cap_vpp_11p5x11p7_pol1m1m2m3m4m5_noshield_base__cor = '5.00000e-02*ic_cap+1.00000e+00'
.include "../parasitics/sky130_fd_pr__model__parasitic__diode_ps2dn.model.spice"
.include "../../../libs.ref/sky130_fd_pr/spice/sky130_fd_pr__pfet_g5v0d16v0__parasitic__diode_pw2dn.model.spice"
.include "../parasitics/sky130_fd_pr__model__parasitic__diode_pw2dn.model.spice"
.include "../../../libs.ref/sky130_fd_pr/spice/sky130_fd_pr__special_nfet_pass_flash.pm3.spice"
.include "../sky130_fd_pr__model__linear.model.spice"
.include "../../../libs.ref/sky130_fd_pr/spice/sky130_fd_pr__diode_pw2nd_05v5.model.spice"
.include "../../../libs.ref/sky130_fd_pr/spice/sky130_fd_pr__diode_pw2nd_11v0.model.spice"
.include "../../../libs.ref/sky130_fd_pr/spice/sky130_fd_pr__diode_pw2nd_05v5_lvt.model.spice"
.include "../../../libs.ref/sky130_fd_pr/spice/sky130_fd_pr__diode_pw2nd_05v5_nvt.model.spice"
.include "../../../libs.ref/sky130_fd_pr/spice/sky130_fd_pr__nfet_g5v0d10v5.pm3.spice"
.include "../../../libs.ref/sky130_fd_pr/spice/sky130_fd_pr__esd_nfet_g5v0d10v5.pm3.spice"
.include "../../../libs.ref/sky130_fd_pr/spice/sky130_fd_pr__nfet_05v0_nvt.pm3.spice"
.include "../../../libs.ref/sky130_fd_pr/spice/sky130_fd_pr__nfet_01v8_lvt.pm3.spice"
.include "../../../libs.ref/sky130_fd_pr/spice/sky130_fd_pr__special_nfet_pass_lvt.pm3.spice"
.include "../../../libs.ref/sky130_fd_pr/spice/sky130_fd_pr__special_nfet_pass.pm3.spice"
.include "../../../libs.ref/sky130_fd_pr/spice/sky130_fd_pr__special_nfet_latch.pm3.spice"
.include "../../../libs.ref/sky130_fd_pr/spice/sky130_fd_pr__npn_05v5_W1p00L1p00.model.spice"
.include "../../../libs.ref/sky130_fd_pr/spice/sky130_fd_pr__npn_05v5_W1p00L2p00.model.spice"
.include "../../../libs.ref/sky130_fd_pr/spice/sky130_fd_pr__npn_11v0_W1p00L1p00.model.spice"
.include "../../../libs.ref/sky130_fd_pr/spice/sky130_fd_pr__nfet_01v8.pm3.spice"
.include "../../../libs.ref/sky130_fd_pr/spice/sky130_fd_pr__esd_nfet_01v8.pm3.spice"
.include "../../../libs.ref/sky130_fd_pr/spice/sky130_fd_pr__nfet_03v3_nvt.pm3.spice"
.include "../../../libs.ref/sky130_fd_pr/spice/sky130_fd_pr__nfet_g5v0d16v0.pm3.spice"
.include "../../../libs.ref/sky130_fd_pr/spice/sky130_fd_pr__nfet_g5v0d16v0__subcircuit.pm3.spice"
.include "../parasitics/sky130_fd_pr__model__parasitic__diode_ps2nw.model.spice"
.include "../../../libs.ref/sky130_fd_pr/spice/sky130_fd_pr__diode_pd2nw_05v5.model.spice"
.include "../../../libs.ref/sky130_fd_pr/spice/sky130_fd_pr__diode_pd2nw_11v0.model.spice"
.include "../../../libs.ref/sky130_fd_pr/spice/sky130_fd_pr__diode_pd2nw_05v5_hvt.model.spice"
.include "../../../libs.ref/sky130_fd_pr/spice/sky130_fd_pr__diode_pd2nw_05v5_lvt.model.spice"
.include "../../../libs.ref/sky130_fd_pr/spice/sky130_fd_pr__pfet_01v8_hvt.pm3.spice"
.include "../../../libs.ref/sky130_fd_pr/spice/sky130_fd_pr__pfet_g5v0d10v5.pm3.spice"
.include "../../../libs.ref/sky130_fd_pr/spice/sky130_fd_pr__esd_pfet_g5v0d10v5.pm3.spice"
.include "../../../libs.ref/sky130_fd_pr/spice/sky130_fd_pr__pfet_01v8_lvt.pm3.spice"
.include "../../../libs.ref/sky130_fd_pr/spice/sky130_fd_pr__pnp_05v5_W3p40L3p40.model.spice"
.include "../../../libs.ref/sky130_fd_pr/spice/sky130_fd_pr__pnp_05v5_W0p68L0p68.model.spice"
.include "../../../libs.ref/sky130_fd_pr/spice/sky130_fd_pr__special_pfet_pass.pm3.spice"
.include "../../../libs.ref/sky130_fd_pr/spice/sky130_fd_pr__pfet_01v8.pm3.spice"
.include "../../../libs.ref/sky130_fd_pr/spice/sky130_fd_pr__pfet_g5v0d16v0.pm3.spice"
.include "../../../libs.ref/sky130_fd_pr/spice/sky130_fd_pr__pfet_g5v0d16v0__subcircuit.pm3.spice"
.include "../sonos_e/begin_of_life.pm3.spice"
.include "../sonos_p/begin_of_life.pm3.spice"
.include "../../../libs.ref/sky130_fd_pr/spice/sky130_fd_pr__cap_vpp_08p6x07p8_l1m1m2_noshield_o1.model.spice"
.include "../capacitors/sky130_fd_pr__model__cap_vpp_only_mos.model.spice"
.include "../capacitors/sky130_fd_pr__model__cap_vpp_only_p.model.spice"
.include "../capacitors/sky130_fd_pr__model__cap_vpp_only_pq.model.spice"
.include "../../../libs.ref/sky130_fd_pr/spice/sky130_fd_pr__cap_var_hvt.model.spice"
.include "../../../libs.ref/sky130_fd_pr/spice/sky130_fd_pr__cap_var_lvt.model.spice"
.include "../../../libs.ref/sky130_fd_pr/spice/sky130_fd_pr__res_iso_pw.model.spice"
.include "../capacitors/sky130_fd_pr__model__cap_mim.model.spice"
.include "../../../libs.ref/sky130_fd_pr/spice/sky130_fd_pr__rf_nfet_g5v0d10v5.pm3.spice"
.include "../../../libs.ref/sky130_fd_pr/spice/sky130_fd_pr__rf_nfet_g5v0d10v5_b.pm3.spice"
.include "../../../libs.ref/sky130_fd_pr/spice/sky130_fd_pr__rf_nfet_01v8_lvt.pm3.spice"
.include "../../../libs.ref/sky130_fd_pr/spice/sky130_fd_pr__rf_nfet_01v8_lvt_b.pm3.spice"
.include "../../../libs.ref/sky130_fd_pr/spice/sky130_fd_pr__rf_nfet_01v8.pm3.spice"
.include "../../../libs.ref/sky130_fd_pr/spice/sky130_fd_pr__rf_nfet_01v8_b.pm3.spice"
.include "../../../libs.ref/sky130_fd_pr/spice/sky130_fd_pr__pfet_01v8_mvt.pm3.spice"
.include "../../../libs.ref/sky130_fd_pr/spice/sky130_fd_pr__rf_pfet_01v8_mvt.pm3.spice"
.include "../../../libs.ref/sky130_fd_pr/spice/sky130_fd_pr__rf_pfet_01v8.pm3.spice"
.include "../../../libs.ref/sky130_fd_pr/spice/sky130_fd_pr__rf_pfet_01v8_b.pm3.spice"
.include "../sky130_fd_pr__model__r+c.model.spice"
.include "../../../libs.ref/sky130_fd_pr/spice/sky130_fd_pr__nfet_20v0_nvt__subcircuit.pm3.spice"
.include "../../../libs.ref/sky130_fd_pr/spice/sky130_fd_pr__nfet_20v0_nvt_iso__subcircuit.pm3.spice"
.include "../../../libs.ref/sky130_fd_pr/spice/sky130_fd_pr__nfet_20v0__subcircuit.pm3.spice"
.include "../../../libs.ref/sky130_fd_pr/spice/sky130_fd_pr__nfet_20v0_iso__subcircuit.pm3.spice"
.include "../../../libs.ref/sky130_fd_pr/spice/sky130_fd_pr__nfet_20v0_zvt__subcircuit.pm3.spice"
.include "../../../libs.ref/sky130_fd_pr/spice/sky130_fd_pr__pfet_20v0__subcircuit.pm3.spice"
