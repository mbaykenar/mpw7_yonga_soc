magic
tech sky130B
magscale 1 2
timestamp 1649977179
<< nwell >>
rect -38 261 2246 582
<< pwell >>
rect 273 157 457 201
rect 1572 181 2198 203
rect 1386 157 2198 181
rect 1 21 2198 157
rect 29 -17 63 21
<< scnmos >>
rect 79 47 109 131
rect 163 47 193 131
rect 351 47 381 175
rect 446 47 476 119
rect 556 47 586 119
rect 652 47 682 131
rect 766 47 796 131
rect 838 47 868 131
rect 1026 47 1056 131
rect 1098 47 1128 131
rect 1194 47 1224 131
rect 1266 47 1296 131
rect 1338 47 1368 131
rect 1462 47 1492 155
rect 1650 47 1680 177
rect 1734 47 1764 177
rect 1922 47 1952 177
rect 2006 47 2036 177
rect 2090 47 2120 177
<< scpmoshvt >>
rect 79 363 109 491
rect 163 363 193 491
rect 351 329 381 497
rect 448 413 478 497
rect 532 413 562 497
rect 652 413 682 497
rect 758 413 788 497
rect 842 413 872 497
rect 926 413 956 497
rect 998 413 1028 497
rect 1106 413 1136 497
rect 1178 413 1208 497
rect 1366 413 1396 497
rect 1462 329 1492 497
rect 1650 297 1680 497
rect 1734 297 1764 497
rect 1922 297 1952 497
rect 2006 297 2036 497
rect 2090 297 2120 497
<< ndiff >>
rect 27 119 79 131
rect 27 85 35 119
rect 69 85 79 119
rect 27 47 79 85
rect 109 93 163 131
rect 109 59 119 93
rect 153 59 163 93
rect 109 47 163 59
rect 193 119 245 131
rect 193 85 203 119
rect 237 85 245 119
rect 193 47 245 85
rect 299 93 351 175
rect 299 59 307 93
rect 341 59 351 93
rect 299 47 351 59
rect 381 119 431 175
rect 1598 165 1650 177
rect 1412 131 1462 155
rect 601 119 652 131
rect 381 111 446 119
rect 381 77 391 111
rect 425 77 446 111
rect 381 47 446 77
rect 476 93 556 119
rect 476 59 501 93
rect 535 59 556 93
rect 476 47 556 59
rect 586 47 652 119
rect 682 89 766 131
rect 682 55 722 89
rect 756 55 766 89
rect 682 47 766 55
rect 796 47 838 131
rect 868 109 920 131
rect 868 75 878 109
rect 912 75 920 109
rect 868 47 920 75
rect 974 93 1026 131
rect 974 59 982 93
rect 1016 59 1026 93
rect 974 47 1026 59
rect 1056 47 1098 131
rect 1128 95 1194 131
rect 1128 61 1144 95
rect 1178 61 1194 95
rect 1128 47 1194 61
rect 1224 47 1266 131
rect 1296 47 1338 131
rect 1368 113 1462 131
rect 1368 79 1398 113
rect 1432 79 1462 113
rect 1368 47 1462 79
rect 1492 120 1544 155
rect 1492 86 1502 120
rect 1536 86 1544 120
rect 1492 47 1544 86
rect 1598 131 1606 165
rect 1640 131 1650 165
rect 1598 97 1650 131
rect 1598 63 1606 97
rect 1640 63 1650 97
rect 1598 47 1650 63
rect 1680 165 1734 177
rect 1680 131 1690 165
rect 1724 131 1734 165
rect 1680 97 1734 131
rect 1680 63 1690 97
rect 1724 63 1734 97
rect 1680 47 1734 63
rect 1764 165 1816 177
rect 1764 131 1774 165
rect 1808 131 1816 165
rect 1764 97 1816 131
rect 1764 63 1774 97
rect 1808 63 1816 97
rect 1764 47 1816 63
rect 1870 119 1922 177
rect 1870 85 1878 119
rect 1912 85 1922 119
rect 1870 47 1922 85
rect 1952 161 2006 177
rect 1952 127 1962 161
rect 1996 127 2006 161
rect 1952 93 2006 127
rect 1952 59 1962 93
rect 1996 59 2006 93
rect 1952 47 2006 59
rect 2036 129 2090 177
rect 2036 95 2046 129
rect 2080 95 2090 129
rect 2036 47 2090 95
rect 2120 94 2172 177
rect 2120 60 2130 94
rect 2164 60 2172 94
rect 2120 47 2172 60
<< pdiff >>
rect 27 477 79 491
rect 27 443 35 477
rect 69 443 79 477
rect 27 409 79 443
rect 27 375 35 409
rect 69 375 79 409
rect 27 363 79 375
rect 109 461 163 491
rect 109 427 119 461
rect 153 427 163 461
rect 109 363 163 427
rect 193 477 245 491
rect 193 443 203 477
rect 237 443 245 477
rect 193 409 245 443
rect 193 375 203 409
rect 237 375 245 409
rect 193 363 245 375
rect 299 461 351 497
rect 299 427 307 461
rect 341 427 351 461
rect 299 329 351 427
rect 381 477 448 497
rect 381 443 391 477
rect 425 443 448 477
rect 381 413 448 443
rect 478 484 532 497
rect 478 450 488 484
rect 522 450 532 484
rect 478 413 532 450
rect 562 413 652 497
rect 682 485 758 497
rect 682 451 702 485
rect 736 451 758 485
rect 682 413 758 451
rect 788 459 842 497
rect 788 425 798 459
rect 832 425 842 459
rect 788 413 842 425
rect 872 485 926 497
rect 872 451 882 485
rect 916 451 926 485
rect 872 413 926 451
rect 956 413 998 497
rect 1028 483 1106 497
rect 1028 449 1038 483
rect 1072 449 1106 483
rect 1028 413 1106 449
rect 1136 413 1178 497
rect 1208 485 1260 497
rect 1208 451 1218 485
rect 1252 451 1260 485
rect 1208 413 1260 451
rect 1314 459 1366 497
rect 1314 425 1322 459
rect 1356 425 1366 459
rect 1314 413 1366 425
rect 1396 459 1462 497
rect 1396 425 1418 459
rect 1452 425 1462 459
rect 1396 413 1462 425
rect 381 409 433 413
rect 381 375 391 409
rect 425 375 433 409
rect 381 329 433 375
rect 1411 329 1462 413
rect 1492 459 1544 497
rect 1492 425 1502 459
rect 1536 425 1544 459
rect 1492 391 1544 425
rect 1492 357 1502 391
rect 1536 357 1544 391
rect 1492 329 1544 357
rect 1598 485 1650 497
rect 1598 451 1606 485
rect 1640 451 1650 485
rect 1598 417 1650 451
rect 1598 383 1606 417
rect 1640 383 1650 417
rect 1598 349 1650 383
rect 1598 315 1606 349
rect 1640 315 1650 349
rect 1598 297 1650 315
rect 1680 485 1734 497
rect 1680 451 1690 485
rect 1724 451 1734 485
rect 1680 417 1734 451
rect 1680 383 1690 417
rect 1724 383 1734 417
rect 1680 349 1734 383
rect 1680 315 1690 349
rect 1724 315 1734 349
rect 1680 297 1734 315
rect 1764 485 1816 497
rect 1764 451 1774 485
rect 1808 451 1816 485
rect 1764 417 1816 451
rect 1764 383 1774 417
rect 1808 383 1816 417
rect 1764 349 1816 383
rect 1764 315 1774 349
rect 1808 315 1816 349
rect 1764 297 1816 315
rect 1870 485 1922 497
rect 1870 451 1878 485
rect 1912 451 1922 485
rect 1870 417 1922 451
rect 1870 383 1878 417
rect 1912 383 1922 417
rect 1870 349 1922 383
rect 1870 315 1878 349
rect 1912 315 1922 349
rect 1870 297 1922 315
rect 1952 485 2006 497
rect 1952 451 1962 485
rect 1996 451 2006 485
rect 1952 417 2006 451
rect 1952 383 1962 417
rect 1996 383 2006 417
rect 1952 349 2006 383
rect 1952 315 1962 349
rect 1996 315 2006 349
rect 1952 297 2006 315
rect 2036 485 2090 497
rect 2036 451 2046 485
rect 2080 451 2090 485
rect 2036 417 2090 451
rect 2036 383 2046 417
rect 2080 383 2090 417
rect 2036 349 2090 383
rect 2036 315 2046 349
rect 2080 315 2090 349
rect 2036 297 2090 315
rect 2120 485 2172 497
rect 2120 451 2130 485
rect 2164 451 2172 485
rect 2120 417 2172 451
rect 2120 383 2130 417
rect 2164 383 2172 417
rect 2120 297 2172 383
<< ndiffc >>
rect 35 85 69 119
rect 119 59 153 93
rect 203 85 237 119
rect 307 59 341 93
rect 391 77 425 111
rect 501 59 535 93
rect 722 55 756 89
rect 878 75 912 109
rect 982 59 1016 93
rect 1144 61 1178 95
rect 1398 79 1432 113
rect 1502 86 1536 120
rect 1606 131 1640 165
rect 1606 63 1640 97
rect 1690 131 1724 165
rect 1690 63 1724 97
rect 1774 131 1808 165
rect 1774 63 1808 97
rect 1878 85 1912 119
rect 1962 127 1996 161
rect 1962 59 1996 93
rect 2046 95 2080 129
rect 2130 60 2164 94
<< pdiffc >>
rect 35 443 69 477
rect 35 375 69 409
rect 119 427 153 461
rect 203 443 237 477
rect 203 375 237 409
rect 307 427 341 461
rect 391 443 425 477
rect 488 450 522 484
rect 702 451 736 485
rect 798 425 832 459
rect 882 451 916 485
rect 1038 449 1072 483
rect 1218 451 1252 485
rect 1322 425 1356 459
rect 1418 425 1452 459
rect 391 375 425 409
rect 1502 425 1536 459
rect 1502 357 1536 391
rect 1606 451 1640 485
rect 1606 383 1640 417
rect 1606 315 1640 349
rect 1690 451 1724 485
rect 1690 383 1724 417
rect 1690 315 1724 349
rect 1774 451 1808 485
rect 1774 383 1808 417
rect 1774 315 1808 349
rect 1878 451 1912 485
rect 1878 383 1912 417
rect 1878 315 1912 349
rect 1962 451 1996 485
rect 1962 383 1996 417
rect 1962 315 1996 349
rect 2046 451 2080 485
rect 2046 383 2080 417
rect 2046 315 2080 349
rect 2130 451 2164 485
rect 2130 383 2164 417
<< poly >>
rect 79 491 109 517
rect 163 491 193 517
rect 351 497 381 523
rect 448 497 478 523
rect 532 497 562 523
rect 652 497 682 523
rect 758 497 788 523
rect 842 497 872 523
rect 926 497 956 523
rect 998 497 1028 523
rect 1106 497 1136 523
rect 1178 497 1208 523
rect 1366 497 1396 523
rect 1462 497 1492 523
rect 1650 497 1680 523
rect 1734 497 1764 523
rect 1922 497 1952 523
rect 2006 497 2036 523
rect 2090 497 2120 523
rect 79 348 109 363
rect 46 318 109 348
rect 46 280 76 318
rect 22 264 76 280
rect 163 274 193 363
rect 22 230 32 264
rect 66 230 76 264
rect 22 214 76 230
rect 118 264 193 274
rect 351 267 381 329
rect 448 279 478 413
rect 532 375 562 413
rect 652 381 682 413
rect 520 365 586 375
rect 520 331 536 365
rect 570 331 586 365
rect 520 321 586 331
rect 652 365 716 381
rect 652 331 672 365
rect 706 331 716 365
rect 652 315 716 331
rect 118 230 134 264
rect 168 230 193 264
rect 118 220 193 230
rect 46 176 76 214
rect 46 146 109 176
rect 79 131 109 146
rect 163 131 193 220
rect 344 251 398 267
rect 344 217 354 251
rect 388 217 398 251
rect 448 249 586 279
rect 344 201 398 217
rect 556 219 586 249
rect 351 175 381 201
rect 446 191 514 207
rect 446 157 470 191
rect 504 157 514 191
rect 446 141 514 157
rect 556 203 610 219
rect 556 169 566 203
rect 600 169 610 203
rect 556 153 610 169
rect 446 119 476 141
rect 556 119 586 153
rect 652 131 682 315
rect 758 229 788 413
rect 842 313 872 413
rect 926 313 956 413
rect 998 375 1028 413
rect 998 365 1064 375
rect 998 331 1014 365
rect 1048 331 1064 365
rect 998 321 1064 331
rect 830 297 956 313
rect 830 263 840 297
rect 874 263 956 297
rect 1106 291 1136 413
rect 1094 279 1136 291
rect 830 247 956 263
rect 1034 269 1136 279
rect 728 213 788 229
rect 728 179 738 213
rect 772 193 788 213
rect 772 179 796 193
rect 728 163 796 179
rect 766 131 796 163
rect 838 183 868 247
rect 1034 235 1050 269
rect 1084 261 1136 269
rect 1178 365 1208 413
rect 1178 349 1246 365
rect 1178 315 1202 349
rect 1236 315 1246 349
rect 1366 337 1396 413
rect 1178 291 1246 315
rect 1362 307 1396 337
rect 1178 261 1296 291
rect 1084 235 1128 261
rect 1034 225 1128 235
rect 838 147 1056 183
rect 838 131 868 147
rect 1026 131 1056 147
rect 1098 131 1128 225
rect 1170 203 1224 219
rect 1170 169 1180 203
rect 1214 169 1224 203
rect 1170 153 1224 169
rect 1194 131 1224 153
rect 1266 131 1296 261
rect 1362 229 1392 307
rect 1462 285 1492 329
rect 1338 213 1392 229
rect 1434 269 1492 285
rect 1434 235 1444 269
rect 1478 259 1492 269
rect 1650 259 1680 297
rect 1734 259 1764 297
rect 1922 259 1952 297
rect 2006 265 2036 297
rect 2090 265 2120 297
rect 1478 235 1952 259
rect 1434 219 1952 235
rect 1338 179 1348 213
rect 1382 179 1392 213
rect 1338 163 1392 179
rect 1462 205 1952 219
rect 1338 131 1368 163
rect 1462 155 1492 205
rect 1650 177 1680 205
rect 1734 177 1764 205
rect 1922 177 1952 205
rect 1994 249 2120 265
rect 1994 215 2004 249
rect 2038 215 2120 249
rect 1994 199 2120 215
rect 2006 177 2036 199
rect 2090 177 2120 199
rect 79 21 109 47
rect 163 21 193 47
rect 351 21 381 47
rect 446 21 476 47
rect 556 21 586 47
rect 652 21 682 47
rect 766 21 796 47
rect 838 21 868 47
rect 1026 21 1056 47
rect 1098 21 1128 47
rect 1194 21 1224 47
rect 1266 21 1296 47
rect 1338 21 1368 47
rect 1462 21 1492 47
rect 1650 21 1680 47
rect 1734 21 1764 47
rect 1922 21 1952 47
rect 2006 21 2036 47
rect 2090 21 2120 47
<< polycont >>
rect 32 230 66 264
rect 536 331 570 365
rect 672 331 706 365
rect 134 230 168 264
rect 354 217 388 251
rect 470 157 504 191
rect 566 169 600 203
rect 1014 331 1048 365
rect 840 263 874 297
rect 738 179 772 213
rect 1050 235 1084 269
rect 1202 315 1236 349
rect 1180 169 1214 203
rect 1444 235 1478 269
rect 1348 179 1382 213
rect 2004 215 2038 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2053 561
rect 2087 527 2145 561
rect 2179 527 2208 561
rect 35 477 69 493
rect 35 409 69 443
rect 103 461 169 527
rect 103 427 119 461
rect 153 427 169 461
rect 203 477 248 493
rect 237 443 248 477
rect 203 409 248 443
rect 291 461 357 527
rect 291 427 307 461
rect 341 427 357 461
rect 391 477 425 493
rect 686 485 762 527
rect 472 450 488 484
rect 522 450 638 484
rect 686 451 702 485
rect 736 451 762 485
rect 866 485 932 527
rect 798 459 832 475
rect 69 391 168 393
rect 69 375 129 391
rect 35 359 129 375
rect 122 357 129 359
rect 163 357 168 391
rect 18 264 88 325
rect 18 230 32 264
rect 66 230 88 264
rect 18 195 88 230
rect 122 264 168 357
rect 122 230 134 264
rect 122 161 168 230
rect 35 127 168 161
rect 237 375 248 409
rect 391 409 425 443
rect 203 187 248 375
rect 203 153 213 187
rect 247 153 248 187
rect 35 119 69 127
rect 203 119 248 153
rect 286 375 391 393
rect 286 359 425 375
rect 286 165 320 359
rect 470 357 489 391
rect 523 365 570 391
rect 523 357 536 365
rect 470 331 536 357
rect 354 251 436 325
rect 388 217 436 251
rect 354 201 436 217
rect 470 315 570 331
rect 470 191 514 315
rect 604 281 638 450
rect 866 451 882 485
rect 916 451 932 485
rect 1186 485 1268 527
rect 1022 449 1038 483
rect 1072 449 1152 483
rect 1186 451 1218 485
rect 1252 451 1268 485
rect 1308 459 1356 475
rect 1022 433 1152 449
rect 798 417 832 425
rect 1118 417 1152 433
rect 1308 425 1322 459
rect 1308 417 1356 425
rect 672 367 942 417
rect 672 365 722 367
rect 706 331 722 365
rect 672 315 722 331
rect 824 297 874 313
rect 824 281 840 297
rect 604 263 840 281
rect 604 247 874 263
rect 604 239 688 247
rect 286 127 425 165
rect 504 157 514 191
rect 470 141 514 157
rect 550 169 566 203
rect 600 187 620 203
rect 550 153 581 169
rect 615 153 620 187
rect 550 129 620 153
rect 35 69 69 85
rect 103 59 119 93
rect 153 59 169 93
rect 237 85 248 119
rect 391 111 425 127
rect 203 69 248 85
rect 103 17 169 59
rect 291 59 307 93
rect 341 59 357 93
rect 654 93 688 239
rect 908 213 942 367
rect 722 179 738 213
rect 772 187 804 213
rect 722 153 765 179
rect 799 153 804 187
rect 722 147 804 153
rect 862 145 942 213
rect 980 391 1080 393
rect 980 365 1041 391
rect 980 179 1014 365
rect 1075 357 1080 391
rect 1048 331 1080 357
rect 1118 383 1356 417
rect 1402 459 1468 527
rect 1604 485 1640 527
rect 1402 425 1418 459
rect 1452 425 1468 459
rect 1402 389 1468 425
rect 1502 459 1536 475
rect 1502 391 1536 425
rect 1048 269 1084 295
rect 1048 255 1050 269
rect 1048 221 1049 255
rect 1118 281 1152 383
rect 1502 353 1536 357
rect 1604 451 1606 485
rect 1604 417 1640 451
rect 1604 383 1606 417
rect 1502 349 1566 353
rect 1186 315 1202 349
rect 1236 315 1566 349
rect 1118 269 1494 281
rect 1118 247 1444 269
rect 1083 221 1084 235
rect 1048 213 1084 221
rect 1164 179 1180 203
rect 980 169 1180 179
rect 1214 169 1230 203
rect 980 145 1230 169
rect 862 109 912 145
rect 391 61 425 77
rect 291 17 357 59
rect 485 59 501 93
rect 535 59 688 93
rect 485 53 688 59
rect 722 89 804 105
rect 756 55 804 89
rect 862 75 878 109
rect 862 59 912 75
rect 948 93 1016 109
rect 1264 95 1298 247
rect 1428 235 1444 247
rect 1478 235 1494 269
rect 1332 179 1348 213
rect 1382 201 1398 213
rect 1382 187 1464 201
rect 1382 179 1409 187
rect 1332 153 1409 179
rect 1443 153 1464 187
rect 1332 147 1464 153
rect 1528 136 1566 315
rect 1604 349 1640 383
rect 1604 315 1606 349
rect 1604 296 1640 315
rect 1674 485 1740 493
rect 1674 451 1690 485
rect 1724 451 1740 485
rect 1674 417 1740 451
rect 1674 383 1690 417
rect 1724 383 1740 417
rect 1674 349 1740 383
rect 1674 315 1690 349
rect 1724 315 1740 349
rect 1502 120 1566 136
rect 948 59 982 93
rect 1128 61 1144 95
rect 1178 61 1298 95
rect 1334 79 1398 113
rect 1432 79 1466 113
rect 722 17 804 55
rect 948 17 1016 59
rect 1334 17 1466 79
rect 1536 86 1566 120
rect 1502 70 1566 86
rect 1604 165 1640 181
rect 1604 131 1606 165
rect 1604 97 1640 131
rect 1604 63 1606 97
rect 1604 17 1640 63
rect 1674 165 1740 315
rect 1774 485 1824 527
rect 1808 451 1824 485
rect 1774 417 1824 451
rect 1808 383 1824 417
rect 1774 349 1824 383
rect 1808 315 1824 349
rect 1774 296 1824 315
rect 1862 485 1928 493
rect 1862 451 1878 485
rect 1912 451 1928 485
rect 1862 417 1928 451
rect 1862 383 1878 417
rect 1912 383 1928 417
rect 1862 349 1928 383
rect 1862 315 1878 349
rect 1912 315 1928 349
rect 1862 265 1928 315
rect 1962 485 1996 527
rect 1962 417 1996 451
rect 1962 349 1996 383
rect 1962 299 1996 315
rect 2030 485 2096 493
rect 2030 451 2046 485
rect 2080 451 2096 485
rect 2030 417 2096 451
rect 2030 383 2046 417
rect 2080 383 2096 417
rect 2030 349 2096 383
rect 2130 485 2183 527
rect 2164 451 2183 485
rect 2130 417 2183 451
rect 2164 383 2183 417
rect 2130 367 2183 383
rect 2030 315 2046 349
rect 2080 333 2096 349
rect 2080 315 2183 333
rect 2030 299 2183 315
rect 1862 249 2038 265
rect 1862 215 2004 249
rect 1862 199 2038 215
rect 1674 131 1690 165
rect 1724 131 1740 165
rect 1674 97 1740 131
rect 1674 63 1690 97
rect 1724 63 1740 97
rect 1674 51 1740 63
rect 1774 165 1824 181
rect 1808 131 1824 165
rect 1774 97 1824 131
rect 1808 63 1824 97
rect 1774 17 1824 63
rect 1862 119 1912 199
rect 2072 169 2183 299
rect 2069 165 2183 169
rect 1862 85 1878 119
rect 1862 51 1912 85
rect 1946 161 2012 165
rect 1946 127 1962 161
rect 1996 127 2012 161
rect 1946 93 2012 127
rect 1946 59 1962 93
rect 1996 59 2012 93
rect 1946 17 2012 59
rect 2046 144 2183 165
rect 2046 129 2096 144
rect 2080 95 2096 129
rect 2046 51 2096 95
rect 2130 94 2183 110
rect 2164 60 2183 94
rect 2130 17 2183 60
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2053 17
rect 2087 -17 2145 17
rect 2179 -17 2208 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 1593 527 1627 561
rect 1685 527 1719 561
rect 1777 527 1811 561
rect 1869 527 1903 561
rect 1961 527 1995 561
rect 2053 527 2087 561
rect 2145 527 2179 561
rect 129 357 163 391
rect 213 153 247 187
rect 489 357 523 391
rect 581 169 600 187
rect 600 169 615 187
rect 581 153 615 169
rect 765 179 772 187
rect 772 179 799 187
rect 765 153 799 179
rect 1041 365 1075 391
rect 1041 357 1048 365
rect 1048 357 1075 365
rect 1049 235 1050 255
rect 1050 235 1083 255
rect 1049 221 1083 235
rect 1409 153 1443 187
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1593 -17 1627 17
rect 1685 -17 1719 17
rect 1777 -17 1811 17
rect 1869 -17 1903 17
rect 1961 -17 1995 17
rect 2053 -17 2087 17
rect 2145 -17 2179 17
<< metal1 >>
rect 0 561 2208 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2053 561
rect 2087 527 2145 561
rect 2179 527 2208 561
rect 0 496 2208 527
rect 117 391 175 397
rect 117 357 129 391
rect 163 388 175 391
rect 477 391 535 397
rect 477 388 489 391
rect 163 360 489 388
rect 163 357 175 360
rect 117 351 175 357
rect 477 357 489 360
rect 523 388 535 391
rect 1029 391 1087 397
rect 1029 388 1041 391
rect 523 360 1041 388
rect 523 357 535 360
rect 477 351 535 357
rect 1029 357 1041 360
rect 1075 357 1087 391
rect 1029 351 1087 357
rect 1037 255 1095 261
rect 1037 252 1049 255
rect 584 224 1049 252
rect 584 193 627 224
rect 1037 221 1049 224
rect 1083 221 1095 255
rect 1037 215 1095 221
rect 201 187 259 193
rect 201 153 213 187
rect 247 184 259 187
rect 569 187 627 193
rect 569 184 581 187
rect 247 156 581 184
rect 247 153 259 156
rect 201 147 259 153
rect 569 153 581 156
rect 615 153 627 187
rect 569 147 627 153
rect 753 187 811 193
rect 753 153 765 187
rect 799 184 811 187
rect 1397 187 1455 193
rect 1397 184 1409 187
rect 799 156 1409 184
rect 799 153 811 156
rect 753 147 811 153
rect 1397 153 1409 156
rect 1443 153 1455 187
rect 1397 147 1455 153
rect 0 17 2208 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2053 17
rect 2087 -17 2145 17
rect 2179 -17 2208 17
rect 0 -48 2208 -17
<< labels >>
flabel locali s 2145 221 2179 255 0 FreeSans 400 0 0 0 Q
port 8 nsew signal output
flabel locali s 1685 85 1719 119 0 FreeSans 400 0 0 0 Q_N
port 9 nsew signal output
flabel locali s 1685 153 1719 187 0 FreeSans 400 0 0 0 Q_N
port 9 nsew signal output
flabel locali s 1685 221 1719 255 0 FreeSans 400 0 0 0 Q_N
port 9 nsew signal output
flabel locali s 1685 289 1719 323 0 FreeSans 400 0 0 0 Q_N
port 9 nsew signal output
flabel locali s 1685 357 1719 391 0 FreeSans 400 0 0 0 Q_N
port 9 nsew signal output
flabel locali s 1685 425 1719 459 0 FreeSans 400 0 0 0 Q_N
port 9 nsew signal output
flabel locali s 397 289 431 323 0 FreeSans 200 0 0 0 D
port 2 nsew signal input
flabel locali s 397 221 431 255 0 FreeSans 200 0 0 0 D
port 2 nsew signal input
flabel locali s 29 527 63 561 3 FreeSans 400 0 0 0 VPWR
port 7 nsew power bidirectional abutment
flabel locali s 2053 425 2087 459 0 FreeSans 400 0 0 0 Q
port 8 nsew signal output
flabel locali s 2053 357 2087 391 0 FreeSans 400 0 0 0 Q
port 8 nsew signal output
flabel locali s 2053 85 2087 119 0 FreeSans 400 0 0 0 Q
port 8 nsew signal output
flabel locali s 765 153 799 187 0 FreeSans 400 0 0 0 SET_B
port 3 nsew signal input
flabel locali s 29 289 63 323 0 FreeSans 400 0 0 0 CLK
port 1 nsew clock input
flabel locali s 29 221 63 255 0 FreeSans 400 0 0 0 CLK
port 1 nsew clock input
flabel locali s 29 -17 63 17 3 FreeSans 400 0 0 0 VGND
port 4 nsew ground bidirectional abutment
flabel nwell s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 6 nsew power bidirectional
flabel nwell s 46 544 46 544 0 FreeSans 200 0 0 0 VPB
port 6 nsew
flabel nwell s 46 544 46 544 3 FreeSans 400 0 0 0 VPB
port 6 nsew
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 5 nsew ground bidirectional
flabel pwell s 46 0 46 0 0 FreeSans 200 0 0 0 VNB
port 5 nsew
flabel pwell s 46 0 46 0 3 FreeSans 400 0 0 0 VNB
port 5 nsew
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 4 nsew ground bidirectional abutment
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 7 nsew power bidirectional abutment
flabel metal1 s 46 544 46 544 0 FreeSans 200 0 0 0 VPWR
port 7 nsew
flabel metal1 s 46 0 46 0 0 FreeSans 200 0 0 0 VGND
port 4 nsew
rlabel comment s 0 0 0 0 4 dfsbp_2
rlabel locali s 1332 201 1398 213 1 SET_B
port 3 nsew signal input
rlabel locali s 1332 147 1464 201 1 SET_B
port 3 nsew signal input
rlabel metal1 s 1397 184 1455 193 1 SET_B
port 3 nsew signal input
rlabel metal1 s 1397 147 1455 156 1 SET_B
port 3 nsew signal input
rlabel metal1 s 753 184 811 193 1 SET_B
port 3 nsew signal input
rlabel metal1 s 753 156 1455 184 1 SET_B
port 3 nsew signal input
rlabel metal1 s 753 147 811 156 1 SET_B
port 3 nsew signal input
rlabel metal1 s 0 -48 2208 48 1 VGND
port 4 nsew ground bidirectional abutment
rlabel metal1 s 0 496 2208 592 1 VPWR
port 7 nsew power bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 2208 544
string GDS_END 2515242
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 2496374
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
<< end >>
