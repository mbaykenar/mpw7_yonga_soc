magic
tech sky130A
timestamp 1649977179
<< properties >>
string GDS_END 39460950
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 39455122
<< end >>
