magic
tech sky130B
magscale 12 1
timestamp 1598786878
<< metal5 >>
rect 0 0 30 30
<< properties >>
string FIXED_BBOX 0 -30 45 105
<< end >>
