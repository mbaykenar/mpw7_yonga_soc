magic
tech sky130B
magscale 1 2
timestamp 1649977179
<< nwell >>
rect -38 261 774 582
<< pwell >>
rect 98 157 717 203
rect 1 67 717 157
rect 1 21 191 67
rect 405 21 717 67
rect 30 -17 64 21
<< scnmos >>
rect 79 47 109 131
rect 180 93 210 177
rect 501 47 531 177
rect 573 47 603 177
<< scpmoshvt >>
rect 79 369 109 497
rect 163 369 193 497
rect 353 297 383 497
rect 573 297 603 497
<< ndiff >>
rect 124 131 180 177
rect 27 106 79 131
rect 27 72 35 106
rect 69 72 79 106
rect 27 47 79 72
rect 109 93 180 131
rect 210 169 333 177
rect 210 135 287 169
rect 321 135 333 169
rect 210 93 333 135
rect 431 93 501 177
rect 109 89 165 93
rect 109 55 119 89
rect 153 55 165 89
rect 109 47 165 55
rect 431 59 439 93
rect 473 59 501 93
rect 431 47 501 59
rect 531 47 573 177
rect 603 157 691 177
rect 603 123 641 157
rect 675 123 691 157
rect 603 89 691 123
rect 603 55 641 89
rect 675 55 691 89
rect 603 47 691 55
<< pdiff >>
rect 27 461 79 497
rect 27 427 35 461
rect 69 427 79 461
rect 27 369 79 427
rect 109 489 163 497
rect 109 455 119 489
rect 153 455 163 489
rect 109 369 163 455
rect 193 470 245 497
rect 193 436 203 470
rect 237 436 245 470
rect 193 369 245 436
rect 299 469 353 497
rect 299 435 307 469
rect 341 435 353 469
rect 299 297 353 435
rect 383 297 573 497
rect 603 448 666 497
rect 603 414 624 448
rect 658 414 666 448
rect 603 380 666 414
rect 603 346 624 380
rect 658 346 666 380
rect 603 297 666 346
<< ndiffc >>
rect 35 72 69 106
rect 287 135 321 169
rect 119 55 153 89
rect 439 59 473 93
rect 641 123 675 157
rect 641 55 675 89
<< pdiffc >>
rect 35 427 69 461
rect 119 455 153 489
rect 203 436 237 470
rect 307 435 341 469
rect 624 414 658 448
rect 624 346 658 380
<< poly >>
rect 79 497 109 523
rect 163 497 193 523
rect 353 497 383 523
rect 573 497 603 523
rect 79 265 109 369
rect 27 249 109 265
rect 27 215 37 249
rect 71 215 109 249
rect 27 199 109 215
rect 163 265 193 369
rect 353 265 383 297
rect 573 265 603 297
rect 163 249 383 265
rect 163 215 198 249
rect 232 215 383 249
rect 163 199 383 215
rect 447 249 531 265
rect 447 215 457 249
rect 491 215 531 249
rect 447 199 531 215
rect 79 131 109 199
rect 180 177 210 199
rect 501 177 531 199
rect 573 249 627 265
rect 573 215 583 249
rect 617 215 627 249
rect 573 199 627 215
rect 573 177 603 199
rect 79 21 109 47
rect 180 39 210 93
rect 501 21 531 47
rect 573 21 603 47
<< polycont >>
rect 37 215 71 249
rect 198 215 232 249
rect 457 215 491 249
rect 583 215 617 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 736 561
rect 17 461 69 493
rect 17 427 35 461
rect 103 489 169 527
rect 103 455 119 489
rect 153 455 169 489
rect 103 435 169 455
rect 203 470 254 492
rect 237 436 254 470
rect 17 401 69 427
rect 203 401 254 436
rect 288 469 361 527
rect 288 435 307 469
rect 341 435 361 469
rect 395 448 719 493
rect 395 414 624 448
rect 658 414 719 448
rect 17 357 148 401
rect 203 360 361 401
rect 17 249 71 323
rect 17 215 37 249
rect 17 199 71 215
rect 105 165 148 357
rect 182 249 248 326
rect 182 215 198 249
rect 232 215 248 249
rect 282 265 361 360
rect 395 380 719 414
rect 395 346 624 380
rect 658 346 719 380
rect 395 299 719 346
rect 282 249 507 265
rect 282 215 457 249
rect 491 215 507 249
rect 541 249 617 265
rect 541 215 583 249
rect 282 177 337 215
rect 541 199 617 215
rect 541 181 591 199
rect 271 169 337 177
rect 17 123 237 165
rect 271 135 287 169
rect 321 135 337 169
rect 271 127 337 135
rect 371 147 591 181
rect 651 165 719 299
rect 625 157 719 165
rect 17 106 69 123
rect 17 72 35 106
rect 203 93 237 123
rect 371 93 405 147
rect 625 123 641 157
rect 675 123 719 157
rect 17 56 69 72
rect 103 55 119 89
rect 153 55 169 89
rect 103 17 169 55
rect 203 51 405 93
rect 439 93 591 113
rect 473 59 591 93
rect 439 17 591 59
rect 625 89 719 123
rect 625 55 641 89
rect 675 55 719 89
rect 625 51 719 55
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 736 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
<< metal1 >>
rect 0 561 736 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 736 561
rect 0 496 736 527
rect 0 17 736 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 736 17
rect 0 -48 736 -17
<< labels >>
rlabel comment s 0 0 0 0 4 ebufn_1
flabel locali s 582 357 616 391 0 FreeSans 200 0 0 0 Z
port 7 nsew signal output
flabel locali s 582 425 616 459 0 FreeSans 200 0 0 0 Z
port 7 nsew signal output
flabel locali s 674 425 708 459 0 FreeSans 200 0 0 0 Z
port 7 nsew signal output
flabel locali s 674 357 708 391 0 FreeSans 200 0 0 0 Z
port 7 nsew signal output
flabel locali s 674 289 708 323 0 FreeSans 200 0 0 0 Z
port 7 nsew signal output
flabel locali s 674 221 708 255 0 FreeSans 200 0 0 0 Z
port 7 nsew signal output
flabel locali s 214 221 248 255 0 FreeSans 200 0 0 0 TE_B
port 2 nsew signal input
flabel locali s 214 289 248 323 0 FreeSans 200 0 0 0 TE_B
port 2 nsew signal input
flabel locali s 30 289 64 323 0 FreeSans 200 0 0 0 A
port 1 nsew signal input
flabel locali s 30 221 64 255 0 FreeSans 200 0 0 0 A
port 1 nsew signal input
flabel locali s 490 357 524 391 0 FreeSans 200 0 0 0 Z
port 7 nsew signal output
flabel locali s 674 85 708 119 0 FreeSans 200 0 0 0 Z
port 7 nsew signal output
flabel locali s 674 153 708 187 0 FreeSans 200 0 0 0 Z
port 7 nsew signal output
flabel locali s 490 425 524 459 0 FreeSans 200 0 0 0 Z
port 7 nsew signal output
flabel locali s 398 425 432 459 0 FreeSans 200 0 0 0 Z
port 7 nsew signal output
flabel locali s 398 357 432 391 0 FreeSans 200 0 0 0 Z
port 7 nsew signal output
flabel pwell s 30 -17 64 17 0 FreeSans 200 0 0 0 VNB
port 4 nsew ground bidirectional
flabel nwell s 30 527 64 561 0 FreeSans 200 0 0 0 VPB
port 5 nsew power bidirectional
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 6 nsew power bidirectional abutment
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 3 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 736 48 1 VGND
port 3 nsew ground bidirectional abutment
rlabel metal1 s 0 496 736 592 1 VPWR
port 6 nsew power bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 736 544
string GDS_END 2924272
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 2917454
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string path 0.000 13.600 18.400 13.600 
<< end >>
