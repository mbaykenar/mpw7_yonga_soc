magic
tech sky130A
magscale 1 2
timestamp 1649977179
<< locali >>
rect 1935 9068 1969 9084
rect 1935 9018 1969 9034
rect 21903 9068 21937 9084
rect 21903 9018 21937 9034
rect 41871 9068 41905 9084
rect 41871 9018 41905 9034
rect 61839 9068 61873 9084
rect 61839 9018 61873 9034
<< viali >>
rect 1935 9034 1969 9068
rect 21903 9034 21937 9068
rect 41871 9034 41905 9068
rect 61839 9034 61873 9068
<< metal1 >>
rect 1923 9068 1981 9074
rect 1923 9034 1935 9068
rect 1969 9065 1981 9068
rect 20701 9065 20707 9077
rect 1969 9037 20707 9065
rect 1969 9034 1981 9037
rect 1923 9028 1981 9034
rect 20701 9025 20707 9037
rect 20759 9025 20765 9077
rect 21891 9068 21949 9074
rect 21891 9034 21903 9068
rect 21937 9065 21949 9068
rect 40669 9065 40675 9077
rect 21937 9037 40675 9065
rect 21937 9034 21949 9037
rect 21891 9028 21949 9034
rect 40669 9025 40675 9037
rect 40727 9025 40733 9077
rect 41859 9068 41917 9074
rect 41859 9034 41871 9068
rect 41905 9065 41917 9068
rect 60637 9065 60643 9077
rect 41905 9037 60643 9065
rect 41905 9034 41917 9037
rect 41859 9028 41917 9034
rect 60637 9025 60643 9037
rect 60695 9025 60701 9077
rect 61827 9068 61885 9074
rect 61827 9034 61839 9068
rect 61873 9065 61885 9068
rect 80605 9065 80611 9077
rect 61873 9037 80611 9065
rect 61873 9034 61885 9037
rect 61827 9028 61885 9034
rect 80605 9025 80611 9037
rect 80663 9025 80669 9077
rect 1629 8153 1689 8209
rect 4125 8153 4185 8209
rect 6621 8153 6681 8209
rect 9117 8153 9177 8209
rect 11613 8153 11673 8209
rect 14109 8153 14169 8209
rect 16605 8153 16665 8209
rect 19101 8153 19161 8209
rect 21597 8153 21657 8209
rect 24093 8153 24153 8209
rect 26589 8153 26649 8209
rect 29085 8153 29145 8209
rect 31581 8153 31641 8209
rect 34077 8153 34137 8209
rect 36573 8153 36633 8209
rect 39069 8153 39129 8209
rect 41565 8153 41625 8209
rect 44061 8153 44121 8209
rect 46557 8153 46617 8209
rect 49053 8153 49113 8209
rect 51549 8153 51609 8209
rect 54045 8153 54105 8209
rect 56541 8153 56601 8209
rect 59037 8153 59097 8209
rect 61533 8153 61593 8209
rect 64029 8153 64089 8209
rect 66525 8153 66585 8209
rect 69021 8153 69081 8209
rect 71517 8153 71577 8209
rect 74013 8153 74073 8209
rect 76509 8153 76569 8209
rect 79005 8153 79065 8209
rect 20701 8119 20707 8128
rect 1473 8085 20707 8119
rect 20701 8076 20707 8085
rect 20759 8119 20765 8128
rect 40669 8119 40675 8128
rect 20759 8085 20817 8119
rect 21441 8085 40675 8119
rect 20759 8076 20765 8085
rect 40669 8076 40675 8085
rect 40727 8119 40733 8128
rect 60637 8119 60643 8128
rect 40727 8085 40785 8119
rect 41409 8085 60643 8119
rect 40727 8076 40733 8085
rect 60637 8076 60643 8085
rect 60695 8119 60701 8128
rect 80605 8119 80611 8128
rect 60695 8085 60753 8119
rect 61377 8085 80611 8119
rect 60695 8076 60701 8085
rect 80605 8076 80611 8085
rect 80663 8119 80669 8128
rect 80663 8085 80721 8119
rect 80663 8076 80669 8085
rect 1501 6136 1529 6202
rect 1501 6108 1601 6136
rect 1478 5696 1524 5950
rect 1573 4820 1601 6108
rect 1703 6056 1731 6202
rect 3997 6136 4025 6202
rect 3997 6108 4097 6136
rect 1646 6028 1731 6056
rect 1646 4808 1674 6028
rect 3974 5696 4020 5950
rect 4069 4820 4097 6108
rect 4199 6056 4227 6202
rect 6493 6136 6521 6202
rect 6493 6108 6593 6136
rect 4142 6028 4227 6056
rect 4142 4808 4170 6028
rect 6470 5696 6516 5950
rect 6565 4820 6593 6108
rect 6695 6056 6723 6202
rect 8989 6136 9017 6202
rect 8989 6108 9089 6136
rect 6638 6028 6723 6056
rect 6638 4808 6666 6028
rect 8966 5696 9012 5950
rect 9061 4820 9089 6108
rect 9191 6056 9219 6202
rect 11485 6136 11513 6202
rect 11485 6108 11585 6136
rect 9134 6028 9219 6056
rect 9134 4808 9162 6028
rect 11462 5696 11508 5950
rect 11557 4820 11585 6108
rect 11687 6056 11715 6202
rect 13981 6136 14009 6202
rect 13981 6108 14081 6136
rect 11630 6028 11715 6056
rect 11630 4808 11658 6028
rect 13958 5696 14004 5950
rect 14053 4820 14081 6108
rect 14183 6056 14211 6202
rect 16477 6136 16505 6202
rect 16477 6108 16577 6136
rect 14126 6028 14211 6056
rect 14126 4808 14154 6028
rect 16454 5696 16500 5950
rect 16549 4820 16577 6108
rect 16679 6056 16707 6202
rect 18973 6136 19001 6202
rect 18973 6108 19073 6136
rect 16622 6028 16707 6056
rect 16622 4808 16650 6028
rect 18950 5696 18996 5950
rect 19045 4820 19073 6108
rect 19175 6056 19203 6202
rect 21469 6136 21497 6202
rect 21469 6108 21569 6136
rect 19118 6028 19203 6056
rect 19118 4808 19146 6028
rect 21446 5696 21492 5950
rect 21541 4820 21569 6108
rect 21671 6056 21699 6202
rect 23965 6136 23993 6202
rect 23965 6108 24065 6136
rect 21614 6028 21699 6056
rect 21614 4808 21642 6028
rect 23942 5696 23988 5950
rect 24037 4820 24065 6108
rect 24167 6056 24195 6202
rect 26461 6136 26489 6202
rect 26461 6108 26561 6136
rect 24110 6028 24195 6056
rect 24110 4808 24138 6028
rect 26438 5696 26484 5950
rect 26533 4820 26561 6108
rect 26663 6056 26691 6202
rect 28957 6136 28985 6202
rect 28957 6108 29057 6136
rect 26606 6028 26691 6056
rect 26606 4808 26634 6028
rect 28934 5696 28980 5950
rect 29029 4820 29057 6108
rect 29159 6056 29187 6202
rect 31453 6136 31481 6202
rect 31453 6108 31553 6136
rect 29102 6028 29187 6056
rect 29102 4808 29130 6028
rect 31430 5696 31476 5950
rect 31525 4820 31553 6108
rect 31655 6056 31683 6202
rect 33949 6136 33977 6202
rect 33949 6108 34049 6136
rect 31598 6028 31683 6056
rect 31598 4808 31626 6028
rect 33926 5696 33972 5950
rect 34021 4820 34049 6108
rect 34151 6056 34179 6202
rect 36445 6136 36473 6202
rect 36445 6108 36545 6136
rect 34094 6028 34179 6056
rect 34094 4808 34122 6028
rect 36422 5696 36468 5950
rect 36517 4820 36545 6108
rect 36647 6056 36675 6202
rect 38941 6136 38969 6202
rect 38941 6108 39041 6136
rect 36590 6028 36675 6056
rect 36590 4808 36618 6028
rect 38918 5696 38964 5950
rect 39013 4820 39041 6108
rect 39143 6056 39171 6202
rect 41437 6136 41465 6202
rect 41437 6108 41537 6136
rect 39086 6028 39171 6056
rect 39086 4808 39114 6028
rect 41414 5696 41460 5950
rect 41509 4820 41537 6108
rect 41639 6056 41667 6202
rect 43933 6136 43961 6202
rect 43933 6108 44033 6136
rect 41582 6028 41667 6056
rect 41582 4808 41610 6028
rect 43910 5696 43956 5950
rect 44005 4820 44033 6108
rect 44135 6056 44163 6202
rect 46429 6136 46457 6202
rect 46429 6108 46529 6136
rect 44078 6028 44163 6056
rect 44078 4808 44106 6028
rect 46406 5696 46452 5950
rect 46501 4820 46529 6108
rect 46631 6056 46659 6202
rect 48925 6136 48953 6202
rect 48925 6108 49025 6136
rect 46574 6028 46659 6056
rect 46574 4808 46602 6028
rect 48902 5696 48948 5950
rect 48997 4820 49025 6108
rect 49127 6056 49155 6202
rect 51421 6136 51449 6202
rect 51421 6108 51521 6136
rect 49070 6028 49155 6056
rect 49070 4808 49098 6028
rect 51398 5696 51444 5950
rect 51493 4820 51521 6108
rect 51623 6056 51651 6202
rect 53917 6136 53945 6202
rect 53917 6108 54017 6136
rect 51566 6028 51651 6056
rect 51566 4808 51594 6028
rect 53894 5696 53940 5950
rect 53989 4820 54017 6108
rect 54119 6056 54147 6202
rect 56413 6136 56441 6202
rect 56413 6108 56513 6136
rect 54062 6028 54147 6056
rect 54062 4808 54090 6028
rect 56390 5696 56436 5950
rect 56485 4820 56513 6108
rect 56615 6056 56643 6202
rect 58909 6136 58937 6202
rect 58909 6108 59009 6136
rect 56558 6028 56643 6056
rect 56558 4808 56586 6028
rect 58886 5696 58932 5950
rect 58981 4820 59009 6108
rect 59111 6056 59139 6202
rect 61405 6136 61433 6202
rect 61405 6108 61505 6136
rect 59054 6028 59139 6056
rect 59054 4808 59082 6028
rect 61382 5696 61428 5950
rect 61477 4820 61505 6108
rect 61607 6056 61635 6202
rect 63901 6136 63929 6202
rect 63901 6108 64001 6136
rect 61550 6028 61635 6056
rect 61550 4808 61578 6028
rect 63878 5696 63924 5950
rect 63973 4820 64001 6108
rect 64103 6056 64131 6202
rect 66397 6136 66425 6202
rect 66397 6108 66497 6136
rect 64046 6028 64131 6056
rect 64046 4808 64074 6028
rect 66374 5696 66420 5950
rect 66469 4820 66497 6108
rect 66599 6056 66627 6202
rect 68893 6136 68921 6202
rect 68893 6108 68993 6136
rect 66542 6028 66627 6056
rect 66542 4808 66570 6028
rect 68870 5696 68916 5950
rect 68965 4820 68993 6108
rect 69095 6056 69123 6202
rect 71389 6136 71417 6202
rect 71389 6108 71489 6136
rect 69038 6028 69123 6056
rect 69038 4808 69066 6028
rect 71366 5696 71412 5950
rect 71461 4820 71489 6108
rect 71591 6056 71619 6202
rect 73885 6136 73913 6202
rect 73885 6108 73985 6136
rect 71534 6028 71619 6056
rect 71534 4808 71562 6028
rect 73862 5696 73908 5950
rect 73957 4820 73985 6108
rect 74087 6056 74115 6202
rect 76381 6136 76409 6202
rect 76381 6108 76481 6136
rect 74030 6028 74115 6056
rect 74030 4808 74058 6028
rect 76358 5696 76404 5950
rect 76453 4820 76481 6108
rect 76583 6056 76611 6202
rect 78877 6136 78905 6202
rect 78877 6108 78977 6136
rect 76526 6028 76611 6056
rect 76526 4808 76554 6028
rect 78854 5696 78900 5950
rect 78949 4820 78977 6108
rect 79079 6056 79107 6202
rect 79022 6028 79107 6056
rect 79022 4808 79050 6028
rect 1573 3628 1601 3694
rect 1454 3600 1601 3628
rect 1454 3194 1482 3600
rect 1646 3548 1674 3694
rect 4069 3628 4097 3694
rect 3950 3600 4097 3628
rect 1646 3520 1946 3548
rect 1918 3318 1946 3520
rect 3950 3194 3978 3600
rect 4142 3548 4170 3694
rect 6565 3628 6593 3694
rect 6446 3600 6593 3628
rect 4142 3520 4442 3548
rect 4414 3318 4442 3520
rect 6446 3194 6474 3600
rect 6638 3548 6666 3694
rect 9061 3628 9089 3694
rect 8942 3600 9089 3628
rect 6638 3520 6938 3548
rect 6910 3318 6938 3520
rect 8942 3194 8970 3600
rect 9134 3548 9162 3694
rect 11557 3628 11585 3694
rect 11438 3600 11585 3628
rect 9134 3520 9434 3548
rect 9406 3318 9434 3520
rect 11438 3194 11466 3600
rect 11630 3548 11658 3694
rect 14053 3628 14081 3694
rect 13934 3600 14081 3628
rect 11630 3520 11930 3548
rect 11902 3318 11930 3520
rect 13934 3194 13962 3600
rect 14126 3548 14154 3694
rect 16549 3628 16577 3694
rect 16430 3600 16577 3628
rect 14126 3520 14426 3548
rect 14398 3318 14426 3520
rect 16430 3194 16458 3600
rect 16622 3548 16650 3694
rect 19045 3628 19073 3694
rect 18926 3600 19073 3628
rect 16622 3520 16922 3548
rect 16894 3318 16922 3520
rect 18926 3194 18954 3600
rect 19118 3548 19146 3694
rect 21541 3628 21569 3694
rect 21422 3600 21569 3628
rect 19118 3520 19418 3548
rect 19390 3318 19418 3520
rect 21422 3194 21450 3600
rect 21614 3548 21642 3694
rect 24037 3628 24065 3694
rect 23918 3600 24065 3628
rect 21614 3520 21914 3548
rect 21886 3318 21914 3520
rect 23918 3194 23946 3600
rect 24110 3548 24138 3694
rect 26533 3628 26561 3694
rect 26414 3600 26561 3628
rect 24110 3520 24410 3548
rect 24382 3318 24410 3520
rect 26414 3194 26442 3600
rect 26606 3548 26634 3694
rect 29029 3628 29057 3694
rect 28910 3600 29057 3628
rect 26606 3520 26906 3548
rect 26878 3318 26906 3520
rect 28910 3194 28938 3600
rect 29102 3548 29130 3694
rect 31525 3628 31553 3694
rect 31406 3600 31553 3628
rect 29102 3520 29402 3548
rect 29374 3318 29402 3520
rect 31406 3194 31434 3600
rect 31598 3548 31626 3694
rect 34021 3628 34049 3694
rect 33902 3600 34049 3628
rect 31598 3520 31898 3548
rect 31870 3318 31898 3520
rect 33902 3194 33930 3600
rect 34094 3548 34122 3694
rect 36517 3628 36545 3694
rect 36398 3600 36545 3628
rect 34094 3520 34394 3548
rect 34366 3318 34394 3520
rect 36398 3194 36426 3600
rect 36590 3548 36618 3694
rect 39013 3628 39041 3694
rect 38894 3600 39041 3628
rect 36590 3520 36890 3548
rect 36862 3318 36890 3520
rect 38894 3194 38922 3600
rect 39086 3548 39114 3694
rect 41509 3628 41537 3694
rect 41390 3600 41537 3628
rect 39086 3520 39386 3548
rect 39358 3318 39386 3520
rect 41390 3194 41418 3600
rect 41582 3548 41610 3694
rect 44005 3628 44033 3694
rect 43886 3600 44033 3628
rect 41582 3520 41882 3548
rect 41854 3318 41882 3520
rect 43886 3194 43914 3600
rect 44078 3548 44106 3694
rect 46501 3628 46529 3694
rect 46382 3600 46529 3628
rect 44078 3520 44378 3548
rect 44350 3318 44378 3520
rect 46382 3194 46410 3600
rect 46574 3548 46602 3694
rect 48997 3628 49025 3694
rect 48878 3600 49025 3628
rect 46574 3520 46874 3548
rect 46846 3318 46874 3520
rect 48878 3194 48906 3600
rect 49070 3548 49098 3694
rect 51493 3628 51521 3694
rect 51374 3600 51521 3628
rect 49070 3520 49370 3548
rect 49342 3318 49370 3520
rect 51374 3194 51402 3600
rect 51566 3548 51594 3694
rect 53989 3628 54017 3694
rect 53870 3600 54017 3628
rect 51566 3520 51866 3548
rect 51838 3318 51866 3520
rect 53870 3194 53898 3600
rect 54062 3548 54090 3694
rect 56485 3628 56513 3694
rect 56366 3600 56513 3628
rect 54062 3520 54362 3548
rect 54334 3318 54362 3520
rect 56366 3194 56394 3600
rect 56558 3548 56586 3694
rect 58981 3628 59009 3694
rect 58862 3600 59009 3628
rect 56558 3520 56858 3548
rect 56830 3318 56858 3520
rect 58862 3194 58890 3600
rect 59054 3548 59082 3694
rect 61477 3628 61505 3694
rect 61358 3600 61505 3628
rect 59054 3520 59354 3548
rect 59326 3318 59354 3520
rect 61358 3194 61386 3600
rect 61550 3548 61578 3694
rect 63973 3628 64001 3694
rect 63854 3600 64001 3628
rect 61550 3520 61850 3548
rect 61822 3318 61850 3520
rect 63854 3194 63882 3600
rect 64046 3548 64074 3694
rect 66469 3628 66497 3694
rect 66350 3600 66497 3628
rect 64046 3520 64346 3548
rect 64318 3318 64346 3520
rect 66350 3194 66378 3600
rect 66542 3548 66570 3694
rect 68965 3628 68993 3694
rect 68846 3600 68993 3628
rect 66542 3520 66842 3548
rect 66814 3318 66842 3520
rect 68846 3194 68874 3600
rect 69038 3548 69066 3694
rect 71461 3628 71489 3694
rect 71342 3600 71489 3628
rect 69038 3520 69338 3548
rect 69310 3318 69338 3520
rect 71342 3194 71370 3600
rect 71534 3548 71562 3694
rect 73957 3628 73985 3694
rect 73838 3600 73985 3628
rect 71534 3520 71834 3548
rect 71806 3318 71834 3520
rect 73838 3194 73866 3600
rect 74030 3548 74058 3694
rect 76453 3628 76481 3694
rect 76334 3600 76481 3628
rect 74030 3520 74330 3548
rect 74302 3318 74330 3520
rect 76334 3194 76362 3600
rect 76526 3548 76554 3694
rect 78949 3628 78977 3694
rect 78830 3600 78977 3628
rect 76526 3520 76826 3548
rect 76798 3318 76826 3520
rect 78830 3194 78858 3600
rect 79022 3548 79050 3694
rect 79022 3520 79322 3548
rect 79294 3318 79322 3520
rect 1454 1192 1482 1258
rect 1440 1164 1482 1192
rect 816 252 844 1006
rect 1280 252 1308 1006
rect 1440 252 1468 1164
rect 1918 1112 1946 1258
rect 1904 1084 1946 1112
rect 2050 1112 2078 1258
rect 2514 1192 2542 1258
rect 2702 1192 2730 1258
rect 2514 1164 2556 1192
rect 2050 1084 2092 1112
rect 1904 252 1932 1084
rect 2064 252 2092 1084
rect 2528 252 2556 1164
rect 2688 1164 2730 1192
rect 2688 252 2716 1164
rect 3166 1112 3194 1258
rect 3152 1084 3194 1112
rect 3298 1112 3326 1258
rect 3762 1192 3790 1258
rect 3950 1192 3978 1258
rect 3762 1164 3804 1192
rect 3298 1084 3340 1112
rect 3152 252 3180 1084
rect 3312 252 3340 1084
rect 3776 252 3804 1164
rect 3936 1164 3978 1192
rect 3936 252 3964 1164
rect 4414 1112 4442 1258
rect 4400 1084 4442 1112
rect 4546 1112 4574 1258
rect 5010 1192 5038 1258
rect 5198 1192 5226 1258
rect 5010 1164 5052 1192
rect 4546 1084 4588 1112
rect 4400 252 4428 1084
rect 4560 252 4588 1084
rect 5024 252 5052 1164
rect 5184 1164 5226 1192
rect 5184 252 5212 1164
rect 5662 1112 5690 1258
rect 5648 1084 5690 1112
rect 5794 1112 5822 1258
rect 6258 1192 6286 1258
rect 6446 1192 6474 1258
rect 6258 1164 6300 1192
rect 5794 1084 5836 1112
rect 5648 252 5676 1084
rect 5808 252 5836 1084
rect 6272 252 6300 1164
rect 6432 1164 6474 1192
rect 6432 252 6460 1164
rect 6910 1112 6938 1258
rect 6896 1084 6938 1112
rect 7042 1112 7070 1258
rect 7506 1192 7534 1258
rect 7694 1192 7722 1258
rect 7506 1164 7548 1192
rect 7042 1084 7084 1112
rect 6896 252 6924 1084
rect 7056 252 7084 1084
rect 7520 252 7548 1164
rect 7680 1164 7722 1192
rect 7680 252 7708 1164
rect 8158 1112 8186 1258
rect 8144 1084 8186 1112
rect 8290 1112 8318 1258
rect 8754 1192 8782 1258
rect 8942 1192 8970 1258
rect 8754 1164 8796 1192
rect 8290 1084 8332 1112
rect 8144 252 8172 1084
rect 8304 252 8332 1084
rect 8768 252 8796 1164
rect 8928 1164 8970 1192
rect 8928 252 8956 1164
rect 9406 1112 9434 1258
rect 9392 1084 9434 1112
rect 9538 1112 9566 1258
rect 10002 1192 10030 1258
rect 10190 1192 10218 1258
rect 10002 1164 10044 1192
rect 9538 1084 9580 1112
rect 9392 252 9420 1084
rect 9552 252 9580 1084
rect 10016 252 10044 1164
rect 10176 1164 10218 1192
rect 10176 252 10204 1164
rect 10654 1112 10682 1258
rect 10640 1084 10682 1112
rect 10786 1112 10814 1258
rect 11250 1192 11278 1258
rect 11438 1192 11466 1258
rect 11250 1164 11292 1192
rect 10786 1084 10828 1112
rect 10640 252 10668 1084
rect 10800 252 10828 1084
rect 11264 252 11292 1164
rect 11424 1164 11466 1192
rect 11424 252 11452 1164
rect 11902 1112 11930 1258
rect 11888 1084 11930 1112
rect 12034 1112 12062 1258
rect 12498 1192 12526 1258
rect 12686 1192 12714 1258
rect 12498 1164 12540 1192
rect 12034 1084 12076 1112
rect 11888 252 11916 1084
rect 12048 252 12076 1084
rect 12512 252 12540 1164
rect 12672 1164 12714 1192
rect 12672 252 12700 1164
rect 13150 1112 13178 1258
rect 13136 1084 13178 1112
rect 13282 1112 13310 1258
rect 13746 1192 13774 1258
rect 13934 1192 13962 1258
rect 13746 1164 13788 1192
rect 13282 1084 13324 1112
rect 13136 252 13164 1084
rect 13296 252 13324 1084
rect 13760 252 13788 1164
rect 13920 1164 13962 1192
rect 13920 252 13948 1164
rect 14398 1112 14426 1258
rect 14384 1084 14426 1112
rect 14530 1112 14558 1258
rect 14994 1192 15022 1258
rect 15182 1192 15210 1258
rect 14994 1164 15036 1192
rect 14530 1084 14572 1112
rect 14384 252 14412 1084
rect 14544 252 14572 1084
rect 15008 252 15036 1164
rect 15168 1164 15210 1192
rect 15168 252 15196 1164
rect 15646 1112 15674 1258
rect 15632 1084 15674 1112
rect 15778 1112 15806 1258
rect 16242 1192 16270 1258
rect 16430 1192 16458 1258
rect 16242 1164 16284 1192
rect 15778 1084 15820 1112
rect 15632 252 15660 1084
rect 15792 252 15820 1084
rect 16256 252 16284 1164
rect 16416 1164 16458 1192
rect 16416 252 16444 1164
rect 16894 1112 16922 1258
rect 16880 1084 16922 1112
rect 17026 1112 17054 1258
rect 17490 1192 17518 1258
rect 17678 1192 17706 1258
rect 17490 1164 17532 1192
rect 17026 1084 17068 1112
rect 16880 252 16908 1084
rect 17040 252 17068 1084
rect 17504 252 17532 1164
rect 17664 1164 17706 1192
rect 17664 252 17692 1164
rect 18142 1112 18170 1258
rect 18128 1084 18170 1112
rect 18274 1112 18302 1258
rect 18738 1192 18766 1258
rect 18926 1192 18954 1258
rect 18738 1164 18780 1192
rect 18274 1084 18316 1112
rect 18128 252 18156 1084
rect 18288 252 18316 1084
rect 18752 252 18780 1164
rect 18912 1164 18954 1192
rect 18912 252 18940 1164
rect 19390 1112 19418 1258
rect 19376 1084 19418 1112
rect 19522 1112 19550 1258
rect 19986 1192 20014 1258
rect 20174 1192 20202 1258
rect 19986 1164 20028 1192
rect 19522 1084 19564 1112
rect 19376 252 19404 1084
rect 19536 252 19564 1084
rect 20000 252 20028 1164
rect 20160 1164 20202 1192
rect 20160 252 20188 1164
rect 20638 1112 20666 1258
rect 20624 1084 20666 1112
rect 20770 1112 20798 1258
rect 21234 1192 21262 1258
rect 21422 1192 21450 1258
rect 21234 1164 21276 1192
rect 20770 1084 20812 1112
rect 20624 252 20652 1084
rect 20784 252 20812 1084
rect 21248 252 21276 1164
rect 21408 1164 21450 1192
rect 21408 252 21436 1164
rect 21886 1112 21914 1258
rect 21872 1084 21914 1112
rect 22018 1112 22046 1258
rect 22482 1192 22510 1258
rect 22670 1192 22698 1258
rect 22482 1164 22524 1192
rect 22018 1084 22060 1112
rect 21872 252 21900 1084
rect 22032 252 22060 1084
rect 22496 252 22524 1164
rect 22656 1164 22698 1192
rect 22656 252 22684 1164
rect 23134 1112 23162 1258
rect 23120 1084 23162 1112
rect 23266 1112 23294 1258
rect 23730 1192 23758 1258
rect 23918 1192 23946 1258
rect 23730 1164 23772 1192
rect 23266 1084 23308 1112
rect 23120 252 23148 1084
rect 23280 252 23308 1084
rect 23744 252 23772 1164
rect 23904 1164 23946 1192
rect 23904 252 23932 1164
rect 24382 1112 24410 1258
rect 24368 1084 24410 1112
rect 24514 1112 24542 1258
rect 24978 1192 25006 1258
rect 25166 1192 25194 1258
rect 24978 1164 25020 1192
rect 24514 1084 24556 1112
rect 24368 252 24396 1084
rect 24528 252 24556 1084
rect 24992 252 25020 1164
rect 25152 1164 25194 1192
rect 25152 252 25180 1164
rect 25630 1112 25658 1258
rect 25616 1084 25658 1112
rect 25762 1112 25790 1258
rect 26226 1192 26254 1258
rect 26414 1192 26442 1258
rect 26226 1164 26268 1192
rect 25762 1084 25804 1112
rect 25616 252 25644 1084
rect 25776 252 25804 1084
rect 26240 252 26268 1164
rect 26400 1164 26442 1192
rect 26400 252 26428 1164
rect 26878 1112 26906 1258
rect 26864 1084 26906 1112
rect 27010 1112 27038 1258
rect 27474 1192 27502 1258
rect 27662 1192 27690 1258
rect 27474 1164 27516 1192
rect 27010 1084 27052 1112
rect 26864 252 26892 1084
rect 27024 252 27052 1084
rect 27488 252 27516 1164
rect 27648 1164 27690 1192
rect 27648 252 27676 1164
rect 28126 1112 28154 1258
rect 28112 1084 28154 1112
rect 28258 1112 28286 1258
rect 28722 1192 28750 1258
rect 28910 1192 28938 1258
rect 28722 1164 28764 1192
rect 28258 1084 28300 1112
rect 28112 252 28140 1084
rect 28272 252 28300 1084
rect 28736 252 28764 1164
rect 28896 1164 28938 1192
rect 28896 252 28924 1164
rect 29374 1112 29402 1258
rect 29360 1084 29402 1112
rect 29506 1112 29534 1258
rect 29970 1192 29998 1258
rect 30158 1192 30186 1258
rect 29970 1164 30012 1192
rect 29506 1084 29548 1112
rect 29360 252 29388 1084
rect 29520 252 29548 1084
rect 29984 252 30012 1164
rect 30144 1164 30186 1192
rect 30144 252 30172 1164
rect 30622 1112 30650 1258
rect 30608 1084 30650 1112
rect 30754 1112 30782 1258
rect 31218 1192 31246 1258
rect 31406 1192 31434 1258
rect 31218 1164 31260 1192
rect 30754 1084 30796 1112
rect 30608 252 30636 1084
rect 30768 252 30796 1084
rect 31232 252 31260 1164
rect 31392 1164 31434 1192
rect 31392 252 31420 1164
rect 31870 1112 31898 1258
rect 31856 1084 31898 1112
rect 32002 1112 32030 1258
rect 32466 1192 32494 1258
rect 32654 1192 32682 1258
rect 32466 1164 32508 1192
rect 32002 1084 32044 1112
rect 31856 252 31884 1084
rect 32016 252 32044 1084
rect 32480 252 32508 1164
rect 32640 1164 32682 1192
rect 32640 252 32668 1164
rect 33118 1112 33146 1258
rect 33104 1084 33146 1112
rect 33250 1112 33278 1258
rect 33714 1192 33742 1258
rect 33902 1192 33930 1258
rect 33714 1164 33756 1192
rect 33250 1084 33292 1112
rect 33104 252 33132 1084
rect 33264 252 33292 1084
rect 33728 252 33756 1164
rect 33888 1164 33930 1192
rect 33888 252 33916 1164
rect 34366 1112 34394 1258
rect 34352 1084 34394 1112
rect 34498 1112 34526 1258
rect 34962 1192 34990 1258
rect 35150 1192 35178 1258
rect 34962 1164 35004 1192
rect 34498 1084 34540 1112
rect 34352 252 34380 1084
rect 34512 252 34540 1084
rect 34976 252 35004 1164
rect 35136 1164 35178 1192
rect 35136 252 35164 1164
rect 35614 1112 35642 1258
rect 35600 1084 35642 1112
rect 35746 1112 35774 1258
rect 36210 1192 36238 1258
rect 36398 1192 36426 1258
rect 36210 1164 36252 1192
rect 35746 1084 35788 1112
rect 35600 252 35628 1084
rect 35760 252 35788 1084
rect 36224 252 36252 1164
rect 36384 1164 36426 1192
rect 36384 252 36412 1164
rect 36862 1112 36890 1258
rect 36848 1084 36890 1112
rect 36994 1112 37022 1258
rect 37458 1192 37486 1258
rect 37646 1192 37674 1258
rect 37458 1164 37500 1192
rect 36994 1084 37036 1112
rect 36848 252 36876 1084
rect 37008 252 37036 1084
rect 37472 252 37500 1164
rect 37632 1164 37674 1192
rect 37632 252 37660 1164
rect 38110 1112 38138 1258
rect 38096 1084 38138 1112
rect 38242 1112 38270 1258
rect 38706 1192 38734 1258
rect 38894 1192 38922 1258
rect 38706 1164 38748 1192
rect 38242 1084 38284 1112
rect 38096 252 38124 1084
rect 38256 252 38284 1084
rect 38720 252 38748 1164
rect 38880 1164 38922 1192
rect 38880 252 38908 1164
rect 39358 1112 39386 1258
rect 39344 1084 39386 1112
rect 39490 1112 39518 1258
rect 39954 1192 39982 1258
rect 40142 1192 40170 1258
rect 39954 1164 39996 1192
rect 39490 1084 39532 1112
rect 39344 252 39372 1084
rect 39504 252 39532 1084
rect 39968 252 39996 1164
rect 40128 1164 40170 1192
rect 40128 252 40156 1164
rect 40606 1112 40634 1258
rect 40592 1084 40634 1112
rect 40738 1112 40766 1258
rect 41202 1192 41230 1258
rect 41390 1192 41418 1258
rect 41202 1164 41244 1192
rect 40738 1084 40780 1112
rect 40592 252 40620 1084
rect 40752 252 40780 1084
rect 41216 252 41244 1164
rect 41376 1164 41418 1192
rect 41376 252 41404 1164
rect 41854 1112 41882 1258
rect 41840 1084 41882 1112
rect 41986 1112 42014 1258
rect 42450 1192 42478 1258
rect 42638 1192 42666 1258
rect 42450 1164 42492 1192
rect 41986 1084 42028 1112
rect 41840 252 41868 1084
rect 42000 252 42028 1084
rect 42464 252 42492 1164
rect 42624 1164 42666 1192
rect 42624 252 42652 1164
rect 43102 1112 43130 1258
rect 43088 1084 43130 1112
rect 43234 1112 43262 1258
rect 43698 1192 43726 1258
rect 43886 1192 43914 1258
rect 43698 1164 43740 1192
rect 43234 1084 43276 1112
rect 43088 252 43116 1084
rect 43248 252 43276 1084
rect 43712 252 43740 1164
rect 43872 1164 43914 1192
rect 43872 252 43900 1164
rect 44350 1112 44378 1258
rect 44336 1084 44378 1112
rect 44482 1112 44510 1258
rect 44946 1192 44974 1258
rect 45134 1192 45162 1258
rect 44946 1164 44988 1192
rect 44482 1084 44524 1112
rect 44336 252 44364 1084
rect 44496 252 44524 1084
rect 44960 252 44988 1164
rect 45120 1164 45162 1192
rect 45120 252 45148 1164
rect 45598 1112 45626 1258
rect 45584 1084 45626 1112
rect 45730 1112 45758 1258
rect 46194 1192 46222 1258
rect 46382 1192 46410 1258
rect 46194 1164 46236 1192
rect 45730 1084 45772 1112
rect 45584 252 45612 1084
rect 45744 252 45772 1084
rect 46208 252 46236 1164
rect 46368 1164 46410 1192
rect 46368 252 46396 1164
rect 46846 1112 46874 1258
rect 46832 1084 46874 1112
rect 46978 1112 47006 1258
rect 47442 1192 47470 1258
rect 47630 1192 47658 1258
rect 47442 1164 47484 1192
rect 46978 1084 47020 1112
rect 46832 252 46860 1084
rect 46992 252 47020 1084
rect 47456 252 47484 1164
rect 47616 1164 47658 1192
rect 47616 252 47644 1164
rect 48094 1112 48122 1258
rect 48080 1084 48122 1112
rect 48226 1112 48254 1258
rect 48690 1192 48718 1258
rect 48878 1192 48906 1258
rect 48690 1164 48732 1192
rect 48226 1084 48268 1112
rect 48080 252 48108 1084
rect 48240 252 48268 1084
rect 48704 252 48732 1164
rect 48864 1164 48906 1192
rect 48864 252 48892 1164
rect 49342 1112 49370 1258
rect 49328 1084 49370 1112
rect 49474 1112 49502 1258
rect 49938 1192 49966 1258
rect 50126 1192 50154 1258
rect 49938 1164 49980 1192
rect 49474 1084 49516 1112
rect 49328 252 49356 1084
rect 49488 252 49516 1084
rect 49952 252 49980 1164
rect 50112 1164 50154 1192
rect 50112 252 50140 1164
rect 50590 1112 50618 1258
rect 50576 1084 50618 1112
rect 50722 1112 50750 1258
rect 51186 1192 51214 1258
rect 51374 1192 51402 1258
rect 51186 1164 51228 1192
rect 50722 1084 50764 1112
rect 50576 252 50604 1084
rect 50736 252 50764 1084
rect 51200 252 51228 1164
rect 51360 1164 51402 1192
rect 51360 252 51388 1164
rect 51838 1112 51866 1258
rect 51824 1084 51866 1112
rect 51970 1112 51998 1258
rect 52434 1192 52462 1258
rect 52622 1192 52650 1258
rect 52434 1164 52476 1192
rect 51970 1084 52012 1112
rect 51824 252 51852 1084
rect 51984 252 52012 1084
rect 52448 252 52476 1164
rect 52608 1164 52650 1192
rect 52608 252 52636 1164
rect 53086 1112 53114 1258
rect 53072 1084 53114 1112
rect 53218 1112 53246 1258
rect 53682 1192 53710 1258
rect 53870 1192 53898 1258
rect 53682 1164 53724 1192
rect 53218 1084 53260 1112
rect 53072 252 53100 1084
rect 53232 252 53260 1084
rect 53696 252 53724 1164
rect 53856 1164 53898 1192
rect 53856 252 53884 1164
rect 54334 1112 54362 1258
rect 54320 1084 54362 1112
rect 54466 1112 54494 1258
rect 54930 1192 54958 1258
rect 55118 1192 55146 1258
rect 54930 1164 54972 1192
rect 54466 1084 54508 1112
rect 54320 252 54348 1084
rect 54480 252 54508 1084
rect 54944 252 54972 1164
rect 55104 1164 55146 1192
rect 55104 252 55132 1164
rect 55582 1112 55610 1258
rect 55568 1084 55610 1112
rect 55714 1112 55742 1258
rect 56178 1192 56206 1258
rect 56366 1192 56394 1258
rect 56178 1164 56220 1192
rect 55714 1084 55756 1112
rect 55568 252 55596 1084
rect 55728 252 55756 1084
rect 56192 252 56220 1164
rect 56352 1164 56394 1192
rect 56352 252 56380 1164
rect 56830 1112 56858 1258
rect 56816 1084 56858 1112
rect 56962 1112 56990 1258
rect 57426 1192 57454 1258
rect 57614 1192 57642 1258
rect 57426 1164 57468 1192
rect 56962 1084 57004 1112
rect 56816 252 56844 1084
rect 56976 252 57004 1084
rect 57440 252 57468 1164
rect 57600 1164 57642 1192
rect 57600 252 57628 1164
rect 58078 1112 58106 1258
rect 58064 1084 58106 1112
rect 58210 1112 58238 1258
rect 58674 1192 58702 1258
rect 58862 1192 58890 1258
rect 58674 1164 58716 1192
rect 58210 1084 58252 1112
rect 58064 252 58092 1084
rect 58224 252 58252 1084
rect 58688 252 58716 1164
rect 58848 1164 58890 1192
rect 58848 252 58876 1164
rect 59326 1112 59354 1258
rect 59312 1084 59354 1112
rect 59458 1112 59486 1258
rect 59922 1192 59950 1258
rect 60110 1192 60138 1258
rect 59922 1164 59964 1192
rect 59458 1084 59500 1112
rect 59312 252 59340 1084
rect 59472 252 59500 1084
rect 59936 252 59964 1164
rect 60096 1164 60138 1192
rect 60096 252 60124 1164
rect 60574 1112 60602 1258
rect 60560 1084 60602 1112
rect 60706 1112 60734 1258
rect 61170 1192 61198 1258
rect 61358 1192 61386 1258
rect 61170 1164 61212 1192
rect 60706 1084 60748 1112
rect 60560 252 60588 1084
rect 60720 252 60748 1084
rect 61184 252 61212 1164
rect 61344 1164 61386 1192
rect 61344 252 61372 1164
rect 61822 1112 61850 1258
rect 61808 1084 61850 1112
rect 61954 1112 61982 1258
rect 62418 1192 62446 1258
rect 62606 1192 62634 1258
rect 62418 1164 62460 1192
rect 61954 1084 61996 1112
rect 61808 252 61836 1084
rect 61968 252 61996 1084
rect 62432 252 62460 1164
rect 62592 1164 62634 1192
rect 62592 252 62620 1164
rect 63070 1112 63098 1258
rect 63056 1084 63098 1112
rect 63202 1112 63230 1258
rect 63666 1192 63694 1258
rect 63854 1192 63882 1258
rect 63666 1164 63708 1192
rect 63202 1084 63244 1112
rect 63056 252 63084 1084
rect 63216 252 63244 1084
rect 63680 252 63708 1164
rect 63840 1164 63882 1192
rect 63840 252 63868 1164
rect 64318 1112 64346 1258
rect 64304 1084 64346 1112
rect 64450 1112 64478 1258
rect 64914 1192 64942 1258
rect 65102 1192 65130 1258
rect 64914 1164 64956 1192
rect 64450 1084 64492 1112
rect 64304 252 64332 1084
rect 64464 252 64492 1084
rect 64928 252 64956 1164
rect 65088 1164 65130 1192
rect 65088 252 65116 1164
rect 65566 1112 65594 1258
rect 65552 1084 65594 1112
rect 65698 1112 65726 1258
rect 66162 1192 66190 1258
rect 66350 1192 66378 1258
rect 66162 1164 66204 1192
rect 65698 1084 65740 1112
rect 65552 252 65580 1084
rect 65712 252 65740 1084
rect 66176 252 66204 1164
rect 66336 1164 66378 1192
rect 66336 252 66364 1164
rect 66814 1112 66842 1258
rect 66800 1084 66842 1112
rect 66946 1112 66974 1258
rect 67410 1192 67438 1258
rect 67598 1192 67626 1258
rect 67410 1164 67452 1192
rect 66946 1084 66988 1112
rect 66800 252 66828 1084
rect 66960 252 66988 1084
rect 67424 252 67452 1164
rect 67584 1164 67626 1192
rect 67584 252 67612 1164
rect 68062 1112 68090 1258
rect 68048 1084 68090 1112
rect 68194 1112 68222 1258
rect 68658 1192 68686 1258
rect 68846 1192 68874 1258
rect 68658 1164 68700 1192
rect 68194 1084 68236 1112
rect 68048 252 68076 1084
rect 68208 252 68236 1084
rect 68672 252 68700 1164
rect 68832 1164 68874 1192
rect 68832 252 68860 1164
rect 69310 1112 69338 1258
rect 69296 1084 69338 1112
rect 69442 1112 69470 1258
rect 69906 1192 69934 1258
rect 70094 1192 70122 1258
rect 69906 1164 69948 1192
rect 69442 1084 69484 1112
rect 69296 252 69324 1084
rect 69456 252 69484 1084
rect 69920 252 69948 1164
rect 70080 1164 70122 1192
rect 70080 252 70108 1164
rect 70558 1112 70586 1258
rect 70544 1084 70586 1112
rect 70690 1112 70718 1258
rect 71154 1192 71182 1258
rect 71342 1192 71370 1258
rect 71154 1164 71196 1192
rect 70690 1084 70732 1112
rect 70544 252 70572 1084
rect 70704 252 70732 1084
rect 71168 252 71196 1164
rect 71328 1164 71370 1192
rect 71328 252 71356 1164
rect 71806 1112 71834 1258
rect 71792 1084 71834 1112
rect 71938 1112 71966 1258
rect 72402 1192 72430 1258
rect 72590 1192 72618 1258
rect 72402 1164 72444 1192
rect 71938 1084 71980 1112
rect 71792 252 71820 1084
rect 71952 252 71980 1084
rect 72416 252 72444 1164
rect 72576 1164 72618 1192
rect 72576 252 72604 1164
rect 73054 1112 73082 1258
rect 73040 1084 73082 1112
rect 73186 1112 73214 1258
rect 73650 1192 73678 1258
rect 73838 1192 73866 1258
rect 73650 1164 73692 1192
rect 73186 1084 73228 1112
rect 73040 252 73068 1084
rect 73200 252 73228 1084
rect 73664 252 73692 1164
rect 73824 1164 73866 1192
rect 73824 252 73852 1164
rect 74302 1112 74330 1258
rect 74288 1084 74330 1112
rect 74434 1112 74462 1258
rect 74898 1192 74926 1258
rect 75086 1192 75114 1258
rect 74898 1164 74940 1192
rect 74434 1084 74476 1112
rect 74288 252 74316 1084
rect 74448 252 74476 1084
rect 74912 252 74940 1164
rect 75072 1164 75114 1192
rect 75072 252 75100 1164
rect 75550 1112 75578 1258
rect 75536 1084 75578 1112
rect 75682 1112 75710 1258
rect 76146 1192 76174 1258
rect 76334 1192 76362 1258
rect 76146 1164 76188 1192
rect 75682 1084 75724 1112
rect 75536 252 75564 1084
rect 75696 252 75724 1084
rect 76160 252 76188 1164
rect 76320 1164 76362 1192
rect 76320 252 76348 1164
rect 76798 1112 76826 1258
rect 76784 1084 76826 1112
rect 76930 1112 76958 1258
rect 77394 1192 77422 1258
rect 77582 1192 77610 1258
rect 77394 1164 77436 1192
rect 76930 1084 76972 1112
rect 76784 252 76812 1084
rect 76944 252 76972 1084
rect 77408 252 77436 1164
rect 77568 1164 77610 1192
rect 77568 252 77596 1164
rect 78046 1112 78074 1258
rect 78032 1084 78074 1112
rect 78178 1112 78206 1258
rect 78642 1192 78670 1258
rect 78830 1192 78858 1258
rect 78642 1164 78684 1192
rect 78178 1084 78220 1112
rect 78032 252 78060 1084
rect 78192 252 78220 1084
rect 78656 252 78684 1164
rect 78816 1164 78858 1192
rect 78816 252 78844 1164
rect 79294 1112 79322 1258
rect 79280 1084 79322 1112
rect 79426 1112 79454 1258
rect 79890 1192 79918 1258
rect 80078 1192 80106 1258
rect 79890 1164 79932 1192
rect 79426 1084 79468 1112
rect 79280 252 79308 1084
rect 79440 252 79468 1084
rect 79904 252 79932 1164
rect 80064 1164 80106 1192
rect 80064 252 80092 1164
rect 80542 1112 80570 1258
rect 80528 1084 80570 1112
rect 80674 1112 80702 1258
rect 81138 1192 81166 1258
rect 81138 1164 81180 1192
rect 80674 1084 80716 1112
rect 80528 252 80556 1084
rect 80688 252 80716 1084
rect 81152 252 81180 1164
<< via1 >>
rect 20707 9025 20759 9077
rect 40675 9025 40727 9077
rect 60643 9025 60695 9077
rect 80611 9025 80663 9077
rect 20707 8076 20759 8128
rect 40675 8076 40727 8128
rect 60643 8076 60695 8128
rect 80611 8076 80663 8128
<< metal2 >>
rect 1360 9301 1388 9329
rect 21328 9301 21356 9329
rect 41296 9301 41324 9329
rect 61264 9301 61292 9329
rect 20707 9077 20759 9083
rect 20707 9019 20759 9025
rect 40675 9077 40727 9083
rect 40675 9019 40727 9025
rect 60643 9077 60695 9083
rect 60643 9019 60695 9025
rect 80611 9077 80663 9083
rect 80611 9019 80663 9025
rect 20719 8134 20747 9019
rect 40687 8134 40715 9019
rect 60655 8134 60683 9019
rect 80623 8134 80651 9019
rect 20707 8128 20759 8134
rect 20707 8070 20759 8076
rect 40675 8128 40727 8134
rect 40675 8070 40727 8076
rect 60643 8128 60695 8134
rect 60643 8070 60695 8076
rect 80611 8128 80663 8134
rect 80611 8070 80663 8076
<< metal3 >>
rect -49 9536 49 9634
rect 81197 9536 81295 9634
rect 0 9037 81246 9097
rect -49 8416 49 8514
rect 81197 8416 81295 8514
rect 1601 7973 1699 8071
rect 4097 7973 4195 8071
rect 6593 7973 6691 8071
rect 9089 7973 9187 8071
rect 11585 7973 11683 8071
rect 14081 7973 14179 8071
rect 16577 7973 16675 8071
rect 19073 7973 19171 8071
rect 21569 7973 21667 8071
rect 24065 7973 24163 8071
rect 26561 7973 26659 8071
rect 29057 7973 29155 8071
rect 31553 7973 31651 8071
rect 34049 7973 34147 8071
rect 36545 7973 36643 8071
rect 39041 7973 39139 8071
rect 41537 7973 41635 8071
rect 44033 7973 44131 8071
rect 46529 7973 46627 8071
rect 49025 7973 49123 8071
rect 51521 7973 51619 8071
rect 54017 7973 54115 8071
rect 56513 7973 56611 8071
rect 59009 7973 59107 8071
rect 61505 7973 61603 8071
rect 64001 7973 64099 8071
rect 66497 7973 66595 8071
rect 68993 7973 69091 8071
rect 71489 7973 71587 8071
rect 73985 7973 74083 8071
rect 76481 7973 76579 8071
rect 78977 7973 79075 8071
rect 1587 7557 1685 7655
rect 4083 7557 4181 7655
rect 6579 7557 6677 7655
rect 9075 7557 9173 7655
rect 11571 7557 11669 7655
rect 14067 7557 14165 7655
rect 16563 7557 16661 7655
rect 19059 7557 19157 7655
rect 21555 7557 21653 7655
rect 24051 7557 24149 7655
rect 26547 7557 26645 7655
rect 29043 7557 29141 7655
rect 31539 7557 31637 7655
rect 34035 7557 34133 7655
rect 36531 7557 36629 7655
rect 39027 7557 39125 7655
rect 41523 7557 41621 7655
rect 44019 7557 44117 7655
rect 46515 7557 46613 7655
rect 49011 7557 49109 7655
rect 51507 7557 51605 7655
rect 54003 7557 54101 7655
rect 56499 7557 56597 7655
rect 58995 7557 59093 7655
rect 61491 7557 61589 7655
rect 63987 7557 64085 7655
rect 66483 7557 66581 7655
rect 68979 7557 69077 7655
rect 71475 7557 71573 7655
rect 73971 7557 74069 7655
rect 76467 7557 76565 7655
rect 78963 7557 79061 7655
rect 1702 7355 1800 7453
rect 4198 7355 4296 7453
rect 6694 7355 6792 7453
rect 9190 7355 9288 7453
rect 11686 7355 11784 7453
rect 14182 7355 14280 7453
rect 16678 7355 16776 7453
rect 19174 7355 19272 7453
rect 21670 7355 21768 7453
rect 24166 7355 24264 7453
rect 26662 7355 26760 7453
rect 29158 7355 29256 7453
rect 31654 7355 31752 7453
rect 34150 7355 34248 7453
rect 36646 7355 36744 7453
rect 39142 7355 39240 7453
rect 41638 7355 41736 7453
rect 44134 7355 44232 7453
rect 46630 7355 46728 7453
rect 49126 7355 49224 7453
rect 51622 7355 51720 7453
rect 54118 7355 54216 7453
rect 56614 7355 56712 7453
rect 59110 7355 59208 7453
rect 61606 7355 61704 7453
rect 64102 7355 64200 7453
rect 66598 7355 66696 7453
rect 69094 7355 69192 7453
rect 71590 7355 71688 7453
rect 74086 7355 74184 7453
rect 76582 7355 76680 7453
rect 79078 7355 79176 7453
rect 1581 7023 1679 7121
rect 4077 7023 4175 7121
rect 6573 7023 6671 7121
rect 9069 7023 9167 7121
rect 11565 7023 11663 7121
rect 14061 7023 14159 7121
rect 16557 7023 16655 7121
rect 19053 7023 19151 7121
rect 21549 7023 21647 7121
rect 24045 7023 24143 7121
rect 26541 7023 26639 7121
rect 29037 7023 29135 7121
rect 31533 7023 31631 7121
rect 34029 7023 34127 7121
rect 36525 7023 36623 7121
rect 39021 7023 39119 7121
rect 41517 7023 41615 7121
rect 44013 7023 44111 7121
rect 46509 7023 46607 7121
rect 49005 7023 49103 7121
rect 51501 7023 51599 7121
rect 53997 7023 54095 7121
rect 56493 7023 56591 7121
rect 58989 7023 59087 7121
rect 61485 7023 61583 7121
rect 63981 7023 64079 7121
rect 66477 7023 66575 7121
rect 68973 7023 69071 7121
rect 71469 7023 71567 7121
rect 73965 7023 74063 7121
rect 76461 7023 76559 7121
rect 78957 7023 79055 7121
rect 1592 6586 1690 6684
rect 4088 6586 4186 6684
rect 6584 6586 6682 6684
rect 9080 6586 9178 6684
rect 11576 6586 11674 6684
rect 14072 6586 14170 6684
rect 16568 6586 16666 6684
rect 19064 6586 19162 6684
rect 21560 6586 21658 6684
rect 24056 6586 24154 6684
rect 26552 6586 26650 6684
rect 29048 6586 29146 6684
rect 31544 6586 31642 6684
rect 34040 6586 34138 6684
rect 36536 6586 36634 6684
rect 39032 6586 39130 6684
rect 41528 6586 41626 6684
rect 44024 6586 44122 6684
rect 46520 6586 46618 6684
rect 49016 6586 49114 6684
rect 51512 6586 51610 6684
rect 54008 6586 54106 6684
rect 56504 6586 56602 6684
rect 59000 6586 59098 6684
rect 61496 6586 61594 6684
rect 63992 6586 64090 6684
rect 66488 6586 66586 6684
rect 68984 6586 69082 6684
rect 71480 6586 71578 6684
rect 73976 6586 74074 6684
rect 76472 6586 76570 6684
rect 78968 6586 79066 6684
rect 1706 5793 1804 5891
rect 4202 5793 4300 5891
rect 6698 5793 6796 5891
rect 9194 5793 9292 5891
rect 11690 5793 11788 5891
rect 14186 5793 14284 5891
rect 16682 5793 16780 5891
rect 19178 5793 19276 5891
rect 21674 5793 21772 5891
rect 24170 5793 24268 5891
rect 26666 5793 26764 5891
rect 29162 5793 29260 5891
rect 31658 5793 31756 5891
rect 34154 5793 34252 5891
rect 36650 5793 36748 5891
rect 39146 5793 39244 5891
rect 41642 5793 41740 5891
rect 44138 5793 44236 5891
rect 46634 5793 46732 5891
rect 49130 5793 49228 5891
rect 51626 5793 51724 5891
rect 54122 5793 54220 5891
rect 56618 5793 56716 5891
rect 59114 5793 59212 5891
rect 61610 5793 61708 5891
rect 64106 5793 64204 5891
rect 66602 5793 66700 5891
rect 69098 5793 69196 5891
rect 71594 5793 71692 5891
rect 74090 5793 74188 5891
rect 76586 5793 76684 5891
rect 79082 5793 79180 5891
rect 1706 5471 1804 5569
rect 4202 5471 4300 5569
rect 6698 5471 6796 5569
rect 9194 5471 9292 5569
rect 11690 5471 11788 5569
rect 14186 5471 14284 5569
rect 16682 5471 16780 5569
rect 19178 5471 19276 5569
rect 21674 5471 21772 5569
rect 24170 5471 24268 5569
rect 26666 5471 26764 5569
rect 29162 5471 29260 5569
rect 31658 5471 31756 5569
rect 34154 5471 34252 5569
rect 36650 5471 36748 5569
rect 39146 5471 39244 5569
rect 41642 5471 41740 5569
rect 44138 5471 44236 5569
rect 46634 5471 46732 5569
rect 49130 5471 49228 5569
rect 51626 5471 51724 5569
rect 54122 5471 54220 5569
rect 56618 5471 56716 5569
rect 59114 5471 59212 5569
rect 61610 5471 61708 5569
rect 64106 5471 64204 5569
rect 66602 5471 66700 5569
rect 69098 5471 69196 5569
rect 71594 5471 71692 5569
rect 74090 5471 74188 5569
rect 76586 5471 76684 5569
rect 79082 5471 79180 5569
rect 1694 4633 1792 4731
rect 4190 4633 4288 4731
rect 6686 4633 6784 4731
rect 9182 4633 9280 4731
rect 11678 4633 11776 4731
rect 14174 4633 14272 4731
rect 16670 4633 16768 4731
rect 19166 4633 19264 4731
rect 21662 4633 21760 4731
rect 24158 4633 24256 4731
rect 26654 4633 26752 4731
rect 29150 4633 29248 4731
rect 31646 4633 31744 4731
rect 34142 4633 34240 4731
rect 36638 4633 36736 4731
rect 39134 4633 39232 4731
rect 41630 4633 41728 4731
rect 44126 4633 44224 4731
rect 46622 4633 46720 4731
rect 49118 4633 49216 4731
rect 51614 4633 51712 4731
rect 54110 4633 54208 4731
rect 56606 4633 56704 4731
rect 59102 4633 59200 4731
rect 61598 4633 61696 4731
rect 64094 4633 64192 4731
rect 66590 4633 66688 4731
rect 69086 4633 69184 4731
rect 71582 4633 71680 4731
rect 74078 4633 74176 4731
rect 76574 4633 76672 4731
rect 79070 4633 79168 4731
rect 1776 3859 1874 3957
rect 4272 3859 4370 3957
rect 6768 3859 6866 3957
rect 9264 3859 9362 3957
rect 11760 3859 11858 3957
rect 14256 3859 14354 3957
rect 16752 3859 16850 3957
rect 19248 3859 19346 3957
rect 21744 3859 21842 3957
rect 24240 3859 24338 3957
rect 26736 3859 26834 3957
rect 29232 3859 29330 3957
rect 31728 3859 31826 3957
rect 34224 3859 34322 3957
rect 36720 3859 36818 3957
rect 39216 3859 39314 3957
rect 41712 3859 41810 3957
rect 44208 3859 44306 3957
rect 46704 3859 46802 3957
rect 49200 3859 49298 3957
rect 51696 3859 51794 3957
rect 54192 3859 54290 3957
rect 56688 3859 56786 3957
rect 59184 3859 59282 3957
rect 61680 3859 61778 3957
rect 64176 3859 64274 3957
rect 66672 3859 66770 3957
rect 69168 3859 69266 3957
rect 71664 3859 71762 3957
rect 74160 3859 74258 3957
rect 76656 3859 76754 3957
rect 79152 3859 79250 3957
rect 0 3726 79250 3786
rect 0 3010 81246 3070
rect 0 2886 81246 2946
rect 0 2762 81246 2822
rect 0 2638 81246 2698
rect 1949 1862 2047 1960
rect 3197 1862 3295 1960
rect 4445 1862 4543 1960
rect 5693 1862 5791 1960
rect 6941 1862 7039 1960
rect 8189 1862 8287 1960
rect 9437 1862 9535 1960
rect 10685 1862 10783 1960
rect 11933 1862 12031 1960
rect 13181 1862 13279 1960
rect 14429 1862 14527 1960
rect 15677 1862 15775 1960
rect 16925 1862 17023 1960
rect 18173 1862 18271 1960
rect 19421 1862 19519 1960
rect 20669 1862 20767 1960
rect 21917 1862 22015 1960
rect 23165 1862 23263 1960
rect 24413 1862 24511 1960
rect 25661 1862 25759 1960
rect 26909 1862 27007 1960
rect 28157 1862 28255 1960
rect 29405 1862 29503 1960
rect 30653 1862 30751 1960
rect 31901 1862 31999 1960
rect 33149 1862 33247 1960
rect 34397 1862 34495 1960
rect 35645 1862 35743 1960
rect 36893 1862 36991 1960
rect 38141 1862 38239 1960
rect 39389 1862 39487 1960
rect 40637 1862 40735 1960
rect 41885 1862 41983 1960
rect 43133 1862 43231 1960
rect 44381 1862 44479 1960
rect 45629 1862 45727 1960
rect 46877 1862 46975 1960
rect 48125 1862 48223 1960
rect 49373 1862 49471 1960
rect 50621 1862 50719 1960
rect 51869 1862 51967 1960
rect 53117 1862 53215 1960
rect 54365 1862 54463 1960
rect 55613 1862 55711 1960
rect 56861 1862 56959 1960
rect 58109 1862 58207 1960
rect 59357 1862 59455 1960
rect 60605 1862 60703 1960
rect 61853 1862 61951 1960
rect 63101 1862 63199 1960
rect 64349 1862 64447 1960
rect 65597 1862 65695 1960
rect 66845 1862 66943 1960
rect 68093 1862 68191 1960
rect 69341 1862 69439 1960
rect 70589 1862 70687 1960
rect 71837 1862 71935 1960
rect 73085 1862 73183 1960
rect 74333 1862 74431 1960
rect 75581 1862 75679 1960
rect 76829 1862 76927 1960
rect 78077 1862 78175 1960
rect 79325 1862 79423 1960
rect 80573 1862 80671 1960
rect 0 951 81246 1011
rect 1132 313 1230 411
rect 1518 313 1616 411
rect 2380 313 2478 411
rect 2766 313 2864 411
rect 3628 313 3726 411
rect 4014 313 4112 411
rect 4876 313 4974 411
rect 5262 313 5360 411
rect 6124 313 6222 411
rect 6510 313 6608 411
rect 7372 313 7470 411
rect 7758 313 7856 411
rect 8620 313 8718 411
rect 9006 313 9104 411
rect 9868 313 9966 411
rect 10254 313 10352 411
rect 11116 313 11214 411
rect 11502 313 11600 411
rect 12364 313 12462 411
rect 12750 313 12848 411
rect 13612 313 13710 411
rect 13998 313 14096 411
rect 14860 313 14958 411
rect 15246 313 15344 411
rect 16108 313 16206 411
rect 16494 313 16592 411
rect 17356 313 17454 411
rect 17742 313 17840 411
rect 18604 313 18702 411
rect 18990 313 19088 411
rect 19852 313 19950 411
rect 20238 313 20336 411
rect 21100 313 21198 411
rect 21486 313 21584 411
rect 22348 313 22446 411
rect 22734 313 22832 411
rect 23596 313 23694 411
rect 23982 313 24080 411
rect 24844 313 24942 411
rect 25230 313 25328 411
rect 26092 313 26190 411
rect 26478 313 26576 411
rect 27340 313 27438 411
rect 27726 313 27824 411
rect 28588 313 28686 411
rect 28974 313 29072 411
rect 29836 313 29934 411
rect 30222 313 30320 411
rect 31084 313 31182 411
rect 31470 313 31568 411
rect 32332 313 32430 411
rect 32718 313 32816 411
rect 33580 313 33678 411
rect 33966 313 34064 411
rect 34828 313 34926 411
rect 35214 313 35312 411
rect 36076 313 36174 411
rect 36462 313 36560 411
rect 37324 313 37422 411
rect 37710 313 37808 411
rect 38572 313 38670 411
rect 38958 313 39056 411
rect 39820 313 39918 411
rect 40206 313 40304 411
rect 41068 313 41166 411
rect 41454 313 41552 411
rect 42316 313 42414 411
rect 42702 313 42800 411
rect 43564 313 43662 411
rect 43950 313 44048 411
rect 44812 313 44910 411
rect 45198 313 45296 411
rect 46060 313 46158 411
rect 46446 313 46544 411
rect 47308 313 47406 411
rect 47694 313 47792 411
rect 48556 313 48654 411
rect 48942 313 49040 411
rect 49804 313 49902 411
rect 50190 313 50288 411
rect 51052 313 51150 411
rect 51438 313 51536 411
rect 52300 313 52398 411
rect 52686 313 52784 411
rect 53548 313 53646 411
rect 53934 313 54032 411
rect 54796 313 54894 411
rect 55182 313 55280 411
rect 56044 313 56142 411
rect 56430 313 56528 411
rect 57292 313 57390 411
rect 57678 313 57776 411
rect 58540 313 58638 411
rect 58926 313 59024 411
rect 59788 313 59886 411
rect 60174 313 60272 411
rect 61036 313 61134 411
rect 61422 313 61520 411
rect 62284 313 62382 411
rect 62670 313 62768 411
rect 63532 313 63630 411
rect 63918 313 64016 411
rect 64780 313 64878 411
rect 65166 313 65264 411
rect 66028 313 66126 411
rect 66414 313 66512 411
rect 67276 313 67374 411
rect 67662 313 67760 411
rect 68524 313 68622 411
rect 68910 313 69008 411
rect 69772 313 69870 411
rect 70158 313 70256 411
rect 71020 313 71118 411
rect 71406 313 71504 411
rect 72268 313 72366 411
rect 72654 313 72752 411
rect 73516 313 73614 411
rect 73902 313 74000 411
rect 74764 313 74862 411
rect 75150 313 75248 411
rect 76012 313 76110 411
rect 76398 313 76496 411
rect 77260 313 77358 411
rect 77646 313 77744 411
rect 78508 313 78606 411
rect 78894 313 78992 411
rect 79756 313 79854 411
rect 80142 313 80240 411
rect 81004 313 81102 411
use sky130_sram_2kbyte_1rw1r_32x512_8_column_mux_array  sky130_sram_2kbyte_1rw1r_32x512_8_column_mux_array_0
timestamp 1649977179
transform 1 0 0 0 -1 3442
box 0 87 81246 2184
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_0
timestamp 1649977179
transform 1 0 61827 0 1 9018
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1
timestamp 1649977179
transform 1 0 41859 0 1 9018
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_2
timestamp 1649977179
transform 1 0 21891 0 1 9018
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_3
timestamp 1649977179
transform 1 0 1923 0 1 9018
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_0
timestamp 1649977179
transform 1 0 80605 0 1 9019
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_1
timestamp 1649977179
transform 1 0 80605 0 1 8070
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_2
timestamp 1649977179
transform 1 0 60637 0 1 9019
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_3
timestamp 1649977179
transform 1 0 60637 0 1 8070
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_4
timestamp 1649977179
transform 1 0 40669 0 1 9019
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_5
timestamp 1649977179
transform 1 0 40669 0 1 8070
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_6
timestamp 1649977179
transform 1 0 20701 0 1 9019
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_7
timestamp 1649977179
transform 1 0 20701 0 1 8070
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_precharge_array  sky130_sram_2kbyte_1rw1r_32x512_8_precharge_array_0
timestamp 1649977179
transform 1 0 0 0 -1 1006
box 0 -12 81246 768
use sky130_sram_2kbyte_1rw1r_32x512_8_sense_amp_array  sky130_sram_2kbyte_1rw1r_32x512_8_sense_amp_array_0
timestamp 1649977179
transform 1 0 0 0 -1 5950
box 0 0 79687 2256
use sky130_sram_2kbyte_1rw1r_32x512_8_write_driver_array  sky130_sram_2kbyte_1rw1r_32x512_8_write_driver_array_0
timestamp 1649977179
transform 1 0 0 0 -1 8213
box 998 4 80721 2011
use sky130_sram_2kbyte_1rw1r_32x512_8_write_mask_and_array  sky130_sram_2kbyte_1rw1r_32x512_8_write_mask_and_array_0
timestamp 1649977179
transform 1 0 0 0 -1 9585
box -49 -49 81295 1177
<< labels >>
rlabel metal3 s 69098 5471 69196 5569 4 vdd
port 1 nsew
rlabel metal3 s 76586 5471 76684 5569 4 vdd
port 1 nsew
rlabel metal3 s 73965 7023 74063 7121 4 vdd
port 1 nsew
rlabel metal3 s 66602 5471 66700 5569 4 vdd
port 1 nsew
rlabel metal3 s 61485 7023 61583 7121 4 vdd
port 1 nsew
rlabel metal3 s 69086 4633 69184 4731 4 vdd
port 1 nsew
rlabel metal3 s 66477 7023 66575 7121 4 vdd
port 1 nsew
rlabel metal3 s 68993 7973 69091 8071 4 vdd
port 1 nsew
rlabel metal3 s 81197 8416 81295 8514 4 vdd
port 1 nsew
rlabel metal3 s 76574 4633 76672 4731 4 vdd
port 1 nsew
rlabel metal3 s 79082 5471 79180 5569 4 vdd
port 1 nsew
rlabel metal3 s 78957 7023 79055 7121 4 vdd
port 1 nsew
rlabel metal3 s 61610 5471 61708 5569 4 vdd
port 1 nsew
rlabel metal3 s 61598 4633 61696 4731 4 vdd
port 1 nsew
rlabel metal3 s 61505 7973 61603 8071 4 vdd
port 1 nsew
rlabel metal3 s 66497 7973 66595 8071 4 vdd
port 1 nsew
rlabel metal3 s 64094 4633 64192 4731 4 vdd
port 1 nsew
rlabel metal3 s 71582 4633 71680 4731 4 vdd
port 1 nsew
rlabel metal3 s 66590 4633 66688 4731 4 vdd
port 1 nsew
rlabel metal3 s 63981 7023 64079 7121 4 vdd
port 1 nsew
rlabel metal3 s 74078 4633 74176 4731 4 vdd
port 1 nsew
rlabel metal3 s 78977 7973 79075 8071 4 vdd
port 1 nsew
rlabel metal3 s 64106 5471 64204 5569 4 vdd
port 1 nsew
rlabel metal3 s 73985 7973 74083 8071 4 vdd
port 1 nsew
rlabel metal3 s 76461 7023 76559 7121 4 vdd
port 1 nsew
rlabel metal3 s 74090 5471 74188 5569 4 vdd
port 1 nsew
rlabel metal3 s 76481 7973 76579 8071 4 vdd
port 1 nsew
rlabel metal3 s 64001 7973 64099 8071 4 vdd
port 1 nsew
rlabel metal3 s 71489 7973 71587 8071 4 vdd
port 1 nsew
rlabel metal3 s 79070 4633 79168 4731 4 vdd
port 1 nsew
rlabel metal3 s 71594 5471 71692 5569 4 vdd
port 1 nsew
rlabel metal3 s 68973 7023 69071 7121 4 vdd
port 1 nsew
rlabel metal3 s 71469 7023 71567 7121 4 vdd
port 1 nsew
rlabel metal3 s 65597 1862 65695 1960 4 gnd
port 2 nsew
rlabel metal3 s 71664 3859 71762 3957 4 gnd
port 2 nsew
rlabel metal3 s 69168 3859 69266 3957 4 gnd
port 2 nsew
rlabel metal3 s 68984 6586 69082 6684 4 gnd
port 2 nsew
rlabel metal3 s 66845 1862 66943 1960 4 gnd
port 2 nsew
rlabel metal3 s 79082 5793 79180 5891 4 gnd
port 2 nsew
rlabel metal3 s 61496 6586 61594 6684 4 gnd
port 2 nsew
rlabel metal3 s 68093 1862 68191 1960 4 gnd
port 2 nsew
rlabel metal3 s 78077 1862 78175 1960 4 gnd
port 2 nsew
rlabel metal3 s 63101 1862 63199 1960 4 gnd
port 2 nsew
rlabel metal3 s 66672 3859 66770 3957 4 gnd
port 2 nsew
rlabel metal3 s 66598 7355 66696 7453 4 gnd
port 2 nsew
rlabel metal3 s 64176 3859 64274 3957 4 gnd
port 2 nsew
rlabel metal3 s 69341 1862 69439 1960 4 gnd
port 2 nsew
rlabel metal3 s 63992 6586 64090 6684 4 gnd
port 2 nsew
rlabel metal3 s 81197 9536 81295 9634 4 gnd
port 2 nsew
rlabel metal3 s 73085 1862 73183 1960 4 gnd
port 2 nsew
rlabel metal3 s 61606 7355 61704 7453 4 gnd
port 2 nsew
rlabel metal3 s 73971 7557 74069 7655 4 gnd
port 2 nsew
rlabel metal3 s 64102 7355 64200 7453 4 gnd
port 2 nsew
rlabel metal3 s 66602 5793 66700 5891 4 gnd
port 2 nsew
rlabel metal3 s 71480 6586 71578 6684 4 gnd
port 2 nsew
rlabel metal3 s 69094 7355 69192 7453 4 gnd
port 2 nsew
rlabel metal3 s 76467 7557 76565 7655 4 gnd
port 2 nsew
rlabel metal3 s 66488 6586 66586 6684 4 gnd
port 2 nsew
rlabel metal3 s 76656 3859 76754 3957 4 gnd
port 2 nsew
rlabel metal3 s 73976 6586 74074 6684 4 gnd
port 2 nsew
rlabel metal3 s 74333 1862 74431 1960 4 gnd
port 2 nsew
rlabel metal3 s 76582 7355 76680 7453 4 gnd
port 2 nsew
rlabel metal3 s 75581 1862 75679 1960 4 gnd
port 2 nsew
rlabel metal3 s 76829 1862 76927 1960 4 gnd
port 2 nsew
rlabel metal3 s 63987 7557 64085 7655 4 gnd
port 2 nsew
rlabel metal3 s 78963 7557 79061 7655 4 gnd
port 2 nsew
rlabel metal3 s 71837 1862 71935 1960 4 gnd
port 2 nsew
rlabel metal3 s 61680 3859 61778 3957 4 gnd
port 2 nsew
rlabel metal3 s 64349 1862 64447 1960 4 gnd
port 2 nsew
rlabel metal3 s 80573 1862 80671 1960 4 gnd
port 2 nsew
rlabel metal3 s 71475 7557 71573 7655 4 gnd
port 2 nsew
rlabel metal3 s 61491 7557 61589 7655 4 gnd
port 2 nsew
rlabel metal3 s 70589 1862 70687 1960 4 gnd
port 2 nsew
rlabel metal3 s 78968 6586 79066 6684 4 gnd
port 2 nsew
rlabel metal3 s 71594 5793 71692 5891 4 gnd
port 2 nsew
rlabel metal3 s 66483 7557 66581 7655 4 gnd
port 2 nsew
rlabel metal3 s 79078 7355 79176 7453 4 gnd
port 2 nsew
rlabel metal3 s 76586 5793 76684 5891 4 gnd
port 2 nsew
rlabel metal3 s 79325 1862 79423 1960 4 gnd
port 2 nsew
rlabel metal3 s 61610 5793 61708 5891 4 gnd
port 2 nsew
rlabel metal3 s 74090 5793 74188 5891 4 gnd
port 2 nsew
rlabel metal3 s 74160 3859 74258 3957 4 gnd
port 2 nsew
rlabel metal3 s 68979 7557 69077 7655 4 gnd
port 2 nsew
rlabel metal3 s 79152 3859 79250 3957 4 gnd
port 2 nsew
rlabel metal3 s 76472 6586 76570 6684 4 gnd
port 2 nsew
rlabel metal3 s 64106 5793 64204 5891 4 gnd
port 2 nsew
rlabel metal3 s 61853 1862 61951 1960 4 gnd
port 2 nsew
rlabel metal3 s 71590 7355 71688 7453 4 gnd
port 2 nsew
rlabel metal3 s 69098 5793 69196 5891 4 gnd
port 2 nsew
rlabel metal3 s 74086 7355 74184 7453 4 gnd
port 2 nsew
rlabel metal3 s 56513 7973 56611 8071 4 vdd
port 1 nsew
rlabel metal3 s 49005 7023 49103 7121 4 vdd
port 1 nsew
rlabel metal3 s 44138 5793 44236 5891 4 gnd
port 2 nsew
rlabel metal3 s 51626 5793 51724 5891 4 gnd
port 2 nsew
rlabel metal3 s 51626 5471 51724 5569 4 vdd
port 1 nsew
rlabel metal3 s 44024 6586 44122 6684 4 gnd
port 2 nsew
rlabel metal3 s 59114 5471 59212 5569 4 vdd
port 1 nsew
rlabel metal3 s 54110 4633 54208 4731 4 vdd
port 1 nsew
rlabel metal3 s 54122 5471 54220 5569 4 vdd
port 1 nsew
rlabel metal3 s 49025 7973 49123 8071 4 vdd
port 1 nsew
rlabel metal3 s 41517 7023 41615 7121 4 vdd
port 1 nsew
rlabel metal3 s 44013 7023 44111 7121 4 vdd
port 1 nsew
rlabel metal3 s 46634 5471 46732 5569 4 vdd
port 1 nsew
rlabel metal3 s 49130 5793 49228 5891 4 gnd
port 2 nsew
rlabel metal3 s 56493 7023 56591 7121 4 vdd
port 1 nsew
rlabel metal3 s 46634 5793 46732 5891 4 gnd
port 2 nsew
rlabel metal3 s 59110 7355 59208 7453 4 gnd
port 2 nsew
rlabel metal3 s 44126 4633 44224 4731 4 vdd
port 1 nsew
rlabel metal3 s 56499 7557 56597 7655 4 gnd
port 2 nsew
rlabel metal3 s 44208 3859 44306 3957 4 gnd
port 2 nsew
rlabel metal3 s 49016 6586 49114 6684 4 gnd
port 2 nsew
rlabel metal3 s 46509 7023 46607 7121 4 vdd
port 1 nsew
rlabel metal3 s 46704 3859 46802 3957 4 gnd
port 2 nsew
rlabel metal3 s 54118 7355 54216 7453 4 gnd
port 2 nsew
rlabel metal3 s 44138 5471 44236 5569 4 vdd
port 1 nsew
rlabel metal3 s 56614 7355 56712 7453 4 gnd
port 2 nsew
rlabel metal3 s 44381 1862 44479 1960 4 gnd
port 2 nsew
rlabel metal3 s 48125 1862 48223 1960 4 gnd
port 2 nsew
rlabel metal3 s 54008 6586 54106 6684 4 gnd
port 2 nsew
rlabel metal3 s 53997 7023 54095 7121 4 vdd
port 1 nsew
rlabel metal3 s 51521 7973 51619 8071 4 vdd
port 1 nsew
rlabel metal3 s 59102 4633 59200 4731 4 vdd
port 1 nsew
rlabel metal3 s 56504 6586 56602 6684 4 gnd
port 2 nsew
rlabel metal3 s 51614 4633 51712 4731 4 vdd
port 1 nsew
rlabel metal3 s 51501 7023 51599 7121 4 vdd
port 1 nsew
rlabel metal3 s 41528 6586 41626 6684 4 gnd
port 2 nsew
rlabel metal3 s 49130 5471 49228 5569 4 vdd
port 1 nsew
rlabel metal3 s 46529 7973 46627 8071 4 vdd
port 1 nsew
rlabel metal3 s 44033 7973 44131 8071 4 vdd
port 1 nsew
rlabel metal3 s 46877 1862 46975 1960 4 gnd
port 2 nsew
rlabel metal3 s 40637 1862 40735 1960 4 gnd
port 2 nsew
rlabel metal3 s 41537 7973 41635 8071 4 vdd
port 1 nsew
rlabel metal3 s 45629 1862 45727 1960 4 gnd
port 2 nsew
rlabel metal3 s 41642 5471 41740 5569 4 vdd
port 1 nsew
rlabel metal3 s 41642 5793 41740 5891 4 gnd
port 2 nsew
rlabel metal3 s 44134 7355 44232 7453 4 gnd
port 2 nsew
rlabel metal3 s 41885 1862 41983 1960 4 gnd
port 2 nsew
rlabel metal3 s 46515 7557 46613 7655 4 gnd
port 2 nsew
rlabel metal3 s 51622 7355 51720 7453 4 gnd
port 2 nsew
rlabel metal3 s 54365 1862 54463 1960 4 gnd
port 2 nsew
rlabel metal3 s 41712 3859 41810 3957 4 gnd
port 2 nsew
rlabel metal3 s 49200 3859 49298 3957 4 gnd
port 2 nsew
rlabel metal3 s 58989 7023 59087 7121 4 vdd
port 1 nsew
rlabel metal3 s 41630 4633 41728 4731 4 vdd
port 1 nsew
rlabel metal3 s 49011 7557 49109 7655 4 gnd
port 2 nsew
rlabel metal3 s 58995 7557 59093 7655 4 gnd
port 2 nsew
rlabel metal3 s 54017 7973 54115 8071 4 vdd
port 1 nsew
rlabel metal3 s 55613 1862 55711 1960 4 gnd
port 2 nsew
rlabel metal3 s 54122 5793 54220 5891 4 gnd
port 2 nsew
rlabel metal3 s 41638 7355 41736 7453 4 gnd
port 2 nsew
rlabel metal3 s 50621 1862 50719 1960 4 gnd
port 2 nsew
rlabel metal3 s 59357 1862 59455 1960 4 gnd
port 2 nsew
rlabel metal3 s 43133 1862 43231 1960 4 gnd
port 2 nsew
rlabel metal3 s 59000 6586 59098 6684 4 gnd
port 2 nsew
rlabel metal3 s 46622 4633 46720 4731 4 vdd
port 1 nsew
rlabel metal3 s 53117 1862 53215 1960 4 gnd
port 2 nsew
rlabel metal3 s 58109 1862 58207 1960 4 gnd
port 2 nsew
rlabel metal3 s 51512 6586 51610 6684 4 gnd
port 2 nsew
rlabel metal3 s 59184 3859 59282 3957 4 gnd
port 2 nsew
rlabel metal3 s 56688 3859 56786 3957 4 gnd
port 2 nsew
rlabel metal3 s 41523 7557 41621 7655 4 gnd
port 2 nsew
rlabel metal3 s 56606 4633 56704 4731 4 vdd
port 1 nsew
rlabel metal3 s 46520 6586 46618 6684 4 gnd
port 2 nsew
rlabel metal3 s 56861 1862 56959 1960 4 gnd
port 2 nsew
rlabel metal3 s 51507 7557 51605 7655 4 gnd
port 2 nsew
rlabel metal3 s 49126 7355 49224 7453 4 gnd
port 2 nsew
rlabel metal3 s 51696 3859 51794 3957 4 gnd
port 2 nsew
rlabel metal3 s 56618 5471 56716 5569 4 vdd
port 1 nsew
rlabel metal3 s 56618 5793 56716 5891 4 gnd
port 2 nsew
rlabel metal3 s 54003 7557 54101 7655 4 gnd
port 2 nsew
rlabel metal3 s 49373 1862 49471 1960 4 gnd
port 2 nsew
rlabel metal3 s 44019 7557 44117 7655 4 gnd
port 2 nsew
rlabel metal3 s 54192 3859 54290 3957 4 gnd
port 2 nsew
rlabel metal3 s 59009 7973 59107 8071 4 vdd
port 1 nsew
rlabel metal3 s 49118 4633 49216 4731 4 vdd
port 1 nsew
rlabel metal3 s 51869 1862 51967 1960 4 gnd
port 2 nsew
rlabel metal3 s 60605 1862 60703 1960 4 gnd
port 2 nsew
rlabel metal3 s 59114 5793 59212 5891 4 gnd
port 2 nsew
rlabel metal3 s 46630 7355 46728 7453 4 gnd
port 2 nsew
rlabel metal3 s 31646 4633 31744 4731 4 vdd
port 1 nsew
rlabel metal3 s 34142 4633 34240 4731 4 vdd
port 1 nsew
rlabel metal3 s 24413 1862 24511 1960 4 gnd
port 2 nsew
rlabel metal3 s 0 2886 81246 2946 4 sel_1
port 3 nsew
rlabel metal3 s 23165 1862 23263 1960 4 gnd
port 2 nsew
rlabel metal3 s 38141 1862 38239 1960 4 gnd
port 2 nsew
rlabel metal3 s 26561 7973 26659 8071 4 vdd
port 1 nsew
rlabel metal3 s 24240 3859 24338 3957 4 gnd
port 2 nsew
rlabel metal3 s 36545 7973 36643 8071 4 vdd
port 1 nsew
rlabel metal3 s 26541 7023 26639 7121 4 vdd
port 1 nsew
rlabel metal3 s 0 2762 81246 2822 4 sel_2
port 4 nsew
rlabel metal3 s 29162 5793 29260 5891 4 gnd
port 2 nsew
rlabel metal3 s 0 2638 81246 2698 4 sel_3
port 5 nsew
rlabel metal3 s 24065 7973 24163 8071 4 vdd
port 1 nsew
rlabel metal3 s 21662 4633 21760 4731 4 vdd
port 1 nsew
rlabel metal3 s 39216 3859 39314 3957 4 gnd
port 2 nsew
rlabel metal3 s 36650 5793 36748 5891 4 gnd
port 2 nsew
rlabel metal3 s 29057 7973 29155 8071 4 vdd
port 1 nsew
rlabel metal3 s 35645 1862 35743 1960 4 gnd
port 2 nsew
rlabel metal3 s 34029 7023 34127 7121 4 vdd
port 1 nsew
rlabel metal3 s 39021 7023 39119 7121 4 vdd
port 1 nsew
rlabel metal3 s 24170 5793 24268 5891 4 gnd
port 2 nsew
rlabel metal3 s 39142 7355 39240 7453 4 gnd
port 2 nsew
rlabel metal3 s 21569 7973 21667 8071 4 vdd
port 1 nsew
rlabel metal3 s 39041 7973 39139 8071 4 vdd
port 1 nsew
rlabel metal3 s 34154 5471 34252 5569 4 vdd
port 1 nsew
rlabel metal3 s 29162 5471 29260 5569 4 vdd
port 1 nsew
rlabel metal3 s 26547 7557 26645 7655 4 gnd
port 2 nsew
rlabel metal3 s 31658 5793 31756 5891 4 gnd
port 2 nsew
rlabel metal3 s 21674 5793 21772 5891 4 gnd
port 2 nsew
rlabel metal3 s 36638 4633 36736 4731 4 vdd
port 1 nsew
rlabel metal3 s 34049 7973 34147 8071 4 vdd
port 1 nsew
rlabel metal3 s 39146 5471 39244 5569 4 vdd
port 1 nsew
rlabel metal3 s 26654 4633 26752 4731 4 vdd
port 1 nsew
rlabel metal3 s 0 3726 79250 3786 4 s_en
port 6 nsew
rlabel metal3 s 34397 1862 34495 1960 4 gnd
port 2 nsew
rlabel metal3 s 20669 1862 20767 1960 4 gnd
port 2 nsew
rlabel metal3 s 36525 7023 36623 7121 4 vdd
port 1 nsew
rlabel metal3 s 24045 7023 24143 7121 4 vdd
port 1 nsew
rlabel metal3 s 21917 1862 22015 1960 4 gnd
port 2 nsew
rlabel metal3 s 30653 1862 30751 1960 4 gnd
port 2 nsew
rlabel metal3 s 0 9037 81246 9097 4 w_en
port 7 nsew
rlabel metal3 s 39032 6586 39130 6684 4 gnd
port 2 nsew
rlabel metal3 s 21549 7023 21647 7121 4 vdd
port 1 nsew
rlabel metal3 s 29037 7023 29135 7121 4 vdd
port 1 nsew
rlabel metal3 s 26552 6586 26650 6684 4 gnd
port 2 nsew
rlabel metal3 s 24170 5471 24268 5569 4 vdd
port 1 nsew
rlabel metal3 s 39134 4633 39232 4731 4 vdd
port 1 nsew
rlabel metal3 s 36720 3859 36818 3957 4 gnd
port 2 nsew
rlabel metal3 s 34224 3859 34322 3957 4 gnd
port 2 nsew
rlabel metal3 s 31658 5471 31756 5569 4 vdd
port 1 nsew
rlabel metal3 s 31901 1862 31999 1960 4 gnd
port 2 nsew
rlabel metal3 s 29048 6586 29146 6684 4 gnd
port 2 nsew
rlabel metal3 s 21670 7355 21768 7453 4 gnd
port 2 nsew
rlabel metal3 s 0 951 81246 1011 4 p_en_bar
port 8 nsew
rlabel metal3 s 24056 6586 24154 6684 4 gnd
port 2 nsew
rlabel metal3 s 21560 6586 21658 6684 4 gnd
port 2 nsew
rlabel metal3 s 26662 7355 26760 7453 4 gnd
port 2 nsew
rlabel metal3 s 34035 7557 34133 7655 4 gnd
port 2 nsew
rlabel metal3 s 29150 4633 29248 4731 4 vdd
port 1 nsew
rlabel metal3 s 24051 7557 24149 7655 4 gnd
port 2 nsew
rlabel metal3 s 31553 7973 31651 8071 4 vdd
port 1 nsew
rlabel metal3 s 36646 7355 36744 7453 4 gnd
port 2 nsew
rlabel metal3 s 34040 6586 34138 6684 4 gnd
port 2 nsew
rlabel metal3 s 21744 3859 21842 3957 4 gnd
port 2 nsew
rlabel metal3 s 24166 7355 24264 7453 4 gnd
port 2 nsew
rlabel metal3 s 31539 7557 31637 7655 4 gnd
port 2 nsew
rlabel metal3 s 31728 3859 31826 3957 4 gnd
port 2 nsew
rlabel metal3 s 24158 4633 24256 4731 4 vdd
port 1 nsew
rlabel metal3 s 29405 1862 29503 1960 4 gnd
port 2 nsew
rlabel metal3 s 29043 7557 29141 7655 4 gnd
port 2 nsew
rlabel metal3 s 26736 3859 26834 3957 4 gnd
port 2 nsew
rlabel metal3 s 39027 7557 39125 7655 4 gnd
port 2 nsew
rlabel metal3 s 33149 1862 33247 1960 4 gnd
port 2 nsew
rlabel metal3 s 34154 5793 34252 5891 4 gnd
port 2 nsew
rlabel metal3 s 28157 1862 28255 1960 4 gnd
port 2 nsew
rlabel metal3 s 0 3010 81246 3070 4 sel_0
port 9 nsew
rlabel metal3 s 31533 7023 31631 7121 4 vdd
port 1 nsew
rlabel metal3 s 29232 3859 29330 3957 4 gnd
port 2 nsew
rlabel metal3 s 26909 1862 27007 1960 4 gnd
port 2 nsew
rlabel metal3 s 31654 7355 31752 7453 4 gnd
port 2 nsew
rlabel metal3 s 21555 7557 21653 7655 4 gnd
port 2 nsew
rlabel metal3 s 36893 1862 36991 1960 4 gnd
port 2 nsew
rlabel metal3 s 36650 5471 36748 5569 4 vdd
port 1 nsew
rlabel metal3 s 36531 7557 36629 7655 4 gnd
port 2 nsew
rlabel metal3 s 26666 5471 26764 5569 4 vdd
port 1 nsew
rlabel metal3 s 26666 5793 26764 5891 4 gnd
port 2 nsew
rlabel metal3 s 29158 7355 29256 7453 4 gnd
port 2 nsew
rlabel metal3 s 25661 1862 25759 1960 4 gnd
port 2 nsew
rlabel metal3 s 31544 6586 31642 6684 4 gnd
port 2 nsew
rlabel metal3 s 34150 7355 34248 7453 4 gnd
port 2 nsew
rlabel metal3 s 21674 5471 21772 5569 4 vdd
port 1 nsew
rlabel metal3 s 39146 5793 39244 5891 4 gnd
port 2 nsew
rlabel metal3 s 39389 1862 39487 1960 4 gnd
port 2 nsew
rlabel metal3 s 36536 6586 36634 6684 4 gnd
port 2 nsew
rlabel metal3 s 6573 7023 6671 7121 4 vdd
port 1 nsew
rlabel metal3 s 9437 1862 9535 1960 4 gnd
port 2 nsew
rlabel metal3 s 6941 1862 7039 1960 4 gnd
port 2 nsew
rlabel metal3 s 4088 6586 4186 6684 4 gnd
port 2 nsew
rlabel metal3 s 1776 3859 1874 3957 4 gnd
port 2 nsew
rlabel metal3 s 4202 5793 4300 5891 4 gnd
port 2 nsew
rlabel metal3 s 3197 1862 3295 1960 4 gnd
port 2 nsew
rlabel metal3 s 14061 7023 14159 7121 4 vdd
port 1 nsew
rlabel metal3 s 5693 1862 5791 1960 4 gnd
port 2 nsew
rlabel metal3 s 6694 7355 6792 7453 4 gnd
port 2 nsew
rlabel metal3 s 16752 3859 16850 3957 4 gnd
port 2 nsew
rlabel metal3 s 16568 6586 16666 6684 4 gnd
port 2 nsew
rlabel metal3 s 14067 7557 14165 7655 4 gnd
port 2 nsew
rlabel metal3 s 8189 1862 8287 1960 4 gnd
port 2 nsew
rlabel metal3 s 1601 7973 1699 8071 4 vdd
port 1 nsew
rlabel metal3 s 11571 7557 11669 7655 4 gnd
port 2 nsew
rlabel metal3 s 4077 7023 4175 7121 4 vdd
port 1 nsew
rlabel metal3 s 16563 7557 16661 7655 4 gnd
port 2 nsew
rlabel metal3 s 1581 7023 1679 7121 4 vdd
port 1 nsew
rlabel metal3 s 1587 7557 1685 7655 4 gnd
port 2 nsew
rlabel metal3 s 1706 5793 1804 5891 4 gnd
port 2 nsew
rlabel metal3 s 9075 7557 9173 7655 4 gnd
port 2 nsew
rlabel metal3 s 11686 7355 11784 7453 4 gnd
port 2 nsew
rlabel metal3 s 9264 3859 9362 3957 4 gnd
port 2 nsew
rlabel metal3 s 11760 3859 11858 3957 4 gnd
port 2 nsew
rlabel metal3 s 11690 5471 11788 5569 4 vdd
port 1 nsew
rlabel metal3 s 11690 5793 11788 5891 4 gnd
port 2 nsew
rlabel metal3 s 14081 7973 14179 8071 4 vdd
port 1 nsew
rlabel metal3 s 16925 1862 17023 1960 4 gnd
port 2 nsew
rlabel metal3 s 9182 4633 9280 4731 4 vdd
port 1 nsew
rlabel metal3 s 15677 1862 15775 1960 4 gnd
port 2 nsew
rlabel metal3 s 19073 7973 19171 8071 4 vdd
port 1 nsew
rlabel metal3 s 6698 5793 6796 5891 4 gnd
port 2 nsew
rlabel metal3 s 11933 1862 12031 1960 4 gnd
port 2 nsew
rlabel metal3 s 1702 7355 1800 7453 4 gnd
port 2 nsew
rlabel metal3 s 14429 1862 14527 1960 4 gnd
port 2 nsew
rlabel metal3 s 14186 5471 14284 5569 4 vdd
port 1 nsew
rlabel metal3 s 1694 4633 1792 4731 4 vdd
port 1 nsew
rlabel metal3 s 6593 7973 6691 8071 4 vdd
port 1 nsew
rlabel metal3 s 16670 4633 16768 4731 4 vdd
port 1 nsew
rlabel metal3 s 18173 1862 18271 1960 4 gnd
port 2 nsew
rlabel metal3 s 1706 5471 1804 5569 4 vdd
port 1 nsew
rlabel metal3 s 16577 7973 16675 8071 4 vdd
port 1 nsew
rlabel metal3 s 9194 5471 9292 5569 4 vdd
port 1 nsew
rlabel metal3 s 11678 4633 11776 4731 4 vdd
port 1 nsew
rlabel metal3 s 19166 4633 19264 4731 4 vdd
port 1 nsew
rlabel metal3 s 10685 1862 10783 1960 4 gnd
port 2 nsew
rlabel metal3 s 14182 7355 14280 7453 4 gnd
port 2 nsew
rlabel metal3 s 6584 6586 6682 6684 4 gnd
port 2 nsew
rlabel metal3 s 9089 7973 9187 8071 4 vdd
port 1 nsew
rlabel metal3 s 14186 5793 14284 5891 4 gnd
port 2 nsew
rlabel metal3 s 19174 7355 19272 7453 4 gnd
port 2 nsew
rlabel metal3 s 9190 7355 9288 7453 4 gnd
port 2 nsew
rlabel metal3 s 4272 3859 4370 3957 4 gnd
port 2 nsew
rlabel metal3 s 13181 1862 13279 1960 4 gnd
port 2 nsew
rlabel metal3 s 14072 6586 14170 6684 4 gnd
port 2 nsew
rlabel metal3 s 9069 7023 9167 7121 4 vdd
port 1 nsew
rlabel metal3 s -49 8416 49 8514 4 vdd
port 1 nsew
rlabel metal3 s 4202 5471 4300 5569 4 vdd
port 1 nsew
rlabel metal3 s 4445 1862 4543 1960 4 gnd
port 2 nsew
rlabel metal3 s 19421 1862 19519 1960 4 gnd
port 2 nsew
rlabel metal3 s 11585 7973 11683 8071 4 vdd
port 1 nsew
rlabel metal3 s 4198 7355 4296 7453 4 gnd
port 2 nsew
rlabel metal3 s 6768 3859 6866 3957 4 gnd
port 2 nsew
rlabel metal3 s 19059 7557 19157 7655 4 gnd
port 2 nsew
rlabel metal3 s 19053 7023 19151 7121 4 vdd
port 1 nsew
rlabel metal3 s 4083 7557 4181 7655 4 gnd
port 2 nsew
rlabel metal3 s 6698 5471 6796 5569 4 vdd
port 1 nsew
rlabel metal3 s 16682 5471 16780 5569 4 vdd
port 1 nsew
rlabel metal3 s 19178 5471 19276 5569 4 vdd
port 1 nsew
rlabel metal3 s 4097 7973 4195 8071 4 vdd
port 1 nsew
rlabel metal3 s 9194 5793 9292 5891 4 gnd
port 2 nsew
rlabel metal3 s 1949 1862 2047 1960 4 gnd
port 2 nsew
rlabel metal3 s 1592 6586 1690 6684 4 gnd
port 2 nsew
rlabel metal3 s 14256 3859 14354 3957 4 gnd
port 2 nsew
rlabel metal3 s 4190 4633 4288 4731 4 vdd
port 1 nsew
rlabel metal3 s 14174 4633 14272 4731 4 vdd
port 1 nsew
rlabel metal3 s 16557 7023 16655 7121 4 vdd
port 1 nsew
rlabel metal3 s 16678 7355 16776 7453 4 gnd
port 2 nsew
rlabel metal3 s 16682 5793 16780 5891 4 gnd
port 2 nsew
rlabel metal3 s 19248 3859 19346 3957 4 gnd
port 2 nsew
rlabel metal3 s 19178 5793 19276 5891 4 gnd
port 2 nsew
rlabel metal3 s 9080 6586 9178 6684 4 gnd
port 2 nsew
rlabel metal3 s 11565 7023 11663 7121 4 vdd
port 1 nsew
rlabel metal3 s 19064 6586 19162 6684 4 gnd
port 2 nsew
rlabel metal3 s 6686 4633 6784 4731 4 vdd
port 1 nsew
rlabel metal3 s 6579 7557 6677 7655 4 gnd
port 2 nsew
rlabel metal3 s -49 9536 49 9634 4 gnd
port 2 nsew
rlabel metal3 s 11576 6586 11674 6684 4 gnd
port 2 nsew
rlabel metal3 s 9868 313 9966 411 4 vdd
port 1 nsew
rlabel metal3 s 34828 313 34926 411 4 vdd
port 1 nsew
rlabel metal3 s 38572 313 38670 411 4 vdd
port 1 nsew
rlabel metal3 s 4014 313 4112 411 4 vdd
port 1 nsew
rlabel metal3 s 31084 313 31182 411 4 vdd
port 1 nsew
rlabel metal3 s 33580 313 33678 411 4 vdd
port 1 nsew
rlabel metal3 s 29836 313 29934 411 4 vdd
port 1 nsew
rlabel metal3 s 16108 313 16206 411 4 vdd
port 1 nsew
rlabel metal3 s 7372 313 7470 411 4 vdd
port 1 nsew
rlabel metal3 s 28974 313 29072 411 4 vdd
port 1 nsew
rlabel metal3 s 13612 313 13710 411 4 vdd
port 1 nsew
rlabel metal3 s 31470 313 31568 411 4 vdd
port 1 nsew
rlabel metal3 s 38958 313 39056 411 4 vdd
port 1 nsew
rlabel metal3 s 24844 313 24942 411 4 vdd
port 1 nsew
rlabel metal3 s 19852 313 19950 411 4 vdd
port 1 nsew
rlabel metal3 s 22734 313 22832 411 4 vdd
port 1 nsew
rlabel metal3 s 17356 313 17454 411 4 vdd
port 1 nsew
rlabel metal3 s 7758 313 7856 411 4 vdd
port 1 nsew
rlabel metal3 s 18604 313 18702 411 4 vdd
port 1 nsew
rlabel metal3 s 22348 313 22446 411 4 vdd
port 1 nsew
rlabel metal3 s 40206 313 40304 411 4 vdd
port 1 nsew
rlabel metal3 s 17742 313 17840 411 4 vdd
port 1 nsew
rlabel metal3 s 5262 313 5360 411 4 vdd
port 1 nsew
rlabel metal3 s 25230 313 25328 411 4 vdd
port 1 nsew
rlabel metal3 s 8620 313 8718 411 4 vdd
port 1 nsew
rlabel metal3 s 35214 313 35312 411 4 vdd
port 1 nsew
rlabel metal3 s 32332 313 32430 411 4 vdd
port 1 nsew
rlabel metal3 s 2380 313 2478 411 4 vdd
port 1 nsew
rlabel metal3 s 27726 313 27824 411 4 vdd
port 1 nsew
rlabel metal3 s 23982 313 24080 411 4 vdd
port 1 nsew
rlabel metal3 s 13998 313 14096 411 4 vdd
port 1 nsew
rlabel metal3 s 18990 313 19088 411 4 vdd
port 1 nsew
rlabel metal3 s 21100 313 21198 411 4 vdd
port 1 nsew
rlabel metal3 s 36462 313 36560 411 4 vdd
port 1 nsew
rlabel metal3 s 26092 313 26190 411 4 vdd
port 1 nsew
rlabel metal3 s 4876 313 4974 411 4 vdd
port 1 nsew
rlabel metal3 s 21486 313 21584 411 4 vdd
port 1 nsew
rlabel metal3 s 33966 313 34064 411 4 vdd
port 1 nsew
rlabel metal3 s 1132 313 1230 411 4 vdd
port 1 nsew
rlabel metal3 s 1518 313 1616 411 4 vdd
port 1 nsew
rlabel metal3 s 3628 313 3726 411 4 vdd
port 1 nsew
rlabel metal3 s 36076 313 36174 411 4 vdd
port 1 nsew
rlabel metal3 s 2766 313 2864 411 4 vdd
port 1 nsew
rlabel metal3 s 6124 313 6222 411 4 vdd
port 1 nsew
rlabel metal3 s 11116 313 11214 411 4 vdd
port 1 nsew
rlabel metal3 s 37710 313 37808 411 4 vdd
port 1 nsew
rlabel metal3 s 28588 313 28686 411 4 vdd
port 1 nsew
rlabel metal3 s 10254 313 10352 411 4 vdd
port 1 nsew
rlabel metal3 s 12750 313 12848 411 4 vdd
port 1 nsew
rlabel metal3 s 30222 313 30320 411 4 vdd
port 1 nsew
rlabel metal3 s 16494 313 16592 411 4 vdd
port 1 nsew
rlabel metal3 s 11502 313 11600 411 4 vdd
port 1 nsew
rlabel metal3 s 6510 313 6608 411 4 vdd
port 1 nsew
rlabel metal3 s 23596 313 23694 411 4 vdd
port 1 nsew
rlabel metal3 s 32718 313 32816 411 4 vdd
port 1 nsew
rlabel metal3 s 20238 313 20336 411 4 vdd
port 1 nsew
rlabel metal3 s 12364 313 12462 411 4 vdd
port 1 nsew
rlabel metal3 s 39820 313 39918 411 4 vdd
port 1 nsew
rlabel metal3 s 26478 313 26576 411 4 vdd
port 1 nsew
rlabel metal3 s 27340 313 27438 411 4 vdd
port 1 nsew
rlabel metal3 s 14860 313 14958 411 4 vdd
port 1 nsew
rlabel metal3 s 37324 313 37422 411 4 vdd
port 1 nsew
rlabel metal3 s 9006 313 9104 411 4 vdd
port 1 nsew
rlabel metal3 s 15246 313 15344 411 4 vdd
port 1 nsew
rlabel metal3 s 80142 313 80240 411 4 vdd
port 1 nsew
rlabel metal3 s 48942 313 49040 411 4 vdd
port 1 nsew
rlabel metal3 s 50190 313 50288 411 4 vdd
port 1 nsew
rlabel metal3 s 78894 313 78992 411 4 vdd
port 1 nsew
rlabel metal3 s 53934 313 54032 411 4 vdd
port 1 nsew
rlabel metal3 s 57678 313 57776 411 4 vdd
port 1 nsew
rlabel metal3 s 61422 313 61520 411 4 vdd
port 1 nsew
rlabel metal3 s 63918 313 64016 411 4 vdd
port 1 nsew
rlabel metal3 s 77646 313 77744 411 4 vdd
port 1 nsew
rlabel metal3 s 58540 313 58638 411 4 vdd
port 1 nsew
rlabel metal3 s 71406 313 71504 411 4 vdd
port 1 nsew
rlabel metal3 s 41068 313 41166 411 4 vdd
port 1 nsew
rlabel metal3 s 51052 313 51150 411 4 vdd
port 1 nsew
rlabel metal3 s 77260 313 77358 411 4 vdd
port 1 nsew
rlabel metal3 s 59788 313 59886 411 4 vdd
port 1 nsew
rlabel metal3 s 73516 313 73614 411 4 vdd
port 1 nsew
rlabel metal3 s 78508 313 78606 411 4 vdd
port 1 nsew
rlabel metal3 s 66414 313 66512 411 4 vdd
port 1 nsew
rlabel metal3 s 56044 313 56142 411 4 vdd
port 1 nsew
rlabel metal3 s 56430 313 56528 411 4 vdd
port 1 nsew
rlabel metal3 s 74764 313 74862 411 4 vdd
port 1 nsew
rlabel metal3 s 67276 313 67374 411 4 vdd
port 1 nsew
rlabel metal3 s 42316 313 42414 411 4 vdd
port 1 nsew
rlabel metal3 s 43950 313 44048 411 4 vdd
port 1 nsew
rlabel metal3 s 71020 313 71118 411 4 vdd
port 1 nsew
rlabel metal3 s 47694 313 47792 411 4 vdd
port 1 nsew
rlabel metal3 s 46060 313 46158 411 4 vdd
port 1 nsew
rlabel metal3 s 69772 313 69870 411 4 vdd
port 1 nsew
rlabel metal3 s 54796 313 54894 411 4 vdd
port 1 nsew
rlabel metal3 s 79756 313 79854 411 4 vdd
port 1 nsew
rlabel metal3 s 68910 313 69008 411 4 vdd
port 1 nsew
rlabel metal3 s 76012 313 76110 411 4 vdd
port 1 nsew
rlabel metal3 s 55182 313 55280 411 4 vdd
port 1 nsew
rlabel metal3 s 52300 313 52398 411 4 vdd
port 1 nsew
rlabel metal3 s 65166 313 65264 411 4 vdd
port 1 nsew
rlabel metal3 s 62284 313 62382 411 4 vdd
port 1 nsew
rlabel metal3 s 66028 313 66126 411 4 vdd
port 1 nsew
rlabel metal3 s 45198 313 45296 411 4 vdd
port 1 nsew
rlabel metal3 s 52686 313 52784 411 4 vdd
port 1 nsew
rlabel metal3 s 58926 313 59024 411 4 vdd
port 1 nsew
rlabel metal3 s 46446 313 46544 411 4 vdd
port 1 nsew
rlabel metal3 s 62670 313 62768 411 4 vdd
port 1 nsew
rlabel metal3 s 43564 313 43662 411 4 vdd
port 1 nsew
rlabel metal3 s 41454 313 41552 411 4 vdd
port 1 nsew
rlabel metal3 s 73902 313 74000 411 4 vdd
port 1 nsew
rlabel metal3 s 72654 313 72752 411 4 vdd
port 1 nsew
rlabel metal3 s 47308 313 47406 411 4 vdd
port 1 nsew
rlabel metal3 s 67662 313 67760 411 4 vdd
port 1 nsew
rlabel metal3 s 61036 313 61134 411 4 vdd
port 1 nsew
rlabel metal3 s 51438 313 51536 411 4 vdd
port 1 nsew
rlabel metal3 s 60174 313 60272 411 4 vdd
port 1 nsew
rlabel metal3 s 48556 313 48654 411 4 vdd
port 1 nsew
rlabel metal3 s 68524 313 68622 411 4 vdd
port 1 nsew
rlabel metal3 s 72268 313 72366 411 4 vdd
port 1 nsew
rlabel metal3 s 63532 313 63630 411 4 vdd
port 1 nsew
rlabel metal3 s 81004 313 81102 411 4 vdd
port 1 nsew
rlabel metal3 s 76398 313 76496 411 4 vdd
port 1 nsew
rlabel metal3 s 49804 313 49902 411 4 vdd
port 1 nsew
rlabel metal3 s 44812 313 44910 411 4 vdd
port 1 nsew
rlabel metal3 s 42702 313 42800 411 4 vdd
port 1 nsew
rlabel metal3 s 64780 313 64878 411 4 vdd
port 1 nsew
rlabel metal3 s 57292 313 57390 411 4 vdd
port 1 nsew
rlabel metal3 s 53548 313 53646 411 4 vdd
port 1 nsew
rlabel metal3 s 70158 313 70256 411 4 vdd
port 1 nsew
rlabel metal3 s 75150 313 75248 411 4 vdd
port 1 nsew
rlabel metal2 s 1360 9301 1388 9329 4 bank_wmask_0
port 10 nsew
rlabel metal2 s 21328 9301 21356 9329 4 bank_wmask_1
port 11 nsew
rlabel metal2 s 41296 9301 41324 9329 4 bank_wmask_2
port 12 nsew
rlabel metal2 s 61264 9301 61292 9329 4 bank_wmask_3
port 13 nsew
rlabel metal1 s 41409 8085 60753 8119 4 wdriver_sel_2
port 14 nsew
rlabel metal1 s 61377 8085 80721 8119 4 wdriver_sel_3
port 15 nsew
rlabel metal1 s 41565 8153 41625 8209 4 din_16
port 16 nsew
rlabel metal1 s 44061 8153 44121 8209 4 din_17
port 17 nsew
rlabel metal1 s 46557 8153 46617 8209 4 din_18
port 18 nsew
rlabel metal1 s 49053 8153 49113 8209 4 din_19
port 19 nsew
rlabel metal1 s 51549 8153 51609 8209 4 din_20
port 20 nsew
rlabel metal1 s 54045 8153 54105 8209 4 din_21
port 21 nsew
rlabel metal1 s 56541 8153 56601 8209 4 din_22
port 22 nsew
rlabel metal1 s 59037 8153 59097 8209 4 din_23
port 23 nsew
rlabel metal1 s 61533 8153 61593 8209 4 din_24
port 24 nsew
rlabel metal1 s 64029 8153 64089 8209 4 din_25
port 25 nsew
rlabel metal1 s 66525 8153 66585 8209 4 din_26
port 26 nsew
rlabel metal1 s 69021 8153 69081 8209 4 din_27
port 27 nsew
rlabel metal1 s 71517 8153 71577 8209 4 din_28
port 28 nsew
rlabel metal1 s 74013 8153 74073 8209 4 din_29
port 29 nsew
rlabel metal1 s 76509 8153 76569 8209 4 din_30
port 30 nsew
rlabel metal1 s 79005 8153 79065 8209 4 din_31
port 31 nsew
rlabel metal1 s 41414 5696 41460 5950 4 dout_16
port 32 nsew
rlabel metal1 s 43910 5696 43956 5950 4 dout_17
port 33 nsew
rlabel metal1 s 46406 5696 46452 5950 4 dout_18
port 34 nsew
rlabel metal1 s 48902 5696 48948 5950 4 dout_19
port 35 nsew
rlabel metal1 s 51398 5696 51444 5950 4 dout_20
port 36 nsew
rlabel metal1 s 53894 5696 53940 5950 4 dout_21
port 37 nsew
rlabel metal1 s 56390 5696 56436 5950 4 dout_22
port 38 nsew
rlabel metal1 s 58886 5696 58932 5950 4 dout_23
port 39 nsew
rlabel metal1 s 61382 5696 61428 5950 4 dout_24
port 40 nsew
rlabel metal1 s 63878 5696 63924 5950 4 dout_25
port 41 nsew
rlabel metal1 s 66374 5696 66420 5950 4 dout_26
port 42 nsew
rlabel metal1 s 68870 5696 68916 5950 4 dout_27
port 43 nsew
rlabel metal1 s 71366 5696 71412 5950 4 dout_28
port 44 nsew
rlabel metal1 s 73862 5696 73908 5950 4 dout_29
port 45 nsew
rlabel metal1 s 76358 5696 76404 5950 4 dout_30
port 46 nsew
rlabel metal1 s 78854 5696 78900 5950 4 dout_31
port 47 nsew
rlabel metal1 s 31581 8153 31641 8209 4 din_12
port 48 nsew
rlabel metal1 s 34077 8153 34137 8209 4 din_13
port 49 nsew
rlabel metal1 s 1478 5696 1524 5950 4 dout_0
port 50 nsew
rlabel metal1 s 3974 5696 4020 5950 4 dout_1
port 51 nsew
rlabel metal1 s 6470 5696 6516 5950 4 dout_2
port 52 nsew
rlabel metal1 s 8966 5696 9012 5950 4 dout_3
port 53 nsew
rlabel metal1 s 11462 5696 11508 5950 4 dout_4
port 54 nsew
rlabel metal1 s 13958 5696 14004 5950 4 dout_5
port 55 nsew
rlabel metal1 s 16454 5696 16500 5950 4 dout_6
port 56 nsew
rlabel metal1 s 18950 5696 18996 5950 4 dout_7
port 57 nsew
rlabel metal1 s 21446 5696 21492 5950 4 dout_8
port 58 nsew
rlabel metal1 s 23942 5696 23988 5950 4 dout_9
port 59 nsew
rlabel metal1 s 26438 5696 26484 5950 4 dout_10
port 60 nsew
rlabel metal1 s 28934 5696 28980 5950 4 dout_11
port 61 nsew
rlabel metal1 s 31430 5696 31476 5950 4 dout_12
port 62 nsew
rlabel metal1 s 33926 5696 33972 5950 4 dout_13
port 63 nsew
rlabel metal1 s 36422 5696 36468 5950 4 dout_14
port 64 nsew
rlabel metal1 s 38918 5696 38964 5950 4 dout_15
port 65 nsew
rlabel metal1 s 36573 8153 36633 8209 4 din_14
port 66 nsew
rlabel metal1 s 39069 8153 39129 8209 4 din_15
port 67 nsew
rlabel metal1 s 1473 8085 20817 8119 4 wdriver_sel_0
port 68 nsew
rlabel metal1 s 21441 8085 40785 8119 4 wdriver_sel_1
port 69 nsew
rlabel metal1 s 1629 8153 1689 8209 4 din_0
port 70 nsew
rlabel metal1 s 4125 8153 4185 8209 4 din_1
port 71 nsew
rlabel metal1 s 6621 8153 6681 8209 4 din_2
port 72 nsew
rlabel metal1 s 9117 8153 9177 8209 4 din_3
port 73 nsew
rlabel metal1 s 11613 8153 11673 8209 4 din_4
port 74 nsew
rlabel metal1 s 14109 8153 14169 8209 4 din_5
port 75 nsew
rlabel metal1 s 16605 8153 16665 8209 4 din_6
port 76 nsew
rlabel metal1 s 19101 8153 19161 8209 4 din_7
port 77 nsew
rlabel metal1 s 21597 8153 21657 8209 4 din_8
port 78 nsew
rlabel metal1 s 24093 8153 24153 8209 4 din_9
port 79 nsew
rlabel metal1 s 26589 8153 26649 8209 4 din_10
port 80 nsew
rlabel metal1 s 29085 8153 29145 8209 4 din_11
port 81 nsew
rlabel metal1 s 1280 252 1308 1006 4 rbl_bl
port 82 nsew
rlabel metal1 s 816 252 844 1006 4 rbl_br
port 83 nsew
rlabel metal1 s 1440 252 1468 1006 4 bl_0
port 84 nsew
rlabel metal1 s 1904 252 1932 1006 4 br_0
port 85 nsew
rlabel metal1 s 2528 252 2556 1006 4 bl_1
port 86 nsew
rlabel metal1 s 2064 252 2092 1006 4 br_1
port 87 nsew
rlabel metal1 s 2688 252 2716 1006 4 bl_2
port 88 nsew
rlabel metal1 s 3152 252 3180 1006 4 br_2
port 89 nsew
rlabel metal1 s 3776 252 3804 1006 4 bl_3
port 90 nsew
rlabel metal1 s 3312 252 3340 1006 4 br_3
port 91 nsew
rlabel metal1 s 3936 252 3964 1006 4 bl_4
port 92 nsew
rlabel metal1 s 4400 252 4428 1006 4 br_4
port 93 nsew
rlabel metal1 s 5024 252 5052 1006 4 bl_5
port 94 nsew
rlabel metal1 s 4560 252 4588 1006 4 br_5
port 95 nsew
rlabel metal1 s 5184 252 5212 1006 4 bl_6
port 96 nsew
rlabel metal1 s 5648 252 5676 1006 4 br_6
port 97 nsew
rlabel metal1 s 6272 252 6300 1006 4 bl_7
port 98 nsew
rlabel metal1 s 5808 252 5836 1006 4 br_7
port 99 nsew
rlabel metal1 s 6432 252 6460 1006 4 bl_8
port 100 nsew
rlabel metal1 s 6896 252 6924 1006 4 br_8
port 101 nsew
rlabel metal1 s 7520 252 7548 1006 4 bl_9
port 102 nsew
rlabel metal1 s 7056 252 7084 1006 4 br_9
port 103 nsew
rlabel metal1 s 7680 252 7708 1006 4 bl_10
port 104 nsew
rlabel metal1 s 8144 252 8172 1006 4 br_10
port 105 nsew
rlabel metal1 s 8768 252 8796 1006 4 bl_11
port 106 nsew
rlabel metal1 s 8304 252 8332 1006 4 br_11
port 107 nsew
rlabel metal1 s 8928 252 8956 1006 4 bl_12
port 108 nsew
rlabel metal1 s 9392 252 9420 1006 4 br_12
port 109 nsew
rlabel metal1 s 10016 252 10044 1006 4 bl_13
port 110 nsew
rlabel metal1 s 9552 252 9580 1006 4 br_13
port 111 nsew
rlabel metal1 s 10176 252 10204 1006 4 bl_14
port 112 nsew
rlabel metal1 s 10640 252 10668 1006 4 br_14
port 113 nsew
rlabel metal1 s 11264 252 11292 1006 4 bl_15
port 114 nsew
rlabel metal1 s 10800 252 10828 1006 4 br_15
port 115 nsew
rlabel metal1 s 11424 252 11452 1006 4 bl_16
port 116 nsew
rlabel metal1 s 11888 252 11916 1006 4 br_16
port 117 nsew
rlabel metal1 s 12512 252 12540 1006 4 bl_17
port 118 nsew
rlabel metal1 s 12048 252 12076 1006 4 br_17
port 119 nsew
rlabel metal1 s 12672 252 12700 1006 4 bl_18
port 120 nsew
rlabel metal1 s 13136 252 13164 1006 4 br_18
port 121 nsew
rlabel metal1 s 13760 252 13788 1006 4 bl_19
port 122 nsew
rlabel metal1 s 13296 252 13324 1006 4 br_19
port 123 nsew
rlabel metal1 s 13920 252 13948 1006 4 bl_20
port 124 nsew
rlabel metal1 s 14384 252 14412 1006 4 br_20
port 125 nsew
rlabel metal1 s 15008 252 15036 1006 4 bl_21
port 126 nsew
rlabel metal1 s 14544 252 14572 1006 4 br_21
port 127 nsew
rlabel metal1 s 15168 252 15196 1006 4 bl_22
port 128 nsew
rlabel metal1 s 15632 252 15660 1006 4 br_22
port 129 nsew
rlabel metal1 s 16256 252 16284 1006 4 bl_23
port 130 nsew
rlabel metal1 s 15792 252 15820 1006 4 br_23
port 131 nsew
rlabel metal1 s 16416 252 16444 1006 4 bl_24
port 132 nsew
rlabel metal1 s 16880 252 16908 1006 4 br_24
port 133 nsew
rlabel metal1 s 17504 252 17532 1006 4 bl_25
port 134 nsew
rlabel metal1 s 17040 252 17068 1006 4 br_25
port 135 nsew
rlabel metal1 s 17664 252 17692 1006 4 bl_26
port 136 nsew
rlabel metal1 s 18128 252 18156 1006 4 br_26
port 137 nsew
rlabel metal1 s 18752 252 18780 1006 4 bl_27
port 138 nsew
rlabel metal1 s 18288 252 18316 1006 4 br_27
port 139 nsew
rlabel metal1 s 18912 252 18940 1006 4 bl_28
port 140 nsew
rlabel metal1 s 19376 252 19404 1006 4 br_28
port 141 nsew
rlabel metal1 s 20000 252 20028 1006 4 bl_29
port 142 nsew
rlabel metal1 s 19536 252 19564 1006 4 br_29
port 143 nsew
rlabel metal1 s 20160 252 20188 1006 4 bl_30
port 144 nsew
rlabel metal1 s 20624 252 20652 1006 4 br_30
port 145 nsew
rlabel metal1 s 20784 252 20812 1006 4 br_31
port 146 nsew
rlabel metal1 s 21248 252 21276 1006 4 bl_31
port 147 nsew
rlabel metal1 s 21408 252 21436 1006 4 bl_32
port 148 nsew
rlabel metal1 s 21872 252 21900 1006 4 br_32
port 149 nsew
rlabel metal1 s 22496 252 22524 1006 4 bl_33
port 150 nsew
rlabel metal1 s 22032 252 22060 1006 4 br_33
port 151 nsew
rlabel metal1 s 22656 252 22684 1006 4 bl_34
port 152 nsew
rlabel metal1 s 23120 252 23148 1006 4 br_34
port 153 nsew
rlabel metal1 s 23744 252 23772 1006 4 bl_35
port 154 nsew
rlabel metal1 s 23280 252 23308 1006 4 br_35
port 155 nsew
rlabel metal1 s 23904 252 23932 1006 4 bl_36
port 156 nsew
rlabel metal1 s 24368 252 24396 1006 4 br_36
port 157 nsew
rlabel metal1 s 24992 252 25020 1006 4 bl_37
port 158 nsew
rlabel metal1 s 24528 252 24556 1006 4 br_37
port 159 nsew
rlabel metal1 s 25152 252 25180 1006 4 bl_38
port 160 nsew
rlabel metal1 s 25616 252 25644 1006 4 br_38
port 161 nsew
rlabel metal1 s 26240 252 26268 1006 4 bl_39
port 162 nsew
rlabel metal1 s 25776 252 25804 1006 4 br_39
port 163 nsew
rlabel metal1 s 26400 252 26428 1006 4 bl_40
port 164 nsew
rlabel metal1 s 26864 252 26892 1006 4 br_40
port 165 nsew
rlabel metal1 s 27488 252 27516 1006 4 bl_41
port 166 nsew
rlabel metal1 s 27024 252 27052 1006 4 br_41
port 167 nsew
rlabel metal1 s 27648 252 27676 1006 4 bl_42
port 168 nsew
rlabel metal1 s 28112 252 28140 1006 4 br_42
port 169 nsew
rlabel metal1 s 28736 252 28764 1006 4 bl_43
port 170 nsew
rlabel metal1 s 28272 252 28300 1006 4 br_43
port 171 nsew
rlabel metal1 s 28896 252 28924 1006 4 bl_44
port 172 nsew
rlabel metal1 s 29360 252 29388 1006 4 br_44
port 173 nsew
rlabel metal1 s 29984 252 30012 1006 4 bl_45
port 174 nsew
rlabel metal1 s 29520 252 29548 1006 4 br_45
port 175 nsew
rlabel metal1 s 30144 252 30172 1006 4 bl_46
port 176 nsew
rlabel metal1 s 30608 252 30636 1006 4 br_46
port 177 nsew
rlabel metal1 s 31232 252 31260 1006 4 bl_47
port 178 nsew
rlabel metal1 s 30768 252 30796 1006 4 br_47
port 179 nsew
rlabel metal1 s 31392 252 31420 1006 4 bl_48
port 180 nsew
rlabel metal1 s 31856 252 31884 1006 4 br_48
port 181 nsew
rlabel metal1 s 32480 252 32508 1006 4 bl_49
port 182 nsew
rlabel metal1 s 32016 252 32044 1006 4 br_49
port 183 nsew
rlabel metal1 s 32640 252 32668 1006 4 bl_50
port 184 nsew
rlabel metal1 s 33104 252 33132 1006 4 br_50
port 185 nsew
rlabel metal1 s 33728 252 33756 1006 4 bl_51
port 186 nsew
rlabel metal1 s 33264 252 33292 1006 4 br_51
port 187 nsew
rlabel metal1 s 33888 252 33916 1006 4 bl_52
port 188 nsew
rlabel metal1 s 34352 252 34380 1006 4 br_52
port 189 nsew
rlabel metal1 s 34976 252 35004 1006 4 bl_53
port 190 nsew
rlabel metal1 s 34512 252 34540 1006 4 br_53
port 191 nsew
rlabel metal1 s 35136 252 35164 1006 4 bl_54
port 192 nsew
rlabel metal1 s 35600 252 35628 1006 4 br_54
port 193 nsew
rlabel metal1 s 36224 252 36252 1006 4 bl_55
port 194 nsew
rlabel metal1 s 35760 252 35788 1006 4 br_55
port 195 nsew
rlabel metal1 s 36384 252 36412 1006 4 bl_56
port 196 nsew
rlabel metal1 s 36848 252 36876 1006 4 br_56
port 197 nsew
rlabel metal1 s 37472 252 37500 1006 4 bl_57
port 198 nsew
rlabel metal1 s 37008 252 37036 1006 4 br_57
port 199 nsew
rlabel metal1 s 37632 252 37660 1006 4 bl_58
port 200 nsew
rlabel metal1 s 38096 252 38124 1006 4 br_58
port 201 nsew
rlabel metal1 s 38720 252 38748 1006 4 bl_59
port 202 nsew
rlabel metal1 s 38256 252 38284 1006 4 br_59
port 203 nsew
rlabel metal1 s 38880 252 38908 1006 4 bl_60
port 204 nsew
rlabel metal1 s 39344 252 39372 1006 4 br_60
port 205 nsew
rlabel metal1 s 39968 252 39996 1006 4 bl_61
port 206 nsew
rlabel metal1 s 39504 252 39532 1006 4 br_61
port 207 nsew
rlabel metal1 s 40128 252 40156 1006 4 bl_62
port 208 nsew
rlabel metal1 s 40592 252 40620 1006 4 br_62
port 209 nsew
rlabel metal1 s 40752 252 40780 1006 4 br_63
port 210 nsew
rlabel metal1 s 41216 252 41244 1006 4 bl_63
port 211 nsew
rlabel metal1 s 41376 252 41404 1006 4 bl_64
port 212 nsew
rlabel metal1 s 41840 252 41868 1006 4 br_64
port 213 nsew
rlabel metal1 s 42464 252 42492 1006 4 bl_65
port 214 nsew
rlabel metal1 s 42000 252 42028 1006 4 br_65
port 215 nsew
rlabel metal1 s 42624 252 42652 1006 4 bl_66
port 216 nsew
rlabel metal1 s 43088 252 43116 1006 4 br_66
port 217 nsew
rlabel metal1 s 43712 252 43740 1006 4 bl_67
port 218 nsew
rlabel metal1 s 43248 252 43276 1006 4 br_67
port 219 nsew
rlabel metal1 s 43872 252 43900 1006 4 bl_68
port 220 nsew
rlabel metal1 s 44336 252 44364 1006 4 br_68
port 221 nsew
rlabel metal1 s 44960 252 44988 1006 4 bl_69
port 222 nsew
rlabel metal1 s 44496 252 44524 1006 4 br_69
port 223 nsew
rlabel metal1 s 45120 252 45148 1006 4 bl_70
port 224 nsew
rlabel metal1 s 45584 252 45612 1006 4 br_70
port 225 nsew
rlabel metal1 s 46208 252 46236 1006 4 bl_71
port 226 nsew
rlabel metal1 s 45744 252 45772 1006 4 br_71
port 227 nsew
rlabel metal1 s 46368 252 46396 1006 4 bl_72
port 228 nsew
rlabel metal1 s 46832 252 46860 1006 4 br_72
port 229 nsew
rlabel metal1 s 47456 252 47484 1006 4 bl_73
port 230 nsew
rlabel metal1 s 46992 252 47020 1006 4 br_73
port 231 nsew
rlabel metal1 s 47616 252 47644 1006 4 bl_74
port 232 nsew
rlabel metal1 s 48080 252 48108 1006 4 br_74
port 233 nsew
rlabel metal1 s 48704 252 48732 1006 4 bl_75
port 234 nsew
rlabel metal1 s 48240 252 48268 1006 4 br_75
port 235 nsew
rlabel metal1 s 48864 252 48892 1006 4 bl_76
port 236 nsew
rlabel metal1 s 49328 252 49356 1006 4 br_76
port 237 nsew
rlabel metal1 s 49952 252 49980 1006 4 bl_77
port 238 nsew
rlabel metal1 s 49488 252 49516 1006 4 br_77
port 239 nsew
rlabel metal1 s 50112 252 50140 1006 4 bl_78
port 240 nsew
rlabel metal1 s 50576 252 50604 1006 4 br_78
port 241 nsew
rlabel metal1 s 51200 252 51228 1006 4 bl_79
port 242 nsew
rlabel metal1 s 50736 252 50764 1006 4 br_79
port 243 nsew
rlabel metal1 s 51360 252 51388 1006 4 bl_80
port 244 nsew
rlabel metal1 s 51824 252 51852 1006 4 br_80
port 245 nsew
rlabel metal1 s 52448 252 52476 1006 4 bl_81
port 246 nsew
rlabel metal1 s 51984 252 52012 1006 4 br_81
port 247 nsew
rlabel metal1 s 52608 252 52636 1006 4 bl_82
port 248 nsew
rlabel metal1 s 53072 252 53100 1006 4 br_82
port 249 nsew
rlabel metal1 s 53696 252 53724 1006 4 bl_83
port 250 nsew
rlabel metal1 s 53232 252 53260 1006 4 br_83
port 251 nsew
rlabel metal1 s 53856 252 53884 1006 4 bl_84
port 252 nsew
rlabel metal1 s 54320 252 54348 1006 4 br_84
port 253 nsew
rlabel metal1 s 54944 252 54972 1006 4 bl_85
port 254 nsew
rlabel metal1 s 54480 252 54508 1006 4 br_85
port 255 nsew
rlabel metal1 s 55104 252 55132 1006 4 bl_86
port 256 nsew
rlabel metal1 s 55568 252 55596 1006 4 br_86
port 257 nsew
rlabel metal1 s 56192 252 56220 1006 4 bl_87
port 258 nsew
rlabel metal1 s 55728 252 55756 1006 4 br_87
port 259 nsew
rlabel metal1 s 56352 252 56380 1006 4 bl_88
port 260 nsew
rlabel metal1 s 56816 252 56844 1006 4 br_88
port 261 nsew
rlabel metal1 s 57440 252 57468 1006 4 bl_89
port 262 nsew
rlabel metal1 s 56976 252 57004 1006 4 br_89
port 263 nsew
rlabel metal1 s 57600 252 57628 1006 4 bl_90
port 264 nsew
rlabel metal1 s 58064 252 58092 1006 4 br_90
port 265 nsew
rlabel metal1 s 58688 252 58716 1006 4 bl_91
port 266 nsew
rlabel metal1 s 58224 252 58252 1006 4 br_91
port 267 nsew
rlabel metal1 s 58848 252 58876 1006 4 bl_92
port 268 nsew
rlabel metal1 s 59312 252 59340 1006 4 br_92
port 269 nsew
rlabel metal1 s 59936 252 59964 1006 4 bl_93
port 270 nsew
rlabel metal1 s 59472 252 59500 1006 4 br_93
port 271 nsew
rlabel metal1 s 60096 252 60124 1006 4 bl_94
port 272 nsew
rlabel metal1 s 60560 252 60588 1006 4 br_94
port 273 nsew
rlabel metal1 s 60720 252 60748 1006 4 br_95
port 274 nsew
rlabel metal1 s 61184 252 61212 1006 4 bl_95
port 275 nsew
rlabel metal1 s 61344 252 61372 1006 4 bl_96
port 276 nsew
rlabel metal1 s 61808 252 61836 1006 4 br_96
port 277 nsew
rlabel metal1 s 62432 252 62460 1006 4 bl_97
port 278 nsew
rlabel metal1 s 61968 252 61996 1006 4 br_97
port 279 nsew
rlabel metal1 s 62592 252 62620 1006 4 bl_98
port 280 nsew
rlabel metal1 s 63056 252 63084 1006 4 br_98
port 281 nsew
rlabel metal1 s 63680 252 63708 1006 4 bl_99
port 282 nsew
rlabel metal1 s 63216 252 63244 1006 4 br_99
port 283 nsew
rlabel metal1 s 63840 252 63868 1006 4 bl_100
port 284 nsew
rlabel metal1 s 64304 252 64332 1006 4 br_100
port 285 nsew
rlabel metal1 s 64928 252 64956 1006 4 bl_101
port 286 nsew
rlabel metal1 s 64464 252 64492 1006 4 br_101
port 287 nsew
rlabel metal1 s 65088 252 65116 1006 4 bl_102
port 288 nsew
rlabel metal1 s 65552 252 65580 1006 4 br_102
port 289 nsew
rlabel metal1 s 66176 252 66204 1006 4 bl_103
port 290 nsew
rlabel metal1 s 65712 252 65740 1006 4 br_103
port 291 nsew
rlabel metal1 s 66336 252 66364 1006 4 bl_104
port 292 nsew
rlabel metal1 s 66800 252 66828 1006 4 br_104
port 293 nsew
rlabel metal1 s 67424 252 67452 1006 4 bl_105
port 294 nsew
rlabel metal1 s 66960 252 66988 1006 4 br_105
port 295 nsew
rlabel metal1 s 67584 252 67612 1006 4 bl_106
port 296 nsew
rlabel metal1 s 68048 252 68076 1006 4 br_106
port 297 nsew
rlabel metal1 s 68672 252 68700 1006 4 bl_107
port 298 nsew
rlabel metal1 s 68208 252 68236 1006 4 br_107
port 299 nsew
rlabel metal1 s 68832 252 68860 1006 4 bl_108
port 300 nsew
rlabel metal1 s 69296 252 69324 1006 4 br_108
port 301 nsew
rlabel metal1 s 69920 252 69948 1006 4 bl_109
port 302 nsew
rlabel metal1 s 69456 252 69484 1006 4 br_109
port 303 nsew
rlabel metal1 s 70080 252 70108 1006 4 bl_110
port 304 nsew
rlabel metal1 s 70544 252 70572 1006 4 br_110
port 305 nsew
rlabel metal1 s 71168 252 71196 1006 4 bl_111
port 306 nsew
rlabel metal1 s 70704 252 70732 1006 4 br_111
port 307 nsew
rlabel metal1 s 71328 252 71356 1006 4 bl_112
port 308 nsew
rlabel metal1 s 71792 252 71820 1006 4 br_112
port 309 nsew
rlabel metal1 s 72416 252 72444 1006 4 bl_113
port 310 nsew
rlabel metal1 s 71952 252 71980 1006 4 br_113
port 311 nsew
rlabel metal1 s 72576 252 72604 1006 4 bl_114
port 312 nsew
rlabel metal1 s 73040 252 73068 1006 4 br_114
port 313 nsew
rlabel metal1 s 73664 252 73692 1006 4 bl_115
port 314 nsew
rlabel metal1 s 73200 252 73228 1006 4 br_115
port 315 nsew
rlabel metal1 s 73824 252 73852 1006 4 bl_116
port 316 nsew
rlabel metal1 s 74288 252 74316 1006 4 br_116
port 317 nsew
rlabel metal1 s 74912 252 74940 1006 4 bl_117
port 318 nsew
rlabel metal1 s 74448 252 74476 1006 4 br_117
port 319 nsew
rlabel metal1 s 75072 252 75100 1006 4 bl_118
port 320 nsew
rlabel metal1 s 75536 252 75564 1006 4 br_118
port 321 nsew
rlabel metal1 s 76160 252 76188 1006 4 bl_119
port 322 nsew
rlabel metal1 s 75696 252 75724 1006 4 br_119
port 323 nsew
rlabel metal1 s 76320 252 76348 1006 4 bl_120
port 324 nsew
rlabel metal1 s 76784 252 76812 1006 4 br_120
port 325 nsew
rlabel metal1 s 77408 252 77436 1006 4 bl_121
port 326 nsew
rlabel metal1 s 76944 252 76972 1006 4 br_121
port 327 nsew
rlabel metal1 s 77568 252 77596 1006 4 bl_122
port 328 nsew
rlabel metal1 s 78032 252 78060 1006 4 br_122
port 329 nsew
rlabel metal1 s 78656 252 78684 1006 4 bl_123
port 330 nsew
rlabel metal1 s 78192 252 78220 1006 4 br_123
port 331 nsew
rlabel metal1 s 78816 252 78844 1006 4 bl_124
port 332 nsew
rlabel metal1 s 79280 252 79308 1006 4 br_124
port 333 nsew
rlabel metal1 s 79904 252 79932 1006 4 bl_125
port 334 nsew
rlabel metal1 s 79440 252 79468 1006 4 br_125
port 335 nsew
rlabel metal1 s 80064 252 80092 1006 4 bl_126
port 336 nsew
rlabel metal1 s 80528 252 80556 1006 4 br_126
port 337 nsew
rlabel metal1 s 81152 252 81180 1006 4 bl_127
port 338 nsew
rlabel metal1 s 80688 252 80716 1006 4 br_127
port 339 nsew
rlabel locali s 1952 9051 1952 9051 4 wdriver_sel_0
port 68 nsew
rlabel locali s 21920 9051 21920 9051 4 wdriver_sel_1
port 69 nsew
rlabel locali s 41888 9051 41888 9051 4 wdriver_sel_2
port 14 nsew
rlabel locali s 61856 9051 61856 9051 4 wdriver_sel_3
port 15 nsew
<< properties >>
string FIXED_BBOX 0 0 81246 9585
string GDS_END 11864444
string GDS_FILE $PDKPATH/libs.ref/sky130_sram_macros/gds/sky130_sram_2kbyte_1rw1r_32x512_8.gds
string GDS_START 11595386
<< end >>
