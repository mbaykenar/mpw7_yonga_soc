magic
tech sky130B
magscale 1 2
timestamp 1649977179
<< nwell >>
rect -38 261 682 582
<< pwell >>
rect 1 163 187 203
rect 454 163 643 203
rect 1 67 643 163
rect 29 27 643 67
rect 29 -17 63 27
rect 454 21 643 27
<< locali >>
rect 117 425 440 491
rect 305 265 354 323
rect 572 299 627 493
rect 18 215 85 265
rect 305 199 470 265
rect 593 152 627 299
rect 572 83 627 152
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 644 561
rect 17 299 69 527
rect 119 265 153 377
rect 205 357 440 391
rect 474 367 530 527
rect 205 299 271 357
rect 406 333 440 357
rect 406 299 538 333
rect 504 265 538 299
rect 119 199 262 265
rect 504 199 559 265
rect 119 181 169 199
rect 17 17 69 181
rect 103 97 169 181
rect 504 165 538 199
rect 205 131 538 165
rect 205 51 257 131
rect 291 17 357 97
rect 391 61 425 131
rect 459 17 534 97
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 644 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
<< metal1 >>
rect 0 561 644 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 644 561
rect 0 496 644 527
rect 0 17 644 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 644 17
rect 0 -48 644 -17
<< labels >>
rlabel locali s 305 199 470 265 6 A
port 1 nsew signal input
rlabel locali s 305 265 354 323 6 A
port 1 nsew signal input
rlabel locali s 117 425 440 491 6 B
port 2 nsew signal input
rlabel locali s 18 215 85 265 6 C_N
port 3 nsew signal input
rlabel metal1 s 0 -48 644 48 8 VGND
port 4 nsew ground bidirectional abutment
rlabel pwell s 454 21 643 27 6 VNB
port 5 nsew ground bidirectional
rlabel pwell s 29 -17 63 27 6 VNB
port 5 nsew ground bidirectional
rlabel pwell s 29 27 643 67 6 VNB
port 5 nsew ground bidirectional
rlabel pwell s 1 67 643 163 6 VNB
port 5 nsew ground bidirectional
rlabel pwell s 454 163 643 203 6 VNB
port 5 nsew ground bidirectional
rlabel pwell s 1 163 187 203 6 VNB
port 5 nsew ground bidirectional
rlabel nwell s -38 261 682 582 6 VPB
port 6 nsew power bidirectional
rlabel metal1 s 0 496 644 592 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 572 83 627 152 6 X
port 8 nsew signal output
rlabel locali s 593 152 627 299 6 X
port 8 nsew signal output
rlabel locali s 572 299 627 493 6 X
port 8 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 644 544
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_END 1057358
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 1051152
<< end >>
