magic
tech sky130B
magscale 1 2
timestamp 1649977179
<< locali >>
rect 1784 3096 1818 3112
rect 1784 3046 1818 3062
rect 3135 2996 3588 3030
rect 1658 2950 1674 2984
rect 1708 2950 1724 2984
rect 1768 2860 1784 2894
rect 1818 2860 1834 2894
rect 1768 2636 1784 2670
rect 1818 2636 1834 2670
rect 1658 2546 1674 2580
rect 1708 2546 1724 2580
rect 3135 2500 3588 2534
rect 1784 2468 1818 2484
rect 1784 2418 1818 2434
rect 1784 2306 1818 2322
rect 1784 2256 1818 2272
rect 3135 2206 3588 2240
rect 1658 2160 1674 2194
rect 1708 2160 1724 2194
rect 1768 2070 1784 2104
rect 1818 2070 1834 2104
rect 1768 1846 1784 1880
rect 1818 1846 1834 1880
rect 1658 1756 1674 1790
rect 1708 1756 1724 1790
rect 3135 1710 3588 1744
rect 1784 1678 1818 1694
rect 1784 1628 1818 1644
rect 1784 1516 1818 1532
rect 1784 1466 1818 1482
rect 3135 1416 3588 1450
rect 1658 1370 1674 1404
rect 1708 1370 1724 1404
rect 1768 1280 1784 1314
rect 1818 1280 1834 1314
rect 1001 1100 1255 1134
rect 1289 1100 1305 1134
rect 460 1004 494 1020
rect 460 954 494 970
rect 1001 920 1035 1100
rect 1768 1056 1784 1090
rect 1818 1056 1834 1090
rect 1658 966 1674 1000
rect 1708 966 1724 1000
rect 3135 920 3588 954
rect 1784 888 1818 904
rect 1784 838 1818 854
rect 1001 705 1175 739
rect 1209 705 1225 739
rect 1784 726 1818 742
rect 1001 626 1035 705
rect 1784 676 1818 692
rect 3135 626 3588 660
rect 460 610 494 626
rect 1658 580 1674 614
rect 1708 580 1724 614
rect 460 560 494 576
rect 1768 490 1784 524
rect 1818 490 1834 524
rect 1001 310 1095 344
rect 1129 310 1145 344
rect 460 214 494 230
rect 460 164 494 180
rect 1001 130 1035 310
rect 1768 266 1784 300
rect 1818 266 1834 300
rect 1658 176 1674 210
rect 1708 176 1724 210
rect 3135 130 3588 164
rect 1784 98 1818 114
rect 1784 48 1818 64
<< viali >>
rect 1784 3062 1818 3096
rect 1674 2950 1708 2984
rect 1784 2860 1818 2894
rect 1784 2636 1818 2670
rect 1674 2546 1708 2580
rect 1784 2434 1818 2468
rect 1784 2272 1818 2306
rect 1674 2160 1708 2194
rect 1784 2070 1818 2104
rect 1784 1846 1818 1880
rect 1674 1756 1708 1790
rect 1784 1644 1818 1678
rect 1784 1482 1818 1516
rect 1674 1370 1708 1404
rect 1784 1280 1818 1314
rect 1255 1100 1289 1134
rect 460 970 494 1004
rect 1784 1056 1818 1090
rect 1674 966 1708 1000
rect 1784 854 1818 888
rect 1175 705 1209 739
rect 1784 692 1818 726
rect 460 576 494 610
rect 1674 580 1708 614
rect 1784 490 1818 524
rect 1095 310 1129 344
rect 460 180 494 214
rect 1784 266 1818 300
rect 1674 176 1708 210
rect 1784 64 1818 98
<< metal1 >>
rect 1326 3105 1378 3111
rect 62 3053 68 3105
rect 120 3053 126 3105
rect 80 229 108 3053
rect 160 2993 188 3080
rect 142 2941 148 2993
rect 200 2941 206 2993
rect 160 625 188 2941
rect 240 2903 268 3080
rect 222 2851 228 2903
rect 280 2851 286 2903
rect 240 1019 268 2851
rect 1098 2483 1126 3080
rect 1086 2477 1138 2483
rect 1086 2419 1138 2425
rect 1098 1693 1126 2419
rect 1178 2209 1206 3080
rect 1166 2203 1218 2209
rect 1166 2145 1218 2151
rect 1178 1805 1206 2145
rect 1166 1799 1218 1805
rect 1166 1741 1218 1747
rect 1086 1687 1138 1693
rect 1086 1629 1138 1635
rect 228 1013 280 1019
rect 222 961 228 1013
rect 280 961 286 1013
rect 445 961 451 1013
rect 503 961 509 1013
rect 228 955 280 961
rect 148 619 200 625
rect 142 567 148 619
rect 200 567 206 619
rect 148 561 200 567
rect 68 223 120 229
rect 62 171 68 223
rect 120 171 126 223
rect 68 165 120 171
rect 80 80 108 165
rect 160 80 188 561
rect 240 80 268 955
rect 445 567 451 619
rect 503 567 509 619
rect 584 421 612 1185
rect 856 421 884 1185
rect 1098 903 1126 1629
rect 1086 897 1138 903
rect 1086 839 1138 845
rect 566 369 572 421
rect 624 369 630 421
rect 838 369 844 421
rect 896 369 902 421
rect 445 171 451 223
rect 503 171 509 223
rect 584 80 612 369
rect 856 80 884 369
rect 1098 356 1126 839
rect 1178 751 1206 1741
rect 1258 1329 1286 3080
rect 1320 3053 1326 3105
rect 1378 3053 1384 3105
rect 1326 3047 1378 3053
rect 1338 2321 1366 3047
rect 1418 2999 1446 3080
rect 1406 2993 1458 2999
rect 1400 2941 1406 2993
rect 1458 2941 1464 2993
rect 1406 2935 1458 2941
rect 1418 2595 1446 2935
rect 1498 2909 1526 3080
rect 1769 3053 1775 3105
rect 1827 3053 1833 3105
rect 1659 2941 1665 2993
rect 1717 2941 1723 2993
rect 1486 2903 1538 2909
rect 1480 2851 1486 2903
rect 1538 2851 1544 2903
rect 1769 2851 1775 2903
rect 1827 2851 1833 2903
rect 1486 2845 1538 2851
rect 1498 2685 1526 2845
rect 1906 2814 1952 3204
rect 2330 2814 2378 3146
rect 2762 2814 2810 3146
rect 1897 2762 1903 2814
rect 1955 2762 1961 2814
rect 2322 2762 2328 2814
rect 2380 2762 2386 2814
rect 2754 2762 2760 2814
rect 2812 2762 2818 2814
rect 3154 2791 3182 3160
rect 3426 2791 3454 3160
rect 1486 2679 1538 2685
rect 1769 2627 1775 2679
rect 1827 2627 1833 2679
rect 1486 2621 1538 2627
rect 1406 2589 1458 2595
rect 1406 2531 1458 2537
rect 1326 2315 1378 2321
rect 1326 2257 1378 2263
rect 1338 1531 1366 2257
rect 1326 1525 1378 1531
rect 1326 1467 1378 1473
rect 1246 1323 1298 1329
rect 1246 1265 1298 1271
rect 1258 1146 1286 1265
rect 1249 1134 1295 1146
rect 1249 1105 1255 1134
rect 1246 1100 1255 1105
rect 1289 1105 1295 1134
rect 1289 1100 1298 1105
rect 1246 1099 1298 1100
rect 1246 1041 1298 1047
rect 1169 739 1215 751
rect 1169 705 1175 739
rect 1209 705 1215 739
rect 1169 693 1215 705
rect 1178 629 1206 693
rect 1166 623 1218 629
rect 1166 565 1218 571
rect 1089 344 1135 356
rect 1089 310 1095 344
rect 1129 310 1135 344
rect 1089 298 1135 310
rect 1098 113 1126 298
rect 1178 225 1206 565
rect 1258 539 1286 1041
rect 1338 741 1366 1467
rect 1418 1419 1446 2531
rect 1498 2119 1526 2621
rect 1659 2537 1665 2589
rect 1717 2537 1723 2589
rect 1769 2425 1775 2477
rect 1827 2425 1833 2477
rect 1769 2263 1775 2315
rect 1827 2263 1833 2315
rect 1659 2151 1665 2203
rect 1717 2151 1723 2203
rect 1486 2113 1538 2119
rect 1769 2061 1775 2113
rect 1827 2061 1833 2113
rect 1486 2055 1538 2061
rect 1498 1895 1526 2055
rect 1906 2024 1952 2762
rect 2330 2024 2378 2762
rect 2762 2024 2810 2762
rect 3136 2739 3142 2791
rect 3194 2739 3200 2791
rect 3408 2739 3414 2791
rect 3466 2739 3472 2791
rect 1897 1972 1903 2024
rect 1955 1972 1961 2024
rect 2322 1972 2328 2024
rect 2380 1972 2386 2024
rect 2754 1972 2760 2024
rect 2812 1972 2818 2024
rect 3154 2001 3182 2739
rect 3426 2001 3454 2739
rect 1486 1889 1538 1895
rect 1769 1837 1775 1889
rect 1827 1837 1833 1889
rect 1486 1831 1538 1837
rect 1406 1413 1458 1419
rect 1406 1355 1458 1361
rect 1418 1015 1446 1355
rect 1406 1009 1458 1015
rect 1406 951 1458 957
rect 1326 735 1378 741
rect 1326 677 1378 683
rect 1246 533 1298 539
rect 1246 475 1298 481
rect 1258 315 1286 475
rect 1246 309 1298 315
rect 1246 251 1298 257
rect 1166 219 1218 225
rect 1166 161 1218 167
rect 1086 107 1138 113
rect 1178 80 1206 161
rect 1258 80 1286 251
rect 1338 80 1366 677
rect 1418 80 1446 951
rect 1498 80 1526 1831
rect 1659 1747 1665 1799
rect 1717 1747 1723 1799
rect 1769 1635 1775 1687
rect 1827 1635 1833 1687
rect 1769 1473 1775 1525
rect 1827 1473 1833 1525
rect 1659 1361 1665 1413
rect 1717 1361 1723 1413
rect 1769 1271 1775 1323
rect 1827 1271 1833 1323
rect 1906 1234 1952 1972
rect 2330 1234 2378 1972
rect 2762 1234 2810 1972
rect 3136 1949 3142 2001
rect 3194 1949 3200 2001
rect 3408 1949 3414 2001
rect 3466 1949 3472 2001
rect 1897 1182 1903 1234
rect 1955 1182 1961 1234
rect 2322 1182 2328 1234
rect 2380 1182 2386 1234
rect 2754 1182 2760 1234
rect 2812 1182 2818 1234
rect 3154 1211 3182 1949
rect 3426 1211 3454 1949
rect 1769 1047 1775 1099
rect 1827 1047 1833 1099
rect 1659 957 1665 1009
rect 1717 957 1723 1009
rect 1769 845 1775 897
rect 1827 845 1833 897
rect 1769 683 1775 735
rect 1827 683 1833 735
rect 1659 571 1665 623
rect 1717 571 1723 623
rect 1769 481 1775 533
rect 1827 481 1833 533
rect 1906 444 1952 1182
rect 2330 444 2378 1182
rect 2762 444 2810 1182
rect 3136 1159 3142 1211
rect 3194 1159 3200 1211
rect 3408 1159 3414 1211
rect 3466 1159 3472 1211
rect 1897 392 1903 444
rect 1955 392 1961 444
rect 2322 392 2328 444
rect 2380 392 2386 444
rect 2754 392 2760 444
rect 2812 392 2818 444
rect 3154 421 3182 1159
rect 3426 421 3454 1159
rect 1769 257 1775 309
rect 1827 257 1833 309
rect 1659 167 1665 219
rect 1717 167 1723 219
rect 1769 55 1775 107
rect 1827 55 1833 107
rect 1906 80 1952 392
rect 2330 80 2378 392
rect 2762 80 2810 392
rect 3136 369 3142 421
rect 3194 369 3200 421
rect 3408 369 3414 421
rect 3466 369 3472 421
rect 3154 80 3182 369
rect 3426 80 3454 369
rect 1086 49 1138 55
<< via1 >>
rect 68 3053 120 3105
rect 148 2941 200 2993
rect 228 2851 280 2903
rect 1086 2425 1138 2477
rect 1166 2151 1218 2203
rect 1166 1747 1218 1799
rect 1086 1635 1138 1687
rect 228 961 280 1013
rect 451 1004 503 1013
rect 451 970 460 1004
rect 460 970 494 1004
rect 494 970 503 1004
rect 451 961 503 970
rect 148 567 200 619
rect 68 171 120 223
rect 451 610 503 619
rect 451 576 460 610
rect 460 576 494 610
rect 494 576 503 610
rect 451 567 503 576
rect 1086 845 1138 897
rect 572 369 624 421
rect 844 369 896 421
rect 451 214 503 223
rect 451 180 460 214
rect 460 180 494 214
rect 494 180 503 214
rect 451 171 503 180
rect 1326 3053 1378 3105
rect 1406 2941 1458 2993
rect 1775 3096 1827 3105
rect 1775 3062 1784 3096
rect 1784 3062 1818 3096
rect 1818 3062 1827 3096
rect 1775 3053 1827 3062
rect 1665 2984 1717 2993
rect 1665 2950 1674 2984
rect 1674 2950 1708 2984
rect 1708 2950 1717 2984
rect 1665 2941 1717 2950
rect 1486 2851 1538 2903
rect 1775 2894 1827 2903
rect 1775 2860 1784 2894
rect 1784 2860 1818 2894
rect 1818 2860 1827 2894
rect 1775 2851 1827 2860
rect 1903 2762 1955 2814
rect 2328 2762 2380 2814
rect 2760 2762 2812 2814
rect 1486 2627 1538 2679
rect 1775 2670 1827 2679
rect 1775 2636 1784 2670
rect 1784 2636 1818 2670
rect 1818 2636 1827 2670
rect 1775 2627 1827 2636
rect 1406 2537 1458 2589
rect 1326 2263 1378 2315
rect 1326 1473 1378 1525
rect 1246 1271 1298 1323
rect 1246 1047 1298 1099
rect 1166 571 1218 623
rect 1665 2580 1717 2589
rect 1665 2546 1674 2580
rect 1674 2546 1708 2580
rect 1708 2546 1717 2580
rect 1665 2537 1717 2546
rect 1775 2468 1827 2477
rect 1775 2434 1784 2468
rect 1784 2434 1818 2468
rect 1818 2434 1827 2468
rect 1775 2425 1827 2434
rect 1775 2306 1827 2315
rect 1775 2272 1784 2306
rect 1784 2272 1818 2306
rect 1818 2272 1827 2306
rect 1775 2263 1827 2272
rect 1665 2194 1717 2203
rect 1665 2160 1674 2194
rect 1674 2160 1708 2194
rect 1708 2160 1717 2194
rect 1665 2151 1717 2160
rect 1486 2061 1538 2113
rect 1775 2104 1827 2113
rect 1775 2070 1784 2104
rect 1784 2070 1818 2104
rect 1818 2070 1827 2104
rect 1775 2061 1827 2070
rect 3142 2739 3194 2791
rect 3414 2739 3466 2791
rect 1903 1972 1955 2024
rect 2328 1972 2380 2024
rect 2760 1972 2812 2024
rect 1486 1837 1538 1889
rect 1775 1880 1827 1889
rect 1775 1846 1784 1880
rect 1784 1846 1818 1880
rect 1818 1846 1827 1880
rect 1775 1837 1827 1846
rect 1406 1361 1458 1413
rect 1406 957 1458 1009
rect 1326 683 1378 735
rect 1246 481 1298 533
rect 1246 257 1298 309
rect 1166 167 1218 219
rect 1086 55 1138 107
rect 1665 1790 1717 1799
rect 1665 1756 1674 1790
rect 1674 1756 1708 1790
rect 1708 1756 1717 1790
rect 1665 1747 1717 1756
rect 1775 1678 1827 1687
rect 1775 1644 1784 1678
rect 1784 1644 1818 1678
rect 1818 1644 1827 1678
rect 1775 1635 1827 1644
rect 1775 1516 1827 1525
rect 1775 1482 1784 1516
rect 1784 1482 1818 1516
rect 1818 1482 1827 1516
rect 1775 1473 1827 1482
rect 1665 1404 1717 1413
rect 1665 1370 1674 1404
rect 1674 1370 1708 1404
rect 1708 1370 1717 1404
rect 1665 1361 1717 1370
rect 1775 1314 1827 1323
rect 1775 1280 1784 1314
rect 1784 1280 1818 1314
rect 1818 1280 1827 1314
rect 1775 1271 1827 1280
rect 3142 1949 3194 2001
rect 3414 1949 3466 2001
rect 1903 1182 1955 1234
rect 2328 1182 2380 1234
rect 2760 1182 2812 1234
rect 1775 1090 1827 1099
rect 1775 1056 1784 1090
rect 1784 1056 1818 1090
rect 1818 1056 1827 1090
rect 1775 1047 1827 1056
rect 1665 1000 1717 1009
rect 1665 966 1674 1000
rect 1674 966 1708 1000
rect 1708 966 1717 1000
rect 1665 957 1717 966
rect 1775 888 1827 897
rect 1775 854 1784 888
rect 1784 854 1818 888
rect 1818 854 1827 888
rect 1775 845 1827 854
rect 1775 726 1827 735
rect 1775 692 1784 726
rect 1784 692 1818 726
rect 1818 692 1827 726
rect 1775 683 1827 692
rect 1665 614 1717 623
rect 1665 580 1674 614
rect 1674 580 1708 614
rect 1708 580 1717 614
rect 1665 571 1717 580
rect 1775 524 1827 533
rect 1775 490 1784 524
rect 1784 490 1818 524
rect 1818 490 1827 524
rect 1775 481 1827 490
rect 3142 1159 3194 1211
rect 3414 1159 3466 1211
rect 1903 392 1955 444
rect 2328 392 2380 444
rect 2760 392 2812 444
rect 1775 300 1827 309
rect 1775 266 1784 300
rect 1784 266 1818 300
rect 1818 266 1827 300
rect 1775 257 1827 266
rect 1665 210 1717 219
rect 1665 176 1674 210
rect 1674 176 1708 210
rect 1708 176 1717 210
rect 1665 167 1717 176
rect 1775 98 1827 107
rect 1775 64 1784 98
rect 1784 64 1818 98
rect 1818 64 1827 98
rect 1775 55 1827 64
rect 3142 369 3194 421
rect 3414 369 3466 421
<< metal2 >>
rect 68 3105 120 3111
rect 1326 3105 1378 3111
rect 1775 3105 1827 3111
rect 1320 3093 1326 3105
rect 120 3065 1326 3093
rect 1320 3053 1326 3065
rect 1378 3093 1384 3105
rect 1378 3065 1775 3093
rect 1378 3053 1384 3065
rect 68 3047 120 3053
rect 1326 3047 1378 3053
rect 1775 3047 1827 3053
rect 148 2993 200 2999
rect 1406 2993 1458 2999
rect 1400 2981 1406 2993
rect 200 2953 1406 2981
rect 1400 2941 1406 2953
rect 1458 2981 1464 2993
rect 1659 2981 1665 2993
rect 1458 2953 1665 2981
rect 1458 2941 1464 2953
rect 1659 2941 1665 2953
rect 1717 2941 1723 2993
rect 148 2935 200 2941
rect 1406 2935 1458 2941
rect 228 2903 280 2909
rect 1486 2903 1538 2909
rect 1480 2891 1486 2903
rect 280 2863 1486 2891
rect 1480 2851 1486 2863
rect 1538 2891 1544 2903
rect 1769 2891 1775 2903
rect 1538 2863 1775 2891
rect 1538 2851 1544 2863
rect 1769 2851 1775 2863
rect 1827 2851 1833 2903
rect 228 2845 280 2851
rect 1486 2845 1538 2851
rect 1901 2816 1957 2825
rect 1901 2751 1957 2760
rect 2326 2816 2382 2825
rect 2326 2751 2382 2760
rect 2758 2816 2814 2825
rect 2758 2751 2814 2760
rect 3140 2793 3196 2802
rect 3140 2728 3196 2737
rect 3412 2793 3468 2802
rect 3412 2728 3468 2737
rect 1480 2627 1486 2679
rect 1538 2667 1544 2679
rect 1769 2667 1775 2679
rect 1538 2639 1775 2667
rect 1538 2627 1544 2639
rect 1769 2627 1775 2639
rect 1827 2627 1833 2679
rect 1400 2537 1406 2589
rect 1458 2577 1464 2589
rect 1659 2577 1665 2589
rect 1458 2549 1665 2577
rect 1458 2537 1464 2549
rect 1659 2537 1665 2549
rect 1717 2537 1723 2589
rect 1775 2477 1827 2483
rect 1080 2425 1086 2477
rect 1138 2465 1144 2477
rect 1138 2437 1775 2465
rect 1138 2425 1144 2437
rect 1775 2419 1827 2425
rect 1775 2315 1827 2321
rect 1320 2263 1326 2315
rect 1378 2303 1384 2315
rect 1378 2275 1775 2303
rect 1378 2263 1384 2275
rect 1775 2257 1827 2263
rect 1160 2151 1166 2203
rect 1218 2191 1224 2203
rect 1659 2191 1665 2203
rect 1218 2163 1665 2191
rect 1218 2151 1224 2163
rect 1659 2151 1665 2163
rect 1717 2151 1723 2203
rect 1480 2061 1486 2113
rect 1538 2101 1544 2113
rect 1769 2101 1775 2113
rect 1538 2073 1775 2101
rect 1538 2061 1544 2073
rect 1769 2061 1775 2073
rect 1827 2061 1833 2113
rect 1901 2026 1957 2035
rect 1901 1961 1957 1970
rect 2326 2026 2382 2035
rect 2326 1961 2382 1970
rect 2758 2026 2814 2035
rect 2758 1961 2814 1970
rect 3140 2003 3196 2012
rect 3140 1938 3196 1947
rect 3412 2003 3468 2012
rect 3412 1938 3468 1947
rect 1480 1837 1486 1889
rect 1538 1877 1544 1889
rect 1769 1877 1775 1889
rect 1538 1849 1775 1877
rect 1538 1837 1544 1849
rect 1769 1837 1775 1849
rect 1827 1837 1833 1889
rect 1160 1747 1166 1799
rect 1218 1787 1224 1799
rect 1659 1787 1665 1799
rect 1218 1759 1665 1787
rect 1218 1747 1224 1759
rect 1659 1747 1665 1759
rect 1717 1747 1723 1799
rect 1775 1687 1827 1693
rect 1080 1635 1086 1687
rect 1138 1675 1144 1687
rect 1138 1647 1775 1675
rect 1138 1635 1144 1647
rect 1775 1629 1827 1635
rect 1775 1525 1827 1531
rect 1320 1473 1326 1525
rect 1378 1513 1384 1525
rect 1378 1485 1775 1513
rect 1378 1473 1384 1485
rect 1775 1467 1827 1473
rect 1400 1361 1406 1413
rect 1458 1401 1464 1413
rect 1659 1401 1665 1413
rect 1458 1373 1665 1401
rect 1458 1361 1464 1373
rect 1659 1361 1665 1373
rect 1717 1361 1723 1413
rect 1240 1271 1246 1323
rect 1298 1311 1304 1323
rect 1769 1311 1775 1323
rect 1298 1283 1775 1311
rect 1298 1271 1304 1283
rect 1769 1271 1775 1283
rect 1827 1271 1833 1323
rect 1901 1236 1957 1245
rect 1901 1171 1957 1180
rect 2326 1236 2382 1245
rect 2326 1171 2382 1180
rect 2758 1236 2814 1245
rect 2758 1171 2814 1180
rect 3140 1213 3196 1222
rect 3140 1148 3196 1157
rect 3412 1213 3468 1222
rect 3412 1148 3468 1157
rect 1240 1047 1246 1099
rect 1298 1087 1304 1099
rect 1769 1087 1775 1099
rect 1298 1059 1775 1087
rect 1298 1047 1304 1059
rect 1769 1047 1775 1059
rect 1827 1047 1833 1099
rect 228 1013 280 1019
rect 451 1013 503 1019
rect 280 973 451 1001
rect 228 955 280 961
rect 451 955 503 961
rect 1400 957 1406 1009
rect 1458 997 1464 1009
rect 1659 997 1665 1009
rect 1458 969 1665 997
rect 1458 957 1464 969
rect 1659 957 1665 969
rect 1717 957 1723 1009
rect 1775 897 1827 903
rect 1080 845 1086 897
rect 1138 885 1144 897
rect 1138 857 1775 885
rect 1138 845 1144 857
rect 1775 839 1827 845
rect 1775 735 1827 741
rect 1320 683 1326 735
rect 1378 723 1384 735
rect 1378 695 1775 723
rect 1378 683 1384 695
rect 1775 677 1827 683
rect 148 619 200 625
rect 451 619 503 625
rect 200 579 451 607
rect 148 561 200 567
rect 1160 571 1166 623
rect 1218 611 1224 623
rect 1659 611 1665 623
rect 1218 583 1665 611
rect 1218 571 1224 583
rect 1659 571 1665 583
rect 1717 571 1723 623
rect 451 561 503 567
rect 1240 481 1246 533
rect 1298 521 1304 533
rect 1769 521 1775 533
rect 1298 493 1775 521
rect 1298 481 1304 493
rect 1769 481 1775 493
rect 1827 481 1833 533
rect 1901 446 1957 455
rect 570 423 626 432
rect 570 358 626 367
rect 842 423 898 432
rect 1901 381 1957 390
rect 2326 446 2382 455
rect 2326 381 2382 390
rect 2758 446 2814 455
rect 2758 381 2814 390
rect 3140 423 3196 432
rect 842 358 898 367
rect 3140 358 3196 367
rect 3412 423 3468 432
rect 3412 358 3468 367
rect 1240 257 1246 309
rect 1298 297 1304 309
rect 1769 297 1775 309
rect 1298 269 1775 297
rect 1298 257 1304 269
rect 1769 257 1775 269
rect 1827 257 1833 309
rect 68 223 120 229
rect 451 223 503 229
rect 120 183 451 211
rect 68 165 120 171
rect 451 165 503 171
rect 1160 167 1166 219
rect 1218 207 1224 219
rect 1659 207 1665 219
rect 1218 179 1665 207
rect 1218 167 1224 179
rect 1659 167 1665 179
rect 1717 167 1723 219
rect 1775 107 1827 113
rect 1080 55 1086 107
rect 1138 95 1144 107
rect 1138 67 1775 95
rect 1138 55 1144 67
rect 1775 49 1827 55
<< via2 >>
rect 1901 2814 1957 2816
rect 1901 2762 1903 2814
rect 1903 2762 1955 2814
rect 1955 2762 1957 2814
rect 1901 2760 1957 2762
rect 2326 2814 2382 2816
rect 2326 2762 2328 2814
rect 2328 2762 2380 2814
rect 2380 2762 2382 2814
rect 2326 2760 2382 2762
rect 2758 2814 2814 2816
rect 2758 2762 2760 2814
rect 2760 2762 2812 2814
rect 2812 2762 2814 2814
rect 2758 2760 2814 2762
rect 3140 2791 3196 2793
rect 3140 2739 3142 2791
rect 3142 2739 3194 2791
rect 3194 2739 3196 2791
rect 3140 2737 3196 2739
rect 3412 2791 3468 2793
rect 3412 2739 3414 2791
rect 3414 2739 3466 2791
rect 3466 2739 3468 2791
rect 3412 2737 3468 2739
rect 1901 2024 1957 2026
rect 1901 1972 1903 2024
rect 1903 1972 1955 2024
rect 1955 1972 1957 2024
rect 1901 1970 1957 1972
rect 2326 2024 2382 2026
rect 2326 1972 2328 2024
rect 2328 1972 2380 2024
rect 2380 1972 2382 2024
rect 2326 1970 2382 1972
rect 2758 2024 2814 2026
rect 2758 1972 2760 2024
rect 2760 1972 2812 2024
rect 2812 1972 2814 2024
rect 2758 1970 2814 1972
rect 3140 2001 3196 2003
rect 3140 1949 3142 2001
rect 3142 1949 3194 2001
rect 3194 1949 3196 2001
rect 3140 1947 3196 1949
rect 3412 2001 3468 2003
rect 3412 1949 3414 2001
rect 3414 1949 3466 2001
rect 3466 1949 3468 2001
rect 3412 1947 3468 1949
rect 1901 1234 1957 1236
rect 1901 1182 1903 1234
rect 1903 1182 1955 1234
rect 1955 1182 1957 1234
rect 1901 1180 1957 1182
rect 2326 1234 2382 1236
rect 2326 1182 2328 1234
rect 2328 1182 2380 1234
rect 2380 1182 2382 1234
rect 2326 1180 2382 1182
rect 2758 1234 2814 1236
rect 2758 1182 2760 1234
rect 2760 1182 2812 1234
rect 2812 1182 2814 1234
rect 2758 1180 2814 1182
rect 3140 1211 3196 1213
rect 3140 1159 3142 1211
rect 3142 1159 3194 1211
rect 3194 1159 3196 1211
rect 3140 1157 3196 1159
rect 3412 1211 3468 1213
rect 3412 1159 3414 1211
rect 3414 1159 3466 1211
rect 3466 1159 3468 1211
rect 3412 1157 3468 1159
rect 1901 444 1957 446
rect 570 421 626 423
rect 570 369 572 421
rect 572 369 624 421
rect 624 369 626 421
rect 570 367 626 369
rect 842 421 898 423
rect 842 369 844 421
rect 844 369 896 421
rect 896 369 898 421
rect 1901 392 1903 444
rect 1903 392 1955 444
rect 1955 392 1957 444
rect 1901 390 1957 392
rect 2326 444 2382 446
rect 2326 392 2328 444
rect 2328 392 2380 444
rect 2380 392 2382 444
rect 2326 390 2382 392
rect 2758 444 2814 446
rect 2758 392 2760 444
rect 2760 392 2812 444
rect 2812 392 2814 444
rect 2758 390 2814 392
rect 3140 421 3196 423
rect 842 367 898 369
rect 3140 369 3142 421
rect 3142 369 3194 421
rect 3194 369 3196 421
rect 3140 367 3196 369
rect 3412 421 3468 423
rect 3412 369 3414 421
rect 3414 369 3466 421
rect 3466 369 3468 421
rect 3412 367 3468 369
<< metal3 >>
rect 1880 2816 1978 2837
rect 1880 2760 1901 2816
rect 1957 2760 1978 2816
rect 1880 2739 1978 2760
rect 2305 2816 2403 2837
rect 2305 2760 2326 2816
rect 2382 2760 2403 2816
rect 2305 2739 2403 2760
rect 2737 2816 2835 2837
rect 2737 2760 2758 2816
rect 2814 2760 2835 2816
rect 2737 2739 2835 2760
rect 3119 2793 3217 2814
rect 3119 2737 3140 2793
rect 3196 2737 3217 2793
rect 3119 2716 3217 2737
rect 3391 2793 3489 2814
rect 3391 2737 3412 2793
rect 3468 2737 3489 2793
rect 3391 2716 3489 2737
rect 1880 2026 1978 2047
rect 1880 1970 1901 2026
rect 1957 1970 1978 2026
rect 1880 1949 1978 1970
rect 2305 2026 2403 2047
rect 2305 1970 2326 2026
rect 2382 1970 2403 2026
rect 2305 1949 2403 1970
rect 2737 2026 2835 2047
rect 2737 1970 2758 2026
rect 2814 1970 2835 2026
rect 2737 1949 2835 1970
rect 3119 2003 3217 2024
rect 3119 1947 3140 2003
rect 3196 1947 3217 2003
rect 3119 1926 3217 1947
rect 3391 2003 3489 2024
rect 3391 1947 3412 2003
rect 3468 1947 3489 2003
rect 3391 1926 3489 1947
rect 1880 1236 1978 1257
rect 1880 1180 1901 1236
rect 1957 1180 1978 1236
rect 1880 1159 1978 1180
rect 2305 1236 2403 1257
rect 2305 1180 2326 1236
rect 2382 1180 2403 1236
rect 2305 1159 2403 1180
rect 2737 1236 2835 1257
rect 2737 1180 2758 1236
rect 2814 1180 2835 1236
rect 2737 1159 2835 1180
rect 3119 1213 3217 1234
rect 3119 1157 3140 1213
rect 3196 1157 3217 1213
rect 3119 1136 3217 1157
rect 3391 1213 3489 1234
rect 3391 1157 3412 1213
rect 3468 1157 3489 1213
rect 3391 1136 3489 1157
rect 1880 446 1978 467
rect 549 423 647 444
rect 549 367 570 423
rect 626 367 647 423
rect 549 346 647 367
rect 821 423 919 444
rect 821 367 842 423
rect 898 367 919 423
rect 1880 390 1901 446
rect 1957 390 1978 446
rect 1880 369 1978 390
rect 2305 446 2403 467
rect 2305 390 2326 446
rect 2382 390 2403 446
rect 2305 369 2403 390
rect 2737 446 2835 467
rect 2737 390 2758 446
rect 2814 390 2835 446
rect 2737 369 2835 390
rect 3119 423 3217 444
rect 821 346 919 367
rect 3119 367 3140 423
rect 3196 367 3217 423
rect 3119 346 3217 367
rect 3391 423 3489 444
rect 3391 367 3412 423
rect 3468 367 3489 423
rect 3391 346 3489 367
use and3_dec  and3_dec_0
timestamp 1649977179
transform 1 0 1658 0 -1 3160
box 0 -60 1948 490
use and3_dec  and3_dec_1
timestamp 1649977179
transform 1 0 1658 0 1 2370
box 0 -60 1948 490
use and3_dec  and3_dec_2
timestamp 1649977179
transform 1 0 1658 0 -1 2370
box 0 -60 1948 490
use and3_dec  and3_dec_3
timestamp 1649977179
transform 1 0 1658 0 1 1580
box 0 -60 1948 490
use and3_dec  and3_dec_4
timestamp 1649977179
transform 1 0 1658 0 -1 1580
box 0 -60 1948 490
use and3_dec  and3_dec_5
timestamp 1649977179
transform 1 0 1658 0 1 790
box 0 -60 1948 490
use and3_dec  and3_dec_6
timestamp 1649977179
transform 1 0 1658 0 -1 790
box 0 -60 1948 490
use and3_dec  and3_dec_7
timestamp 1649977179
transform 1 0 1658 0 1 0
box 0 -60 1948 490
use contact_7  contact_7_0
timestamp 1649977179
transform 1 0 1772 0 1 48
box 0 0 1 1
use contact_7  contact_7_1
timestamp 1649977179
transform 1 0 448 0 1 164
box 0 0 1 1
use contact_7  contact_7_2
timestamp 1649977179
transform 1 0 448 0 1 954
box 0 0 1 1
use contact_7  contact_7_3
timestamp 1649977179
transform 1 0 448 0 1 560
box 0 0 1 1
use contact_7  contact_7_4
timestamp 1649977179
transform 1 0 1772 0 1 1466
box 0 0 1 1
use contact_7  contact_7_5
timestamp 1649977179
transform 1 0 1772 0 1 838
box 0 0 1 1
use contact_7  contact_7_6
timestamp 1649977179
transform 1 0 1772 0 1 676
box 0 0 1 1
use contact_7  contact_7_7
timestamp 1649977179
transform 1 0 1772 0 1 3046
box 0 0 1 1
use contact_7  contact_7_8
timestamp 1649977179
transform 1 0 1772 0 1 2418
box 0 0 1 1
use contact_7  contact_7_9
timestamp 1649977179
transform 1 0 1772 0 1 2256
box 0 0 1 1
use contact_7  contact_7_10
timestamp 1649977179
transform 1 0 1772 0 1 1628
box 0 0 1 1
use contact_8  contact_8_0
timestamp 1649977179
transform 1 0 2754 0 1 1176
box 0 0 1 1
use contact_8  contact_8_1
timestamp 1649977179
transform 1 0 2754 0 1 1176
box 0 0 1 1
use contact_8  contact_8_2
timestamp 1649977179
transform 1 0 3408 0 1 1153
box 0 0 1 1
use contact_8  contact_8_3
timestamp 1649977179
transform 1 0 3408 0 1 1153
box 0 0 1 1
use contact_8  contact_8_4
timestamp 1649977179
transform 1 0 2322 0 1 386
box 0 0 1 1
use contact_8  contact_8_5
timestamp 1649977179
transform 1 0 2322 0 1 386
box 0 0 1 1
use contact_8  contact_8_6
timestamp 1649977179
transform 1 0 2754 0 1 386
box 0 0 1 1
use contact_8  contact_8_7
timestamp 1649977179
transform 1 0 2754 0 1 386
box 0 0 1 1
use contact_8  contact_8_8
timestamp 1649977179
transform 1 0 1897 0 1 1176
box 0 0 1 1
use contact_8  contact_8_9
timestamp 1649977179
transform 1 0 1897 0 1 1176
box 0 0 1 1
use contact_8  contact_8_10
timestamp 1649977179
transform 1 0 3136 0 1 1153
box 0 0 1 1
use contact_8  contact_8_11
timestamp 1649977179
transform 1 0 3136 0 1 1153
box 0 0 1 1
use contact_8  contact_8_12
timestamp 1649977179
transform 1 0 1897 0 1 386
box 0 0 1 1
use contact_8  contact_8_13
timestamp 1649977179
transform 1 0 1897 0 1 386
box 0 0 1 1
use contact_8  contact_8_14
timestamp 1649977179
transform 1 0 3136 0 1 363
box 0 0 1 1
use contact_8  contact_8_15
timestamp 1649977179
transform 1 0 3136 0 1 363
box 0 0 1 1
use contact_8  contact_8_16
timestamp 1649977179
transform 1 0 3408 0 1 363
box 0 0 1 1
use contact_8  contact_8_17
timestamp 1649977179
transform 1 0 3408 0 1 363
box 0 0 1 1
use contact_8  contact_8_18
timestamp 1649977179
transform 1 0 2322 0 1 1176
box 0 0 1 1
use contact_8  contact_8_19
timestamp 1649977179
transform 1 0 2322 0 1 1176
box 0 0 1 1
use contact_8  contact_8_20
timestamp 1649977179
transform 1 0 1769 0 1 49
box 0 0 1 1
use contact_8  contact_8_21
timestamp 1649977179
transform 1 0 445 0 1 165
box 0 0 1 1
use contact_8  contact_8_22
timestamp 1649977179
transform 1 0 566 0 1 363
box 0 0 1 1
use contact_8  contact_8_23
timestamp 1649977179
transform 1 0 566 0 1 363
box 0 0 1 1
use contact_8  contact_8_24
timestamp 1649977179
transform 1 0 222 0 1 955
box 0 0 1 1
use contact_8  contact_8_25
timestamp 1649977179
transform 1 0 445 0 1 955
box 0 0 1 1
use contact_8  contact_8_26
timestamp 1649977179
transform 1 0 142 0 1 561
box 0 0 1 1
use contact_8  contact_8_27
timestamp 1649977179
transform 1 0 445 0 1 561
box 0 0 1 1
use contact_8  contact_8_28
timestamp 1649977179
transform 1 0 62 0 1 165
box 0 0 1 1
use contact_8  contact_8_29
timestamp 1649977179
transform 1 0 1769 0 1 1467
box 0 0 1 1
use contact_8  contact_8_30
timestamp 1649977179
transform 1 0 838 0 1 363
box 0 0 1 1
use contact_8  contact_8_31
timestamp 1649977179
transform 1 0 838 0 1 363
box 0 0 1 1
use contact_8  contact_8_32
timestamp 1649977179
transform 1 0 1769 0 1 839
box 0 0 1 1
use contact_8  contact_8_33
timestamp 1649977179
transform 1 0 1769 0 1 677
box 0 0 1 1
use contact_8  contact_8_34
timestamp 1649977179
transform 1 0 1769 0 1 3047
box 0 0 1 1
use contact_8  contact_8_35
timestamp 1649977179
transform 1 0 1769 0 1 2419
box 0 0 1 1
use contact_8  contact_8_36
timestamp 1649977179
transform 1 0 1769 0 1 2257
box 0 0 1 1
use contact_8  contact_8_37
timestamp 1649977179
transform 1 0 1769 0 1 1629
box 0 0 1 1
use contact_8  contact_8_38
timestamp 1649977179
transform 1 0 1480 0 1 2845
box 0 0 1 1
use contact_8  contact_8_39
timestamp 1649977179
transform 1 0 222 0 1 2845
box 0 0 1 1
use contact_8  contact_8_40
timestamp 1649977179
transform 1 0 1400 0 1 2935
box 0 0 1 1
use contact_8  contact_8_41
timestamp 1649977179
transform 1 0 142 0 1 2935
box 0 0 1 1
use contact_8  contact_8_42
timestamp 1649977179
transform 1 0 1320 0 1 3047
box 0 0 1 1
use contact_8  contact_8_43
timestamp 1649977179
transform 1 0 62 0 1 3047
box 0 0 1 1
use contact_8  contact_8_44
timestamp 1649977179
transform 1 0 1897 0 1 2756
box 0 0 1 1
use contact_8  contact_8_45
timestamp 1649977179
transform 1 0 1897 0 1 2756
box 0 0 1 1
use contact_8  contact_8_46
timestamp 1649977179
transform 1 0 3136 0 1 2733
box 0 0 1 1
use contact_8  contact_8_47
timestamp 1649977179
transform 1 0 3136 0 1 2733
box 0 0 1 1
use contact_8  contact_8_48
timestamp 1649977179
transform 1 0 1897 0 1 1966
box 0 0 1 1
use contact_8  contact_8_49
timestamp 1649977179
transform 1 0 1897 0 1 1966
box 0 0 1 1
use contact_8  contact_8_50
timestamp 1649977179
transform 1 0 3136 0 1 1943
box 0 0 1 1
use contact_8  contact_8_51
timestamp 1649977179
transform 1 0 3136 0 1 1943
box 0 0 1 1
use contact_8  contact_8_52
timestamp 1649977179
transform 1 0 2322 0 1 2756
box 0 0 1 1
use contact_8  contact_8_53
timestamp 1649977179
transform 1 0 2322 0 1 2756
box 0 0 1 1
use contact_8  contact_8_54
timestamp 1649977179
transform 1 0 2754 0 1 2756
box 0 0 1 1
use contact_8  contact_8_55
timestamp 1649977179
transform 1 0 2754 0 1 2756
box 0 0 1 1
use contact_8  contact_8_56
timestamp 1649977179
transform 1 0 3408 0 1 2733
box 0 0 1 1
use contact_8  contact_8_57
timestamp 1649977179
transform 1 0 3408 0 1 2733
box 0 0 1 1
use contact_8  contact_8_58
timestamp 1649977179
transform 1 0 2322 0 1 1966
box 0 0 1 1
use contact_8  contact_8_59
timestamp 1649977179
transform 1 0 2322 0 1 1966
box 0 0 1 1
use contact_8  contact_8_60
timestamp 1649977179
transform 1 0 2754 0 1 1966
box 0 0 1 1
use contact_8  contact_8_61
timestamp 1649977179
transform 1 0 2754 0 1 1966
box 0 0 1 1
use contact_8  contact_8_62
timestamp 1649977179
transform 1 0 3408 0 1 1943
box 0 0 1 1
use contact_8  contact_8_63
timestamp 1649977179
transform 1 0 3408 0 1 1943
box 0 0 1 1
use contact_9  contact_9_0
timestamp 1649977179
transform 1 0 2753 0 1 1171
box 0 0 1 1
use contact_9  contact_9_1
timestamp 1649977179
transform 1 0 2753 0 1 1171
box 0 0 1 1
use contact_9  contact_9_2
timestamp 1649977179
transform 1 0 3407 0 1 1148
box 0 0 1 1
use contact_9  contact_9_3
timestamp 1649977179
transform 1 0 3407 0 1 1148
box 0 0 1 1
use contact_9  contact_9_4
timestamp 1649977179
transform 1 0 2321 0 1 381
box 0 0 1 1
use contact_9  contact_9_5
timestamp 1649977179
transform 1 0 2321 0 1 381
box 0 0 1 1
use contact_9  contact_9_6
timestamp 1649977179
transform 1 0 2753 0 1 381
box 0 0 1 1
use contact_9  contact_9_7
timestamp 1649977179
transform 1 0 2753 0 1 381
box 0 0 1 1
use contact_9  contact_9_8
timestamp 1649977179
transform 1 0 1896 0 1 1171
box 0 0 1 1
use contact_9  contact_9_9
timestamp 1649977179
transform 1 0 1896 0 1 1171
box 0 0 1 1
use contact_9  contact_9_10
timestamp 1649977179
transform 1 0 3135 0 1 1148
box 0 0 1 1
use contact_9  contact_9_11
timestamp 1649977179
transform 1 0 3135 0 1 1148
box 0 0 1 1
use contact_9  contact_9_12
timestamp 1649977179
transform 1 0 1896 0 1 381
box 0 0 1 1
use contact_9  contact_9_13
timestamp 1649977179
transform 1 0 1896 0 1 381
box 0 0 1 1
use contact_9  contact_9_14
timestamp 1649977179
transform 1 0 3135 0 1 358
box 0 0 1 1
use contact_9  contact_9_15
timestamp 1649977179
transform 1 0 3135 0 1 358
box 0 0 1 1
use contact_9  contact_9_16
timestamp 1649977179
transform 1 0 3407 0 1 358
box 0 0 1 1
use contact_9  contact_9_17
timestamp 1649977179
transform 1 0 3407 0 1 358
box 0 0 1 1
use contact_9  contact_9_18
timestamp 1649977179
transform 1 0 2321 0 1 1171
box 0 0 1 1
use contact_9  contact_9_19
timestamp 1649977179
transform 1 0 2321 0 1 1171
box 0 0 1 1
use contact_9  contact_9_20
timestamp 1649977179
transform 1 0 565 0 1 358
box 0 0 1 1
use contact_9  contact_9_21
timestamp 1649977179
transform 1 0 565 0 1 358
box 0 0 1 1
use contact_9  contact_9_22
timestamp 1649977179
transform 1 0 837 0 1 358
box 0 0 1 1
use contact_9  contact_9_23
timestamp 1649977179
transform 1 0 837 0 1 358
box 0 0 1 1
use contact_9  contact_9_24
timestamp 1649977179
transform 1 0 1896 0 1 2751
box 0 0 1 1
use contact_9  contact_9_25
timestamp 1649977179
transform 1 0 1896 0 1 2751
box 0 0 1 1
use contact_9  contact_9_26
timestamp 1649977179
transform 1 0 3135 0 1 2728
box 0 0 1 1
use contact_9  contact_9_27
timestamp 1649977179
transform 1 0 3135 0 1 2728
box 0 0 1 1
use contact_9  contact_9_28
timestamp 1649977179
transform 1 0 1896 0 1 1961
box 0 0 1 1
use contact_9  contact_9_29
timestamp 1649977179
transform 1 0 1896 0 1 1961
box 0 0 1 1
use contact_9  contact_9_30
timestamp 1649977179
transform 1 0 3135 0 1 1938
box 0 0 1 1
use contact_9  contact_9_31
timestamp 1649977179
transform 1 0 3135 0 1 1938
box 0 0 1 1
use contact_9  contact_9_32
timestamp 1649977179
transform 1 0 2321 0 1 2751
box 0 0 1 1
use contact_9  contact_9_33
timestamp 1649977179
transform 1 0 2321 0 1 2751
box 0 0 1 1
use contact_9  contact_9_34
timestamp 1649977179
transform 1 0 2753 0 1 2751
box 0 0 1 1
use contact_9  contact_9_35
timestamp 1649977179
transform 1 0 2753 0 1 2751
box 0 0 1 1
use contact_9  contact_9_36
timestamp 1649977179
transform 1 0 3407 0 1 2728
box 0 0 1 1
use contact_9  contact_9_37
timestamp 1649977179
transform 1 0 3407 0 1 2728
box 0 0 1 1
use contact_9  contact_9_38
timestamp 1649977179
transform 1 0 2321 0 1 1961
box 0 0 1 1
use contact_9  contact_9_39
timestamp 1649977179
transform 1 0 2321 0 1 1961
box 0 0 1 1
use contact_9  contact_9_40
timestamp 1649977179
transform 1 0 2753 0 1 1961
box 0 0 1 1
use contact_9  contact_9_41
timestamp 1649977179
transform 1 0 2753 0 1 1961
box 0 0 1 1
use contact_9  contact_9_42
timestamp 1649977179
transform 1 0 3407 0 1 1938
box 0 0 1 1
use contact_9  contact_9_43
timestamp 1649977179
transform 1 0 3407 0 1 1938
box 0 0 1 1
use contact_26  contact_26_0
timestamp 1649977179
transform 1 0 1079 0 1 298
box 0 0 1 1
use contact_26  contact_26_1
timestamp 1649977179
transform 1 0 1239 0 1 1088
box 0 0 1 1
use contact_26  contact_26_2
timestamp 1649977179
transform 1 0 1159 0 1 693
box 0 0 1 1
use contact_27  contact_27_0
timestamp 1649977179
transform 1 0 1320 0 1 677
box 0 0 1 1
use contact_27  contact_27_1
timestamp 1649977179
transform 1 0 1240 0 1 251
box 0 0 1 1
use contact_27  contact_27_2
timestamp 1649977179
transform 1 0 1160 0 1 161
box 0 0 1 1
use contact_27  contact_27_3
timestamp 1649977179
transform 1 0 1080 0 1 49
box 0 0 1 1
use contact_27  contact_27_4
timestamp 1649977179
transform 1 0 1240 0 1 1265
box 0 0 1 1
use contact_27  contact_27_5
timestamp 1649977179
transform 1 0 1400 0 1 1355
box 0 0 1 1
use contact_27  contact_27_6
timestamp 1649977179
transform 1 0 1320 0 1 1467
box 0 0 1 1
use contact_27  contact_27_7
timestamp 1649977179
transform 1 0 1240 0 1 1041
box 0 0 1 1
use contact_27  contact_27_8
timestamp 1649977179
transform 1 0 1400 0 1 951
box 0 0 1 1
use contact_27  contact_27_9
timestamp 1649977179
transform 1 0 1080 0 1 839
box 0 0 1 1
use contact_27  contact_27_10
timestamp 1649977179
transform 1 0 1240 0 1 475
box 0 0 1 1
use contact_27  contact_27_11
timestamp 1649977179
transform 1 0 1160 0 1 565
box 0 0 1 1
use contact_27  contact_27_12
timestamp 1649977179
transform 1 0 1480 0 1 2845
box 0 0 1 1
use contact_27  contact_27_13
timestamp 1649977179
transform 1 0 1400 0 1 2935
box 0 0 1 1
use contact_27  contact_27_14
timestamp 1649977179
transform 1 0 1320 0 1 3047
box 0 0 1 1
use contact_27  contact_27_15
timestamp 1649977179
transform 1 0 1480 0 1 2621
box 0 0 1 1
use contact_27  contact_27_16
timestamp 1649977179
transform 1 0 1400 0 1 2531
box 0 0 1 1
use contact_27  contact_27_17
timestamp 1649977179
transform 1 0 1080 0 1 2419
box 0 0 1 1
use contact_27  contact_27_18
timestamp 1649977179
transform 1 0 1480 0 1 2055
box 0 0 1 1
use contact_27  contact_27_19
timestamp 1649977179
transform 1 0 1160 0 1 2145
box 0 0 1 1
use contact_27  contact_27_20
timestamp 1649977179
transform 1 0 1320 0 1 2257
box 0 0 1 1
use contact_27  contact_27_21
timestamp 1649977179
transform 1 0 1480 0 1 1831
box 0 0 1 1
use contact_27  contact_27_22
timestamp 1649977179
transform 1 0 1160 0 1 1741
box 0 0 1 1
use contact_27  contact_27_23
timestamp 1649977179
transform 1 0 1080 0 1 1629
box 0 0 1 1
use contact_28  contact_28_0
timestamp 1649977179
transform 1 0 1768 0 1 260
box 0 0 1 1
use contact_28  contact_28_1
timestamp 1649977179
transform 1 0 1658 0 1 170
box 0 0 1 1
use contact_28  contact_28_2
timestamp 1649977179
transform 1 0 1768 0 1 1274
box 0 0 1 1
use contact_28  contact_28_3
timestamp 1649977179
transform 1 0 1658 0 1 1364
box 0 0 1 1
use contact_28  contact_28_4
timestamp 1649977179
transform 1 0 1768 0 1 1050
box 0 0 1 1
use contact_28  contact_28_5
timestamp 1649977179
transform 1 0 1658 0 1 960
box 0 0 1 1
use contact_28  contact_28_6
timestamp 1649977179
transform 1 0 1768 0 1 484
box 0 0 1 1
use contact_28  contact_28_7
timestamp 1649977179
transform 1 0 1658 0 1 574
box 0 0 1 1
use contact_28  contact_28_8
timestamp 1649977179
transform 1 0 1658 0 1 2944
box 0 0 1 1
use contact_28  contact_28_9
timestamp 1649977179
transform 1 0 1768 0 1 2630
box 0 0 1 1
use contact_28  contact_28_10
timestamp 1649977179
transform 1 0 1658 0 1 2540
box 0 0 1 1
use contact_28  contact_28_11
timestamp 1649977179
transform 1 0 1768 0 1 2064
box 0 0 1 1
use contact_28  contact_28_12
timestamp 1649977179
transform 1 0 1658 0 1 2154
box 0 0 1 1
use contact_28  contact_28_13
timestamp 1649977179
transform 1 0 1768 0 1 1840
box 0 0 1 1
use contact_28  contact_28_14
timestamp 1649977179
transform 1 0 1658 0 1 1750
box 0 0 1 1
use contact_28  contact_28_15
timestamp 1649977179
transform 1 0 1768 0 1 2854
box 0 0 1 1
use contact_29  contact_29_0
timestamp 1649977179
transform 1 0 1769 0 1 257
box 0 0 1 1
use contact_29  contact_29_1
timestamp 1649977179
transform 1 0 1659 0 1 167
box 0 0 1 1
use contact_29  contact_29_2
timestamp 1649977179
transform 1 0 1769 0 1 1271
box 0 0 1 1
use contact_29  contact_29_3
timestamp 1649977179
transform 1 0 1659 0 1 1361
box 0 0 1 1
use contact_29  contact_29_4
timestamp 1649977179
transform 1 0 1769 0 1 1047
box 0 0 1 1
use contact_29  contact_29_5
timestamp 1649977179
transform 1 0 1659 0 1 957
box 0 0 1 1
use contact_29  contact_29_6
timestamp 1649977179
transform 1 0 1769 0 1 481
box 0 0 1 1
use contact_29  contact_29_7
timestamp 1649977179
transform 1 0 1659 0 1 571
box 0 0 1 1
use contact_29  contact_29_8
timestamp 1649977179
transform 1 0 1659 0 1 2941
box 0 0 1 1
use contact_29  contact_29_9
timestamp 1649977179
transform 1 0 1769 0 1 2627
box 0 0 1 1
use contact_29  contact_29_10
timestamp 1649977179
transform 1 0 1659 0 1 2537
box 0 0 1 1
use contact_29  contact_29_11
timestamp 1649977179
transform 1 0 1769 0 1 2061
box 0 0 1 1
use contact_29  contact_29_12
timestamp 1649977179
transform 1 0 1659 0 1 2151
box 0 0 1 1
use contact_29  contact_29_13
timestamp 1649977179
transform 1 0 1769 0 1 1837
box 0 0 1 1
use contact_29  contact_29_14
timestamp 1649977179
transform 1 0 1659 0 1 1747
box 0 0 1 1
use contact_29  contact_29_15
timestamp 1649977179
transform 1 0 1769 0 1 2851
box 0 0 1 1
use pinv_dec  pinv_dec_0
timestamp 1649977179
transform 1 0 400 0 -1 790
box 44 0 636 490
use pinv_dec  pinv_dec_1
timestamp 1649977179
transform 1 0 400 0 1 0
box 44 0 636 490
use pinv_dec  pinv_dec_2
timestamp 1649977179
transform 1 0 400 0 1 790
box 44 0 636 490
<< labels >>
rlabel locali s 3361 2223 3361 2223 4 out_5
port 9 nsew
rlabel locali s 3361 1433 3361 1433 4 out_3
port 7 nsew
rlabel locali s 3361 937 3361 937 4 out_2
port 6 nsew
rlabel locali s 3361 2517 3361 2517 4 out_6
port 10 nsew
rlabel locali s 3361 1727 3361 1727 4 out_4
port 8 nsew
rlabel locali s 3361 3013 3361 3013 4 out_7
port 11 nsew
rlabel locali s 3361 147 3361 147 4 out_0
port 4 nsew
rlabel locali s 3361 643 3361 643 4 out_1
port 5 nsew
rlabel metal1 s 254 987 254 987 4 in_2
port 3 nsew
rlabel metal1 s 94 197 94 197 4 in_0
port 1 nsew
rlabel metal1 s 174 593 174 593 4 in_1
port 2 nsew
rlabel metal3 s 3440 2765 3440 2765 4 vdd
port 12 nsew
rlabel metal3 s 2786 2788 2786 2788 4 vdd
port 12 nsew
rlabel metal3 s 2786 418 2786 418 4 vdd
port 12 nsew
rlabel metal3 s 3440 1975 3440 1975 4 vdd
port 12 nsew
rlabel metal3 s 870 395 870 395 4 vdd
port 12 nsew
rlabel metal3 s 2354 418 2354 418 4 vdd
port 12 nsew
rlabel metal3 s 3440 1185 3440 1185 4 vdd
port 12 nsew
rlabel metal3 s 2786 1208 2786 1208 4 vdd
port 12 nsew
rlabel metal3 s 3440 395 3440 395 4 vdd
port 12 nsew
rlabel metal3 s 2786 1998 2786 1998 4 vdd
port 12 nsew
rlabel metal3 s 2354 1998 2354 1998 4 vdd
port 12 nsew
rlabel metal3 s 2354 1208 2354 1208 4 vdd
port 12 nsew
rlabel metal3 s 2354 2788 2354 2788 4 vdd
port 12 nsew
rlabel metal3 s 1929 418 1929 418 4 gnd
port 13 nsew
rlabel metal3 s 3168 1975 3168 1975 4 gnd
port 13 nsew
rlabel metal3 s 1929 1208 1929 1208 4 gnd
port 13 nsew
rlabel metal3 s 3168 1185 3168 1185 4 gnd
port 13 nsew
rlabel metal3 s 598 395 598 395 4 gnd
port 13 nsew
rlabel metal3 s 1929 1998 1929 1998 4 gnd
port 13 nsew
rlabel metal3 s 3168 395 3168 395 4 gnd
port 13 nsew
rlabel metal3 s 3168 2765 3168 2765 4 gnd
port 13 nsew
rlabel metal3 s 1929 2788 1929 2788 4 gnd
port 13 nsew
<< properties >>
string FIXED_BBOX 0 0 3588 3160
string GDS_END 131580
string GDS_FILE $PDKPATH/libs.ref/sky130_sram_macros/gds/sram_1rw1r_32_256_8_sky130.gds
string GDS_START 112716
<< end >>
