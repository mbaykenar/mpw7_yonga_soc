magic
tech sky130B
magscale 12 1
timestamp 1598786981
<< metal5 >>
rect 0 90 45 105
rect 0 15 15 90
rect 30 15 45 90
rect 0 0 45 15
<< properties >>
string FIXED_BBOX 0 -30 60 105
<< end >>
