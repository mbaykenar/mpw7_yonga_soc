magic
tech sky130A
magscale 1 2
timestamp 1649977179
use sky130_fd_pr__hvdfm1sd2__example_55959141808243  sky130_fd_pr__hvdfm1sd2__example_55959141808243_0
timestamp 1649977179
transform 1 0 180 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfm1sd2__example_55959141808243  sky130_fd_pr__hvdfm1sd2__example_55959141808243_1
timestamp 1649977179
transform 1 0 416 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfm1sd2__example_55959141808243  sky130_fd_pr__hvdfm1sd2__example_55959141808243_2
timestamp 1649977179
transform 1 0 652 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfm1sd__example_55959141808242  sky130_fd_pr__hvdfm1sd__example_55959141808242_0
timestamp 1649977179
transform -1 0 0 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfm1sd__example_55959141808242  sky130_fd_pr__hvdfm1sd__example_55959141808242_1
timestamp 1649977179
transform 1 0 888 0 1 0
box 0 0 1 1
<< labels >>
flabel comment s 916 85 916 85 0 FreeSans 300 0 0 0 S
flabel comment s 680 85 680 85 0 FreeSans 300 0 0 0 D
flabel comment s 444 85 444 85 0 FreeSans 300 0 0 0 S
flabel comment s 208 85 208 85 0 FreeSans 300 0 0 0 D
flabel comment s -28 85 -28 85 0 FreeSans 300 0 0 0 S
<< properties >>
string GDS_END 37240046
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 37237502
<< end >>
