magic
tech sky130A
timestamp 1649977179
<< properties >>
string GDS_END 39433700
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 39433440
<< end >>
