magic
tech sky130A
magscale 1 2
timestamp 1649977179
<< nwell >>
rect 0 415 534 1116
<< pwell >>
rect 40 118 497 310
<< mvnmos >>
rect 119 144 239 284
rect 295 144 415 284
<< mvpmos >>
rect 119 750 239 950
rect 295 750 415 950
rect 119 482 239 682
rect 295 482 415 682
<< mvndiff >>
rect 66 272 119 284
rect 66 238 74 272
rect 108 238 119 272
rect 66 204 119 238
rect 66 170 74 204
rect 108 170 119 204
rect 66 144 119 170
rect 239 272 295 284
rect 239 238 250 272
rect 284 238 295 272
rect 239 204 295 238
rect 239 170 250 204
rect 284 170 295 204
rect 239 144 295 170
rect 415 272 471 284
rect 415 238 426 272
rect 460 238 471 272
rect 415 204 471 238
rect 415 170 426 204
rect 460 170 471 204
rect 415 144 471 170
<< mvpdiff >>
rect 66 932 119 950
rect 66 898 74 932
rect 108 898 119 932
rect 66 864 119 898
rect 66 830 74 864
rect 108 830 119 864
rect 66 796 119 830
rect 66 762 74 796
rect 108 762 119 796
rect 66 750 119 762
rect 239 932 295 950
rect 239 898 250 932
rect 284 898 295 932
rect 239 864 295 898
rect 239 830 250 864
rect 284 830 295 864
rect 239 796 295 830
rect 239 762 250 796
rect 284 762 295 796
rect 239 750 295 762
rect 415 932 468 950
rect 415 898 426 932
rect 460 898 468 932
rect 415 864 468 898
rect 415 830 426 864
rect 460 830 468 864
rect 415 796 468 830
rect 415 762 426 796
rect 460 762 468 796
rect 415 750 468 762
rect 66 670 119 682
rect 66 636 74 670
rect 108 636 119 670
rect 66 602 119 636
rect 66 568 74 602
rect 108 568 119 602
rect 66 534 119 568
rect 66 500 74 534
rect 108 500 119 534
rect 66 482 119 500
rect 239 670 295 682
rect 239 636 250 670
rect 284 636 295 670
rect 239 602 295 636
rect 239 568 250 602
rect 284 568 295 602
rect 239 482 295 568
rect 415 670 468 682
rect 415 636 426 670
rect 460 636 468 670
rect 415 602 468 636
rect 415 568 426 602
rect 460 568 468 602
rect 415 534 468 568
rect 415 500 426 534
rect 460 500 468 534
rect 415 482 468 500
<< mvndiffc >>
rect 74 238 108 272
rect 74 170 108 204
rect 250 238 284 272
rect 250 170 284 204
rect 426 238 460 272
rect 426 170 460 204
<< mvpdiffc >>
rect 74 898 108 932
rect 74 830 108 864
rect 74 762 108 796
rect 250 898 284 932
rect 250 830 284 864
rect 250 762 284 796
rect 426 898 460 932
rect 426 830 460 864
rect 426 762 460 796
rect 74 636 108 670
rect 74 568 108 602
rect 74 500 108 534
rect 250 636 284 670
rect 250 568 284 602
rect 426 636 460 670
rect 426 568 460 602
rect 426 500 460 534
<< poly >>
rect 119 950 239 976
rect 295 950 415 976
rect 119 682 239 750
rect 295 682 415 750
rect 119 434 239 482
rect 119 400 162 434
rect 196 400 239 434
rect 119 366 239 400
rect 119 332 162 366
rect 196 332 239 366
rect 119 284 239 332
rect 295 434 415 482
rect 295 400 340 434
rect 374 400 415 434
rect 295 366 415 400
rect 295 332 340 366
rect 374 332 415 366
rect 295 284 415 332
rect 119 118 239 144
rect 295 118 415 144
<< polycont >>
rect 162 400 196 434
rect 162 332 196 366
rect 340 400 374 434
rect 340 332 374 366
<< locali >>
rect 74 932 108 944
rect 74 864 108 872
rect 74 796 108 830
rect 74 670 108 762
rect 74 602 108 636
rect 74 534 108 568
rect 250 932 284 948
rect 250 864 284 898
rect 250 796 284 830
rect 250 670 284 762
rect 250 602 284 636
rect 250 552 284 568
rect 426 932 460 978
rect 426 864 460 898
rect 426 796 460 830
rect 426 670 460 762
rect 426 602 460 636
rect 426 534 460 568
rect 74 484 108 500
rect 250 500 426 518
rect 250 484 460 500
rect 146 400 162 434
rect 196 400 212 434
rect 146 366 212 400
rect 146 332 162 366
rect 196 332 212 366
rect 74 272 108 288
rect 74 227 108 238
rect 74 155 108 170
rect 250 272 284 484
rect 324 400 340 434
rect 374 400 390 434
rect 324 366 390 400
rect 324 332 340 366
rect 374 332 390 366
rect 250 204 284 238
rect 250 154 284 170
rect 426 272 460 288
rect 426 227 460 238
rect 426 155 460 170
<< viali >>
rect 74 944 108 978
rect 74 898 108 906
rect 74 872 108 898
rect 74 204 108 227
rect 74 193 108 204
rect 74 121 108 155
rect 426 204 460 227
rect 426 193 460 204
rect 426 121 460 155
<< metal1 >>
rect 62 978 472 1062
rect 62 944 74 978
rect 108 944 472 978
rect 62 906 472 944
rect 62 872 74 906
rect 108 872 472 906
rect 62 859 472 872
rect 41 227 472 239
rect 41 193 74 227
rect 108 193 426 227
rect 460 193 472 227
rect 41 155 472 193
rect 41 121 74 155
rect 108 121 426 155
rect 460 121 472 155
rect 41 24 472 121
use sky130_fd_pr__hvdfl1sd__example_55959141808418  sky130_fd_pr__hvdfl1sd__example_55959141808418_0
timestamp 1649977179
transform -1 0 295 0 -1 682
box 0 0 1 1
use sky130_fd_pr__model__nfet_highvoltage__example_55959141808419  sky130_fd_pr__model__nfet_highvoltage__example_55959141808419_0
timestamp 1649977179
transform 1 0 119 0 -1 284
box -28 0 324 63
use sky130_fd_pr__model__pfet_highvoltage__example_55959141808420  sky130_fd_pr__model__pfet_highvoltage__example_55959141808420_0
timestamp 1649977179
transform -1 0 415 0 -1 682
box -28 0 145 100
use sky130_fd_pr__model__pfet_highvoltage__example_55959141808420  sky130_fd_pr__model__pfet_highvoltage__example_55959141808420_1
timestamp 1649977179
transform 1 0 119 0 -1 682
box -28 0 145 100
use sky130_fd_pr__model__pfet_highvoltage__example_55959141808421  sky130_fd_pr__model__pfet_highvoltage__example_55959141808421_0
timestamp 1649977179
transform 1 0 119 0 1 750
box -28 0 324 97
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_0
timestamp 1649977179
transform 0 -1 460 -1 0 227
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_1
timestamp 1649977179
transform 0 -1 108 1 0 872
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_2
timestamp 1649977179
transform 0 -1 108 -1 0 227
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_559591418083  sky130_fd_pr__via_pol1__example_559591418083_0
timestamp 1649977179
transform 0 -1 390 1 0 316
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_559591418083  sky130_fd_pr__via_pol1__example_559591418083_1
timestamp 1649977179
transform 0 -1 212 1 0 316
box 0 0 1 1
<< labels >>
flabel locali s 149 355 200 396 0 FreeSans 400 0 0 0 IN0
port 1 nsew
<< properties >>
string GDS_END 35743774
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 35741646
<< end >>
