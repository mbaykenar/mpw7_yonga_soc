magic
tech sky130B
magscale 1 2
timestamp 1649977179
<< nwell >>
rect -36 679 1700 1471
<< pwell >>
rect 1528 25 1630 159
<< psubdiff >>
rect 1554 109 1604 133
rect 1554 75 1562 109
rect 1596 75 1604 109
rect 1554 51 1604 75
<< nsubdiff >>
rect 1554 1339 1604 1363
rect 1554 1305 1562 1339
rect 1596 1305 1604 1339
rect 1554 1281 1604 1305
<< psubdiffcont >>
rect 1562 75 1596 109
<< nsubdiffcont >>
rect 1562 1305 1596 1339
<< poly >>
rect 114 740 144 907
rect 48 724 144 740
rect 48 690 64 724
rect 98 690 144 724
rect 48 674 144 690
rect 114 507 144 674
<< polycont >>
rect 64 690 98 724
<< locali >>
rect 0 1397 1664 1431
rect 62 1130 96 1397
rect 274 1130 308 1397
rect 490 1130 524 1397
rect 706 1130 740 1397
rect 922 1130 956 1397
rect 1138 1130 1172 1397
rect 1354 1130 1388 1397
rect 1562 1339 1596 1397
rect 1562 1289 1596 1305
rect 64 724 98 740
rect 64 674 98 690
rect 812 724 846 1096
rect 812 690 863 724
rect 812 318 846 690
rect 62 17 96 218
rect 274 17 308 218
rect 490 17 524 218
rect 706 17 740 218
rect 922 17 956 218
rect 1138 17 1172 218
rect 1354 17 1388 218
rect 1562 109 1596 125
rect 1562 17 1596 75
rect 0 -17 1664 17
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_16  sky130_sram_1kbyte_1rw1r_32x256_8_contact_16_0
timestamp 1649977179
transform 1 0 48 0 1 674
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_28  sky130_sram_1kbyte_1rw1r_32x256_8_contact_28_0
timestamp 1649977179
transform 1 0 1554 0 1 1281
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_29  sky130_sram_1kbyte_1rw1r_32x256_8_contact_29_0
timestamp 1649977179
transform 1 0 1554 0 1 51
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_nmos_m13_w2_000_sli_dli_da_p  sky130_sram_1kbyte_1rw1r_32x256_8_nmos_m13_w2_000_sli_dli_da_p_0
timestamp 1649977179
transform 1 0 54 0 1 51
box -26 -26 1472 456
use sky130_sram_1kbyte_1rw1r_32x256_8_pmos_m13_w2_000_sli_dli_da_p  sky130_sram_1kbyte_1rw1r_32x256_8_pmos_m13_w2_000_sli_dli_da_p_0
timestamp 1649977179
transform 1 0 54 0 1 963
box -59 -56 1505 454
<< labels >>
rlabel locali s 81 707 81 707 4 A
port 1 nsew
rlabel locali s 846 707 846 707 4 Z
port 2 nsew
rlabel locali s 832 0 832 0 4 gnd
port 3 nsew
rlabel locali s 832 1414 832 1414 4 vdd
port 4 nsew
<< properties >>
string FIXED_BBOX 0 0 1664 1414
string GDS_END 382704
string GDS_FILE $PDKPATH/libs.ref/sky130_sram_macros/gds/sky130_sram_1kbyte_1rw1r_32x256_8.gds
string GDS_START 380066
<< end >>
