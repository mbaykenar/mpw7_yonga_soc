magic
tech sky130B
magscale 1 2
timestamp 1662552610
<< viali >>
rect 2053 27557 2087 27591
rect 3985 27557 4019 27591
rect 5181 27557 5215 27591
rect 5825 27557 5859 27591
rect 7757 27557 7791 27591
rect 8401 27557 8435 27591
rect 10333 27557 10367 27591
rect 10977 27557 11011 27591
rect 14105 27557 14139 27591
rect 14933 27557 14967 27591
rect 15577 27557 15611 27591
rect 18061 27557 18095 27591
rect 18705 27557 18739 27591
rect 19993 27557 20027 27591
rect 20637 27557 20671 27591
rect 21281 27557 21315 27591
rect 23213 27557 23247 27591
rect 24593 27557 24627 27591
rect 25237 27557 25271 27591
rect 25881 27557 25915 27591
rect 26985 27557 27019 27591
rect 30389 27557 30423 27591
rect 31033 27557 31067 27591
rect 32321 27557 32355 27591
rect 33609 27557 33643 27591
rect 34713 27557 34747 27591
rect 37289 27557 37323 27591
rect 37933 27557 37967 27591
rect 38577 27557 38611 27591
rect 40049 27557 40083 27591
rect 41337 27557 41371 27591
rect 43913 27557 43947 27591
rect 45201 27557 45235 27591
rect 45845 27557 45879 27591
rect 46489 27557 46523 27591
rect 1409 27489 1443 27523
rect 7113 27489 7147 27523
rect 9689 27489 9723 27523
rect 11713 27489 11747 27523
rect 12357 27489 12391 27523
rect 13001 27489 13035 27523
rect 16681 27489 16715 27523
rect 22569 27489 22603 27523
rect 23857 27489 23891 27523
rect 27813 27489 27847 27523
rect 28457 27489 28491 27523
rect 29561 27489 29595 27523
rect 35357 27489 35391 27523
rect 36001 27489 36035 27523
rect 40693 27489 40727 27523
rect 42625 27489 42659 27523
rect 2697 27421 2731 27455
rect 42901 27421 42935 27455
rect 47869 27421 47903 27455
rect 48053 27285 48087 27319
rect 2697 27081 2731 27115
rect 47593 27081 47627 27115
rect 2053 27013 2087 27047
rect 1409 26945 1443 26979
rect 6561 26945 6595 26979
rect 9137 26945 9171 26979
rect 19441 26945 19475 26979
rect 22017 26945 22051 26979
rect 36185 26945 36219 26979
rect 38761 26945 38795 26979
rect 42441 26945 42475 26979
rect 43913 26945 43947 26979
rect 45753 26945 45787 26979
rect 47041 26945 47075 26979
rect 46397 26877 46431 26911
rect 2053 26537 2087 26571
rect 47501 26537 47535 26571
rect 46857 26401 46891 26435
rect 1409 26333 1443 26367
rect 48145 26197 48179 26231
rect 1409 25857 1443 25891
rect 48145 25857 48179 25891
rect 47041 25789 47075 25823
rect 1409 25245 1443 25279
rect 48145 25245 48179 25279
rect 1409 24565 1443 24599
rect 48145 24565 48179 24599
rect 48145 24157 48179 24191
rect 1409 24021 1443 24055
rect 1409 23477 1443 23511
rect 48145 23477 48179 23511
rect 48145 22389 48179 22423
rect 1409 21981 1443 22015
rect 48145 21981 48179 22015
rect 1409 21301 1443 21335
rect 1409 20893 1443 20927
rect 48145 20893 48179 20927
rect 1409 19805 1443 19839
rect 1409 19125 1443 19159
rect 48145 19125 48179 19159
rect 1409 18717 1443 18751
rect 48145 18581 48179 18615
rect 48145 18037 48179 18071
rect 48145 16949 48179 16983
rect 48145 16541 48179 16575
rect 1409 15861 1443 15895
rect 48145 15861 48179 15895
rect 1409 15453 1443 15487
rect 22937 14977 22971 15011
rect 22753 14773 22787 14807
rect 41613 14433 41647 14467
rect 42625 14433 42659 14467
rect 1409 14365 1443 14399
rect 38393 14365 38427 14399
rect 39865 14365 39899 14399
rect 48145 14365 48179 14399
rect 39037 14297 39071 14331
rect 40141 14297 40175 14331
rect 25145 14229 25179 14263
rect 43269 14229 43303 14263
rect 24961 13957 24995 13991
rect 43545 13957 43579 13991
rect 34805 13889 34839 13923
rect 24685 13821 24719 13855
rect 27905 13821 27939 13855
rect 29653 13821 29687 13855
rect 43269 13821 43303 13855
rect 45017 13821 45051 13855
rect 1409 13685 1443 13719
rect 26433 13685 26467 13719
rect 28162 13685 28196 13719
rect 33333 13685 33367 13719
rect 48145 13685 48179 13719
rect 27997 13481 28031 13515
rect 36645 13481 36679 13515
rect 27353 13345 27387 13379
rect 32413 13345 32447 13379
rect 22661 13277 22695 13311
rect 34897 13277 34931 13311
rect 48145 13277 48179 13311
rect 33057 13209 33091 13243
rect 35173 13209 35207 13243
rect 22477 13141 22511 13175
rect 29101 12937 29135 12971
rect 45109 12937 45143 12971
rect 46397 12937 46431 12971
rect 47685 12937 47719 12971
rect 30389 12869 30423 12903
rect 33793 12869 33827 12903
rect 41061 12801 41095 12835
rect 45201 12801 45235 12835
rect 45845 12801 45879 12835
rect 46489 12801 46523 12835
rect 47593 12801 47627 12835
rect 45753 12733 45787 12767
rect 40969 12665 41003 12699
rect 1409 12597 1443 12631
rect 35265 12597 35299 12631
rect 48145 12189 48179 12223
rect 1409 11645 1443 11679
rect 48145 11509 48179 11543
rect 47409 11305 47443 11339
rect 46949 11169 46983 11203
rect 47041 11169 47075 11203
rect 47225 11101 47259 11135
rect 1409 11033 1443 11067
rect 47593 10761 47627 10795
rect 47593 10625 47627 10659
rect 47777 10625 47811 10659
rect 48145 10013 48179 10047
rect 46305 9537 46339 9571
rect 46121 9401 46155 9435
rect 1409 8925 1443 8959
rect 48145 8925 48179 8959
rect 1409 8313 1443 8347
rect 47961 8041 47995 8075
rect 48145 7837 48179 7871
rect 1409 7701 1443 7735
rect 1409 7293 1443 7327
rect 48145 7293 48179 7327
rect 1409 6205 1443 6239
rect 48145 6069 48179 6103
rect 1409 5661 1443 5695
rect 1409 4981 1443 5015
rect 48145 4981 48179 5015
rect 48145 4573 48179 4607
rect 1409 3893 1443 3927
rect 47041 3893 47075 3927
rect 48145 3893 48179 3927
rect 2053 3553 2087 3587
rect 1409 3485 1443 3519
rect 2697 3485 2731 3519
rect 46857 3485 46891 3519
rect 48145 3485 48179 3519
rect 47501 3349 47535 3383
rect 45753 3145 45787 3179
rect 45569 3009 45603 3043
rect 2697 2941 2731 2975
rect 3985 2941 4019 2975
rect 31033 2941 31067 2975
rect 36185 2941 36219 2975
rect 47041 2941 47075 2975
rect 47777 2941 47811 2975
rect 2053 2873 2087 2907
rect 1409 2805 1443 2839
rect 9137 2805 9171 2839
rect 16865 2805 16899 2839
rect 19441 2805 19475 2839
rect 23305 2805 23339 2839
rect 28457 2805 28491 2839
rect 43913 2805 43947 2839
rect 46397 2805 46431 2839
rect 1409 2397 1443 2431
rect 2605 2397 2639 2431
rect 3249 2397 3283 2431
rect 5181 2397 5215 2431
rect 5825 2397 5859 2431
rect 7113 2397 7147 2431
rect 7757 2397 7791 2431
rect 8401 2397 8435 2431
rect 10333 2397 10367 2431
rect 10977 2397 11011 2431
rect 13001 2397 13035 2431
rect 14105 2397 14139 2431
rect 14933 2397 14967 2431
rect 17417 2397 17451 2431
rect 18061 2397 18095 2431
rect 18705 2397 18739 2431
rect 19993 2397 20027 2431
rect 20637 2397 20671 2431
rect 22201 2397 22235 2431
rect 22937 2397 22971 2431
rect 23857 2397 23891 2431
rect 24593 2397 24627 2431
rect 25237 2397 25271 2431
rect 25881 2397 25915 2431
rect 26985 2397 27019 2431
rect 29561 2397 29595 2431
rect 30205 2397 30239 2431
rect 30849 2397 30883 2431
rect 33609 2397 33643 2431
rect 34713 2397 34747 2431
rect 35357 2397 35391 2431
rect 37473 2397 37507 2431
rect 38761 2397 38795 2431
rect 39865 2397 39899 2431
rect 40693 2397 40727 2431
rect 41337 2397 41371 2431
rect 43085 2397 43119 2431
rect 46489 2397 46523 2431
rect 47593 2397 47627 2431
rect 4537 2261 4571 2295
rect 9689 2261 9723 2295
rect 11713 2261 11747 2295
rect 12357 2261 12391 2295
rect 16129 2261 16163 2295
rect 21281 2261 21315 2295
rect 22017 2261 22051 2295
rect 22753 2261 22787 2295
rect 27629 2261 27663 2295
rect 28273 2261 28307 2295
rect 32321 2261 32355 2295
rect 32965 2261 32999 2295
rect 36001 2261 36035 2295
rect 42441 2261 42475 2295
rect 43729 2261 43763 2295
rect 45017 2261 45051 2295
rect 45661 2261 45695 2295
<< metal1 >>
rect 1104 27770 48852 27792
rect 1104 27718 6924 27770
rect 6976 27718 6988 27770
rect 7040 27718 7052 27770
rect 7104 27718 7116 27770
rect 7168 27718 7180 27770
rect 7232 27718 18872 27770
rect 18924 27718 18936 27770
rect 18988 27718 19000 27770
rect 19052 27718 19064 27770
rect 19116 27718 19128 27770
rect 19180 27718 30820 27770
rect 30872 27718 30884 27770
rect 30936 27718 30948 27770
rect 31000 27718 31012 27770
rect 31064 27718 31076 27770
rect 31128 27718 42768 27770
rect 42820 27718 42832 27770
rect 42884 27718 42896 27770
rect 42948 27718 42960 27770
rect 43012 27718 43024 27770
rect 43076 27718 48852 27770
rect 1104 27696 48852 27718
rect 2038 27588 2044 27600
rect 1999 27560 2044 27588
rect 2038 27548 2044 27560
rect 2096 27548 2102 27600
rect 3970 27588 3976 27600
rect 3931 27560 3976 27588
rect 3970 27548 3976 27560
rect 4028 27548 4034 27600
rect 5166 27588 5172 27600
rect 5127 27560 5172 27588
rect 5166 27548 5172 27560
rect 5224 27548 5230 27600
rect 5810 27588 5816 27600
rect 5771 27560 5816 27588
rect 5810 27548 5816 27560
rect 5868 27548 5874 27600
rect 7742 27588 7748 27600
rect 7703 27560 7748 27588
rect 7742 27548 7748 27560
rect 7800 27548 7806 27600
rect 8386 27588 8392 27600
rect 8347 27560 8392 27588
rect 8386 27548 8392 27560
rect 8444 27548 8450 27600
rect 10318 27588 10324 27600
rect 10279 27560 10324 27588
rect 10318 27548 10324 27560
rect 10376 27548 10382 27600
rect 10962 27588 10968 27600
rect 10923 27560 10968 27588
rect 10962 27548 10968 27560
rect 11020 27548 11026 27600
rect 13814 27548 13820 27600
rect 13872 27588 13878 27600
rect 14093 27591 14151 27597
rect 14093 27588 14105 27591
rect 13872 27560 14105 27588
rect 13872 27548 13878 27560
rect 14093 27557 14105 27560
rect 14139 27557 14151 27591
rect 14918 27588 14924 27600
rect 14879 27560 14924 27588
rect 14093 27551 14151 27557
rect 14918 27548 14924 27560
rect 14976 27548 14982 27600
rect 15562 27588 15568 27600
rect 15523 27560 15568 27588
rect 15562 27548 15568 27560
rect 15620 27548 15626 27600
rect 18046 27588 18052 27600
rect 18007 27560 18052 27588
rect 18046 27548 18052 27560
rect 18104 27548 18110 27600
rect 18690 27588 18696 27600
rect 18651 27560 18696 27588
rect 18690 27548 18696 27560
rect 18748 27548 18754 27600
rect 19978 27588 19984 27600
rect 19939 27560 19984 27588
rect 19978 27548 19984 27560
rect 20036 27548 20042 27600
rect 20622 27588 20628 27600
rect 20583 27560 20628 27588
rect 20622 27548 20628 27560
rect 20680 27548 20686 27600
rect 21266 27588 21272 27600
rect 21227 27560 21272 27588
rect 21266 27548 21272 27560
rect 21324 27548 21330 27600
rect 23198 27588 23204 27600
rect 23159 27560 23204 27588
rect 23198 27548 23204 27560
rect 23256 27548 23262 27600
rect 24578 27588 24584 27600
rect 24539 27560 24584 27588
rect 24578 27548 24584 27560
rect 24636 27548 24642 27600
rect 25222 27588 25228 27600
rect 25183 27560 25228 27588
rect 25222 27548 25228 27560
rect 25280 27548 25286 27600
rect 25866 27588 25872 27600
rect 25827 27560 25872 27588
rect 25866 27548 25872 27560
rect 25924 27548 25930 27600
rect 26418 27548 26424 27600
rect 26476 27588 26482 27600
rect 26973 27591 27031 27597
rect 26973 27588 26985 27591
rect 26476 27560 26985 27588
rect 26476 27548 26482 27560
rect 26973 27557 26985 27560
rect 27019 27557 27031 27591
rect 30374 27588 30380 27600
rect 30335 27560 30380 27588
rect 26973 27551 27031 27557
rect 30374 27548 30380 27560
rect 30432 27548 30438 27600
rect 31021 27591 31079 27597
rect 31021 27557 31033 27591
rect 31067 27588 31079 27591
rect 31202 27588 31208 27600
rect 31067 27560 31208 27588
rect 31067 27557 31079 27560
rect 31021 27551 31079 27557
rect 31202 27548 31208 27560
rect 31260 27548 31266 27600
rect 32306 27588 32312 27600
rect 32267 27560 32312 27588
rect 32306 27548 32312 27560
rect 32364 27548 32370 27600
rect 33594 27588 33600 27600
rect 33555 27560 33600 27588
rect 33594 27548 33600 27560
rect 33652 27548 33658 27600
rect 34514 27548 34520 27600
rect 34572 27588 34578 27600
rect 34701 27591 34759 27597
rect 34701 27588 34713 27591
rect 34572 27560 34713 27588
rect 34572 27548 34578 27560
rect 34701 27557 34713 27560
rect 34747 27557 34759 27591
rect 37274 27588 37280 27600
rect 37235 27560 37280 27588
rect 34701 27551 34759 27557
rect 37274 27548 37280 27560
rect 37332 27548 37338 27600
rect 37366 27548 37372 27600
rect 37424 27588 37430 27600
rect 37921 27591 37979 27597
rect 37921 27588 37933 27591
rect 37424 27560 37933 27588
rect 37424 27548 37430 27560
rect 37921 27557 37933 27560
rect 37967 27557 37979 27591
rect 37921 27551 37979 27557
rect 38010 27548 38016 27600
rect 38068 27588 38074 27600
rect 38565 27591 38623 27597
rect 38565 27588 38577 27591
rect 38068 27560 38577 27588
rect 38068 27548 38074 27560
rect 38565 27557 38577 27560
rect 38611 27557 38623 27591
rect 40034 27588 40040 27600
rect 39995 27560 40040 27588
rect 38565 27551 38623 27557
rect 40034 27548 40040 27560
rect 40092 27548 40098 27600
rect 41322 27588 41328 27600
rect 41283 27560 41328 27588
rect 41322 27548 41328 27560
rect 41380 27548 41386 27600
rect 43162 27548 43168 27600
rect 43220 27588 43226 27600
rect 43901 27591 43959 27597
rect 43901 27588 43913 27591
rect 43220 27560 43913 27588
rect 43220 27548 43226 27560
rect 43901 27557 43913 27560
rect 43947 27557 43959 27591
rect 45186 27588 45192 27600
rect 45147 27560 45192 27588
rect 43901 27551 43959 27557
rect 45186 27548 45192 27560
rect 45244 27548 45250 27600
rect 45830 27588 45836 27600
rect 45791 27560 45836 27588
rect 45830 27548 45836 27560
rect 45888 27548 45894 27600
rect 46474 27588 46480 27600
rect 46435 27560 46480 27588
rect 46474 27548 46480 27560
rect 46532 27548 46538 27600
rect 1302 27480 1308 27532
rect 1360 27520 1366 27532
rect 1397 27523 1455 27529
rect 1397 27520 1409 27523
rect 1360 27492 1409 27520
rect 1360 27480 1366 27492
rect 1397 27489 1409 27492
rect 1443 27489 1455 27523
rect 1397 27483 1455 27489
rect 7101 27523 7159 27529
rect 7101 27489 7113 27523
rect 7147 27520 7159 27523
rect 7282 27520 7288 27532
rect 7147 27492 7288 27520
rect 7147 27489 7159 27492
rect 7101 27483 7159 27489
rect 7282 27480 7288 27492
rect 7340 27480 7346 27532
rect 9674 27480 9680 27532
rect 9732 27520 9738 27532
rect 11698 27520 11704 27532
rect 9732 27492 9777 27520
rect 11659 27492 11704 27520
rect 9732 27480 9738 27492
rect 11698 27480 11704 27492
rect 11756 27480 11762 27532
rect 12342 27520 12348 27532
rect 12303 27492 12348 27520
rect 12342 27480 12348 27492
rect 12400 27480 12406 27532
rect 12986 27520 12992 27532
rect 12947 27492 12992 27520
rect 12986 27480 12992 27492
rect 13044 27480 13050 27532
rect 16574 27480 16580 27532
rect 16632 27520 16638 27532
rect 16669 27523 16727 27529
rect 16669 27520 16681 27523
rect 16632 27492 16681 27520
rect 16632 27480 16638 27492
rect 16669 27489 16681 27492
rect 16715 27489 16727 27523
rect 22554 27520 22560 27532
rect 22515 27492 22560 27520
rect 16669 27483 16727 27489
rect 22554 27480 22560 27492
rect 22612 27480 22618 27532
rect 23842 27520 23848 27532
rect 23803 27492 23848 27520
rect 23842 27480 23848 27492
rect 23900 27480 23906 27532
rect 27798 27520 27804 27532
rect 27759 27492 27804 27520
rect 27798 27480 27804 27492
rect 27856 27480 27862 27532
rect 28442 27520 28448 27532
rect 28403 27492 28448 27520
rect 28442 27480 28448 27492
rect 28500 27480 28506 27532
rect 28994 27480 29000 27532
rect 29052 27520 29058 27532
rect 29549 27523 29607 27529
rect 29549 27520 29561 27523
rect 29052 27492 29561 27520
rect 29052 27480 29058 27492
rect 29549 27489 29561 27492
rect 29595 27489 29607 27523
rect 29549 27483 29607 27489
rect 34790 27480 34796 27532
rect 34848 27520 34854 27532
rect 35345 27523 35403 27529
rect 35345 27520 35357 27523
rect 34848 27492 35357 27520
rect 34848 27480 34854 27492
rect 35345 27489 35357 27492
rect 35391 27489 35403 27523
rect 35345 27483 35403 27489
rect 35894 27480 35900 27532
rect 35952 27520 35958 27532
rect 35989 27523 36047 27529
rect 35989 27520 36001 27523
rect 35952 27492 36001 27520
rect 35952 27480 35958 27492
rect 35989 27489 36001 27492
rect 36035 27489 36047 27523
rect 40678 27520 40684 27532
rect 40639 27492 40684 27520
rect 35989 27483 36047 27489
rect 40678 27480 40684 27492
rect 40736 27480 40742 27532
rect 42610 27520 42616 27532
rect 42571 27492 42616 27520
rect 42610 27480 42616 27492
rect 42668 27480 42674 27532
rect 14 27412 20 27464
rect 72 27452 78 27464
rect 2685 27455 2743 27461
rect 2685 27452 2697 27455
rect 72 27424 2697 27452
rect 72 27412 78 27424
rect 2685 27421 2697 27424
rect 2731 27421 2743 27455
rect 42889 27455 42947 27461
rect 42889 27452 42901 27455
rect 2685 27415 2743 27421
rect 38626 27424 42901 27452
rect 22922 27344 22928 27396
rect 22980 27384 22986 27396
rect 38626 27384 38654 27424
rect 42889 27421 42901 27424
rect 42935 27421 42947 27455
rect 42889 27415 42947 27421
rect 47394 27412 47400 27464
rect 47452 27452 47458 27464
rect 47857 27455 47915 27461
rect 47857 27452 47869 27455
rect 47452 27424 47869 27452
rect 47452 27412 47458 27424
rect 47857 27421 47869 27424
rect 47903 27421 47915 27455
rect 47857 27415 47915 27421
rect 22980 27356 38654 27384
rect 22980 27344 22986 27356
rect 48041 27319 48099 27325
rect 48041 27285 48053 27319
rect 48087 27316 48099 27319
rect 48314 27316 48320 27328
rect 48087 27288 48320 27316
rect 48087 27285 48099 27288
rect 48041 27279 48099 27285
rect 48314 27276 48320 27288
rect 48372 27276 48378 27328
rect 1104 27226 48852 27248
rect 1104 27174 12898 27226
rect 12950 27174 12962 27226
rect 13014 27174 13026 27226
rect 13078 27174 13090 27226
rect 13142 27174 13154 27226
rect 13206 27174 24846 27226
rect 24898 27174 24910 27226
rect 24962 27174 24974 27226
rect 25026 27174 25038 27226
rect 25090 27174 25102 27226
rect 25154 27174 36794 27226
rect 36846 27174 36858 27226
rect 36910 27174 36922 27226
rect 36974 27174 36986 27226
rect 37038 27174 37050 27226
rect 37102 27174 48852 27226
rect 1104 27152 48852 27174
rect 658 27072 664 27124
rect 716 27112 722 27124
rect 2685 27115 2743 27121
rect 2685 27112 2697 27115
rect 716 27084 2697 27112
rect 716 27072 722 27084
rect 2685 27081 2697 27084
rect 2731 27081 2743 27115
rect 2685 27075 2743 27081
rect 47026 27072 47032 27124
rect 47084 27112 47090 27124
rect 47581 27115 47639 27121
rect 47581 27112 47593 27115
rect 47084 27084 47593 27112
rect 47084 27072 47090 27084
rect 47581 27081 47593 27084
rect 47627 27081 47639 27115
rect 47581 27075 47639 27081
rect 2041 27047 2099 27053
rect 2041 27013 2053 27047
rect 2087 27044 2099 27047
rect 2866 27044 2872 27056
rect 2087 27016 2872 27044
rect 2087 27013 2099 27016
rect 2041 27007 2099 27013
rect 2866 27004 2872 27016
rect 2924 27004 2930 27056
rect 1394 26976 1400 26988
rect 1355 26948 1400 26976
rect 1394 26936 1400 26948
rect 1452 26936 1458 26988
rect 6546 26976 6552 26988
rect 6507 26948 6552 26976
rect 6546 26936 6552 26948
rect 6604 26936 6610 26988
rect 9122 26976 9128 26988
rect 9083 26948 9128 26976
rect 9122 26936 9128 26948
rect 9180 26936 9186 26988
rect 19426 26976 19432 26988
rect 19387 26948 19432 26976
rect 19426 26936 19432 26948
rect 19484 26936 19490 26988
rect 22002 26976 22008 26988
rect 21963 26948 22008 26976
rect 22002 26936 22008 26948
rect 22060 26936 22066 26988
rect 36170 26976 36176 26988
rect 36131 26948 36176 26976
rect 36170 26936 36176 26948
rect 36228 26936 36234 26988
rect 38746 26976 38752 26988
rect 38707 26948 38752 26976
rect 38746 26936 38752 26948
rect 38804 26936 38810 26988
rect 41874 26936 41880 26988
rect 41932 26976 41938 26988
rect 42429 26979 42487 26985
rect 42429 26976 42441 26979
rect 41932 26948 42441 26976
rect 41932 26936 41938 26948
rect 42429 26945 42441 26948
rect 42475 26945 42487 26979
rect 43898 26976 43904 26988
rect 43859 26948 43904 26976
rect 42429 26939 42487 26945
rect 43898 26936 43904 26948
rect 43956 26936 43962 26988
rect 45738 26976 45744 26988
rect 45699 26948 45744 26976
rect 45738 26936 45744 26948
rect 45796 26936 45802 26988
rect 47029 26979 47087 26985
rect 47029 26945 47041 26979
rect 47075 26976 47087 26979
rect 47670 26976 47676 26988
rect 47075 26948 47676 26976
rect 47075 26945 47087 26948
rect 47029 26939 47087 26945
rect 47670 26936 47676 26948
rect 47728 26936 47734 26988
rect 46385 26911 46443 26917
rect 46385 26877 46397 26911
rect 46431 26908 46443 26911
rect 48958 26908 48964 26920
rect 46431 26880 48964 26908
rect 46431 26877 46443 26880
rect 46385 26871 46443 26877
rect 48958 26868 48964 26880
rect 49016 26868 49022 26920
rect 1104 26682 48852 26704
rect 1104 26630 6924 26682
rect 6976 26630 6988 26682
rect 7040 26630 7052 26682
rect 7104 26630 7116 26682
rect 7168 26630 7180 26682
rect 7232 26630 18872 26682
rect 18924 26630 18936 26682
rect 18988 26630 19000 26682
rect 19052 26630 19064 26682
rect 19116 26630 19128 26682
rect 19180 26630 30820 26682
rect 30872 26630 30884 26682
rect 30936 26630 30948 26682
rect 31000 26630 31012 26682
rect 31064 26630 31076 26682
rect 31128 26630 42768 26682
rect 42820 26630 42832 26682
rect 42884 26630 42896 26682
rect 42948 26630 42960 26682
rect 43012 26630 43024 26682
rect 43076 26630 48852 26682
rect 1104 26608 48852 26630
rect 2041 26571 2099 26577
rect 2041 26537 2053 26571
rect 2087 26568 2099 26571
rect 2774 26568 2780 26580
rect 2087 26540 2780 26568
rect 2087 26537 2099 26540
rect 2041 26531 2099 26537
rect 2774 26528 2780 26540
rect 2832 26528 2838 26580
rect 47486 26568 47492 26580
rect 47447 26540 47492 26568
rect 47486 26528 47492 26540
rect 47544 26528 47550 26580
rect 46842 26432 46848 26444
rect 46803 26404 46848 26432
rect 46842 26392 46848 26404
rect 46900 26392 46906 26444
rect 1394 26364 1400 26376
rect 1355 26336 1400 26364
rect 1394 26324 1400 26336
rect 1452 26324 1458 26376
rect 48133 26231 48191 26237
rect 48133 26197 48145 26231
rect 48179 26228 48191 26231
rect 48222 26228 48228 26240
rect 48179 26200 48228 26228
rect 48179 26197 48191 26200
rect 48133 26191 48191 26197
rect 48222 26188 48228 26200
rect 48280 26188 48286 26240
rect 1104 26138 48852 26160
rect 1104 26086 12898 26138
rect 12950 26086 12962 26138
rect 13014 26086 13026 26138
rect 13078 26086 13090 26138
rect 13142 26086 13154 26138
rect 13206 26086 24846 26138
rect 24898 26086 24910 26138
rect 24962 26086 24974 26138
rect 25026 26086 25038 26138
rect 25090 26086 25102 26138
rect 25154 26086 36794 26138
rect 36846 26086 36858 26138
rect 36910 26086 36922 26138
rect 36974 26086 36986 26138
rect 37038 26086 37050 26138
rect 37102 26086 48852 26138
rect 1104 26064 48852 26086
rect 1397 25891 1455 25897
rect 1397 25857 1409 25891
rect 1443 25888 1455 25891
rect 1486 25888 1492 25900
rect 1443 25860 1492 25888
rect 1443 25857 1455 25860
rect 1397 25851 1455 25857
rect 1486 25848 1492 25860
rect 1544 25848 1550 25900
rect 48130 25888 48136 25900
rect 48091 25860 48136 25888
rect 48130 25848 48136 25860
rect 48188 25848 48194 25900
rect 47029 25823 47087 25829
rect 47029 25789 47041 25823
rect 47075 25820 47087 25823
rect 49602 25820 49608 25832
rect 47075 25792 49608 25820
rect 47075 25789 47087 25792
rect 47029 25783 47087 25789
rect 49602 25780 49608 25792
rect 49660 25780 49666 25832
rect 1104 25594 48852 25616
rect 1104 25542 6924 25594
rect 6976 25542 6988 25594
rect 7040 25542 7052 25594
rect 7104 25542 7116 25594
rect 7168 25542 7180 25594
rect 7232 25542 18872 25594
rect 18924 25542 18936 25594
rect 18988 25542 19000 25594
rect 19052 25542 19064 25594
rect 19116 25542 19128 25594
rect 19180 25542 30820 25594
rect 30872 25542 30884 25594
rect 30936 25542 30948 25594
rect 31000 25542 31012 25594
rect 31064 25542 31076 25594
rect 31128 25542 42768 25594
rect 42820 25542 42832 25594
rect 42884 25542 42896 25594
rect 42948 25542 42960 25594
rect 43012 25542 43024 25594
rect 43076 25542 48852 25594
rect 1104 25520 48852 25542
rect 1394 25276 1400 25288
rect 1355 25248 1400 25276
rect 1394 25236 1400 25248
rect 1452 25236 1458 25288
rect 48130 25276 48136 25288
rect 48091 25248 48136 25276
rect 48130 25236 48136 25248
rect 48188 25236 48194 25288
rect 1104 25050 48852 25072
rect 1104 24998 12898 25050
rect 12950 24998 12962 25050
rect 13014 24998 13026 25050
rect 13078 24998 13090 25050
rect 13142 24998 13154 25050
rect 13206 24998 24846 25050
rect 24898 24998 24910 25050
rect 24962 24998 24974 25050
rect 25026 24998 25038 25050
rect 25090 24998 25102 25050
rect 25154 24998 36794 25050
rect 36846 24998 36858 25050
rect 36910 24998 36922 25050
rect 36974 24998 36986 25050
rect 37038 24998 37050 25050
rect 37102 24998 48852 25050
rect 1104 24976 48852 24998
rect 1394 24596 1400 24608
rect 1355 24568 1400 24596
rect 1394 24556 1400 24568
rect 1452 24556 1458 24608
rect 48130 24596 48136 24608
rect 48091 24568 48136 24596
rect 48130 24556 48136 24568
rect 48188 24556 48194 24608
rect 1104 24506 48852 24528
rect 1104 24454 6924 24506
rect 6976 24454 6988 24506
rect 7040 24454 7052 24506
rect 7104 24454 7116 24506
rect 7168 24454 7180 24506
rect 7232 24454 18872 24506
rect 18924 24454 18936 24506
rect 18988 24454 19000 24506
rect 19052 24454 19064 24506
rect 19116 24454 19128 24506
rect 19180 24454 30820 24506
rect 30872 24454 30884 24506
rect 30936 24454 30948 24506
rect 31000 24454 31012 24506
rect 31064 24454 31076 24506
rect 31128 24454 42768 24506
rect 42820 24454 42832 24506
rect 42884 24454 42896 24506
rect 42948 24454 42960 24506
rect 43012 24454 43024 24506
rect 43076 24454 48852 24506
rect 1104 24432 48852 24454
rect 48133 24191 48191 24197
rect 48133 24157 48145 24191
rect 48179 24188 48191 24191
rect 48222 24188 48228 24200
rect 48179 24160 48228 24188
rect 48179 24157 48191 24160
rect 48133 24151 48191 24157
rect 48222 24148 48228 24160
rect 48280 24148 48286 24200
rect 1394 24052 1400 24064
rect 1355 24024 1400 24052
rect 1394 24012 1400 24024
rect 1452 24012 1458 24064
rect 1104 23962 48852 23984
rect 1104 23910 12898 23962
rect 12950 23910 12962 23962
rect 13014 23910 13026 23962
rect 13078 23910 13090 23962
rect 13142 23910 13154 23962
rect 13206 23910 24846 23962
rect 24898 23910 24910 23962
rect 24962 23910 24974 23962
rect 25026 23910 25038 23962
rect 25090 23910 25102 23962
rect 25154 23910 36794 23962
rect 36846 23910 36858 23962
rect 36910 23910 36922 23962
rect 36974 23910 36986 23962
rect 37038 23910 37050 23962
rect 37102 23910 48852 23962
rect 1104 23888 48852 23910
rect 1394 23508 1400 23520
rect 1355 23480 1400 23508
rect 1394 23468 1400 23480
rect 1452 23468 1458 23520
rect 48130 23508 48136 23520
rect 48091 23480 48136 23508
rect 48130 23468 48136 23480
rect 48188 23468 48194 23520
rect 1104 23418 48852 23440
rect 1104 23366 6924 23418
rect 6976 23366 6988 23418
rect 7040 23366 7052 23418
rect 7104 23366 7116 23418
rect 7168 23366 7180 23418
rect 7232 23366 18872 23418
rect 18924 23366 18936 23418
rect 18988 23366 19000 23418
rect 19052 23366 19064 23418
rect 19116 23366 19128 23418
rect 19180 23366 30820 23418
rect 30872 23366 30884 23418
rect 30936 23366 30948 23418
rect 31000 23366 31012 23418
rect 31064 23366 31076 23418
rect 31128 23366 42768 23418
rect 42820 23366 42832 23418
rect 42884 23366 42896 23418
rect 42948 23366 42960 23418
rect 43012 23366 43024 23418
rect 43076 23366 48852 23418
rect 1104 23344 48852 23366
rect 1104 22874 48852 22896
rect 1104 22822 12898 22874
rect 12950 22822 12962 22874
rect 13014 22822 13026 22874
rect 13078 22822 13090 22874
rect 13142 22822 13154 22874
rect 13206 22822 24846 22874
rect 24898 22822 24910 22874
rect 24962 22822 24974 22874
rect 25026 22822 25038 22874
rect 25090 22822 25102 22874
rect 25154 22822 36794 22874
rect 36846 22822 36858 22874
rect 36910 22822 36922 22874
rect 36974 22822 36986 22874
rect 37038 22822 37050 22874
rect 37102 22822 48852 22874
rect 1104 22800 48852 22822
rect 48130 22420 48136 22432
rect 48091 22392 48136 22420
rect 48130 22380 48136 22392
rect 48188 22380 48194 22432
rect 1104 22330 48852 22352
rect 1104 22278 6924 22330
rect 6976 22278 6988 22330
rect 7040 22278 7052 22330
rect 7104 22278 7116 22330
rect 7168 22278 7180 22330
rect 7232 22278 18872 22330
rect 18924 22278 18936 22330
rect 18988 22278 19000 22330
rect 19052 22278 19064 22330
rect 19116 22278 19128 22330
rect 19180 22278 30820 22330
rect 30872 22278 30884 22330
rect 30936 22278 30948 22330
rect 31000 22278 31012 22330
rect 31064 22278 31076 22330
rect 31128 22278 42768 22330
rect 42820 22278 42832 22330
rect 42884 22278 42896 22330
rect 42948 22278 42960 22330
rect 43012 22278 43024 22330
rect 43076 22278 48852 22330
rect 1104 22256 48852 22278
rect 1394 22012 1400 22024
rect 1355 21984 1400 22012
rect 1394 21972 1400 21984
rect 1452 21972 1458 22024
rect 48130 22012 48136 22024
rect 48091 21984 48136 22012
rect 48130 21972 48136 21984
rect 48188 21972 48194 22024
rect 1104 21786 48852 21808
rect 1104 21734 12898 21786
rect 12950 21734 12962 21786
rect 13014 21734 13026 21786
rect 13078 21734 13090 21786
rect 13142 21734 13154 21786
rect 13206 21734 24846 21786
rect 24898 21734 24910 21786
rect 24962 21734 24974 21786
rect 25026 21734 25038 21786
rect 25090 21734 25102 21786
rect 25154 21734 36794 21786
rect 36846 21734 36858 21786
rect 36910 21734 36922 21786
rect 36974 21734 36986 21786
rect 37038 21734 37050 21786
rect 37102 21734 48852 21786
rect 1104 21712 48852 21734
rect 1394 21332 1400 21344
rect 1355 21304 1400 21332
rect 1394 21292 1400 21304
rect 1452 21292 1458 21344
rect 1104 21242 48852 21264
rect 1104 21190 6924 21242
rect 6976 21190 6988 21242
rect 7040 21190 7052 21242
rect 7104 21190 7116 21242
rect 7168 21190 7180 21242
rect 7232 21190 18872 21242
rect 18924 21190 18936 21242
rect 18988 21190 19000 21242
rect 19052 21190 19064 21242
rect 19116 21190 19128 21242
rect 19180 21190 30820 21242
rect 30872 21190 30884 21242
rect 30936 21190 30948 21242
rect 31000 21190 31012 21242
rect 31064 21190 31076 21242
rect 31128 21190 42768 21242
rect 42820 21190 42832 21242
rect 42884 21190 42896 21242
rect 42948 21190 42960 21242
rect 43012 21190 43024 21242
rect 43076 21190 48852 21242
rect 1104 21168 48852 21190
rect 1394 20924 1400 20936
rect 1355 20896 1400 20924
rect 1394 20884 1400 20896
rect 1452 20884 1458 20936
rect 48133 20927 48191 20933
rect 48133 20893 48145 20927
rect 48179 20924 48191 20927
rect 48222 20924 48228 20936
rect 48179 20896 48228 20924
rect 48179 20893 48191 20896
rect 48133 20887 48191 20893
rect 48222 20884 48228 20896
rect 48280 20884 48286 20936
rect 1104 20698 48852 20720
rect 1104 20646 12898 20698
rect 12950 20646 12962 20698
rect 13014 20646 13026 20698
rect 13078 20646 13090 20698
rect 13142 20646 13154 20698
rect 13206 20646 24846 20698
rect 24898 20646 24910 20698
rect 24962 20646 24974 20698
rect 25026 20646 25038 20698
rect 25090 20646 25102 20698
rect 25154 20646 36794 20698
rect 36846 20646 36858 20698
rect 36910 20646 36922 20698
rect 36974 20646 36986 20698
rect 37038 20646 37050 20698
rect 37102 20646 48852 20698
rect 1104 20624 48852 20646
rect 1104 20154 48852 20176
rect 1104 20102 6924 20154
rect 6976 20102 6988 20154
rect 7040 20102 7052 20154
rect 7104 20102 7116 20154
rect 7168 20102 7180 20154
rect 7232 20102 18872 20154
rect 18924 20102 18936 20154
rect 18988 20102 19000 20154
rect 19052 20102 19064 20154
rect 19116 20102 19128 20154
rect 19180 20102 30820 20154
rect 30872 20102 30884 20154
rect 30936 20102 30948 20154
rect 31000 20102 31012 20154
rect 31064 20102 31076 20154
rect 31128 20102 42768 20154
rect 42820 20102 42832 20154
rect 42884 20102 42896 20154
rect 42948 20102 42960 20154
rect 43012 20102 43024 20154
rect 43076 20102 48852 20154
rect 1104 20080 48852 20102
rect 1394 19836 1400 19848
rect 1355 19808 1400 19836
rect 1394 19796 1400 19808
rect 1452 19796 1458 19848
rect 1104 19610 48852 19632
rect 1104 19558 12898 19610
rect 12950 19558 12962 19610
rect 13014 19558 13026 19610
rect 13078 19558 13090 19610
rect 13142 19558 13154 19610
rect 13206 19558 24846 19610
rect 24898 19558 24910 19610
rect 24962 19558 24974 19610
rect 25026 19558 25038 19610
rect 25090 19558 25102 19610
rect 25154 19558 36794 19610
rect 36846 19558 36858 19610
rect 36910 19558 36922 19610
rect 36974 19558 36986 19610
rect 37038 19558 37050 19610
rect 37102 19558 48852 19610
rect 1104 19536 48852 19558
rect 1394 19156 1400 19168
rect 1355 19128 1400 19156
rect 1394 19116 1400 19128
rect 1452 19116 1458 19168
rect 48130 19156 48136 19168
rect 48091 19128 48136 19156
rect 48130 19116 48136 19128
rect 48188 19116 48194 19168
rect 1104 19066 48852 19088
rect 1104 19014 6924 19066
rect 6976 19014 6988 19066
rect 7040 19014 7052 19066
rect 7104 19014 7116 19066
rect 7168 19014 7180 19066
rect 7232 19014 18872 19066
rect 18924 19014 18936 19066
rect 18988 19014 19000 19066
rect 19052 19014 19064 19066
rect 19116 19014 19128 19066
rect 19180 19014 30820 19066
rect 30872 19014 30884 19066
rect 30936 19014 30948 19066
rect 31000 19014 31012 19066
rect 31064 19014 31076 19066
rect 31128 19014 42768 19066
rect 42820 19014 42832 19066
rect 42884 19014 42896 19066
rect 42948 19014 42960 19066
rect 43012 19014 43024 19066
rect 43076 19014 48852 19066
rect 1104 18992 48852 19014
rect 1394 18748 1400 18760
rect 1355 18720 1400 18748
rect 1394 18708 1400 18720
rect 1452 18708 1458 18760
rect 48133 18615 48191 18621
rect 48133 18581 48145 18615
rect 48179 18612 48191 18615
rect 48222 18612 48228 18624
rect 48179 18584 48228 18612
rect 48179 18581 48191 18584
rect 48133 18575 48191 18581
rect 48222 18572 48228 18584
rect 48280 18572 48286 18624
rect 1104 18522 48852 18544
rect 1104 18470 12898 18522
rect 12950 18470 12962 18522
rect 13014 18470 13026 18522
rect 13078 18470 13090 18522
rect 13142 18470 13154 18522
rect 13206 18470 24846 18522
rect 24898 18470 24910 18522
rect 24962 18470 24974 18522
rect 25026 18470 25038 18522
rect 25090 18470 25102 18522
rect 25154 18470 36794 18522
rect 36846 18470 36858 18522
rect 36910 18470 36922 18522
rect 36974 18470 36986 18522
rect 37038 18470 37050 18522
rect 37102 18470 48852 18522
rect 1104 18448 48852 18470
rect 48130 18068 48136 18080
rect 48091 18040 48136 18068
rect 48130 18028 48136 18040
rect 48188 18028 48194 18080
rect 1104 17978 48852 18000
rect 1104 17926 6924 17978
rect 6976 17926 6988 17978
rect 7040 17926 7052 17978
rect 7104 17926 7116 17978
rect 7168 17926 7180 17978
rect 7232 17926 18872 17978
rect 18924 17926 18936 17978
rect 18988 17926 19000 17978
rect 19052 17926 19064 17978
rect 19116 17926 19128 17978
rect 19180 17926 30820 17978
rect 30872 17926 30884 17978
rect 30936 17926 30948 17978
rect 31000 17926 31012 17978
rect 31064 17926 31076 17978
rect 31128 17926 42768 17978
rect 42820 17926 42832 17978
rect 42884 17926 42896 17978
rect 42948 17926 42960 17978
rect 43012 17926 43024 17978
rect 43076 17926 48852 17978
rect 1104 17904 48852 17926
rect 1104 17434 48852 17456
rect 1104 17382 12898 17434
rect 12950 17382 12962 17434
rect 13014 17382 13026 17434
rect 13078 17382 13090 17434
rect 13142 17382 13154 17434
rect 13206 17382 24846 17434
rect 24898 17382 24910 17434
rect 24962 17382 24974 17434
rect 25026 17382 25038 17434
rect 25090 17382 25102 17434
rect 25154 17382 36794 17434
rect 36846 17382 36858 17434
rect 36910 17382 36922 17434
rect 36974 17382 36986 17434
rect 37038 17382 37050 17434
rect 37102 17382 48852 17434
rect 1104 17360 48852 17382
rect 48130 16980 48136 16992
rect 48091 16952 48136 16980
rect 48130 16940 48136 16952
rect 48188 16940 48194 16992
rect 1104 16890 48852 16912
rect 1104 16838 6924 16890
rect 6976 16838 6988 16890
rect 7040 16838 7052 16890
rect 7104 16838 7116 16890
rect 7168 16838 7180 16890
rect 7232 16838 18872 16890
rect 18924 16838 18936 16890
rect 18988 16838 19000 16890
rect 19052 16838 19064 16890
rect 19116 16838 19128 16890
rect 19180 16838 30820 16890
rect 30872 16838 30884 16890
rect 30936 16838 30948 16890
rect 31000 16838 31012 16890
rect 31064 16838 31076 16890
rect 31128 16838 42768 16890
rect 42820 16838 42832 16890
rect 42884 16838 42896 16890
rect 42948 16838 42960 16890
rect 43012 16838 43024 16890
rect 43076 16838 48852 16890
rect 1104 16816 48852 16838
rect 48133 16575 48191 16581
rect 48133 16541 48145 16575
rect 48179 16572 48191 16575
rect 48222 16572 48228 16584
rect 48179 16544 48228 16572
rect 48179 16541 48191 16544
rect 48133 16535 48191 16541
rect 48222 16532 48228 16544
rect 48280 16532 48286 16584
rect 1104 16346 48852 16368
rect 1104 16294 12898 16346
rect 12950 16294 12962 16346
rect 13014 16294 13026 16346
rect 13078 16294 13090 16346
rect 13142 16294 13154 16346
rect 13206 16294 24846 16346
rect 24898 16294 24910 16346
rect 24962 16294 24974 16346
rect 25026 16294 25038 16346
rect 25090 16294 25102 16346
rect 25154 16294 36794 16346
rect 36846 16294 36858 16346
rect 36910 16294 36922 16346
rect 36974 16294 36986 16346
rect 37038 16294 37050 16346
rect 37102 16294 48852 16346
rect 1104 16272 48852 16294
rect 1394 15892 1400 15904
rect 1355 15864 1400 15892
rect 1394 15852 1400 15864
rect 1452 15852 1458 15904
rect 48130 15892 48136 15904
rect 48091 15864 48136 15892
rect 48130 15852 48136 15864
rect 48188 15852 48194 15904
rect 1104 15802 48852 15824
rect 1104 15750 6924 15802
rect 6976 15750 6988 15802
rect 7040 15750 7052 15802
rect 7104 15750 7116 15802
rect 7168 15750 7180 15802
rect 7232 15750 18872 15802
rect 18924 15750 18936 15802
rect 18988 15750 19000 15802
rect 19052 15750 19064 15802
rect 19116 15750 19128 15802
rect 19180 15750 30820 15802
rect 30872 15750 30884 15802
rect 30936 15750 30948 15802
rect 31000 15750 31012 15802
rect 31064 15750 31076 15802
rect 31128 15750 42768 15802
rect 42820 15750 42832 15802
rect 42884 15750 42896 15802
rect 42948 15750 42960 15802
rect 43012 15750 43024 15802
rect 43076 15750 48852 15802
rect 1104 15728 48852 15750
rect 1394 15484 1400 15496
rect 1355 15456 1400 15484
rect 1394 15444 1400 15456
rect 1452 15444 1458 15496
rect 1104 15258 48852 15280
rect 1104 15206 12898 15258
rect 12950 15206 12962 15258
rect 13014 15206 13026 15258
rect 13078 15206 13090 15258
rect 13142 15206 13154 15258
rect 13206 15206 24846 15258
rect 24898 15206 24910 15258
rect 24962 15206 24974 15258
rect 25026 15206 25038 15258
rect 25090 15206 25102 15258
rect 25154 15206 36794 15258
rect 36846 15206 36858 15258
rect 36910 15206 36922 15258
rect 36974 15206 36986 15258
rect 37038 15206 37050 15258
rect 37102 15206 48852 15258
rect 1104 15184 48852 15206
rect 22922 15008 22928 15020
rect 22883 14980 22928 15008
rect 22922 14968 22928 14980
rect 22980 14968 22986 15020
rect 22741 14807 22799 14813
rect 22741 14773 22753 14807
rect 22787 14804 22799 14807
rect 22922 14804 22928 14816
rect 22787 14776 22928 14804
rect 22787 14773 22799 14776
rect 22741 14767 22799 14773
rect 22922 14764 22928 14776
rect 22980 14764 22986 14816
rect 1104 14714 48852 14736
rect 1104 14662 6924 14714
rect 6976 14662 6988 14714
rect 7040 14662 7052 14714
rect 7104 14662 7116 14714
rect 7168 14662 7180 14714
rect 7232 14662 18872 14714
rect 18924 14662 18936 14714
rect 18988 14662 19000 14714
rect 19052 14662 19064 14714
rect 19116 14662 19128 14714
rect 19180 14662 30820 14714
rect 30872 14662 30884 14714
rect 30936 14662 30948 14714
rect 31000 14662 31012 14714
rect 31064 14662 31076 14714
rect 31128 14662 42768 14714
rect 42820 14662 42832 14714
rect 42884 14662 42896 14714
rect 42948 14662 42960 14714
rect 43012 14662 43024 14714
rect 43076 14662 48852 14714
rect 1104 14640 48852 14662
rect 41601 14467 41659 14473
rect 41601 14433 41613 14467
rect 41647 14464 41659 14467
rect 42613 14467 42671 14473
rect 42613 14464 42625 14467
rect 41647 14436 42625 14464
rect 41647 14433 41659 14436
rect 41601 14427 41659 14433
rect 42613 14433 42625 14436
rect 42659 14433 42671 14467
rect 42613 14427 42671 14433
rect 1394 14396 1400 14408
rect 1355 14368 1400 14396
rect 1394 14356 1400 14368
rect 1452 14356 1458 14408
rect 38378 14396 38384 14408
rect 38339 14368 38384 14396
rect 38378 14356 38384 14368
rect 38436 14356 38442 14408
rect 39850 14396 39856 14408
rect 39811 14368 39856 14396
rect 39850 14356 39856 14368
rect 39908 14356 39914 14408
rect 48130 14396 48136 14408
rect 48091 14368 48136 14396
rect 48130 14356 48136 14368
rect 48188 14356 48194 14408
rect 39025 14331 39083 14337
rect 39025 14297 39037 14331
rect 39071 14328 39083 14331
rect 40129 14331 40187 14337
rect 40129 14328 40141 14331
rect 39071 14300 40141 14328
rect 39071 14297 39083 14300
rect 39025 14291 39083 14297
rect 40129 14297 40141 14300
rect 40175 14297 40187 14331
rect 45094 14328 45100 14340
rect 41354 14300 45100 14328
rect 40129 14291 40187 14297
rect 45094 14288 45100 14300
rect 45152 14288 45158 14340
rect 25133 14263 25191 14269
rect 25133 14229 25145 14263
rect 25179 14260 25191 14263
rect 25222 14260 25228 14272
rect 25179 14232 25228 14260
rect 25179 14229 25191 14232
rect 25133 14223 25191 14229
rect 25222 14220 25228 14232
rect 25280 14220 25286 14272
rect 43254 14260 43260 14272
rect 43215 14232 43260 14260
rect 43254 14220 43260 14232
rect 43312 14220 43318 14272
rect 1104 14170 48852 14192
rect 1104 14118 12898 14170
rect 12950 14118 12962 14170
rect 13014 14118 13026 14170
rect 13078 14118 13090 14170
rect 13142 14118 13154 14170
rect 13206 14118 24846 14170
rect 24898 14118 24910 14170
rect 24962 14118 24974 14170
rect 25026 14118 25038 14170
rect 25090 14118 25102 14170
rect 25154 14118 36794 14170
rect 36846 14118 36858 14170
rect 36910 14118 36922 14170
rect 36974 14118 36986 14170
rect 37038 14118 37050 14170
rect 37102 14118 48852 14170
rect 1104 14096 48852 14118
rect 45554 14056 45560 14068
rect 38626 14028 45560 14056
rect 24949 13991 25007 13997
rect 24949 13957 24961 13991
rect 24995 13988 25007 13991
rect 25222 13988 25228 14000
rect 24995 13960 25228 13988
rect 24995 13957 25007 13960
rect 24949 13951 25007 13957
rect 25222 13948 25228 13960
rect 25280 13948 25286 14000
rect 30282 13988 30288 14000
rect 29394 13960 30288 13988
rect 30282 13948 30288 13960
rect 30340 13948 30346 14000
rect 26050 13880 26056 13932
rect 26108 13880 26114 13932
rect 34793 13923 34851 13929
rect 34793 13889 34805 13923
rect 34839 13920 34851 13923
rect 38626 13920 38654 14028
rect 45554 14016 45560 14028
rect 45612 14016 45618 14068
rect 43254 13948 43260 14000
rect 43312 13988 43318 14000
rect 43533 13991 43591 13997
rect 43533 13988 43545 13991
rect 43312 13960 43545 13988
rect 43312 13948 43318 13960
rect 43533 13957 43545 13960
rect 43579 13957 43591 13991
rect 47670 13988 47676 14000
rect 44758 13960 47676 13988
rect 43533 13951 43591 13957
rect 47670 13948 47676 13960
rect 47728 13948 47734 14000
rect 34839 13892 38654 13920
rect 34839 13889 34851 13892
rect 34793 13883 34851 13889
rect 24670 13852 24676 13864
rect 24631 13824 24676 13852
rect 24670 13812 24676 13824
rect 24728 13852 24734 13864
rect 27893 13855 27951 13861
rect 27893 13852 27905 13855
rect 24728 13824 27905 13852
rect 24728 13812 24734 13824
rect 27893 13821 27905 13824
rect 27939 13852 27951 13855
rect 29178 13852 29184 13864
rect 27939 13824 29184 13852
rect 27939 13821 27951 13824
rect 27893 13815 27951 13821
rect 29178 13812 29184 13824
rect 29236 13812 29242 13864
rect 29641 13855 29699 13861
rect 29641 13821 29653 13855
rect 29687 13852 29699 13855
rect 32398 13852 32404 13864
rect 29687 13824 32404 13852
rect 29687 13821 29699 13824
rect 29641 13815 29699 13821
rect 32398 13812 32404 13824
rect 32456 13812 32462 13864
rect 39850 13812 39856 13864
rect 39908 13852 39914 13864
rect 43257 13855 43315 13861
rect 43257 13852 43269 13855
rect 39908 13824 43269 13852
rect 39908 13812 39914 13824
rect 43257 13821 43269 13824
rect 43303 13821 43315 13855
rect 43257 13815 43315 13821
rect 45005 13855 45063 13861
rect 45005 13821 45017 13855
rect 45051 13852 45063 13855
rect 46934 13852 46940 13864
rect 45051 13824 46940 13852
rect 45051 13821 45063 13824
rect 45005 13815 45063 13821
rect 46934 13812 46940 13824
rect 46992 13812 46998 13864
rect 1394 13716 1400 13728
rect 1355 13688 1400 13716
rect 1394 13676 1400 13688
rect 1452 13676 1458 13728
rect 26418 13716 26424 13728
rect 26379 13688 26424 13716
rect 26418 13676 26424 13688
rect 26476 13676 26482 13728
rect 27982 13676 27988 13728
rect 28040 13716 28046 13728
rect 28150 13719 28208 13725
rect 28150 13716 28162 13719
rect 28040 13688 28162 13716
rect 28040 13676 28046 13688
rect 28150 13685 28162 13688
rect 28196 13685 28208 13719
rect 33318 13716 33324 13728
rect 33279 13688 33324 13716
rect 28150 13679 28208 13685
rect 33318 13676 33324 13688
rect 33376 13676 33382 13728
rect 48133 13719 48191 13725
rect 48133 13685 48145 13719
rect 48179 13716 48191 13719
rect 48222 13716 48228 13728
rect 48179 13688 48228 13716
rect 48179 13685 48191 13688
rect 48133 13679 48191 13685
rect 48222 13676 48228 13688
rect 48280 13676 48286 13728
rect 1104 13626 48852 13648
rect 1104 13574 6924 13626
rect 6976 13574 6988 13626
rect 7040 13574 7052 13626
rect 7104 13574 7116 13626
rect 7168 13574 7180 13626
rect 7232 13574 18872 13626
rect 18924 13574 18936 13626
rect 18988 13574 19000 13626
rect 19052 13574 19064 13626
rect 19116 13574 19128 13626
rect 19180 13574 30820 13626
rect 30872 13574 30884 13626
rect 30936 13574 30948 13626
rect 31000 13574 31012 13626
rect 31064 13574 31076 13626
rect 31128 13574 42768 13626
rect 42820 13574 42832 13626
rect 42884 13574 42896 13626
rect 42948 13574 42960 13626
rect 43012 13574 43024 13626
rect 43076 13574 48852 13626
rect 1104 13552 48852 13574
rect 27982 13512 27988 13524
rect 27943 13484 27988 13512
rect 27982 13472 27988 13484
rect 28040 13472 28046 13524
rect 36633 13515 36691 13521
rect 36633 13481 36645 13515
rect 36679 13512 36691 13515
rect 38378 13512 38384 13524
rect 36679 13484 38384 13512
rect 36679 13481 36691 13484
rect 36633 13475 36691 13481
rect 38378 13472 38384 13484
rect 38436 13472 38442 13524
rect 26418 13336 26424 13388
rect 26476 13376 26482 13388
rect 27341 13379 27399 13385
rect 27341 13376 27353 13379
rect 26476 13348 27353 13376
rect 26476 13336 26482 13348
rect 27341 13345 27353 13348
rect 27387 13345 27399 13379
rect 32398 13376 32404 13388
rect 32359 13348 32404 13376
rect 27341 13339 27399 13345
rect 32398 13336 32404 13348
rect 32456 13336 32462 13388
rect 22649 13311 22707 13317
rect 22649 13277 22661 13311
rect 22695 13308 22707 13311
rect 24670 13308 24676 13320
rect 22695 13280 24676 13308
rect 22695 13277 22707 13280
rect 22649 13271 22707 13277
rect 24670 13268 24676 13280
rect 24728 13268 24734 13320
rect 34882 13308 34888 13320
rect 34843 13280 34888 13308
rect 34882 13268 34888 13280
rect 34940 13268 34946 13320
rect 48130 13308 48136 13320
rect 48091 13280 48136 13308
rect 48130 13268 48136 13280
rect 48188 13268 48194 13320
rect 33045 13243 33103 13249
rect 33045 13209 33057 13243
rect 33091 13240 33103 13243
rect 35161 13243 35219 13249
rect 35161 13240 35173 13243
rect 33091 13212 35173 13240
rect 33091 13209 33103 13212
rect 33045 13203 33103 13209
rect 35161 13209 35173 13212
rect 35207 13209 35219 13243
rect 46382 13240 46388 13252
rect 36386 13212 46388 13240
rect 35161 13203 35219 13209
rect 46382 13200 46388 13212
rect 46440 13200 46446 13252
rect 22186 13132 22192 13184
rect 22244 13172 22250 13184
rect 22465 13175 22523 13181
rect 22465 13172 22477 13175
rect 22244 13144 22477 13172
rect 22244 13132 22250 13144
rect 22465 13141 22477 13144
rect 22511 13141 22523 13175
rect 22465 13135 22523 13141
rect 1104 13082 48852 13104
rect 1104 13030 12898 13082
rect 12950 13030 12962 13082
rect 13014 13030 13026 13082
rect 13078 13030 13090 13082
rect 13142 13030 13154 13082
rect 13206 13030 24846 13082
rect 24898 13030 24910 13082
rect 24962 13030 24974 13082
rect 25026 13030 25038 13082
rect 25090 13030 25102 13082
rect 25154 13030 36794 13082
rect 36846 13030 36858 13082
rect 36910 13030 36922 13082
rect 36974 13030 36986 13082
rect 37038 13030 37050 13082
rect 37102 13030 48852 13082
rect 1104 13008 48852 13030
rect 29089 12971 29147 12977
rect 29089 12937 29101 12971
rect 29135 12968 29147 12971
rect 29178 12968 29184 12980
rect 29135 12940 29184 12968
rect 29135 12937 29147 12940
rect 29089 12931 29147 12937
rect 29178 12928 29184 12940
rect 29236 12928 29242 12980
rect 45094 12968 45100 12980
rect 45055 12940 45100 12968
rect 45094 12928 45100 12940
rect 45152 12928 45158 12980
rect 46382 12968 46388 12980
rect 46343 12940 46388 12968
rect 46382 12928 46388 12940
rect 46440 12928 46446 12980
rect 47670 12968 47676 12980
rect 47631 12940 47676 12968
rect 47670 12928 47676 12940
rect 47728 12928 47734 12980
rect 30377 12903 30435 12909
rect 30377 12869 30389 12903
rect 30423 12900 30435 12903
rect 33318 12900 33324 12912
rect 30423 12872 33324 12900
rect 30423 12869 30435 12872
rect 30377 12863 30435 12869
rect 33318 12860 33324 12872
rect 33376 12900 33382 12912
rect 33781 12903 33839 12909
rect 33781 12900 33793 12903
rect 33376 12872 33793 12900
rect 33376 12860 33382 12872
rect 33781 12869 33793 12872
rect 33827 12869 33839 12903
rect 33781 12863 33839 12869
rect 41049 12835 41107 12841
rect 41049 12801 41061 12835
rect 41095 12832 41107 12835
rect 45189 12835 45247 12841
rect 45189 12832 45201 12835
rect 41095 12804 45201 12832
rect 41095 12801 41107 12804
rect 41049 12795 41107 12801
rect 45189 12801 45201 12804
rect 45235 12832 45247 12835
rect 45833 12835 45891 12841
rect 45833 12832 45845 12835
rect 45235 12804 45845 12832
rect 45235 12801 45247 12804
rect 45189 12795 45247 12801
rect 45833 12801 45845 12804
rect 45879 12832 45891 12835
rect 46106 12832 46112 12844
rect 45879 12804 46112 12832
rect 45879 12801 45891 12804
rect 45833 12795 45891 12801
rect 46106 12792 46112 12804
rect 46164 12832 46170 12844
rect 46477 12835 46535 12841
rect 46477 12832 46489 12835
rect 46164 12804 46489 12832
rect 46164 12792 46170 12804
rect 46477 12801 46489 12804
rect 46523 12832 46535 12835
rect 47581 12835 47639 12841
rect 47581 12832 47593 12835
rect 46523 12804 47593 12832
rect 46523 12801 46535 12804
rect 46477 12795 46535 12801
rect 47581 12801 47593 12804
rect 47627 12801 47639 12835
rect 47581 12795 47639 12801
rect 30282 12724 30288 12776
rect 30340 12764 30346 12776
rect 45741 12767 45799 12773
rect 45741 12764 45753 12767
rect 30340 12736 45753 12764
rect 30340 12724 30346 12736
rect 45741 12733 45753 12736
rect 45787 12733 45799 12767
rect 45741 12727 45799 12733
rect 26050 12656 26056 12708
rect 26108 12696 26114 12708
rect 40957 12699 41015 12705
rect 40957 12696 40969 12699
rect 26108 12668 40969 12696
rect 26108 12656 26114 12668
rect 40957 12665 40969 12668
rect 41003 12665 41015 12699
rect 40957 12659 41015 12665
rect 1394 12628 1400 12640
rect 1355 12600 1400 12628
rect 1394 12588 1400 12600
rect 1452 12588 1458 12640
rect 34882 12588 34888 12640
rect 34940 12628 34946 12640
rect 35253 12631 35311 12637
rect 35253 12628 35265 12631
rect 34940 12600 35265 12628
rect 34940 12588 34946 12600
rect 35253 12597 35265 12600
rect 35299 12628 35311 12631
rect 39850 12628 39856 12640
rect 35299 12600 39856 12628
rect 35299 12597 35311 12600
rect 35253 12591 35311 12597
rect 39850 12588 39856 12600
rect 39908 12588 39914 12640
rect 1104 12538 48852 12560
rect 1104 12486 6924 12538
rect 6976 12486 6988 12538
rect 7040 12486 7052 12538
rect 7104 12486 7116 12538
rect 7168 12486 7180 12538
rect 7232 12486 18872 12538
rect 18924 12486 18936 12538
rect 18988 12486 19000 12538
rect 19052 12486 19064 12538
rect 19116 12486 19128 12538
rect 19180 12486 30820 12538
rect 30872 12486 30884 12538
rect 30936 12486 30948 12538
rect 31000 12486 31012 12538
rect 31064 12486 31076 12538
rect 31128 12486 42768 12538
rect 42820 12486 42832 12538
rect 42884 12486 42896 12538
rect 42948 12486 42960 12538
rect 43012 12486 43024 12538
rect 43076 12486 48852 12538
rect 1104 12464 48852 12486
rect 48133 12223 48191 12229
rect 48133 12189 48145 12223
rect 48179 12220 48191 12223
rect 48222 12220 48228 12232
rect 48179 12192 48228 12220
rect 48179 12189 48191 12192
rect 48133 12183 48191 12189
rect 48222 12180 48228 12192
rect 48280 12180 48286 12232
rect 1104 11994 48852 12016
rect 1104 11942 12898 11994
rect 12950 11942 12962 11994
rect 13014 11942 13026 11994
rect 13078 11942 13090 11994
rect 13142 11942 13154 11994
rect 13206 11942 24846 11994
rect 24898 11942 24910 11994
rect 24962 11942 24974 11994
rect 25026 11942 25038 11994
rect 25090 11942 25102 11994
rect 25154 11942 36794 11994
rect 36846 11942 36858 11994
rect 36910 11942 36922 11994
rect 36974 11942 36986 11994
rect 37038 11942 37050 11994
rect 37102 11942 48852 11994
rect 1104 11920 48852 11942
rect 1394 11676 1400 11688
rect 1355 11648 1400 11676
rect 1394 11636 1400 11648
rect 1452 11636 1458 11688
rect 48130 11540 48136 11552
rect 48091 11512 48136 11540
rect 48130 11500 48136 11512
rect 48188 11500 48194 11552
rect 1104 11450 48852 11472
rect 1104 11398 6924 11450
rect 6976 11398 6988 11450
rect 7040 11398 7052 11450
rect 7104 11398 7116 11450
rect 7168 11398 7180 11450
rect 7232 11398 18872 11450
rect 18924 11398 18936 11450
rect 18988 11398 19000 11450
rect 19052 11398 19064 11450
rect 19116 11398 19128 11450
rect 19180 11398 30820 11450
rect 30872 11398 30884 11450
rect 30936 11398 30948 11450
rect 31000 11398 31012 11450
rect 31064 11398 31076 11450
rect 31128 11398 42768 11450
rect 42820 11398 42832 11450
rect 42884 11398 42896 11450
rect 42948 11398 42960 11450
rect 43012 11398 43024 11450
rect 43076 11398 48852 11450
rect 1104 11376 48852 11398
rect 47394 11336 47400 11348
rect 47355 11308 47400 11336
rect 47394 11296 47400 11308
rect 47452 11296 47458 11348
rect 46934 11200 46940 11212
rect 46895 11172 46940 11200
rect 46934 11160 46940 11172
rect 46992 11160 46998 11212
rect 47029 11203 47087 11209
rect 47029 11169 47041 11203
rect 47075 11200 47087 11203
rect 47762 11200 47768 11212
rect 47075 11172 47768 11200
rect 47075 11169 47087 11172
rect 47029 11163 47087 11169
rect 47762 11160 47768 11172
rect 47820 11160 47826 11212
rect 47210 11132 47216 11144
rect 47171 11104 47216 11132
rect 47210 11092 47216 11104
rect 47268 11092 47274 11144
rect 1394 11064 1400 11076
rect 1355 11036 1400 11064
rect 1394 11024 1400 11036
rect 1452 11024 1458 11076
rect 1104 10906 48852 10928
rect 1104 10854 12898 10906
rect 12950 10854 12962 10906
rect 13014 10854 13026 10906
rect 13078 10854 13090 10906
rect 13142 10854 13154 10906
rect 13206 10854 24846 10906
rect 24898 10854 24910 10906
rect 24962 10854 24974 10906
rect 25026 10854 25038 10906
rect 25090 10854 25102 10906
rect 25154 10854 36794 10906
rect 36846 10854 36858 10906
rect 36910 10854 36922 10906
rect 36974 10854 36986 10906
rect 37038 10854 37050 10906
rect 37102 10854 48852 10906
rect 1104 10832 48852 10854
rect 47210 10752 47216 10804
rect 47268 10792 47274 10804
rect 47581 10795 47639 10801
rect 47581 10792 47593 10795
rect 47268 10764 47593 10792
rect 47268 10752 47274 10764
rect 47581 10761 47593 10764
rect 47627 10761 47639 10795
rect 47581 10755 47639 10761
rect 47578 10656 47584 10668
rect 47539 10628 47584 10656
rect 47578 10616 47584 10628
rect 47636 10616 47642 10668
rect 47762 10656 47768 10668
rect 47723 10628 47768 10656
rect 47762 10616 47768 10628
rect 47820 10616 47826 10668
rect 1104 10362 48852 10384
rect 1104 10310 6924 10362
rect 6976 10310 6988 10362
rect 7040 10310 7052 10362
rect 7104 10310 7116 10362
rect 7168 10310 7180 10362
rect 7232 10310 18872 10362
rect 18924 10310 18936 10362
rect 18988 10310 19000 10362
rect 19052 10310 19064 10362
rect 19116 10310 19128 10362
rect 19180 10310 30820 10362
rect 30872 10310 30884 10362
rect 30936 10310 30948 10362
rect 31000 10310 31012 10362
rect 31064 10310 31076 10362
rect 31128 10310 42768 10362
rect 42820 10310 42832 10362
rect 42884 10310 42896 10362
rect 42948 10310 42960 10362
rect 43012 10310 43024 10362
rect 43076 10310 48852 10362
rect 1104 10288 48852 10310
rect 48130 10044 48136 10056
rect 48091 10016 48136 10044
rect 48130 10004 48136 10016
rect 48188 10004 48194 10056
rect 1104 9818 48852 9840
rect 1104 9766 12898 9818
rect 12950 9766 12962 9818
rect 13014 9766 13026 9818
rect 13078 9766 13090 9818
rect 13142 9766 13154 9818
rect 13206 9766 24846 9818
rect 24898 9766 24910 9818
rect 24962 9766 24974 9818
rect 25026 9766 25038 9818
rect 25090 9766 25102 9818
rect 25154 9766 36794 9818
rect 36846 9766 36858 9818
rect 36910 9766 36922 9818
rect 36974 9766 36986 9818
rect 37038 9766 37050 9818
rect 37102 9766 48852 9818
rect 1104 9744 48852 9766
rect 45738 9528 45744 9580
rect 45796 9568 45802 9580
rect 46293 9571 46351 9577
rect 46293 9568 46305 9571
rect 45796 9540 46305 9568
rect 45796 9528 45802 9540
rect 46293 9537 46305 9540
rect 46339 9568 46351 9571
rect 47578 9568 47584 9580
rect 46339 9540 47584 9568
rect 46339 9537 46351 9540
rect 46293 9531 46351 9537
rect 47578 9528 47584 9540
rect 47636 9528 47642 9580
rect 46106 9432 46112 9444
rect 46067 9404 46112 9432
rect 46106 9392 46112 9404
rect 46164 9392 46170 9444
rect 1104 9274 48852 9296
rect 1104 9222 6924 9274
rect 6976 9222 6988 9274
rect 7040 9222 7052 9274
rect 7104 9222 7116 9274
rect 7168 9222 7180 9274
rect 7232 9222 18872 9274
rect 18924 9222 18936 9274
rect 18988 9222 19000 9274
rect 19052 9222 19064 9274
rect 19116 9222 19128 9274
rect 19180 9222 30820 9274
rect 30872 9222 30884 9274
rect 30936 9222 30948 9274
rect 31000 9222 31012 9274
rect 31064 9222 31076 9274
rect 31128 9222 42768 9274
rect 42820 9222 42832 9274
rect 42884 9222 42896 9274
rect 42948 9222 42960 9274
rect 43012 9222 43024 9274
rect 43076 9222 48852 9274
rect 1104 9200 48852 9222
rect 1394 8956 1400 8968
rect 1355 8928 1400 8956
rect 1394 8916 1400 8928
rect 1452 8916 1458 8968
rect 48130 8956 48136 8968
rect 48091 8928 48136 8956
rect 48130 8916 48136 8928
rect 48188 8916 48194 8968
rect 1104 8730 48852 8752
rect 1104 8678 12898 8730
rect 12950 8678 12962 8730
rect 13014 8678 13026 8730
rect 13078 8678 13090 8730
rect 13142 8678 13154 8730
rect 13206 8678 24846 8730
rect 24898 8678 24910 8730
rect 24962 8678 24974 8730
rect 25026 8678 25038 8730
rect 25090 8678 25102 8730
rect 25154 8678 36794 8730
rect 36846 8678 36858 8730
rect 36910 8678 36922 8730
rect 36974 8678 36986 8730
rect 37038 8678 37050 8730
rect 37102 8678 48852 8730
rect 1104 8656 48852 8678
rect 1394 8344 1400 8356
rect 1355 8316 1400 8344
rect 1394 8304 1400 8316
rect 1452 8304 1458 8356
rect 1104 8186 48852 8208
rect 1104 8134 6924 8186
rect 6976 8134 6988 8186
rect 7040 8134 7052 8186
rect 7104 8134 7116 8186
rect 7168 8134 7180 8186
rect 7232 8134 18872 8186
rect 18924 8134 18936 8186
rect 18988 8134 19000 8186
rect 19052 8134 19064 8186
rect 19116 8134 19128 8186
rect 19180 8134 30820 8186
rect 30872 8134 30884 8186
rect 30936 8134 30948 8186
rect 31000 8134 31012 8186
rect 31064 8134 31076 8186
rect 31128 8134 42768 8186
rect 42820 8134 42832 8186
rect 42884 8134 42896 8186
rect 42948 8134 42960 8186
rect 43012 8134 43024 8186
rect 43076 8134 48852 8186
rect 1104 8112 48852 8134
rect 47946 8072 47952 8084
rect 47907 8044 47952 8072
rect 47946 8032 47952 8044
rect 48004 8032 48010 8084
rect 48130 7868 48136 7880
rect 48091 7840 48136 7868
rect 48130 7828 48136 7840
rect 48188 7828 48194 7880
rect 1394 7732 1400 7744
rect 1355 7704 1400 7732
rect 1394 7692 1400 7704
rect 1452 7692 1458 7744
rect 1104 7642 48852 7664
rect 1104 7590 12898 7642
rect 12950 7590 12962 7642
rect 13014 7590 13026 7642
rect 13078 7590 13090 7642
rect 13142 7590 13154 7642
rect 13206 7590 24846 7642
rect 24898 7590 24910 7642
rect 24962 7590 24974 7642
rect 25026 7590 25038 7642
rect 25090 7590 25102 7642
rect 25154 7590 36794 7642
rect 36846 7590 36858 7642
rect 36910 7590 36922 7642
rect 36974 7590 36986 7642
rect 37038 7590 37050 7642
rect 37102 7590 48852 7642
rect 1104 7568 48852 7590
rect 1394 7324 1400 7336
rect 1355 7296 1400 7324
rect 1394 7284 1400 7296
rect 1452 7284 1458 7336
rect 48133 7327 48191 7333
rect 48133 7293 48145 7327
rect 48179 7324 48191 7327
rect 48222 7324 48228 7336
rect 48179 7296 48228 7324
rect 48179 7293 48191 7296
rect 48133 7287 48191 7293
rect 48222 7284 48228 7296
rect 48280 7284 48286 7336
rect 1104 7098 48852 7120
rect 1104 7046 6924 7098
rect 6976 7046 6988 7098
rect 7040 7046 7052 7098
rect 7104 7046 7116 7098
rect 7168 7046 7180 7098
rect 7232 7046 18872 7098
rect 18924 7046 18936 7098
rect 18988 7046 19000 7098
rect 19052 7046 19064 7098
rect 19116 7046 19128 7098
rect 19180 7046 30820 7098
rect 30872 7046 30884 7098
rect 30936 7046 30948 7098
rect 31000 7046 31012 7098
rect 31064 7046 31076 7098
rect 31128 7046 42768 7098
rect 42820 7046 42832 7098
rect 42884 7046 42896 7098
rect 42948 7046 42960 7098
rect 43012 7046 43024 7098
rect 43076 7046 48852 7098
rect 1104 7024 48852 7046
rect 1104 6554 48852 6576
rect 1104 6502 12898 6554
rect 12950 6502 12962 6554
rect 13014 6502 13026 6554
rect 13078 6502 13090 6554
rect 13142 6502 13154 6554
rect 13206 6502 24846 6554
rect 24898 6502 24910 6554
rect 24962 6502 24974 6554
rect 25026 6502 25038 6554
rect 25090 6502 25102 6554
rect 25154 6502 36794 6554
rect 36846 6502 36858 6554
rect 36910 6502 36922 6554
rect 36974 6502 36986 6554
rect 37038 6502 37050 6554
rect 37102 6502 48852 6554
rect 1104 6480 48852 6502
rect 1394 6236 1400 6248
rect 1355 6208 1400 6236
rect 1394 6196 1400 6208
rect 1452 6196 1458 6248
rect 48130 6100 48136 6112
rect 48091 6072 48136 6100
rect 48130 6060 48136 6072
rect 48188 6060 48194 6112
rect 1104 6010 48852 6032
rect 1104 5958 6924 6010
rect 6976 5958 6988 6010
rect 7040 5958 7052 6010
rect 7104 5958 7116 6010
rect 7168 5958 7180 6010
rect 7232 5958 18872 6010
rect 18924 5958 18936 6010
rect 18988 5958 19000 6010
rect 19052 5958 19064 6010
rect 19116 5958 19128 6010
rect 19180 5958 30820 6010
rect 30872 5958 30884 6010
rect 30936 5958 30948 6010
rect 31000 5958 31012 6010
rect 31064 5958 31076 6010
rect 31128 5958 42768 6010
rect 42820 5958 42832 6010
rect 42884 5958 42896 6010
rect 42948 5958 42960 6010
rect 43012 5958 43024 6010
rect 43076 5958 48852 6010
rect 1104 5936 48852 5958
rect 1394 5692 1400 5704
rect 1355 5664 1400 5692
rect 1394 5652 1400 5664
rect 1452 5652 1458 5704
rect 1104 5466 48852 5488
rect 1104 5414 12898 5466
rect 12950 5414 12962 5466
rect 13014 5414 13026 5466
rect 13078 5414 13090 5466
rect 13142 5414 13154 5466
rect 13206 5414 24846 5466
rect 24898 5414 24910 5466
rect 24962 5414 24974 5466
rect 25026 5414 25038 5466
rect 25090 5414 25102 5466
rect 25154 5414 36794 5466
rect 36846 5414 36858 5466
rect 36910 5414 36922 5466
rect 36974 5414 36986 5466
rect 37038 5414 37050 5466
rect 37102 5414 48852 5466
rect 1104 5392 48852 5414
rect 1394 5012 1400 5024
rect 1355 4984 1400 5012
rect 1394 4972 1400 4984
rect 1452 4972 1458 5024
rect 48133 5015 48191 5021
rect 48133 4981 48145 5015
rect 48179 5012 48191 5015
rect 48222 5012 48228 5024
rect 48179 4984 48228 5012
rect 48179 4981 48191 4984
rect 48133 4975 48191 4981
rect 48222 4972 48228 4984
rect 48280 4972 48286 5024
rect 1104 4922 48852 4944
rect 1104 4870 6924 4922
rect 6976 4870 6988 4922
rect 7040 4870 7052 4922
rect 7104 4870 7116 4922
rect 7168 4870 7180 4922
rect 7232 4870 18872 4922
rect 18924 4870 18936 4922
rect 18988 4870 19000 4922
rect 19052 4870 19064 4922
rect 19116 4870 19128 4922
rect 19180 4870 30820 4922
rect 30872 4870 30884 4922
rect 30936 4870 30948 4922
rect 31000 4870 31012 4922
rect 31064 4870 31076 4922
rect 31128 4870 42768 4922
rect 42820 4870 42832 4922
rect 42884 4870 42896 4922
rect 42948 4870 42960 4922
rect 43012 4870 43024 4922
rect 43076 4870 48852 4922
rect 1104 4848 48852 4870
rect 48130 4604 48136 4616
rect 48091 4576 48136 4604
rect 48130 4564 48136 4576
rect 48188 4564 48194 4616
rect 1104 4378 48852 4400
rect 1104 4326 12898 4378
rect 12950 4326 12962 4378
rect 13014 4326 13026 4378
rect 13078 4326 13090 4378
rect 13142 4326 13154 4378
rect 13206 4326 24846 4378
rect 24898 4326 24910 4378
rect 24962 4326 24974 4378
rect 25026 4326 25038 4378
rect 25090 4326 25102 4378
rect 25154 4326 36794 4378
rect 36846 4326 36858 4378
rect 36910 4326 36922 4378
rect 36974 4326 36986 4378
rect 37038 4326 37050 4378
rect 37102 4326 48852 4378
rect 1104 4304 48852 4326
rect 1397 3927 1455 3933
rect 1397 3893 1409 3927
rect 1443 3924 1455 3927
rect 2866 3924 2872 3936
rect 1443 3896 2872 3924
rect 1443 3893 1455 3896
rect 1397 3887 1455 3893
rect 2866 3884 2872 3896
rect 2924 3884 2930 3936
rect 47029 3927 47087 3933
rect 47029 3893 47041 3927
rect 47075 3924 47087 3927
rect 47762 3924 47768 3936
rect 47075 3896 47768 3924
rect 47075 3893 47087 3896
rect 47029 3887 47087 3893
rect 47762 3884 47768 3896
rect 47820 3884 47826 3936
rect 48133 3927 48191 3933
rect 48133 3893 48145 3927
rect 48179 3924 48191 3927
rect 48958 3924 48964 3936
rect 48179 3896 48964 3924
rect 48179 3893 48191 3896
rect 48133 3887 48191 3893
rect 48958 3884 48964 3896
rect 49016 3884 49022 3936
rect 1104 3834 48852 3856
rect 1104 3782 6924 3834
rect 6976 3782 6988 3834
rect 7040 3782 7052 3834
rect 7104 3782 7116 3834
rect 7168 3782 7180 3834
rect 7232 3782 18872 3834
rect 18924 3782 18936 3834
rect 18988 3782 19000 3834
rect 19052 3782 19064 3834
rect 19116 3782 19128 3834
rect 19180 3782 30820 3834
rect 30872 3782 30884 3834
rect 30936 3782 30948 3834
rect 31000 3782 31012 3834
rect 31064 3782 31076 3834
rect 31128 3782 42768 3834
rect 42820 3782 42832 3834
rect 42884 3782 42896 3834
rect 42948 3782 42960 3834
rect 43012 3782 43024 3834
rect 43076 3782 48852 3834
rect 1104 3760 48852 3782
rect 2041 3587 2099 3593
rect 2041 3553 2053 3587
rect 2087 3584 2099 3587
rect 2774 3584 2780 3596
rect 2087 3556 2780 3584
rect 2087 3553 2099 3556
rect 2041 3547 2099 3553
rect 2774 3544 2780 3556
rect 2832 3544 2838 3596
rect 1394 3516 1400 3528
rect 1355 3488 1400 3516
rect 1394 3476 1400 3488
rect 1452 3476 1458 3528
rect 2685 3519 2743 3525
rect 2685 3485 2697 3519
rect 2731 3516 2743 3519
rect 2958 3516 2964 3528
rect 2731 3488 2964 3516
rect 2731 3485 2743 3488
rect 2685 3479 2743 3485
rect 2958 3476 2964 3488
rect 3016 3476 3022 3528
rect 46658 3476 46664 3528
rect 46716 3516 46722 3528
rect 46845 3519 46903 3525
rect 46845 3516 46857 3519
rect 46716 3488 46857 3516
rect 46716 3476 46722 3488
rect 46845 3485 46857 3488
rect 46891 3485 46903 3519
rect 48130 3516 48136 3528
rect 48091 3488 48136 3516
rect 46845 3479 46903 3485
rect 48130 3476 48136 3488
rect 48188 3476 48194 3528
rect 47489 3383 47547 3389
rect 47489 3349 47501 3383
rect 47535 3380 47547 3383
rect 49602 3380 49608 3392
rect 47535 3352 49608 3380
rect 47535 3349 47547 3352
rect 47489 3343 47547 3349
rect 49602 3340 49608 3352
rect 49660 3340 49666 3392
rect 1104 3290 48852 3312
rect 1104 3238 12898 3290
rect 12950 3238 12962 3290
rect 13014 3238 13026 3290
rect 13078 3238 13090 3290
rect 13142 3238 13154 3290
rect 13206 3238 24846 3290
rect 24898 3238 24910 3290
rect 24962 3238 24974 3290
rect 25026 3238 25038 3290
rect 25090 3238 25102 3290
rect 25154 3238 36794 3290
rect 36846 3238 36858 3290
rect 36910 3238 36922 3290
rect 36974 3238 36986 3290
rect 37038 3238 37050 3290
rect 37102 3238 48852 3290
rect 1104 3216 48852 3238
rect 45738 3176 45744 3188
rect 45699 3148 45744 3176
rect 45738 3136 45744 3148
rect 45796 3136 45802 3188
rect 45554 3040 45560 3052
rect 45515 3012 45560 3040
rect 45554 3000 45560 3012
rect 45612 3000 45618 3052
rect 2685 2975 2743 2981
rect 2685 2941 2697 2975
rect 2731 2972 2743 2975
rect 3050 2972 3056 2984
rect 2731 2944 3056 2972
rect 2731 2941 2743 2944
rect 2685 2935 2743 2941
rect 3050 2932 3056 2944
rect 3108 2932 3114 2984
rect 3878 2932 3884 2984
rect 3936 2972 3942 2984
rect 3973 2975 4031 2981
rect 3973 2972 3985 2975
rect 3936 2944 3985 2972
rect 3936 2932 3942 2944
rect 3973 2941 3985 2944
rect 4019 2941 4031 2975
rect 3973 2935 4031 2941
rect 30742 2932 30748 2984
rect 30800 2972 30806 2984
rect 31021 2975 31079 2981
rect 31021 2972 31033 2975
rect 30800 2944 31033 2972
rect 30800 2932 30806 2944
rect 31021 2941 31033 2944
rect 31067 2941 31079 2975
rect 31021 2935 31079 2941
rect 36078 2932 36084 2984
rect 36136 2972 36142 2984
rect 36173 2975 36231 2981
rect 36173 2972 36185 2975
rect 36136 2944 36185 2972
rect 36136 2932 36142 2944
rect 36173 2941 36185 2944
rect 36219 2941 36231 2975
rect 36173 2935 36231 2941
rect 46842 2932 46848 2984
rect 46900 2972 46906 2984
rect 47029 2975 47087 2981
rect 47029 2972 47041 2975
rect 46900 2944 47041 2972
rect 46900 2932 46906 2944
rect 47029 2941 47041 2944
rect 47075 2941 47087 2975
rect 47029 2935 47087 2941
rect 47670 2932 47676 2984
rect 47728 2972 47734 2984
rect 47765 2975 47823 2981
rect 47765 2972 47777 2975
rect 47728 2944 47777 2972
rect 47728 2932 47734 2944
rect 47765 2941 47777 2944
rect 47811 2941 47823 2975
rect 47765 2935 47823 2941
rect 14 2864 20 2916
rect 72 2904 78 2916
rect 2041 2907 2099 2913
rect 2041 2904 2053 2907
rect 72 2876 2053 2904
rect 72 2864 78 2876
rect 2041 2873 2053 2876
rect 2087 2873 2099 2907
rect 2041 2867 2099 2873
rect 658 2796 664 2848
rect 716 2836 722 2848
rect 1397 2839 1455 2845
rect 1397 2836 1409 2839
rect 716 2808 1409 2836
rect 716 2796 722 2808
rect 1397 2805 1409 2808
rect 1443 2805 1455 2839
rect 1397 2799 1455 2805
rect 9030 2796 9036 2848
rect 9088 2836 9094 2848
rect 9125 2839 9183 2845
rect 9125 2836 9137 2839
rect 9088 2808 9137 2836
rect 9088 2796 9094 2808
rect 9125 2805 9137 2808
rect 9171 2805 9183 2839
rect 9125 2799 9183 2805
rect 16758 2796 16764 2848
rect 16816 2836 16822 2848
rect 16853 2839 16911 2845
rect 16853 2836 16865 2839
rect 16816 2808 16865 2836
rect 16816 2796 16822 2808
rect 16853 2805 16865 2808
rect 16899 2805 16911 2839
rect 16853 2799 16911 2805
rect 19334 2796 19340 2848
rect 19392 2836 19398 2848
rect 19429 2839 19487 2845
rect 19429 2836 19441 2839
rect 19392 2808 19441 2836
rect 19392 2796 19398 2808
rect 19429 2805 19441 2808
rect 19475 2805 19487 2839
rect 19429 2799 19487 2805
rect 23198 2796 23204 2848
rect 23256 2836 23262 2848
rect 23293 2839 23351 2845
rect 23293 2836 23305 2839
rect 23256 2808 23305 2836
rect 23256 2796 23262 2808
rect 23293 2805 23305 2808
rect 23339 2805 23351 2839
rect 23293 2799 23351 2805
rect 28350 2796 28356 2848
rect 28408 2836 28414 2848
rect 28445 2839 28503 2845
rect 28445 2836 28457 2839
rect 28408 2808 28457 2836
rect 28408 2796 28414 2808
rect 28445 2805 28457 2808
rect 28491 2805 28503 2839
rect 28445 2799 28503 2805
rect 43806 2796 43812 2848
rect 43864 2836 43870 2848
rect 43901 2839 43959 2845
rect 43901 2836 43913 2839
rect 43864 2808 43913 2836
rect 43864 2796 43870 2808
rect 43901 2805 43913 2808
rect 43947 2805 43959 2839
rect 43901 2799 43959 2805
rect 46385 2839 46443 2845
rect 46385 2805 46397 2839
rect 46431 2836 46443 2839
rect 46750 2836 46756 2848
rect 46431 2808 46756 2836
rect 46431 2805 46443 2808
rect 46385 2799 46443 2805
rect 46750 2796 46756 2808
rect 46808 2796 46814 2848
rect 1104 2746 48852 2768
rect 1104 2694 6924 2746
rect 6976 2694 6988 2746
rect 7040 2694 7052 2746
rect 7104 2694 7116 2746
rect 7168 2694 7180 2746
rect 7232 2694 18872 2746
rect 18924 2694 18936 2746
rect 18988 2694 19000 2746
rect 19052 2694 19064 2746
rect 19116 2694 19128 2746
rect 19180 2694 30820 2746
rect 30872 2694 30884 2746
rect 30936 2694 30948 2746
rect 31000 2694 31012 2746
rect 31064 2694 31076 2746
rect 31128 2694 42768 2746
rect 42820 2694 42832 2746
rect 42884 2694 42896 2746
rect 42948 2694 42960 2746
rect 43012 2694 43024 2746
rect 43076 2694 48852 2746
rect 1104 2672 48852 2694
rect 1302 2388 1308 2440
rect 1360 2428 1366 2440
rect 1397 2431 1455 2437
rect 1397 2428 1409 2431
rect 1360 2400 1409 2428
rect 1360 2388 1366 2400
rect 1397 2397 1409 2400
rect 1443 2397 1455 2431
rect 2590 2428 2596 2440
rect 2551 2400 2596 2428
rect 1397 2391 1455 2397
rect 2590 2388 2596 2400
rect 2648 2388 2654 2440
rect 3234 2428 3240 2440
rect 3195 2400 3240 2428
rect 3234 2388 3240 2400
rect 3292 2388 3298 2440
rect 5166 2428 5172 2440
rect 5127 2400 5172 2428
rect 5166 2388 5172 2400
rect 5224 2388 5230 2440
rect 5810 2428 5816 2440
rect 5771 2400 5816 2428
rect 5810 2388 5816 2400
rect 5868 2388 5874 2440
rect 7098 2428 7104 2440
rect 7059 2400 7104 2428
rect 7098 2388 7104 2400
rect 7156 2388 7162 2440
rect 7742 2428 7748 2440
rect 7703 2400 7748 2428
rect 7742 2388 7748 2400
rect 7800 2388 7806 2440
rect 8386 2428 8392 2440
rect 8347 2400 8392 2428
rect 8386 2388 8392 2400
rect 8444 2388 8450 2440
rect 10318 2428 10324 2440
rect 10279 2400 10324 2428
rect 10318 2388 10324 2400
rect 10376 2388 10382 2440
rect 10962 2428 10968 2440
rect 10923 2400 10968 2428
rect 10962 2388 10968 2400
rect 11020 2388 11026 2440
rect 12802 2388 12808 2440
rect 12860 2428 12866 2440
rect 12989 2431 13047 2437
rect 12989 2428 13001 2431
rect 12860 2400 13001 2428
rect 12860 2388 12866 2400
rect 12989 2397 13001 2400
rect 13035 2397 13047 2431
rect 12989 2391 13047 2397
rect 13538 2388 13544 2440
rect 13596 2428 13602 2440
rect 14093 2431 14151 2437
rect 14093 2428 14105 2431
rect 13596 2400 14105 2428
rect 13596 2388 13602 2400
rect 14093 2397 14105 2400
rect 14139 2397 14151 2431
rect 14093 2391 14151 2397
rect 14826 2388 14832 2440
rect 14884 2428 14890 2440
rect 14921 2431 14979 2437
rect 14921 2428 14933 2431
rect 14884 2400 14933 2428
rect 14884 2388 14890 2400
rect 14921 2397 14933 2400
rect 14967 2397 14979 2431
rect 17402 2428 17408 2440
rect 17363 2400 17408 2428
rect 14921 2391 14979 2397
rect 17402 2388 17408 2400
rect 17460 2388 17466 2440
rect 18046 2428 18052 2440
rect 18007 2400 18052 2428
rect 18046 2388 18052 2400
rect 18104 2388 18110 2440
rect 18690 2428 18696 2440
rect 18651 2400 18696 2428
rect 18690 2388 18696 2400
rect 18748 2388 18754 2440
rect 19978 2428 19984 2440
rect 19939 2400 19984 2428
rect 19978 2388 19984 2400
rect 20036 2388 20042 2440
rect 20622 2428 20628 2440
rect 20583 2400 20628 2428
rect 20622 2388 20628 2400
rect 20680 2388 20686 2440
rect 22186 2428 22192 2440
rect 22147 2400 22192 2428
rect 22186 2388 22192 2400
rect 22244 2388 22250 2440
rect 22922 2428 22928 2440
rect 22883 2400 22928 2428
rect 22922 2388 22928 2400
rect 22980 2388 22986 2440
rect 23842 2428 23848 2440
rect 23803 2400 23848 2428
rect 23842 2388 23848 2400
rect 23900 2388 23906 2440
rect 24486 2388 24492 2440
rect 24544 2428 24550 2440
rect 24581 2431 24639 2437
rect 24581 2428 24593 2431
rect 24544 2400 24593 2428
rect 24544 2388 24550 2400
rect 24581 2397 24593 2400
rect 24627 2397 24639 2431
rect 25222 2428 25228 2440
rect 25183 2400 25228 2428
rect 24581 2391 24639 2397
rect 25222 2388 25228 2400
rect 25280 2388 25286 2440
rect 25774 2388 25780 2440
rect 25832 2428 25838 2440
rect 25869 2431 25927 2437
rect 25869 2428 25881 2431
rect 25832 2400 25881 2428
rect 25832 2388 25838 2400
rect 25869 2397 25881 2400
rect 25915 2397 25927 2431
rect 25869 2391 25927 2397
rect 26418 2388 26424 2440
rect 26476 2428 26482 2440
rect 26973 2431 27031 2437
rect 26973 2428 26985 2431
rect 26476 2400 26985 2428
rect 26476 2388 26482 2400
rect 26973 2397 26985 2400
rect 27019 2397 27031 2431
rect 26973 2391 27031 2397
rect 28994 2388 29000 2440
rect 29052 2428 29058 2440
rect 29549 2431 29607 2437
rect 29549 2428 29561 2431
rect 29052 2400 29561 2428
rect 29052 2388 29058 2400
rect 29549 2397 29561 2400
rect 29595 2397 29607 2431
rect 29549 2391 29607 2397
rect 29638 2388 29644 2440
rect 29696 2428 29702 2440
rect 30193 2431 30251 2437
rect 30193 2428 30205 2431
rect 29696 2400 30205 2428
rect 29696 2388 29702 2400
rect 30193 2397 30205 2400
rect 30239 2397 30251 2431
rect 30193 2391 30251 2397
rect 30282 2388 30288 2440
rect 30340 2428 30346 2440
rect 30837 2431 30895 2437
rect 30837 2428 30849 2431
rect 30340 2400 30849 2428
rect 30340 2388 30346 2400
rect 30837 2397 30849 2400
rect 30883 2397 30895 2431
rect 30837 2391 30895 2397
rect 33502 2388 33508 2440
rect 33560 2428 33566 2440
rect 33597 2431 33655 2437
rect 33597 2428 33609 2431
rect 33560 2400 33609 2428
rect 33560 2388 33566 2400
rect 33597 2397 33609 2400
rect 33643 2397 33655 2431
rect 33597 2391 33655 2397
rect 34146 2388 34152 2440
rect 34204 2428 34210 2440
rect 34701 2431 34759 2437
rect 34701 2428 34713 2431
rect 34204 2400 34713 2428
rect 34204 2388 34210 2400
rect 34701 2397 34713 2400
rect 34747 2397 34759 2431
rect 34701 2391 34759 2397
rect 34790 2388 34796 2440
rect 34848 2428 34854 2440
rect 35345 2431 35403 2437
rect 35345 2428 35357 2431
rect 34848 2400 35357 2428
rect 34848 2388 34854 2400
rect 35345 2397 35357 2400
rect 35391 2397 35403 2431
rect 35345 2391 35403 2397
rect 37366 2388 37372 2440
rect 37424 2428 37430 2440
rect 37461 2431 37519 2437
rect 37461 2428 37473 2431
rect 37424 2400 37473 2428
rect 37424 2388 37430 2400
rect 37461 2397 37473 2400
rect 37507 2397 37519 2431
rect 37461 2391 37519 2397
rect 38654 2388 38660 2440
rect 38712 2428 38718 2440
rect 38749 2431 38807 2437
rect 38749 2428 38761 2431
rect 38712 2400 38761 2428
rect 38712 2388 38718 2400
rect 38749 2397 38761 2400
rect 38795 2397 38807 2431
rect 38749 2391 38807 2397
rect 39298 2388 39304 2440
rect 39356 2428 39362 2440
rect 39853 2431 39911 2437
rect 39853 2428 39865 2431
rect 39356 2400 39865 2428
rect 39356 2388 39362 2400
rect 39853 2397 39865 2400
rect 39899 2397 39911 2431
rect 39853 2391 39911 2397
rect 40586 2388 40592 2440
rect 40644 2428 40650 2440
rect 40681 2431 40739 2437
rect 40681 2428 40693 2431
rect 40644 2400 40693 2428
rect 40644 2388 40650 2400
rect 40681 2397 40693 2400
rect 40727 2397 40739 2431
rect 40681 2391 40739 2397
rect 41230 2388 41236 2440
rect 41288 2428 41294 2440
rect 41325 2431 41383 2437
rect 41325 2428 41337 2431
rect 41288 2400 41337 2428
rect 41288 2388 41294 2400
rect 41325 2397 41337 2400
rect 41371 2397 41383 2431
rect 41325 2391 41383 2397
rect 42518 2388 42524 2440
rect 42576 2428 42582 2440
rect 43073 2431 43131 2437
rect 43073 2428 43085 2431
rect 42576 2400 43085 2428
rect 42576 2388 42582 2400
rect 43073 2397 43085 2400
rect 43119 2397 43131 2431
rect 43073 2391 43131 2397
rect 46382 2388 46388 2440
rect 46440 2428 46446 2440
rect 46477 2431 46535 2437
rect 46477 2428 46489 2431
rect 46440 2400 46489 2428
rect 46440 2388 46446 2400
rect 46477 2397 46489 2400
rect 46523 2397 46535 2431
rect 46477 2391 46535 2397
rect 47026 2388 47032 2440
rect 47084 2428 47090 2440
rect 47581 2431 47639 2437
rect 47581 2428 47593 2431
rect 47084 2400 47593 2428
rect 47084 2388 47090 2400
rect 47581 2397 47593 2400
rect 47627 2397 47639 2431
rect 47581 2391 47639 2397
rect 4522 2292 4528 2304
rect 4483 2264 4528 2292
rect 4522 2252 4528 2264
rect 4580 2252 4586 2304
rect 9674 2252 9680 2304
rect 9732 2292 9738 2304
rect 9732 2264 9777 2292
rect 9732 2252 9738 2264
rect 11606 2252 11612 2304
rect 11664 2292 11670 2304
rect 11701 2295 11759 2301
rect 11701 2292 11713 2295
rect 11664 2264 11713 2292
rect 11664 2252 11670 2264
rect 11701 2261 11713 2264
rect 11747 2261 11759 2295
rect 11701 2255 11759 2261
rect 12250 2252 12256 2304
rect 12308 2292 12314 2304
rect 12345 2295 12403 2301
rect 12345 2292 12357 2295
rect 12308 2264 12357 2292
rect 12308 2252 12314 2264
rect 12345 2261 12357 2264
rect 12391 2261 12403 2295
rect 16114 2292 16120 2304
rect 16075 2264 16120 2292
rect 12345 2255 12403 2261
rect 16114 2252 16120 2264
rect 16172 2252 16178 2304
rect 21266 2292 21272 2304
rect 21227 2264 21272 2292
rect 21266 2252 21272 2264
rect 21324 2252 21330 2304
rect 21910 2252 21916 2304
rect 21968 2292 21974 2304
rect 22005 2295 22063 2301
rect 22005 2292 22017 2295
rect 21968 2264 22017 2292
rect 21968 2252 21974 2264
rect 22005 2261 22017 2264
rect 22051 2261 22063 2295
rect 22005 2255 22063 2261
rect 22554 2252 22560 2304
rect 22612 2292 22618 2304
rect 22741 2295 22799 2301
rect 22741 2292 22753 2295
rect 22612 2264 22753 2292
rect 22612 2252 22618 2264
rect 22741 2261 22753 2264
rect 22787 2261 22799 2295
rect 22741 2255 22799 2261
rect 27062 2252 27068 2304
rect 27120 2292 27126 2304
rect 27617 2295 27675 2301
rect 27617 2292 27629 2295
rect 27120 2264 27629 2292
rect 27120 2252 27126 2264
rect 27617 2261 27629 2264
rect 27663 2261 27675 2295
rect 27617 2255 27675 2261
rect 27706 2252 27712 2304
rect 27764 2292 27770 2304
rect 28261 2295 28319 2301
rect 28261 2292 28273 2295
rect 27764 2264 28273 2292
rect 27764 2252 27770 2264
rect 28261 2261 28273 2264
rect 28307 2261 28319 2295
rect 28261 2255 28319 2261
rect 32214 2252 32220 2304
rect 32272 2292 32278 2304
rect 32309 2295 32367 2301
rect 32309 2292 32321 2295
rect 32272 2264 32321 2292
rect 32272 2252 32278 2264
rect 32309 2261 32321 2264
rect 32355 2261 32367 2295
rect 32309 2255 32367 2261
rect 32858 2252 32864 2304
rect 32916 2292 32922 2304
rect 32953 2295 33011 2301
rect 32953 2292 32965 2295
rect 32916 2264 32965 2292
rect 32916 2252 32922 2264
rect 32953 2261 32965 2264
rect 32999 2261 33011 2295
rect 32953 2255 33011 2261
rect 35434 2252 35440 2304
rect 35492 2292 35498 2304
rect 35989 2295 36047 2301
rect 35989 2292 36001 2295
rect 35492 2264 36001 2292
rect 35492 2252 35498 2264
rect 35989 2261 36001 2264
rect 36035 2261 36047 2295
rect 35989 2255 36047 2261
rect 41874 2252 41880 2304
rect 41932 2292 41938 2304
rect 42429 2295 42487 2301
rect 42429 2292 42441 2295
rect 41932 2264 42441 2292
rect 41932 2252 41938 2264
rect 42429 2261 42441 2264
rect 42475 2261 42487 2295
rect 42429 2255 42487 2261
rect 43162 2252 43168 2304
rect 43220 2292 43226 2304
rect 43717 2295 43775 2301
rect 43717 2292 43729 2295
rect 43220 2264 43729 2292
rect 43220 2252 43226 2264
rect 43717 2261 43729 2264
rect 43763 2261 43775 2295
rect 43717 2255 43775 2261
rect 44450 2252 44456 2304
rect 44508 2292 44514 2304
rect 45005 2295 45063 2301
rect 45005 2292 45017 2295
rect 44508 2264 45017 2292
rect 44508 2252 44514 2264
rect 45005 2261 45017 2264
rect 45051 2261 45063 2295
rect 45005 2255 45063 2261
rect 45094 2252 45100 2304
rect 45152 2292 45158 2304
rect 45649 2295 45707 2301
rect 45649 2292 45661 2295
rect 45152 2264 45661 2292
rect 45152 2252 45158 2264
rect 45649 2261 45661 2264
rect 45695 2261 45707 2295
rect 45649 2255 45707 2261
rect 1104 2202 48852 2224
rect 1104 2150 12898 2202
rect 12950 2150 12962 2202
rect 13014 2150 13026 2202
rect 13078 2150 13090 2202
rect 13142 2150 13154 2202
rect 13206 2150 24846 2202
rect 24898 2150 24910 2202
rect 24962 2150 24974 2202
rect 25026 2150 25038 2202
rect 25090 2150 25102 2202
rect 25154 2150 36794 2202
rect 36846 2150 36858 2202
rect 36910 2150 36922 2202
rect 36974 2150 36986 2202
rect 37038 2150 37050 2202
rect 37102 2150 48852 2202
rect 1104 2128 48852 2150
<< via1 >>
rect 6924 27718 6976 27770
rect 6988 27718 7040 27770
rect 7052 27718 7104 27770
rect 7116 27718 7168 27770
rect 7180 27718 7232 27770
rect 18872 27718 18924 27770
rect 18936 27718 18988 27770
rect 19000 27718 19052 27770
rect 19064 27718 19116 27770
rect 19128 27718 19180 27770
rect 30820 27718 30872 27770
rect 30884 27718 30936 27770
rect 30948 27718 31000 27770
rect 31012 27718 31064 27770
rect 31076 27718 31128 27770
rect 42768 27718 42820 27770
rect 42832 27718 42884 27770
rect 42896 27718 42948 27770
rect 42960 27718 43012 27770
rect 43024 27718 43076 27770
rect 2044 27591 2096 27600
rect 2044 27557 2053 27591
rect 2053 27557 2087 27591
rect 2087 27557 2096 27591
rect 2044 27548 2096 27557
rect 3976 27591 4028 27600
rect 3976 27557 3985 27591
rect 3985 27557 4019 27591
rect 4019 27557 4028 27591
rect 3976 27548 4028 27557
rect 5172 27591 5224 27600
rect 5172 27557 5181 27591
rect 5181 27557 5215 27591
rect 5215 27557 5224 27591
rect 5172 27548 5224 27557
rect 5816 27591 5868 27600
rect 5816 27557 5825 27591
rect 5825 27557 5859 27591
rect 5859 27557 5868 27591
rect 5816 27548 5868 27557
rect 7748 27591 7800 27600
rect 7748 27557 7757 27591
rect 7757 27557 7791 27591
rect 7791 27557 7800 27591
rect 7748 27548 7800 27557
rect 8392 27591 8444 27600
rect 8392 27557 8401 27591
rect 8401 27557 8435 27591
rect 8435 27557 8444 27591
rect 8392 27548 8444 27557
rect 10324 27591 10376 27600
rect 10324 27557 10333 27591
rect 10333 27557 10367 27591
rect 10367 27557 10376 27591
rect 10324 27548 10376 27557
rect 10968 27591 11020 27600
rect 10968 27557 10977 27591
rect 10977 27557 11011 27591
rect 11011 27557 11020 27591
rect 10968 27548 11020 27557
rect 13820 27548 13872 27600
rect 14924 27591 14976 27600
rect 14924 27557 14933 27591
rect 14933 27557 14967 27591
rect 14967 27557 14976 27591
rect 14924 27548 14976 27557
rect 15568 27591 15620 27600
rect 15568 27557 15577 27591
rect 15577 27557 15611 27591
rect 15611 27557 15620 27591
rect 15568 27548 15620 27557
rect 18052 27591 18104 27600
rect 18052 27557 18061 27591
rect 18061 27557 18095 27591
rect 18095 27557 18104 27591
rect 18052 27548 18104 27557
rect 18696 27591 18748 27600
rect 18696 27557 18705 27591
rect 18705 27557 18739 27591
rect 18739 27557 18748 27591
rect 18696 27548 18748 27557
rect 19984 27591 20036 27600
rect 19984 27557 19993 27591
rect 19993 27557 20027 27591
rect 20027 27557 20036 27591
rect 19984 27548 20036 27557
rect 20628 27591 20680 27600
rect 20628 27557 20637 27591
rect 20637 27557 20671 27591
rect 20671 27557 20680 27591
rect 20628 27548 20680 27557
rect 21272 27591 21324 27600
rect 21272 27557 21281 27591
rect 21281 27557 21315 27591
rect 21315 27557 21324 27591
rect 21272 27548 21324 27557
rect 23204 27591 23256 27600
rect 23204 27557 23213 27591
rect 23213 27557 23247 27591
rect 23247 27557 23256 27591
rect 23204 27548 23256 27557
rect 24584 27591 24636 27600
rect 24584 27557 24593 27591
rect 24593 27557 24627 27591
rect 24627 27557 24636 27591
rect 24584 27548 24636 27557
rect 25228 27591 25280 27600
rect 25228 27557 25237 27591
rect 25237 27557 25271 27591
rect 25271 27557 25280 27591
rect 25228 27548 25280 27557
rect 25872 27591 25924 27600
rect 25872 27557 25881 27591
rect 25881 27557 25915 27591
rect 25915 27557 25924 27591
rect 25872 27548 25924 27557
rect 26424 27548 26476 27600
rect 30380 27591 30432 27600
rect 30380 27557 30389 27591
rect 30389 27557 30423 27591
rect 30423 27557 30432 27591
rect 30380 27548 30432 27557
rect 31208 27548 31260 27600
rect 32312 27591 32364 27600
rect 32312 27557 32321 27591
rect 32321 27557 32355 27591
rect 32355 27557 32364 27591
rect 32312 27548 32364 27557
rect 33600 27591 33652 27600
rect 33600 27557 33609 27591
rect 33609 27557 33643 27591
rect 33643 27557 33652 27591
rect 33600 27548 33652 27557
rect 34520 27548 34572 27600
rect 37280 27591 37332 27600
rect 37280 27557 37289 27591
rect 37289 27557 37323 27591
rect 37323 27557 37332 27591
rect 37280 27548 37332 27557
rect 37372 27548 37424 27600
rect 38016 27548 38068 27600
rect 40040 27591 40092 27600
rect 40040 27557 40049 27591
rect 40049 27557 40083 27591
rect 40083 27557 40092 27591
rect 40040 27548 40092 27557
rect 41328 27591 41380 27600
rect 41328 27557 41337 27591
rect 41337 27557 41371 27591
rect 41371 27557 41380 27591
rect 41328 27548 41380 27557
rect 43168 27548 43220 27600
rect 45192 27591 45244 27600
rect 45192 27557 45201 27591
rect 45201 27557 45235 27591
rect 45235 27557 45244 27591
rect 45192 27548 45244 27557
rect 45836 27591 45888 27600
rect 45836 27557 45845 27591
rect 45845 27557 45879 27591
rect 45879 27557 45888 27591
rect 45836 27548 45888 27557
rect 46480 27591 46532 27600
rect 46480 27557 46489 27591
rect 46489 27557 46523 27591
rect 46523 27557 46532 27591
rect 46480 27548 46532 27557
rect 1308 27480 1360 27532
rect 7288 27480 7340 27532
rect 9680 27523 9732 27532
rect 9680 27489 9689 27523
rect 9689 27489 9723 27523
rect 9723 27489 9732 27523
rect 11704 27523 11756 27532
rect 9680 27480 9732 27489
rect 11704 27489 11713 27523
rect 11713 27489 11747 27523
rect 11747 27489 11756 27523
rect 11704 27480 11756 27489
rect 12348 27523 12400 27532
rect 12348 27489 12357 27523
rect 12357 27489 12391 27523
rect 12391 27489 12400 27523
rect 12348 27480 12400 27489
rect 12992 27523 13044 27532
rect 12992 27489 13001 27523
rect 13001 27489 13035 27523
rect 13035 27489 13044 27523
rect 12992 27480 13044 27489
rect 16580 27480 16632 27532
rect 22560 27523 22612 27532
rect 22560 27489 22569 27523
rect 22569 27489 22603 27523
rect 22603 27489 22612 27523
rect 22560 27480 22612 27489
rect 23848 27523 23900 27532
rect 23848 27489 23857 27523
rect 23857 27489 23891 27523
rect 23891 27489 23900 27523
rect 23848 27480 23900 27489
rect 27804 27523 27856 27532
rect 27804 27489 27813 27523
rect 27813 27489 27847 27523
rect 27847 27489 27856 27523
rect 27804 27480 27856 27489
rect 28448 27523 28500 27532
rect 28448 27489 28457 27523
rect 28457 27489 28491 27523
rect 28491 27489 28500 27523
rect 28448 27480 28500 27489
rect 29000 27480 29052 27532
rect 34796 27480 34848 27532
rect 35900 27480 35952 27532
rect 40684 27523 40736 27532
rect 40684 27489 40693 27523
rect 40693 27489 40727 27523
rect 40727 27489 40736 27523
rect 40684 27480 40736 27489
rect 42616 27523 42668 27532
rect 42616 27489 42625 27523
rect 42625 27489 42659 27523
rect 42659 27489 42668 27523
rect 42616 27480 42668 27489
rect 20 27412 72 27464
rect 22928 27344 22980 27396
rect 47400 27412 47452 27464
rect 48320 27276 48372 27328
rect 12898 27174 12950 27226
rect 12962 27174 13014 27226
rect 13026 27174 13078 27226
rect 13090 27174 13142 27226
rect 13154 27174 13206 27226
rect 24846 27174 24898 27226
rect 24910 27174 24962 27226
rect 24974 27174 25026 27226
rect 25038 27174 25090 27226
rect 25102 27174 25154 27226
rect 36794 27174 36846 27226
rect 36858 27174 36910 27226
rect 36922 27174 36974 27226
rect 36986 27174 37038 27226
rect 37050 27174 37102 27226
rect 664 27072 716 27124
rect 47032 27072 47084 27124
rect 2872 27004 2924 27056
rect 1400 26979 1452 26988
rect 1400 26945 1409 26979
rect 1409 26945 1443 26979
rect 1443 26945 1452 26979
rect 1400 26936 1452 26945
rect 6552 26979 6604 26988
rect 6552 26945 6561 26979
rect 6561 26945 6595 26979
rect 6595 26945 6604 26979
rect 6552 26936 6604 26945
rect 9128 26979 9180 26988
rect 9128 26945 9137 26979
rect 9137 26945 9171 26979
rect 9171 26945 9180 26979
rect 9128 26936 9180 26945
rect 19432 26979 19484 26988
rect 19432 26945 19441 26979
rect 19441 26945 19475 26979
rect 19475 26945 19484 26979
rect 19432 26936 19484 26945
rect 22008 26979 22060 26988
rect 22008 26945 22017 26979
rect 22017 26945 22051 26979
rect 22051 26945 22060 26979
rect 22008 26936 22060 26945
rect 36176 26979 36228 26988
rect 36176 26945 36185 26979
rect 36185 26945 36219 26979
rect 36219 26945 36228 26979
rect 36176 26936 36228 26945
rect 38752 26979 38804 26988
rect 38752 26945 38761 26979
rect 38761 26945 38795 26979
rect 38795 26945 38804 26979
rect 38752 26936 38804 26945
rect 41880 26936 41932 26988
rect 43904 26979 43956 26988
rect 43904 26945 43913 26979
rect 43913 26945 43947 26979
rect 43947 26945 43956 26979
rect 43904 26936 43956 26945
rect 45744 26979 45796 26988
rect 45744 26945 45753 26979
rect 45753 26945 45787 26979
rect 45787 26945 45796 26979
rect 45744 26936 45796 26945
rect 47676 26936 47728 26988
rect 48964 26868 49016 26920
rect 6924 26630 6976 26682
rect 6988 26630 7040 26682
rect 7052 26630 7104 26682
rect 7116 26630 7168 26682
rect 7180 26630 7232 26682
rect 18872 26630 18924 26682
rect 18936 26630 18988 26682
rect 19000 26630 19052 26682
rect 19064 26630 19116 26682
rect 19128 26630 19180 26682
rect 30820 26630 30872 26682
rect 30884 26630 30936 26682
rect 30948 26630 31000 26682
rect 31012 26630 31064 26682
rect 31076 26630 31128 26682
rect 42768 26630 42820 26682
rect 42832 26630 42884 26682
rect 42896 26630 42948 26682
rect 42960 26630 43012 26682
rect 43024 26630 43076 26682
rect 2780 26528 2832 26580
rect 47492 26571 47544 26580
rect 47492 26537 47501 26571
rect 47501 26537 47535 26571
rect 47535 26537 47544 26571
rect 47492 26528 47544 26537
rect 46848 26435 46900 26444
rect 46848 26401 46857 26435
rect 46857 26401 46891 26435
rect 46891 26401 46900 26435
rect 46848 26392 46900 26401
rect 1400 26367 1452 26376
rect 1400 26333 1409 26367
rect 1409 26333 1443 26367
rect 1443 26333 1452 26367
rect 1400 26324 1452 26333
rect 48228 26188 48280 26240
rect 12898 26086 12950 26138
rect 12962 26086 13014 26138
rect 13026 26086 13078 26138
rect 13090 26086 13142 26138
rect 13154 26086 13206 26138
rect 24846 26086 24898 26138
rect 24910 26086 24962 26138
rect 24974 26086 25026 26138
rect 25038 26086 25090 26138
rect 25102 26086 25154 26138
rect 36794 26086 36846 26138
rect 36858 26086 36910 26138
rect 36922 26086 36974 26138
rect 36986 26086 37038 26138
rect 37050 26086 37102 26138
rect 1492 25848 1544 25900
rect 48136 25891 48188 25900
rect 48136 25857 48145 25891
rect 48145 25857 48179 25891
rect 48179 25857 48188 25891
rect 48136 25848 48188 25857
rect 49608 25780 49660 25832
rect 6924 25542 6976 25594
rect 6988 25542 7040 25594
rect 7052 25542 7104 25594
rect 7116 25542 7168 25594
rect 7180 25542 7232 25594
rect 18872 25542 18924 25594
rect 18936 25542 18988 25594
rect 19000 25542 19052 25594
rect 19064 25542 19116 25594
rect 19128 25542 19180 25594
rect 30820 25542 30872 25594
rect 30884 25542 30936 25594
rect 30948 25542 31000 25594
rect 31012 25542 31064 25594
rect 31076 25542 31128 25594
rect 42768 25542 42820 25594
rect 42832 25542 42884 25594
rect 42896 25542 42948 25594
rect 42960 25542 43012 25594
rect 43024 25542 43076 25594
rect 1400 25279 1452 25288
rect 1400 25245 1409 25279
rect 1409 25245 1443 25279
rect 1443 25245 1452 25279
rect 1400 25236 1452 25245
rect 48136 25279 48188 25288
rect 48136 25245 48145 25279
rect 48145 25245 48179 25279
rect 48179 25245 48188 25279
rect 48136 25236 48188 25245
rect 12898 24998 12950 25050
rect 12962 24998 13014 25050
rect 13026 24998 13078 25050
rect 13090 24998 13142 25050
rect 13154 24998 13206 25050
rect 24846 24998 24898 25050
rect 24910 24998 24962 25050
rect 24974 24998 25026 25050
rect 25038 24998 25090 25050
rect 25102 24998 25154 25050
rect 36794 24998 36846 25050
rect 36858 24998 36910 25050
rect 36922 24998 36974 25050
rect 36986 24998 37038 25050
rect 37050 24998 37102 25050
rect 1400 24599 1452 24608
rect 1400 24565 1409 24599
rect 1409 24565 1443 24599
rect 1443 24565 1452 24599
rect 1400 24556 1452 24565
rect 48136 24599 48188 24608
rect 48136 24565 48145 24599
rect 48145 24565 48179 24599
rect 48179 24565 48188 24599
rect 48136 24556 48188 24565
rect 6924 24454 6976 24506
rect 6988 24454 7040 24506
rect 7052 24454 7104 24506
rect 7116 24454 7168 24506
rect 7180 24454 7232 24506
rect 18872 24454 18924 24506
rect 18936 24454 18988 24506
rect 19000 24454 19052 24506
rect 19064 24454 19116 24506
rect 19128 24454 19180 24506
rect 30820 24454 30872 24506
rect 30884 24454 30936 24506
rect 30948 24454 31000 24506
rect 31012 24454 31064 24506
rect 31076 24454 31128 24506
rect 42768 24454 42820 24506
rect 42832 24454 42884 24506
rect 42896 24454 42948 24506
rect 42960 24454 43012 24506
rect 43024 24454 43076 24506
rect 48228 24148 48280 24200
rect 1400 24055 1452 24064
rect 1400 24021 1409 24055
rect 1409 24021 1443 24055
rect 1443 24021 1452 24055
rect 1400 24012 1452 24021
rect 12898 23910 12950 23962
rect 12962 23910 13014 23962
rect 13026 23910 13078 23962
rect 13090 23910 13142 23962
rect 13154 23910 13206 23962
rect 24846 23910 24898 23962
rect 24910 23910 24962 23962
rect 24974 23910 25026 23962
rect 25038 23910 25090 23962
rect 25102 23910 25154 23962
rect 36794 23910 36846 23962
rect 36858 23910 36910 23962
rect 36922 23910 36974 23962
rect 36986 23910 37038 23962
rect 37050 23910 37102 23962
rect 1400 23511 1452 23520
rect 1400 23477 1409 23511
rect 1409 23477 1443 23511
rect 1443 23477 1452 23511
rect 1400 23468 1452 23477
rect 48136 23511 48188 23520
rect 48136 23477 48145 23511
rect 48145 23477 48179 23511
rect 48179 23477 48188 23511
rect 48136 23468 48188 23477
rect 6924 23366 6976 23418
rect 6988 23366 7040 23418
rect 7052 23366 7104 23418
rect 7116 23366 7168 23418
rect 7180 23366 7232 23418
rect 18872 23366 18924 23418
rect 18936 23366 18988 23418
rect 19000 23366 19052 23418
rect 19064 23366 19116 23418
rect 19128 23366 19180 23418
rect 30820 23366 30872 23418
rect 30884 23366 30936 23418
rect 30948 23366 31000 23418
rect 31012 23366 31064 23418
rect 31076 23366 31128 23418
rect 42768 23366 42820 23418
rect 42832 23366 42884 23418
rect 42896 23366 42948 23418
rect 42960 23366 43012 23418
rect 43024 23366 43076 23418
rect 12898 22822 12950 22874
rect 12962 22822 13014 22874
rect 13026 22822 13078 22874
rect 13090 22822 13142 22874
rect 13154 22822 13206 22874
rect 24846 22822 24898 22874
rect 24910 22822 24962 22874
rect 24974 22822 25026 22874
rect 25038 22822 25090 22874
rect 25102 22822 25154 22874
rect 36794 22822 36846 22874
rect 36858 22822 36910 22874
rect 36922 22822 36974 22874
rect 36986 22822 37038 22874
rect 37050 22822 37102 22874
rect 48136 22423 48188 22432
rect 48136 22389 48145 22423
rect 48145 22389 48179 22423
rect 48179 22389 48188 22423
rect 48136 22380 48188 22389
rect 6924 22278 6976 22330
rect 6988 22278 7040 22330
rect 7052 22278 7104 22330
rect 7116 22278 7168 22330
rect 7180 22278 7232 22330
rect 18872 22278 18924 22330
rect 18936 22278 18988 22330
rect 19000 22278 19052 22330
rect 19064 22278 19116 22330
rect 19128 22278 19180 22330
rect 30820 22278 30872 22330
rect 30884 22278 30936 22330
rect 30948 22278 31000 22330
rect 31012 22278 31064 22330
rect 31076 22278 31128 22330
rect 42768 22278 42820 22330
rect 42832 22278 42884 22330
rect 42896 22278 42948 22330
rect 42960 22278 43012 22330
rect 43024 22278 43076 22330
rect 1400 22015 1452 22024
rect 1400 21981 1409 22015
rect 1409 21981 1443 22015
rect 1443 21981 1452 22015
rect 1400 21972 1452 21981
rect 48136 22015 48188 22024
rect 48136 21981 48145 22015
rect 48145 21981 48179 22015
rect 48179 21981 48188 22015
rect 48136 21972 48188 21981
rect 12898 21734 12950 21786
rect 12962 21734 13014 21786
rect 13026 21734 13078 21786
rect 13090 21734 13142 21786
rect 13154 21734 13206 21786
rect 24846 21734 24898 21786
rect 24910 21734 24962 21786
rect 24974 21734 25026 21786
rect 25038 21734 25090 21786
rect 25102 21734 25154 21786
rect 36794 21734 36846 21786
rect 36858 21734 36910 21786
rect 36922 21734 36974 21786
rect 36986 21734 37038 21786
rect 37050 21734 37102 21786
rect 1400 21335 1452 21344
rect 1400 21301 1409 21335
rect 1409 21301 1443 21335
rect 1443 21301 1452 21335
rect 1400 21292 1452 21301
rect 6924 21190 6976 21242
rect 6988 21190 7040 21242
rect 7052 21190 7104 21242
rect 7116 21190 7168 21242
rect 7180 21190 7232 21242
rect 18872 21190 18924 21242
rect 18936 21190 18988 21242
rect 19000 21190 19052 21242
rect 19064 21190 19116 21242
rect 19128 21190 19180 21242
rect 30820 21190 30872 21242
rect 30884 21190 30936 21242
rect 30948 21190 31000 21242
rect 31012 21190 31064 21242
rect 31076 21190 31128 21242
rect 42768 21190 42820 21242
rect 42832 21190 42884 21242
rect 42896 21190 42948 21242
rect 42960 21190 43012 21242
rect 43024 21190 43076 21242
rect 1400 20927 1452 20936
rect 1400 20893 1409 20927
rect 1409 20893 1443 20927
rect 1443 20893 1452 20927
rect 1400 20884 1452 20893
rect 48228 20884 48280 20936
rect 12898 20646 12950 20698
rect 12962 20646 13014 20698
rect 13026 20646 13078 20698
rect 13090 20646 13142 20698
rect 13154 20646 13206 20698
rect 24846 20646 24898 20698
rect 24910 20646 24962 20698
rect 24974 20646 25026 20698
rect 25038 20646 25090 20698
rect 25102 20646 25154 20698
rect 36794 20646 36846 20698
rect 36858 20646 36910 20698
rect 36922 20646 36974 20698
rect 36986 20646 37038 20698
rect 37050 20646 37102 20698
rect 6924 20102 6976 20154
rect 6988 20102 7040 20154
rect 7052 20102 7104 20154
rect 7116 20102 7168 20154
rect 7180 20102 7232 20154
rect 18872 20102 18924 20154
rect 18936 20102 18988 20154
rect 19000 20102 19052 20154
rect 19064 20102 19116 20154
rect 19128 20102 19180 20154
rect 30820 20102 30872 20154
rect 30884 20102 30936 20154
rect 30948 20102 31000 20154
rect 31012 20102 31064 20154
rect 31076 20102 31128 20154
rect 42768 20102 42820 20154
rect 42832 20102 42884 20154
rect 42896 20102 42948 20154
rect 42960 20102 43012 20154
rect 43024 20102 43076 20154
rect 1400 19839 1452 19848
rect 1400 19805 1409 19839
rect 1409 19805 1443 19839
rect 1443 19805 1452 19839
rect 1400 19796 1452 19805
rect 12898 19558 12950 19610
rect 12962 19558 13014 19610
rect 13026 19558 13078 19610
rect 13090 19558 13142 19610
rect 13154 19558 13206 19610
rect 24846 19558 24898 19610
rect 24910 19558 24962 19610
rect 24974 19558 25026 19610
rect 25038 19558 25090 19610
rect 25102 19558 25154 19610
rect 36794 19558 36846 19610
rect 36858 19558 36910 19610
rect 36922 19558 36974 19610
rect 36986 19558 37038 19610
rect 37050 19558 37102 19610
rect 1400 19159 1452 19168
rect 1400 19125 1409 19159
rect 1409 19125 1443 19159
rect 1443 19125 1452 19159
rect 1400 19116 1452 19125
rect 48136 19159 48188 19168
rect 48136 19125 48145 19159
rect 48145 19125 48179 19159
rect 48179 19125 48188 19159
rect 48136 19116 48188 19125
rect 6924 19014 6976 19066
rect 6988 19014 7040 19066
rect 7052 19014 7104 19066
rect 7116 19014 7168 19066
rect 7180 19014 7232 19066
rect 18872 19014 18924 19066
rect 18936 19014 18988 19066
rect 19000 19014 19052 19066
rect 19064 19014 19116 19066
rect 19128 19014 19180 19066
rect 30820 19014 30872 19066
rect 30884 19014 30936 19066
rect 30948 19014 31000 19066
rect 31012 19014 31064 19066
rect 31076 19014 31128 19066
rect 42768 19014 42820 19066
rect 42832 19014 42884 19066
rect 42896 19014 42948 19066
rect 42960 19014 43012 19066
rect 43024 19014 43076 19066
rect 1400 18751 1452 18760
rect 1400 18717 1409 18751
rect 1409 18717 1443 18751
rect 1443 18717 1452 18751
rect 1400 18708 1452 18717
rect 48228 18572 48280 18624
rect 12898 18470 12950 18522
rect 12962 18470 13014 18522
rect 13026 18470 13078 18522
rect 13090 18470 13142 18522
rect 13154 18470 13206 18522
rect 24846 18470 24898 18522
rect 24910 18470 24962 18522
rect 24974 18470 25026 18522
rect 25038 18470 25090 18522
rect 25102 18470 25154 18522
rect 36794 18470 36846 18522
rect 36858 18470 36910 18522
rect 36922 18470 36974 18522
rect 36986 18470 37038 18522
rect 37050 18470 37102 18522
rect 48136 18071 48188 18080
rect 48136 18037 48145 18071
rect 48145 18037 48179 18071
rect 48179 18037 48188 18071
rect 48136 18028 48188 18037
rect 6924 17926 6976 17978
rect 6988 17926 7040 17978
rect 7052 17926 7104 17978
rect 7116 17926 7168 17978
rect 7180 17926 7232 17978
rect 18872 17926 18924 17978
rect 18936 17926 18988 17978
rect 19000 17926 19052 17978
rect 19064 17926 19116 17978
rect 19128 17926 19180 17978
rect 30820 17926 30872 17978
rect 30884 17926 30936 17978
rect 30948 17926 31000 17978
rect 31012 17926 31064 17978
rect 31076 17926 31128 17978
rect 42768 17926 42820 17978
rect 42832 17926 42884 17978
rect 42896 17926 42948 17978
rect 42960 17926 43012 17978
rect 43024 17926 43076 17978
rect 12898 17382 12950 17434
rect 12962 17382 13014 17434
rect 13026 17382 13078 17434
rect 13090 17382 13142 17434
rect 13154 17382 13206 17434
rect 24846 17382 24898 17434
rect 24910 17382 24962 17434
rect 24974 17382 25026 17434
rect 25038 17382 25090 17434
rect 25102 17382 25154 17434
rect 36794 17382 36846 17434
rect 36858 17382 36910 17434
rect 36922 17382 36974 17434
rect 36986 17382 37038 17434
rect 37050 17382 37102 17434
rect 48136 16983 48188 16992
rect 48136 16949 48145 16983
rect 48145 16949 48179 16983
rect 48179 16949 48188 16983
rect 48136 16940 48188 16949
rect 6924 16838 6976 16890
rect 6988 16838 7040 16890
rect 7052 16838 7104 16890
rect 7116 16838 7168 16890
rect 7180 16838 7232 16890
rect 18872 16838 18924 16890
rect 18936 16838 18988 16890
rect 19000 16838 19052 16890
rect 19064 16838 19116 16890
rect 19128 16838 19180 16890
rect 30820 16838 30872 16890
rect 30884 16838 30936 16890
rect 30948 16838 31000 16890
rect 31012 16838 31064 16890
rect 31076 16838 31128 16890
rect 42768 16838 42820 16890
rect 42832 16838 42884 16890
rect 42896 16838 42948 16890
rect 42960 16838 43012 16890
rect 43024 16838 43076 16890
rect 48228 16532 48280 16584
rect 12898 16294 12950 16346
rect 12962 16294 13014 16346
rect 13026 16294 13078 16346
rect 13090 16294 13142 16346
rect 13154 16294 13206 16346
rect 24846 16294 24898 16346
rect 24910 16294 24962 16346
rect 24974 16294 25026 16346
rect 25038 16294 25090 16346
rect 25102 16294 25154 16346
rect 36794 16294 36846 16346
rect 36858 16294 36910 16346
rect 36922 16294 36974 16346
rect 36986 16294 37038 16346
rect 37050 16294 37102 16346
rect 1400 15895 1452 15904
rect 1400 15861 1409 15895
rect 1409 15861 1443 15895
rect 1443 15861 1452 15895
rect 1400 15852 1452 15861
rect 48136 15895 48188 15904
rect 48136 15861 48145 15895
rect 48145 15861 48179 15895
rect 48179 15861 48188 15895
rect 48136 15852 48188 15861
rect 6924 15750 6976 15802
rect 6988 15750 7040 15802
rect 7052 15750 7104 15802
rect 7116 15750 7168 15802
rect 7180 15750 7232 15802
rect 18872 15750 18924 15802
rect 18936 15750 18988 15802
rect 19000 15750 19052 15802
rect 19064 15750 19116 15802
rect 19128 15750 19180 15802
rect 30820 15750 30872 15802
rect 30884 15750 30936 15802
rect 30948 15750 31000 15802
rect 31012 15750 31064 15802
rect 31076 15750 31128 15802
rect 42768 15750 42820 15802
rect 42832 15750 42884 15802
rect 42896 15750 42948 15802
rect 42960 15750 43012 15802
rect 43024 15750 43076 15802
rect 1400 15487 1452 15496
rect 1400 15453 1409 15487
rect 1409 15453 1443 15487
rect 1443 15453 1452 15487
rect 1400 15444 1452 15453
rect 12898 15206 12950 15258
rect 12962 15206 13014 15258
rect 13026 15206 13078 15258
rect 13090 15206 13142 15258
rect 13154 15206 13206 15258
rect 24846 15206 24898 15258
rect 24910 15206 24962 15258
rect 24974 15206 25026 15258
rect 25038 15206 25090 15258
rect 25102 15206 25154 15258
rect 36794 15206 36846 15258
rect 36858 15206 36910 15258
rect 36922 15206 36974 15258
rect 36986 15206 37038 15258
rect 37050 15206 37102 15258
rect 22928 15011 22980 15020
rect 22928 14977 22937 15011
rect 22937 14977 22971 15011
rect 22971 14977 22980 15011
rect 22928 14968 22980 14977
rect 22928 14764 22980 14816
rect 6924 14662 6976 14714
rect 6988 14662 7040 14714
rect 7052 14662 7104 14714
rect 7116 14662 7168 14714
rect 7180 14662 7232 14714
rect 18872 14662 18924 14714
rect 18936 14662 18988 14714
rect 19000 14662 19052 14714
rect 19064 14662 19116 14714
rect 19128 14662 19180 14714
rect 30820 14662 30872 14714
rect 30884 14662 30936 14714
rect 30948 14662 31000 14714
rect 31012 14662 31064 14714
rect 31076 14662 31128 14714
rect 42768 14662 42820 14714
rect 42832 14662 42884 14714
rect 42896 14662 42948 14714
rect 42960 14662 43012 14714
rect 43024 14662 43076 14714
rect 1400 14399 1452 14408
rect 1400 14365 1409 14399
rect 1409 14365 1443 14399
rect 1443 14365 1452 14399
rect 1400 14356 1452 14365
rect 38384 14399 38436 14408
rect 38384 14365 38393 14399
rect 38393 14365 38427 14399
rect 38427 14365 38436 14399
rect 38384 14356 38436 14365
rect 39856 14399 39908 14408
rect 39856 14365 39865 14399
rect 39865 14365 39899 14399
rect 39899 14365 39908 14399
rect 39856 14356 39908 14365
rect 48136 14399 48188 14408
rect 48136 14365 48145 14399
rect 48145 14365 48179 14399
rect 48179 14365 48188 14399
rect 48136 14356 48188 14365
rect 45100 14288 45152 14340
rect 25228 14220 25280 14272
rect 43260 14263 43312 14272
rect 43260 14229 43269 14263
rect 43269 14229 43303 14263
rect 43303 14229 43312 14263
rect 43260 14220 43312 14229
rect 12898 14118 12950 14170
rect 12962 14118 13014 14170
rect 13026 14118 13078 14170
rect 13090 14118 13142 14170
rect 13154 14118 13206 14170
rect 24846 14118 24898 14170
rect 24910 14118 24962 14170
rect 24974 14118 25026 14170
rect 25038 14118 25090 14170
rect 25102 14118 25154 14170
rect 36794 14118 36846 14170
rect 36858 14118 36910 14170
rect 36922 14118 36974 14170
rect 36986 14118 37038 14170
rect 37050 14118 37102 14170
rect 25228 13948 25280 14000
rect 30288 13948 30340 14000
rect 26056 13880 26108 13932
rect 45560 14016 45612 14068
rect 43260 13948 43312 14000
rect 47676 13948 47728 14000
rect 24676 13855 24728 13864
rect 24676 13821 24685 13855
rect 24685 13821 24719 13855
rect 24719 13821 24728 13855
rect 24676 13812 24728 13821
rect 29184 13812 29236 13864
rect 32404 13812 32456 13864
rect 39856 13812 39908 13864
rect 46940 13812 46992 13864
rect 1400 13719 1452 13728
rect 1400 13685 1409 13719
rect 1409 13685 1443 13719
rect 1443 13685 1452 13719
rect 1400 13676 1452 13685
rect 26424 13719 26476 13728
rect 26424 13685 26433 13719
rect 26433 13685 26467 13719
rect 26467 13685 26476 13719
rect 26424 13676 26476 13685
rect 27988 13676 28040 13728
rect 33324 13719 33376 13728
rect 33324 13685 33333 13719
rect 33333 13685 33367 13719
rect 33367 13685 33376 13719
rect 33324 13676 33376 13685
rect 48228 13676 48280 13728
rect 6924 13574 6976 13626
rect 6988 13574 7040 13626
rect 7052 13574 7104 13626
rect 7116 13574 7168 13626
rect 7180 13574 7232 13626
rect 18872 13574 18924 13626
rect 18936 13574 18988 13626
rect 19000 13574 19052 13626
rect 19064 13574 19116 13626
rect 19128 13574 19180 13626
rect 30820 13574 30872 13626
rect 30884 13574 30936 13626
rect 30948 13574 31000 13626
rect 31012 13574 31064 13626
rect 31076 13574 31128 13626
rect 42768 13574 42820 13626
rect 42832 13574 42884 13626
rect 42896 13574 42948 13626
rect 42960 13574 43012 13626
rect 43024 13574 43076 13626
rect 27988 13515 28040 13524
rect 27988 13481 27997 13515
rect 27997 13481 28031 13515
rect 28031 13481 28040 13515
rect 27988 13472 28040 13481
rect 38384 13472 38436 13524
rect 26424 13336 26476 13388
rect 32404 13379 32456 13388
rect 32404 13345 32413 13379
rect 32413 13345 32447 13379
rect 32447 13345 32456 13379
rect 32404 13336 32456 13345
rect 24676 13268 24728 13320
rect 34888 13311 34940 13320
rect 34888 13277 34897 13311
rect 34897 13277 34931 13311
rect 34931 13277 34940 13311
rect 34888 13268 34940 13277
rect 48136 13311 48188 13320
rect 48136 13277 48145 13311
rect 48145 13277 48179 13311
rect 48179 13277 48188 13311
rect 48136 13268 48188 13277
rect 46388 13200 46440 13252
rect 22192 13132 22244 13184
rect 12898 13030 12950 13082
rect 12962 13030 13014 13082
rect 13026 13030 13078 13082
rect 13090 13030 13142 13082
rect 13154 13030 13206 13082
rect 24846 13030 24898 13082
rect 24910 13030 24962 13082
rect 24974 13030 25026 13082
rect 25038 13030 25090 13082
rect 25102 13030 25154 13082
rect 36794 13030 36846 13082
rect 36858 13030 36910 13082
rect 36922 13030 36974 13082
rect 36986 13030 37038 13082
rect 37050 13030 37102 13082
rect 29184 12928 29236 12980
rect 45100 12971 45152 12980
rect 45100 12937 45109 12971
rect 45109 12937 45143 12971
rect 45143 12937 45152 12971
rect 45100 12928 45152 12937
rect 46388 12971 46440 12980
rect 46388 12937 46397 12971
rect 46397 12937 46431 12971
rect 46431 12937 46440 12971
rect 46388 12928 46440 12937
rect 47676 12971 47728 12980
rect 47676 12937 47685 12971
rect 47685 12937 47719 12971
rect 47719 12937 47728 12971
rect 47676 12928 47728 12937
rect 33324 12860 33376 12912
rect 46112 12792 46164 12844
rect 30288 12724 30340 12776
rect 26056 12656 26108 12708
rect 1400 12631 1452 12640
rect 1400 12597 1409 12631
rect 1409 12597 1443 12631
rect 1443 12597 1452 12631
rect 1400 12588 1452 12597
rect 34888 12588 34940 12640
rect 39856 12588 39908 12640
rect 6924 12486 6976 12538
rect 6988 12486 7040 12538
rect 7052 12486 7104 12538
rect 7116 12486 7168 12538
rect 7180 12486 7232 12538
rect 18872 12486 18924 12538
rect 18936 12486 18988 12538
rect 19000 12486 19052 12538
rect 19064 12486 19116 12538
rect 19128 12486 19180 12538
rect 30820 12486 30872 12538
rect 30884 12486 30936 12538
rect 30948 12486 31000 12538
rect 31012 12486 31064 12538
rect 31076 12486 31128 12538
rect 42768 12486 42820 12538
rect 42832 12486 42884 12538
rect 42896 12486 42948 12538
rect 42960 12486 43012 12538
rect 43024 12486 43076 12538
rect 48228 12180 48280 12232
rect 12898 11942 12950 11994
rect 12962 11942 13014 11994
rect 13026 11942 13078 11994
rect 13090 11942 13142 11994
rect 13154 11942 13206 11994
rect 24846 11942 24898 11994
rect 24910 11942 24962 11994
rect 24974 11942 25026 11994
rect 25038 11942 25090 11994
rect 25102 11942 25154 11994
rect 36794 11942 36846 11994
rect 36858 11942 36910 11994
rect 36922 11942 36974 11994
rect 36986 11942 37038 11994
rect 37050 11942 37102 11994
rect 1400 11679 1452 11688
rect 1400 11645 1409 11679
rect 1409 11645 1443 11679
rect 1443 11645 1452 11679
rect 1400 11636 1452 11645
rect 48136 11543 48188 11552
rect 48136 11509 48145 11543
rect 48145 11509 48179 11543
rect 48179 11509 48188 11543
rect 48136 11500 48188 11509
rect 6924 11398 6976 11450
rect 6988 11398 7040 11450
rect 7052 11398 7104 11450
rect 7116 11398 7168 11450
rect 7180 11398 7232 11450
rect 18872 11398 18924 11450
rect 18936 11398 18988 11450
rect 19000 11398 19052 11450
rect 19064 11398 19116 11450
rect 19128 11398 19180 11450
rect 30820 11398 30872 11450
rect 30884 11398 30936 11450
rect 30948 11398 31000 11450
rect 31012 11398 31064 11450
rect 31076 11398 31128 11450
rect 42768 11398 42820 11450
rect 42832 11398 42884 11450
rect 42896 11398 42948 11450
rect 42960 11398 43012 11450
rect 43024 11398 43076 11450
rect 47400 11339 47452 11348
rect 47400 11305 47409 11339
rect 47409 11305 47443 11339
rect 47443 11305 47452 11339
rect 47400 11296 47452 11305
rect 46940 11203 46992 11212
rect 46940 11169 46949 11203
rect 46949 11169 46983 11203
rect 46983 11169 46992 11203
rect 46940 11160 46992 11169
rect 47768 11160 47820 11212
rect 47216 11135 47268 11144
rect 47216 11101 47225 11135
rect 47225 11101 47259 11135
rect 47259 11101 47268 11135
rect 47216 11092 47268 11101
rect 1400 11067 1452 11076
rect 1400 11033 1409 11067
rect 1409 11033 1443 11067
rect 1443 11033 1452 11067
rect 1400 11024 1452 11033
rect 12898 10854 12950 10906
rect 12962 10854 13014 10906
rect 13026 10854 13078 10906
rect 13090 10854 13142 10906
rect 13154 10854 13206 10906
rect 24846 10854 24898 10906
rect 24910 10854 24962 10906
rect 24974 10854 25026 10906
rect 25038 10854 25090 10906
rect 25102 10854 25154 10906
rect 36794 10854 36846 10906
rect 36858 10854 36910 10906
rect 36922 10854 36974 10906
rect 36986 10854 37038 10906
rect 37050 10854 37102 10906
rect 47216 10752 47268 10804
rect 47584 10659 47636 10668
rect 47584 10625 47593 10659
rect 47593 10625 47627 10659
rect 47627 10625 47636 10659
rect 47584 10616 47636 10625
rect 47768 10659 47820 10668
rect 47768 10625 47777 10659
rect 47777 10625 47811 10659
rect 47811 10625 47820 10659
rect 47768 10616 47820 10625
rect 6924 10310 6976 10362
rect 6988 10310 7040 10362
rect 7052 10310 7104 10362
rect 7116 10310 7168 10362
rect 7180 10310 7232 10362
rect 18872 10310 18924 10362
rect 18936 10310 18988 10362
rect 19000 10310 19052 10362
rect 19064 10310 19116 10362
rect 19128 10310 19180 10362
rect 30820 10310 30872 10362
rect 30884 10310 30936 10362
rect 30948 10310 31000 10362
rect 31012 10310 31064 10362
rect 31076 10310 31128 10362
rect 42768 10310 42820 10362
rect 42832 10310 42884 10362
rect 42896 10310 42948 10362
rect 42960 10310 43012 10362
rect 43024 10310 43076 10362
rect 48136 10047 48188 10056
rect 48136 10013 48145 10047
rect 48145 10013 48179 10047
rect 48179 10013 48188 10047
rect 48136 10004 48188 10013
rect 12898 9766 12950 9818
rect 12962 9766 13014 9818
rect 13026 9766 13078 9818
rect 13090 9766 13142 9818
rect 13154 9766 13206 9818
rect 24846 9766 24898 9818
rect 24910 9766 24962 9818
rect 24974 9766 25026 9818
rect 25038 9766 25090 9818
rect 25102 9766 25154 9818
rect 36794 9766 36846 9818
rect 36858 9766 36910 9818
rect 36922 9766 36974 9818
rect 36986 9766 37038 9818
rect 37050 9766 37102 9818
rect 45744 9528 45796 9580
rect 47584 9528 47636 9580
rect 46112 9435 46164 9444
rect 46112 9401 46121 9435
rect 46121 9401 46155 9435
rect 46155 9401 46164 9435
rect 46112 9392 46164 9401
rect 6924 9222 6976 9274
rect 6988 9222 7040 9274
rect 7052 9222 7104 9274
rect 7116 9222 7168 9274
rect 7180 9222 7232 9274
rect 18872 9222 18924 9274
rect 18936 9222 18988 9274
rect 19000 9222 19052 9274
rect 19064 9222 19116 9274
rect 19128 9222 19180 9274
rect 30820 9222 30872 9274
rect 30884 9222 30936 9274
rect 30948 9222 31000 9274
rect 31012 9222 31064 9274
rect 31076 9222 31128 9274
rect 42768 9222 42820 9274
rect 42832 9222 42884 9274
rect 42896 9222 42948 9274
rect 42960 9222 43012 9274
rect 43024 9222 43076 9274
rect 1400 8959 1452 8968
rect 1400 8925 1409 8959
rect 1409 8925 1443 8959
rect 1443 8925 1452 8959
rect 1400 8916 1452 8925
rect 48136 8959 48188 8968
rect 48136 8925 48145 8959
rect 48145 8925 48179 8959
rect 48179 8925 48188 8959
rect 48136 8916 48188 8925
rect 12898 8678 12950 8730
rect 12962 8678 13014 8730
rect 13026 8678 13078 8730
rect 13090 8678 13142 8730
rect 13154 8678 13206 8730
rect 24846 8678 24898 8730
rect 24910 8678 24962 8730
rect 24974 8678 25026 8730
rect 25038 8678 25090 8730
rect 25102 8678 25154 8730
rect 36794 8678 36846 8730
rect 36858 8678 36910 8730
rect 36922 8678 36974 8730
rect 36986 8678 37038 8730
rect 37050 8678 37102 8730
rect 1400 8347 1452 8356
rect 1400 8313 1409 8347
rect 1409 8313 1443 8347
rect 1443 8313 1452 8347
rect 1400 8304 1452 8313
rect 6924 8134 6976 8186
rect 6988 8134 7040 8186
rect 7052 8134 7104 8186
rect 7116 8134 7168 8186
rect 7180 8134 7232 8186
rect 18872 8134 18924 8186
rect 18936 8134 18988 8186
rect 19000 8134 19052 8186
rect 19064 8134 19116 8186
rect 19128 8134 19180 8186
rect 30820 8134 30872 8186
rect 30884 8134 30936 8186
rect 30948 8134 31000 8186
rect 31012 8134 31064 8186
rect 31076 8134 31128 8186
rect 42768 8134 42820 8186
rect 42832 8134 42884 8186
rect 42896 8134 42948 8186
rect 42960 8134 43012 8186
rect 43024 8134 43076 8186
rect 47952 8075 48004 8084
rect 47952 8041 47961 8075
rect 47961 8041 47995 8075
rect 47995 8041 48004 8075
rect 47952 8032 48004 8041
rect 48136 7871 48188 7880
rect 48136 7837 48145 7871
rect 48145 7837 48179 7871
rect 48179 7837 48188 7871
rect 48136 7828 48188 7837
rect 1400 7735 1452 7744
rect 1400 7701 1409 7735
rect 1409 7701 1443 7735
rect 1443 7701 1452 7735
rect 1400 7692 1452 7701
rect 12898 7590 12950 7642
rect 12962 7590 13014 7642
rect 13026 7590 13078 7642
rect 13090 7590 13142 7642
rect 13154 7590 13206 7642
rect 24846 7590 24898 7642
rect 24910 7590 24962 7642
rect 24974 7590 25026 7642
rect 25038 7590 25090 7642
rect 25102 7590 25154 7642
rect 36794 7590 36846 7642
rect 36858 7590 36910 7642
rect 36922 7590 36974 7642
rect 36986 7590 37038 7642
rect 37050 7590 37102 7642
rect 1400 7327 1452 7336
rect 1400 7293 1409 7327
rect 1409 7293 1443 7327
rect 1443 7293 1452 7327
rect 1400 7284 1452 7293
rect 48228 7284 48280 7336
rect 6924 7046 6976 7098
rect 6988 7046 7040 7098
rect 7052 7046 7104 7098
rect 7116 7046 7168 7098
rect 7180 7046 7232 7098
rect 18872 7046 18924 7098
rect 18936 7046 18988 7098
rect 19000 7046 19052 7098
rect 19064 7046 19116 7098
rect 19128 7046 19180 7098
rect 30820 7046 30872 7098
rect 30884 7046 30936 7098
rect 30948 7046 31000 7098
rect 31012 7046 31064 7098
rect 31076 7046 31128 7098
rect 42768 7046 42820 7098
rect 42832 7046 42884 7098
rect 42896 7046 42948 7098
rect 42960 7046 43012 7098
rect 43024 7046 43076 7098
rect 12898 6502 12950 6554
rect 12962 6502 13014 6554
rect 13026 6502 13078 6554
rect 13090 6502 13142 6554
rect 13154 6502 13206 6554
rect 24846 6502 24898 6554
rect 24910 6502 24962 6554
rect 24974 6502 25026 6554
rect 25038 6502 25090 6554
rect 25102 6502 25154 6554
rect 36794 6502 36846 6554
rect 36858 6502 36910 6554
rect 36922 6502 36974 6554
rect 36986 6502 37038 6554
rect 37050 6502 37102 6554
rect 1400 6239 1452 6248
rect 1400 6205 1409 6239
rect 1409 6205 1443 6239
rect 1443 6205 1452 6239
rect 1400 6196 1452 6205
rect 48136 6103 48188 6112
rect 48136 6069 48145 6103
rect 48145 6069 48179 6103
rect 48179 6069 48188 6103
rect 48136 6060 48188 6069
rect 6924 5958 6976 6010
rect 6988 5958 7040 6010
rect 7052 5958 7104 6010
rect 7116 5958 7168 6010
rect 7180 5958 7232 6010
rect 18872 5958 18924 6010
rect 18936 5958 18988 6010
rect 19000 5958 19052 6010
rect 19064 5958 19116 6010
rect 19128 5958 19180 6010
rect 30820 5958 30872 6010
rect 30884 5958 30936 6010
rect 30948 5958 31000 6010
rect 31012 5958 31064 6010
rect 31076 5958 31128 6010
rect 42768 5958 42820 6010
rect 42832 5958 42884 6010
rect 42896 5958 42948 6010
rect 42960 5958 43012 6010
rect 43024 5958 43076 6010
rect 1400 5695 1452 5704
rect 1400 5661 1409 5695
rect 1409 5661 1443 5695
rect 1443 5661 1452 5695
rect 1400 5652 1452 5661
rect 12898 5414 12950 5466
rect 12962 5414 13014 5466
rect 13026 5414 13078 5466
rect 13090 5414 13142 5466
rect 13154 5414 13206 5466
rect 24846 5414 24898 5466
rect 24910 5414 24962 5466
rect 24974 5414 25026 5466
rect 25038 5414 25090 5466
rect 25102 5414 25154 5466
rect 36794 5414 36846 5466
rect 36858 5414 36910 5466
rect 36922 5414 36974 5466
rect 36986 5414 37038 5466
rect 37050 5414 37102 5466
rect 1400 5015 1452 5024
rect 1400 4981 1409 5015
rect 1409 4981 1443 5015
rect 1443 4981 1452 5015
rect 1400 4972 1452 4981
rect 48228 4972 48280 5024
rect 6924 4870 6976 4922
rect 6988 4870 7040 4922
rect 7052 4870 7104 4922
rect 7116 4870 7168 4922
rect 7180 4870 7232 4922
rect 18872 4870 18924 4922
rect 18936 4870 18988 4922
rect 19000 4870 19052 4922
rect 19064 4870 19116 4922
rect 19128 4870 19180 4922
rect 30820 4870 30872 4922
rect 30884 4870 30936 4922
rect 30948 4870 31000 4922
rect 31012 4870 31064 4922
rect 31076 4870 31128 4922
rect 42768 4870 42820 4922
rect 42832 4870 42884 4922
rect 42896 4870 42948 4922
rect 42960 4870 43012 4922
rect 43024 4870 43076 4922
rect 48136 4607 48188 4616
rect 48136 4573 48145 4607
rect 48145 4573 48179 4607
rect 48179 4573 48188 4607
rect 48136 4564 48188 4573
rect 12898 4326 12950 4378
rect 12962 4326 13014 4378
rect 13026 4326 13078 4378
rect 13090 4326 13142 4378
rect 13154 4326 13206 4378
rect 24846 4326 24898 4378
rect 24910 4326 24962 4378
rect 24974 4326 25026 4378
rect 25038 4326 25090 4378
rect 25102 4326 25154 4378
rect 36794 4326 36846 4378
rect 36858 4326 36910 4378
rect 36922 4326 36974 4378
rect 36986 4326 37038 4378
rect 37050 4326 37102 4378
rect 2872 3884 2924 3936
rect 47768 3884 47820 3936
rect 48964 3884 49016 3936
rect 6924 3782 6976 3834
rect 6988 3782 7040 3834
rect 7052 3782 7104 3834
rect 7116 3782 7168 3834
rect 7180 3782 7232 3834
rect 18872 3782 18924 3834
rect 18936 3782 18988 3834
rect 19000 3782 19052 3834
rect 19064 3782 19116 3834
rect 19128 3782 19180 3834
rect 30820 3782 30872 3834
rect 30884 3782 30936 3834
rect 30948 3782 31000 3834
rect 31012 3782 31064 3834
rect 31076 3782 31128 3834
rect 42768 3782 42820 3834
rect 42832 3782 42884 3834
rect 42896 3782 42948 3834
rect 42960 3782 43012 3834
rect 43024 3782 43076 3834
rect 2780 3544 2832 3596
rect 1400 3519 1452 3528
rect 1400 3485 1409 3519
rect 1409 3485 1443 3519
rect 1443 3485 1452 3519
rect 1400 3476 1452 3485
rect 2964 3476 3016 3528
rect 46664 3476 46716 3528
rect 48136 3519 48188 3528
rect 48136 3485 48145 3519
rect 48145 3485 48179 3519
rect 48179 3485 48188 3519
rect 48136 3476 48188 3485
rect 49608 3340 49660 3392
rect 12898 3238 12950 3290
rect 12962 3238 13014 3290
rect 13026 3238 13078 3290
rect 13090 3238 13142 3290
rect 13154 3238 13206 3290
rect 24846 3238 24898 3290
rect 24910 3238 24962 3290
rect 24974 3238 25026 3290
rect 25038 3238 25090 3290
rect 25102 3238 25154 3290
rect 36794 3238 36846 3290
rect 36858 3238 36910 3290
rect 36922 3238 36974 3290
rect 36986 3238 37038 3290
rect 37050 3238 37102 3290
rect 45744 3179 45796 3188
rect 45744 3145 45753 3179
rect 45753 3145 45787 3179
rect 45787 3145 45796 3179
rect 45744 3136 45796 3145
rect 45560 3043 45612 3052
rect 45560 3009 45569 3043
rect 45569 3009 45603 3043
rect 45603 3009 45612 3043
rect 45560 3000 45612 3009
rect 3056 2932 3108 2984
rect 3884 2932 3936 2984
rect 30748 2932 30800 2984
rect 36084 2932 36136 2984
rect 46848 2932 46900 2984
rect 47676 2932 47728 2984
rect 20 2864 72 2916
rect 664 2796 716 2848
rect 9036 2796 9088 2848
rect 16764 2796 16816 2848
rect 19340 2796 19392 2848
rect 23204 2796 23256 2848
rect 28356 2796 28408 2848
rect 43812 2796 43864 2848
rect 46756 2796 46808 2848
rect 6924 2694 6976 2746
rect 6988 2694 7040 2746
rect 7052 2694 7104 2746
rect 7116 2694 7168 2746
rect 7180 2694 7232 2746
rect 18872 2694 18924 2746
rect 18936 2694 18988 2746
rect 19000 2694 19052 2746
rect 19064 2694 19116 2746
rect 19128 2694 19180 2746
rect 30820 2694 30872 2746
rect 30884 2694 30936 2746
rect 30948 2694 31000 2746
rect 31012 2694 31064 2746
rect 31076 2694 31128 2746
rect 42768 2694 42820 2746
rect 42832 2694 42884 2746
rect 42896 2694 42948 2746
rect 42960 2694 43012 2746
rect 43024 2694 43076 2746
rect 1308 2388 1360 2440
rect 2596 2431 2648 2440
rect 2596 2397 2605 2431
rect 2605 2397 2639 2431
rect 2639 2397 2648 2431
rect 2596 2388 2648 2397
rect 3240 2431 3292 2440
rect 3240 2397 3249 2431
rect 3249 2397 3283 2431
rect 3283 2397 3292 2431
rect 3240 2388 3292 2397
rect 5172 2431 5224 2440
rect 5172 2397 5181 2431
rect 5181 2397 5215 2431
rect 5215 2397 5224 2431
rect 5172 2388 5224 2397
rect 5816 2431 5868 2440
rect 5816 2397 5825 2431
rect 5825 2397 5859 2431
rect 5859 2397 5868 2431
rect 5816 2388 5868 2397
rect 7104 2431 7156 2440
rect 7104 2397 7113 2431
rect 7113 2397 7147 2431
rect 7147 2397 7156 2431
rect 7104 2388 7156 2397
rect 7748 2431 7800 2440
rect 7748 2397 7757 2431
rect 7757 2397 7791 2431
rect 7791 2397 7800 2431
rect 7748 2388 7800 2397
rect 8392 2431 8444 2440
rect 8392 2397 8401 2431
rect 8401 2397 8435 2431
rect 8435 2397 8444 2431
rect 8392 2388 8444 2397
rect 10324 2431 10376 2440
rect 10324 2397 10333 2431
rect 10333 2397 10367 2431
rect 10367 2397 10376 2431
rect 10324 2388 10376 2397
rect 10968 2431 11020 2440
rect 10968 2397 10977 2431
rect 10977 2397 11011 2431
rect 11011 2397 11020 2431
rect 10968 2388 11020 2397
rect 12808 2388 12860 2440
rect 13544 2388 13596 2440
rect 14832 2388 14884 2440
rect 17408 2431 17460 2440
rect 17408 2397 17417 2431
rect 17417 2397 17451 2431
rect 17451 2397 17460 2431
rect 17408 2388 17460 2397
rect 18052 2431 18104 2440
rect 18052 2397 18061 2431
rect 18061 2397 18095 2431
rect 18095 2397 18104 2431
rect 18052 2388 18104 2397
rect 18696 2431 18748 2440
rect 18696 2397 18705 2431
rect 18705 2397 18739 2431
rect 18739 2397 18748 2431
rect 18696 2388 18748 2397
rect 19984 2431 20036 2440
rect 19984 2397 19993 2431
rect 19993 2397 20027 2431
rect 20027 2397 20036 2431
rect 19984 2388 20036 2397
rect 20628 2431 20680 2440
rect 20628 2397 20637 2431
rect 20637 2397 20671 2431
rect 20671 2397 20680 2431
rect 20628 2388 20680 2397
rect 22192 2431 22244 2440
rect 22192 2397 22201 2431
rect 22201 2397 22235 2431
rect 22235 2397 22244 2431
rect 22192 2388 22244 2397
rect 22928 2431 22980 2440
rect 22928 2397 22937 2431
rect 22937 2397 22971 2431
rect 22971 2397 22980 2431
rect 22928 2388 22980 2397
rect 23848 2431 23900 2440
rect 23848 2397 23857 2431
rect 23857 2397 23891 2431
rect 23891 2397 23900 2431
rect 23848 2388 23900 2397
rect 24492 2388 24544 2440
rect 25228 2431 25280 2440
rect 25228 2397 25237 2431
rect 25237 2397 25271 2431
rect 25271 2397 25280 2431
rect 25228 2388 25280 2397
rect 25780 2388 25832 2440
rect 26424 2388 26476 2440
rect 29000 2388 29052 2440
rect 29644 2388 29696 2440
rect 30288 2388 30340 2440
rect 33508 2388 33560 2440
rect 34152 2388 34204 2440
rect 34796 2388 34848 2440
rect 37372 2388 37424 2440
rect 38660 2388 38712 2440
rect 39304 2388 39356 2440
rect 40592 2388 40644 2440
rect 41236 2388 41288 2440
rect 42524 2388 42576 2440
rect 46388 2388 46440 2440
rect 47032 2388 47084 2440
rect 4528 2295 4580 2304
rect 4528 2261 4537 2295
rect 4537 2261 4571 2295
rect 4571 2261 4580 2295
rect 4528 2252 4580 2261
rect 9680 2295 9732 2304
rect 9680 2261 9689 2295
rect 9689 2261 9723 2295
rect 9723 2261 9732 2295
rect 9680 2252 9732 2261
rect 11612 2252 11664 2304
rect 12256 2252 12308 2304
rect 16120 2295 16172 2304
rect 16120 2261 16129 2295
rect 16129 2261 16163 2295
rect 16163 2261 16172 2295
rect 16120 2252 16172 2261
rect 21272 2295 21324 2304
rect 21272 2261 21281 2295
rect 21281 2261 21315 2295
rect 21315 2261 21324 2295
rect 21272 2252 21324 2261
rect 21916 2252 21968 2304
rect 22560 2252 22612 2304
rect 27068 2252 27120 2304
rect 27712 2252 27764 2304
rect 32220 2252 32272 2304
rect 32864 2252 32916 2304
rect 35440 2252 35492 2304
rect 41880 2252 41932 2304
rect 43168 2252 43220 2304
rect 44456 2252 44508 2304
rect 45100 2252 45152 2304
rect 12898 2150 12950 2202
rect 12962 2150 13014 2202
rect 13026 2150 13078 2202
rect 13090 2150 13142 2202
rect 13154 2150 13206 2202
rect 24846 2150 24898 2202
rect 24910 2150 24962 2202
rect 24974 2150 25026 2202
rect 25038 2150 25090 2202
rect 25102 2150 25154 2202
rect 36794 2150 36846 2202
rect 36858 2150 36910 2202
rect 36922 2150 36974 2202
rect 36986 2150 37038 2202
rect 37050 2150 37102 2202
<< metal2 >>
rect 18 29200 74 30000
rect 662 29200 718 30000
rect 1306 29200 1362 30000
rect 1950 29322 2006 30000
rect 1950 29294 2084 29322
rect 1950 29200 2006 29294
rect 32 27470 60 29200
rect 20 27464 72 27470
rect 20 27406 72 27412
rect 676 27130 704 29200
rect 1320 27538 1348 29200
rect 1398 27976 1454 27985
rect 1398 27911 1454 27920
rect 1308 27532 1360 27538
rect 1308 27474 1360 27480
rect 664 27124 716 27130
rect 664 27066 716 27072
rect 1412 26994 1440 27911
rect 2056 27606 2084 29294
rect 2594 29200 2650 30000
rect 2870 29336 2926 29345
rect 2870 29271 2926 29280
rect 2778 28656 2834 28665
rect 2778 28591 2834 28600
rect 2044 27600 2096 27606
rect 2044 27542 2096 27548
rect 1490 27296 1546 27305
rect 1490 27231 1546 27240
rect 1400 26988 1452 26994
rect 1400 26930 1452 26936
rect 1400 26376 1452 26382
rect 1400 26318 1452 26324
rect 1412 25945 1440 26318
rect 1398 25936 1454 25945
rect 1504 25906 1532 27231
rect 2792 26586 2820 28591
rect 2884 27062 2912 29271
rect 3238 29200 3294 30000
rect 3882 29322 3938 30000
rect 3882 29294 4016 29322
rect 3882 29200 3938 29294
rect 3988 27606 4016 29294
rect 4526 29200 4582 30000
rect 5170 29200 5226 30000
rect 5814 29200 5870 30000
rect 6458 29322 6514 30000
rect 7102 29322 7158 30000
rect 6458 29294 6592 29322
rect 6458 29200 6514 29294
rect 5184 27606 5212 29200
rect 5828 27606 5856 29200
rect 3976 27600 4028 27606
rect 3976 27542 4028 27548
rect 5172 27600 5224 27606
rect 5172 27542 5224 27548
rect 5816 27600 5868 27606
rect 5816 27542 5868 27548
rect 2872 27056 2924 27062
rect 2872 26998 2924 27004
rect 6564 26994 6592 29294
rect 7102 29294 7328 29322
rect 7102 29200 7158 29294
rect 6924 27772 7232 27781
rect 6924 27770 6930 27772
rect 6986 27770 7010 27772
rect 7066 27770 7090 27772
rect 7146 27770 7170 27772
rect 7226 27770 7232 27772
rect 6986 27718 6988 27770
rect 7168 27718 7170 27770
rect 6924 27716 6930 27718
rect 6986 27716 7010 27718
rect 7066 27716 7090 27718
rect 7146 27716 7170 27718
rect 7226 27716 7232 27718
rect 6924 27707 7232 27716
rect 7300 27538 7328 29294
rect 7746 29200 7802 30000
rect 8390 29200 8446 30000
rect 9034 29322 9090 30000
rect 9034 29294 9168 29322
rect 9034 29200 9090 29294
rect 7760 27606 7788 29200
rect 8404 27606 8432 29200
rect 7748 27600 7800 27606
rect 7748 27542 7800 27548
rect 8392 27600 8444 27606
rect 8392 27542 8444 27548
rect 7288 27532 7340 27538
rect 7288 27474 7340 27480
rect 9140 26994 9168 29294
rect 9678 29200 9734 30000
rect 10322 29200 10378 30000
rect 10966 29200 11022 30000
rect 11610 29322 11666 30000
rect 12254 29322 12310 30000
rect 12898 29322 12954 30000
rect 13542 29322 13598 30000
rect 11610 29294 11744 29322
rect 11610 29200 11666 29294
rect 9692 27538 9720 29200
rect 10336 27606 10364 29200
rect 10980 27606 11008 29200
rect 10324 27600 10376 27606
rect 10324 27542 10376 27548
rect 10968 27600 11020 27606
rect 10968 27542 11020 27548
rect 11716 27538 11744 29294
rect 12254 29294 12388 29322
rect 12254 29200 12310 29294
rect 12360 27538 12388 29294
rect 12898 29294 13032 29322
rect 12898 29200 12954 29294
rect 13004 27538 13032 29294
rect 13542 29294 13768 29322
rect 13542 29200 13598 29294
rect 13740 27554 13768 29294
rect 14186 29200 14242 30000
rect 14830 29322 14886 30000
rect 15474 29322 15530 30000
rect 16118 29322 16174 30000
rect 14830 29294 14964 29322
rect 14830 29200 14886 29294
rect 14936 27606 14964 29294
rect 15474 29294 15608 29322
rect 15474 29200 15530 29294
rect 15580 27606 15608 29294
rect 16118 29294 16528 29322
rect 16118 29200 16174 29294
rect 13820 27600 13872 27606
rect 13740 27548 13820 27554
rect 13740 27542 13872 27548
rect 14924 27600 14976 27606
rect 14924 27542 14976 27548
rect 15568 27600 15620 27606
rect 15568 27542 15620 27548
rect 16500 27554 16528 29294
rect 16762 29200 16818 30000
rect 17406 29200 17462 30000
rect 18050 29200 18106 30000
rect 18694 29200 18750 30000
rect 19338 29322 19394 30000
rect 19338 29294 19472 29322
rect 19338 29200 19394 29294
rect 18064 27606 18092 29200
rect 18708 27606 18736 29200
rect 18872 27772 19180 27781
rect 18872 27770 18878 27772
rect 18934 27770 18958 27772
rect 19014 27770 19038 27772
rect 19094 27770 19118 27772
rect 19174 27770 19180 27772
rect 18934 27718 18936 27770
rect 19116 27718 19118 27770
rect 18872 27716 18878 27718
rect 18934 27716 18958 27718
rect 19014 27716 19038 27718
rect 19094 27716 19118 27718
rect 19174 27716 19180 27718
rect 18872 27707 19180 27716
rect 18052 27600 18104 27606
rect 9680 27532 9732 27538
rect 9680 27474 9732 27480
rect 11704 27532 11756 27538
rect 11704 27474 11756 27480
rect 12348 27532 12400 27538
rect 12348 27474 12400 27480
rect 12992 27532 13044 27538
rect 13740 27526 13860 27542
rect 16500 27538 16620 27554
rect 18052 27542 18104 27548
rect 18696 27600 18748 27606
rect 18696 27542 18748 27548
rect 16500 27532 16632 27538
rect 16500 27526 16580 27532
rect 12992 27474 13044 27480
rect 16580 27474 16632 27480
rect 12898 27228 13206 27237
rect 12898 27226 12904 27228
rect 12960 27226 12984 27228
rect 13040 27226 13064 27228
rect 13120 27226 13144 27228
rect 13200 27226 13206 27228
rect 12960 27174 12962 27226
rect 13142 27174 13144 27226
rect 12898 27172 12904 27174
rect 12960 27172 12984 27174
rect 13040 27172 13064 27174
rect 13120 27172 13144 27174
rect 13200 27172 13206 27174
rect 12898 27163 13206 27172
rect 19444 26994 19472 29294
rect 19982 29200 20038 30000
rect 20626 29200 20682 30000
rect 21270 29200 21326 30000
rect 21914 29322 21970 30000
rect 21914 29294 22048 29322
rect 21914 29200 21970 29294
rect 19996 27606 20024 29200
rect 20640 27606 20668 29200
rect 21284 27606 21312 29200
rect 19984 27600 20036 27606
rect 19984 27542 20036 27548
rect 20628 27600 20680 27606
rect 20628 27542 20680 27548
rect 21272 27600 21324 27606
rect 21272 27542 21324 27548
rect 22020 26994 22048 29294
rect 22558 29200 22614 30000
rect 23202 29200 23258 30000
rect 23846 29200 23902 30000
rect 24490 29322 24546 30000
rect 25134 29322 25190 30000
rect 25778 29322 25834 30000
rect 24490 29294 24624 29322
rect 24490 29200 24546 29294
rect 22572 27538 22600 29200
rect 23216 27606 23244 29200
rect 23204 27600 23256 27606
rect 23204 27542 23256 27548
rect 23860 27538 23888 29200
rect 24596 27606 24624 29294
rect 25134 29294 25268 29322
rect 25134 29200 25190 29294
rect 25240 27606 25268 29294
rect 25778 29294 25912 29322
rect 25778 29200 25834 29294
rect 25884 27606 25912 29294
rect 26422 29200 26478 30000
rect 27066 29200 27122 30000
rect 27710 29322 27766 30000
rect 28354 29322 28410 30000
rect 27710 29294 27844 29322
rect 27710 29200 27766 29294
rect 26436 27606 26464 29200
rect 24584 27600 24636 27606
rect 24584 27542 24636 27548
rect 25228 27600 25280 27606
rect 25228 27542 25280 27548
rect 25872 27600 25924 27606
rect 25872 27542 25924 27548
rect 26424 27600 26476 27606
rect 26424 27542 26476 27548
rect 27816 27538 27844 29294
rect 28354 29294 28488 29322
rect 28354 29200 28410 29294
rect 28460 27538 28488 29294
rect 28998 29200 29054 30000
rect 29642 29200 29698 30000
rect 30286 29200 30342 30000
rect 30930 29322 30986 30000
rect 30930 29294 31248 29322
rect 30930 29200 30986 29294
rect 29012 27538 29040 29200
rect 30300 27554 30328 29200
rect 30820 27772 31128 27781
rect 30820 27770 30826 27772
rect 30882 27770 30906 27772
rect 30962 27770 30986 27772
rect 31042 27770 31066 27772
rect 31122 27770 31128 27772
rect 30882 27718 30884 27770
rect 31064 27718 31066 27770
rect 30820 27716 30826 27718
rect 30882 27716 30906 27718
rect 30962 27716 30986 27718
rect 31042 27716 31066 27718
rect 31122 27716 31128 27718
rect 30820 27707 31128 27716
rect 31220 27606 31248 29294
rect 31574 29200 31630 30000
rect 32218 29322 32274 30000
rect 32218 29294 32352 29322
rect 32218 29200 32274 29294
rect 32324 27606 32352 29294
rect 32862 29200 32918 30000
rect 33506 29322 33562 30000
rect 34150 29322 34206 30000
rect 33506 29294 33640 29322
rect 33506 29200 33562 29294
rect 33612 27606 33640 29294
rect 34150 29294 34468 29322
rect 34150 29200 34206 29294
rect 30380 27600 30432 27606
rect 30300 27548 30380 27554
rect 30300 27542 30432 27548
rect 31208 27600 31260 27606
rect 31208 27542 31260 27548
rect 32312 27600 32364 27606
rect 32312 27542 32364 27548
rect 33600 27600 33652 27606
rect 33600 27542 33652 27548
rect 34440 27554 34468 29294
rect 34794 29200 34850 30000
rect 35438 29322 35494 30000
rect 36082 29322 36138 30000
rect 36726 29322 36782 30000
rect 35438 29294 35848 29322
rect 35438 29200 35494 29294
rect 34520 27600 34572 27606
rect 34440 27548 34520 27554
rect 34440 27542 34572 27548
rect 22560 27532 22612 27538
rect 22560 27474 22612 27480
rect 23848 27532 23900 27538
rect 23848 27474 23900 27480
rect 27804 27532 27856 27538
rect 27804 27474 27856 27480
rect 28448 27532 28500 27538
rect 28448 27474 28500 27480
rect 29000 27532 29052 27538
rect 30300 27526 30420 27542
rect 34440 27526 34560 27542
rect 34808 27538 34836 29200
rect 35820 27554 35848 29294
rect 36082 29294 36216 29322
rect 36082 29200 36138 29294
rect 35820 27538 35940 27554
rect 34796 27532 34848 27538
rect 29000 27474 29052 27480
rect 35820 27532 35952 27538
rect 35820 27526 35900 27532
rect 34796 27474 34848 27480
rect 35900 27474 35952 27480
rect 22928 27396 22980 27402
rect 22928 27338 22980 27344
rect 6552 26988 6604 26994
rect 6552 26930 6604 26936
rect 9128 26988 9180 26994
rect 9128 26930 9180 26936
rect 19432 26988 19484 26994
rect 19432 26930 19484 26936
rect 22008 26988 22060 26994
rect 22008 26930 22060 26936
rect 6924 26684 7232 26693
rect 6924 26682 6930 26684
rect 6986 26682 7010 26684
rect 7066 26682 7090 26684
rect 7146 26682 7170 26684
rect 7226 26682 7232 26684
rect 6986 26630 6988 26682
rect 7168 26630 7170 26682
rect 6924 26628 6930 26630
rect 6986 26628 7010 26630
rect 7066 26628 7090 26630
rect 7146 26628 7170 26630
rect 7226 26628 7232 26630
rect 6924 26619 7232 26628
rect 18872 26684 19180 26693
rect 18872 26682 18878 26684
rect 18934 26682 18958 26684
rect 19014 26682 19038 26684
rect 19094 26682 19118 26684
rect 19174 26682 19180 26684
rect 18934 26630 18936 26682
rect 19116 26630 19118 26682
rect 18872 26628 18878 26630
rect 18934 26628 18958 26630
rect 19014 26628 19038 26630
rect 19094 26628 19118 26630
rect 19174 26628 19180 26630
rect 18872 26619 19180 26628
rect 2780 26580 2832 26586
rect 2780 26522 2832 26528
rect 12898 26140 13206 26149
rect 12898 26138 12904 26140
rect 12960 26138 12984 26140
rect 13040 26138 13064 26140
rect 13120 26138 13144 26140
rect 13200 26138 13206 26140
rect 12960 26086 12962 26138
rect 13142 26086 13144 26138
rect 12898 26084 12904 26086
rect 12960 26084 12984 26086
rect 13040 26084 13064 26086
rect 13120 26084 13144 26086
rect 13200 26084 13206 26086
rect 12898 26075 13206 26084
rect 1398 25871 1454 25880
rect 1492 25900 1544 25906
rect 1492 25842 1544 25848
rect 6924 25596 7232 25605
rect 6924 25594 6930 25596
rect 6986 25594 7010 25596
rect 7066 25594 7090 25596
rect 7146 25594 7170 25596
rect 7226 25594 7232 25596
rect 6986 25542 6988 25594
rect 7168 25542 7170 25594
rect 6924 25540 6930 25542
rect 6986 25540 7010 25542
rect 7066 25540 7090 25542
rect 7146 25540 7170 25542
rect 7226 25540 7232 25542
rect 6924 25531 7232 25540
rect 18872 25596 19180 25605
rect 18872 25594 18878 25596
rect 18934 25594 18958 25596
rect 19014 25594 19038 25596
rect 19094 25594 19118 25596
rect 19174 25594 19180 25596
rect 18934 25542 18936 25594
rect 19116 25542 19118 25594
rect 18872 25540 18878 25542
rect 18934 25540 18958 25542
rect 19014 25540 19038 25542
rect 19094 25540 19118 25542
rect 19174 25540 19180 25542
rect 18872 25531 19180 25540
rect 1400 25288 1452 25294
rect 1398 25256 1400 25265
rect 1452 25256 1454 25265
rect 1398 25191 1454 25200
rect 12898 25052 13206 25061
rect 12898 25050 12904 25052
rect 12960 25050 12984 25052
rect 13040 25050 13064 25052
rect 13120 25050 13144 25052
rect 13200 25050 13206 25052
rect 12960 24998 12962 25050
rect 13142 24998 13144 25050
rect 12898 24996 12904 24998
rect 12960 24996 12984 24998
rect 13040 24996 13064 24998
rect 13120 24996 13144 24998
rect 13200 24996 13206 24998
rect 12898 24987 13206 24996
rect 1400 24608 1452 24614
rect 1398 24576 1400 24585
rect 1452 24576 1454 24585
rect 1398 24511 1454 24520
rect 6924 24508 7232 24517
rect 6924 24506 6930 24508
rect 6986 24506 7010 24508
rect 7066 24506 7090 24508
rect 7146 24506 7170 24508
rect 7226 24506 7232 24508
rect 6986 24454 6988 24506
rect 7168 24454 7170 24506
rect 6924 24452 6930 24454
rect 6986 24452 7010 24454
rect 7066 24452 7090 24454
rect 7146 24452 7170 24454
rect 7226 24452 7232 24454
rect 6924 24443 7232 24452
rect 18872 24508 19180 24517
rect 18872 24506 18878 24508
rect 18934 24506 18958 24508
rect 19014 24506 19038 24508
rect 19094 24506 19118 24508
rect 19174 24506 19180 24508
rect 18934 24454 18936 24506
rect 19116 24454 19118 24506
rect 18872 24452 18878 24454
rect 18934 24452 18958 24454
rect 19014 24452 19038 24454
rect 19094 24452 19118 24454
rect 19174 24452 19180 24454
rect 18872 24443 19180 24452
rect 1400 24064 1452 24070
rect 1400 24006 1452 24012
rect 1412 23905 1440 24006
rect 12898 23964 13206 23973
rect 12898 23962 12904 23964
rect 12960 23962 12984 23964
rect 13040 23962 13064 23964
rect 13120 23962 13144 23964
rect 13200 23962 13206 23964
rect 12960 23910 12962 23962
rect 13142 23910 13144 23962
rect 12898 23908 12904 23910
rect 12960 23908 12984 23910
rect 13040 23908 13064 23910
rect 13120 23908 13144 23910
rect 13200 23908 13206 23910
rect 1398 23896 1454 23905
rect 12898 23899 13206 23908
rect 1398 23831 1454 23840
rect 1400 23520 1452 23526
rect 1400 23462 1452 23468
rect 1412 23225 1440 23462
rect 6924 23420 7232 23429
rect 6924 23418 6930 23420
rect 6986 23418 7010 23420
rect 7066 23418 7090 23420
rect 7146 23418 7170 23420
rect 7226 23418 7232 23420
rect 6986 23366 6988 23418
rect 7168 23366 7170 23418
rect 6924 23364 6930 23366
rect 6986 23364 7010 23366
rect 7066 23364 7090 23366
rect 7146 23364 7170 23366
rect 7226 23364 7232 23366
rect 6924 23355 7232 23364
rect 18872 23420 19180 23429
rect 18872 23418 18878 23420
rect 18934 23418 18958 23420
rect 19014 23418 19038 23420
rect 19094 23418 19118 23420
rect 19174 23418 19180 23420
rect 18934 23366 18936 23418
rect 19116 23366 19118 23418
rect 18872 23364 18878 23366
rect 18934 23364 18958 23366
rect 19014 23364 19038 23366
rect 19094 23364 19118 23366
rect 19174 23364 19180 23366
rect 18872 23355 19180 23364
rect 1398 23216 1454 23225
rect 1398 23151 1454 23160
rect 12898 22876 13206 22885
rect 12898 22874 12904 22876
rect 12960 22874 12984 22876
rect 13040 22874 13064 22876
rect 13120 22874 13144 22876
rect 13200 22874 13206 22876
rect 12960 22822 12962 22874
rect 13142 22822 13144 22874
rect 12898 22820 12904 22822
rect 12960 22820 12984 22822
rect 13040 22820 13064 22822
rect 13120 22820 13144 22822
rect 13200 22820 13206 22822
rect 12898 22811 13206 22820
rect 6924 22332 7232 22341
rect 6924 22330 6930 22332
rect 6986 22330 7010 22332
rect 7066 22330 7090 22332
rect 7146 22330 7170 22332
rect 7226 22330 7232 22332
rect 6986 22278 6988 22330
rect 7168 22278 7170 22330
rect 6924 22276 6930 22278
rect 6986 22276 7010 22278
rect 7066 22276 7090 22278
rect 7146 22276 7170 22278
rect 7226 22276 7232 22278
rect 6924 22267 7232 22276
rect 18872 22332 19180 22341
rect 18872 22330 18878 22332
rect 18934 22330 18958 22332
rect 19014 22330 19038 22332
rect 19094 22330 19118 22332
rect 19174 22330 19180 22332
rect 18934 22278 18936 22330
rect 19116 22278 19118 22330
rect 18872 22276 18878 22278
rect 18934 22276 18958 22278
rect 19014 22276 19038 22278
rect 19094 22276 19118 22278
rect 19174 22276 19180 22278
rect 18872 22267 19180 22276
rect 1400 22024 1452 22030
rect 1400 21966 1452 21972
rect 1412 21865 1440 21966
rect 1398 21856 1454 21865
rect 1398 21791 1454 21800
rect 12898 21788 13206 21797
rect 12898 21786 12904 21788
rect 12960 21786 12984 21788
rect 13040 21786 13064 21788
rect 13120 21786 13144 21788
rect 13200 21786 13206 21788
rect 12960 21734 12962 21786
rect 13142 21734 13144 21786
rect 12898 21732 12904 21734
rect 12960 21732 12984 21734
rect 13040 21732 13064 21734
rect 13120 21732 13144 21734
rect 13200 21732 13206 21734
rect 12898 21723 13206 21732
rect 1400 21344 1452 21350
rect 1400 21286 1452 21292
rect 1412 21185 1440 21286
rect 6924 21244 7232 21253
rect 6924 21242 6930 21244
rect 6986 21242 7010 21244
rect 7066 21242 7090 21244
rect 7146 21242 7170 21244
rect 7226 21242 7232 21244
rect 6986 21190 6988 21242
rect 7168 21190 7170 21242
rect 6924 21188 6930 21190
rect 6986 21188 7010 21190
rect 7066 21188 7090 21190
rect 7146 21188 7170 21190
rect 7226 21188 7232 21190
rect 1398 21176 1454 21185
rect 6924 21179 7232 21188
rect 18872 21244 19180 21253
rect 18872 21242 18878 21244
rect 18934 21242 18958 21244
rect 19014 21242 19038 21244
rect 19094 21242 19118 21244
rect 19174 21242 19180 21244
rect 18934 21190 18936 21242
rect 19116 21190 19118 21242
rect 18872 21188 18878 21190
rect 18934 21188 18958 21190
rect 19014 21188 19038 21190
rect 19094 21188 19118 21190
rect 19174 21188 19180 21190
rect 18872 21179 19180 21188
rect 1398 21111 1454 21120
rect 1400 20936 1452 20942
rect 1400 20878 1452 20884
rect 1412 20505 1440 20878
rect 12898 20700 13206 20709
rect 12898 20698 12904 20700
rect 12960 20698 12984 20700
rect 13040 20698 13064 20700
rect 13120 20698 13144 20700
rect 13200 20698 13206 20700
rect 12960 20646 12962 20698
rect 13142 20646 13144 20698
rect 12898 20644 12904 20646
rect 12960 20644 12984 20646
rect 13040 20644 13064 20646
rect 13120 20644 13144 20646
rect 13200 20644 13206 20646
rect 12898 20635 13206 20644
rect 1398 20496 1454 20505
rect 1398 20431 1454 20440
rect 6924 20156 7232 20165
rect 6924 20154 6930 20156
rect 6986 20154 7010 20156
rect 7066 20154 7090 20156
rect 7146 20154 7170 20156
rect 7226 20154 7232 20156
rect 6986 20102 6988 20154
rect 7168 20102 7170 20154
rect 6924 20100 6930 20102
rect 6986 20100 7010 20102
rect 7066 20100 7090 20102
rect 7146 20100 7170 20102
rect 7226 20100 7232 20102
rect 6924 20091 7232 20100
rect 18872 20156 19180 20165
rect 18872 20154 18878 20156
rect 18934 20154 18958 20156
rect 19014 20154 19038 20156
rect 19094 20154 19118 20156
rect 19174 20154 19180 20156
rect 18934 20102 18936 20154
rect 19116 20102 19118 20154
rect 18872 20100 18878 20102
rect 18934 20100 18958 20102
rect 19014 20100 19038 20102
rect 19094 20100 19118 20102
rect 19174 20100 19180 20102
rect 18872 20091 19180 20100
rect 1400 19848 1452 19854
rect 1398 19816 1400 19825
rect 1452 19816 1454 19825
rect 1398 19751 1454 19760
rect 12898 19612 13206 19621
rect 12898 19610 12904 19612
rect 12960 19610 12984 19612
rect 13040 19610 13064 19612
rect 13120 19610 13144 19612
rect 13200 19610 13206 19612
rect 12960 19558 12962 19610
rect 13142 19558 13144 19610
rect 12898 19556 12904 19558
rect 12960 19556 12984 19558
rect 13040 19556 13064 19558
rect 13120 19556 13144 19558
rect 13200 19556 13206 19558
rect 12898 19547 13206 19556
rect 1400 19168 1452 19174
rect 1398 19136 1400 19145
rect 1452 19136 1454 19145
rect 1398 19071 1454 19080
rect 6924 19068 7232 19077
rect 6924 19066 6930 19068
rect 6986 19066 7010 19068
rect 7066 19066 7090 19068
rect 7146 19066 7170 19068
rect 7226 19066 7232 19068
rect 6986 19014 6988 19066
rect 7168 19014 7170 19066
rect 6924 19012 6930 19014
rect 6986 19012 7010 19014
rect 7066 19012 7090 19014
rect 7146 19012 7170 19014
rect 7226 19012 7232 19014
rect 6924 19003 7232 19012
rect 18872 19068 19180 19077
rect 18872 19066 18878 19068
rect 18934 19066 18958 19068
rect 19014 19066 19038 19068
rect 19094 19066 19118 19068
rect 19174 19066 19180 19068
rect 18934 19014 18936 19066
rect 19116 19014 19118 19066
rect 18872 19012 18878 19014
rect 18934 19012 18958 19014
rect 19014 19012 19038 19014
rect 19094 19012 19118 19014
rect 19174 19012 19180 19014
rect 18872 19003 19180 19012
rect 1400 18760 1452 18766
rect 1400 18702 1452 18708
rect 1412 18465 1440 18702
rect 12898 18524 13206 18533
rect 12898 18522 12904 18524
rect 12960 18522 12984 18524
rect 13040 18522 13064 18524
rect 13120 18522 13144 18524
rect 13200 18522 13206 18524
rect 12960 18470 12962 18522
rect 13142 18470 13144 18522
rect 12898 18468 12904 18470
rect 12960 18468 12984 18470
rect 13040 18468 13064 18470
rect 13120 18468 13144 18470
rect 13200 18468 13206 18470
rect 1398 18456 1454 18465
rect 12898 18459 13206 18468
rect 1398 18391 1454 18400
rect 6924 17980 7232 17989
rect 6924 17978 6930 17980
rect 6986 17978 7010 17980
rect 7066 17978 7090 17980
rect 7146 17978 7170 17980
rect 7226 17978 7232 17980
rect 6986 17926 6988 17978
rect 7168 17926 7170 17978
rect 6924 17924 6930 17926
rect 6986 17924 7010 17926
rect 7066 17924 7090 17926
rect 7146 17924 7170 17926
rect 7226 17924 7232 17926
rect 6924 17915 7232 17924
rect 18872 17980 19180 17989
rect 18872 17978 18878 17980
rect 18934 17978 18958 17980
rect 19014 17978 19038 17980
rect 19094 17978 19118 17980
rect 19174 17978 19180 17980
rect 18934 17926 18936 17978
rect 19116 17926 19118 17978
rect 18872 17924 18878 17926
rect 18934 17924 18958 17926
rect 19014 17924 19038 17926
rect 19094 17924 19118 17926
rect 19174 17924 19180 17926
rect 18872 17915 19180 17924
rect 12898 17436 13206 17445
rect 12898 17434 12904 17436
rect 12960 17434 12984 17436
rect 13040 17434 13064 17436
rect 13120 17434 13144 17436
rect 13200 17434 13206 17436
rect 12960 17382 12962 17434
rect 13142 17382 13144 17434
rect 12898 17380 12904 17382
rect 12960 17380 12984 17382
rect 13040 17380 13064 17382
rect 13120 17380 13144 17382
rect 13200 17380 13206 17382
rect 12898 17371 13206 17380
rect 6924 16892 7232 16901
rect 6924 16890 6930 16892
rect 6986 16890 7010 16892
rect 7066 16890 7090 16892
rect 7146 16890 7170 16892
rect 7226 16890 7232 16892
rect 6986 16838 6988 16890
rect 7168 16838 7170 16890
rect 6924 16836 6930 16838
rect 6986 16836 7010 16838
rect 7066 16836 7090 16838
rect 7146 16836 7170 16838
rect 7226 16836 7232 16838
rect 6924 16827 7232 16836
rect 18872 16892 19180 16901
rect 18872 16890 18878 16892
rect 18934 16890 18958 16892
rect 19014 16890 19038 16892
rect 19094 16890 19118 16892
rect 19174 16890 19180 16892
rect 18934 16838 18936 16890
rect 19116 16838 19118 16890
rect 18872 16836 18878 16838
rect 18934 16836 18958 16838
rect 19014 16836 19038 16838
rect 19094 16836 19118 16838
rect 19174 16836 19180 16838
rect 18872 16827 19180 16836
rect 12898 16348 13206 16357
rect 12898 16346 12904 16348
rect 12960 16346 12984 16348
rect 13040 16346 13064 16348
rect 13120 16346 13144 16348
rect 13200 16346 13206 16348
rect 12960 16294 12962 16346
rect 13142 16294 13144 16346
rect 12898 16292 12904 16294
rect 12960 16292 12984 16294
rect 13040 16292 13064 16294
rect 13120 16292 13144 16294
rect 13200 16292 13206 16294
rect 12898 16283 13206 16292
rect 1400 15904 1452 15910
rect 1400 15846 1452 15852
rect 1412 15745 1440 15846
rect 6924 15804 7232 15813
rect 6924 15802 6930 15804
rect 6986 15802 7010 15804
rect 7066 15802 7090 15804
rect 7146 15802 7170 15804
rect 7226 15802 7232 15804
rect 6986 15750 6988 15802
rect 7168 15750 7170 15802
rect 6924 15748 6930 15750
rect 6986 15748 7010 15750
rect 7066 15748 7090 15750
rect 7146 15748 7170 15750
rect 7226 15748 7232 15750
rect 1398 15736 1454 15745
rect 6924 15739 7232 15748
rect 18872 15804 19180 15813
rect 18872 15802 18878 15804
rect 18934 15802 18958 15804
rect 19014 15802 19038 15804
rect 19094 15802 19118 15804
rect 19174 15802 19180 15804
rect 18934 15750 18936 15802
rect 19116 15750 19118 15802
rect 18872 15748 18878 15750
rect 18934 15748 18958 15750
rect 19014 15748 19038 15750
rect 19094 15748 19118 15750
rect 19174 15748 19180 15750
rect 18872 15739 19180 15748
rect 1398 15671 1454 15680
rect 1400 15496 1452 15502
rect 1400 15438 1452 15444
rect 1412 15065 1440 15438
rect 12898 15260 13206 15269
rect 12898 15258 12904 15260
rect 12960 15258 12984 15260
rect 13040 15258 13064 15260
rect 13120 15258 13144 15260
rect 13200 15258 13206 15260
rect 12960 15206 12962 15258
rect 13142 15206 13144 15258
rect 12898 15204 12904 15206
rect 12960 15204 12984 15206
rect 13040 15204 13064 15206
rect 13120 15204 13144 15206
rect 13200 15204 13206 15206
rect 12898 15195 13206 15204
rect 1398 15056 1454 15065
rect 22940 15026 22968 27338
rect 24846 27228 25154 27237
rect 24846 27226 24852 27228
rect 24908 27226 24932 27228
rect 24988 27226 25012 27228
rect 25068 27226 25092 27228
rect 25148 27226 25154 27228
rect 24908 27174 24910 27226
rect 25090 27174 25092 27226
rect 24846 27172 24852 27174
rect 24908 27172 24932 27174
rect 24988 27172 25012 27174
rect 25068 27172 25092 27174
rect 25148 27172 25154 27174
rect 24846 27163 25154 27172
rect 36188 26994 36216 29294
rect 36726 29294 37228 29322
rect 36726 29200 36782 29294
rect 37200 27554 37228 29294
rect 37370 29200 37426 30000
rect 38014 29200 38070 30000
rect 38658 29322 38714 30000
rect 38658 29294 38792 29322
rect 38658 29200 38714 29294
rect 37384 27606 37412 29200
rect 38028 27606 38056 29200
rect 37280 27600 37332 27606
rect 37200 27548 37280 27554
rect 37200 27542 37332 27548
rect 37372 27600 37424 27606
rect 37372 27542 37424 27548
rect 38016 27600 38068 27606
rect 38016 27542 38068 27548
rect 37200 27526 37320 27542
rect 36794 27228 37102 27237
rect 36794 27226 36800 27228
rect 36856 27226 36880 27228
rect 36936 27226 36960 27228
rect 37016 27226 37040 27228
rect 37096 27226 37102 27228
rect 36856 27174 36858 27226
rect 37038 27174 37040 27226
rect 36794 27172 36800 27174
rect 36856 27172 36880 27174
rect 36936 27172 36960 27174
rect 37016 27172 37040 27174
rect 37096 27172 37102 27174
rect 36794 27163 37102 27172
rect 38764 26994 38792 29294
rect 39302 29200 39358 30000
rect 39946 29200 40002 30000
rect 40590 29322 40646 30000
rect 41234 29322 41290 30000
rect 40590 29294 40724 29322
rect 40590 29200 40646 29294
rect 39960 27554 39988 29200
rect 40040 27600 40092 27606
rect 39960 27548 40040 27554
rect 39960 27542 40092 27548
rect 39960 27526 40080 27542
rect 40696 27538 40724 29294
rect 41234 29294 41368 29322
rect 41234 29200 41290 29294
rect 41340 27606 41368 29294
rect 41878 29200 41934 30000
rect 42522 29322 42578 30000
rect 42522 29294 42656 29322
rect 42522 29200 42578 29294
rect 41328 27600 41380 27606
rect 41328 27542 41380 27548
rect 40684 27532 40736 27538
rect 40684 27474 40736 27480
rect 41892 26994 41920 29200
rect 42628 27538 42656 29294
rect 43166 29200 43222 30000
rect 43810 29322 43866 30000
rect 43810 29294 43944 29322
rect 43810 29200 43866 29294
rect 42768 27772 43076 27781
rect 42768 27770 42774 27772
rect 42830 27770 42854 27772
rect 42910 27770 42934 27772
rect 42990 27770 43014 27772
rect 43070 27770 43076 27772
rect 42830 27718 42832 27770
rect 43012 27718 43014 27770
rect 42768 27716 42774 27718
rect 42830 27716 42854 27718
rect 42910 27716 42934 27718
rect 42990 27716 43014 27718
rect 43070 27716 43076 27718
rect 42768 27707 43076 27716
rect 43180 27606 43208 29200
rect 43168 27600 43220 27606
rect 43168 27542 43220 27548
rect 42616 27532 42668 27538
rect 42616 27474 42668 27480
rect 43916 26994 43944 29294
rect 44454 29200 44510 30000
rect 45098 29322 45154 30000
rect 45742 29322 45798 30000
rect 46386 29322 46442 30000
rect 45098 29294 45232 29322
rect 45098 29200 45154 29294
rect 45204 27606 45232 29294
rect 45742 29294 45876 29322
rect 45742 29200 45798 29294
rect 45742 28248 45798 28257
rect 45742 28183 45798 28192
rect 45192 27600 45244 27606
rect 45192 27542 45244 27548
rect 45756 26994 45784 28183
rect 45848 27606 45876 29294
rect 46386 29294 46520 29322
rect 46386 29200 46442 29294
rect 46492 27606 46520 29294
rect 47030 29200 47086 30000
rect 47674 29200 47730 30000
rect 48318 29200 48374 30000
rect 48962 29200 49018 30000
rect 49606 29200 49662 30000
rect 45836 27600 45888 27606
rect 45836 27542 45888 27548
rect 46480 27600 46532 27606
rect 46480 27542 46532 27548
rect 47044 27130 47072 29200
rect 47490 27704 47546 27713
rect 47490 27639 47546 27648
rect 47400 27464 47452 27470
rect 47400 27406 47452 27412
rect 47032 27124 47084 27130
rect 47032 27066 47084 27072
rect 36176 26988 36228 26994
rect 36176 26930 36228 26936
rect 38752 26988 38804 26994
rect 38752 26930 38804 26936
rect 41880 26988 41932 26994
rect 41880 26930 41932 26936
rect 43904 26988 43956 26994
rect 43904 26930 43956 26936
rect 45744 26988 45796 26994
rect 45744 26930 45796 26936
rect 46846 26888 46902 26897
rect 46846 26823 46902 26832
rect 30820 26684 31128 26693
rect 30820 26682 30826 26684
rect 30882 26682 30906 26684
rect 30962 26682 30986 26684
rect 31042 26682 31066 26684
rect 31122 26682 31128 26684
rect 30882 26630 30884 26682
rect 31064 26630 31066 26682
rect 30820 26628 30826 26630
rect 30882 26628 30906 26630
rect 30962 26628 30986 26630
rect 31042 26628 31066 26630
rect 31122 26628 31128 26630
rect 30820 26619 31128 26628
rect 42768 26684 43076 26693
rect 42768 26682 42774 26684
rect 42830 26682 42854 26684
rect 42910 26682 42934 26684
rect 42990 26682 43014 26684
rect 43070 26682 43076 26684
rect 42830 26630 42832 26682
rect 43012 26630 43014 26682
rect 42768 26628 42774 26630
rect 42830 26628 42854 26630
rect 42910 26628 42934 26630
rect 42990 26628 43014 26630
rect 43070 26628 43076 26630
rect 42768 26619 43076 26628
rect 46860 26450 46888 26823
rect 46848 26444 46900 26450
rect 46848 26386 46900 26392
rect 24846 26140 25154 26149
rect 24846 26138 24852 26140
rect 24908 26138 24932 26140
rect 24988 26138 25012 26140
rect 25068 26138 25092 26140
rect 25148 26138 25154 26140
rect 24908 26086 24910 26138
rect 25090 26086 25092 26138
rect 24846 26084 24852 26086
rect 24908 26084 24932 26086
rect 24988 26084 25012 26086
rect 25068 26084 25092 26086
rect 25148 26084 25154 26086
rect 24846 26075 25154 26084
rect 36794 26140 37102 26149
rect 36794 26138 36800 26140
rect 36856 26138 36880 26140
rect 36936 26138 36960 26140
rect 37016 26138 37040 26140
rect 37096 26138 37102 26140
rect 36856 26086 36858 26138
rect 37038 26086 37040 26138
rect 36794 26084 36800 26086
rect 36856 26084 36880 26086
rect 36936 26084 36960 26086
rect 37016 26084 37040 26086
rect 37096 26084 37102 26086
rect 36794 26075 37102 26084
rect 30820 25596 31128 25605
rect 30820 25594 30826 25596
rect 30882 25594 30906 25596
rect 30962 25594 30986 25596
rect 31042 25594 31066 25596
rect 31122 25594 31128 25596
rect 30882 25542 30884 25594
rect 31064 25542 31066 25594
rect 30820 25540 30826 25542
rect 30882 25540 30906 25542
rect 30962 25540 30986 25542
rect 31042 25540 31066 25542
rect 31122 25540 31128 25542
rect 30820 25531 31128 25540
rect 42768 25596 43076 25605
rect 42768 25594 42774 25596
rect 42830 25594 42854 25596
rect 42910 25594 42934 25596
rect 42990 25594 43014 25596
rect 43070 25594 43076 25596
rect 42830 25542 42832 25594
rect 43012 25542 43014 25594
rect 42768 25540 42774 25542
rect 42830 25540 42854 25542
rect 42910 25540 42934 25542
rect 42990 25540 43014 25542
rect 43070 25540 43076 25542
rect 42768 25531 43076 25540
rect 24846 25052 25154 25061
rect 24846 25050 24852 25052
rect 24908 25050 24932 25052
rect 24988 25050 25012 25052
rect 25068 25050 25092 25052
rect 25148 25050 25154 25052
rect 24908 24998 24910 25050
rect 25090 24998 25092 25050
rect 24846 24996 24852 24998
rect 24908 24996 24932 24998
rect 24988 24996 25012 24998
rect 25068 24996 25092 24998
rect 25148 24996 25154 24998
rect 24846 24987 25154 24996
rect 36794 25052 37102 25061
rect 36794 25050 36800 25052
rect 36856 25050 36880 25052
rect 36936 25050 36960 25052
rect 37016 25050 37040 25052
rect 37096 25050 37102 25052
rect 36856 24998 36858 25050
rect 37038 24998 37040 25050
rect 36794 24996 36800 24998
rect 36856 24996 36880 24998
rect 36936 24996 36960 24998
rect 37016 24996 37040 24998
rect 37096 24996 37102 24998
rect 36794 24987 37102 24996
rect 30820 24508 31128 24517
rect 30820 24506 30826 24508
rect 30882 24506 30906 24508
rect 30962 24506 30986 24508
rect 31042 24506 31066 24508
rect 31122 24506 31128 24508
rect 30882 24454 30884 24506
rect 31064 24454 31066 24506
rect 30820 24452 30826 24454
rect 30882 24452 30906 24454
rect 30962 24452 30986 24454
rect 31042 24452 31066 24454
rect 31122 24452 31128 24454
rect 30820 24443 31128 24452
rect 42768 24508 43076 24517
rect 42768 24506 42774 24508
rect 42830 24506 42854 24508
rect 42910 24506 42934 24508
rect 42990 24506 43014 24508
rect 43070 24506 43076 24508
rect 42830 24454 42832 24506
rect 43012 24454 43014 24506
rect 42768 24452 42774 24454
rect 42830 24452 42854 24454
rect 42910 24452 42934 24454
rect 42990 24452 43014 24454
rect 43070 24452 43076 24454
rect 42768 24443 43076 24452
rect 24846 23964 25154 23973
rect 24846 23962 24852 23964
rect 24908 23962 24932 23964
rect 24988 23962 25012 23964
rect 25068 23962 25092 23964
rect 25148 23962 25154 23964
rect 24908 23910 24910 23962
rect 25090 23910 25092 23962
rect 24846 23908 24852 23910
rect 24908 23908 24932 23910
rect 24988 23908 25012 23910
rect 25068 23908 25092 23910
rect 25148 23908 25154 23910
rect 24846 23899 25154 23908
rect 36794 23964 37102 23973
rect 36794 23962 36800 23964
rect 36856 23962 36880 23964
rect 36936 23962 36960 23964
rect 37016 23962 37040 23964
rect 37096 23962 37102 23964
rect 36856 23910 36858 23962
rect 37038 23910 37040 23962
rect 36794 23908 36800 23910
rect 36856 23908 36880 23910
rect 36936 23908 36960 23910
rect 37016 23908 37040 23910
rect 37096 23908 37102 23910
rect 36794 23899 37102 23908
rect 30820 23420 31128 23429
rect 30820 23418 30826 23420
rect 30882 23418 30906 23420
rect 30962 23418 30986 23420
rect 31042 23418 31066 23420
rect 31122 23418 31128 23420
rect 30882 23366 30884 23418
rect 31064 23366 31066 23418
rect 30820 23364 30826 23366
rect 30882 23364 30906 23366
rect 30962 23364 30986 23366
rect 31042 23364 31066 23366
rect 31122 23364 31128 23366
rect 30820 23355 31128 23364
rect 42768 23420 43076 23429
rect 42768 23418 42774 23420
rect 42830 23418 42854 23420
rect 42910 23418 42934 23420
rect 42990 23418 43014 23420
rect 43070 23418 43076 23420
rect 42830 23366 42832 23418
rect 43012 23366 43014 23418
rect 42768 23364 42774 23366
rect 42830 23364 42854 23366
rect 42910 23364 42934 23366
rect 42990 23364 43014 23366
rect 43070 23364 43076 23366
rect 42768 23355 43076 23364
rect 24846 22876 25154 22885
rect 24846 22874 24852 22876
rect 24908 22874 24932 22876
rect 24988 22874 25012 22876
rect 25068 22874 25092 22876
rect 25148 22874 25154 22876
rect 24908 22822 24910 22874
rect 25090 22822 25092 22874
rect 24846 22820 24852 22822
rect 24908 22820 24932 22822
rect 24988 22820 25012 22822
rect 25068 22820 25092 22822
rect 25148 22820 25154 22822
rect 24846 22811 25154 22820
rect 36794 22876 37102 22885
rect 36794 22874 36800 22876
rect 36856 22874 36880 22876
rect 36936 22874 36960 22876
rect 37016 22874 37040 22876
rect 37096 22874 37102 22876
rect 36856 22822 36858 22874
rect 37038 22822 37040 22874
rect 36794 22820 36800 22822
rect 36856 22820 36880 22822
rect 36936 22820 36960 22822
rect 37016 22820 37040 22822
rect 37096 22820 37102 22822
rect 36794 22811 37102 22820
rect 30820 22332 31128 22341
rect 30820 22330 30826 22332
rect 30882 22330 30906 22332
rect 30962 22330 30986 22332
rect 31042 22330 31066 22332
rect 31122 22330 31128 22332
rect 30882 22278 30884 22330
rect 31064 22278 31066 22330
rect 30820 22276 30826 22278
rect 30882 22276 30906 22278
rect 30962 22276 30986 22278
rect 31042 22276 31066 22278
rect 31122 22276 31128 22278
rect 30820 22267 31128 22276
rect 42768 22332 43076 22341
rect 42768 22330 42774 22332
rect 42830 22330 42854 22332
rect 42910 22330 42934 22332
rect 42990 22330 43014 22332
rect 43070 22330 43076 22332
rect 42830 22278 42832 22330
rect 43012 22278 43014 22330
rect 42768 22276 42774 22278
rect 42830 22276 42854 22278
rect 42910 22276 42934 22278
rect 42990 22276 43014 22278
rect 43070 22276 43076 22278
rect 42768 22267 43076 22276
rect 24846 21788 25154 21797
rect 24846 21786 24852 21788
rect 24908 21786 24932 21788
rect 24988 21786 25012 21788
rect 25068 21786 25092 21788
rect 25148 21786 25154 21788
rect 24908 21734 24910 21786
rect 25090 21734 25092 21786
rect 24846 21732 24852 21734
rect 24908 21732 24932 21734
rect 24988 21732 25012 21734
rect 25068 21732 25092 21734
rect 25148 21732 25154 21734
rect 24846 21723 25154 21732
rect 36794 21788 37102 21797
rect 36794 21786 36800 21788
rect 36856 21786 36880 21788
rect 36936 21786 36960 21788
rect 37016 21786 37040 21788
rect 37096 21786 37102 21788
rect 36856 21734 36858 21786
rect 37038 21734 37040 21786
rect 36794 21732 36800 21734
rect 36856 21732 36880 21734
rect 36936 21732 36960 21734
rect 37016 21732 37040 21734
rect 37096 21732 37102 21734
rect 36794 21723 37102 21732
rect 30820 21244 31128 21253
rect 30820 21242 30826 21244
rect 30882 21242 30906 21244
rect 30962 21242 30986 21244
rect 31042 21242 31066 21244
rect 31122 21242 31128 21244
rect 30882 21190 30884 21242
rect 31064 21190 31066 21242
rect 30820 21188 30826 21190
rect 30882 21188 30906 21190
rect 30962 21188 30986 21190
rect 31042 21188 31066 21190
rect 31122 21188 31128 21190
rect 30820 21179 31128 21188
rect 42768 21244 43076 21253
rect 42768 21242 42774 21244
rect 42830 21242 42854 21244
rect 42910 21242 42934 21244
rect 42990 21242 43014 21244
rect 43070 21242 43076 21244
rect 42830 21190 42832 21242
rect 43012 21190 43014 21242
rect 42768 21188 42774 21190
rect 42830 21188 42854 21190
rect 42910 21188 42934 21190
rect 42990 21188 43014 21190
rect 43070 21188 43076 21190
rect 42768 21179 43076 21188
rect 24846 20700 25154 20709
rect 24846 20698 24852 20700
rect 24908 20698 24932 20700
rect 24988 20698 25012 20700
rect 25068 20698 25092 20700
rect 25148 20698 25154 20700
rect 24908 20646 24910 20698
rect 25090 20646 25092 20698
rect 24846 20644 24852 20646
rect 24908 20644 24932 20646
rect 24988 20644 25012 20646
rect 25068 20644 25092 20646
rect 25148 20644 25154 20646
rect 24846 20635 25154 20644
rect 36794 20700 37102 20709
rect 36794 20698 36800 20700
rect 36856 20698 36880 20700
rect 36936 20698 36960 20700
rect 37016 20698 37040 20700
rect 37096 20698 37102 20700
rect 36856 20646 36858 20698
rect 37038 20646 37040 20698
rect 36794 20644 36800 20646
rect 36856 20644 36880 20646
rect 36936 20644 36960 20646
rect 37016 20644 37040 20646
rect 37096 20644 37102 20646
rect 36794 20635 37102 20644
rect 30820 20156 31128 20165
rect 30820 20154 30826 20156
rect 30882 20154 30906 20156
rect 30962 20154 30986 20156
rect 31042 20154 31066 20156
rect 31122 20154 31128 20156
rect 30882 20102 30884 20154
rect 31064 20102 31066 20154
rect 30820 20100 30826 20102
rect 30882 20100 30906 20102
rect 30962 20100 30986 20102
rect 31042 20100 31066 20102
rect 31122 20100 31128 20102
rect 30820 20091 31128 20100
rect 42768 20156 43076 20165
rect 42768 20154 42774 20156
rect 42830 20154 42854 20156
rect 42910 20154 42934 20156
rect 42990 20154 43014 20156
rect 43070 20154 43076 20156
rect 42830 20102 42832 20154
rect 43012 20102 43014 20154
rect 42768 20100 42774 20102
rect 42830 20100 42854 20102
rect 42910 20100 42934 20102
rect 42990 20100 43014 20102
rect 43070 20100 43076 20102
rect 42768 20091 43076 20100
rect 24846 19612 25154 19621
rect 24846 19610 24852 19612
rect 24908 19610 24932 19612
rect 24988 19610 25012 19612
rect 25068 19610 25092 19612
rect 25148 19610 25154 19612
rect 24908 19558 24910 19610
rect 25090 19558 25092 19610
rect 24846 19556 24852 19558
rect 24908 19556 24932 19558
rect 24988 19556 25012 19558
rect 25068 19556 25092 19558
rect 25148 19556 25154 19558
rect 24846 19547 25154 19556
rect 36794 19612 37102 19621
rect 36794 19610 36800 19612
rect 36856 19610 36880 19612
rect 36936 19610 36960 19612
rect 37016 19610 37040 19612
rect 37096 19610 37102 19612
rect 36856 19558 36858 19610
rect 37038 19558 37040 19610
rect 36794 19556 36800 19558
rect 36856 19556 36880 19558
rect 36936 19556 36960 19558
rect 37016 19556 37040 19558
rect 37096 19556 37102 19558
rect 36794 19547 37102 19556
rect 30820 19068 31128 19077
rect 30820 19066 30826 19068
rect 30882 19066 30906 19068
rect 30962 19066 30986 19068
rect 31042 19066 31066 19068
rect 31122 19066 31128 19068
rect 30882 19014 30884 19066
rect 31064 19014 31066 19066
rect 30820 19012 30826 19014
rect 30882 19012 30906 19014
rect 30962 19012 30986 19014
rect 31042 19012 31066 19014
rect 31122 19012 31128 19014
rect 30820 19003 31128 19012
rect 42768 19068 43076 19077
rect 42768 19066 42774 19068
rect 42830 19066 42854 19068
rect 42910 19066 42934 19068
rect 42990 19066 43014 19068
rect 43070 19066 43076 19068
rect 42830 19014 42832 19066
rect 43012 19014 43014 19066
rect 42768 19012 42774 19014
rect 42830 19012 42854 19014
rect 42910 19012 42934 19014
rect 42990 19012 43014 19014
rect 43070 19012 43076 19014
rect 42768 19003 43076 19012
rect 24846 18524 25154 18533
rect 24846 18522 24852 18524
rect 24908 18522 24932 18524
rect 24988 18522 25012 18524
rect 25068 18522 25092 18524
rect 25148 18522 25154 18524
rect 24908 18470 24910 18522
rect 25090 18470 25092 18522
rect 24846 18468 24852 18470
rect 24908 18468 24932 18470
rect 24988 18468 25012 18470
rect 25068 18468 25092 18470
rect 25148 18468 25154 18470
rect 24846 18459 25154 18468
rect 36794 18524 37102 18533
rect 36794 18522 36800 18524
rect 36856 18522 36880 18524
rect 36936 18522 36960 18524
rect 37016 18522 37040 18524
rect 37096 18522 37102 18524
rect 36856 18470 36858 18522
rect 37038 18470 37040 18522
rect 36794 18468 36800 18470
rect 36856 18468 36880 18470
rect 36936 18468 36960 18470
rect 37016 18468 37040 18470
rect 37096 18468 37102 18470
rect 36794 18459 37102 18468
rect 30820 17980 31128 17989
rect 30820 17978 30826 17980
rect 30882 17978 30906 17980
rect 30962 17978 30986 17980
rect 31042 17978 31066 17980
rect 31122 17978 31128 17980
rect 30882 17926 30884 17978
rect 31064 17926 31066 17978
rect 30820 17924 30826 17926
rect 30882 17924 30906 17926
rect 30962 17924 30986 17926
rect 31042 17924 31066 17926
rect 31122 17924 31128 17926
rect 30820 17915 31128 17924
rect 42768 17980 43076 17989
rect 42768 17978 42774 17980
rect 42830 17978 42854 17980
rect 42910 17978 42934 17980
rect 42990 17978 43014 17980
rect 43070 17978 43076 17980
rect 42830 17926 42832 17978
rect 43012 17926 43014 17978
rect 42768 17924 42774 17926
rect 42830 17924 42854 17926
rect 42910 17924 42934 17926
rect 42990 17924 43014 17926
rect 43070 17924 43076 17926
rect 42768 17915 43076 17924
rect 24846 17436 25154 17445
rect 24846 17434 24852 17436
rect 24908 17434 24932 17436
rect 24988 17434 25012 17436
rect 25068 17434 25092 17436
rect 25148 17434 25154 17436
rect 24908 17382 24910 17434
rect 25090 17382 25092 17434
rect 24846 17380 24852 17382
rect 24908 17380 24932 17382
rect 24988 17380 25012 17382
rect 25068 17380 25092 17382
rect 25148 17380 25154 17382
rect 24846 17371 25154 17380
rect 36794 17436 37102 17445
rect 36794 17434 36800 17436
rect 36856 17434 36880 17436
rect 36936 17434 36960 17436
rect 37016 17434 37040 17436
rect 37096 17434 37102 17436
rect 36856 17382 36858 17434
rect 37038 17382 37040 17434
rect 36794 17380 36800 17382
rect 36856 17380 36880 17382
rect 36936 17380 36960 17382
rect 37016 17380 37040 17382
rect 37096 17380 37102 17382
rect 36794 17371 37102 17380
rect 30820 16892 31128 16901
rect 30820 16890 30826 16892
rect 30882 16890 30906 16892
rect 30962 16890 30986 16892
rect 31042 16890 31066 16892
rect 31122 16890 31128 16892
rect 30882 16838 30884 16890
rect 31064 16838 31066 16890
rect 30820 16836 30826 16838
rect 30882 16836 30906 16838
rect 30962 16836 30986 16838
rect 31042 16836 31066 16838
rect 31122 16836 31128 16838
rect 30820 16827 31128 16836
rect 42768 16892 43076 16901
rect 42768 16890 42774 16892
rect 42830 16890 42854 16892
rect 42910 16890 42934 16892
rect 42990 16890 43014 16892
rect 43070 16890 43076 16892
rect 42830 16838 42832 16890
rect 43012 16838 43014 16890
rect 42768 16836 42774 16838
rect 42830 16836 42854 16838
rect 42910 16836 42934 16838
rect 42990 16836 43014 16838
rect 43070 16836 43076 16838
rect 42768 16827 43076 16836
rect 24846 16348 25154 16357
rect 24846 16346 24852 16348
rect 24908 16346 24932 16348
rect 24988 16346 25012 16348
rect 25068 16346 25092 16348
rect 25148 16346 25154 16348
rect 24908 16294 24910 16346
rect 25090 16294 25092 16346
rect 24846 16292 24852 16294
rect 24908 16292 24932 16294
rect 24988 16292 25012 16294
rect 25068 16292 25092 16294
rect 25148 16292 25154 16294
rect 24846 16283 25154 16292
rect 36794 16348 37102 16357
rect 36794 16346 36800 16348
rect 36856 16346 36880 16348
rect 36936 16346 36960 16348
rect 37016 16346 37040 16348
rect 37096 16346 37102 16348
rect 36856 16294 36858 16346
rect 37038 16294 37040 16346
rect 36794 16292 36800 16294
rect 36856 16292 36880 16294
rect 36936 16292 36960 16294
rect 37016 16292 37040 16294
rect 37096 16292 37102 16294
rect 36794 16283 37102 16292
rect 30820 15804 31128 15813
rect 30820 15802 30826 15804
rect 30882 15802 30906 15804
rect 30962 15802 30986 15804
rect 31042 15802 31066 15804
rect 31122 15802 31128 15804
rect 30882 15750 30884 15802
rect 31064 15750 31066 15802
rect 30820 15748 30826 15750
rect 30882 15748 30906 15750
rect 30962 15748 30986 15750
rect 31042 15748 31066 15750
rect 31122 15748 31128 15750
rect 30820 15739 31128 15748
rect 42768 15804 43076 15813
rect 42768 15802 42774 15804
rect 42830 15802 42854 15804
rect 42910 15802 42934 15804
rect 42990 15802 43014 15804
rect 43070 15802 43076 15804
rect 42830 15750 42832 15802
rect 43012 15750 43014 15802
rect 42768 15748 42774 15750
rect 42830 15748 42854 15750
rect 42910 15748 42934 15750
rect 42990 15748 43014 15750
rect 43070 15748 43076 15750
rect 42768 15739 43076 15748
rect 24846 15260 25154 15269
rect 24846 15258 24852 15260
rect 24908 15258 24932 15260
rect 24988 15258 25012 15260
rect 25068 15258 25092 15260
rect 25148 15258 25154 15260
rect 24908 15206 24910 15258
rect 25090 15206 25092 15258
rect 24846 15204 24852 15206
rect 24908 15204 24932 15206
rect 24988 15204 25012 15206
rect 25068 15204 25092 15206
rect 25148 15204 25154 15206
rect 24846 15195 25154 15204
rect 36794 15260 37102 15269
rect 36794 15258 36800 15260
rect 36856 15258 36880 15260
rect 36936 15258 36960 15260
rect 37016 15258 37040 15260
rect 37096 15258 37102 15260
rect 36856 15206 36858 15258
rect 37038 15206 37040 15258
rect 36794 15204 36800 15206
rect 36856 15204 36880 15206
rect 36936 15204 36960 15206
rect 37016 15204 37040 15206
rect 37096 15204 37102 15206
rect 36794 15195 37102 15204
rect 1398 14991 1454 15000
rect 22928 15020 22980 15026
rect 22928 14962 22980 14968
rect 22928 14816 22980 14822
rect 22928 14758 22980 14764
rect 6924 14716 7232 14725
rect 6924 14714 6930 14716
rect 6986 14714 7010 14716
rect 7066 14714 7090 14716
rect 7146 14714 7170 14716
rect 7226 14714 7232 14716
rect 6986 14662 6988 14714
rect 7168 14662 7170 14714
rect 6924 14660 6930 14662
rect 6986 14660 7010 14662
rect 7066 14660 7090 14662
rect 7146 14660 7170 14662
rect 7226 14660 7232 14662
rect 6924 14651 7232 14660
rect 18872 14716 19180 14725
rect 18872 14714 18878 14716
rect 18934 14714 18958 14716
rect 19014 14714 19038 14716
rect 19094 14714 19118 14716
rect 19174 14714 19180 14716
rect 18934 14662 18936 14714
rect 19116 14662 19118 14714
rect 18872 14660 18878 14662
rect 18934 14660 18958 14662
rect 19014 14660 19038 14662
rect 19094 14660 19118 14662
rect 19174 14660 19180 14662
rect 18872 14651 19180 14660
rect 1400 14408 1452 14414
rect 1398 14376 1400 14385
rect 1452 14376 1454 14385
rect 1398 14311 1454 14320
rect 12898 14172 13206 14181
rect 12898 14170 12904 14172
rect 12960 14170 12984 14172
rect 13040 14170 13064 14172
rect 13120 14170 13144 14172
rect 13200 14170 13206 14172
rect 12960 14118 12962 14170
rect 13142 14118 13144 14170
rect 12898 14116 12904 14118
rect 12960 14116 12984 14118
rect 13040 14116 13064 14118
rect 13120 14116 13144 14118
rect 13200 14116 13206 14118
rect 12898 14107 13206 14116
rect 1400 13728 1452 13734
rect 1398 13696 1400 13705
rect 1452 13696 1454 13705
rect 1398 13631 1454 13640
rect 6924 13628 7232 13637
rect 6924 13626 6930 13628
rect 6986 13626 7010 13628
rect 7066 13626 7090 13628
rect 7146 13626 7170 13628
rect 7226 13626 7232 13628
rect 6986 13574 6988 13626
rect 7168 13574 7170 13626
rect 6924 13572 6930 13574
rect 6986 13572 7010 13574
rect 7066 13572 7090 13574
rect 7146 13572 7170 13574
rect 7226 13572 7232 13574
rect 6924 13563 7232 13572
rect 18872 13628 19180 13637
rect 18872 13626 18878 13628
rect 18934 13626 18958 13628
rect 19014 13626 19038 13628
rect 19094 13626 19118 13628
rect 19174 13626 19180 13628
rect 18934 13574 18936 13626
rect 19116 13574 19118 13626
rect 18872 13572 18878 13574
rect 18934 13572 18958 13574
rect 19014 13572 19038 13574
rect 19094 13572 19118 13574
rect 19174 13572 19180 13574
rect 18872 13563 19180 13572
rect 22192 13184 22244 13190
rect 22192 13126 22244 13132
rect 12898 13084 13206 13093
rect 12898 13082 12904 13084
rect 12960 13082 12984 13084
rect 13040 13082 13064 13084
rect 13120 13082 13144 13084
rect 13200 13082 13206 13084
rect 12960 13030 12962 13082
rect 13142 13030 13144 13082
rect 12898 13028 12904 13030
rect 12960 13028 12984 13030
rect 13040 13028 13064 13030
rect 13120 13028 13144 13030
rect 13200 13028 13206 13030
rect 12898 13019 13206 13028
rect 1400 12640 1452 12646
rect 1400 12582 1452 12588
rect 1412 12345 1440 12582
rect 6924 12540 7232 12549
rect 6924 12538 6930 12540
rect 6986 12538 7010 12540
rect 7066 12538 7090 12540
rect 7146 12538 7170 12540
rect 7226 12538 7232 12540
rect 6986 12486 6988 12538
rect 7168 12486 7170 12538
rect 6924 12484 6930 12486
rect 6986 12484 7010 12486
rect 7066 12484 7090 12486
rect 7146 12484 7170 12486
rect 7226 12484 7232 12486
rect 6924 12475 7232 12484
rect 18872 12540 19180 12549
rect 18872 12538 18878 12540
rect 18934 12538 18958 12540
rect 19014 12538 19038 12540
rect 19094 12538 19118 12540
rect 19174 12538 19180 12540
rect 18934 12486 18936 12538
rect 19116 12486 19118 12538
rect 18872 12484 18878 12486
rect 18934 12484 18958 12486
rect 19014 12484 19038 12486
rect 19094 12484 19118 12486
rect 19174 12484 19180 12486
rect 18872 12475 19180 12484
rect 1398 12336 1454 12345
rect 1398 12271 1454 12280
rect 12898 11996 13206 12005
rect 12898 11994 12904 11996
rect 12960 11994 12984 11996
rect 13040 11994 13064 11996
rect 13120 11994 13144 11996
rect 13200 11994 13206 11996
rect 12960 11942 12962 11994
rect 13142 11942 13144 11994
rect 12898 11940 12904 11942
rect 12960 11940 12984 11942
rect 13040 11940 13064 11942
rect 13120 11940 13144 11942
rect 13200 11940 13206 11942
rect 12898 11931 13206 11940
rect 1400 11688 1452 11694
rect 1398 11656 1400 11665
rect 1452 11656 1454 11665
rect 1398 11591 1454 11600
rect 6924 11452 7232 11461
rect 6924 11450 6930 11452
rect 6986 11450 7010 11452
rect 7066 11450 7090 11452
rect 7146 11450 7170 11452
rect 7226 11450 7232 11452
rect 6986 11398 6988 11450
rect 7168 11398 7170 11450
rect 6924 11396 6930 11398
rect 6986 11396 7010 11398
rect 7066 11396 7090 11398
rect 7146 11396 7170 11398
rect 7226 11396 7232 11398
rect 6924 11387 7232 11396
rect 18872 11452 19180 11461
rect 18872 11450 18878 11452
rect 18934 11450 18958 11452
rect 19014 11450 19038 11452
rect 19094 11450 19118 11452
rect 19174 11450 19180 11452
rect 18934 11398 18936 11450
rect 19116 11398 19118 11450
rect 18872 11396 18878 11398
rect 18934 11396 18958 11398
rect 19014 11396 19038 11398
rect 19094 11396 19118 11398
rect 19174 11396 19180 11398
rect 18872 11387 19180 11396
rect 1400 11076 1452 11082
rect 1400 11018 1452 11024
rect 1412 10985 1440 11018
rect 1398 10976 1454 10985
rect 1398 10911 1454 10920
rect 12898 10908 13206 10917
rect 12898 10906 12904 10908
rect 12960 10906 12984 10908
rect 13040 10906 13064 10908
rect 13120 10906 13144 10908
rect 13200 10906 13206 10908
rect 12960 10854 12962 10906
rect 13142 10854 13144 10906
rect 12898 10852 12904 10854
rect 12960 10852 12984 10854
rect 13040 10852 13064 10854
rect 13120 10852 13144 10854
rect 13200 10852 13206 10854
rect 12898 10843 13206 10852
rect 6924 10364 7232 10373
rect 6924 10362 6930 10364
rect 6986 10362 7010 10364
rect 7066 10362 7090 10364
rect 7146 10362 7170 10364
rect 7226 10362 7232 10364
rect 6986 10310 6988 10362
rect 7168 10310 7170 10362
rect 6924 10308 6930 10310
rect 6986 10308 7010 10310
rect 7066 10308 7090 10310
rect 7146 10308 7170 10310
rect 7226 10308 7232 10310
rect 6924 10299 7232 10308
rect 18872 10364 19180 10373
rect 18872 10362 18878 10364
rect 18934 10362 18958 10364
rect 19014 10362 19038 10364
rect 19094 10362 19118 10364
rect 19174 10362 19180 10364
rect 18934 10310 18936 10362
rect 19116 10310 19118 10362
rect 18872 10308 18878 10310
rect 18934 10308 18958 10310
rect 19014 10308 19038 10310
rect 19094 10308 19118 10310
rect 19174 10308 19180 10310
rect 18872 10299 19180 10308
rect 12898 9820 13206 9829
rect 12898 9818 12904 9820
rect 12960 9818 12984 9820
rect 13040 9818 13064 9820
rect 13120 9818 13144 9820
rect 13200 9818 13206 9820
rect 12960 9766 12962 9818
rect 13142 9766 13144 9818
rect 12898 9764 12904 9766
rect 12960 9764 12984 9766
rect 13040 9764 13064 9766
rect 13120 9764 13144 9766
rect 13200 9764 13206 9766
rect 12898 9755 13206 9764
rect 6924 9276 7232 9285
rect 6924 9274 6930 9276
rect 6986 9274 7010 9276
rect 7066 9274 7090 9276
rect 7146 9274 7170 9276
rect 7226 9274 7232 9276
rect 6986 9222 6988 9274
rect 7168 9222 7170 9274
rect 6924 9220 6930 9222
rect 6986 9220 7010 9222
rect 7066 9220 7090 9222
rect 7146 9220 7170 9222
rect 7226 9220 7232 9222
rect 6924 9211 7232 9220
rect 18872 9276 19180 9285
rect 18872 9274 18878 9276
rect 18934 9274 18958 9276
rect 19014 9274 19038 9276
rect 19094 9274 19118 9276
rect 19174 9274 19180 9276
rect 18934 9222 18936 9274
rect 19116 9222 19118 9274
rect 18872 9220 18878 9222
rect 18934 9220 18958 9222
rect 19014 9220 19038 9222
rect 19094 9220 19118 9222
rect 19174 9220 19180 9222
rect 18872 9211 19180 9220
rect 1400 8968 1452 8974
rect 1398 8936 1400 8945
rect 1452 8936 1454 8945
rect 1398 8871 1454 8880
rect 12898 8732 13206 8741
rect 12898 8730 12904 8732
rect 12960 8730 12984 8732
rect 13040 8730 13064 8732
rect 13120 8730 13144 8732
rect 13200 8730 13206 8732
rect 12960 8678 12962 8730
rect 13142 8678 13144 8730
rect 12898 8676 12904 8678
rect 12960 8676 12984 8678
rect 13040 8676 13064 8678
rect 13120 8676 13144 8678
rect 13200 8676 13206 8678
rect 12898 8667 13206 8676
rect 1400 8356 1452 8362
rect 1400 8298 1452 8304
rect 1412 8265 1440 8298
rect 1398 8256 1454 8265
rect 1398 8191 1454 8200
rect 6924 8188 7232 8197
rect 6924 8186 6930 8188
rect 6986 8186 7010 8188
rect 7066 8186 7090 8188
rect 7146 8186 7170 8188
rect 7226 8186 7232 8188
rect 6986 8134 6988 8186
rect 7168 8134 7170 8186
rect 6924 8132 6930 8134
rect 6986 8132 7010 8134
rect 7066 8132 7090 8134
rect 7146 8132 7170 8134
rect 7226 8132 7232 8134
rect 6924 8123 7232 8132
rect 18872 8188 19180 8197
rect 18872 8186 18878 8188
rect 18934 8186 18958 8188
rect 19014 8186 19038 8188
rect 19094 8186 19118 8188
rect 19174 8186 19180 8188
rect 18934 8134 18936 8186
rect 19116 8134 19118 8186
rect 18872 8132 18878 8134
rect 18934 8132 18958 8134
rect 19014 8132 19038 8134
rect 19094 8132 19118 8134
rect 19174 8132 19180 8134
rect 18872 8123 19180 8132
rect 1400 7744 1452 7750
rect 1400 7686 1452 7692
rect 1412 7585 1440 7686
rect 12898 7644 13206 7653
rect 12898 7642 12904 7644
rect 12960 7642 12984 7644
rect 13040 7642 13064 7644
rect 13120 7642 13144 7644
rect 13200 7642 13206 7644
rect 12960 7590 12962 7642
rect 13142 7590 13144 7642
rect 12898 7588 12904 7590
rect 12960 7588 12984 7590
rect 13040 7588 13064 7590
rect 13120 7588 13144 7590
rect 13200 7588 13206 7590
rect 1398 7576 1454 7585
rect 12898 7579 13206 7588
rect 1398 7511 1454 7520
rect 1400 7336 1452 7342
rect 1400 7278 1452 7284
rect 1412 6905 1440 7278
rect 6924 7100 7232 7109
rect 6924 7098 6930 7100
rect 6986 7098 7010 7100
rect 7066 7098 7090 7100
rect 7146 7098 7170 7100
rect 7226 7098 7232 7100
rect 6986 7046 6988 7098
rect 7168 7046 7170 7098
rect 6924 7044 6930 7046
rect 6986 7044 7010 7046
rect 7066 7044 7090 7046
rect 7146 7044 7170 7046
rect 7226 7044 7232 7046
rect 6924 7035 7232 7044
rect 18872 7100 19180 7109
rect 18872 7098 18878 7100
rect 18934 7098 18958 7100
rect 19014 7098 19038 7100
rect 19094 7098 19118 7100
rect 19174 7098 19180 7100
rect 18934 7046 18936 7098
rect 19116 7046 19118 7098
rect 18872 7044 18878 7046
rect 18934 7044 18958 7046
rect 19014 7044 19038 7046
rect 19094 7044 19118 7046
rect 19174 7044 19180 7046
rect 18872 7035 19180 7044
rect 1398 6896 1454 6905
rect 1398 6831 1454 6840
rect 12898 6556 13206 6565
rect 12898 6554 12904 6556
rect 12960 6554 12984 6556
rect 13040 6554 13064 6556
rect 13120 6554 13144 6556
rect 13200 6554 13206 6556
rect 12960 6502 12962 6554
rect 13142 6502 13144 6554
rect 12898 6500 12904 6502
rect 12960 6500 12984 6502
rect 13040 6500 13064 6502
rect 13120 6500 13144 6502
rect 13200 6500 13206 6502
rect 12898 6491 13206 6500
rect 1400 6248 1452 6254
rect 1398 6216 1400 6225
rect 1452 6216 1454 6225
rect 1398 6151 1454 6160
rect 6924 6012 7232 6021
rect 6924 6010 6930 6012
rect 6986 6010 7010 6012
rect 7066 6010 7090 6012
rect 7146 6010 7170 6012
rect 7226 6010 7232 6012
rect 6986 5958 6988 6010
rect 7168 5958 7170 6010
rect 6924 5956 6930 5958
rect 6986 5956 7010 5958
rect 7066 5956 7090 5958
rect 7146 5956 7170 5958
rect 7226 5956 7232 5958
rect 6924 5947 7232 5956
rect 18872 6012 19180 6021
rect 18872 6010 18878 6012
rect 18934 6010 18958 6012
rect 19014 6010 19038 6012
rect 19094 6010 19118 6012
rect 19174 6010 19180 6012
rect 18934 5958 18936 6010
rect 19116 5958 19118 6010
rect 18872 5956 18878 5958
rect 18934 5956 18958 5958
rect 19014 5956 19038 5958
rect 19094 5956 19118 5958
rect 19174 5956 19180 5958
rect 18872 5947 19180 5956
rect 1400 5704 1452 5710
rect 1400 5646 1452 5652
rect 1412 5545 1440 5646
rect 1398 5536 1454 5545
rect 1398 5471 1454 5480
rect 12898 5468 13206 5477
rect 12898 5466 12904 5468
rect 12960 5466 12984 5468
rect 13040 5466 13064 5468
rect 13120 5466 13144 5468
rect 13200 5466 13206 5468
rect 12960 5414 12962 5466
rect 13142 5414 13144 5466
rect 12898 5412 12904 5414
rect 12960 5412 12984 5414
rect 13040 5412 13064 5414
rect 13120 5412 13144 5414
rect 13200 5412 13206 5414
rect 12898 5403 13206 5412
rect 1400 5024 1452 5030
rect 1400 4966 1452 4972
rect 1412 4865 1440 4966
rect 6924 4924 7232 4933
rect 6924 4922 6930 4924
rect 6986 4922 7010 4924
rect 7066 4922 7090 4924
rect 7146 4922 7170 4924
rect 7226 4922 7232 4924
rect 6986 4870 6988 4922
rect 7168 4870 7170 4922
rect 6924 4868 6930 4870
rect 6986 4868 7010 4870
rect 7066 4868 7090 4870
rect 7146 4868 7170 4870
rect 7226 4868 7232 4870
rect 1398 4856 1454 4865
rect 6924 4859 7232 4868
rect 18872 4924 19180 4933
rect 18872 4922 18878 4924
rect 18934 4922 18958 4924
rect 19014 4922 19038 4924
rect 19094 4922 19118 4924
rect 19174 4922 19180 4924
rect 18934 4870 18936 4922
rect 19116 4870 19118 4922
rect 18872 4868 18878 4870
rect 18934 4868 18958 4870
rect 19014 4868 19038 4870
rect 19094 4868 19118 4870
rect 19174 4868 19180 4870
rect 18872 4859 19180 4868
rect 1398 4791 1454 4800
rect 12898 4380 13206 4389
rect 12898 4378 12904 4380
rect 12960 4378 12984 4380
rect 13040 4378 13064 4380
rect 13120 4378 13144 4380
rect 13200 4378 13206 4380
rect 12960 4326 12962 4378
rect 13142 4326 13144 4378
rect 12898 4324 12904 4326
rect 12960 4324 12984 4326
rect 13040 4324 13064 4326
rect 13120 4324 13144 4326
rect 13200 4324 13206 4326
rect 12898 4315 13206 4324
rect 2872 3936 2924 3942
rect 2872 3878 2924 3884
rect 2780 3596 2832 3602
rect 2780 3538 2832 3544
rect 1400 3528 1452 3534
rect 1398 3496 1400 3505
rect 1452 3496 1454 3505
rect 1398 3431 1454 3440
rect 20 2916 72 2922
rect 20 2858 72 2864
rect 32 800 60 2858
rect 664 2848 716 2854
rect 664 2790 716 2796
rect 676 800 704 2790
rect 1308 2440 1360 2446
rect 1308 2382 1360 2388
rect 2596 2440 2648 2446
rect 2596 2382 2648 2388
rect 1320 800 1348 2382
rect 2608 800 2636 2382
rect 2792 2145 2820 3538
rect 2778 2136 2834 2145
rect 2778 2071 2834 2080
rect 2884 1465 2912 3878
rect 6924 3836 7232 3845
rect 6924 3834 6930 3836
rect 6986 3834 7010 3836
rect 7066 3834 7090 3836
rect 7146 3834 7170 3836
rect 7226 3834 7232 3836
rect 6986 3782 6988 3834
rect 7168 3782 7170 3834
rect 6924 3780 6930 3782
rect 6986 3780 7010 3782
rect 7066 3780 7090 3782
rect 7146 3780 7170 3782
rect 7226 3780 7232 3782
rect 6924 3771 7232 3780
rect 18872 3836 19180 3845
rect 18872 3834 18878 3836
rect 18934 3834 18958 3836
rect 19014 3834 19038 3836
rect 19094 3834 19118 3836
rect 19174 3834 19180 3836
rect 18934 3782 18936 3834
rect 19116 3782 19118 3834
rect 18872 3780 18878 3782
rect 18934 3780 18958 3782
rect 19014 3780 19038 3782
rect 19094 3780 19118 3782
rect 19174 3780 19180 3782
rect 18872 3771 19180 3780
rect 2964 3528 3016 3534
rect 2964 3470 3016 3476
rect 2870 1456 2926 1465
rect 2870 1391 2926 1400
rect 18 0 74 800
rect 662 0 718 800
rect 1306 0 1362 800
rect 1950 0 2006 800
rect 2594 0 2650 800
rect 2976 785 3004 3470
rect 12898 3292 13206 3301
rect 12898 3290 12904 3292
rect 12960 3290 12984 3292
rect 13040 3290 13064 3292
rect 13120 3290 13144 3292
rect 13200 3290 13206 3292
rect 12960 3238 12962 3290
rect 13142 3238 13144 3290
rect 12898 3236 12904 3238
rect 12960 3236 12984 3238
rect 13040 3236 13064 3238
rect 13120 3236 13144 3238
rect 13200 3236 13206 3238
rect 12898 3227 13206 3236
rect 3056 2984 3108 2990
rect 3056 2926 3108 2932
rect 3884 2984 3936 2990
rect 3884 2926 3936 2932
rect 2962 776 3018 785
rect 2962 711 3018 720
rect 2962 96 3018 105
rect 3068 82 3096 2926
rect 3240 2440 3292 2446
rect 3240 2382 3292 2388
rect 3252 800 3280 2382
rect 3896 800 3924 2926
rect 9036 2848 9088 2854
rect 9036 2790 9088 2796
rect 16764 2848 16816 2854
rect 16764 2790 16816 2796
rect 19340 2848 19392 2854
rect 19340 2790 19392 2796
rect 6924 2748 7232 2757
rect 6924 2746 6930 2748
rect 6986 2746 7010 2748
rect 7066 2746 7090 2748
rect 7146 2746 7170 2748
rect 7226 2746 7232 2748
rect 6986 2694 6988 2746
rect 7168 2694 7170 2746
rect 6924 2692 6930 2694
rect 6986 2692 7010 2694
rect 7066 2692 7090 2694
rect 7146 2692 7170 2694
rect 7226 2692 7232 2694
rect 6924 2683 7232 2692
rect 5172 2440 5224 2446
rect 5172 2382 5224 2388
rect 5816 2440 5868 2446
rect 5816 2382 5868 2388
rect 7104 2440 7156 2446
rect 7104 2382 7156 2388
rect 7748 2440 7800 2446
rect 7748 2382 7800 2388
rect 8392 2440 8444 2446
rect 8392 2382 8444 2388
rect 4528 2304 4580 2310
rect 4528 2246 4580 2252
rect 4540 800 4568 2246
rect 5184 800 5212 2382
rect 5828 800 5856 2382
rect 7116 800 7144 2382
rect 7760 800 7788 2382
rect 8404 800 8432 2382
rect 9048 800 9076 2790
rect 10324 2440 10376 2446
rect 10324 2382 10376 2388
rect 10968 2440 11020 2446
rect 10968 2382 11020 2388
rect 12808 2440 12860 2446
rect 12808 2382 12860 2388
rect 13544 2440 13596 2446
rect 13544 2382 13596 2388
rect 14832 2440 14884 2446
rect 14832 2382 14884 2388
rect 9680 2304 9732 2310
rect 9680 2246 9732 2252
rect 9692 800 9720 2246
rect 10336 800 10364 2382
rect 10980 800 11008 2382
rect 11612 2304 11664 2310
rect 11612 2246 11664 2252
rect 12256 2304 12308 2310
rect 12256 2246 12308 2252
rect 11624 800 11652 2246
rect 12268 800 12296 2246
rect 12820 1306 12848 2382
rect 12898 2204 13206 2213
rect 12898 2202 12904 2204
rect 12960 2202 12984 2204
rect 13040 2202 13064 2204
rect 13120 2202 13144 2204
rect 13200 2202 13206 2204
rect 12960 2150 12962 2202
rect 13142 2150 13144 2202
rect 12898 2148 12904 2150
rect 12960 2148 12984 2150
rect 13040 2148 13064 2150
rect 13120 2148 13144 2150
rect 13200 2148 13206 2150
rect 12898 2139 13206 2148
rect 12820 1278 12940 1306
rect 12912 800 12940 1278
rect 13556 800 13584 2382
rect 14844 800 14872 2382
rect 16120 2304 16172 2310
rect 16120 2246 16172 2252
rect 16132 800 16160 2246
rect 16776 800 16804 2790
rect 18872 2748 19180 2757
rect 18872 2746 18878 2748
rect 18934 2746 18958 2748
rect 19014 2746 19038 2748
rect 19094 2746 19118 2748
rect 19174 2746 19180 2748
rect 18934 2694 18936 2746
rect 19116 2694 19118 2746
rect 18872 2692 18878 2694
rect 18934 2692 18958 2694
rect 19014 2692 19038 2694
rect 19094 2692 19118 2694
rect 19174 2692 19180 2694
rect 18872 2683 19180 2692
rect 17408 2440 17460 2446
rect 17408 2382 17460 2388
rect 18052 2440 18104 2446
rect 18052 2382 18104 2388
rect 18696 2440 18748 2446
rect 18696 2382 18748 2388
rect 17420 800 17448 2382
rect 18064 800 18092 2382
rect 18708 800 18736 2382
rect 19352 800 19380 2790
rect 22204 2446 22232 13126
rect 22940 2446 22968 14758
rect 30820 14716 31128 14725
rect 30820 14714 30826 14716
rect 30882 14714 30906 14716
rect 30962 14714 30986 14716
rect 31042 14714 31066 14716
rect 31122 14714 31128 14716
rect 30882 14662 30884 14714
rect 31064 14662 31066 14714
rect 30820 14660 30826 14662
rect 30882 14660 30906 14662
rect 30962 14660 30986 14662
rect 31042 14660 31066 14662
rect 31122 14660 31128 14662
rect 30820 14651 31128 14660
rect 42768 14716 43076 14725
rect 42768 14714 42774 14716
rect 42830 14714 42854 14716
rect 42910 14714 42934 14716
rect 42990 14714 43014 14716
rect 43070 14714 43076 14716
rect 42830 14662 42832 14714
rect 43012 14662 43014 14714
rect 42768 14660 42774 14662
rect 42830 14660 42854 14662
rect 42910 14660 42934 14662
rect 42990 14660 43014 14662
rect 43070 14660 43076 14662
rect 42768 14651 43076 14660
rect 38384 14408 38436 14414
rect 38384 14350 38436 14356
rect 39856 14408 39908 14414
rect 39856 14350 39908 14356
rect 25228 14272 25280 14278
rect 25228 14214 25280 14220
rect 24846 14172 25154 14181
rect 24846 14170 24852 14172
rect 24908 14170 24932 14172
rect 24988 14170 25012 14172
rect 25068 14170 25092 14172
rect 25148 14170 25154 14172
rect 24908 14118 24910 14170
rect 25090 14118 25092 14170
rect 24846 14116 24852 14118
rect 24908 14116 24932 14118
rect 24988 14116 25012 14118
rect 25068 14116 25092 14118
rect 25148 14116 25154 14118
rect 24846 14107 25154 14116
rect 25240 14006 25268 14214
rect 36794 14172 37102 14181
rect 36794 14170 36800 14172
rect 36856 14170 36880 14172
rect 36936 14170 36960 14172
rect 37016 14170 37040 14172
rect 37096 14170 37102 14172
rect 36856 14118 36858 14170
rect 37038 14118 37040 14170
rect 36794 14116 36800 14118
rect 36856 14116 36880 14118
rect 36936 14116 36960 14118
rect 37016 14116 37040 14118
rect 37096 14116 37102 14118
rect 36794 14107 37102 14116
rect 25228 14000 25280 14006
rect 25228 13942 25280 13948
rect 30288 14000 30340 14006
rect 30288 13942 30340 13948
rect 26056 13932 26108 13938
rect 26056 13874 26108 13880
rect 24676 13864 24728 13870
rect 24676 13806 24728 13812
rect 24688 13326 24716 13806
rect 24676 13320 24728 13326
rect 24676 13262 24728 13268
rect 24846 13084 25154 13093
rect 24846 13082 24852 13084
rect 24908 13082 24932 13084
rect 24988 13082 25012 13084
rect 25068 13082 25092 13084
rect 25148 13082 25154 13084
rect 24908 13030 24910 13082
rect 25090 13030 25092 13082
rect 24846 13028 24852 13030
rect 24908 13028 24932 13030
rect 24988 13028 25012 13030
rect 25068 13028 25092 13030
rect 25148 13028 25154 13030
rect 24846 13019 25154 13028
rect 26068 12714 26096 13874
rect 29184 13864 29236 13870
rect 29184 13806 29236 13812
rect 26424 13728 26476 13734
rect 26424 13670 26476 13676
rect 27988 13728 28040 13734
rect 27988 13670 28040 13676
rect 26436 13394 26464 13670
rect 28000 13530 28028 13670
rect 27988 13524 28040 13530
rect 27988 13466 28040 13472
rect 26424 13388 26476 13394
rect 26424 13330 26476 13336
rect 29196 12986 29224 13806
rect 29184 12980 29236 12986
rect 29184 12922 29236 12928
rect 30300 12782 30328 13942
rect 32404 13864 32456 13870
rect 32404 13806 32456 13812
rect 30820 13628 31128 13637
rect 30820 13626 30826 13628
rect 30882 13626 30906 13628
rect 30962 13626 30986 13628
rect 31042 13626 31066 13628
rect 31122 13626 31128 13628
rect 30882 13574 30884 13626
rect 31064 13574 31066 13626
rect 30820 13572 30826 13574
rect 30882 13572 30906 13574
rect 30962 13572 30986 13574
rect 31042 13572 31066 13574
rect 31122 13572 31128 13574
rect 30820 13563 31128 13572
rect 32416 13394 32444 13806
rect 33324 13728 33376 13734
rect 33324 13670 33376 13676
rect 32404 13388 32456 13394
rect 32404 13330 32456 13336
rect 33336 12918 33364 13670
rect 38396 13530 38424 14350
rect 39868 13870 39896 14350
rect 45100 14340 45152 14346
rect 45100 14282 45152 14288
rect 43260 14272 43312 14278
rect 43260 14214 43312 14220
rect 43272 14006 43300 14214
rect 43260 14000 43312 14006
rect 43260 13942 43312 13948
rect 39856 13864 39908 13870
rect 39856 13806 39908 13812
rect 38384 13524 38436 13530
rect 38384 13466 38436 13472
rect 34888 13320 34940 13326
rect 34888 13262 34940 13268
rect 33324 12912 33376 12918
rect 33324 12854 33376 12860
rect 30288 12776 30340 12782
rect 30288 12718 30340 12724
rect 26056 12708 26108 12714
rect 26056 12650 26108 12656
rect 34900 12646 34928 13262
rect 36794 13084 37102 13093
rect 36794 13082 36800 13084
rect 36856 13082 36880 13084
rect 36936 13082 36960 13084
rect 37016 13082 37040 13084
rect 37096 13082 37102 13084
rect 36856 13030 36858 13082
rect 37038 13030 37040 13082
rect 36794 13028 36800 13030
rect 36856 13028 36880 13030
rect 36936 13028 36960 13030
rect 37016 13028 37040 13030
rect 37096 13028 37102 13030
rect 36794 13019 37102 13028
rect 39868 12646 39896 13806
rect 42768 13628 43076 13637
rect 42768 13626 42774 13628
rect 42830 13626 42854 13628
rect 42910 13626 42934 13628
rect 42990 13626 43014 13628
rect 43070 13626 43076 13628
rect 42830 13574 42832 13626
rect 43012 13574 43014 13626
rect 42768 13572 42774 13574
rect 42830 13572 42854 13574
rect 42910 13572 42934 13574
rect 42990 13572 43014 13574
rect 43070 13572 43076 13574
rect 42768 13563 43076 13572
rect 45112 12986 45140 14282
rect 45560 14068 45612 14074
rect 45560 14010 45612 14016
rect 45572 13841 45600 14010
rect 46940 13864 46992 13870
rect 45558 13832 45614 13841
rect 46940 13806 46992 13812
rect 45558 13767 45614 13776
rect 46388 13252 46440 13258
rect 46388 13194 46440 13200
rect 46400 12986 46428 13194
rect 45100 12980 45152 12986
rect 45100 12922 45152 12928
rect 46388 12980 46440 12986
rect 46388 12922 46440 12928
rect 46112 12844 46164 12850
rect 46112 12786 46164 12792
rect 34888 12640 34940 12646
rect 34888 12582 34940 12588
rect 39856 12640 39908 12646
rect 39856 12582 39908 12588
rect 30820 12540 31128 12549
rect 30820 12538 30826 12540
rect 30882 12538 30906 12540
rect 30962 12538 30986 12540
rect 31042 12538 31066 12540
rect 31122 12538 31128 12540
rect 30882 12486 30884 12538
rect 31064 12486 31066 12538
rect 30820 12484 30826 12486
rect 30882 12484 30906 12486
rect 30962 12484 30986 12486
rect 31042 12484 31066 12486
rect 31122 12484 31128 12486
rect 30820 12475 31128 12484
rect 42768 12540 43076 12549
rect 42768 12538 42774 12540
rect 42830 12538 42854 12540
rect 42910 12538 42934 12540
rect 42990 12538 43014 12540
rect 43070 12538 43076 12540
rect 42830 12486 42832 12538
rect 43012 12486 43014 12538
rect 42768 12484 42774 12486
rect 42830 12484 42854 12486
rect 42910 12484 42934 12486
rect 42990 12484 43014 12486
rect 43070 12484 43076 12486
rect 42768 12475 43076 12484
rect 24846 11996 25154 12005
rect 24846 11994 24852 11996
rect 24908 11994 24932 11996
rect 24988 11994 25012 11996
rect 25068 11994 25092 11996
rect 25148 11994 25154 11996
rect 24908 11942 24910 11994
rect 25090 11942 25092 11994
rect 24846 11940 24852 11942
rect 24908 11940 24932 11942
rect 24988 11940 25012 11942
rect 25068 11940 25092 11942
rect 25148 11940 25154 11942
rect 24846 11931 25154 11940
rect 36794 11996 37102 12005
rect 36794 11994 36800 11996
rect 36856 11994 36880 11996
rect 36936 11994 36960 11996
rect 37016 11994 37040 11996
rect 37096 11994 37102 11996
rect 36856 11942 36858 11994
rect 37038 11942 37040 11994
rect 36794 11940 36800 11942
rect 36856 11940 36880 11942
rect 36936 11940 36960 11942
rect 37016 11940 37040 11942
rect 37096 11940 37102 11942
rect 36794 11931 37102 11940
rect 30820 11452 31128 11461
rect 30820 11450 30826 11452
rect 30882 11450 30906 11452
rect 30962 11450 30986 11452
rect 31042 11450 31066 11452
rect 31122 11450 31128 11452
rect 30882 11398 30884 11450
rect 31064 11398 31066 11450
rect 30820 11396 30826 11398
rect 30882 11396 30906 11398
rect 30962 11396 30986 11398
rect 31042 11396 31066 11398
rect 31122 11396 31128 11398
rect 30820 11387 31128 11396
rect 42768 11452 43076 11461
rect 42768 11450 42774 11452
rect 42830 11450 42854 11452
rect 42910 11450 42934 11452
rect 42990 11450 43014 11452
rect 43070 11450 43076 11452
rect 42830 11398 42832 11450
rect 43012 11398 43014 11450
rect 42768 11396 42774 11398
rect 42830 11396 42854 11398
rect 42910 11396 42934 11398
rect 42990 11396 43014 11398
rect 43070 11396 43076 11398
rect 42768 11387 43076 11396
rect 24846 10908 25154 10917
rect 24846 10906 24852 10908
rect 24908 10906 24932 10908
rect 24988 10906 25012 10908
rect 25068 10906 25092 10908
rect 25148 10906 25154 10908
rect 24908 10854 24910 10906
rect 25090 10854 25092 10906
rect 24846 10852 24852 10854
rect 24908 10852 24932 10854
rect 24988 10852 25012 10854
rect 25068 10852 25092 10854
rect 25148 10852 25154 10854
rect 24846 10843 25154 10852
rect 36794 10908 37102 10917
rect 36794 10906 36800 10908
rect 36856 10906 36880 10908
rect 36936 10906 36960 10908
rect 37016 10906 37040 10908
rect 37096 10906 37102 10908
rect 36856 10854 36858 10906
rect 37038 10854 37040 10906
rect 36794 10852 36800 10854
rect 36856 10852 36880 10854
rect 36936 10852 36960 10854
rect 37016 10852 37040 10854
rect 37096 10852 37102 10854
rect 36794 10843 37102 10852
rect 30820 10364 31128 10373
rect 30820 10362 30826 10364
rect 30882 10362 30906 10364
rect 30962 10362 30986 10364
rect 31042 10362 31066 10364
rect 31122 10362 31128 10364
rect 30882 10310 30884 10362
rect 31064 10310 31066 10362
rect 30820 10308 30826 10310
rect 30882 10308 30906 10310
rect 30962 10308 30986 10310
rect 31042 10308 31066 10310
rect 31122 10308 31128 10310
rect 30820 10299 31128 10308
rect 42768 10364 43076 10373
rect 42768 10362 42774 10364
rect 42830 10362 42854 10364
rect 42910 10362 42934 10364
rect 42990 10362 43014 10364
rect 43070 10362 43076 10364
rect 42830 10310 42832 10362
rect 43012 10310 43014 10362
rect 42768 10308 42774 10310
rect 42830 10308 42854 10310
rect 42910 10308 42934 10310
rect 42990 10308 43014 10310
rect 43070 10308 43076 10310
rect 42768 10299 43076 10308
rect 24846 9820 25154 9829
rect 24846 9818 24852 9820
rect 24908 9818 24932 9820
rect 24988 9818 25012 9820
rect 25068 9818 25092 9820
rect 25148 9818 25154 9820
rect 24908 9766 24910 9818
rect 25090 9766 25092 9818
rect 24846 9764 24852 9766
rect 24908 9764 24932 9766
rect 24988 9764 25012 9766
rect 25068 9764 25092 9766
rect 25148 9764 25154 9766
rect 24846 9755 25154 9764
rect 36794 9820 37102 9829
rect 36794 9818 36800 9820
rect 36856 9818 36880 9820
rect 36936 9818 36960 9820
rect 37016 9818 37040 9820
rect 37096 9818 37102 9820
rect 36856 9766 36858 9818
rect 37038 9766 37040 9818
rect 36794 9764 36800 9766
rect 36856 9764 36880 9766
rect 36936 9764 36960 9766
rect 37016 9764 37040 9766
rect 37096 9764 37102 9766
rect 36794 9755 37102 9764
rect 45744 9580 45796 9586
rect 45744 9522 45796 9528
rect 30820 9276 31128 9285
rect 30820 9274 30826 9276
rect 30882 9274 30906 9276
rect 30962 9274 30986 9276
rect 31042 9274 31066 9276
rect 31122 9274 31128 9276
rect 30882 9222 30884 9274
rect 31064 9222 31066 9274
rect 30820 9220 30826 9222
rect 30882 9220 30906 9222
rect 30962 9220 30986 9222
rect 31042 9220 31066 9222
rect 31122 9220 31128 9222
rect 30820 9211 31128 9220
rect 42768 9276 43076 9285
rect 42768 9274 42774 9276
rect 42830 9274 42854 9276
rect 42910 9274 42934 9276
rect 42990 9274 43014 9276
rect 43070 9274 43076 9276
rect 42830 9222 42832 9274
rect 43012 9222 43014 9274
rect 42768 9220 42774 9222
rect 42830 9220 42854 9222
rect 42910 9220 42934 9222
rect 42990 9220 43014 9222
rect 43070 9220 43076 9222
rect 42768 9211 43076 9220
rect 24846 8732 25154 8741
rect 24846 8730 24852 8732
rect 24908 8730 24932 8732
rect 24988 8730 25012 8732
rect 25068 8730 25092 8732
rect 25148 8730 25154 8732
rect 24908 8678 24910 8730
rect 25090 8678 25092 8730
rect 24846 8676 24852 8678
rect 24908 8676 24932 8678
rect 24988 8676 25012 8678
rect 25068 8676 25092 8678
rect 25148 8676 25154 8678
rect 24846 8667 25154 8676
rect 36794 8732 37102 8741
rect 36794 8730 36800 8732
rect 36856 8730 36880 8732
rect 36936 8730 36960 8732
rect 37016 8730 37040 8732
rect 37096 8730 37102 8732
rect 36856 8678 36858 8730
rect 37038 8678 37040 8730
rect 36794 8676 36800 8678
rect 36856 8676 36880 8678
rect 36936 8676 36960 8678
rect 37016 8676 37040 8678
rect 37096 8676 37102 8678
rect 36794 8667 37102 8676
rect 30820 8188 31128 8197
rect 30820 8186 30826 8188
rect 30882 8186 30906 8188
rect 30962 8186 30986 8188
rect 31042 8186 31066 8188
rect 31122 8186 31128 8188
rect 30882 8134 30884 8186
rect 31064 8134 31066 8186
rect 30820 8132 30826 8134
rect 30882 8132 30906 8134
rect 30962 8132 30986 8134
rect 31042 8132 31066 8134
rect 31122 8132 31128 8134
rect 30820 8123 31128 8132
rect 42768 8188 43076 8197
rect 42768 8186 42774 8188
rect 42830 8186 42854 8188
rect 42910 8186 42934 8188
rect 42990 8186 43014 8188
rect 43070 8186 43076 8188
rect 42830 8134 42832 8186
rect 43012 8134 43014 8186
rect 42768 8132 42774 8134
rect 42830 8132 42854 8134
rect 42910 8132 42934 8134
rect 42990 8132 43014 8134
rect 43070 8132 43076 8134
rect 42768 8123 43076 8132
rect 24846 7644 25154 7653
rect 24846 7642 24852 7644
rect 24908 7642 24932 7644
rect 24988 7642 25012 7644
rect 25068 7642 25092 7644
rect 25148 7642 25154 7644
rect 24908 7590 24910 7642
rect 25090 7590 25092 7642
rect 24846 7588 24852 7590
rect 24908 7588 24932 7590
rect 24988 7588 25012 7590
rect 25068 7588 25092 7590
rect 25148 7588 25154 7590
rect 24846 7579 25154 7588
rect 36794 7644 37102 7653
rect 36794 7642 36800 7644
rect 36856 7642 36880 7644
rect 36936 7642 36960 7644
rect 37016 7642 37040 7644
rect 37096 7642 37102 7644
rect 36856 7590 36858 7642
rect 37038 7590 37040 7642
rect 36794 7588 36800 7590
rect 36856 7588 36880 7590
rect 36936 7588 36960 7590
rect 37016 7588 37040 7590
rect 37096 7588 37102 7590
rect 36794 7579 37102 7588
rect 30820 7100 31128 7109
rect 30820 7098 30826 7100
rect 30882 7098 30906 7100
rect 30962 7098 30986 7100
rect 31042 7098 31066 7100
rect 31122 7098 31128 7100
rect 30882 7046 30884 7098
rect 31064 7046 31066 7098
rect 30820 7044 30826 7046
rect 30882 7044 30906 7046
rect 30962 7044 30986 7046
rect 31042 7044 31066 7046
rect 31122 7044 31128 7046
rect 30820 7035 31128 7044
rect 42768 7100 43076 7109
rect 42768 7098 42774 7100
rect 42830 7098 42854 7100
rect 42910 7098 42934 7100
rect 42990 7098 43014 7100
rect 43070 7098 43076 7100
rect 42830 7046 42832 7098
rect 43012 7046 43014 7098
rect 42768 7044 42774 7046
rect 42830 7044 42854 7046
rect 42910 7044 42934 7046
rect 42990 7044 43014 7046
rect 43070 7044 43076 7046
rect 42768 7035 43076 7044
rect 24846 6556 25154 6565
rect 24846 6554 24852 6556
rect 24908 6554 24932 6556
rect 24988 6554 25012 6556
rect 25068 6554 25092 6556
rect 25148 6554 25154 6556
rect 24908 6502 24910 6554
rect 25090 6502 25092 6554
rect 24846 6500 24852 6502
rect 24908 6500 24932 6502
rect 24988 6500 25012 6502
rect 25068 6500 25092 6502
rect 25148 6500 25154 6502
rect 24846 6491 25154 6500
rect 36794 6556 37102 6565
rect 36794 6554 36800 6556
rect 36856 6554 36880 6556
rect 36936 6554 36960 6556
rect 37016 6554 37040 6556
rect 37096 6554 37102 6556
rect 36856 6502 36858 6554
rect 37038 6502 37040 6554
rect 36794 6500 36800 6502
rect 36856 6500 36880 6502
rect 36936 6500 36960 6502
rect 37016 6500 37040 6502
rect 37096 6500 37102 6502
rect 36794 6491 37102 6500
rect 30820 6012 31128 6021
rect 30820 6010 30826 6012
rect 30882 6010 30906 6012
rect 30962 6010 30986 6012
rect 31042 6010 31066 6012
rect 31122 6010 31128 6012
rect 30882 5958 30884 6010
rect 31064 5958 31066 6010
rect 30820 5956 30826 5958
rect 30882 5956 30906 5958
rect 30962 5956 30986 5958
rect 31042 5956 31066 5958
rect 31122 5956 31128 5958
rect 30820 5947 31128 5956
rect 42768 6012 43076 6021
rect 42768 6010 42774 6012
rect 42830 6010 42854 6012
rect 42910 6010 42934 6012
rect 42990 6010 43014 6012
rect 43070 6010 43076 6012
rect 42830 5958 42832 6010
rect 43012 5958 43014 6010
rect 42768 5956 42774 5958
rect 42830 5956 42854 5958
rect 42910 5956 42934 5958
rect 42990 5956 43014 5958
rect 43070 5956 43076 5958
rect 42768 5947 43076 5956
rect 24846 5468 25154 5477
rect 24846 5466 24852 5468
rect 24908 5466 24932 5468
rect 24988 5466 25012 5468
rect 25068 5466 25092 5468
rect 25148 5466 25154 5468
rect 24908 5414 24910 5466
rect 25090 5414 25092 5466
rect 24846 5412 24852 5414
rect 24908 5412 24932 5414
rect 24988 5412 25012 5414
rect 25068 5412 25092 5414
rect 25148 5412 25154 5414
rect 24846 5403 25154 5412
rect 36794 5468 37102 5477
rect 36794 5466 36800 5468
rect 36856 5466 36880 5468
rect 36936 5466 36960 5468
rect 37016 5466 37040 5468
rect 37096 5466 37102 5468
rect 36856 5414 36858 5466
rect 37038 5414 37040 5466
rect 36794 5412 36800 5414
rect 36856 5412 36880 5414
rect 36936 5412 36960 5414
rect 37016 5412 37040 5414
rect 37096 5412 37102 5414
rect 36794 5403 37102 5412
rect 30820 4924 31128 4933
rect 30820 4922 30826 4924
rect 30882 4922 30906 4924
rect 30962 4922 30986 4924
rect 31042 4922 31066 4924
rect 31122 4922 31128 4924
rect 30882 4870 30884 4922
rect 31064 4870 31066 4922
rect 30820 4868 30826 4870
rect 30882 4868 30906 4870
rect 30962 4868 30986 4870
rect 31042 4868 31066 4870
rect 31122 4868 31128 4870
rect 30820 4859 31128 4868
rect 42768 4924 43076 4933
rect 42768 4922 42774 4924
rect 42830 4922 42854 4924
rect 42910 4922 42934 4924
rect 42990 4922 43014 4924
rect 43070 4922 43076 4924
rect 42830 4870 42832 4922
rect 43012 4870 43014 4922
rect 42768 4868 42774 4870
rect 42830 4868 42854 4870
rect 42910 4868 42934 4870
rect 42990 4868 43014 4870
rect 43070 4868 43076 4870
rect 42768 4859 43076 4868
rect 24846 4380 25154 4389
rect 24846 4378 24852 4380
rect 24908 4378 24932 4380
rect 24988 4378 25012 4380
rect 25068 4378 25092 4380
rect 25148 4378 25154 4380
rect 24908 4326 24910 4378
rect 25090 4326 25092 4378
rect 24846 4324 24852 4326
rect 24908 4324 24932 4326
rect 24988 4324 25012 4326
rect 25068 4324 25092 4326
rect 25148 4324 25154 4326
rect 24846 4315 25154 4324
rect 36794 4380 37102 4389
rect 36794 4378 36800 4380
rect 36856 4378 36880 4380
rect 36936 4378 36960 4380
rect 37016 4378 37040 4380
rect 37096 4378 37102 4380
rect 36856 4326 36858 4378
rect 37038 4326 37040 4378
rect 36794 4324 36800 4326
rect 36856 4324 36880 4326
rect 36936 4324 36960 4326
rect 37016 4324 37040 4326
rect 37096 4324 37102 4326
rect 36794 4315 37102 4324
rect 30820 3836 31128 3845
rect 30820 3834 30826 3836
rect 30882 3834 30906 3836
rect 30962 3834 30986 3836
rect 31042 3834 31066 3836
rect 31122 3834 31128 3836
rect 30882 3782 30884 3834
rect 31064 3782 31066 3834
rect 30820 3780 30826 3782
rect 30882 3780 30906 3782
rect 30962 3780 30986 3782
rect 31042 3780 31066 3782
rect 31122 3780 31128 3782
rect 30820 3771 31128 3780
rect 42768 3836 43076 3845
rect 42768 3834 42774 3836
rect 42830 3834 42854 3836
rect 42910 3834 42934 3836
rect 42990 3834 43014 3836
rect 43070 3834 43076 3836
rect 42830 3782 42832 3834
rect 43012 3782 43014 3834
rect 42768 3780 42774 3782
rect 42830 3780 42854 3782
rect 42910 3780 42934 3782
rect 42990 3780 43014 3782
rect 43070 3780 43076 3782
rect 42768 3771 43076 3780
rect 24846 3292 25154 3301
rect 24846 3290 24852 3292
rect 24908 3290 24932 3292
rect 24988 3290 25012 3292
rect 25068 3290 25092 3292
rect 25148 3290 25154 3292
rect 24908 3238 24910 3290
rect 25090 3238 25092 3290
rect 24846 3236 24852 3238
rect 24908 3236 24932 3238
rect 24988 3236 25012 3238
rect 25068 3236 25092 3238
rect 25148 3236 25154 3238
rect 24846 3227 25154 3236
rect 36794 3292 37102 3301
rect 36794 3290 36800 3292
rect 36856 3290 36880 3292
rect 36936 3290 36960 3292
rect 37016 3290 37040 3292
rect 37096 3290 37102 3292
rect 36856 3238 36858 3290
rect 37038 3238 37040 3290
rect 36794 3236 36800 3238
rect 36856 3236 36880 3238
rect 36936 3236 36960 3238
rect 37016 3236 37040 3238
rect 37096 3236 37102 3238
rect 36794 3227 37102 3236
rect 45756 3194 45784 9522
rect 46124 9450 46152 12786
rect 46952 11218 46980 13806
rect 47412 11354 47440 27406
rect 47504 26586 47532 27639
rect 47688 26994 47716 29200
rect 48332 27334 48360 29200
rect 48320 27328 48372 27334
rect 48320 27270 48372 27276
rect 47676 26988 47728 26994
rect 47676 26930 47728 26936
rect 48976 26926 49004 29200
rect 48964 26920 49016 26926
rect 48964 26862 49016 26868
rect 47492 26580 47544 26586
rect 47492 26522 47544 26528
rect 48134 26344 48190 26353
rect 48134 26279 48190 26288
rect 48148 25906 48176 26279
rect 48228 26240 48280 26246
rect 48228 26182 48280 26188
rect 48136 25900 48188 25906
rect 48136 25842 48188 25848
rect 48240 25537 48268 26182
rect 49620 25838 49648 29200
rect 49608 25832 49660 25838
rect 49608 25774 49660 25780
rect 48226 25528 48282 25537
rect 48226 25463 48282 25472
rect 48136 25288 48188 25294
rect 48136 25230 48188 25236
rect 48148 24993 48176 25230
rect 48134 24984 48190 24993
rect 48134 24919 48190 24928
rect 48136 24608 48188 24614
rect 48136 24550 48188 24556
rect 48148 23633 48176 24550
rect 48228 24200 48280 24206
rect 48228 24142 48280 24148
rect 48134 23624 48190 23633
rect 48134 23559 48190 23568
rect 48136 23520 48188 23526
rect 48240 23497 48268 24142
rect 48136 23462 48188 23468
rect 48226 23488 48282 23497
rect 48148 22522 48176 23462
rect 48226 23423 48282 23432
rect 48148 22494 48268 22522
rect 48136 22432 48188 22438
rect 48136 22374 48188 22380
rect 48148 22137 48176 22374
rect 48240 22273 48268 22494
rect 48226 22264 48282 22273
rect 48226 22199 48282 22208
rect 48134 22128 48190 22137
rect 48134 22063 48190 22072
rect 48136 22024 48188 22030
rect 48136 21966 48188 21972
rect 48148 20777 48176 21966
rect 48228 20936 48280 20942
rect 48228 20878 48280 20884
rect 48134 20768 48190 20777
rect 48134 20703 48190 20712
rect 48240 19417 48268 20878
rect 48226 19408 48282 19417
rect 48226 19343 48282 19352
rect 48136 19168 48188 19174
rect 48136 19110 48188 19116
rect 48148 18193 48176 19110
rect 48228 18624 48280 18630
rect 48228 18566 48280 18572
rect 48134 18184 48190 18193
rect 48134 18119 48190 18128
rect 48136 18080 48188 18086
rect 48240 18057 48268 18566
rect 48136 18022 48188 18028
rect 48226 18048 48282 18057
rect 48148 17082 48176 18022
rect 48226 17983 48282 17992
rect 48148 17054 48268 17082
rect 48136 16992 48188 16998
rect 48136 16934 48188 16940
rect 48148 16697 48176 16934
rect 48240 16833 48268 17054
rect 48226 16824 48282 16833
rect 48226 16759 48282 16768
rect 48134 16688 48190 16697
rect 48134 16623 48190 16632
rect 48228 16584 48280 16590
rect 48228 16526 48280 16532
rect 48136 15904 48188 15910
rect 48136 15846 48188 15852
rect 48148 15337 48176 15846
rect 48240 15473 48268 16526
rect 48226 15464 48282 15473
rect 48226 15399 48282 15408
rect 48134 15328 48190 15337
rect 48134 15263 48190 15272
rect 48778 15056 48834 15065
rect 48778 14991 48834 15000
rect 48136 14408 48188 14414
rect 48136 14350 48188 14356
rect 47676 14000 47728 14006
rect 48148 13977 48176 14350
rect 47676 13942 47728 13948
rect 48134 13968 48190 13977
rect 47688 12986 47716 13942
rect 48134 13903 48190 13912
rect 48792 13841 48820 14991
rect 48778 13832 48834 13841
rect 48778 13767 48834 13776
rect 48228 13728 48280 13734
rect 48228 13670 48280 13676
rect 48778 13696 48834 13705
rect 48136 13320 48188 13326
rect 48136 13262 48188 13268
rect 47676 12980 47728 12986
rect 47676 12922 47728 12928
rect 48148 12753 48176 13262
rect 48134 12744 48190 12753
rect 48134 12679 48190 12688
rect 48240 12617 48268 13670
rect 48778 13631 48834 13640
rect 48792 12617 48820 13631
rect 48226 12608 48282 12617
rect 48226 12543 48282 12552
rect 48778 12608 48834 12617
rect 48778 12543 48834 12552
rect 48778 12336 48834 12345
rect 48778 12271 48834 12280
rect 48228 12232 48280 12238
rect 48228 12174 48280 12180
rect 48136 11552 48188 11558
rect 48136 11494 48188 11500
rect 48148 11393 48176 11494
rect 48134 11384 48190 11393
rect 47400 11348 47452 11354
rect 48134 11319 48190 11328
rect 47400 11290 47452 11296
rect 48240 11257 48268 12174
rect 48792 11257 48820 12271
rect 48226 11248 48282 11257
rect 46940 11212 46992 11218
rect 46940 11154 46992 11160
rect 47768 11212 47820 11218
rect 48226 11183 48282 11192
rect 48778 11248 48834 11257
rect 48778 11183 48834 11192
rect 47768 11154 47820 11160
rect 47216 11144 47268 11150
rect 47216 11086 47268 11092
rect 47228 10810 47256 11086
rect 47216 10804 47268 10810
rect 47216 10746 47268 10752
rect 47780 10674 47808 11154
rect 47584 10668 47636 10674
rect 47584 10610 47636 10616
rect 47768 10668 47820 10674
rect 47768 10610 47820 10616
rect 47596 9586 47624 10610
rect 47780 9674 47808 10610
rect 48136 10056 48188 10062
rect 48136 9998 48188 10004
rect 48148 9674 48176 9998
rect 47780 9646 47992 9674
rect 48148 9646 48268 9674
rect 47584 9580 47636 9586
rect 47584 9522 47636 9528
rect 46112 9444 46164 9450
rect 46112 9386 46164 9392
rect 47964 8090 47992 9646
rect 48136 8968 48188 8974
rect 48136 8910 48188 8916
rect 48148 8673 48176 8910
rect 48134 8664 48190 8673
rect 48134 8599 48190 8608
rect 48240 8537 48268 9646
rect 48778 9616 48834 9625
rect 48778 9551 48834 9560
rect 48792 8537 48820 9551
rect 48226 8528 48282 8537
rect 48226 8463 48282 8472
rect 48778 8528 48834 8537
rect 48778 8463 48834 8472
rect 47952 8084 48004 8090
rect 47952 8026 48004 8032
rect 48136 7880 48188 7886
rect 48136 7822 48188 7828
rect 48148 7177 48176 7822
rect 48228 7336 48280 7342
rect 48228 7278 48280 7284
rect 48134 7168 48190 7177
rect 48134 7103 48190 7112
rect 48136 6112 48188 6118
rect 48136 6054 48188 6060
rect 48148 5953 48176 6054
rect 48134 5944 48190 5953
rect 48134 5879 48190 5888
rect 48240 5817 48268 7278
rect 48778 6896 48834 6905
rect 48778 6831 48834 6840
rect 48792 5817 48820 6831
rect 48226 5808 48282 5817
rect 48226 5743 48282 5752
rect 48778 5808 48834 5817
rect 48778 5743 48834 5752
rect 48228 5024 48280 5030
rect 48228 4966 48280 4972
rect 48136 4616 48188 4622
rect 48136 4558 48188 4564
rect 48148 4185 48176 4558
rect 48240 4457 48268 4966
rect 48226 4448 48282 4457
rect 48226 4383 48282 4392
rect 48134 4176 48190 4185
rect 48134 4111 48190 4120
rect 47768 3936 47820 3942
rect 47768 3878 47820 3884
rect 48964 3936 49016 3942
rect 48964 3878 49016 3884
rect 46664 3528 46716 3534
rect 46664 3470 46716 3476
rect 45744 3188 45796 3194
rect 45744 3130 45796 3136
rect 45560 3052 45612 3058
rect 45560 2994 45612 3000
rect 30748 2984 30800 2990
rect 30748 2926 30800 2932
rect 36084 2984 36136 2990
rect 36084 2926 36136 2932
rect 23204 2848 23256 2854
rect 23204 2790 23256 2796
rect 28356 2848 28408 2854
rect 28356 2790 28408 2796
rect 19984 2440 20036 2446
rect 19984 2382 20036 2388
rect 20628 2440 20680 2446
rect 20628 2382 20680 2388
rect 22192 2440 22244 2446
rect 22192 2382 22244 2388
rect 22928 2440 22980 2446
rect 22928 2382 22980 2388
rect 19996 800 20024 2382
rect 20640 800 20668 2382
rect 21272 2304 21324 2310
rect 21272 2246 21324 2252
rect 21916 2304 21968 2310
rect 21916 2246 21968 2252
rect 22560 2304 22612 2310
rect 22560 2246 22612 2252
rect 21284 800 21312 2246
rect 21928 800 21956 2246
rect 22572 800 22600 2246
rect 23216 800 23244 2790
rect 23848 2440 23900 2446
rect 23848 2382 23900 2388
rect 24492 2440 24544 2446
rect 24492 2382 24544 2388
rect 25228 2440 25280 2446
rect 25228 2382 25280 2388
rect 25780 2440 25832 2446
rect 25780 2382 25832 2388
rect 26424 2440 26476 2446
rect 26424 2382 26476 2388
rect 23860 800 23888 2382
rect 24504 800 24532 2382
rect 24846 2204 25154 2213
rect 24846 2202 24852 2204
rect 24908 2202 24932 2204
rect 24988 2202 25012 2204
rect 25068 2202 25092 2204
rect 25148 2202 25154 2204
rect 24908 2150 24910 2202
rect 25090 2150 25092 2202
rect 24846 2148 24852 2150
rect 24908 2148 24932 2150
rect 24988 2148 25012 2150
rect 25068 2148 25092 2150
rect 25148 2148 25154 2150
rect 24846 2139 25154 2148
rect 25240 1306 25268 2382
rect 25148 1278 25268 1306
rect 25148 800 25176 1278
rect 25792 800 25820 2382
rect 26436 800 26464 2382
rect 27068 2304 27120 2310
rect 27068 2246 27120 2252
rect 27712 2304 27764 2310
rect 27712 2246 27764 2252
rect 27080 800 27108 2246
rect 27724 800 27752 2246
rect 28368 800 28396 2790
rect 29000 2440 29052 2446
rect 29000 2382 29052 2388
rect 29644 2440 29696 2446
rect 29644 2382 29696 2388
rect 30288 2440 30340 2446
rect 30288 2382 30340 2388
rect 29012 800 29040 2382
rect 29656 800 29684 2382
rect 30300 800 30328 2382
rect 30760 1578 30788 2926
rect 30820 2748 31128 2757
rect 30820 2746 30826 2748
rect 30882 2746 30906 2748
rect 30962 2746 30986 2748
rect 31042 2746 31066 2748
rect 31122 2746 31128 2748
rect 30882 2694 30884 2746
rect 31064 2694 31066 2746
rect 30820 2692 30826 2694
rect 30882 2692 30906 2694
rect 30962 2692 30986 2694
rect 31042 2692 31066 2694
rect 31122 2692 31128 2694
rect 30820 2683 31128 2692
rect 33508 2440 33560 2446
rect 33508 2382 33560 2388
rect 34152 2440 34204 2446
rect 34152 2382 34204 2388
rect 34796 2440 34848 2446
rect 34796 2382 34848 2388
rect 32220 2304 32272 2310
rect 32220 2246 32272 2252
rect 32864 2304 32916 2310
rect 32864 2246 32916 2252
rect 30760 1550 30972 1578
rect 30944 800 30972 1550
rect 32232 800 32260 2246
rect 32876 800 32904 2246
rect 33520 800 33548 2382
rect 34164 800 34192 2382
rect 34808 800 34836 2382
rect 35440 2304 35492 2310
rect 35440 2246 35492 2252
rect 35452 800 35480 2246
rect 36096 800 36124 2926
rect 43812 2848 43864 2854
rect 43812 2790 43864 2796
rect 42768 2748 43076 2757
rect 42768 2746 42774 2748
rect 42830 2746 42854 2748
rect 42910 2746 42934 2748
rect 42990 2746 43014 2748
rect 43070 2746 43076 2748
rect 42830 2694 42832 2746
rect 43012 2694 43014 2746
rect 42768 2692 42774 2694
rect 42830 2692 42854 2694
rect 42910 2692 42934 2694
rect 42990 2692 43014 2694
rect 43070 2692 43076 2694
rect 42768 2683 43076 2692
rect 37372 2440 37424 2446
rect 37372 2382 37424 2388
rect 38660 2440 38712 2446
rect 38660 2382 38712 2388
rect 39304 2440 39356 2446
rect 39304 2382 39356 2388
rect 40592 2440 40644 2446
rect 40592 2382 40644 2388
rect 41236 2440 41288 2446
rect 41236 2382 41288 2388
rect 42524 2440 42576 2446
rect 42524 2382 42576 2388
rect 36794 2204 37102 2213
rect 36794 2202 36800 2204
rect 36856 2202 36880 2204
rect 36936 2202 36960 2204
rect 37016 2202 37040 2204
rect 37096 2202 37102 2204
rect 36856 2150 36858 2202
rect 37038 2150 37040 2202
rect 36794 2148 36800 2150
rect 36856 2148 36880 2150
rect 36936 2148 36960 2150
rect 37016 2148 37040 2150
rect 37096 2148 37102 2150
rect 36794 2139 37102 2148
rect 37384 800 37412 2382
rect 38672 800 38700 2382
rect 39316 800 39344 2382
rect 40604 800 40632 2382
rect 41248 800 41276 2382
rect 41880 2304 41932 2310
rect 41880 2246 41932 2252
rect 41892 800 41920 2246
rect 42536 800 42564 2382
rect 43168 2304 43220 2310
rect 43168 2246 43220 2252
rect 43180 800 43208 2246
rect 43824 800 43852 2790
rect 44456 2304 44508 2310
rect 44456 2246 44508 2252
rect 45100 2304 45152 2310
rect 45100 2246 45152 2252
rect 44468 800 44496 2246
rect 45112 800 45140 2246
rect 45572 1737 45600 2994
rect 46388 2440 46440 2446
rect 46388 2382 46440 2388
rect 45558 1728 45614 1737
rect 45558 1663 45614 1672
rect 46400 800 46428 2382
rect 3018 54 3096 82
rect 2962 31 3018 40
rect 3238 0 3294 800
rect 3882 0 3938 800
rect 4526 0 4582 800
rect 5170 0 5226 800
rect 5814 0 5870 800
rect 6458 0 6514 800
rect 7102 0 7158 800
rect 7746 0 7802 800
rect 8390 0 8446 800
rect 9034 0 9090 800
rect 9678 0 9734 800
rect 10322 0 10378 800
rect 10966 0 11022 800
rect 11610 0 11666 800
rect 12254 0 12310 800
rect 12898 0 12954 800
rect 13542 0 13598 800
rect 14186 0 14242 800
rect 14830 0 14886 800
rect 15474 0 15530 800
rect 16118 0 16174 800
rect 16762 0 16818 800
rect 17406 0 17462 800
rect 18050 0 18106 800
rect 18694 0 18750 800
rect 19338 0 19394 800
rect 19982 0 20038 800
rect 20626 0 20682 800
rect 21270 0 21326 800
rect 21914 0 21970 800
rect 22558 0 22614 800
rect 23202 0 23258 800
rect 23846 0 23902 800
rect 24490 0 24546 800
rect 25134 0 25190 800
rect 25778 0 25834 800
rect 26422 0 26478 800
rect 27066 0 27122 800
rect 27710 0 27766 800
rect 28354 0 28410 800
rect 28998 0 29054 800
rect 29642 0 29698 800
rect 30286 0 30342 800
rect 30930 0 30986 800
rect 31574 0 31630 800
rect 32218 0 32274 800
rect 32862 0 32918 800
rect 33506 0 33562 800
rect 34150 0 34206 800
rect 34794 0 34850 800
rect 35438 0 35494 800
rect 36082 0 36138 800
rect 36726 0 36782 800
rect 37370 0 37426 800
rect 38014 0 38070 800
rect 38658 0 38714 800
rect 39302 0 39358 800
rect 39946 0 40002 800
rect 40590 0 40646 800
rect 41234 0 41290 800
rect 41878 0 41934 800
rect 42522 0 42578 800
rect 43166 0 43222 800
rect 43810 0 43866 800
rect 44454 0 44510 800
rect 45098 0 45154 800
rect 45742 0 45798 800
rect 46386 0 46442 800
rect 46676 105 46704 3470
rect 46848 2984 46900 2990
rect 46848 2926 46900 2932
rect 47676 2984 47728 2990
rect 47676 2926 47728 2932
rect 46756 2848 46808 2854
rect 46860 2825 46888 2926
rect 46756 2790 46808 2796
rect 46846 2816 46902 2825
rect 46768 377 46796 2790
rect 46846 2751 46902 2760
rect 47032 2440 47084 2446
rect 47032 2382 47084 2388
rect 47044 800 47072 2382
rect 47688 800 47716 2926
rect 47780 1465 47808 3878
rect 48136 3528 48188 3534
rect 48136 3470 48188 3476
rect 48148 3097 48176 3470
rect 48134 3088 48190 3097
rect 48134 3023 48190 3032
rect 47766 1456 47822 1465
rect 47766 1391 47822 1400
rect 48976 800 49004 3878
rect 49608 3392 49660 3398
rect 49608 3334 49660 3340
rect 49620 800 49648 3334
rect 46754 368 46810 377
rect 46754 303 46810 312
rect 46662 96 46718 105
rect 46662 31 46718 40
rect 47030 0 47086 800
rect 47674 0 47730 800
rect 48318 0 48374 800
rect 48962 0 49018 800
rect 49606 0 49662 800
<< via2 >>
rect 1398 27920 1454 27976
rect 2870 29280 2926 29336
rect 2778 28600 2834 28656
rect 1490 27240 1546 27296
rect 1398 25880 1454 25936
rect 6930 27770 6986 27772
rect 7010 27770 7066 27772
rect 7090 27770 7146 27772
rect 7170 27770 7226 27772
rect 6930 27718 6976 27770
rect 6976 27718 6986 27770
rect 7010 27718 7040 27770
rect 7040 27718 7052 27770
rect 7052 27718 7066 27770
rect 7090 27718 7104 27770
rect 7104 27718 7116 27770
rect 7116 27718 7146 27770
rect 7170 27718 7180 27770
rect 7180 27718 7226 27770
rect 6930 27716 6986 27718
rect 7010 27716 7066 27718
rect 7090 27716 7146 27718
rect 7170 27716 7226 27718
rect 18878 27770 18934 27772
rect 18958 27770 19014 27772
rect 19038 27770 19094 27772
rect 19118 27770 19174 27772
rect 18878 27718 18924 27770
rect 18924 27718 18934 27770
rect 18958 27718 18988 27770
rect 18988 27718 19000 27770
rect 19000 27718 19014 27770
rect 19038 27718 19052 27770
rect 19052 27718 19064 27770
rect 19064 27718 19094 27770
rect 19118 27718 19128 27770
rect 19128 27718 19174 27770
rect 18878 27716 18934 27718
rect 18958 27716 19014 27718
rect 19038 27716 19094 27718
rect 19118 27716 19174 27718
rect 12904 27226 12960 27228
rect 12984 27226 13040 27228
rect 13064 27226 13120 27228
rect 13144 27226 13200 27228
rect 12904 27174 12950 27226
rect 12950 27174 12960 27226
rect 12984 27174 13014 27226
rect 13014 27174 13026 27226
rect 13026 27174 13040 27226
rect 13064 27174 13078 27226
rect 13078 27174 13090 27226
rect 13090 27174 13120 27226
rect 13144 27174 13154 27226
rect 13154 27174 13200 27226
rect 12904 27172 12960 27174
rect 12984 27172 13040 27174
rect 13064 27172 13120 27174
rect 13144 27172 13200 27174
rect 30826 27770 30882 27772
rect 30906 27770 30962 27772
rect 30986 27770 31042 27772
rect 31066 27770 31122 27772
rect 30826 27718 30872 27770
rect 30872 27718 30882 27770
rect 30906 27718 30936 27770
rect 30936 27718 30948 27770
rect 30948 27718 30962 27770
rect 30986 27718 31000 27770
rect 31000 27718 31012 27770
rect 31012 27718 31042 27770
rect 31066 27718 31076 27770
rect 31076 27718 31122 27770
rect 30826 27716 30882 27718
rect 30906 27716 30962 27718
rect 30986 27716 31042 27718
rect 31066 27716 31122 27718
rect 6930 26682 6986 26684
rect 7010 26682 7066 26684
rect 7090 26682 7146 26684
rect 7170 26682 7226 26684
rect 6930 26630 6976 26682
rect 6976 26630 6986 26682
rect 7010 26630 7040 26682
rect 7040 26630 7052 26682
rect 7052 26630 7066 26682
rect 7090 26630 7104 26682
rect 7104 26630 7116 26682
rect 7116 26630 7146 26682
rect 7170 26630 7180 26682
rect 7180 26630 7226 26682
rect 6930 26628 6986 26630
rect 7010 26628 7066 26630
rect 7090 26628 7146 26630
rect 7170 26628 7226 26630
rect 18878 26682 18934 26684
rect 18958 26682 19014 26684
rect 19038 26682 19094 26684
rect 19118 26682 19174 26684
rect 18878 26630 18924 26682
rect 18924 26630 18934 26682
rect 18958 26630 18988 26682
rect 18988 26630 19000 26682
rect 19000 26630 19014 26682
rect 19038 26630 19052 26682
rect 19052 26630 19064 26682
rect 19064 26630 19094 26682
rect 19118 26630 19128 26682
rect 19128 26630 19174 26682
rect 18878 26628 18934 26630
rect 18958 26628 19014 26630
rect 19038 26628 19094 26630
rect 19118 26628 19174 26630
rect 12904 26138 12960 26140
rect 12984 26138 13040 26140
rect 13064 26138 13120 26140
rect 13144 26138 13200 26140
rect 12904 26086 12950 26138
rect 12950 26086 12960 26138
rect 12984 26086 13014 26138
rect 13014 26086 13026 26138
rect 13026 26086 13040 26138
rect 13064 26086 13078 26138
rect 13078 26086 13090 26138
rect 13090 26086 13120 26138
rect 13144 26086 13154 26138
rect 13154 26086 13200 26138
rect 12904 26084 12960 26086
rect 12984 26084 13040 26086
rect 13064 26084 13120 26086
rect 13144 26084 13200 26086
rect 6930 25594 6986 25596
rect 7010 25594 7066 25596
rect 7090 25594 7146 25596
rect 7170 25594 7226 25596
rect 6930 25542 6976 25594
rect 6976 25542 6986 25594
rect 7010 25542 7040 25594
rect 7040 25542 7052 25594
rect 7052 25542 7066 25594
rect 7090 25542 7104 25594
rect 7104 25542 7116 25594
rect 7116 25542 7146 25594
rect 7170 25542 7180 25594
rect 7180 25542 7226 25594
rect 6930 25540 6986 25542
rect 7010 25540 7066 25542
rect 7090 25540 7146 25542
rect 7170 25540 7226 25542
rect 18878 25594 18934 25596
rect 18958 25594 19014 25596
rect 19038 25594 19094 25596
rect 19118 25594 19174 25596
rect 18878 25542 18924 25594
rect 18924 25542 18934 25594
rect 18958 25542 18988 25594
rect 18988 25542 19000 25594
rect 19000 25542 19014 25594
rect 19038 25542 19052 25594
rect 19052 25542 19064 25594
rect 19064 25542 19094 25594
rect 19118 25542 19128 25594
rect 19128 25542 19174 25594
rect 18878 25540 18934 25542
rect 18958 25540 19014 25542
rect 19038 25540 19094 25542
rect 19118 25540 19174 25542
rect 1398 25236 1400 25256
rect 1400 25236 1452 25256
rect 1452 25236 1454 25256
rect 1398 25200 1454 25236
rect 12904 25050 12960 25052
rect 12984 25050 13040 25052
rect 13064 25050 13120 25052
rect 13144 25050 13200 25052
rect 12904 24998 12950 25050
rect 12950 24998 12960 25050
rect 12984 24998 13014 25050
rect 13014 24998 13026 25050
rect 13026 24998 13040 25050
rect 13064 24998 13078 25050
rect 13078 24998 13090 25050
rect 13090 24998 13120 25050
rect 13144 24998 13154 25050
rect 13154 24998 13200 25050
rect 12904 24996 12960 24998
rect 12984 24996 13040 24998
rect 13064 24996 13120 24998
rect 13144 24996 13200 24998
rect 1398 24556 1400 24576
rect 1400 24556 1452 24576
rect 1452 24556 1454 24576
rect 1398 24520 1454 24556
rect 6930 24506 6986 24508
rect 7010 24506 7066 24508
rect 7090 24506 7146 24508
rect 7170 24506 7226 24508
rect 6930 24454 6976 24506
rect 6976 24454 6986 24506
rect 7010 24454 7040 24506
rect 7040 24454 7052 24506
rect 7052 24454 7066 24506
rect 7090 24454 7104 24506
rect 7104 24454 7116 24506
rect 7116 24454 7146 24506
rect 7170 24454 7180 24506
rect 7180 24454 7226 24506
rect 6930 24452 6986 24454
rect 7010 24452 7066 24454
rect 7090 24452 7146 24454
rect 7170 24452 7226 24454
rect 18878 24506 18934 24508
rect 18958 24506 19014 24508
rect 19038 24506 19094 24508
rect 19118 24506 19174 24508
rect 18878 24454 18924 24506
rect 18924 24454 18934 24506
rect 18958 24454 18988 24506
rect 18988 24454 19000 24506
rect 19000 24454 19014 24506
rect 19038 24454 19052 24506
rect 19052 24454 19064 24506
rect 19064 24454 19094 24506
rect 19118 24454 19128 24506
rect 19128 24454 19174 24506
rect 18878 24452 18934 24454
rect 18958 24452 19014 24454
rect 19038 24452 19094 24454
rect 19118 24452 19174 24454
rect 12904 23962 12960 23964
rect 12984 23962 13040 23964
rect 13064 23962 13120 23964
rect 13144 23962 13200 23964
rect 12904 23910 12950 23962
rect 12950 23910 12960 23962
rect 12984 23910 13014 23962
rect 13014 23910 13026 23962
rect 13026 23910 13040 23962
rect 13064 23910 13078 23962
rect 13078 23910 13090 23962
rect 13090 23910 13120 23962
rect 13144 23910 13154 23962
rect 13154 23910 13200 23962
rect 12904 23908 12960 23910
rect 12984 23908 13040 23910
rect 13064 23908 13120 23910
rect 13144 23908 13200 23910
rect 1398 23840 1454 23896
rect 6930 23418 6986 23420
rect 7010 23418 7066 23420
rect 7090 23418 7146 23420
rect 7170 23418 7226 23420
rect 6930 23366 6976 23418
rect 6976 23366 6986 23418
rect 7010 23366 7040 23418
rect 7040 23366 7052 23418
rect 7052 23366 7066 23418
rect 7090 23366 7104 23418
rect 7104 23366 7116 23418
rect 7116 23366 7146 23418
rect 7170 23366 7180 23418
rect 7180 23366 7226 23418
rect 6930 23364 6986 23366
rect 7010 23364 7066 23366
rect 7090 23364 7146 23366
rect 7170 23364 7226 23366
rect 18878 23418 18934 23420
rect 18958 23418 19014 23420
rect 19038 23418 19094 23420
rect 19118 23418 19174 23420
rect 18878 23366 18924 23418
rect 18924 23366 18934 23418
rect 18958 23366 18988 23418
rect 18988 23366 19000 23418
rect 19000 23366 19014 23418
rect 19038 23366 19052 23418
rect 19052 23366 19064 23418
rect 19064 23366 19094 23418
rect 19118 23366 19128 23418
rect 19128 23366 19174 23418
rect 18878 23364 18934 23366
rect 18958 23364 19014 23366
rect 19038 23364 19094 23366
rect 19118 23364 19174 23366
rect 1398 23160 1454 23216
rect 12904 22874 12960 22876
rect 12984 22874 13040 22876
rect 13064 22874 13120 22876
rect 13144 22874 13200 22876
rect 12904 22822 12950 22874
rect 12950 22822 12960 22874
rect 12984 22822 13014 22874
rect 13014 22822 13026 22874
rect 13026 22822 13040 22874
rect 13064 22822 13078 22874
rect 13078 22822 13090 22874
rect 13090 22822 13120 22874
rect 13144 22822 13154 22874
rect 13154 22822 13200 22874
rect 12904 22820 12960 22822
rect 12984 22820 13040 22822
rect 13064 22820 13120 22822
rect 13144 22820 13200 22822
rect 6930 22330 6986 22332
rect 7010 22330 7066 22332
rect 7090 22330 7146 22332
rect 7170 22330 7226 22332
rect 6930 22278 6976 22330
rect 6976 22278 6986 22330
rect 7010 22278 7040 22330
rect 7040 22278 7052 22330
rect 7052 22278 7066 22330
rect 7090 22278 7104 22330
rect 7104 22278 7116 22330
rect 7116 22278 7146 22330
rect 7170 22278 7180 22330
rect 7180 22278 7226 22330
rect 6930 22276 6986 22278
rect 7010 22276 7066 22278
rect 7090 22276 7146 22278
rect 7170 22276 7226 22278
rect 18878 22330 18934 22332
rect 18958 22330 19014 22332
rect 19038 22330 19094 22332
rect 19118 22330 19174 22332
rect 18878 22278 18924 22330
rect 18924 22278 18934 22330
rect 18958 22278 18988 22330
rect 18988 22278 19000 22330
rect 19000 22278 19014 22330
rect 19038 22278 19052 22330
rect 19052 22278 19064 22330
rect 19064 22278 19094 22330
rect 19118 22278 19128 22330
rect 19128 22278 19174 22330
rect 18878 22276 18934 22278
rect 18958 22276 19014 22278
rect 19038 22276 19094 22278
rect 19118 22276 19174 22278
rect 1398 21800 1454 21856
rect 12904 21786 12960 21788
rect 12984 21786 13040 21788
rect 13064 21786 13120 21788
rect 13144 21786 13200 21788
rect 12904 21734 12950 21786
rect 12950 21734 12960 21786
rect 12984 21734 13014 21786
rect 13014 21734 13026 21786
rect 13026 21734 13040 21786
rect 13064 21734 13078 21786
rect 13078 21734 13090 21786
rect 13090 21734 13120 21786
rect 13144 21734 13154 21786
rect 13154 21734 13200 21786
rect 12904 21732 12960 21734
rect 12984 21732 13040 21734
rect 13064 21732 13120 21734
rect 13144 21732 13200 21734
rect 6930 21242 6986 21244
rect 7010 21242 7066 21244
rect 7090 21242 7146 21244
rect 7170 21242 7226 21244
rect 6930 21190 6976 21242
rect 6976 21190 6986 21242
rect 7010 21190 7040 21242
rect 7040 21190 7052 21242
rect 7052 21190 7066 21242
rect 7090 21190 7104 21242
rect 7104 21190 7116 21242
rect 7116 21190 7146 21242
rect 7170 21190 7180 21242
rect 7180 21190 7226 21242
rect 6930 21188 6986 21190
rect 7010 21188 7066 21190
rect 7090 21188 7146 21190
rect 7170 21188 7226 21190
rect 18878 21242 18934 21244
rect 18958 21242 19014 21244
rect 19038 21242 19094 21244
rect 19118 21242 19174 21244
rect 18878 21190 18924 21242
rect 18924 21190 18934 21242
rect 18958 21190 18988 21242
rect 18988 21190 19000 21242
rect 19000 21190 19014 21242
rect 19038 21190 19052 21242
rect 19052 21190 19064 21242
rect 19064 21190 19094 21242
rect 19118 21190 19128 21242
rect 19128 21190 19174 21242
rect 18878 21188 18934 21190
rect 18958 21188 19014 21190
rect 19038 21188 19094 21190
rect 19118 21188 19174 21190
rect 1398 21120 1454 21176
rect 12904 20698 12960 20700
rect 12984 20698 13040 20700
rect 13064 20698 13120 20700
rect 13144 20698 13200 20700
rect 12904 20646 12950 20698
rect 12950 20646 12960 20698
rect 12984 20646 13014 20698
rect 13014 20646 13026 20698
rect 13026 20646 13040 20698
rect 13064 20646 13078 20698
rect 13078 20646 13090 20698
rect 13090 20646 13120 20698
rect 13144 20646 13154 20698
rect 13154 20646 13200 20698
rect 12904 20644 12960 20646
rect 12984 20644 13040 20646
rect 13064 20644 13120 20646
rect 13144 20644 13200 20646
rect 1398 20440 1454 20496
rect 6930 20154 6986 20156
rect 7010 20154 7066 20156
rect 7090 20154 7146 20156
rect 7170 20154 7226 20156
rect 6930 20102 6976 20154
rect 6976 20102 6986 20154
rect 7010 20102 7040 20154
rect 7040 20102 7052 20154
rect 7052 20102 7066 20154
rect 7090 20102 7104 20154
rect 7104 20102 7116 20154
rect 7116 20102 7146 20154
rect 7170 20102 7180 20154
rect 7180 20102 7226 20154
rect 6930 20100 6986 20102
rect 7010 20100 7066 20102
rect 7090 20100 7146 20102
rect 7170 20100 7226 20102
rect 18878 20154 18934 20156
rect 18958 20154 19014 20156
rect 19038 20154 19094 20156
rect 19118 20154 19174 20156
rect 18878 20102 18924 20154
rect 18924 20102 18934 20154
rect 18958 20102 18988 20154
rect 18988 20102 19000 20154
rect 19000 20102 19014 20154
rect 19038 20102 19052 20154
rect 19052 20102 19064 20154
rect 19064 20102 19094 20154
rect 19118 20102 19128 20154
rect 19128 20102 19174 20154
rect 18878 20100 18934 20102
rect 18958 20100 19014 20102
rect 19038 20100 19094 20102
rect 19118 20100 19174 20102
rect 1398 19796 1400 19816
rect 1400 19796 1452 19816
rect 1452 19796 1454 19816
rect 1398 19760 1454 19796
rect 12904 19610 12960 19612
rect 12984 19610 13040 19612
rect 13064 19610 13120 19612
rect 13144 19610 13200 19612
rect 12904 19558 12950 19610
rect 12950 19558 12960 19610
rect 12984 19558 13014 19610
rect 13014 19558 13026 19610
rect 13026 19558 13040 19610
rect 13064 19558 13078 19610
rect 13078 19558 13090 19610
rect 13090 19558 13120 19610
rect 13144 19558 13154 19610
rect 13154 19558 13200 19610
rect 12904 19556 12960 19558
rect 12984 19556 13040 19558
rect 13064 19556 13120 19558
rect 13144 19556 13200 19558
rect 1398 19116 1400 19136
rect 1400 19116 1452 19136
rect 1452 19116 1454 19136
rect 1398 19080 1454 19116
rect 6930 19066 6986 19068
rect 7010 19066 7066 19068
rect 7090 19066 7146 19068
rect 7170 19066 7226 19068
rect 6930 19014 6976 19066
rect 6976 19014 6986 19066
rect 7010 19014 7040 19066
rect 7040 19014 7052 19066
rect 7052 19014 7066 19066
rect 7090 19014 7104 19066
rect 7104 19014 7116 19066
rect 7116 19014 7146 19066
rect 7170 19014 7180 19066
rect 7180 19014 7226 19066
rect 6930 19012 6986 19014
rect 7010 19012 7066 19014
rect 7090 19012 7146 19014
rect 7170 19012 7226 19014
rect 18878 19066 18934 19068
rect 18958 19066 19014 19068
rect 19038 19066 19094 19068
rect 19118 19066 19174 19068
rect 18878 19014 18924 19066
rect 18924 19014 18934 19066
rect 18958 19014 18988 19066
rect 18988 19014 19000 19066
rect 19000 19014 19014 19066
rect 19038 19014 19052 19066
rect 19052 19014 19064 19066
rect 19064 19014 19094 19066
rect 19118 19014 19128 19066
rect 19128 19014 19174 19066
rect 18878 19012 18934 19014
rect 18958 19012 19014 19014
rect 19038 19012 19094 19014
rect 19118 19012 19174 19014
rect 12904 18522 12960 18524
rect 12984 18522 13040 18524
rect 13064 18522 13120 18524
rect 13144 18522 13200 18524
rect 12904 18470 12950 18522
rect 12950 18470 12960 18522
rect 12984 18470 13014 18522
rect 13014 18470 13026 18522
rect 13026 18470 13040 18522
rect 13064 18470 13078 18522
rect 13078 18470 13090 18522
rect 13090 18470 13120 18522
rect 13144 18470 13154 18522
rect 13154 18470 13200 18522
rect 12904 18468 12960 18470
rect 12984 18468 13040 18470
rect 13064 18468 13120 18470
rect 13144 18468 13200 18470
rect 1398 18400 1454 18456
rect 6930 17978 6986 17980
rect 7010 17978 7066 17980
rect 7090 17978 7146 17980
rect 7170 17978 7226 17980
rect 6930 17926 6976 17978
rect 6976 17926 6986 17978
rect 7010 17926 7040 17978
rect 7040 17926 7052 17978
rect 7052 17926 7066 17978
rect 7090 17926 7104 17978
rect 7104 17926 7116 17978
rect 7116 17926 7146 17978
rect 7170 17926 7180 17978
rect 7180 17926 7226 17978
rect 6930 17924 6986 17926
rect 7010 17924 7066 17926
rect 7090 17924 7146 17926
rect 7170 17924 7226 17926
rect 18878 17978 18934 17980
rect 18958 17978 19014 17980
rect 19038 17978 19094 17980
rect 19118 17978 19174 17980
rect 18878 17926 18924 17978
rect 18924 17926 18934 17978
rect 18958 17926 18988 17978
rect 18988 17926 19000 17978
rect 19000 17926 19014 17978
rect 19038 17926 19052 17978
rect 19052 17926 19064 17978
rect 19064 17926 19094 17978
rect 19118 17926 19128 17978
rect 19128 17926 19174 17978
rect 18878 17924 18934 17926
rect 18958 17924 19014 17926
rect 19038 17924 19094 17926
rect 19118 17924 19174 17926
rect 12904 17434 12960 17436
rect 12984 17434 13040 17436
rect 13064 17434 13120 17436
rect 13144 17434 13200 17436
rect 12904 17382 12950 17434
rect 12950 17382 12960 17434
rect 12984 17382 13014 17434
rect 13014 17382 13026 17434
rect 13026 17382 13040 17434
rect 13064 17382 13078 17434
rect 13078 17382 13090 17434
rect 13090 17382 13120 17434
rect 13144 17382 13154 17434
rect 13154 17382 13200 17434
rect 12904 17380 12960 17382
rect 12984 17380 13040 17382
rect 13064 17380 13120 17382
rect 13144 17380 13200 17382
rect 6930 16890 6986 16892
rect 7010 16890 7066 16892
rect 7090 16890 7146 16892
rect 7170 16890 7226 16892
rect 6930 16838 6976 16890
rect 6976 16838 6986 16890
rect 7010 16838 7040 16890
rect 7040 16838 7052 16890
rect 7052 16838 7066 16890
rect 7090 16838 7104 16890
rect 7104 16838 7116 16890
rect 7116 16838 7146 16890
rect 7170 16838 7180 16890
rect 7180 16838 7226 16890
rect 6930 16836 6986 16838
rect 7010 16836 7066 16838
rect 7090 16836 7146 16838
rect 7170 16836 7226 16838
rect 18878 16890 18934 16892
rect 18958 16890 19014 16892
rect 19038 16890 19094 16892
rect 19118 16890 19174 16892
rect 18878 16838 18924 16890
rect 18924 16838 18934 16890
rect 18958 16838 18988 16890
rect 18988 16838 19000 16890
rect 19000 16838 19014 16890
rect 19038 16838 19052 16890
rect 19052 16838 19064 16890
rect 19064 16838 19094 16890
rect 19118 16838 19128 16890
rect 19128 16838 19174 16890
rect 18878 16836 18934 16838
rect 18958 16836 19014 16838
rect 19038 16836 19094 16838
rect 19118 16836 19174 16838
rect 12904 16346 12960 16348
rect 12984 16346 13040 16348
rect 13064 16346 13120 16348
rect 13144 16346 13200 16348
rect 12904 16294 12950 16346
rect 12950 16294 12960 16346
rect 12984 16294 13014 16346
rect 13014 16294 13026 16346
rect 13026 16294 13040 16346
rect 13064 16294 13078 16346
rect 13078 16294 13090 16346
rect 13090 16294 13120 16346
rect 13144 16294 13154 16346
rect 13154 16294 13200 16346
rect 12904 16292 12960 16294
rect 12984 16292 13040 16294
rect 13064 16292 13120 16294
rect 13144 16292 13200 16294
rect 6930 15802 6986 15804
rect 7010 15802 7066 15804
rect 7090 15802 7146 15804
rect 7170 15802 7226 15804
rect 6930 15750 6976 15802
rect 6976 15750 6986 15802
rect 7010 15750 7040 15802
rect 7040 15750 7052 15802
rect 7052 15750 7066 15802
rect 7090 15750 7104 15802
rect 7104 15750 7116 15802
rect 7116 15750 7146 15802
rect 7170 15750 7180 15802
rect 7180 15750 7226 15802
rect 6930 15748 6986 15750
rect 7010 15748 7066 15750
rect 7090 15748 7146 15750
rect 7170 15748 7226 15750
rect 18878 15802 18934 15804
rect 18958 15802 19014 15804
rect 19038 15802 19094 15804
rect 19118 15802 19174 15804
rect 18878 15750 18924 15802
rect 18924 15750 18934 15802
rect 18958 15750 18988 15802
rect 18988 15750 19000 15802
rect 19000 15750 19014 15802
rect 19038 15750 19052 15802
rect 19052 15750 19064 15802
rect 19064 15750 19094 15802
rect 19118 15750 19128 15802
rect 19128 15750 19174 15802
rect 18878 15748 18934 15750
rect 18958 15748 19014 15750
rect 19038 15748 19094 15750
rect 19118 15748 19174 15750
rect 1398 15680 1454 15736
rect 12904 15258 12960 15260
rect 12984 15258 13040 15260
rect 13064 15258 13120 15260
rect 13144 15258 13200 15260
rect 12904 15206 12950 15258
rect 12950 15206 12960 15258
rect 12984 15206 13014 15258
rect 13014 15206 13026 15258
rect 13026 15206 13040 15258
rect 13064 15206 13078 15258
rect 13078 15206 13090 15258
rect 13090 15206 13120 15258
rect 13144 15206 13154 15258
rect 13154 15206 13200 15258
rect 12904 15204 12960 15206
rect 12984 15204 13040 15206
rect 13064 15204 13120 15206
rect 13144 15204 13200 15206
rect 1398 15000 1454 15056
rect 24852 27226 24908 27228
rect 24932 27226 24988 27228
rect 25012 27226 25068 27228
rect 25092 27226 25148 27228
rect 24852 27174 24898 27226
rect 24898 27174 24908 27226
rect 24932 27174 24962 27226
rect 24962 27174 24974 27226
rect 24974 27174 24988 27226
rect 25012 27174 25026 27226
rect 25026 27174 25038 27226
rect 25038 27174 25068 27226
rect 25092 27174 25102 27226
rect 25102 27174 25148 27226
rect 24852 27172 24908 27174
rect 24932 27172 24988 27174
rect 25012 27172 25068 27174
rect 25092 27172 25148 27174
rect 36800 27226 36856 27228
rect 36880 27226 36936 27228
rect 36960 27226 37016 27228
rect 37040 27226 37096 27228
rect 36800 27174 36846 27226
rect 36846 27174 36856 27226
rect 36880 27174 36910 27226
rect 36910 27174 36922 27226
rect 36922 27174 36936 27226
rect 36960 27174 36974 27226
rect 36974 27174 36986 27226
rect 36986 27174 37016 27226
rect 37040 27174 37050 27226
rect 37050 27174 37096 27226
rect 36800 27172 36856 27174
rect 36880 27172 36936 27174
rect 36960 27172 37016 27174
rect 37040 27172 37096 27174
rect 42774 27770 42830 27772
rect 42854 27770 42910 27772
rect 42934 27770 42990 27772
rect 43014 27770 43070 27772
rect 42774 27718 42820 27770
rect 42820 27718 42830 27770
rect 42854 27718 42884 27770
rect 42884 27718 42896 27770
rect 42896 27718 42910 27770
rect 42934 27718 42948 27770
rect 42948 27718 42960 27770
rect 42960 27718 42990 27770
rect 43014 27718 43024 27770
rect 43024 27718 43070 27770
rect 42774 27716 42830 27718
rect 42854 27716 42910 27718
rect 42934 27716 42990 27718
rect 43014 27716 43070 27718
rect 45742 28192 45798 28248
rect 47490 27648 47546 27704
rect 46846 26832 46902 26888
rect 30826 26682 30882 26684
rect 30906 26682 30962 26684
rect 30986 26682 31042 26684
rect 31066 26682 31122 26684
rect 30826 26630 30872 26682
rect 30872 26630 30882 26682
rect 30906 26630 30936 26682
rect 30936 26630 30948 26682
rect 30948 26630 30962 26682
rect 30986 26630 31000 26682
rect 31000 26630 31012 26682
rect 31012 26630 31042 26682
rect 31066 26630 31076 26682
rect 31076 26630 31122 26682
rect 30826 26628 30882 26630
rect 30906 26628 30962 26630
rect 30986 26628 31042 26630
rect 31066 26628 31122 26630
rect 42774 26682 42830 26684
rect 42854 26682 42910 26684
rect 42934 26682 42990 26684
rect 43014 26682 43070 26684
rect 42774 26630 42820 26682
rect 42820 26630 42830 26682
rect 42854 26630 42884 26682
rect 42884 26630 42896 26682
rect 42896 26630 42910 26682
rect 42934 26630 42948 26682
rect 42948 26630 42960 26682
rect 42960 26630 42990 26682
rect 43014 26630 43024 26682
rect 43024 26630 43070 26682
rect 42774 26628 42830 26630
rect 42854 26628 42910 26630
rect 42934 26628 42990 26630
rect 43014 26628 43070 26630
rect 24852 26138 24908 26140
rect 24932 26138 24988 26140
rect 25012 26138 25068 26140
rect 25092 26138 25148 26140
rect 24852 26086 24898 26138
rect 24898 26086 24908 26138
rect 24932 26086 24962 26138
rect 24962 26086 24974 26138
rect 24974 26086 24988 26138
rect 25012 26086 25026 26138
rect 25026 26086 25038 26138
rect 25038 26086 25068 26138
rect 25092 26086 25102 26138
rect 25102 26086 25148 26138
rect 24852 26084 24908 26086
rect 24932 26084 24988 26086
rect 25012 26084 25068 26086
rect 25092 26084 25148 26086
rect 36800 26138 36856 26140
rect 36880 26138 36936 26140
rect 36960 26138 37016 26140
rect 37040 26138 37096 26140
rect 36800 26086 36846 26138
rect 36846 26086 36856 26138
rect 36880 26086 36910 26138
rect 36910 26086 36922 26138
rect 36922 26086 36936 26138
rect 36960 26086 36974 26138
rect 36974 26086 36986 26138
rect 36986 26086 37016 26138
rect 37040 26086 37050 26138
rect 37050 26086 37096 26138
rect 36800 26084 36856 26086
rect 36880 26084 36936 26086
rect 36960 26084 37016 26086
rect 37040 26084 37096 26086
rect 30826 25594 30882 25596
rect 30906 25594 30962 25596
rect 30986 25594 31042 25596
rect 31066 25594 31122 25596
rect 30826 25542 30872 25594
rect 30872 25542 30882 25594
rect 30906 25542 30936 25594
rect 30936 25542 30948 25594
rect 30948 25542 30962 25594
rect 30986 25542 31000 25594
rect 31000 25542 31012 25594
rect 31012 25542 31042 25594
rect 31066 25542 31076 25594
rect 31076 25542 31122 25594
rect 30826 25540 30882 25542
rect 30906 25540 30962 25542
rect 30986 25540 31042 25542
rect 31066 25540 31122 25542
rect 42774 25594 42830 25596
rect 42854 25594 42910 25596
rect 42934 25594 42990 25596
rect 43014 25594 43070 25596
rect 42774 25542 42820 25594
rect 42820 25542 42830 25594
rect 42854 25542 42884 25594
rect 42884 25542 42896 25594
rect 42896 25542 42910 25594
rect 42934 25542 42948 25594
rect 42948 25542 42960 25594
rect 42960 25542 42990 25594
rect 43014 25542 43024 25594
rect 43024 25542 43070 25594
rect 42774 25540 42830 25542
rect 42854 25540 42910 25542
rect 42934 25540 42990 25542
rect 43014 25540 43070 25542
rect 24852 25050 24908 25052
rect 24932 25050 24988 25052
rect 25012 25050 25068 25052
rect 25092 25050 25148 25052
rect 24852 24998 24898 25050
rect 24898 24998 24908 25050
rect 24932 24998 24962 25050
rect 24962 24998 24974 25050
rect 24974 24998 24988 25050
rect 25012 24998 25026 25050
rect 25026 24998 25038 25050
rect 25038 24998 25068 25050
rect 25092 24998 25102 25050
rect 25102 24998 25148 25050
rect 24852 24996 24908 24998
rect 24932 24996 24988 24998
rect 25012 24996 25068 24998
rect 25092 24996 25148 24998
rect 36800 25050 36856 25052
rect 36880 25050 36936 25052
rect 36960 25050 37016 25052
rect 37040 25050 37096 25052
rect 36800 24998 36846 25050
rect 36846 24998 36856 25050
rect 36880 24998 36910 25050
rect 36910 24998 36922 25050
rect 36922 24998 36936 25050
rect 36960 24998 36974 25050
rect 36974 24998 36986 25050
rect 36986 24998 37016 25050
rect 37040 24998 37050 25050
rect 37050 24998 37096 25050
rect 36800 24996 36856 24998
rect 36880 24996 36936 24998
rect 36960 24996 37016 24998
rect 37040 24996 37096 24998
rect 30826 24506 30882 24508
rect 30906 24506 30962 24508
rect 30986 24506 31042 24508
rect 31066 24506 31122 24508
rect 30826 24454 30872 24506
rect 30872 24454 30882 24506
rect 30906 24454 30936 24506
rect 30936 24454 30948 24506
rect 30948 24454 30962 24506
rect 30986 24454 31000 24506
rect 31000 24454 31012 24506
rect 31012 24454 31042 24506
rect 31066 24454 31076 24506
rect 31076 24454 31122 24506
rect 30826 24452 30882 24454
rect 30906 24452 30962 24454
rect 30986 24452 31042 24454
rect 31066 24452 31122 24454
rect 42774 24506 42830 24508
rect 42854 24506 42910 24508
rect 42934 24506 42990 24508
rect 43014 24506 43070 24508
rect 42774 24454 42820 24506
rect 42820 24454 42830 24506
rect 42854 24454 42884 24506
rect 42884 24454 42896 24506
rect 42896 24454 42910 24506
rect 42934 24454 42948 24506
rect 42948 24454 42960 24506
rect 42960 24454 42990 24506
rect 43014 24454 43024 24506
rect 43024 24454 43070 24506
rect 42774 24452 42830 24454
rect 42854 24452 42910 24454
rect 42934 24452 42990 24454
rect 43014 24452 43070 24454
rect 24852 23962 24908 23964
rect 24932 23962 24988 23964
rect 25012 23962 25068 23964
rect 25092 23962 25148 23964
rect 24852 23910 24898 23962
rect 24898 23910 24908 23962
rect 24932 23910 24962 23962
rect 24962 23910 24974 23962
rect 24974 23910 24988 23962
rect 25012 23910 25026 23962
rect 25026 23910 25038 23962
rect 25038 23910 25068 23962
rect 25092 23910 25102 23962
rect 25102 23910 25148 23962
rect 24852 23908 24908 23910
rect 24932 23908 24988 23910
rect 25012 23908 25068 23910
rect 25092 23908 25148 23910
rect 36800 23962 36856 23964
rect 36880 23962 36936 23964
rect 36960 23962 37016 23964
rect 37040 23962 37096 23964
rect 36800 23910 36846 23962
rect 36846 23910 36856 23962
rect 36880 23910 36910 23962
rect 36910 23910 36922 23962
rect 36922 23910 36936 23962
rect 36960 23910 36974 23962
rect 36974 23910 36986 23962
rect 36986 23910 37016 23962
rect 37040 23910 37050 23962
rect 37050 23910 37096 23962
rect 36800 23908 36856 23910
rect 36880 23908 36936 23910
rect 36960 23908 37016 23910
rect 37040 23908 37096 23910
rect 30826 23418 30882 23420
rect 30906 23418 30962 23420
rect 30986 23418 31042 23420
rect 31066 23418 31122 23420
rect 30826 23366 30872 23418
rect 30872 23366 30882 23418
rect 30906 23366 30936 23418
rect 30936 23366 30948 23418
rect 30948 23366 30962 23418
rect 30986 23366 31000 23418
rect 31000 23366 31012 23418
rect 31012 23366 31042 23418
rect 31066 23366 31076 23418
rect 31076 23366 31122 23418
rect 30826 23364 30882 23366
rect 30906 23364 30962 23366
rect 30986 23364 31042 23366
rect 31066 23364 31122 23366
rect 42774 23418 42830 23420
rect 42854 23418 42910 23420
rect 42934 23418 42990 23420
rect 43014 23418 43070 23420
rect 42774 23366 42820 23418
rect 42820 23366 42830 23418
rect 42854 23366 42884 23418
rect 42884 23366 42896 23418
rect 42896 23366 42910 23418
rect 42934 23366 42948 23418
rect 42948 23366 42960 23418
rect 42960 23366 42990 23418
rect 43014 23366 43024 23418
rect 43024 23366 43070 23418
rect 42774 23364 42830 23366
rect 42854 23364 42910 23366
rect 42934 23364 42990 23366
rect 43014 23364 43070 23366
rect 24852 22874 24908 22876
rect 24932 22874 24988 22876
rect 25012 22874 25068 22876
rect 25092 22874 25148 22876
rect 24852 22822 24898 22874
rect 24898 22822 24908 22874
rect 24932 22822 24962 22874
rect 24962 22822 24974 22874
rect 24974 22822 24988 22874
rect 25012 22822 25026 22874
rect 25026 22822 25038 22874
rect 25038 22822 25068 22874
rect 25092 22822 25102 22874
rect 25102 22822 25148 22874
rect 24852 22820 24908 22822
rect 24932 22820 24988 22822
rect 25012 22820 25068 22822
rect 25092 22820 25148 22822
rect 36800 22874 36856 22876
rect 36880 22874 36936 22876
rect 36960 22874 37016 22876
rect 37040 22874 37096 22876
rect 36800 22822 36846 22874
rect 36846 22822 36856 22874
rect 36880 22822 36910 22874
rect 36910 22822 36922 22874
rect 36922 22822 36936 22874
rect 36960 22822 36974 22874
rect 36974 22822 36986 22874
rect 36986 22822 37016 22874
rect 37040 22822 37050 22874
rect 37050 22822 37096 22874
rect 36800 22820 36856 22822
rect 36880 22820 36936 22822
rect 36960 22820 37016 22822
rect 37040 22820 37096 22822
rect 30826 22330 30882 22332
rect 30906 22330 30962 22332
rect 30986 22330 31042 22332
rect 31066 22330 31122 22332
rect 30826 22278 30872 22330
rect 30872 22278 30882 22330
rect 30906 22278 30936 22330
rect 30936 22278 30948 22330
rect 30948 22278 30962 22330
rect 30986 22278 31000 22330
rect 31000 22278 31012 22330
rect 31012 22278 31042 22330
rect 31066 22278 31076 22330
rect 31076 22278 31122 22330
rect 30826 22276 30882 22278
rect 30906 22276 30962 22278
rect 30986 22276 31042 22278
rect 31066 22276 31122 22278
rect 42774 22330 42830 22332
rect 42854 22330 42910 22332
rect 42934 22330 42990 22332
rect 43014 22330 43070 22332
rect 42774 22278 42820 22330
rect 42820 22278 42830 22330
rect 42854 22278 42884 22330
rect 42884 22278 42896 22330
rect 42896 22278 42910 22330
rect 42934 22278 42948 22330
rect 42948 22278 42960 22330
rect 42960 22278 42990 22330
rect 43014 22278 43024 22330
rect 43024 22278 43070 22330
rect 42774 22276 42830 22278
rect 42854 22276 42910 22278
rect 42934 22276 42990 22278
rect 43014 22276 43070 22278
rect 24852 21786 24908 21788
rect 24932 21786 24988 21788
rect 25012 21786 25068 21788
rect 25092 21786 25148 21788
rect 24852 21734 24898 21786
rect 24898 21734 24908 21786
rect 24932 21734 24962 21786
rect 24962 21734 24974 21786
rect 24974 21734 24988 21786
rect 25012 21734 25026 21786
rect 25026 21734 25038 21786
rect 25038 21734 25068 21786
rect 25092 21734 25102 21786
rect 25102 21734 25148 21786
rect 24852 21732 24908 21734
rect 24932 21732 24988 21734
rect 25012 21732 25068 21734
rect 25092 21732 25148 21734
rect 36800 21786 36856 21788
rect 36880 21786 36936 21788
rect 36960 21786 37016 21788
rect 37040 21786 37096 21788
rect 36800 21734 36846 21786
rect 36846 21734 36856 21786
rect 36880 21734 36910 21786
rect 36910 21734 36922 21786
rect 36922 21734 36936 21786
rect 36960 21734 36974 21786
rect 36974 21734 36986 21786
rect 36986 21734 37016 21786
rect 37040 21734 37050 21786
rect 37050 21734 37096 21786
rect 36800 21732 36856 21734
rect 36880 21732 36936 21734
rect 36960 21732 37016 21734
rect 37040 21732 37096 21734
rect 30826 21242 30882 21244
rect 30906 21242 30962 21244
rect 30986 21242 31042 21244
rect 31066 21242 31122 21244
rect 30826 21190 30872 21242
rect 30872 21190 30882 21242
rect 30906 21190 30936 21242
rect 30936 21190 30948 21242
rect 30948 21190 30962 21242
rect 30986 21190 31000 21242
rect 31000 21190 31012 21242
rect 31012 21190 31042 21242
rect 31066 21190 31076 21242
rect 31076 21190 31122 21242
rect 30826 21188 30882 21190
rect 30906 21188 30962 21190
rect 30986 21188 31042 21190
rect 31066 21188 31122 21190
rect 42774 21242 42830 21244
rect 42854 21242 42910 21244
rect 42934 21242 42990 21244
rect 43014 21242 43070 21244
rect 42774 21190 42820 21242
rect 42820 21190 42830 21242
rect 42854 21190 42884 21242
rect 42884 21190 42896 21242
rect 42896 21190 42910 21242
rect 42934 21190 42948 21242
rect 42948 21190 42960 21242
rect 42960 21190 42990 21242
rect 43014 21190 43024 21242
rect 43024 21190 43070 21242
rect 42774 21188 42830 21190
rect 42854 21188 42910 21190
rect 42934 21188 42990 21190
rect 43014 21188 43070 21190
rect 24852 20698 24908 20700
rect 24932 20698 24988 20700
rect 25012 20698 25068 20700
rect 25092 20698 25148 20700
rect 24852 20646 24898 20698
rect 24898 20646 24908 20698
rect 24932 20646 24962 20698
rect 24962 20646 24974 20698
rect 24974 20646 24988 20698
rect 25012 20646 25026 20698
rect 25026 20646 25038 20698
rect 25038 20646 25068 20698
rect 25092 20646 25102 20698
rect 25102 20646 25148 20698
rect 24852 20644 24908 20646
rect 24932 20644 24988 20646
rect 25012 20644 25068 20646
rect 25092 20644 25148 20646
rect 36800 20698 36856 20700
rect 36880 20698 36936 20700
rect 36960 20698 37016 20700
rect 37040 20698 37096 20700
rect 36800 20646 36846 20698
rect 36846 20646 36856 20698
rect 36880 20646 36910 20698
rect 36910 20646 36922 20698
rect 36922 20646 36936 20698
rect 36960 20646 36974 20698
rect 36974 20646 36986 20698
rect 36986 20646 37016 20698
rect 37040 20646 37050 20698
rect 37050 20646 37096 20698
rect 36800 20644 36856 20646
rect 36880 20644 36936 20646
rect 36960 20644 37016 20646
rect 37040 20644 37096 20646
rect 30826 20154 30882 20156
rect 30906 20154 30962 20156
rect 30986 20154 31042 20156
rect 31066 20154 31122 20156
rect 30826 20102 30872 20154
rect 30872 20102 30882 20154
rect 30906 20102 30936 20154
rect 30936 20102 30948 20154
rect 30948 20102 30962 20154
rect 30986 20102 31000 20154
rect 31000 20102 31012 20154
rect 31012 20102 31042 20154
rect 31066 20102 31076 20154
rect 31076 20102 31122 20154
rect 30826 20100 30882 20102
rect 30906 20100 30962 20102
rect 30986 20100 31042 20102
rect 31066 20100 31122 20102
rect 42774 20154 42830 20156
rect 42854 20154 42910 20156
rect 42934 20154 42990 20156
rect 43014 20154 43070 20156
rect 42774 20102 42820 20154
rect 42820 20102 42830 20154
rect 42854 20102 42884 20154
rect 42884 20102 42896 20154
rect 42896 20102 42910 20154
rect 42934 20102 42948 20154
rect 42948 20102 42960 20154
rect 42960 20102 42990 20154
rect 43014 20102 43024 20154
rect 43024 20102 43070 20154
rect 42774 20100 42830 20102
rect 42854 20100 42910 20102
rect 42934 20100 42990 20102
rect 43014 20100 43070 20102
rect 24852 19610 24908 19612
rect 24932 19610 24988 19612
rect 25012 19610 25068 19612
rect 25092 19610 25148 19612
rect 24852 19558 24898 19610
rect 24898 19558 24908 19610
rect 24932 19558 24962 19610
rect 24962 19558 24974 19610
rect 24974 19558 24988 19610
rect 25012 19558 25026 19610
rect 25026 19558 25038 19610
rect 25038 19558 25068 19610
rect 25092 19558 25102 19610
rect 25102 19558 25148 19610
rect 24852 19556 24908 19558
rect 24932 19556 24988 19558
rect 25012 19556 25068 19558
rect 25092 19556 25148 19558
rect 36800 19610 36856 19612
rect 36880 19610 36936 19612
rect 36960 19610 37016 19612
rect 37040 19610 37096 19612
rect 36800 19558 36846 19610
rect 36846 19558 36856 19610
rect 36880 19558 36910 19610
rect 36910 19558 36922 19610
rect 36922 19558 36936 19610
rect 36960 19558 36974 19610
rect 36974 19558 36986 19610
rect 36986 19558 37016 19610
rect 37040 19558 37050 19610
rect 37050 19558 37096 19610
rect 36800 19556 36856 19558
rect 36880 19556 36936 19558
rect 36960 19556 37016 19558
rect 37040 19556 37096 19558
rect 30826 19066 30882 19068
rect 30906 19066 30962 19068
rect 30986 19066 31042 19068
rect 31066 19066 31122 19068
rect 30826 19014 30872 19066
rect 30872 19014 30882 19066
rect 30906 19014 30936 19066
rect 30936 19014 30948 19066
rect 30948 19014 30962 19066
rect 30986 19014 31000 19066
rect 31000 19014 31012 19066
rect 31012 19014 31042 19066
rect 31066 19014 31076 19066
rect 31076 19014 31122 19066
rect 30826 19012 30882 19014
rect 30906 19012 30962 19014
rect 30986 19012 31042 19014
rect 31066 19012 31122 19014
rect 42774 19066 42830 19068
rect 42854 19066 42910 19068
rect 42934 19066 42990 19068
rect 43014 19066 43070 19068
rect 42774 19014 42820 19066
rect 42820 19014 42830 19066
rect 42854 19014 42884 19066
rect 42884 19014 42896 19066
rect 42896 19014 42910 19066
rect 42934 19014 42948 19066
rect 42948 19014 42960 19066
rect 42960 19014 42990 19066
rect 43014 19014 43024 19066
rect 43024 19014 43070 19066
rect 42774 19012 42830 19014
rect 42854 19012 42910 19014
rect 42934 19012 42990 19014
rect 43014 19012 43070 19014
rect 24852 18522 24908 18524
rect 24932 18522 24988 18524
rect 25012 18522 25068 18524
rect 25092 18522 25148 18524
rect 24852 18470 24898 18522
rect 24898 18470 24908 18522
rect 24932 18470 24962 18522
rect 24962 18470 24974 18522
rect 24974 18470 24988 18522
rect 25012 18470 25026 18522
rect 25026 18470 25038 18522
rect 25038 18470 25068 18522
rect 25092 18470 25102 18522
rect 25102 18470 25148 18522
rect 24852 18468 24908 18470
rect 24932 18468 24988 18470
rect 25012 18468 25068 18470
rect 25092 18468 25148 18470
rect 36800 18522 36856 18524
rect 36880 18522 36936 18524
rect 36960 18522 37016 18524
rect 37040 18522 37096 18524
rect 36800 18470 36846 18522
rect 36846 18470 36856 18522
rect 36880 18470 36910 18522
rect 36910 18470 36922 18522
rect 36922 18470 36936 18522
rect 36960 18470 36974 18522
rect 36974 18470 36986 18522
rect 36986 18470 37016 18522
rect 37040 18470 37050 18522
rect 37050 18470 37096 18522
rect 36800 18468 36856 18470
rect 36880 18468 36936 18470
rect 36960 18468 37016 18470
rect 37040 18468 37096 18470
rect 30826 17978 30882 17980
rect 30906 17978 30962 17980
rect 30986 17978 31042 17980
rect 31066 17978 31122 17980
rect 30826 17926 30872 17978
rect 30872 17926 30882 17978
rect 30906 17926 30936 17978
rect 30936 17926 30948 17978
rect 30948 17926 30962 17978
rect 30986 17926 31000 17978
rect 31000 17926 31012 17978
rect 31012 17926 31042 17978
rect 31066 17926 31076 17978
rect 31076 17926 31122 17978
rect 30826 17924 30882 17926
rect 30906 17924 30962 17926
rect 30986 17924 31042 17926
rect 31066 17924 31122 17926
rect 42774 17978 42830 17980
rect 42854 17978 42910 17980
rect 42934 17978 42990 17980
rect 43014 17978 43070 17980
rect 42774 17926 42820 17978
rect 42820 17926 42830 17978
rect 42854 17926 42884 17978
rect 42884 17926 42896 17978
rect 42896 17926 42910 17978
rect 42934 17926 42948 17978
rect 42948 17926 42960 17978
rect 42960 17926 42990 17978
rect 43014 17926 43024 17978
rect 43024 17926 43070 17978
rect 42774 17924 42830 17926
rect 42854 17924 42910 17926
rect 42934 17924 42990 17926
rect 43014 17924 43070 17926
rect 24852 17434 24908 17436
rect 24932 17434 24988 17436
rect 25012 17434 25068 17436
rect 25092 17434 25148 17436
rect 24852 17382 24898 17434
rect 24898 17382 24908 17434
rect 24932 17382 24962 17434
rect 24962 17382 24974 17434
rect 24974 17382 24988 17434
rect 25012 17382 25026 17434
rect 25026 17382 25038 17434
rect 25038 17382 25068 17434
rect 25092 17382 25102 17434
rect 25102 17382 25148 17434
rect 24852 17380 24908 17382
rect 24932 17380 24988 17382
rect 25012 17380 25068 17382
rect 25092 17380 25148 17382
rect 36800 17434 36856 17436
rect 36880 17434 36936 17436
rect 36960 17434 37016 17436
rect 37040 17434 37096 17436
rect 36800 17382 36846 17434
rect 36846 17382 36856 17434
rect 36880 17382 36910 17434
rect 36910 17382 36922 17434
rect 36922 17382 36936 17434
rect 36960 17382 36974 17434
rect 36974 17382 36986 17434
rect 36986 17382 37016 17434
rect 37040 17382 37050 17434
rect 37050 17382 37096 17434
rect 36800 17380 36856 17382
rect 36880 17380 36936 17382
rect 36960 17380 37016 17382
rect 37040 17380 37096 17382
rect 30826 16890 30882 16892
rect 30906 16890 30962 16892
rect 30986 16890 31042 16892
rect 31066 16890 31122 16892
rect 30826 16838 30872 16890
rect 30872 16838 30882 16890
rect 30906 16838 30936 16890
rect 30936 16838 30948 16890
rect 30948 16838 30962 16890
rect 30986 16838 31000 16890
rect 31000 16838 31012 16890
rect 31012 16838 31042 16890
rect 31066 16838 31076 16890
rect 31076 16838 31122 16890
rect 30826 16836 30882 16838
rect 30906 16836 30962 16838
rect 30986 16836 31042 16838
rect 31066 16836 31122 16838
rect 42774 16890 42830 16892
rect 42854 16890 42910 16892
rect 42934 16890 42990 16892
rect 43014 16890 43070 16892
rect 42774 16838 42820 16890
rect 42820 16838 42830 16890
rect 42854 16838 42884 16890
rect 42884 16838 42896 16890
rect 42896 16838 42910 16890
rect 42934 16838 42948 16890
rect 42948 16838 42960 16890
rect 42960 16838 42990 16890
rect 43014 16838 43024 16890
rect 43024 16838 43070 16890
rect 42774 16836 42830 16838
rect 42854 16836 42910 16838
rect 42934 16836 42990 16838
rect 43014 16836 43070 16838
rect 24852 16346 24908 16348
rect 24932 16346 24988 16348
rect 25012 16346 25068 16348
rect 25092 16346 25148 16348
rect 24852 16294 24898 16346
rect 24898 16294 24908 16346
rect 24932 16294 24962 16346
rect 24962 16294 24974 16346
rect 24974 16294 24988 16346
rect 25012 16294 25026 16346
rect 25026 16294 25038 16346
rect 25038 16294 25068 16346
rect 25092 16294 25102 16346
rect 25102 16294 25148 16346
rect 24852 16292 24908 16294
rect 24932 16292 24988 16294
rect 25012 16292 25068 16294
rect 25092 16292 25148 16294
rect 36800 16346 36856 16348
rect 36880 16346 36936 16348
rect 36960 16346 37016 16348
rect 37040 16346 37096 16348
rect 36800 16294 36846 16346
rect 36846 16294 36856 16346
rect 36880 16294 36910 16346
rect 36910 16294 36922 16346
rect 36922 16294 36936 16346
rect 36960 16294 36974 16346
rect 36974 16294 36986 16346
rect 36986 16294 37016 16346
rect 37040 16294 37050 16346
rect 37050 16294 37096 16346
rect 36800 16292 36856 16294
rect 36880 16292 36936 16294
rect 36960 16292 37016 16294
rect 37040 16292 37096 16294
rect 30826 15802 30882 15804
rect 30906 15802 30962 15804
rect 30986 15802 31042 15804
rect 31066 15802 31122 15804
rect 30826 15750 30872 15802
rect 30872 15750 30882 15802
rect 30906 15750 30936 15802
rect 30936 15750 30948 15802
rect 30948 15750 30962 15802
rect 30986 15750 31000 15802
rect 31000 15750 31012 15802
rect 31012 15750 31042 15802
rect 31066 15750 31076 15802
rect 31076 15750 31122 15802
rect 30826 15748 30882 15750
rect 30906 15748 30962 15750
rect 30986 15748 31042 15750
rect 31066 15748 31122 15750
rect 42774 15802 42830 15804
rect 42854 15802 42910 15804
rect 42934 15802 42990 15804
rect 43014 15802 43070 15804
rect 42774 15750 42820 15802
rect 42820 15750 42830 15802
rect 42854 15750 42884 15802
rect 42884 15750 42896 15802
rect 42896 15750 42910 15802
rect 42934 15750 42948 15802
rect 42948 15750 42960 15802
rect 42960 15750 42990 15802
rect 43014 15750 43024 15802
rect 43024 15750 43070 15802
rect 42774 15748 42830 15750
rect 42854 15748 42910 15750
rect 42934 15748 42990 15750
rect 43014 15748 43070 15750
rect 24852 15258 24908 15260
rect 24932 15258 24988 15260
rect 25012 15258 25068 15260
rect 25092 15258 25148 15260
rect 24852 15206 24898 15258
rect 24898 15206 24908 15258
rect 24932 15206 24962 15258
rect 24962 15206 24974 15258
rect 24974 15206 24988 15258
rect 25012 15206 25026 15258
rect 25026 15206 25038 15258
rect 25038 15206 25068 15258
rect 25092 15206 25102 15258
rect 25102 15206 25148 15258
rect 24852 15204 24908 15206
rect 24932 15204 24988 15206
rect 25012 15204 25068 15206
rect 25092 15204 25148 15206
rect 36800 15258 36856 15260
rect 36880 15258 36936 15260
rect 36960 15258 37016 15260
rect 37040 15258 37096 15260
rect 36800 15206 36846 15258
rect 36846 15206 36856 15258
rect 36880 15206 36910 15258
rect 36910 15206 36922 15258
rect 36922 15206 36936 15258
rect 36960 15206 36974 15258
rect 36974 15206 36986 15258
rect 36986 15206 37016 15258
rect 37040 15206 37050 15258
rect 37050 15206 37096 15258
rect 36800 15204 36856 15206
rect 36880 15204 36936 15206
rect 36960 15204 37016 15206
rect 37040 15204 37096 15206
rect 6930 14714 6986 14716
rect 7010 14714 7066 14716
rect 7090 14714 7146 14716
rect 7170 14714 7226 14716
rect 6930 14662 6976 14714
rect 6976 14662 6986 14714
rect 7010 14662 7040 14714
rect 7040 14662 7052 14714
rect 7052 14662 7066 14714
rect 7090 14662 7104 14714
rect 7104 14662 7116 14714
rect 7116 14662 7146 14714
rect 7170 14662 7180 14714
rect 7180 14662 7226 14714
rect 6930 14660 6986 14662
rect 7010 14660 7066 14662
rect 7090 14660 7146 14662
rect 7170 14660 7226 14662
rect 18878 14714 18934 14716
rect 18958 14714 19014 14716
rect 19038 14714 19094 14716
rect 19118 14714 19174 14716
rect 18878 14662 18924 14714
rect 18924 14662 18934 14714
rect 18958 14662 18988 14714
rect 18988 14662 19000 14714
rect 19000 14662 19014 14714
rect 19038 14662 19052 14714
rect 19052 14662 19064 14714
rect 19064 14662 19094 14714
rect 19118 14662 19128 14714
rect 19128 14662 19174 14714
rect 18878 14660 18934 14662
rect 18958 14660 19014 14662
rect 19038 14660 19094 14662
rect 19118 14660 19174 14662
rect 1398 14356 1400 14376
rect 1400 14356 1452 14376
rect 1452 14356 1454 14376
rect 1398 14320 1454 14356
rect 12904 14170 12960 14172
rect 12984 14170 13040 14172
rect 13064 14170 13120 14172
rect 13144 14170 13200 14172
rect 12904 14118 12950 14170
rect 12950 14118 12960 14170
rect 12984 14118 13014 14170
rect 13014 14118 13026 14170
rect 13026 14118 13040 14170
rect 13064 14118 13078 14170
rect 13078 14118 13090 14170
rect 13090 14118 13120 14170
rect 13144 14118 13154 14170
rect 13154 14118 13200 14170
rect 12904 14116 12960 14118
rect 12984 14116 13040 14118
rect 13064 14116 13120 14118
rect 13144 14116 13200 14118
rect 1398 13676 1400 13696
rect 1400 13676 1452 13696
rect 1452 13676 1454 13696
rect 1398 13640 1454 13676
rect 6930 13626 6986 13628
rect 7010 13626 7066 13628
rect 7090 13626 7146 13628
rect 7170 13626 7226 13628
rect 6930 13574 6976 13626
rect 6976 13574 6986 13626
rect 7010 13574 7040 13626
rect 7040 13574 7052 13626
rect 7052 13574 7066 13626
rect 7090 13574 7104 13626
rect 7104 13574 7116 13626
rect 7116 13574 7146 13626
rect 7170 13574 7180 13626
rect 7180 13574 7226 13626
rect 6930 13572 6986 13574
rect 7010 13572 7066 13574
rect 7090 13572 7146 13574
rect 7170 13572 7226 13574
rect 18878 13626 18934 13628
rect 18958 13626 19014 13628
rect 19038 13626 19094 13628
rect 19118 13626 19174 13628
rect 18878 13574 18924 13626
rect 18924 13574 18934 13626
rect 18958 13574 18988 13626
rect 18988 13574 19000 13626
rect 19000 13574 19014 13626
rect 19038 13574 19052 13626
rect 19052 13574 19064 13626
rect 19064 13574 19094 13626
rect 19118 13574 19128 13626
rect 19128 13574 19174 13626
rect 18878 13572 18934 13574
rect 18958 13572 19014 13574
rect 19038 13572 19094 13574
rect 19118 13572 19174 13574
rect 12904 13082 12960 13084
rect 12984 13082 13040 13084
rect 13064 13082 13120 13084
rect 13144 13082 13200 13084
rect 12904 13030 12950 13082
rect 12950 13030 12960 13082
rect 12984 13030 13014 13082
rect 13014 13030 13026 13082
rect 13026 13030 13040 13082
rect 13064 13030 13078 13082
rect 13078 13030 13090 13082
rect 13090 13030 13120 13082
rect 13144 13030 13154 13082
rect 13154 13030 13200 13082
rect 12904 13028 12960 13030
rect 12984 13028 13040 13030
rect 13064 13028 13120 13030
rect 13144 13028 13200 13030
rect 6930 12538 6986 12540
rect 7010 12538 7066 12540
rect 7090 12538 7146 12540
rect 7170 12538 7226 12540
rect 6930 12486 6976 12538
rect 6976 12486 6986 12538
rect 7010 12486 7040 12538
rect 7040 12486 7052 12538
rect 7052 12486 7066 12538
rect 7090 12486 7104 12538
rect 7104 12486 7116 12538
rect 7116 12486 7146 12538
rect 7170 12486 7180 12538
rect 7180 12486 7226 12538
rect 6930 12484 6986 12486
rect 7010 12484 7066 12486
rect 7090 12484 7146 12486
rect 7170 12484 7226 12486
rect 18878 12538 18934 12540
rect 18958 12538 19014 12540
rect 19038 12538 19094 12540
rect 19118 12538 19174 12540
rect 18878 12486 18924 12538
rect 18924 12486 18934 12538
rect 18958 12486 18988 12538
rect 18988 12486 19000 12538
rect 19000 12486 19014 12538
rect 19038 12486 19052 12538
rect 19052 12486 19064 12538
rect 19064 12486 19094 12538
rect 19118 12486 19128 12538
rect 19128 12486 19174 12538
rect 18878 12484 18934 12486
rect 18958 12484 19014 12486
rect 19038 12484 19094 12486
rect 19118 12484 19174 12486
rect 1398 12280 1454 12336
rect 12904 11994 12960 11996
rect 12984 11994 13040 11996
rect 13064 11994 13120 11996
rect 13144 11994 13200 11996
rect 12904 11942 12950 11994
rect 12950 11942 12960 11994
rect 12984 11942 13014 11994
rect 13014 11942 13026 11994
rect 13026 11942 13040 11994
rect 13064 11942 13078 11994
rect 13078 11942 13090 11994
rect 13090 11942 13120 11994
rect 13144 11942 13154 11994
rect 13154 11942 13200 11994
rect 12904 11940 12960 11942
rect 12984 11940 13040 11942
rect 13064 11940 13120 11942
rect 13144 11940 13200 11942
rect 1398 11636 1400 11656
rect 1400 11636 1452 11656
rect 1452 11636 1454 11656
rect 1398 11600 1454 11636
rect 6930 11450 6986 11452
rect 7010 11450 7066 11452
rect 7090 11450 7146 11452
rect 7170 11450 7226 11452
rect 6930 11398 6976 11450
rect 6976 11398 6986 11450
rect 7010 11398 7040 11450
rect 7040 11398 7052 11450
rect 7052 11398 7066 11450
rect 7090 11398 7104 11450
rect 7104 11398 7116 11450
rect 7116 11398 7146 11450
rect 7170 11398 7180 11450
rect 7180 11398 7226 11450
rect 6930 11396 6986 11398
rect 7010 11396 7066 11398
rect 7090 11396 7146 11398
rect 7170 11396 7226 11398
rect 18878 11450 18934 11452
rect 18958 11450 19014 11452
rect 19038 11450 19094 11452
rect 19118 11450 19174 11452
rect 18878 11398 18924 11450
rect 18924 11398 18934 11450
rect 18958 11398 18988 11450
rect 18988 11398 19000 11450
rect 19000 11398 19014 11450
rect 19038 11398 19052 11450
rect 19052 11398 19064 11450
rect 19064 11398 19094 11450
rect 19118 11398 19128 11450
rect 19128 11398 19174 11450
rect 18878 11396 18934 11398
rect 18958 11396 19014 11398
rect 19038 11396 19094 11398
rect 19118 11396 19174 11398
rect 1398 10920 1454 10976
rect 12904 10906 12960 10908
rect 12984 10906 13040 10908
rect 13064 10906 13120 10908
rect 13144 10906 13200 10908
rect 12904 10854 12950 10906
rect 12950 10854 12960 10906
rect 12984 10854 13014 10906
rect 13014 10854 13026 10906
rect 13026 10854 13040 10906
rect 13064 10854 13078 10906
rect 13078 10854 13090 10906
rect 13090 10854 13120 10906
rect 13144 10854 13154 10906
rect 13154 10854 13200 10906
rect 12904 10852 12960 10854
rect 12984 10852 13040 10854
rect 13064 10852 13120 10854
rect 13144 10852 13200 10854
rect 6930 10362 6986 10364
rect 7010 10362 7066 10364
rect 7090 10362 7146 10364
rect 7170 10362 7226 10364
rect 6930 10310 6976 10362
rect 6976 10310 6986 10362
rect 7010 10310 7040 10362
rect 7040 10310 7052 10362
rect 7052 10310 7066 10362
rect 7090 10310 7104 10362
rect 7104 10310 7116 10362
rect 7116 10310 7146 10362
rect 7170 10310 7180 10362
rect 7180 10310 7226 10362
rect 6930 10308 6986 10310
rect 7010 10308 7066 10310
rect 7090 10308 7146 10310
rect 7170 10308 7226 10310
rect 18878 10362 18934 10364
rect 18958 10362 19014 10364
rect 19038 10362 19094 10364
rect 19118 10362 19174 10364
rect 18878 10310 18924 10362
rect 18924 10310 18934 10362
rect 18958 10310 18988 10362
rect 18988 10310 19000 10362
rect 19000 10310 19014 10362
rect 19038 10310 19052 10362
rect 19052 10310 19064 10362
rect 19064 10310 19094 10362
rect 19118 10310 19128 10362
rect 19128 10310 19174 10362
rect 18878 10308 18934 10310
rect 18958 10308 19014 10310
rect 19038 10308 19094 10310
rect 19118 10308 19174 10310
rect 12904 9818 12960 9820
rect 12984 9818 13040 9820
rect 13064 9818 13120 9820
rect 13144 9818 13200 9820
rect 12904 9766 12950 9818
rect 12950 9766 12960 9818
rect 12984 9766 13014 9818
rect 13014 9766 13026 9818
rect 13026 9766 13040 9818
rect 13064 9766 13078 9818
rect 13078 9766 13090 9818
rect 13090 9766 13120 9818
rect 13144 9766 13154 9818
rect 13154 9766 13200 9818
rect 12904 9764 12960 9766
rect 12984 9764 13040 9766
rect 13064 9764 13120 9766
rect 13144 9764 13200 9766
rect 6930 9274 6986 9276
rect 7010 9274 7066 9276
rect 7090 9274 7146 9276
rect 7170 9274 7226 9276
rect 6930 9222 6976 9274
rect 6976 9222 6986 9274
rect 7010 9222 7040 9274
rect 7040 9222 7052 9274
rect 7052 9222 7066 9274
rect 7090 9222 7104 9274
rect 7104 9222 7116 9274
rect 7116 9222 7146 9274
rect 7170 9222 7180 9274
rect 7180 9222 7226 9274
rect 6930 9220 6986 9222
rect 7010 9220 7066 9222
rect 7090 9220 7146 9222
rect 7170 9220 7226 9222
rect 18878 9274 18934 9276
rect 18958 9274 19014 9276
rect 19038 9274 19094 9276
rect 19118 9274 19174 9276
rect 18878 9222 18924 9274
rect 18924 9222 18934 9274
rect 18958 9222 18988 9274
rect 18988 9222 19000 9274
rect 19000 9222 19014 9274
rect 19038 9222 19052 9274
rect 19052 9222 19064 9274
rect 19064 9222 19094 9274
rect 19118 9222 19128 9274
rect 19128 9222 19174 9274
rect 18878 9220 18934 9222
rect 18958 9220 19014 9222
rect 19038 9220 19094 9222
rect 19118 9220 19174 9222
rect 1398 8916 1400 8936
rect 1400 8916 1452 8936
rect 1452 8916 1454 8936
rect 1398 8880 1454 8916
rect 12904 8730 12960 8732
rect 12984 8730 13040 8732
rect 13064 8730 13120 8732
rect 13144 8730 13200 8732
rect 12904 8678 12950 8730
rect 12950 8678 12960 8730
rect 12984 8678 13014 8730
rect 13014 8678 13026 8730
rect 13026 8678 13040 8730
rect 13064 8678 13078 8730
rect 13078 8678 13090 8730
rect 13090 8678 13120 8730
rect 13144 8678 13154 8730
rect 13154 8678 13200 8730
rect 12904 8676 12960 8678
rect 12984 8676 13040 8678
rect 13064 8676 13120 8678
rect 13144 8676 13200 8678
rect 1398 8200 1454 8256
rect 6930 8186 6986 8188
rect 7010 8186 7066 8188
rect 7090 8186 7146 8188
rect 7170 8186 7226 8188
rect 6930 8134 6976 8186
rect 6976 8134 6986 8186
rect 7010 8134 7040 8186
rect 7040 8134 7052 8186
rect 7052 8134 7066 8186
rect 7090 8134 7104 8186
rect 7104 8134 7116 8186
rect 7116 8134 7146 8186
rect 7170 8134 7180 8186
rect 7180 8134 7226 8186
rect 6930 8132 6986 8134
rect 7010 8132 7066 8134
rect 7090 8132 7146 8134
rect 7170 8132 7226 8134
rect 18878 8186 18934 8188
rect 18958 8186 19014 8188
rect 19038 8186 19094 8188
rect 19118 8186 19174 8188
rect 18878 8134 18924 8186
rect 18924 8134 18934 8186
rect 18958 8134 18988 8186
rect 18988 8134 19000 8186
rect 19000 8134 19014 8186
rect 19038 8134 19052 8186
rect 19052 8134 19064 8186
rect 19064 8134 19094 8186
rect 19118 8134 19128 8186
rect 19128 8134 19174 8186
rect 18878 8132 18934 8134
rect 18958 8132 19014 8134
rect 19038 8132 19094 8134
rect 19118 8132 19174 8134
rect 12904 7642 12960 7644
rect 12984 7642 13040 7644
rect 13064 7642 13120 7644
rect 13144 7642 13200 7644
rect 12904 7590 12950 7642
rect 12950 7590 12960 7642
rect 12984 7590 13014 7642
rect 13014 7590 13026 7642
rect 13026 7590 13040 7642
rect 13064 7590 13078 7642
rect 13078 7590 13090 7642
rect 13090 7590 13120 7642
rect 13144 7590 13154 7642
rect 13154 7590 13200 7642
rect 12904 7588 12960 7590
rect 12984 7588 13040 7590
rect 13064 7588 13120 7590
rect 13144 7588 13200 7590
rect 1398 7520 1454 7576
rect 6930 7098 6986 7100
rect 7010 7098 7066 7100
rect 7090 7098 7146 7100
rect 7170 7098 7226 7100
rect 6930 7046 6976 7098
rect 6976 7046 6986 7098
rect 7010 7046 7040 7098
rect 7040 7046 7052 7098
rect 7052 7046 7066 7098
rect 7090 7046 7104 7098
rect 7104 7046 7116 7098
rect 7116 7046 7146 7098
rect 7170 7046 7180 7098
rect 7180 7046 7226 7098
rect 6930 7044 6986 7046
rect 7010 7044 7066 7046
rect 7090 7044 7146 7046
rect 7170 7044 7226 7046
rect 18878 7098 18934 7100
rect 18958 7098 19014 7100
rect 19038 7098 19094 7100
rect 19118 7098 19174 7100
rect 18878 7046 18924 7098
rect 18924 7046 18934 7098
rect 18958 7046 18988 7098
rect 18988 7046 19000 7098
rect 19000 7046 19014 7098
rect 19038 7046 19052 7098
rect 19052 7046 19064 7098
rect 19064 7046 19094 7098
rect 19118 7046 19128 7098
rect 19128 7046 19174 7098
rect 18878 7044 18934 7046
rect 18958 7044 19014 7046
rect 19038 7044 19094 7046
rect 19118 7044 19174 7046
rect 1398 6840 1454 6896
rect 12904 6554 12960 6556
rect 12984 6554 13040 6556
rect 13064 6554 13120 6556
rect 13144 6554 13200 6556
rect 12904 6502 12950 6554
rect 12950 6502 12960 6554
rect 12984 6502 13014 6554
rect 13014 6502 13026 6554
rect 13026 6502 13040 6554
rect 13064 6502 13078 6554
rect 13078 6502 13090 6554
rect 13090 6502 13120 6554
rect 13144 6502 13154 6554
rect 13154 6502 13200 6554
rect 12904 6500 12960 6502
rect 12984 6500 13040 6502
rect 13064 6500 13120 6502
rect 13144 6500 13200 6502
rect 1398 6196 1400 6216
rect 1400 6196 1452 6216
rect 1452 6196 1454 6216
rect 1398 6160 1454 6196
rect 6930 6010 6986 6012
rect 7010 6010 7066 6012
rect 7090 6010 7146 6012
rect 7170 6010 7226 6012
rect 6930 5958 6976 6010
rect 6976 5958 6986 6010
rect 7010 5958 7040 6010
rect 7040 5958 7052 6010
rect 7052 5958 7066 6010
rect 7090 5958 7104 6010
rect 7104 5958 7116 6010
rect 7116 5958 7146 6010
rect 7170 5958 7180 6010
rect 7180 5958 7226 6010
rect 6930 5956 6986 5958
rect 7010 5956 7066 5958
rect 7090 5956 7146 5958
rect 7170 5956 7226 5958
rect 18878 6010 18934 6012
rect 18958 6010 19014 6012
rect 19038 6010 19094 6012
rect 19118 6010 19174 6012
rect 18878 5958 18924 6010
rect 18924 5958 18934 6010
rect 18958 5958 18988 6010
rect 18988 5958 19000 6010
rect 19000 5958 19014 6010
rect 19038 5958 19052 6010
rect 19052 5958 19064 6010
rect 19064 5958 19094 6010
rect 19118 5958 19128 6010
rect 19128 5958 19174 6010
rect 18878 5956 18934 5958
rect 18958 5956 19014 5958
rect 19038 5956 19094 5958
rect 19118 5956 19174 5958
rect 1398 5480 1454 5536
rect 12904 5466 12960 5468
rect 12984 5466 13040 5468
rect 13064 5466 13120 5468
rect 13144 5466 13200 5468
rect 12904 5414 12950 5466
rect 12950 5414 12960 5466
rect 12984 5414 13014 5466
rect 13014 5414 13026 5466
rect 13026 5414 13040 5466
rect 13064 5414 13078 5466
rect 13078 5414 13090 5466
rect 13090 5414 13120 5466
rect 13144 5414 13154 5466
rect 13154 5414 13200 5466
rect 12904 5412 12960 5414
rect 12984 5412 13040 5414
rect 13064 5412 13120 5414
rect 13144 5412 13200 5414
rect 6930 4922 6986 4924
rect 7010 4922 7066 4924
rect 7090 4922 7146 4924
rect 7170 4922 7226 4924
rect 6930 4870 6976 4922
rect 6976 4870 6986 4922
rect 7010 4870 7040 4922
rect 7040 4870 7052 4922
rect 7052 4870 7066 4922
rect 7090 4870 7104 4922
rect 7104 4870 7116 4922
rect 7116 4870 7146 4922
rect 7170 4870 7180 4922
rect 7180 4870 7226 4922
rect 6930 4868 6986 4870
rect 7010 4868 7066 4870
rect 7090 4868 7146 4870
rect 7170 4868 7226 4870
rect 18878 4922 18934 4924
rect 18958 4922 19014 4924
rect 19038 4922 19094 4924
rect 19118 4922 19174 4924
rect 18878 4870 18924 4922
rect 18924 4870 18934 4922
rect 18958 4870 18988 4922
rect 18988 4870 19000 4922
rect 19000 4870 19014 4922
rect 19038 4870 19052 4922
rect 19052 4870 19064 4922
rect 19064 4870 19094 4922
rect 19118 4870 19128 4922
rect 19128 4870 19174 4922
rect 18878 4868 18934 4870
rect 18958 4868 19014 4870
rect 19038 4868 19094 4870
rect 19118 4868 19174 4870
rect 1398 4800 1454 4856
rect 12904 4378 12960 4380
rect 12984 4378 13040 4380
rect 13064 4378 13120 4380
rect 13144 4378 13200 4380
rect 12904 4326 12950 4378
rect 12950 4326 12960 4378
rect 12984 4326 13014 4378
rect 13014 4326 13026 4378
rect 13026 4326 13040 4378
rect 13064 4326 13078 4378
rect 13078 4326 13090 4378
rect 13090 4326 13120 4378
rect 13144 4326 13154 4378
rect 13154 4326 13200 4378
rect 12904 4324 12960 4326
rect 12984 4324 13040 4326
rect 13064 4324 13120 4326
rect 13144 4324 13200 4326
rect 1398 3476 1400 3496
rect 1400 3476 1452 3496
rect 1452 3476 1454 3496
rect 1398 3440 1454 3476
rect 2778 2080 2834 2136
rect 6930 3834 6986 3836
rect 7010 3834 7066 3836
rect 7090 3834 7146 3836
rect 7170 3834 7226 3836
rect 6930 3782 6976 3834
rect 6976 3782 6986 3834
rect 7010 3782 7040 3834
rect 7040 3782 7052 3834
rect 7052 3782 7066 3834
rect 7090 3782 7104 3834
rect 7104 3782 7116 3834
rect 7116 3782 7146 3834
rect 7170 3782 7180 3834
rect 7180 3782 7226 3834
rect 6930 3780 6986 3782
rect 7010 3780 7066 3782
rect 7090 3780 7146 3782
rect 7170 3780 7226 3782
rect 18878 3834 18934 3836
rect 18958 3834 19014 3836
rect 19038 3834 19094 3836
rect 19118 3834 19174 3836
rect 18878 3782 18924 3834
rect 18924 3782 18934 3834
rect 18958 3782 18988 3834
rect 18988 3782 19000 3834
rect 19000 3782 19014 3834
rect 19038 3782 19052 3834
rect 19052 3782 19064 3834
rect 19064 3782 19094 3834
rect 19118 3782 19128 3834
rect 19128 3782 19174 3834
rect 18878 3780 18934 3782
rect 18958 3780 19014 3782
rect 19038 3780 19094 3782
rect 19118 3780 19174 3782
rect 2870 1400 2926 1456
rect 12904 3290 12960 3292
rect 12984 3290 13040 3292
rect 13064 3290 13120 3292
rect 13144 3290 13200 3292
rect 12904 3238 12950 3290
rect 12950 3238 12960 3290
rect 12984 3238 13014 3290
rect 13014 3238 13026 3290
rect 13026 3238 13040 3290
rect 13064 3238 13078 3290
rect 13078 3238 13090 3290
rect 13090 3238 13120 3290
rect 13144 3238 13154 3290
rect 13154 3238 13200 3290
rect 12904 3236 12960 3238
rect 12984 3236 13040 3238
rect 13064 3236 13120 3238
rect 13144 3236 13200 3238
rect 2962 720 3018 776
rect 2962 40 3018 96
rect 6930 2746 6986 2748
rect 7010 2746 7066 2748
rect 7090 2746 7146 2748
rect 7170 2746 7226 2748
rect 6930 2694 6976 2746
rect 6976 2694 6986 2746
rect 7010 2694 7040 2746
rect 7040 2694 7052 2746
rect 7052 2694 7066 2746
rect 7090 2694 7104 2746
rect 7104 2694 7116 2746
rect 7116 2694 7146 2746
rect 7170 2694 7180 2746
rect 7180 2694 7226 2746
rect 6930 2692 6986 2694
rect 7010 2692 7066 2694
rect 7090 2692 7146 2694
rect 7170 2692 7226 2694
rect 12904 2202 12960 2204
rect 12984 2202 13040 2204
rect 13064 2202 13120 2204
rect 13144 2202 13200 2204
rect 12904 2150 12950 2202
rect 12950 2150 12960 2202
rect 12984 2150 13014 2202
rect 13014 2150 13026 2202
rect 13026 2150 13040 2202
rect 13064 2150 13078 2202
rect 13078 2150 13090 2202
rect 13090 2150 13120 2202
rect 13144 2150 13154 2202
rect 13154 2150 13200 2202
rect 12904 2148 12960 2150
rect 12984 2148 13040 2150
rect 13064 2148 13120 2150
rect 13144 2148 13200 2150
rect 18878 2746 18934 2748
rect 18958 2746 19014 2748
rect 19038 2746 19094 2748
rect 19118 2746 19174 2748
rect 18878 2694 18924 2746
rect 18924 2694 18934 2746
rect 18958 2694 18988 2746
rect 18988 2694 19000 2746
rect 19000 2694 19014 2746
rect 19038 2694 19052 2746
rect 19052 2694 19064 2746
rect 19064 2694 19094 2746
rect 19118 2694 19128 2746
rect 19128 2694 19174 2746
rect 18878 2692 18934 2694
rect 18958 2692 19014 2694
rect 19038 2692 19094 2694
rect 19118 2692 19174 2694
rect 30826 14714 30882 14716
rect 30906 14714 30962 14716
rect 30986 14714 31042 14716
rect 31066 14714 31122 14716
rect 30826 14662 30872 14714
rect 30872 14662 30882 14714
rect 30906 14662 30936 14714
rect 30936 14662 30948 14714
rect 30948 14662 30962 14714
rect 30986 14662 31000 14714
rect 31000 14662 31012 14714
rect 31012 14662 31042 14714
rect 31066 14662 31076 14714
rect 31076 14662 31122 14714
rect 30826 14660 30882 14662
rect 30906 14660 30962 14662
rect 30986 14660 31042 14662
rect 31066 14660 31122 14662
rect 42774 14714 42830 14716
rect 42854 14714 42910 14716
rect 42934 14714 42990 14716
rect 43014 14714 43070 14716
rect 42774 14662 42820 14714
rect 42820 14662 42830 14714
rect 42854 14662 42884 14714
rect 42884 14662 42896 14714
rect 42896 14662 42910 14714
rect 42934 14662 42948 14714
rect 42948 14662 42960 14714
rect 42960 14662 42990 14714
rect 43014 14662 43024 14714
rect 43024 14662 43070 14714
rect 42774 14660 42830 14662
rect 42854 14660 42910 14662
rect 42934 14660 42990 14662
rect 43014 14660 43070 14662
rect 24852 14170 24908 14172
rect 24932 14170 24988 14172
rect 25012 14170 25068 14172
rect 25092 14170 25148 14172
rect 24852 14118 24898 14170
rect 24898 14118 24908 14170
rect 24932 14118 24962 14170
rect 24962 14118 24974 14170
rect 24974 14118 24988 14170
rect 25012 14118 25026 14170
rect 25026 14118 25038 14170
rect 25038 14118 25068 14170
rect 25092 14118 25102 14170
rect 25102 14118 25148 14170
rect 24852 14116 24908 14118
rect 24932 14116 24988 14118
rect 25012 14116 25068 14118
rect 25092 14116 25148 14118
rect 36800 14170 36856 14172
rect 36880 14170 36936 14172
rect 36960 14170 37016 14172
rect 37040 14170 37096 14172
rect 36800 14118 36846 14170
rect 36846 14118 36856 14170
rect 36880 14118 36910 14170
rect 36910 14118 36922 14170
rect 36922 14118 36936 14170
rect 36960 14118 36974 14170
rect 36974 14118 36986 14170
rect 36986 14118 37016 14170
rect 37040 14118 37050 14170
rect 37050 14118 37096 14170
rect 36800 14116 36856 14118
rect 36880 14116 36936 14118
rect 36960 14116 37016 14118
rect 37040 14116 37096 14118
rect 24852 13082 24908 13084
rect 24932 13082 24988 13084
rect 25012 13082 25068 13084
rect 25092 13082 25148 13084
rect 24852 13030 24898 13082
rect 24898 13030 24908 13082
rect 24932 13030 24962 13082
rect 24962 13030 24974 13082
rect 24974 13030 24988 13082
rect 25012 13030 25026 13082
rect 25026 13030 25038 13082
rect 25038 13030 25068 13082
rect 25092 13030 25102 13082
rect 25102 13030 25148 13082
rect 24852 13028 24908 13030
rect 24932 13028 24988 13030
rect 25012 13028 25068 13030
rect 25092 13028 25148 13030
rect 30826 13626 30882 13628
rect 30906 13626 30962 13628
rect 30986 13626 31042 13628
rect 31066 13626 31122 13628
rect 30826 13574 30872 13626
rect 30872 13574 30882 13626
rect 30906 13574 30936 13626
rect 30936 13574 30948 13626
rect 30948 13574 30962 13626
rect 30986 13574 31000 13626
rect 31000 13574 31012 13626
rect 31012 13574 31042 13626
rect 31066 13574 31076 13626
rect 31076 13574 31122 13626
rect 30826 13572 30882 13574
rect 30906 13572 30962 13574
rect 30986 13572 31042 13574
rect 31066 13572 31122 13574
rect 36800 13082 36856 13084
rect 36880 13082 36936 13084
rect 36960 13082 37016 13084
rect 37040 13082 37096 13084
rect 36800 13030 36846 13082
rect 36846 13030 36856 13082
rect 36880 13030 36910 13082
rect 36910 13030 36922 13082
rect 36922 13030 36936 13082
rect 36960 13030 36974 13082
rect 36974 13030 36986 13082
rect 36986 13030 37016 13082
rect 37040 13030 37050 13082
rect 37050 13030 37096 13082
rect 36800 13028 36856 13030
rect 36880 13028 36936 13030
rect 36960 13028 37016 13030
rect 37040 13028 37096 13030
rect 42774 13626 42830 13628
rect 42854 13626 42910 13628
rect 42934 13626 42990 13628
rect 43014 13626 43070 13628
rect 42774 13574 42820 13626
rect 42820 13574 42830 13626
rect 42854 13574 42884 13626
rect 42884 13574 42896 13626
rect 42896 13574 42910 13626
rect 42934 13574 42948 13626
rect 42948 13574 42960 13626
rect 42960 13574 42990 13626
rect 43014 13574 43024 13626
rect 43024 13574 43070 13626
rect 42774 13572 42830 13574
rect 42854 13572 42910 13574
rect 42934 13572 42990 13574
rect 43014 13572 43070 13574
rect 45558 13776 45614 13832
rect 30826 12538 30882 12540
rect 30906 12538 30962 12540
rect 30986 12538 31042 12540
rect 31066 12538 31122 12540
rect 30826 12486 30872 12538
rect 30872 12486 30882 12538
rect 30906 12486 30936 12538
rect 30936 12486 30948 12538
rect 30948 12486 30962 12538
rect 30986 12486 31000 12538
rect 31000 12486 31012 12538
rect 31012 12486 31042 12538
rect 31066 12486 31076 12538
rect 31076 12486 31122 12538
rect 30826 12484 30882 12486
rect 30906 12484 30962 12486
rect 30986 12484 31042 12486
rect 31066 12484 31122 12486
rect 42774 12538 42830 12540
rect 42854 12538 42910 12540
rect 42934 12538 42990 12540
rect 43014 12538 43070 12540
rect 42774 12486 42820 12538
rect 42820 12486 42830 12538
rect 42854 12486 42884 12538
rect 42884 12486 42896 12538
rect 42896 12486 42910 12538
rect 42934 12486 42948 12538
rect 42948 12486 42960 12538
rect 42960 12486 42990 12538
rect 43014 12486 43024 12538
rect 43024 12486 43070 12538
rect 42774 12484 42830 12486
rect 42854 12484 42910 12486
rect 42934 12484 42990 12486
rect 43014 12484 43070 12486
rect 24852 11994 24908 11996
rect 24932 11994 24988 11996
rect 25012 11994 25068 11996
rect 25092 11994 25148 11996
rect 24852 11942 24898 11994
rect 24898 11942 24908 11994
rect 24932 11942 24962 11994
rect 24962 11942 24974 11994
rect 24974 11942 24988 11994
rect 25012 11942 25026 11994
rect 25026 11942 25038 11994
rect 25038 11942 25068 11994
rect 25092 11942 25102 11994
rect 25102 11942 25148 11994
rect 24852 11940 24908 11942
rect 24932 11940 24988 11942
rect 25012 11940 25068 11942
rect 25092 11940 25148 11942
rect 36800 11994 36856 11996
rect 36880 11994 36936 11996
rect 36960 11994 37016 11996
rect 37040 11994 37096 11996
rect 36800 11942 36846 11994
rect 36846 11942 36856 11994
rect 36880 11942 36910 11994
rect 36910 11942 36922 11994
rect 36922 11942 36936 11994
rect 36960 11942 36974 11994
rect 36974 11942 36986 11994
rect 36986 11942 37016 11994
rect 37040 11942 37050 11994
rect 37050 11942 37096 11994
rect 36800 11940 36856 11942
rect 36880 11940 36936 11942
rect 36960 11940 37016 11942
rect 37040 11940 37096 11942
rect 30826 11450 30882 11452
rect 30906 11450 30962 11452
rect 30986 11450 31042 11452
rect 31066 11450 31122 11452
rect 30826 11398 30872 11450
rect 30872 11398 30882 11450
rect 30906 11398 30936 11450
rect 30936 11398 30948 11450
rect 30948 11398 30962 11450
rect 30986 11398 31000 11450
rect 31000 11398 31012 11450
rect 31012 11398 31042 11450
rect 31066 11398 31076 11450
rect 31076 11398 31122 11450
rect 30826 11396 30882 11398
rect 30906 11396 30962 11398
rect 30986 11396 31042 11398
rect 31066 11396 31122 11398
rect 42774 11450 42830 11452
rect 42854 11450 42910 11452
rect 42934 11450 42990 11452
rect 43014 11450 43070 11452
rect 42774 11398 42820 11450
rect 42820 11398 42830 11450
rect 42854 11398 42884 11450
rect 42884 11398 42896 11450
rect 42896 11398 42910 11450
rect 42934 11398 42948 11450
rect 42948 11398 42960 11450
rect 42960 11398 42990 11450
rect 43014 11398 43024 11450
rect 43024 11398 43070 11450
rect 42774 11396 42830 11398
rect 42854 11396 42910 11398
rect 42934 11396 42990 11398
rect 43014 11396 43070 11398
rect 24852 10906 24908 10908
rect 24932 10906 24988 10908
rect 25012 10906 25068 10908
rect 25092 10906 25148 10908
rect 24852 10854 24898 10906
rect 24898 10854 24908 10906
rect 24932 10854 24962 10906
rect 24962 10854 24974 10906
rect 24974 10854 24988 10906
rect 25012 10854 25026 10906
rect 25026 10854 25038 10906
rect 25038 10854 25068 10906
rect 25092 10854 25102 10906
rect 25102 10854 25148 10906
rect 24852 10852 24908 10854
rect 24932 10852 24988 10854
rect 25012 10852 25068 10854
rect 25092 10852 25148 10854
rect 36800 10906 36856 10908
rect 36880 10906 36936 10908
rect 36960 10906 37016 10908
rect 37040 10906 37096 10908
rect 36800 10854 36846 10906
rect 36846 10854 36856 10906
rect 36880 10854 36910 10906
rect 36910 10854 36922 10906
rect 36922 10854 36936 10906
rect 36960 10854 36974 10906
rect 36974 10854 36986 10906
rect 36986 10854 37016 10906
rect 37040 10854 37050 10906
rect 37050 10854 37096 10906
rect 36800 10852 36856 10854
rect 36880 10852 36936 10854
rect 36960 10852 37016 10854
rect 37040 10852 37096 10854
rect 30826 10362 30882 10364
rect 30906 10362 30962 10364
rect 30986 10362 31042 10364
rect 31066 10362 31122 10364
rect 30826 10310 30872 10362
rect 30872 10310 30882 10362
rect 30906 10310 30936 10362
rect 30936 10310 30948 10362
rect 30948 10310 30962 10362
rect 30986 10310 31000 10362
rect 31000 10310 31012 10362
rect 31012 10310 31042 10362
rect 31066 10310 31076 10362
rect 31076 10310 31122 10362
rect 30826 10308 30882 10310
rect 30906 10308 30962 10310
rect 30986 10308 31042 10310
rect 31066 10308 31122 10310
rect 42774 10362 42830 10364
rect 42854 10362 42910 10364
rect 42934 10362 42990 10364
rect 43014 10362 43070 10364
rect 42774 10310 42820 10362
rect 42820 10310 42830 10362
rect 42854 10310 42884 10362
rect 42884 10310 42896 10362
rect 42896 10310 42910 10362
rect 42934 10310 42948 10362
rect 42948 10310 42960 10362
rect 42960 10310 42990 10362
rect 43014 10310 43024 10362
rect 43024 10310 43070 10362
rect 42774 10308 42830 10310
rect 42854 10308 42910 10310
rect 42934 10308 42990 10310
rect 43014 10308 43070 10310
rect 24852 9818 24908 9820
rect 24932 9818 24988 9820
rect 25012 9818 25068 9820
rect 25092 9818 25148 9820
rect 24852 9766 24898 9818
rect 24898 9766 24908 9818
rect 24932 9766 24962 9818
rect 24962 9766 24974 9818
rect 24974 9766 24988 9818
rect 25012 9766 25026 9818
rect 25026 9766 25038 9818
rect 25038 9766 25068 9818
rect 25092 9766 25102 9818
rect 25102 9766 25148 9818
rect 24852 9764 24908 9766
rect 24932 9764 24988 9766
rect 25012 9764 25068 9766
rect 25092 9764 25148 9766
rect 36800 9818 36856 9820
rect 36880 9818 36936 9820
rect 36960 9818 37016 9820
rect 37040 9818 37096 9820
rect 36800 9766 36846 9818
rect 36846 9766 36856 9818
rect 36880 9766 36910 9818
rect 36910 9766 36922 9818
rect 36922 9766 36936 9818
rect 36960 9766 36974 9818
rect 36974 9766 36986 9818
rect 36986 9766 37016 9818
rect 37040 9766 37050 9818
rect 37050 9766 37096 9818
rect 36800 9764 36856 9766
rect 36880 9764 36936 9766
rect 36960 9764 37016 9766
rect 37040 9764 37096 9766
rect 30826 9274 30882 9276
rect 30906 9274 30962 9276
rect 30986 9274 31042 9276
rect 31066 9274 31122 9276
rect 30826 9222 30872 9274
rect 30872 9222 30882 9274
rect 30906 9222 30936 9274
rect 30936 9222 30948 9274
rect 30948 9222 30962 9274
rect 30986 9222 31000 9274
rect 31000 9222 31012 9274
rect 31012 9222 31042 9274
rect 31066 9222 31076 9274
rect 31076 9222 31122 9274
rect 30826 9220 30882 9222
rect 30906 9220 30962 9222
rect 30986 9220 31042 9222
rect 31066 9220 31122 9222
rect 42774 9274 42830 9276
rect 42854 9274 42910 9276
rect 42934 9274 42990 9276
rect 43014 9274 43070 9276
rect 42774 9222 42820 9274
rect 42820 9222 42830 9274
rect 42854 9222 42884 9274
rect 42884 9222 42896 9274
rect 42896 9222 42910 9274
rect 42934 9222 42948 9274
rect 42948 9222 42960 9274
rect 42960 9222 42990 9274
rect 43014 9222 43024 9274
rect 43024 9222 43070 9274
rect 42774 9220 42830 9222
rect 42854 9220 42910 9222
rect 42934 9220 42990 9222
rect 43014 9220 43070 9222
rect 24852 8730 24908 8732
rect 24932 8730 24988 8732
rect 25012 8730 25068 8732
rect 25092 8730 25148 8732
rect 24852 8678 24898 8730
rect 24898 8678 24908 8730
rect 24932 8678 24962 8730
rect 24962 8678 24974 8730
rect 24974 8678 24988 8730
rect 25012 8678 25026 8730
rect 25026 8678 25038 8730
rect 25038 8678 25068 8730
rect 25092 8678 25102 8730
rect 25102 8678 25148 8730
rect 24852 8676 24908 8678
rect 24932 8676 24988 8678
rect 25012 8676 25068 8678
rect 25092 8676 25148 8678
rect 36800 8730 36856 8732
rect 36880 8730 36936 8732
rect 36960 8730 37016 8732
rect 37040 8730 37096 8732
rect 36800 8678 36846 8730
rect 36846 8678 36856 8730
rect 36880 8678 36910 8730
rect 36910 8678 36922 8730
rect 36922 8678 36936 8730
rect 36960 8678 36974 8730
rect 36974 8678 36986 8730
rect 36986 8678 37016 8730
rect 37040 8678 37050 8730
rect 37050 8678 37096 8730
rect 36800 8676 36856 8678
rect 36880 8676 36936 8678
rect 36960 8676 37016 8678
rect 37040 8676 37096 8678
rect 30826 8186 30882 8188
rect 30906 8186 30962 8188
rect 30986 8186 31042 8188
rect 31066 8186 31122 8188
rect 30826 8134 30872 8186
rect 30872 8134 30882 8186
rect 30906 8134 30936 8186
rect 30936 8134 30948 8186
rect 30948 8134 30962 8186
rect 30986 8134 31000 8186
rect 31000 8134 31012 8186
rect 31012 8134 31042 8186
rect 31066 8134 31076 8186
rect 31076 8134 31122 8186
rect 30826 8132 30882 8134
rect 30906 8132 30962 8134
rect 30986 8132 31042 8134
rect 31066 8132 31122 8134
rect 42774 8186 42830 8188
rect 42854 8186 42910 8188
rect 42934 8186 42990 8188
rect 43014 8186 43070 8188
rect 42774 8134 42820 8186
rect 42820 8134 42830 8186
rect 42854 8134 42884 8186
rect 42884 8134 42896 8186
rect 42896 8134 42910 8186
rect 42934 8134 42948 8186
rect 42948 8134 42960 8186
rect 42960 8134 42990 8186
rect 43014 8134 43024 8186
rect 43024 8134 43070 8186
rect 42774 8132 42830 8134
rect 42854 8132 42910 8134
rect 42934 8132 42990 8134
rect 43014 8132 43070 8134
rect 24852 7642 24908 7644
rect 24932 7642 24988 7644
rect 25012 7642 25068 7644
rect 25092 7642 25148 7644
rect 24852 7590 24898 7642
rect 24898 7590 24908 7642
rect 24932 7590 24962 7642
rect 24962 7590 24974 7642
rect 24974 7590 24988 7642
rect 25012 7590 25026 7642
rect 25026 7590 25038 7642
rect 25038 7590 25068 7642
rect 25092 7590 25102 7642
rect 25102 7590 25148 7642
rect 24852 7588 24908 7590
rect 24932 7588 24988 7590
rect 25012 7588 25068 7590
rect 25092 7588 25148 7590
rect 36800 7642 36856 7644
rect 36880 7642 36936 7644
rect 36960 7642 37016 7644
rect 37040 7642 37096 7644
rect 36800 7590 36846 7642
rect 36846 7590 36856 7642
rect 36880 7590 36910 7642
rect 36910 7590 36922 7642
rect 36922 7590 36936 7642
rect 36960 7590 36974 7642
rect 36974 7590 36986 7642
rect 36986 7590 37016 7642
rect 37040 7590 37050 7642
rect 37050 7590 37096 7642
rect 36800 7588 36856 7590
rect 36880 7588 36936 7590
rect 36960 7588 37016 7590
rect 37040 7588 37096 7590
rect 30826 7098 30882 7100
rect 30906 7098 30962 7100
rect 30986 7098 31042 7100
rect 31066 7098 31122 7100
rect 30826 7046 30872 7098
rect 30872 7046 30882 7098
rect 30906 7046 30936 7098
rect 30936 7046 30948 7098
rect 30948 7046 30962 7098
rect 30986 7046 31000 7098
rect 31000 7046 31012 7098
rect 31012 7046 31042 7098
rect 31066 7046 31076 7098
rect 31076 7046 31122 7098
rect 30826 7044 30882 7046
rect 30906 7044 30962 7046
rect 30986 7044 31042 7046
rect 31066 7044 31122 7046
rect 42774 7098 42830 7100
rect 42854 7098 42910 7100
rect 42934 7098 42990 7100
rect 43014 7098 43070 7100
rect 42774 7046 42820 7098
rect 42820 7046 42830 7098
rect 42854 7046 42884 7098
rect 42884 7046 42896 7098
rect 42896 7046 42910 7098
rect 42934 7046 42948 7098
rect 42948 7046 42960 7098
rect 42960 7046 42990 7098
rect 43014 7046 43024 7098
rect 43024 7046 43070 7098
rect 42774 7044 42830 7046
rect 42854 7044 42910 7046
rect 42934 7044 42990 7046
rect 43014 7044 43070 7046
rect 24852 6554 24908 6556
rect 24932 6554 24988 6556
rect 25012 6554 25068 6556
rect 25092 6554 25148 6556
rect 24852 6502 24898 6554
rect 24898 6502 24908 6554
rect 24932 6502 24962 6554
rect 24962 6502 24974 6554
rect 24974 6502 24988 6554
rect 25012 6502 25026 6554
rect 25026 6502 25038 6554
rect 25038 6502 25068 6554
rect 25092 6502 25102 6554
rect 25102 6502 25148 6554
rect 24852 6500 24908 6502
rect 24932 6500 24988 6502
rect 25012 6500 25068 6502
rect 25092 6500 25148 6502
rect 36800 6554 36856 6556
rect 36880 6554 36936 6556
rect 36960 6554 37016 6556
rect 37040 6554 37096 6556
rect 36800 6502 36846 6554
rect 36846 6502 36856 6554
rect 36880 6502 36910 6554
rect 36910 6502 36922 6554
rect 36922 6502 36936 6554
rect 36960 6502 36974 6554
rect 36974 6502 36986 6554
rect 36986 6502 37016 6554
rect 37040 6502 37050 6554
rect 37050 6502 37096 6554
rect 36800 6500 36856 6502
rect 36880 6500 36936 6502
rect 36960 6500 37016 6502
rect 37040 6500 37096 6502
rect 30826 6010 30882 6012
rect 30906 6010 30962 6012
rect 30986 6010 31042 6012
rect 31066 6010 31122 6012
rect 30826 5958 30872 6010
rect 30872 5958 30882 6010
rect 30906 5958 30936 6010
rect 30936 5958 30948 6010
rect 30948 5958 30962 6010
rect 30986 5958 31000 6010
rect 31000 5958 31012 6010
rect 31012 5958 31042 6010
rect 31066 5958 31076 6010
rect 31076 5958 31122 6010
rect 30826 5956 30882 5958
rect 30906 5956 30962 5958
rect 30986 5956 31042 5958
rect 31066 5956 31122 5958
rect 42774 6010 42830 6012
rect 42854 6010 42910 6012
rect 42934 6010 42990 6012
rect 43014 6010 43070 6012
rect 42774 5958 42820 6010
rect 42820 5958 42830 6010
rect 42854 5958 42884 6010
rect 42884 5958 42896 6010
rect 42896 5958 42910 6010
rect 42934 5958 42948 6010
rect 42948 5958 42960 6010
rect 42960 5958 42990 6010
rect 43014 5958 43024 6010
rect 43024 5958 43070 6010
rect 42774 5956 42830 5958
rect 42854 5956 42910 5958
rect 42934 5956 42990 5958
rect 43014 5956 43070 5958
rect 24852 5466 24908 5468
rect 24932 5466 24988 5468
rect 25012 5466 25068 5468
rect 25092 5466 25148 5468
rect 24852 5414 24898 5466
rect 24898 5414 24908 5466
rect 24932 5414 24962 5466
rect 24962 5414 24974 5466
rect 24974 5414 24988 5466
rect 25012 5414 25026 5466
rect 25026 5414 25038 5466
rect 25038 5414 25068 5466
rect 25092 5414 25102 5466
rect 25102 5414 25148 5466
rect 24852 5412 24908 5414
rect 24932 5412 24988 5414
rect 25012 5412 25068 5414
rect 25092 5412 25148 5414
rect 36800 5466 36856 5468
rect 36880 5466 36936 5468
rect 36960 5466 37016 5468
rect 37040 5466 37096 5468
rect 36800 5414 36846 5466
rect 36846 5414 36856 5466
rect 36880 5414 36910 5466
rect 36910 5414 36922 5466
rect 36922 5414 36936 5466
rect 36960 5414 36974 5466
rect 36974 5414 36986 5466
rect 36986 5414 37016 5466
rect 37040 5414 37050 5466
rect 37050 5414 37096 5466
rect 36800 5412 36856 5414
rect 36880 5412 36936 5414
rect 36960 5412 37016 5414
rect 37040 5412 37096 5414
rect 30826 4922 30882 4924
rect 30906 4922 30962 4924
rect 30986 4922 31042 4924
rect 31066 4922 31122 4924
rect 30826 4870 30872 4922
rect 30872 4870 30882 4922
rect 30906 4870 30936 4922
rect 30936 4870 30948 4922
rect 30948 4870 30962 4922
rect 30986 4870 31000 4922
rect 31000 4870 31012 4922
rect 31012 4870 31042 4922
rect 31066 4870 31076 4922
rect 31076 4870 31122 4922
rect 30826 4868 30882 4870
rect 30906 4868 30962 4870
rect 30986 4868 31042 4870
rect 31066 4868 31122 4870
rect 42774 4922 42830 4924
rect 42854 4922 42910 4924
rect 42934 4922 42990 4924
rect 43014 4922 43070 4924
rect 42774 4870 42820 4922
rect 42820 4870 42830 4922
rect 42854 4870 42884 4922
rect 42884 4870 42896 4922
rect 42896 4870 42910 4922
rect 42934 4870 42948 4922
rect 42948 4870 42960 4922
rect 42960 4870 42990 4922
rect 43014 4870 43024 4922
rect 43024 4870 43070 4922
rect 42774 4868 42830 4870
rect 42854 4868 42910 4870
rect 42934 4868 42990 4870
rect 43014 4868 43070 4870
rect 24852 4378 24908 4380
rect 24932 4378 24988 4380
rect 25012 4378 25068 4380
rect 25092 4378 25148 4380
rect 24852 4326 24898 4378
rect 24898 4326 24908 4378
rect 24932 4326 24962 4378
rect 24962 4326 24974 4378
rect 24974 4326 24988 4378
rect 25012 4326 25026 4378
rect 25026 4326 25038 4378
rect 25038 4326 25068 4378
rect 25092 4326 25102 4378
rect 25102 4326 25148 4378
rect 24852 4324 24908 4326
rect 24932 4324 24988 4326
rect 25012 4324 25068 4326
rect 25092 4324 25148 4326
rect 36800 4378 36856 4380
rect 36880 4378 36936 4380
rect 36960 4378 37016 4380
rect 37040 4378 37096 4380
rect 36800 4326 36846 4378
rect 36846 4326 36856 4378
rect 36880 4326 36910 4378
rect 36910 4326 36922 4378
rect 36922 4326 36936 4378
rect 36960 4326 36974 4378
rect 36974 4326 36986 4378
rect 36986 4326 37016 4378
rect 37040 4326 37050 4378
rect 37050 4326 37096 4378
rect 36800 4324 36856 4326
rect 36880 4324 36936 4326
rect 36960 4324 37016 4326
rect 37040 4324 37096 4326
rect 30826 3834 30882 3836
rect 30906 3834 30962 3836
rect 30986 3834 31042 3836
rect 31066 3834 31122 3836
rect 30826 3782 30872 3834
rect 30872 3782 30882 3834
rect 30906 3782 30936 3834
rect 30936 3782 30948 3834
rect 30948 3782 30962 3834
rect 30986 3782 31000 3834
rect 31000 3782 31012 3834
rect 31012 3782 31042 3834
rect 31066 3782 31076 3834
rect 31076 3782 31122 3834
rect 30826 3780 30882 3782
rect 30906 3780 30962 3782
rect 30986 3780 31042 3782
rect 31066 3780 31122 3782
rect 42774 3834 42830 3836
rect 42854 3834 42910 3836
rect 42934 3834 42990 3836
rect 43014 3834 43070 3836
rect 42774 3782 42820 3834
rect 42820 3782 42830 3834
rect 42854 3782 42884 3834
rect 42884 3782 42896 3834
rect 42896 3782 42910 3834
rect 42934 3782 42948 3834
rect 42948 3782 42960 3834
rect 42960 3782 42990 3834
rect 43014 3782 43024 3834
rect 43024 3782 43070 3834
rect 42774 3780 42830 3782
rect 42854 3780 42910 3782
rect 42934 3780 42990 3782
rect 43014 3780 43070 3782
rect 24852 3290 24908 3292
rect 24932 3290 24988 3292
rect 25012 3290 25068 3292
rect 25092 3290 25148 3292
rect 24852 3238 24898 3290
rect 24898 3238 24908 3290
rect 24932 3238 24962 3290
rect 24962 3238 24974 3290
rect 24974 3238 24988 3290
rect 25012 3238 25026 3290
rect 25026 3238 25038 3290
rect 25038 3238 25068 3290
rect 25092 3238 25102 3290
rect 25102 3238 25148 3290
rect 24852 3236 24908 3238
rect 24932 3236 24988 3238
rect 25012 3236 25068 3238
rect 25092 3236 25148 3238
rect 36800 3290 36856 3292
rect 36880 3290 36936 3292
rect 36960 3290 37016 3292
rect 37040 3290 37096 3292
rect 36800 3238 36846 3290
rect 36846 3238 36856 3290
rect 36880 3238 36910 3290
rect 36910 3238 36922 3290
rect 36922 3238 36936 3290
rect 36960 3238 36974 3290
rect 36974 3238 36986 3290
rect 36986 3238 37016 3290
rect 37040 3238 37050 3290
rect 37050 3238 37096 3290
rect 36800 3236 36856 3238
rect 36880 3236 36936 3238
rect 36960 3236 37016 3238
rect 37040 3236 37096 3238
rect 48134 26288 48190 26344
rect 48226 25472 48282 25528
rect 48134 24928 48190 24984
rect 48134 23568 48190 23624
rect 48226 23432 48282 23488
rect 48226 22208 48282 22264
rect 48134 22072 48190 22128
rect 48134 20712 48190 20768
rect 48226 19352 48282 19408
rect 48134 18128 48190 18184
rect 48226 17992 48282 18048
rect 48226 16768 48282 16824
rect 48134 16632 48190 16688
rect 48226 15408 48282 15464
rect 48134 15272 48190 15328
rect 48778 15000 48834 15056
rect 48134 13912 48190 13968
rect 48778 13776 48834 13832
rect 48134 12688 48190 12744
rect 48778 13640 48834 13696
rect 48226 12552 48282 12608
rect 48778 12552 48834 12608
rect 48778 12280 48834 12336
rect 48134 11328 48190 11384
rect 48226 11192 48282 11248
rect 48778 11192 48834 11248
rect 48134 8608 48190 8664
rect 48778 9560 48834 9616
rect 48226 8472 48282 8528
rect 48778 8472 48834 8528
rect 48134 7112 48190 7168
rect 48134 5888 48190 5944
rect 48778 6840 48834 6896
rect 48226 5752 48282 5808
rect 48778 5752 48834 5808
rect 48226 4392 48282 4448
rect 48134 4120 48190 4176
rect 24852 2202 24908 2204
rect 24932 2202 24988 2204
rect 25012 2202 25068 2204
rect 25092 2202 25148 2204
rect 24852 2150 24898 2202
rect 24898 2150 24908 2202
rect 24932 2150 24962 2202
rect 24962 2150 24974 2202
rect 24974 2150 24988 2202
rect 25012 2150 25026 2202
rect 25026 2150 25038 2202
rect 25038 2150 25068 2202
rect 25092 2150 25102 2202
rect 25102 2150 25148 2202
rect 24852 2148 24908 2150
rect 24932 2148 24988 2150
rect 25012 2148 25068 2150
rect 25092 2148 25148 2150
rect 30826 2746 30882 2748
rect 30906 2746 30962 2748
rect 30986 2746 31042 2748
rect 31066 2746 31122 2748
rect 30826 2694 30872 2746
rect 30872 2694 30882 2746
rect 30906 2694 30936 2746
rect 30936 2694 30948 2746
rect 30948 2694 30962 2746
rect 30986 2694 31000 2746
rect 31000 2694 31012 2746
rect 31012 2694 31042 2746
rect 31066 2694 31076 2746
rect 31076 2694 31122 2746
rect 30826 2692 30882 2694
rect 30906 2692 30962 2694
rect 30986 2692 31042 2694
rect 31066 2692 31122 2694
rect 42774 2746 42830 2748
rect 42854 2746 42910 2748
rect 42934 2746 42990 2748
rect 43014 2746 43070 2748
rect 42774 2694 42820 2746
rect 42820 2694 42830 2746
rect 42854 2694 42884 2746
rect 42884 2694 42896 2746
rect 42896 2694 42910 2746
rect 42934 2694 42948 2746
rect 42948 2694 42960 2746
rect 42960 2694 42990 2746
rect 43014 2694 43024 2746
rect 43024 2694 43070 2746
rect 42774 2692 42830 2694
rect 42854 2692 42910 2694
rect 42934 2692 42990 2694
rect 43014 2692 43070 2694
rect 36800 2202 36856 2204
rect 36880 2202 36936 2204
rect 36960 2202 37016 2204
rect 37040 2202 37096 2204
rect 36800 2150 36846 2202
rect 36846 2150 36856 2202
rect 36880 2150 36910 2202
rect 36910 2150 36922 2202
rect 36922 2150 36936 2202
rect 36960 2150 36974 2202
rect 36974 2150 36986 2202
rect 36986 2150 37016 2202
rect 37040 2150 37050 2202
rect 37050 2150 37096 2202
rect 36800 2148 36856 2150
rect 36880 2148 36936 2150
rect 36960 2148 37016 2150
rect 37040 2148 37096 2150
rect 45558 1672 45614 1728
rect 46846 2760 46902 2816
rect 48134 3032 48190 3088
rect 47766 1400 47822 1456
rect 46754 312 46810 368
rect 46662 40 46718 96
<< metal3 >>
rect 0 29338 800 29368
rect 2865 29338 2931 29341
rect 0 29336 2931 29338
rect 0 29280 2870 29336
rect 2926 29280 2931 29336
rect 0 29278 2931 29280
rect 0 29248 800 29278
rect 2865 29275 2931 29278
rect 49200 29248 50000 29368
rect 0 28658 800 28688
rect 2773 28658 2839 28661
rect 49200 28658 50000 28688
rect 0 28656 2839 28658
rect 0 28600 2778 28656
rect 2834 28600 2839 28656
rect 0 28598 2839 28600
rect 0 28568 800 28598
rect 2773 28595 2839 28598
rect 48270 28598 50000 28658
rect 45737 28250 45803 28253
rect 48270 28250 48330 28598
rect 49200 28568 50000 28598
rect 45737 28248 48330 28250
rect 45737 28192 45742 28248
rect 45798 28192 48330 28248
rect 45737 28190 48330 28192
rect 45737 28187 45803 28190
rect 0 27978 800 28008
rect 1393 27978 1459 27981
rect 49200 27978 50000 28008
rect 0 27976 1459 27978
rect 0 27920 1398 27976
rect 1454 27920 1459 27976
rect 0 27918 1459 27920
rect 0 27888 800 27918
rect 1393 27915 1459 27918
rect 48270 27918 50000 27978
rect 6920 27776 7236 27777
rect 6920 27712 6926 27776
rect 6990 27712 7006 27776
rect 7070 27712 7086 27776
rect 7150 27712 7166 27776
rect 7230 27712 7236 27776
rect 6920 27711 7236 27712
rect 18868 27776 19184 27777
rect 18868 27712 18874 27776
rect 18938 27712 18954 27776
rect 19018 27712 19034 27776
rect 19098 27712 19114 27776
rect 19178 27712 19184 27776
rect 18868 27711 19184 27712
rect 30816 27776 31132 27777
rect 30816 27712 30822 27776
rect 30886 27712 30902 27776
rect 30966 27712 30982 27776
rect 31046 27712 31062 27776
rect 31126 27712 31132 27776
rect 30816 27711 31132 27712
rect 42764 27776 43080 27777
rect 42764 27712 42770 27776
rect 42834 27712 42850 27776
rect 42914 27712 42930 27776
rect 42994 27712 43010 27776
rect 43074 27712 43080 27776
rect 42764 27711 43080 27712
rect 47485 27706 47551 27709
rect 48270 27706 48330 27918
rect 49200 27888 50000 27918
rect 47485 27704 48330 27706
rect 47485 27648 47490 27704
rect 47546 27648 48330 27704
rect 47485 27646 48330 27648
rect 47485 27643 47551 27646
rect 0 27298 800 27328
rect 1485 27298 1551 27301
rect 49200 27298 50000 27328
rect 0 27296 1551 27298
rect 0 27240 1490 27296
rect 1546 27240 1551 27296
rect 0 27238 1551 27240
rect 0 27208 800 27238
rect 1485 27235 1551 27238
rect 48270 27238 50000 27298
rect 12894 27232 13210 27233
rect 12894 27168 12900 27232
rect 12964 27168 12980 27232
rect 13044 27168 13060 27232
rect 13124 27168 13140 27232
rect 13204 27168 13210 27232
rect 12894 27167 13210 27168
rect 24842 27232 25158 27233
rect 24842 27168 24848 27232
rect 24912 27168 24928 27232
rect 24992 27168 25008 27232
rect 25072 27168 25088 27232
rect 25152 27168 25158 27232
rect 24842 27167 25158 27168
rect 36790 27232 37106 27233
rect 36790 27168 36796 27232
rect 36860 27168 36876 27232
rect 36940 27168 36956 27232
rect 37020 27168 37036 27232
rect 37100 27168 37106 27232
rect 36790 27167 37106 27168
rect 46841 26890 46907 26893
rect 48270 26890 48330 27238
rect 49200 27208 50000 27238
rect 46841 26888 48330 26890
rect 46841 26832 46846 26888
rect 46902 26832 48330 26888
rect 46841 26830 48330 26832
rect 46841 26827 46907 26830
rect 6920 26688 7236 26689
rect 0 26528 800 26648
rect 6920 26624 6926 26688
rect 6990 26624 7006 26688
rect 7070 26624 7086 26688
rect 7150 26624 7166 26688
rect 7230 26624 7236 26688
rect 6920 26623 7236 26624
rect 18868 26688 19184 26689
rect 18868 26624 18874 26688
rect 18938 26624 18954 26688
rect 19018 26624 19034 26688
rect 19098 26624 19114 26688
rect 19178 26624 19184 26688
rect 18868 26623 19184 26624
rect 30816 26688 31132 26689
rect 30816 26624 30822 26688
rect 30886 26624 30902 26688
rect 30966 26624 30982 26688
rect 31046 26624 31062 26688
rect 31126 26624 31132 26688
rect 30816 26623 31132 26624
rect 42764 26688 43080 26689
rect 42764 26624 42770 26688
rect 42834 26624 42850 26688
rect 42914 26624 42930 26688
rect 42994 26624 43010 26688
rect 43074 26624 43080 26688
rect 42764 26623 43080 26624
rect 49200 26618 50000 26648
rect 48270 26558 50000 26618
rect 48129 26346 48195 26349
rect 48270 26346 48330 26558
rect 49200 26528 50000 26558
rect 48129 26344 48330 26346
rect 48129 26288 48134 26344
rect 48190 26288 48330 26344
rect 48129 26286 48330 26288
rect 48129 26283 48195 26286
rect 12894 26144 13210 26145
rect 12894 26080 12900 26144
rect 12964 26080 12980 26144
rect 13044 26080 13060 26144
rect 13124 26080 13140 26144
rect 13204 26080 13210 26144
rect 12894 26079 13210 26080
rect 24842 26144 25158 26145
rect 24842 26080 24848 26144
rect 24912 26080 24928 26144
rect 24992 26080 25008 26144
rect 25072 26080 25088 26144
rect 25152 26080 25158 26144
rect 24842 26079 25158 26080
rect 36790 26144 37106 26145
rect 36790 26080 36796 26144
rect 36860 26080 36876 26144
rect 36940 26080 36956 26144
rect 37020 26080 37036 26144
rect 37100 26080 37106 26144
rect 36790 26079 37106 26080
rect 0 25938 800 25968
rect 1393 25938 1459 25941
rect 49200 25938 50000 25968
rect 0 25936 1459 25938
rect 0 25880 1398 25936
rect 1454 25880 1459 25936
rect 0 25878 1459 25880
rect 0 25848 800 25878
rect 1393 25875 1459 25878
rect 48270 25878 50000 25938
rect 6920 25600 7236 25601
rect 6920 25536 6926 25600
rect 6990 25536 7006 25600
rect 7070 25536 7086 25600
rect 7150 25536 7166 25600
rect 7230 25536 7236 25600
rect 6920 25535 7236 25536
rect 18868 25600 19184 25601
rect 18868 25536 18874 25600
rect 18938 25536 18954 25600
rect 19018 25536 19034 25600
rect 19098 25536 19114 25600
rect 19178 25536 19184 25600
rect 18868 25535 19184 25536
rect 30816 25600 31132 25601
rect 30816 25536 30822 25600
rect 30886 25536 30902 25600
rect 30966 25536 30982 25600
rect 31046 25536 31062 25600
rect 31126 25536 31132 25600
rect 30816 25535 31132 25536
rect 42764 25600 43080 25601
rect 42764 25536 42770 25600
rect 42834 25536 42850 25600
rect 42914 25536 42930 25600
rect 42994 25536 43010 25600
rect 43074 25536 43080 25600
rect 42764 25535 43080 25536
rect 48270 25533 48330 25878
rect 49200 25848 50000 25878
rect 48221 25530 48330 25533
rect 48140 25528 48330 25530
rect 48140 25472 48226 25528
rect 48282 25472 48330 25528
rect 48140 25470 48330 25472
rect 48221 25467 48287 25470
rect 0 25258 800 25288
rect 1393 25258 1459 25261
rect 49200 25258 50000 25288
rect 0 25256 1459 25258
rect 0 25200 1398 25256
rect 1454 25200 1459 25256
rect 0 25198 1459 25200
rect 0 25168 800 25198
rect 1393 25195 1459 25198
rect 48270 25198 50000 25258
rect 12894 25056 13210 25057
rect 12894 24992 12900 25056
rect 12964 24992 12980 25056
rect 13044 24992 13060 25056
rect 13124 24992 13140 25056
rect 13204 24992 13210 25056
rect 12894 24991 13210 24992
rect 24842 25056 25158 25057
rect 24842 24992 24848 25056
rect 24912 24992 24928 25056
rect 24992 24992 25008 25056
rect 25072 24992 25088 25056
rect 25152 24992 25158 25056
rect 24842 24991 25158 24992
rect 36790 25056 37106 25057
rect 36790 24992 36796 25056
rect 36860 24992 36876 25056
rect 36940 24992 36956 25056
rect 37020 24992 37036 25056
rect 37100 24992 37106 25056
rect 36790 24991 37106 24992
rect 48129 24986 48195 24989
rect 48270 24986 48330 25198
rect 49200 25168 50000 25198
rect 48129 24984 48330 24986
rect 48129 24928 48134 24984
rect 48190 24928 48330 24984
rect 48129 24926 48330 24928
rect 48129 24923 48195 24926
rect 0 24578 800 24608
rect 1393 24578 1459 24581
rect 49200 24578 50000 24608
rect 0 24576 1459 24578
rect 0 24520 1398 24576
rect 1454 24520 1459 24576
rect 0 24518 1459 24520
rect 0 24488 800 24518
rect 1393 24515 1459 24518
rect 48270 24518 50000 24578
rect 6920 24512 7236 24513
rect 6920 24448 6926 24512
rect 6990 24448 7006 24512
rect 7070 24448 7086 24512
rect 7150 24448 7166 24512
rect 7230 24448 7236 24512
rect 6920 24447 7236 24448
rect 18868 24512 19184 24513
rect 18868 24448 18874 24512
rect 18938 24448 18954 24512
rect 19018 24448 19034 24512
rect 19098 24448 19114 24512
rect 19178 24448 19184 24512
rect 18868 24447 19184 24448
rect 30816 24512 31132 24513
rect 30816 24448 30822 24512
rect 30886 24448 30902 24512
rect 30966 24448 30982 24512
rect 31046 24448 31062 24512
rect 31126 24448 31132 24512
rect 30816 24447 31132 24448
rect 42764 24512 43080 24513
rect 42764 24448 42770 24512
rect 42834 24448 42850 24512
rect 42914 24448 42930 24512
rect 42994 24448 43010 24512
rect 43074 24448 43080 24512
rect 42764 24447 43080 24448
rect 12894 23968 13210 23969
rect 0 23898 800 23928
rect 12894 23904 12900 23968
rect 12964 23904 12980 23968
rect 13044 23904 13060 23968
rect 13124 23904 13140 23968
rect 13204 23904 13210 23968
rect 12894 23903 13210 23904
rect 24842 23968 25158 23969
rect 24842 23904 24848 23968
rect 24912 23904 24928 23968
rect 24992 23904 25008 23968
rect 25072 23904 25088 23968
rect 25152 23904 25158 23968
rect 24842 23903 25158 23904
rect 36790 23968 37106 23969
rect 36790 23904 36796 23968
rect 36860 23904 36876 23968
rect 36940 23904 36956 23968
rect 37020 23904 37036 23968
rect 37100 23904 37106 23968
rect 36790 23903 37106 23904
rect 1393 23898 1459 23901
rect 0 23896 1459 23898
rect 0 23840 1398 23896
rect 1454 23840 1459 23896
rect 0 23838 1459 23840
rect 0 23808 800 23838
rect 1393 23835 1459 23838
rect 48129 23626 48195 23629
rect 48270 23626 48330 24518
rect 49200 24488 50000 24518
rect 49200 23898 50000 23928
rect 48129 23624 48330 23626
rect 48129 23568 48134 23624
rect 48190 23568 48330 23624
rect 48129 23566 48330 23568
rect 48822 23838 50000 23898
rect 48129 23563 48195 23566
rect 48221 23490 48287 23493
rect 48822 23490 48882 23838
rect 49200 23808 50000 23838
rect 48140 23488 48882 23490
rect 48140 23432 48226 23488
rect 48282 23432 48882 23488
rect 48140 23430 48882 23432
rect 48221 23427 48287 23430
rect 6920 23424 7236 23425
rect 6920 23360 6926 23424
rect 6990 23360 7006 23424
rect 7070 23360 7086 23424
rect 7150 23360 7166 23424
rect 7230 23360 7236 23424
rect 6920 23359 7236 23360
rect 18868 23424 19184 23425
rect 18868 23360 18874 23424
rect 18938 23360 18954 23424
rect 19018 23360 19034 23424
rect 19098 23360 19114 23424
rect 19178 23360 19184 23424
rect 18868 23359 19184 23360
rect 30816 23424 31132 23425
rect 30816 23360 30822 23424
rect 30886 23360 30902 23424
rect 30966 23360 30982 23424
rect 31046 23360 31062 23424
rect 31126 23360 31132 23424
rect 30816 23359 31132 23360
rect 42764 23424 43080 23425
rect 42764 23360 42770 23424
rect 42834 23360 42850 23424
rect 42914 23360 42930 23424
rect 42994 23360 43010 23424
rect 43074 23360 43080 23424
rect 42764 23359 43080 23360
rect 0 23218 800 23248
rect 1393 23218 1459 23221
rect 49200 23218 50000 23248
rect 0 23216 1459 23218
rect 0 23160 1398 23216
rect 1454 23160 1459 23216
rect 0 23158 1459 23160
rect 0 23128 800 23158
rect 1393 23155 1459 23158
rect 48270 23158 50000 23218
rect 12894 22880 13210 22881
rect 12894 22816 12900 22880
rect 12964 22816 12980 22880
rect 13044 22816 13060 22880
rect 13124 22816 13140 22880
rect 13204 22816 13210 22880
rect 12894 22815 13210 22816
rect 24842 22880 25158 22881
rect 24842 22816 24848 22880
rect 24912 22816 24928 22880
rect 24992 22816 25008 22880
rect 25072 22816 25088 22880
rect 25152 22816 25158 22880
rect 24842 22815 25158 22816
rect 36790 22880 37106 22881
rect 36790 22816 36796 22880
rect 36860 22816 36876 22880
rect 36940 22816 36956 22880
rect 37020 22816 37036 22880
rect 37100 22816 37106 22880
rect 36790 22815 37106 22816
rect 0 22448 800 22568
rect 6920 22336 7236 22337
rect 6920 22272 6926 22336
rect 6990 22272 7006 22336
rect 7070 22272 7086 22336
rect 7150 22272 7166 22336
rect 7230 22272 7236 22336
rect 6920 22271 7236 22272
rect 18868 22336 19184 22337
rect 18868 22272 18874 22336
rect 18938 22272 18954 22336
rect 19018 22272 19034 22336
rect 19098 22272 19114 22336
rect 19178 22272 19184 22336
rect 18868 22271 19184 22272
rect 30816 22336 31132 22337
rect 30816 22272 30822 22336
rect 30886 22272 30902 22336
rect 30966 22272 30982 22336
rect 31046 22272 31062 22336
rect 31126 22272 31132 22336
rect 30816 22271 31132 22272
rect 42764 22336 43080 22337
rect 42764 22272 42770 22336
rect 42834 22272 42850 22336
rect 42914 22272 42930 22336
rect 42994 22272 43010 22336
rect 43074 22272 43080 22336
rect 42764 22271 43080 22272
rect 48270 22269 48330 23158
rect 49200 23128 50000 23158
rect 49200 22538 50000 22568
rect 48221 22266 48330 22269
rect 48140 22264 48330 22266
rect 48140 22208 48226 22264
rect 48282 22208 48330 22264
rect 48140 22206 48330 22208
rect 48822 22478 50000 22538
rect 48221 22203 48287 22206
rect 48129 22130 48195 22133
rect 48822 22130 48882 22478
rect 49200 22448 50000 22478
rect 48129 22128 48882 22130
rect 48129 22072 48134 22128
rect 48190 22072 48882 22128
rect 48129 22070 48882 22072
rect 48129 22067 48195 22070
rect 0 21858 800 21888
rect 1393 21858 1459 21861
rect 49200 21858 50000 21888
rect 0 21856 1459 21858
rect 0 21800 1398 21856
rect 1454 21800 1459 21856
rect 0 21798 1459 21800
rect 0 21768 800 21798
rect 1393 21795 1459 21798
rect 48270 21798 50000 21858
rect 12894 21792 13210 21793
rect 12894 21728 12900 21792
rect 12964 21728 12980 21792
rect 13044 21728 13060 21792
rect 13124 21728 13140 21792
rect 13204 21728 13210 21792
rect 12894 21727 13210 21728
rect 24842 21792 25158 21793
rect 24842 21728 24848 21792
rect 24912 21728 24928 21792
rect 24992 21728 25008 21792
rect 25072 21728 25088 21792
rect 25152 21728 25158 21792
rect 24842 21727 25158 21728
rect 36790 21792 37106 21793
rect 36790 21728 36796 21792
rect 36860 21728 36876 21792
rect 36940 21728 36956 21792
rect 37020 21728 37036 21792
rect 37100 21728 37106 21792
rect 36790 21727 37106 21728
rect 6920 21248 7236 21249
rect 0 21178 800 21208
rect 6920 21184 6926 21248
rect 6990 21184 7006 21248
rect 7070 21184 7086 21248
rect 7150 21184 7166 21248
rect 7230 21184 7236 21248
rect 6920 21183 7236 21184
rect 18868 21248 19184 21249
rect 18868 21184 18874 21248
rect 18938 21184 18954 21248
rect 19018 21184 19034 21248
rect 19098 21184 19114 21248
rect 19178 21184 19184 21248
rect 18868 21183 19184 21184
rect 30816 21248 31132 21249
rect 30816 21184 30822 21248
rect 30886 21184 30902 21248
rect 30966 21184 30982 21248
rect 31046 21184 31062 21248
rect 31126 21184 31132 21248
rect 30816 21183 31132 21184
rect 42764 21248 43080 21249
rect 42764 21184 42770 21248
rect 42834 21184 42850 21248
rect 42914 21184 42930 21248
rect 42994 21184 43010 21248
rect 43074 21184 43080 21248
rect 42764 21183 43080 21184
rect 1393 21178 1459 21181
rect 0 21176 1459 21178
rect 0 21120 1398 21176
rect 1454 21120 1459 21176
rect 0 21118 1459 21120
rect 0 21088 800 21118
rect 1393 21115 1459 21118
rect 48129 20770 48195 20773
rect 48270 20770 48330 21798
rect 49200 21768 50000 21798
rect 49200 21088 50000 21208
rect 48129 20768 48330 20770
rect 48129 20712 48134 20768
rect 48190 20712 48330 20768
rect 48129 20710 48330 20712
rect 48129 20707 48195 20710
rect 12894 20704 13210 20705
rect 12894 20640 12900 20704
rect 12964 20640 12980 20704
rect 13044 20640 13060 20704
rect 13124 20640 13140 20704
rect 13204 20640 13210 20704
rect 12894 20639 13210 20640
rect 24842 20704 25158 20705
rect 24842 20640 24848 20704
rect 24912 20640 24928 20704
rect 24992 20640 25008 20704
rect 25072 20640 25088 20704
rect 25152 20640 25158 20704
rect 24842 20639 25158 20640
rect 36790 20704 37106 20705
rect 36790 20640 36796 20704
rect 36860 20640 36876 20704
rect 36940 20640 36956 20704
rect 37020 20640 37036 20704
rect 37100 20640 37106 20704
rect 36790 20639 37106 20640
rect 0 20498 800 20528
rect 1393 20498 1459 20501
rect 49200 20498 50000 20528
rect 0 20496 1459 20498
rect 0 20440 1398 20496
rect 1454 20440 1459 20496
rect 0 20438 1459 20440
rect 0 20408 800 20438
rect 1393 20435 1459 20438
rect 48270 20438 50000 20498
rect 6920 20160 7236 20161
rect 6920 20096 6926 20160
rect 6990 20096 7006 20160
rect 7070 20096 7086 20160
rect 7150 20096 7166 20160
rect 7230 20096 7236 20160
rect 6920 20095 7236 20096
rect 18868 20160 19184 20161
rect 18868 20096 18874 20160
rect 18938 20096 18954 20160
rect 19018 20096 19034 20160
rect 19098 20096 19114 20160
rect 19178 20096 19184 20160
rect 18868 20095 19184 20096
rect 30816 20160 31132 20161
rect 30816 20096 30822 20160
rect 30886 20096 30902 20160
rect 30966 20096 30982 20160
rect 31046 20096 31062 20160
rect 31126 20096 31132 20160
rect 30816 20095 31132 20096
rect 42764 20160 43080 20161
rect 42764 20096 42770 20160
rect 42834 20096 42850 20160
rect 42914 20096 42930 20160
rect 42994 20096 43010 20160
rect 43074 20096 43080 20160
rect 42764 20095 43080 20096
rect 0 19818 800 19848
rect 1393 19818 1459 19821
rect 0 19816 1459 19818
rect 0 19760 1398 19816
rect 1454 19760 1459 19816
rect 0 19758 1459 19760
rect 0 19728 800 19758
rect 1393 19755 1459 19758
rect 12894 19616 13210 19617
rect 12894 19552 12900 19616
rect 12964 19552 12980 19616
rect 13044 19552 13060 19616
rect 13124 19552 13140 19616
rect 13204 19552 13210 19616
rect 12894 19551 13210 19552
rect 24842 19616 25158 19617
rect 24842 19552 24848 19616
rect 24912 19552 24928 19616
rect 24992 19552 25008 19616
rect 25072 19552 25088 19616
rect 25152 19552 25158 19616
rect 24842 19551 25158 19552
rect 36790 19616 37106 19617
rect 36790 19552 36796 19616
rect 36860 19552 36876 19616
rect 36940 19552 36956 19616
rect 37020 19552 37036 19616
rect 37100 19552 37106 19616
rect 36790 19551 37106 19552
rect 48270 19413 48330 20438
rect 49200 20408 50000 20438
rect 49200 19728 50000 19848
rect 48221 19410 48330 19413
rect 48140 19408 48330 19410
rect 48140 19352 48226 19408
rect 48282 19352 48330 19408
rect 48140 19350 48330 19352
rect 48221 19347 48287 19350
rect 0 19138 800 19168
rect 1393 19138 1459 19141
rect 49200 19138 50000 19168
rect 0 19136 1459 19138
rect 0 19080 1398 19136
rect 1454 19080 1459 19136
rect 0 19078 1459 19080
rect 0 19048 800 19078
rect 1393 19075 1459 19078
rect 48270 19078 50000 19138
rect 6920 19072 7236 19073
rect 6920 19008 6926 19072
rect 6990 19008 7006 19072
rect 7070 19008 7086 19072
rect 7150 19008 7166 19072
rect 7230 19008 7236 19072
rect 6920 19007 7236 19008
rect 18868 19072 19184 19073
rect 18868 19008 18874 19072
rect 18938 19008 18954 19072
rect 19018 19008 19034 19072
rect 19098 19008 19114 19072
rect 19178 19008 19184 19072
rect 18868 19007 19184 19008
rect 30816 19072 31132 19073
rect 30816 19008 30822 19072
rect 30886 19008 30902 19072
rect 30966 19008 30982 19072
rect 31046 19008 31062 19072
rect 31126 19008 31132 19072
rect 30816 19007 31132 19008
rect 42764 19072 43080 19073
rect 42764 19008 42770 19072
rect 42834 19008 42850 19072
rect 42914 19008 42930 19072
rect 42994 19008 43010 19072
rect 43074 19008 43080 19072
rect 42764 19007 43080 19008
rect 12894 18528 13210 18529
rect 0 18458 800 18488
rect 12894 18464 12900 18528
rect 12964 18464 12980 18528
rect 13044 18464 13060 18528
rect 13124 18464 13140 18528
rect 13204 18464 13210 18528
rect 12894 18463 13210 18464
rect 24842 18528 25158 18529
rect 24842 18464 24848 18528
rect 24912 18464 24928 18528
rect 24992 18464 25008 18528
rect 25072 18464 25088 18528
rect 25152 18464 25158 18528
rect 24842 18463 25158 18464
rect 36790 18528 37106 18529
rect 36790 18464 36796 18528
rect 36860 18464 36876 18528
rect 36940 18464 36956 18528
rect 37020 18464 37036 18528
rect 37100 18464 37106 18528
rect 36790 18463 37106 18464
rect 1393 18458 1459 18461
rect 0 18456 1459 18458
rect 0 18400 1398 18456
rect 1454 18400 1459 18456
rect 0 18398 1459 18400
rect 0 18368 800 18398
rect 1393 18395 1459 18398
rect 48129 18186 48195 18189
rect 48270 18186 48330 19078
rect 49200 19048 50000 19078
rect 49200 18458 50000 18488
rect 48129 18184 48330 18186
rect 48129 18128 48134 18184
rect 48190 18128 48330 18184
rect 48129 18126 48330 18128
rect 48822 18398 50000 18458
rect 48129 18123 48195 18126
rect 48221 18050 48287 18053
rect 48822 18050 48882 18398
rect 49200 18368 50000 18398
rect 48140 18048 48882 18050
rect 48140 17992 48226 18048
rect 48282 17992 48882 18048
rect 48140 17990 48882 17992
rect 48221 17987 48287 17990
rect 6920 17984 7236 17985
rect 6920 17920 6926 17984
rect 6990 17920 7006 17984
rect 7070 17920 7086 17984
rect 7150 17920 7166 17984
rect 7230 17920 7236 17984
rect 6920 17919 7236 17920
rect 18868 17984 19184 17985
rect 18868 17920 18874 17984
rect 18938 17920 18954 17984
rect 19018 17920 19034 17984
rect 19098 17920 19114 17984
rect 19178 17920 19184 17984
rect 18868 17919 19184 17920
rect 30816 17984 31132 17985
rect 30816 17920 30822 17984
rect 30886 17920 30902 17984
rect 30966 17920 30982 17984
rect 31046 17920 31062 17984
rect 31126 17920 31132 17984
rect 30816 17919 31132 17920
rect 42764 17984 43080 17985
rect 42764 17920 42770 17984
rect 42834 17920 42850 17984
rect 42914 17920 42930 17984
rect 42994 17920 43010 17984
rect 43074 17920 43080 17984
rect 42764 17919 43080 17920
rect 0 17688 800 17808
rect 49200 17778 50000 17808
rect 48270 17718 50000 17778
rect 12894 17440 13210 17441
rect 12894 17376 12900 17440
rect 12964 17376 12980 17440
rect 13044 17376 13060 17440
rect 13124 17376 13140 17440
rect 13204 17376 13210 17440
rect 12894 17375 13210 17376
rect 24842 17440 25158 17441
rect 24842 17376 24848 17440
rect 24912 17376 24928 17440
rect 24992 17376 25008 17440
rect 25072 17376 25088 17440
rect 25152 17376 25158 17440
rect 24842 17375 25158 17376
rect 36790 17440 37106 17441
rect 36790 17376 36796 17440
rect 36860 17376 36876 17440
rect 36940 17376 36956 17440
rect 37020 17376 37036 17440
rect 37100 17376 37106 17440
rect 36790 17375 37106 17376
rect 0 17008 800 17128
rect 6920 16896 7236 16897
rect 6920 16832 6926 16896
rect 6990 16832 7006 16896
rect 7070 16832 7086 16896
rect 7150 16832 7166 16896
rect 7230 16832 7236 16896
rect 6920 16831 7236 16832
rect 18868 16896 19184 16897
rect 18868 16832 18874 16896
rect 18938 16832 18954 16896
rect 19018 16832 19034 16896
rect 19098 16832 19114 16896
rect 19178 16832 19184 16896
rect 18868 16831 19184 16832
rect 30816 16896 31132 16897
rect 30816 16832 30822 16896
rect 30886 16832 30902 16896
rect 30966 16832 30982 16896
rect 31046 16832 31062 16896
rect 31126 16832 31132 16896
rect 30816 16831 31132 16832
rect 42764 16896 43080 16897
rect 42764 16832 42770 16896
rect 42834 16832 42850 16896
rect 42914 16832 42930 16896
rect 42994 16832 43010 16896
rect 43074 16832 43080 16896
rect 42764 16831 43080 16832
rect 48270 16829 48330 17718
rect 49200 17688 50000 17718
rect 49200 17098 50000 17128
rect 48221 16826 48330 16829
rect 48140 16824 48330 16826
rect 48140 16768 48226 16824
rect 48282 16768 48330 16824
rect 48140 16766 48330 16768
rect 48822 17038 50000 17098
rect 48221 16763 48287 16766
rect 48129 16690 48195 16693
rect 48822 16690 48882 17038
rect 49200 17008 50000 17038
rect 48129 16688 48882 16690
rect 48129 16632 48134 16688
rect 48190 16632 48882 16688
rect 48129 16630 48882 16632
rect 48129 16627 48195 16630
rect 0 16328 800 16448
rect 49200 16418 50000 16448
rect 48270 16358 50000 16418
rect 12894 16352 13210 16353
rect 12894 16288 12900 16352
rect 12964 16288 12980 16352
rect 13044 16288 13060 16352
rect 13124 16288 13140 16352
rect 13204 16288 13210 16352
rect 12894 16287 13210 16288
rect 24842 16352 25158 16353
rect 24842 16288 24848 16352
rect 24912 16288 24928 16352
rect 24992 16288 25008 16352
rect 25072 16288 25088 16352
rect 25152 16288 25158 16352
rect 24842 16287 25158 16288
rect 36790 16352 37106 16353
rect 36790 16288 36796 16352
rect 36860 16288 36876 16352
rect 36940 16288 36956 16352
rect 37020 16288 37036 16352
rect 37100 16288 37106 16352
rect 36790 16287 37106 16288
rect 6920 15808 7236 15809
rect 0 15738 800 15768
rect 6920 15744 6926 15808
rect 6990 15744 7006 15808
rect 7070 15744 7086 15808
rect 7150 15744 7166 15808
rect 7230 15744 7236 15808
rect 6920 15743 7236 15744
rect 18868 15808 19184 15809
rect 18868 15744 18874 15808
rect 18938 15744 18954 15808
rect 19018 15744 19034 15808
rect 19098 15744 19114 15808
rect 19178 15744 19184 15808
rect 18868 15743 19184 15744
rect 30816 15808 31132 15809
rect 30816 15744 30822 15808
rect 30886 15744 30902 15808
rect 30966 15744 30982 15808
rect 31046 15744 31062 15808
rect 31126 15744 31132 15808
rect 30816 15743 31132 15744
rect 42764 15808 43080 15809
rect 42764 15744 42770 15808
rect 42834 15744 42850 15808
rect 42914 15744 42930 15808
rect 42994 15744 43010 15808
rect 43074 15744 43080 15808
rect 42764 15743 43080 15744
rect 1393 15738 1459 15741
rect 0 15736 1459 15738
rect 0 15680 1398 15736
rect 1454 15680 1459 15736
rect 0 15678 1459 15680
rect 0 15648 800 15678
rect 1393 15675 1459 15678
rect 48270 15469 48330 16358
rect 49200 16328 50000 16358
rect 49200 15738 50000 15768
rect 48221 15466 48330 15469
rect 48140 15464 48330 15466
rect 48140 15408 48226 15464
rect 48282 15408 48330 15464
rect 48140 15406 48330 15408
rect 48822 15678 50000 15738
rect 48221 15403 48287 15406
rect 48129 15330 48195 15333
rect 48822 15330 48882 15678
rect 49200 15648 50000 15678
rect 48129 15328 48882 15330
rect 48129 15272 48134 15328
rect 48190 15272 48882 15328
rect 48129 15270 48882 15272
rect 48129 15267 48195 15270
rect 12894 15264 13210 15265
rect 12894 15200 12900 15264
rect 12964 15200 12980 15264
rect 13044 15200 13060 15264
rect 13124 15200 13140 15264
rect 13204 15200 13210 15264
rect 12894 15199 13210 15200
rect 24842 15264 25158 15265
rect 24842 15200 24848 15264
rect 24912 15200 24928 15264
rect 24992 15200 25008 15264
rect 25072 15200 25088 15264
rect 25152 15200 25158 15264
rect 24842 15199 25158 15200
rect 36790 15264 37106 15265
rect 36790 15200 36796 15264
rect 36860 15200 36876 15264
rect 36940 15200 36956 15264
rect 37020 15200 37036 15264
rect 37100 15200 37106 15264
rect 36790 15199 37106 15200
rect 0 15058 800 15088
rect 1393 15058 1459 15061
rect 0 15056 1459 15058
rect 0 15000 1398 15056
rect 1454 15000 1459 15056
rect 0 14998 1459 15000
rect 0 14968 800 14998
rect 1393 14995 1459 14998
rect 48773 15058 48839 15061
rect 49200 15058 50000 15088
rect 48773 15056 50000 15058
rect 48773 15000 48778 15056
rect 48834 15000 50000 15056
rect 48773 14998 50000 15000
rect 48773 14995 48839 14998
rect 49200 14968 50000 14998
rect 6920 14720 7236 14721
rect 6920 14656 6926 14720
rect 6990 14656 7006 14720
rect 7070 14656 7086 14720
rect 7150 14656 7166 14720
rect 7230 14656 7236 14720
rect 6920 14655 7236 14656
rect 18868 14720 19184 14721
rect 18868 14656 18874 14720
rect 18938 14656 18954 14720
rect 19018 14656 19034 14720
rect 19098 14656 19114 14720
rect 19178 14656 19184 14720
rect 18868 14655 19184 14656
rect 30816 14720 31132 14721
rect 30816 14656 30822 14720
rect 30886 14656 30902 14720
rect 30966 14656 30982 14720
rect 31046 14656 31062 14720
rect 31126 14656 31132 14720
rect 30816 14655 31132 14656
rect 42764 14720 43080 14721
rect 42764 14656 42770 14720
rect 42834 14656 42850 14720
rect 42914 14656 42930 14720
rect 42994 14656 43010 14720
rect 43074 14656 43080 14720
rect 42764 14655 43080 14656
rect 0 14378 800 14408
rect 1393 14378 1459 14381
rect 49200 14378 50000 14408
rect 0 14376 1459 14378
rect 0 14320 1398 14376
rect 1454 14320 1459 14376
rect 0 14318 1459 14320
rect 0 14288 800 14318
rect 1393 14315 1459 14318
rect 48270 14318 50000 14378
rect 12894 14176 13210 14177
rect 12894 14112 12900 14176
rect 12964 14112 12980 14176
rect 13044 14112 13060 14176
rect 13124 14112 13140 14176
rect 13204 14112 13210 14176
rect 12894 14111 13210 14112
rect 24842 14176 25158 14177
rect 24842 14112 24848 14176
rect 24912 14112 24928 14176
rect 24992 14112 25008 14176
rect 25072 14112 25088 14176
rect 25152 14112 25158 14176
rect 24842 14111 25158 14112
rect 36790 14176 37106 14177
rect 36790 14112 36796 14176
rect 36860 14112 36876 14176
rect 36940 14112 36956 14176
rect 37020 14112 37036 14176
rect 37100 14112 37106 14176
rect 36790 14111 37106 14112
rect 48129 13970 48195 13973
rect 48270 13970 48330 14318
rect 49200 14288 50000 14318
rect 48129 13968 48330 13970
rect 48129 13912 48134 13968
rect 48190 13912 48330 13968
rect 48129 13910 48330 13912
rect 48129 13907 48195 13910
rect 45553 13834 45619 13837
rect 48773 13834 48839 13837
rect 45553 13832 48839 13834
rect 45553 13776 45558 13832
rect 45614 13776 48778 13832
rect 48834 13776 48839 13832
rect 45553 13774 48839 13776
rect 45553 13771 45619 13774
rect 48773 13771 48839 13774
rect 0 13698 800 13728
rect 1393 13698 1459 13701
rect 0 13696 1459 13698
rect 0 13640 1398 13696
rect 1454 13640 1459 13696
rect 0 13638 1459 13640
rect 0 13608 800 13638
rect 1393 13635 1459 13638
rect 48773 13698 48839 13701
rect 49200 13698 50000 13728
rect 48773 13696 50000 13698
rect 48773 13640 48778 13696
rect 48834 13640 50000 13696
rect 48773 13638 50000 13640
rect 48773 13635 48839 13638
rect 6920 13632 7236 13633
rect 6920 13568 6926 13632
rect 6990 13568 7006 13632
rect 7070 13568 7086 13632
rect 7150 13568 7166 13632
rect 7230 13568 7236 13632
rect 6920 13567 7236 13568
rect 18868 13632 19184 13633
rect 18868 13568 18874 13632
rect 18938 13568 18954 13632
rect 19018 13568 19034 13632
rect 19098 13568 19114 13632
rect 19178 13568 19184 13632
rect 18868 13567 19184 13568
rect 30816 13632 31132 13633
rect 30816 13568 30822 13632
rect 30886 13568 30902 13632
rect 30966 13568 30982 13632
rect 31046 13568 31062 13632
rect 31126 13568 31132 13632
rect 30816 13567 31132 13568
rect 42764 13632 43080 13633
rect 42764 13568 42770 13632
rect 42834 13568 42850 13632
rect 42914 13568 42930 13632
rect 42994 13568 43010 13632
rect 43074 13568 43080 13632
rect 49200 13608 50000 13638
rect 42764 13567 43080 13568
rect 12894 13088 13210 13089
rect 0 12928 800 13048
rect 12894 13024 12900 13088
rect 12964 13024 12980 13088
rect 13044 13024 13060 13088
rect 13124 13024 13140 13088
rect 13204 13024 13210 13088
rect 12894 13023 13210 13024
rect 24842 13088 25158 13089
rect 24842 13024 24848 13088
rect 24912 13024 24928 13088
rect 24992 13024 25008 13088
rect 25072 13024 25088 13088
rect 25152 13024 25158 13088
rect 24842 13023 25158 13024
rect 36790 13088 37106 13089
rect 36790 13024 36796 13088
rect 36860 13024 36876 13088
rect 36940 13024 36956 13088
rect 37020 13024 37036 13088
rect 37100 13024 37106 13088
rect 36790 13023 37106 13024
rect 49200 13018 50000 13048
rect 48270 12958 50000 13018
rect 48129 12746 48195 12749
rect 48270 12746 48330 12958
rect 49200 12928 50000 12958
rect 48129 12744 48330 12746
rect 48129 12688 48134 12744
rect 48190 12688 48330 12744
rect 48129 12686 48330 12688
rect 48129 12683 48195 12686
rect 48221 12610 48287 12613
rect 48773 12610 48839 12613
rect 48140 12608 48839 12610
rect 48140 12552 48226 12608
rect 48282 12552 48778 12608
rect 48834 12552 48839 12608
rect 48140 12550 48839 12552
rect 48221 12547 48287 12550
rect 48773 12547 48839 12550
rect 6920 12544 7236 12545
rect 6920 12480 6926 12544
rect 6990 12480 7006 12544
rect 7070 12480 7086 12544
rect 7150 12480 7166 12544
rect 7230 12480 7236 12544
rect 6920 12479 7236 12480
rect 18868 12544 19184 12545
rect 18868 12480 18874 12544
rect 18938 12480 18954 12544
rect 19018 12480 19034 12544
rect 19098 12480 19114 12544
rect 19178 12480 19184 12544
rect 18868 12479 19184 12480
rect 30816 12544 31132 12545
rect 30816 12480 30822 12544
rect 30886 12480 30902 12544
rect 30966 12480 30982 12544
rect 31046 12480 31062 12544
rect 31126 12480 31132 12544
rect 30816 12479 31132 12480
rect 42764 12544 43080 12545
rect 42764 12480 42770 12544
rect 42834 12480 42850 12544
rect 42914 12480 42930 12544
rect 42994 12480 43010 12544
rect 43074 12480 43080 12544
rect 42764 12479 43080 12480
rect 0 12338 800 12368
rect 1393 12338 1459 12341
rect 0 12336 1459 12338
rect 0 12280 1398 12336
rect 1454 12280 1459 12336
rect 0 12278 1459 12280
rect 0 12248 800 12278
rect 1393 12275 1459 12278
rect 48773 12338 48839 12341
rect 49200 12338 50000 12368
rect 48773 12336 50000 12338
rect 48773 12280 48778 12336
rect 48834 12280 50000 12336
rect 48773 12278 50000 12280
rect 48773 12275 48839 12278
rect 49200 12248 50000 12278
rect 12894 12000 13210 12001
rect 12894 11936 12900 12000
rect 12964 11936 12980 12000
rect 13044 11936 13060 12000
rect 13124 11936 13140 12000
rect 13204 11936 13210 12000
rect 12894 11935 13210 11936
rect 24842 12000 25158 12001
rect 24842 11936 24848 12000
rect 24912 11936 24928 12000
rect 24992 11936 25008 12000
rect 25072 11936 25088 12000
rect 25152 11936 25158 12000
rect 24842 11935 25158 11936
rect 36790 12000 37106 12001
rect 36790 11936 36796 12000
rect 36860 11936 36876 12000
rect 36940 11936 36956 12000
rect 37020 11936 37036 12000
rect 37100 11936 37106 12000
rect 36790 11935 37106 11936
rect 0 11658 800 11688
rect 1393 11658 1459 11661
rect 49200 11658 50000 11688
rect 0 11656 1459 11658
rect 0 11600 1398 11656
rect 1454 11600 1459 11656
rect 0 11598 1459 11600
rect 0 11568 800 11598
rect 1393 11595 1459 11598
rect 48270 11598 50000 11658
rect 6920 11456 7236 11457
rect 6920 11392 6926 11456
rect 6990 11392 7006 11456
rect 7070 11392 7086 11456
rect 7150 11392 7166 11456
rect 7230 11392 7236 11456
rect 6920 11391 7236 11392
rect 18868 11456 19184 11457
rect 18868 11392 18874 11456
rect 18938 11392 18954 11456
rect 19018 11392 19034 11456
rect 19098 11392 19114 11456
rect 19178 11392 19184 11456
rect 18868 11391 19184 11392
rect 30816 11456 31132 11457
rect 30816 11392 30822 11456
rect 30886 11392 30902 11456
rect 30966 11392 30982 11456
rect 31046 11392 31062 11456
rect 31126 11392 31132 11456
rect 30816 11391 31132 11392
rect 42764 11456 43080 11457
rect 42764 11392 42770 11456
rect 42834 11392 42850 11456
rect 42914 11392 42930 11456
rect 42994 11392 43010 11456
rect 43074 11392 43080 11456
rect 42764 11391 43080 11392
rect 48129 11386 48195 11389
rect 48270 11386 48330 11598
rect 49200 11568 50000 11598
rect 48129 11384 48330 11386
rect 48129 11328 48134 11384
rect 48190 11328 48330 11384
rect 48129 11326 48330 11328
rect 48129 11323 48195 11326
rect 48221 11250 48287 11253
rect 48773 11250 48839 11253
rect 48140 11248 48839 11250
rect 48140 11192 48226 11248
rect 48282 11192 48778 11248
rect 48834 11192 48839 11248
rect 48140 11190 48839 11192
rect 48221 11187 48287 11190
rect 48773 11187 48839 11190
rect 0 10978 800 11008
rect 1393 10978 1459 10981
rect 0 10976 1459 10978
rect 0 10920 1398 10976
rect 1454 10920 1459 10976
rect 0 10918 1459 10920
rect 0 10888 800 10918
rect 1393 10915 1459 10918
rect 12894 10912 13210 10913
rect 12894 10848 12900 10912
rect 12964 10848 12980 10912
rect 13044 10848 13060 10912
rect 13124 10848 13140 10912
rect 13204 10848 13210 10912
rect 12894 10847 13210 10848
rect 24842 10912 25158 10913
rect 24842 10848 24848 10912
rect 24912 10848 24928 10912
rect 24992 10848 25008 10912
rect 25072 10848 25088 10912
rect 25152 10848 25158 10912
rect 24842 10847 25158 10848
rect 36790 10912 37106 10913
rect 36790 10848 36796 10912
rect 36860 10848 36876 10912
rect 36940 10848 36956 10912
rect 37020 10848 37036 10912
rect 37100 10848 37106 10912
rect 49200 10888 50000 11008
rect 36790 10847 37106 10848
rect 6920 10368 7236 10369
rect 0 10208 800 10328
rect 6920 10304 6926 10368
rect 6990 10304 7006 10368
rect 7070 10304 7086 10368
rect 7150 10304 7166 10368
rect 7230 10304 7236 10368
rect 6920 10303 7236 10304
rect 18868 10368 19184 10369
rect 18868 10304 18874 10368
rect 18938 10304 18954 10368
rect 19018 10304 19034 10368
rect 19098 10304 19114 10368
rect 19178 10304 19184 10368
rect 18868 10303 19184 10304
rect 30816 10368 31132 10369
rect 30816 10304 30822 10368
rect 30886 10304 30902 10368
rect 30966 10304 30982 10368
rect 31046 10304 31062 10368
rect 31126 10304 31132 10368
rect 30816 10303 31132 10304
rect 42764 10368 43080 10369
rect 42764 10304 42770 10368
rect 42834 10304 42850 10368
rect 42914 10304 42930 10368
rect 42994 10304 43010 10368
rect 43074 10304 43080 10368
rect 42764 10303 43080 10304
rect 49200 10208 50000 10328
rect 12894 9824 13210 9825
rect 12894 9760 12900 9824
rect 12964 9760 12980 9824
rect 13044 9760 13060 9824
rect 13124 9760 13140 9824
rect 13204 9760 13210 9824
rect 12894 9759 13210 9760
rect 24842 9824 25158 9825
rect 24842 9760 24848 9824
rect 24912 9760 24928 9824
rect 24992 9760 25008 9824
rect 25072 9760 25088 9824
rect 25152 9760 25158 9824
rect 24842 9759 25158 9760
rect 36790 9824 37106 9825
rect 36790 9760 36796 9824
rect 36860 9760 36876 9824
rect 36940 9760 36956 9824
rect 37020 9760 37036 9824
rect 37100 9760 37106 9824
rect 36790 9759 37106 9760
rect 0 9528 800 9648
rect 48773 9618 48839 9621
rect 49200 9618 50000 9648
rect 48773 9616 50000 9618
rect 48773 9560 48778 9616
rect 48834 9560 50000 9616
rect 48773 9558 50000 9560
rect 48773 9555 48839 9558
rect 49200 9528 50000 9558
rect 6920 9280 7236 9281
rect 6920 9216 6926 9280
rect 6990 9216 7006 9280
rect 7070 9216 7086 9280
rect 7150 9216 7166 9280
rect 7230 9216 7236 9280
rect 6920 9215 7236 9216
rect 18868 9280 19184 9281
rect 18868 9216 18874 9280
rect 18938 9216 18954 9280
rect 19018 9216 19034 9280
rect 19098 9216 19114 9280
rect 19178 9216 19184 9280
rect 18868 9215 19184 9216
rect 30816 9280 31132 9281
rect 30816 9216 30822 9280
rect 30886 9216 30902 9280
rect 30966 9216 30982 9280
rect 31046 9216 31062 9280
rect 31126 9216 31132 9280
rect 30816 9215 31132 9216
rect 42764 9280 43080 9281
rect 42764 9216 42770 9280
rect 42834 9216 42850 9280
rect 42914 9216 42930 9280
rect 42994 9216 43010 9280
rect 43074 9216 43080 9280
rect 42764 9215 43080 9216
rect 0 8938 800 8968
rect 1393 8938 1459 8941
rect 49200 8938 50000 8968
rect 0 8936 1459 8938
rect 0 8880 1398 8936
rect 1454 8880 1459 8936
rect 0 8878 1459 8880
rect 0 8848 800 8878
rect 1393 8875 1459 8878
rect 48270 8878 50000 8938
rect 12894 8736 13210 8737
rect 12894 8672 12900 8736
rect 12964 8672 12980 8736
rect 13044 8672 13060 8736
rect 13124 8672 13140 8736
rect 13204 8672 13210 8736
rect 12894 8671 13210 8672
rect 24842 8736 25158 8737
rect 24842 8672 24848 8736
rect 24912 8672 24928 8736
rect 24992 8672 25008 8736
rect 25072 8672 25088 8736
rect 25152 8672 25158 8736
rect 24842 8671 25158 8672
rect 36790 8736 37106 8737
rect 36790 8672 36796 8736
rect 36860 8672 36876 8736
rect 36940 8672 36956 8736
rect 37020 8672 37036 8736
rect 37100 8672 37106 8736
rect 36790 8671 37106 8672
rect 48129 8666 48195 8669
rect 48270 8666 48330 8878
rect 49200 8848 50000 8878
rect 48129 8664 48330 8666
rect 48129 8608 48134 8664
rect 48190 8608 48330 8664
rect 48129 8606 48330 8608
rect 48129 8603 48195 8606
rect 48221 8530 48287 8533
rect 48773 8530 48839 8533
rect 48140 8528 48839 8530
rect 48140 8472 48226 8528
rect 48282 8472 48778 8528
rect 48834 8472 48839 8528
rect 48140 8470 48839 8472
rect 48221 8467 48287 8470
rect 48773 8467 48839 8470
rect 0 8258 800 8288
rect 1393 8258 1459 8261
rect 0 8256 1459 8258
rect 0 8200 1398 8256
rect 1454 8200 1459 8256
rect 0 8198 1459 8200
rect 0 8168 800 8198
rect 1393 8195 1459 8198
rect 6920 8192 7236 8193
rect 6920 8128 6926 8192
rect 6990 8128 7006 8192
rect 7070 8128 7086 8192
rect 7150 8128 7166 8192
rect 7230 8128 7236 8192
rect 6920 8127 7236 8128
rect 18868 8192 19184 8193
rect 18868 8128 18874 8192
rect 18938 8128 18954 8192
rect 19018 8128 19034 8192
rect 19098 8128 19114 8192
rect 19178 8128 19184 8192
rect 18868 8127 19184 8128
rect 30816 8192 31132 8193
rect 30816 8128 30822 8192
rect 30886 8128 30902 8192
rect 30966 8128 30982 8192
rect 31046 8128 31062 8192
rect 31126 8128 31132 8192
rect 30816 8127 31132 8128
rect 42764 8192 43080 8193
rect 42764 8128 42770 8192
rect 42834 8128 42850 8192
rect 42914 8128 42930 8192
rect 42994 8128 43010 8192
rect 43074 8128 43080 8192
rect 49200 8168 50000 8288
rect 42764 8127 43080 8128
rect 12894 7648 13210 7649
rect 0 7578 800 7608
rect 12894 7584 12900 7648
rect 12964 7584 12980 7648
rect 13044 7584 13060 7648
rect 13124 7584 13140 7648
rect 13204 7584 13210 7648
rect 12894 7583 13210 7584
rect 24842 7648 25158 7649
rect 24842 7584 24848 7648
rect 24912 7584 24928 7648
rect 24992 7584 25008 7648
rect 25072 7584 25088 7648
rect 25152 7584 25158 7648
rect 24842 7583 25158 7584
rect 36790 7648 37106 7649
rect 36790 7584 36796 7648
rect 36860 7584 36876 7648
rect 36940 7584 36956 7648
rect 37020 7584 37036 7648
rect 37100 7584 37106 7648
rect 36790 7583 37106 7584
rect 1393 7578 1459 7581
rect 49200 7578 50000 7608
rect 0 7576 1459 7578
rect 0 7520 1398 7576
rect 1454 7520 1459 7576
rect 0 7518 1459 7520
rect 0 7488 800 7518
rect 1393 7515 1459 7518
rect 48270 7518 50000 7578
rect 48129 7170 48195 7173
rect 48270 7170 48330 7518
rect 49200 7488 50000 7518
rect 48129 7168 48330 7170
rect 48129 7112 48134 7168
rect 48190 7112 48330 7168
rect 48129 7110 48330 7112
rect 48129 7107 48195 7110
rect 6920 7104 7236 7105
rect 6920 7040 6926 7104
rect 6990 7040 7006 7104
rect 7070 7040 7086 7104
rect 7150 7040 7166 7104
rect 7230 7040 7236 7104
rect 6920 7039 7236 7040
rect 18868 7104 19184 7105
rect 18868 7040 18874 7104
rect 18938 7040 18954 7104
rect 19018 7040 19034 7104
rect 19098 7040 19114 7104
rect 19178 7040 19184 7104
rect 18868 7039 19184 7040
rect 30816 7104 31132 7105
rect 30816 7040 30822 7104
rect 30886 7040 30902 7104
rect 30966 7040 30982 7104
rect 31046 7040 31062 7104
rect 31126 7040 31132 7104
rect 30816 7039 31132 7040
rect 42764 7104 43080 7105
rect 42764 7040 42770 7104
rect 42834 7040 42850 7104
rect 42914 7040 42930 7104
rect 42994 7040 43010 7104
rect 43074 7040 43080 7104
rect 42764 7039 43080 7040
rect 0 6898 800 6928
rect 1393 6898 1459 6901
rect 0 6896 1459 6898
rect 0 6840 1398 6896
rect 1454 6840 1459 6896
rect 0 6838 1459 6840
rect 0 6808 800 6838
rect 1393 6835 1459 6838
rect 48773 6898 48839 6901
rect 49200 6898 50000 6928
rect 48773 6896 50000 6898
rect 48773 6840 48778 6896
rect 48834 6840 50000 6896
rect 48773 6838 50000 6840
rect 48773 6835 48839 6838
rect 49200 6808 50000 6838
rect 12894 6560 13210 6561
rect 12894 6496 12900 6560
rect 12964 6496 12980 6560
rect 13044 6496 13060 6560
rect 13124 6496 13140 6560
rect 13204 6496 13210 6560
rect 12894 6495 13210 6496
rect 24842 6560 25158 6561
rect 24842 6496 24848 6560
rect 24912 6496 24928 6560
rect 24992 6496 25008 6560
rect 25072 6496 25088 6560
rect 25152 6496 25158 6560
rect 24842 6495 25158 6496
rect 36790 6560 37106 6561
rect 36790 6496 36796 6560
rect 36860 6496 36876 6560
rect 36940 6496 36956 6560
rect 37020 6496 37036 6560
rect 37100 6496 37106 6560
rect 36790 6495 37106 6496
rect 0 6218 800 6248
rect 1393 6218 1459 6221
rect 49200 6218 50000 6248
rect 0 6216 1459 6218
rect 0 6160 1398 6216
rect 1454 6160 1459 6216
rect 0 6158 1459 6160
rect 0 6128 800 6158
rect 1393 6155 1459 6158
rect 48270 6158 50000 6218
rect 6920 6016 7236 6017
rect 6920 5952 6926 6016
rect 6990 5952 7006 6016
rect 7070 5952 7086 6016
rect 7150 5952 7166 6016
rect 7230 5952 7236 6016
rect 6920 5951 7236 5952
rect 18868 6016 19184 6017
rect 18868 5952 18874 6016
rect 18938 5952 18954 6016
rect 19018 5952 19034 6016
rect 19098 5952 19114 6016
rect 19178 5952 19184 6016
rect 18868 5951 19184 5952
rect 30816 6016 31132 6017
rect 30816 5952 30822 6016
rect 30886 5952 30902 6016
rect 30966 5952 30982 6016
rect 31046 5952 31062 6016
rect 31126 5952 31132 6016
rect 30816 5951 31132 5952
rect 42764 6016 43080 6017
rect 42764 5952 42770 6016
rect 42834 5952 42850 6016
rect 42914 5952 42930 6016
rect 42994 5952 43010 6016
rect 43074 5952 43080 6016
rect 42764 5951 43080 5952
rect 48129 5946 48195 5949
rect 48270 5946 48330 6158
rect 49200 6128 50000 6158
rect 48129 5944 48330 5946
rect 48129 5888 48134 5944
rect 48190 5888 48330 5944
rect 48129 5886 48330 5888
rect 48129 5883 48195 5886
rect 48221 5810 48287 5813
rect 48773 5810 48839 5813
rect 48140 5808 48839 5810
rect 48140 5752 48226 5808
rect 48282 5752 48778 5808
rect 48834 5752 48839 5808
rect 48140 5750 48839 5752
rect 48221 5747 48287 5750
rect 48773 5747 48839 5750
rect 0 5538 800 5568
rect 1393 5538 1459 5541
rect 0 5536 1459 5538
rect 0 5480 1398 5536
rect 1454 5480 1459 5536
rect 0 5478 1459 5480
rect 0 5448 800 5478
rect 1393 5475 1459 5478
rect 12894 5472 13210 5473
rect 12894 5408 12900 5472
rect 12964 5408 12980 5472
rect 13044 5408 13060 5472
rect 13124 5408 13140 5472
rect 13204 5408 13210 5472
rect 12894 5407 13210 5408
rect 24842 5472 25158 5473
rect 24842 5408 24848 5472
rect 24912 5408 24928 5472
rect 24992 5408 25008 5472
rect 25072 5408 25088 5472
rect 25152 5408 25158 5472
rect 24842 5407 25158 5408
rect 36790 5472 37106 5473
rect 36790 5408 36796 5472
rect 36860 5408 36876 5472
rect 36940 5408 36956 5472
rect 37020 5408 37036 5472
rect 37100 5408 37106 5472
rect 49200 5448 50000 5568
rect 36790 5407 37106 5408
rect 6920 4928 7236 4929
rect 0 4858 800 4888
rect 6920 4864 6926 4928
rect 6990 4864 7006 4928
rect 7070 4864 7086 4928
rect 7150 4864 7166 4928
rect 7230 4864 7236 4928
rect 6920 4863 7236 4864
rect 18868 4928 19184 4929
rect 18868 4864 18874 4928
rect 18938 4864 18954 4928
rect 19018 4864 19034 4928
rect 19098 4864 19114 4928
rect 19178 4864 19184 4928
rect 18868 4863 19184 4864
rect 30816 4928 31132 4929
rect 30816 4864 30822 4928
rect 30886 4864 30902 4928
rect 30966 4864 30982 4928
rect 31046 4864 31062 4928
rect 31126 4864 31132 4928
rect 30816 4863 31132 4864
rect 42764 4928 43080 4929
rect 42764 4864 42770 4928
rect 42834 4864 42850 4928
rect 42914 4864 42930 4928
rect 42994 4864 43010 4928
rect 43074 4864 43080 4928
rect 42764 4863 43080 4864
rect 1393 4858 1459 4861
rect 49200 4858 50000 4888
rect 0 4856 1459 4858
rect 0 4800 1398 4856
rect 1454 4800 1459 4856
rect 0 4798 1459 4800
rect 0 4768 800 4798
rect 1393 4795 1459 4798
rect 48270 4798 50000 4858
rect 48270 4453 48330 4798
rect 49200 4768 50000 4798
rect 48221 4450 48330 4453
rect 48140 4448 48330 4450
rect 48140 4392 48226 4448
rect 48282 4392 48330 4448
rect 48140 4390 48330 4392
rect 48221 4387 48287 4390
rect 12894 4384 13210 4385
rect 12894 4320 12900 4384
rect 12964 4320 12980 4384
rect 13044 4320 13060 4384
rect 13124 4320 13140 4384
rect 13204 4320 13210 4384
rect 12894 4319 13210 4320
rect 24842 4384 25158 4385
rect 24842 4320 24848 4384
rect 24912 4320 24928 4384
rect 24992 4320 25008 4384
rect 25072 4320 25088 4384
rect 25152 4320 25158 4384
rect 24842 4319 25158 4320
rect 36790 4384 37106 4385
rect 36790 4320 36796 4384
rect 36860 4320 36876 4384
rect 36940 4320 36956 4384
rect 37020 4320 37036 4384
rect 37100 4320 37106 4384
rect 36790 4319 37106 4320
rect 0 4088 800 4208
rect 48129 4178 48195 4181
rect 49200 4178 50000 4208
rect 48129 4176 50000 4178
rect 48129 4120 48134 4176
rect 48190 4120 50000 4176
rect 48129 4118 50000 4120
rect 48129 4115 48195 4118
rect 49200 4088 50000 4118
rect 6920 3840 7236 3841
rect 6920 3776 6926 3840
rect 6990 3776 7006 3840
rect 7070 3776 7086 3840
rect 7150 3776 7166 3840
rect 7230 3776 7236 3840
rect 6920 3775 7236 3776
rect 18868 3840 19184 3841
rect 18868 3776 18874 3840
rect 18938 3776 18954 3840
rect 19018 3776 19034 3840
rect 19098 3776 19114 3840
rect 19178 3776 19184 3840
rect 18868 3775 19184 3776
rect 30816 3840 31132 3841
rect 30816 3776 30822 3840
rect 30886 3776 30902 3840
rect 30966 3776 30982 3840
rect 31046 3776 31062 3840
rect 31126 3776 31132 3840
rect 30816 3775 31132 3776
rect 42764 3840 43080 3841
rect 42764 3776 42770 3840
rect 42834 3776 42850 3840
rect 42914 3776 42930 3840
rect 42994 3776 43010 3840
rect 43074 3776 43080 3840
rect 42764 3775 43080 3776
rect 0 3498 800 3528
rect 1393 3498 1459 3501
rect 49200 3498 50000 3528
rect 0 3496 1459 3498
rect 0 3440 1398 3496
rect 1454 3440 1459 3496
rect 0 3438 1459 3440
rect 0 3408 800 3438
rect 1393 3435 1459 3438
rect 48270 3438 50000 3498
rect 12894 3296 13210 3297
rect 12894 3232 12900 3296
rect 12964 3232 12980 3296
rect 13044 3232 13060 3296
rect 13124 3232 13140 3296
rect 13204 3232 13210 3296
rect 12894 3231 13210 3232
rect 24842 3296 25158 3297
rect 24842 3232 24848 3296
rect 24912 3232 24928 3296
rect 24992 3232 25008 3296
rect 25072 3232 25088 3296
rect 25152 3232 25158 3296
rect 24842 3231 25158 3232
rect 36790 3296 37106 3297
rect 36790 3232 36796 3296
rect 36860 3232 36876 3296
rect 36940 3232 36956 3296
rect 37020 3232 37036 3296
rect 37100 3232 37106 3296
rect 36790 3231 37106 3232
rect 48129 3090 48195 3093
rect 48270 3090 48330 3438
rect 49200 3408 50000 3438
rect 48129 3088 48330 3090
rect 48129 3032 48134 3088
rect 48190 3032 48330 3088
rect 48129 3030 48330 3032
rect 48129 3027 48195 3030
rect 0 2728 800 2848
rect 46841 2818 46907 2821
rect 49200 2818 50000 2848
rect 46841 2816 50000 2818
rect 46841 2760 46846 2816
rect 46902 2760 50000 2816
rect 46841 2758 50000 2760
rect 46841 2755 46907 2758
rect 6920 2752 7236 2753
rect 6920 2688 6926 2752
rect 6990 2688 7006 2752
rect 7070 2688 7086 2752
rect 7150 2688 7166 2752
rect 7230 2688 7236 2752
rect 6920 2687 7236 2688
rect 18868 2752 19184 2753
rect 18868 2688 18874 2752
rect 18938 2688 18954 2752
rect 19018 2688 19034 2752
rect 19098 2688 19114 2752
rect 19178 2688 19184 2752
rect 18868 2687 19184 2688
rect 30816 2752 31132 2753
rect 30816 2688 30822 2752
rect 30886 2688 30902 2752
rect 30966 2688 30982 2752
rect 31046 2688 31062 2752
rect 31126 2688 31132 2752
rect 30816 2687 31132 2688
rect 42764 2752 43080 2753
rect 42764 2688 42770 2752
rect 42834 2688 42850 2752
rect 42914 2688 42930 2752
rect 42994 2688 43010 2752
rect 43074 2688 43080 2752
rect 49200 2728 50000 2758
rect 42764 2687 43080 2688
rect 12894 2208 13210 2209
rect 0 2138 800 2168
rect 12894 2144 12900 2208
rect 12964 2144 12980 2208
rect 13044 2144 13060 2208
rect 13124 2144 13140 2208
rect 13204 2144 13210 2208
rect 12894 2143 13210 2144
rect 24842 2208 25158 2209
rect 24842 2144 24848 2208
rect 24912 2144 24928 2208
rect 24992 2144 25008 2208
rect 25072 2144 25088 2208
rect 25152 2144 25158 2208
rect 24842 2143 25158 2144
rect 36790 2208 37106 2209
rect 36790 2144 36796 2208
rect 36860 2144 36876 2208
rect 36940 2144 36956 2208
rect 37020 2144 37036 2208
rect 37100 2144 37106 2208
rect 36790 2143 37106 2144
rect 2773 2138 2839 2141
rect 49200 2138 50000 2168
rect 0 2136 2839 2138
rect 0 2080 2778 2136
rect 2834 2080 2839 2136
rect 0 2078 2839 2080
rect 0 2048 800 2078
rect 2773 2075 2839 2078
rect 48270 2078 50000 2138
rect 45553 1730 45619 1733
rect 48270 1730 48330 2078
rect 49200 2048 50000 2078
rect 45553 1728 48330 1730
rect 45553 1672 45558 1728
rect 45614 1672 48330 1728
rect 45553 1670 48330 1672
rect 45553 1667 45619 1670
rect 0 1458 800 1488
rect 2865 1458 2931 1461
rect 0 1456 2931 1458
rect 0 1400 2870 1456
rect 2926 1400 2931 1456
rect 0 1398 2931 1400
rect 0 1368 800 1398
rect 2865 1395 2931 1398
rect 47761 1458 47827 1461
rect 49200 1458 50000 1488
rect 47761 1456 50000 1458
rect 47761 1400 47766 1456
rect 47822 1400 50000 1456
rect 47761 1398 50000 1400
rect 47761 1395 47827 1398
rect 49200 1368 50000 1398
rect 0 778 800 808
rect 2957 778 3023 781
rect 49200 778 50000 808
rect 0 776 3023 778
rect 0 720 2962 776
rect 3018 720 3023 776
rect 0 718 3023 720
rect 0 688 800 718
rect 2957 715 3023 718
rect 48270 718 50000 778
rect 46749 370 46815 373
rect 48270 370 48330 718
rect 49200 688 50000 718
rect 46749 368 48330 370
rect 46749 312 46754 368
rect 46810 312 48330 368
rect 46749 310 48330 312
rect 46749 307 46815 310
rect 0 98 800 128
rect 2957 98 3023 101
rect 0 96 3023 98
rect 0 40 2962 96
rect 3018 40 3023 96
rect 0 38 3023 40
rect 0 8 800 38
rect 2957 35 3023 38
rect 46657 98 46723 101
rect 49200 98 50000 128
rect 46657 96 50000 98
rect 46657 40 46662 96
rect 46718 40 50000 96
rect 46657 38 50000 40
rect 46657 35 46723 38
rect 49200 8 50000 38
<< via3 >>
rect 6926 27772 6990 27776
rect 6926 27716 6930 27772
rect 6930 27716 6986 27772
rect 6986 27716 6990 27772
rect 6926 27712 6990 27716
rect 7006 27772 7070 27776
rect 7006 27716 7010 27772
rect 7010 27716 7066 27772
rect 7066 27716 7070 27772
rect 7006 27712 7070 27716
rect 7086 27772 7150 27776
rect 7086 27716 7090 27772
rect 7090 27716 7146 27772
rect 7146 27716 7150 27772
rect 7086 27712 7150 27716
rect 7166 27772 7230 27776
rect 7166 27716 7170 27772
rect 7170 27716 7226 27772
rect 7226 27716 7230 27772
rect 7166 27712 7230 27716
rect 18874 27772 18938 27776
rect 18874 27716 18878 27772
rect 18878 27716 18934 27772
rect 18934 27716 18938 27772
rect 18874 27712 18938 27716
rect 18954 27772 19018 27776
rect 18954 27716 18958 27772
rect 18958 27716 19014 27772
rect 19014 27716 19018 27772
rect 18954 27712 19018 27716
rect 19034 27772 19098 27776
rect 19034 27716 19038 27772
rect 19038 27716 19094 27772
rect 19094 27716 19098 27772
rect 19034 27712 19098 27716
rect 19114 27772 19178 27776
rect 19114 27716 19118 27772
rect 19118 27716 19174 27772
rect 19174 27716 19178 27772
rect 19114 27712 19178 27716
rect 30822 27772 30886 27776
rect 30822 27716 30826 27772
rect 30826 27716 30882 27772
rect 30882 27716 30886 27772
rect 30822 27712 30886 27716
rect 30902 27772 30966 27776
rect 30902 27716 30906 27772
rect 30906 27716 30962 27772
rect 30962 27716 30966 27772
rect 30902 27712 30966 27716
rect 30982 27772 31046 27776
rect 30982 27716 30986 27772
rect 30986 27716 31042 27772
rect 31042 27716 31046 27772
rect 30982 27712 31046 27716
rect 31062 27772 31126 27776
rect 31062 27716 31066 27772
rect 31066 27716 31122 27772
rect 31122 27716 31126 27772
rect 31062 27712 31126 27716
rect 42770 27772 42834 27776
rect 42770 27716 42774 27772
rect 42774 27716 42830 27772
rect 42830 27716 42834 27772
rect 42770 27712 42834 27716
rect 42850 27772 42914 27776
rect 42850 27716 42854 27772
rect 42854 27716 42910 27772
rect 42910 27716 42914 27772
rect 42850 27712 42914 27716
rect 42930 27772 42994 27776
rect 42930 27716 42934 27772
rect 42934 27716 42990 27772
rect 42990 27716 42994 27772
rect 42930 27712 42994 27716
rect 43010 27772 43074 27776
rect 43010 27716 43014 27772
rect 43014 27716 43070 27772
rect 43070 27716 43074 27772
rect 43010 27712 43074 27716
rect 12900 27228 12964 27232
rect 12900 27172 12904 27228
rect 12904 27172 12960 27228
rect 12960 27172 12964 27228
rect 12900 27168 12964 27172
rect 12980 27228 13044 27232
rect 12980 27172 12984 27228
rect 12984 27172 13040 27228
rect 13040 27172 13044 27228
rect 12980 27168 13044 27172
rect 13060 27228 13124 27232
rect 13060 27172 13064 27228
rect 13064 27172 13120 27228
rect 13120 27172 13124 27228
rect 13060 27168 13124 27172
rect 13140 27228 13204 27232
rect 13140 27172 13144 27228
rect 13144 27172 13200 27228
rect 13200 27172 13204 27228
rect 13140 27168 13204 27172
rect 24848 27228 24912 27232
rect 24848 27172 24852 27228
rect 24852 27172 24908 27228
rect 24908 27172 24912 27228
rect 24848 27168 24912 27172
rect 24928 27228 24992 27232
rect 24928 27172 24932 27228
rect 24932 27172 24988 27228
rect 24988 27172 24992 27228
rect 24928 27168 24992 27172
rect 25008 27228 25072 27232
rect 25008 27172 25012 27228
rect 25012 27172 25068 27228
rect 25068 27172 25072 27228
rect 25008 27168 25072 27172
rect 25088 27228 25152 27232
rect 25088 27172 25092 27228
rect 25092 27172 25148 27228
rect 25148 27172 25152 27228
rect 25088 27168 25152 27172
rect 36796 27228 36860 27232
rect 36796 27172 36800 27228
rect 36800 27172 36856 27228
rect 36856 27172 36860 27228
rect 36796 27168 36860 27172
rect 36876 27228 36940 27232
rect 36876 27172 36880 27228
rect 36880 27172 36936 27228
rect 36936 27172 36940 27228
rect 36876 27168 36940 27172
rect 36956 27228 37020 27232
rect 36956 27172 36960 27228
rect 36960 27172 37016 27228
rect 37016 27172 37020 27228
rect 36956 27168 37020 27172
rect 37036 27228 37100 27232
rect 37036 27172 37040 27228
rect 37040 27172 37096 27228
rect 37096 27172 37100 27228
rect 37036 27168 37100 27172
rect 6926 26684 6990 26688
rect 6926 26628 6930 26684
rect 6930 26628 6986 26684
rect 6986 26628 6990 26684
rect 6926 26624 6990 26628
rect 7006 26684 7070 26688
rect 7006 26628 7010 26684
rect 7010 26628 7066 26684
rect 7066 26628 7070 26684
rect 7006 26624 7070 26628
rect 7086 26684 7150 26688
rect 7086 26628 7090 26684
rect 7090 26628 7146 26684
rect 7146 26628 7150 26684
rect 7086 26624 7150 26628
rect 7166 26684 7230 26688
rect 7166 26628 7170 26684
rect 7170 26628 7226 26684
rect 7226 26628 7230 26684
rect 7166 26624 7230 26628
rect 18874 26684 18938 26688
rect 18874 26628 18878 26684
rect 18878 26628 18934 26684
rect 18934 26628 18938 26684
rect 18874 26624 18938 26628
rect 18954 26684 19018 26688
rect 18954 26628 18958 26684
rect 18958 26628 19014 26684
rect 19014 26628 19018 26684
rect 18954 26624 19018 26628
rect 19034 26684 19098 26688
rect 19034 26628 19038 26684
rect 19038 26628 19094 26684
rect 19094 26628 19098 26684
rect 19034 26624 19098 26628
rect 19114 26684 19178 26688
rect 19114 26628 19118 26684
rect 19118 26628 19174 26684
rect 19174 26628 19178 26684
rect 19114 26624 19178 26628
rect 30822 26684 30886 26688
rect 30822 26628 30826 26684
rect 30826 26628 30882 26684
rect 30882 26628 30886 26684
rect 30822 26624 30886 26628
rect 30902 26684 30966 26688
rect 30902 26628 30906 26684
rect 30906 26628 30962 26684
rect 30962 26628 30966 26684
rect 30902 26624 30966 26628
rect 30982 26684 31046 26688
rect 30982 26628 30986 26684
rect 30986 26628 31042 26684
rect 31042 26628 31046 26684
rect 30982 26624 31046 26628
rect 31062 26684 31126 26688
rect 31062 26628 31066 26684
rect 31066 26628 31122 26684
rect 31122 26628 31126 26684
rect 31062 26624 31126 26628
rect 42770 26684 42834 26688
rect 42770 26628 42774 26684
rect 42774 26628 42830 26684
rect 42830 26628 42834 26684
rect 42770 26624 42834 26628
rect 42850 26684 42914 26688
rect 42850 26628 42854 26684
rect 42854 26628 42910 26684
rect 42910 26628 42914 26684
rect 42850 26624 42914 26628
rect 42930 26684 42994 26688
rect 42930 26628 42934 26684
rect 42934 26628 42990 26684
rect 42990 26628 42994 26684
rect 42930 26624 42994 26628
rect 43010 26684 43074 26688
rect 43010 26628 43014 26684
rect 43014 26628 43070 26684
rect 43070 26628 43074 26684
rect 43010 26624 43074 26628
rect 12900 26140 12964 26144
rect 12900 26084 12904 26140
rect 12904 26084 12960 26140
rect 12960 26084 12964 26140
rect 12900 26080 12964 26084
rect 12980 26140 13044 26144
rect 12980 26084 12984 26140
rect 12984 26084 13040 26140
rect 13040 26084 13044 26140
rect 12980 26080 13044 26084
rect 13060 26140 13124 26144
rect 13060 26084 13064 26140
rect 13064 26084 13120 26140
rect 13120 26084 13124 26140
rect 13060 26080 13124 26084
rect 13140 26140 13204 26144
rect 13140 26084 13144 26140
rect 13144 26084 13200 26140
rect 13200 26084 13204 26140
rect 13140 26080 13204 26084
rect 24848 26140 24912 26144
rect 24848 26084 24852 26140
rect 24852 26084 24908 26140
rect 24908 26084 24912 26140
rect 24848 26080 24912 26084
rect 24928 26140 24992 26144
rect 24928 26084 24932 26140
rect 24932 26084 24988 26140
rect 24988 26084 24992 26140
rect 24928 26080 24992 26084
rect 25008 26140 25072 26144
rect 25008 26084 25012 26140
rect 25012 26084 25068 26140
rect 25068 26084 25072 26140
rect 25008 26080 25072 26084
rect 25088 26140 25152 26144
rect 25088 26084 25092 26140
rect 25092 26084 25148 26140
rect 25148 26084 25152 26140
rect 25088 26080 25152 26084
rect 36796 26140 36860 26144
rect 36796 26084 36800 26140
rect 36800 26084 36856 26140
rect 36856 26084 36860 26140
rect 36796 26080 36860 26084
rect 36876 26140 36940 26144
rect 36876 26084 36880 26140
rect 36880 26084 36936 26140
rect 36936 26084 36940 26140
rect 36876 26080 36940 26084
rect 36956 26140 37020 26144
rect 36956 26084 36960 26140
rect 36960 26084 37016 26140
rect 37016 26084 37020 26140
rect 36956 26080 37020 26084
rect 37036 26140 37100 26144
rect 37036 26084 37040 26140
rect 37040 26084 37096 26140
rect 37096 26084 37100 26140
rect 37036 26080 37100 26084
rect 6926 25596 6990 25600
rect 6926 25540 6930 25596
rect 6930 25540 6986 25596
rect 6986 25540 6990 25596
rect 6926 25536 6990 25540
rect 7006 25596 7070 25600
rect 7006 25540 7010 25596
rect 7010 25540 7066 25596
rect 7066 25540 7070 25596
rect 7006 25536 7070 25540
rect 7086 25596 7150 25600
rect 7086 25540 7090 25596
rect 7090 25540 7146 25596
rect 7146 25540 7150 25596
rect 7086 25536 7150 25540
rect 7166 25596 7230 25600
rect 7166 25540 7170 25596
rect 7170 25540 7226 25596
rect 7226 25540 7230 25596
rect 7166 25536 7230 25540
rect 18874 25596 18938 25600
rect 18874 25540 18878 25596
rect 18878 25540 18934 25596
rect 18934 25540 18938 25596
rect 18874 25536 18938 25540
rect 18954 25596 19018 25600
rect 18954 25540 18958 25596
rect 18958 25540 19014 25596
rect 19014 25540 19018 25596
rect 18954 25536 19018 25540
rect 19034 25596 19098 25600
rect 19034 25540 19038 25596
rect 19038 25540 19094 25596
rect 19094 25540 19098 25596
rect 19034 25536 19098 25540
rect 19114 25596 19178 25600
rect 19114 25540 19118 25596
rect 19118 25540 19174 25596
rect 19174 25540 19178 25596
rect 19114 25536 19178 25540
rect 30822 25596 30886 25600
rect 30822 25540 30826 25596
rect 30826 25540 30882 25596
rect 30882 25540 30886 25596
rect 30822 25536 30886 25540
rect 30902 25596 30966 25600
rect 30902 25540 30906 25596
rect 30906 25540 30962 25596
rect 30962 25540 30966 25596
rect 30902 25536 30966 25540
rect 30982 25596 31046 25600
rect 30982 25540 30986 25596
rect 30986 25540 31042 25596
rect 31042 25540 31046 25596
rect 30982 25536 31046 25540
rect 31062 25596 31126 25600
rect 31062 25540 31066 25596
rect 31066 25540 31122 25596
rect 31122 25540 31126 25596
rect 31062 25536 31126 25540
rect 42770 25596 42834 25600
rect 42770 25540 42774 25596
rect 42774 25540 42830 25596
rect 42830 25540 42834 25596
rect 42770 25536 42834 25540
rect 42850 25596 42914 25600
rect 42850 25540 42854 25596
rect 42854 25540 42910 25596
rect 42910 25540 42914 25596
rect 42850 25536 42914 25540
rect 42930 25596 42994 25600
rect 42930 25540 42934 25596
rect 42934 25540 42990 25596
rect 42990 25540 42994 25596
rect 42930 25536 42994 25540
rect 43010 25596 43074 25600
rect 43010 25540 43014 25596
rect 43014 25540 43070 25596
rect 43070 25540 43074 25596
rect 43010 25536 43074 25540
rect 12900 25052 12964 25056
rect 12900 24996 12904 25052
rect 12904 24996 12960 25052
rect 12960 24996 12964 25052
rect 12900 24992 12964 24996
rect 12980 25052 13044 25056
rect 12980 24996 12984 25052
rect 12984 24996 13040 25052
rect 13040 24996 13044 25052
rect 12980 24992 13044 24996
rect 13060 25052 13124 25056
rect 13060 24996 13064 25052
rect 13064 24996 13120 25052
rect 13120 24996 13124 25052
rect 13060 24992 13124 24996
rect 13140 25052 13204 25056
rect 13140 24996 13144 25052
rect 13144 24996 13200 25052
rect 13200 24996 13204 25052
rect 13140 24992 13204 24996
rect 24848 25052 24912 25056
rect 24848 24996 24852 25052
rect 24852 24996 24908 25052
rect 24908 24996 24912 25052
rect 24848 24992 24912 24996
rect 24928 25052 24992 25056
rect 24928 24996 24932 25052
rect 24932 24996 24988 25052
rect 24988 24996 24992 25052
rect 24928 24992 24992 24996
rect 25008 25052 25072 25056
rect 25008 24996 25012 25052
rect 25012 24996 25068 25052
rect 25068 24996 25072 25052
rect 25008 24992 25072 24996
rect 25088 25052 25152 25056
rect 25088 24996 25092 25052
rect 25092 24996 25148 25052
rect 25148 24996 25152 25052
rect 25088 24992 25152 24996
rect 36796 25052 36860 25056
rect 36796 24996 36800 25052
rect 36800 24996 36856 25052
rect 36856 24996 36860 25052
rect 36796 24992 36860 24996
rect 36876 25052 36940 25056
rect 36876 24996 36880 25052
rect 36880 24996 36936 25052
rect 36936 24996 36940 25052
rect 36876 24992 36940 24996
rect 36956 25052 37020 25056
rect 36956 24996 36960 25052
rect 36960 24996 37016 25052
rect 37016 24996 37020 25052
rect 36956 24992 37020 24996
rect 37036 25052 37100 25056
rect 37036 24996 37040 25052
rect 37040 24996 37096 25052
rect 37096 24996 37100 25052
rect 37036 24992 37100 24996
rect 6926 24508 6990 24512
rect 6926 24452 6930 24508
rect 6930 24452 6986 24508
rect 6986 24452 6990 24508
rect 6926 24448 6990 24452
rect 7006 24508 7070 24512
rect 7006 24452 7010 24508
rect 7010 24452 7066 24508
rect 7066 24452 7070 24508
rect 7006 24448 7070 24452
rect 7086 24508 7150 24512
rect 7086 24452 7090 24508
rect 7090 24452 7146 24508
rect 7146 24452 7150 24508
rect 7086 24448 7150 24452
rect 7166 24508 7230 24512
rect 7166 24452 7170 24508
rect 7170 24452 7226 24508
rect 7226 24452 7230 24508
rect 7166 24448 7230 24452
rect 18874 24508 18938 24512
rect 18874 24452 18878 24508
rect 18878 24452 18934 24508
rect 18934 24452 18938 24508
rect 18874 24448 18938 24452
rect 18954 24508 19018 24512
rect 18954 24452 18958 24508
rect 18958 24452 19014 24508
rect 19014 24452 19018 24508
rect 18954 24448 19018 24452
rect 19034 24508 19098 24512
rect 19034 24452 19038 24508
rect 19038 24452 19094 24508
rect 19094 24452 19098 24508
rect 19034 24448 19098 24452
rect 19114 24508 19178 24512
rect 19114 24452 19118 24508
rect 19118 24452 19174 24508
rect 19174 24452 19178 24508
rect 19114 24448 19178 24452
rect 30822 24508 30886 24512
rect 30822 24452 30826 24508
rect 30826 24452 30882 24508
rect 30882 24452 30886 24508
rect 30822 24448 30886 24452
rect 30902 24508 30966 24512
rect 30902 24452 30906 24508
rect 30906 24452 30962 24508
rect 30962 24452 30966 24508
rect 30902 24448 30966 24452
rect 30982 24508 31046 24512
rect 30982 24452 30986 24508
rect 30986 24452 31042 24508
rect 31042 24452 31046 24508
rect 30982 24448 31046 24452
rect 31062 24508 31126 24512
rect 31062 24452 31066 24508
rect 31066 24452 31122 24508
rect 31122 24452 31126 24508
rect 31062 24448 31126 24452
rect 42770 24508 42834 24512
rect 42770 24452 42774 24508
rect 42774 24452 42830 24508
rect 42830 24452 42834 24508
rect 42770 24448 42834 24452
rect 42850 24508 42914 24512
rect 42850 24452 42854 24508
rect 42854 24452 42910 24508
rect 42910 24452 42914 24508
rect 42850 24448 42914 24452
rect 42930 24508 42994 24512
rect 42930 24452 42934 24508
rect 42934 24452 42990 24508
rect 42990 24452 42994 24508
rect 42930 24448 42994 24452
rect 43010 24508 43074 24512
rect 43010 24452 43014 24508
rect 43014 24452 43070 24508
rect 43070 24452 43074 24508
rect 43010 24448 43074 24452
rect 12900 23964 12964 23968
rect 12900 23908 12904 23964
rect 12904 23908 12960 23964
rect 12960 23908 12964 23964
rect 12900 23904 12964 23908
rect 12980 23964 13044 23968
rect 12980 23908 12984 23964
rect 12984 23908 13040 23964
rect 13040 23908 13044 23964
rect 12980 23904 13044 23908
rect 13060 23964 13124 23968
rect 13060 23908 13064 23964
rect 13064 23908 13120 23964
rect 13120 23908 13124 23964
rect 13060 23904 13124 23908
rect 13140 23964 13204 23968
rect 13140 23908 13144 23964
rect 13144 23908 13200 23964
rect 13200 23908 13204 23964
rect 13140 23904 13204 23908
rect 24848 23964 24912 23968
rect 24848 23908 24852 23964
rect 24852 23908 24908 23964
rect 24908 23908 24912 23964
rect 24848 23904 24912 23908
rect 24928 23964 24992 23968
rect 24928 23908 24932 23964
rect 24932 23908 24988 23964
rect 24988 23908 24992 23964
rect 24928 23904 24992 23908
rect 25008 23964 25072 23968
rect 25008 23908 25012 23964
rect 25012 23908 25068 23964
rect 25068 23908 25072 23964
rect 25008 23904 25072 23908
rect 25088 23964 25152 23968
rect 25088 23908 25092 23964
rect 25092 23908 25148 23964
rect 25148 23908 25152 23964
rect 25088 23904 25152 23908
rect 36796 23964 36860 23968
rect 36796 23908 36800 23964
rect 36800 23908 36856 23964
rect 36856 23908 36860 23964
rect 36796 23904 36860 23908
rect 36876 23964 36940 23968
rect 36876 23908 36880 23964
rect 36880 23908 36936 23964
rect 36936 23908 36940 23964
rect 36876 23904 36940 23908
rect 36956 23964 37020 23968
rect 36956 23908 36960 23964
rect 36960 23908 37016 23964
rect 37016 23908 37020 23964
rect 36956 23904 37020 23908
rect 37036 23964 37100 23968
rect 37036 23908 37040 23964
rect 37040 23908 37096 23964
rect 37096 23908 37100 23964
rect 37036 23904 37100 23908
rect 6926 23420 6990 23424
rect 6926 23364 6930 23420
rect 6930 23364 6986 23420
rect 6986 23364 6990 23420
rect 6926 23360 6990 23364
rect 7006 23420 7070 23424
rect 7006 23364 7010 23420
rect 7010 23364 7066 23420
rect 7066 23364 7070 23420
rect 7006 23360 7070 23364
rect 7086 23420 7150 23424
rect 7086 23364 7090 23420
rect 7090 23364 7146 23420
rect 7146 23364 7150 23420
rect 7086 23360 7150 23364
rect 7166 23420 7230 23424
rect 7166 23364 7170 23420
rect 7170 23364 7226 23420
rect 7226 23364 7230 23420
rect 7166 23360 7230 23364
rect 18874 23420 18938 23424
rect 18874 23364 18878 23420
rect 18878 23364 18934 23420
rect 18934 23364 18938 23420
rect 18874 23360 18938 23364
rect 18954 23420 19018 23424
rect 18954 23364 18958 23420
rect 18958 23364 19014 23420
rect 19014 23364 19018 23420
rect 18954 23360 19018 23364
rect 19034 23420 19098 23424
rect 19034 23364 19038 23420
rect 19038 23364 19094 23420
rect 19094 23364 19098 23420
rect 19034 23360 19098 23364
rect 19114 23420 19178 23424
rect 19114 23364 19118 23420
rect 19118 23364 19174 23420
rect 19174 23364 19178 23420
rect 19114 23360 19178 23364
rect 30822 23420 30886 23424
rect 30822 23364 30826 23420
rect 30826 23364 30882 23420
rect 30882 23364 30886 23420
rect 30822 23360 30886 23364
rect 30902 23420 30966 23424
rect 30902 23364 30906 23420
rect 30906 23364 30962 23420
rect 30962 23364 30966 23420
rect 30902 23360 30966 23364
rect 30982 23420 31046 23424
rect 30982 23364 30986 23420
rect 30986 23364 31042 23420
rect 31042 23364 31046 23420
rect 30982 23360 31046 23364
rect 31062 23420 31126 23424
rect 31062 23364 31066 23420
rect 31066 23364 31122 23420
rect 31122 23364 31126 23420
rect 31062 23360 31126 23364
rect 42770 23420 42834 23424
rect 42770 23364 42774 23420
rect 42774 23364 42830 23420
rect 42830 23364 42834 23420
rect 42770 23360 42834 23364
rect 42850 23420 42914 23424
rect 42850 23364 42854 23420
rect 42854 23364 42910 23420
rect 42910 23364 42914 23420
rect 42850 23360 42914 23364
rect 42930 23420 42994 23424
rect 42930 23364 42934 23420
rect 42934 23364 42990 23420
rect 42990 23364 42994 23420
rect 42930 23360 42994 23364
rect 43010 23420 43074 23424
rect 43010 23364 43014 23420
rect 43014 23364 43070 23420
rect 43070 23364 43074 23420
rect 43010 23360 43074 23364
rect 12900 22876 12964 22880
rect 12900 22820 12904 22876
rect 12904 22820 12960 22876
rect 12960 22820 12964 22876
rect 12900 22816 12964 22820
rect 12980 22876 13044 22880
rect 12980 22820 12984 22876
rect 12984 22820 13040 22876
rect 13040 22820 13044 22876
rect 12980 22816 13044 22820
rect 13060 22876 13124 22880
rect 13060 22820 13064 22876
rect 13064 22820 13120 22876
rect 13120 22820 13124 22876
rect 13060 22816 13124 22820
rect 13140 22876 13204 22880
rect 13140 22820 13144 22876
rect 13144 22820 13200 22876
rect 13200 22820 13204 22876
rect 13140 22816 13204 22820
rect 24848 22876 24912 22880
rect 24848 22820 24852 22876
rect 24852 22820 24908 22876
rect 24908 22820 24912 22876
rect 24848 22816 24912 22820
rect 24928 22876 24992 22880
rect 24928 22820 24932 22876
rect 24932 22820 24988 22876
rect 24988 22820 24992 22876
rect 24928 22816 24992 22820
rect 25008 22876 25072 22880
rect 25008 22820 25012 22876
rect 25012 22820 25068 22876
rect 25068 22820 25072 22876
rect 25008 22816 25072 22820
rect 25088 22876 25152 22880
rect 25088 22820 25092 22876
rect 25092 22820 25148 22876
rect 25148 22820 25152 22876
rect 25088 22816 25152 22820
rect 36796 22876 36860 22880
rect 36796 22820 36800 22876
rect 36800 22820 36856 22876
rect 36856 22820 36860 22876
rect 36796 22816 36860 22820
rect 36876 22876 36940 22880
rect 36876 22820 36880 22876
rect 36880 22820 36936 22876
rect 36936 22820 36940 22876
rect 36876 22816 36940 22820
rect 36956 22876 37020 22880
rect 36956 22820 36960 22876
rect 36960 22820 37016 22876
rect 37016 22820 37020 22876
rect 36956 22816 37020 22820
rect 37036 22876 37100 22880
rect 37036 22820 37040 22876
rect 37040 22820 37096 22876
rect 37096 22820 37100 22876
rect 37036 22816 37100 22820
rect 6926 22332 6990 22336
rect 6926 22276 6930 22332
rect 6930 22276 6986 22332
rect 6986 22276 6990 22332
rect 6926 22272 6990 22276
rect 7006 22332 7070 22336
rect 7006 22276 7010 22332
rect 7010 22276 7066 22332
rect 7066 22276 7070 22332
rect 7006 22272 7070 22276
rect 7086 22332 7150 22336
rect 7086 22276 7090 22332
rect 7090 22276 7146 22332
rect 7146 22276 7150 22332
rect 7086 22272 7150 22276
rect 7166 22332 7230 22336
rect 7166 22276 7170 22332
rect 7170 22276 7226 22332
rect 7226 22276 7230 22332
rect 7166 22272 7230 22276
rect 18874 22332 18938 22336
rect 18874 22276 18878 22332
rect 18878 22276 18934 22332
rect 18934 22276 18938 22332
rect 18874 22272 18938 22276
rect 18954 22332 19018 22336
rect 18954 22276 18958 22332
rect 18958 22276 19014 22332
rect 19014 22276 19018 22332
rect 18954 22272 19018 22276
rect 19034 22332 19098 22336
rect 19034 22276 19038 22332
rect 19038 22276 19094 22332
rect 19094 22276 19098 22332
rect 19034 22272 19098 22276
rect 19114 22332 19178 22336
rect 19114 22276 19118 22332
rect 19118 22276 19174 22332
rect 19174 22276 19178 22332
rect 19114 22272 19178 22276
rect 30822 22332 30886 22336
rect 30822 22276 30826 22332
rect 30826 22276 30882 22332
rect 30882 22276 30886 22332
rect 30822 22272 30886 22276
rect 30902 22332 30966 22336
rect 30902 22276 30906 22332
rect 30906 22276 30962 22332
rect 30962 22276 30966 22332
rect 30902 22272 30966 22276
rect 30982 22332 31046 22336
rect 30982 22276 30986 22332
rect 30986 22276 31042 22332
rect 31042 22276 31046 22332
rect 30982 22272 31046 22276
rect 31062 22332 31126 22336
rect 31062 22276 31066 22332
rect 31066 22276 31122 22332
rect 31122 22276 31126 22332
rect 31062 22272 31126 22276
rect 42770 22332 42834 22336
rect 42770 22276 42774 22332
rect 42774 22276 42830 22332
rect 42830 22276 42834 22332
rect 42770 22272 42834 22276
rect 42850 22332 42914 22336
rect 42850 22276 42854 22332
rect 42854 22276 42910 22332
rect 42910 22276 42914 22332
rect 42850 22272 42914 22276
rect 42930 22332 42994 22336
rect 42930 22276 42934 22332
rect 42934 22276 42990 22332
rect 42990 22276 42994 22332
rect 42930 22272 42994 22276
rect 43010 22332 43074 22336
rect 43010 22276 43014 22332
rect 43014 22276 43070 22332
rect 43070 22276 43074 22332
rect 43010 22272 43074 22276
rect 12900 21788 12964 21792
rect 12900 21732 12904 21788
rect 12904 21732 12960 21788
rect 12960 21732 12964 21788
rect 12900 21728 12964 21732
rect 12980 21788 13044 21792
rect 12980 21732 12984 21788
rect 12984 21732 13040 21788
rect 13040 21732 13044 21788
rect 12980 21728 13044 21732
rect 13060 21788 13124 21792
rect 13060 21732 13064 21788
rect 13064 21732 13120 21788
rect 13120 21732 13124 21788
rect 13060 21728 13124 21732
rect 13140 21788 13204 21792
rect 13140 21732 13144 21788
rect 13144 21732 13200 21788
rect 13200 21732 13204 21788
rect 13140 21728 13204 21732
rect 24848 21788 24912 21792
rect 24848 21732 24852 21788
rect 24852 21732 24908 21788
rect 24908 21732 24912 21788
rect 24848 21728 24912 21732
rect 24928 21788 24992 21792
rect 24928 21732 24932 21788
rect 24932 21732 24988 21788
rect 24988 21732 24992 21788
rect 24928 21728 24992 21732
rect 25008 21788 25072 21792
rect 25008 21732 25012 21788
rect 25012 21732 25068 21788
rect 25068 21732 25072 21788
rect 25008 21728 25072 21732
rect 25088 21788 25152 21792
rect 25088 21732 25092 21788
rect 25092 21732 25148 21788
rect 25148 21732 25152 21788
rect 25088 21728 25152 21732
rect 36796 21788 36860 21792
rect 36796 21732 36800 21788
rect 36800 21732 36856 21788
rect 36856 21732 36860 21788
rect 36796 21728 36860 21732
rect 36876 21788 36940 21792
rect 36876 21732 36880 21788
rect 36880 21732 36936 21788
rect 36936 21732 36940 21788
rect 36876 21728 36940 21732
rect 36956 21788 37020 21792
rect 36956 21732 36960 21788
rect 36960 21732 37016 21788
rect 37016 21732 37020 21788
rect 36956 21728 37020 21732
rect 37036 21788 37100 21792
rect 37036 21732 37040 21788
rect 37040 21732 37096 21788
rect 37096 21732 37100 21788
rect 37036 21728 37100 21732
rect 6926 21244 6990 21248
rect 6926 21188 6930 21244
rect 6930 21188 6986 21244
rect 6986 21188 6990 21244
rect 6926 21184 6990 21188
rect 7006 21244 7070 21248
rect 7006 21188 7010 21244
rect 7010 21188 7066 21244
rect 7066 21188 7070 21244
rect 7006 21184 7070 21188
rect 7086 21244 7150 21248
rect 7086 21188 7090 21244
rect 7090 21188 7146 21244
rect 7146 21188 7150 21244
rect 7086 21184 7150 21188
rect 7166 21244 7230 21248
rect 7166 21188 7170 21244
rect 7170 21188 7226 21244
rect 7226 21188 7230 21244
rect 7166 21184 7230 21188
rect 18874 21244 18938 21248
rect 18874 21188 18878 21244
rect 18878 21188 18934 21244
rect 18934 21188 18938 21244
rect 18874 21184 18938 21188
rect 18954 21244 19018 21248
rect 18954 21188 18958 21244
rect 18958 21188 19014 21244
rect 19014 21188 19018 21244
rect 18954 21184 19018 21188
rect 19034 21244 19098 21248
rect 19034 21188 19038 21244
rect 19038 21188 19094 21244
rect 19094 21188 19098 21244
rect 19034 21184 19098 21188
rect 19114 21244 19178 21248
rect 19114 21188 19118 21244
rect 19118 21188 19174 21244
rect 19174 21188 19178 21244
rect 19114 21184 19178 21188
rect 30822 21244 30886 21248
rect 30822 21188 30826 21244
rect 30826 21188 30882 21244
rect 30882 21188 30886 21244
rect 30822 21184 30886 21188
rect 30902 21244 30966 21248
rect 30902 21188 30906 21244
rect 30906 21188 30962 21244
rect 30962 21188 30966 21244
rect 30902 21184 30966 21188
rect 30982 21244 31046 21248
rect 30982 21188 30986 21244
rect 30986 21188 31042 21244
rect 31042 21188 31046 21244
rect 30982 21184 31046 21188
rect 31062 21244 31126 21248
rect 31062 21188 31066 21244
rect 31066 21188 31122 21244
rect 31122 21188 31126 21244
rect 31062 21184 31126 21188
rect 42770 21244 42834 21248
rect 42770 21188 42774 21244
rect 42774 21188 42830 21244
rect 42830 21188 42834 21244
rect 42770 21184 42834 21188
rect 42850 21244 42914 21248
rect 42850 21188 42854 21244
rect 42854 21188 42910 21244
rect 42910 21188 42914 21244
rect 42850 21184 42914 21188
rect 42930 21244 42994 21248
rect 42930 21188 42934 21244
rect 42934 21188 42990 21244
rect 42990 21188 42994 21244
rect 42930 21184 42994 21188
rect 43010 21244 43074 21248
rect 43010 21188 43014 21244
rect 43014 21188 43070 21244
rect 43070 21188 43074 21244
rect 43010 21184 43074 21188
rect 12900 20700 12964 20704
rect 12900 20644 12904 20700
rect 12904 20644 12960 20700
rect 12960 20644 12964 20700
rect 12900 20640 12964 20644
rect 12980 20700 13044 20704
rect 12980 20644 12984 20700
rect 12984 20644 13040 20700
rect 13040 20644 13044 20700
rect 12980 20640 13044 20644
rect 13060 20700 13124 20704
rect 13060 20644 13064 20700
rect 13064 20644 13120 20700
rect 13120 20644 13124 20700
rect 13060 20640 13124 20644
rect 13140 20700 13204 20704
rect 13140 20644 13144 20700
rect 13144 20644 13200 20700
rect 13200 20644 13204 20700
rect 13140 20640 13204 20644
rect 24848 20700 24912 20704
rect 24848 20644 24852 20700
rect 24852 20644 24908 20700
rect 24908 20644 24912 20700
rect 24848 20640 24912 20644
rect 24928 20700 24992 20704
rect 24928 20644 24932 20700
rect 24932 20644 24988 20700
rect 24988 20644 24992 20700
rect 24928 20640 24992 20644
rect 25008 20700 25072 20704
rect 25008 20644 25012 20700
rect 25012 20644 25068 20700
rect 25068 20644 25072 20700
rect 25008 20640 25072 20644
rect 25088 20700 25152 20704
rect 25088 20644 25092 20700
rect 25092 20644 25148 20700
rect 25148 20644 25152 20700
rect 25088 20640 25152 20644
rect 36796 20700 36860 20704
rect 36796 20644 36800 20700
rect 36800 20644 36856 20700
rect 36856 20644 36860 20700
rect 36796 20640 36860 20644
rect 36876 20700 36940 20704
rect 36876 20644 36880 20700
rect 36880 20644 36936 20700
rect 36936 20644 36940 20700
rect 36876 20640 36940 20644
rect 36956 20700 37020 20704
rect 36956 20644 36960 20700
rect 36960 20644 37016 20700
rect 37016 20644 37020 20700
rect 36956 20640 37020 20644
rect 37036 20700 37100 20704
rect 37036 20644 37040 20700
rect 37040 20644 37096 20700
rect 37096 20644 37100 20700
rect 37036 20640 37100 20644
rect 6926 20156 6990 20160
rect 6926 20100 6930 20156
rect 6930 20100 6986 20156
rect 6986 20100 6990 20156
rect 6926 20096 6990 20100
rect 7006 20156 7070 20160
rect 7006 20100 7010 20156
rect 7010 20100 7066 20156
rect 7066 20100 7070 20156
rect 7006 20096 7070 20100
rect 7086 20156 7150 20160
rect 7086 20100 7090 20156
rect 7090 20100 7146 20156
rect 7146 20100 7150 20156
rect 7086 20096 7150 20100
rect 7166 20156 7230 20160
rect 7166 20100 7170 20156
rect 7170 20100 7226 20156
rect 7226 20100 7230 20156
rect 7166 20096 7230 20100
rect 18874 20156 18938 20160
rect 18874 20100 18878 20156
rect 18878 20100 18934 20156
rect 18934 20100 18938 20156
rect 18874 20096 18938 20100
rect 18954 20156 19018 20160
rect 18954 20100 18958 20156
rect 18958 20100 19014 20156
rect 19014 20100 19018 20156
rect 18954 20096 19018 20100
rect 19034 20156 19098 20160
rect 19034 20100 19038 20156
rect 19038 20100 19094 20156
rect 19094 20100 19098 20156
rect 19034 20096 19098 20100
rect 19114 20156 19178 20160
rect 19114 20100 19118 20156
rect 19118 20100 19174 20156
rect 19174 20100 19178 20156
rect 19114 20096 19178 20100
rect 30822 20156 30886 20160
rect 30822 20100 30826 20156
rect 30826 20100 30882 20156
rect 30882 20100 30886 20156
rect 30822 20096 30886 20100
rect 30902 20156 30966 20160
rect 30902 20100 30906 20156
rect 30906 20100 30962 20156
rect 30962 20100 30966 20156
rect 30902 20096 30966 20100
rect 30982 20156 31046 20160
rect 30982 20100 30986 20156
rect 30986 20100 31042 20156
rect 31042 20100 31046 20156
rect 30982 20096 31046 20100
rect 31062 20156 31126 20160
rect 31062 20100 31066 20156
rect 31066 20100 31122 20156
rect 31122 20100 31126 20156
rect 31062 20096 31126 20100
rect 42770 20156 42834 20160
rect 42770 20100 42774 20156
rect 42774 20100 42830 20156
rect 42830 20100 42834 20156
rect 42770 20096 42834 20100
rect 42850 20156 42914 20160
rect 42850 20100 42854 20156
rect 42854 20100 42910 20156
rect 42910 20100 42914 20156
rect 42850 20096 42914 20100
rect 42930 20156 42994 20160
rect 42930 20100 42934 20156
rect 42934 20100 42990 20156
rect 42990 20100 42994 20156
rect 42930 20096 42994 20100
rect 43010 20156 43074 20160
rect 43010 20100 43014 20156
rect 43014 20100 43070 20156
rect 43070 20100 43074 20156
rect 43010 20096 43074 20100
rect 12900 19612 12964 19616
rect 12900 19556 12904 19612
rect 12904 19556 12960 19612
rect 12960 19556 12964 19612
rect 12900 19552 12964 19556
rect 12980 19612 13044 19616
rect 12980 19556 12984 19612
rect 12984 19556 13040 19612
rect 13040 19556 13044 19612
rect 12980 19552 13044 19556
rect 13060 19612 13124 19616
rect 13060 19556 13064 19612
rect 13064 19556 13120 19612
rect 13120 19556 13124 19612
rect 13060 19552 13124 19556
rect 13140 19612 13204 19616
rect 13140 19556 13144 19612
rect 13144 19556 13200 19612
rect 13200 19556 13204 19612
rect 13140 19552 13204 19556
rect 24848 19612 24912 19616
rect 24848 19556 24852 19612
rect 24852 19556 24908 19612
rect 24908 19556 24912 19612
rect 24848 19552 24912 19556
rect 24928 19612 24992 19616
rect 24928 19556 24932 19612
rect 24932 19556 24988 19612
rect 24988 19556 24992 19612
rect 24928 19552 24992 19556
rect 25008 19612 25072 19616
rect 25008 19556 25012 19612
rect 25012 19556 25068 19612
rect 25068 19556 25072 19612
rect 25008 19552 25072 19556
rect 25088 19612 25152 19616
rect 25088 19556 25092 19612
rect 25092 19556 25148 19612
rect 25148 19556 25152 19612
rect 25088 19552 25152 19556
rect 36796 19612 36860 19616
rect 36796 19556 36800 19612
rect 36800 19556 36856 19612
rect 36856 19556 36860 19612
rect 36796 19552 36860 19556
rect 36876 19612 36940 19616
rect 36876 19556 36880 19612
rect 36880 19556 36936 19612
rect 36936 19556 36940 19612
rect 36876 19552 36940 19556
rect 36956 19612 37020 19616
rect 36956 19556 36960 19612
rect 36960 19556 37016 19612
rect 37016 19556 37020 19612
rect 36956 19552 37020 19556
rect 37036 19612 37100 19616
rect 37036 19556 37040 19612
rect 37040 19556 37096 19612
rect 37096 19556 37100 19612
rect 37036 19552 37100 19556
rect 6926 19068 6990 19072
rect 6926 19012 6930 19068
rect 6930 19012 6986 19068
rect 6986 19012 6990 19068
rect 6926 19008 6990 19012
rect 7006 19068 7070 19072
rect 7006 19012 7010 19068
rect 7010 19012 7066 19068
rect 7066 19012 7070 19068
rect 7006 19008 7070 19012
rect 7086 19068 7150 19072
rect 7086 19012 7090 19068
rect 7090 19012 7146 19068
rect 7146 19012 7150 19068
rect 7086 19008 7150 19012
rect 7166 19068 7230 19072
rect 7166 19012 7170 19068
rect 7170 19012 7226 19068
rect 7226 19012 7230 19068
rect 7166 19008 7230 19012
rect 18874 19068 18938 19072
rect 18874 19012 18878 19068
rect 18878 19012 18934 19068
rect 18934 19012 18938 19068
rect 18874 19008 18938 19012
rect 18954 19068 19018 19072
rect 18954 19012 18958 19068
rect 18958 19012 19014 19068
rect 19014 19012 19018 19068
rect 18954 19008 19018 19012
rect 19034 19068 19098 19072
rect 19034 19012 19038 19068
rect 19038 19012 19094 19068
rect 19094 19012 19098 19068
rect 19034 19008 19098 19012
rect 19114 19068 19178 19072
rect 19114 19012 19118 19068
rect 19118 19012 19174 19068
rect 19174 19012 19178 19068
rect 19114 19008 19178 19012
rect 30822 19068 30886 19072
rect 30822 19012 30826 19068
rect 30826 19012 30882 19068
rect 30882 19012 30886 19068
rect 30822 19008 30886 19012
rect 30902 19068 30966 19072
rect 30902 19012 30906 19068
rect 30906 19012 30962 19068
rect 30962 19012 30966 19068
rect 30902 19008 30966 19012
rect 30982 19068 31046 19072
rect 30982 19012 30986 19068
rect 30986 19012 31042 19068
rect 31042 19012 31046 19068
rect 30982 19008 31046 19012
rect 31062 19068 31126 19072
rect 31062 19012 31066 19068
rect 31066 19012 31122 19068
rect 31122 19012 31126 19068
rect 31062 19008 31126 19012
rect 42770 19068 42834 19072
rect 42770 19012 42774 19068
rect 42774 19012 42830 19068
rect 42830 19012 42834 19068
rect 42770 19008 42834 19012
rect 42850 19068 42914 19072
rect 42850 19012 42854 19068
rect 42854 19012 42910 19068
rect 42910 19012 42914 19068
rect 42850 19008 42914 19012
rect 42930 19068 42994 19072
rect 42930 19012 42934 19068
rect 42934 19012 42990 19068
rect 42990 19012 42994 19068
rect 42930 19008 42994 19012
rect 43010 19068 43074 19072
rect 43010 19012 43014 19068
rect 43014 19012 43070 19068
rect 43070 19012 43074 19068
rect 43010 19008 43074 19012
rect 12900 18524 12964 18528
rect 12900 18468 12904 18524
rect 12904 18468 12960 18524
rect 12960 18468 12964 18524
rect 12900 18464 12964 18468
rect 12980 18524 13044 18528
rect 12980 18468 12984 18524
rect 12984 18468 13040 18524
rect 13040 18468 13044 18524
rect 12980 18464 13044 18468
rect 13060 18524 13124 18528
rect 13060 18468 13064 18524
rect 13064 18468 13120 18524
rect 13120 18468 13124 18524
rect 13060 18464 13124 18468
rect 13140 18524 13204 18528
rect 13140 18468 13144 18524
rect 13144 18468 13200 18524
rect 13200 18468 13204 18524
rect 13140 18464 13204 18468
rect 24848 18524 24912 18528
rect 24848 18468 24852 18524
rect 24852 18468 24908 18524
rect 24908 18468 24912 18524
rect 24848 18464 24912 18468
rect 24928 18524 24992 18528
rect 24928 18468 24932 18524
rect 24932 18468 24988 18524
rect 24988 18468 24992 18524
rect 24928 18464 24992 18468
rect 25008 18524 25072 18528
rect 25008 18468 25012 18524
rect 25012 18468 25068 18524
rect 25068 18468 25072 18524
rect 25008 18464 25072 18468
rect 25088 18524 25152 18528
rect 25088 18468 25092 18524
rect 25092 18468 25148 18524
rect 25148 18468 25152 18524
rect 25088 18464 25152 18468
rect 36796 18524 36860 18528
rect 36796 18468 36800 18524
rect 36800 18468 36856 18524
rect 36856 18468 36860 18524
rect 36796 18464 36860 18468
rect 36876 18524 36940 18528
rect 36876 18468 36880 18524
rect 36880 18468 36936 18524
rect 36936 18468 36940 18524
rect 36876 18464 36940 18468
rect 36956 18524 37020 18528
rect 36956 18468 36960 18524
rect 36960 18468 37016 18524
rect 37016 18468 37020 18524
rect 36956 18464 37020 18468
rect 37036 18524 37100 18528
rect 37036 18468 37040 18524
rect 37040 18468 37096 18524
rect 37096 18468 37100 18524
rect 37036 18464 37100 18468
rect 6926 17980 6990 17984
rect 6926 17924 6930 17980
rect 6930 17924 6986 17980
rect 6986 17924 6990 17980
rect 6926 17920 6990 17924
rect 7006 17980 7070 17984
rect 7006 17924 7010 17980
rect 7010 17924 7066 17980
rect 7066 17924 7070 17980
rect 7006 17920 7070 17924
rect 7086 17980 7150 17984
rect 7086 17924 7090 17980
rect 7090 17924 7146 17980
rect 7146 17924 7150 17980
rect 7086 17920 7150 17924
rect 7166 17980 7230 17984
rect 7166 17924 7170 17980
rect 7170 17924 7226 17980
rect 7226 17924 7230 17980
rect 7166 17920 7230 17924
rect 18874 17980 18938 17984
rect 18874 17924 18878 17980
rect 18878 17924 18934 17980
rect 18934 17924 18938 17980
rect 18874 17920 18938 17924
rect 18954 17980 19018 17984
rect 18954 17924 18958 17980
rect 18958 17924 19014 17980
rect 19014 17924 19018 17980
rect 18954 17920 19018 17924
rect 19034 17980 19098 17984
rect 19034 17924 19038 17980
rect 19038 17924 19094 17980
rect 19094 17924 19098 17980
rect 19034 17920 19098 17924
rect 19114 17980 19178 17984
rect 19114 17924 19118 17980
rect 19118 17924 19174 17980
rect 19174 17924 19178 17980
rect 19114 17920 19178 17924
rect 30822 17980 30886 17984
rect 30822 17924 30826 17980
rect 30826 17924 30882 17980
rect 30882 17924 30886 17980
rect 30822 17920 30886 17924
rect 30902 17980 30966 17984
rect 30902 17924 30906 17980
rect 30906 17924 30962 17980
rect 30962 17924 30966 17980
rect 30902 17920 30966 17924
rect 30982 17980 31046 17984
rect 30982 17924 30986 17980
rect 30986 17924 31042 17980
rect 31042 17924 31046 17980
rect 30982 17920 31046 17924
rect 31062 17980 31126 17984
rect 31062 17924 31066 17980
rect 31066 17924 31122 17980
rect 31122 17924 31126 17980
rect 31062 17920 31126 17924
rect 42770 17980 42834 17984
rect 42770 17924 42774 17980
rect 42774 17924 42830 17980
rect 42830 17924 42834 17980
rect 42770 17920 42834 17924
rect 42850 17980 42914 17984
rect 42850 17924 42854 17980
rect 42854 17924 42910 17980
rect 42910 17924 42914 17980
rect 42850 17920 42914 17924
rect 42930 17980 42994 17984
rect 42930 17924 42934 17980
rect 42934 17924 42990 17980
rect 42990 17924 42994 17980
rect 42930 17920 42994 17924
rect 43010 17980 43074 17984
rect 43010 17924 43014 17980
rect 43014 17924 43070 17980
rect 43070 17924 43074 17980
rect 43010 17920 43074 17924
rect 12900 17436 12964 17440
rect 12900 17380 12904 17436
rect 12904 17380 12960 17436
rect 12960 17380 12964 17436
rect 12900 17376 12964 17380
rect 12980 17436 13044 17440
rect 12980 17380 12984 17436
rect 12984 17380 13040 17436
rect 13040 17380 13044 17436
rect 12980 17376 13044 17380
rect 13060 17436 13124 17440
rect 13060 17380 13064 17436
rect 13064 17380 13120 17436
rect 13120 17380 13124 17436
rect 13060 17376 13124 17380
rect 13140 17436 13204 17440
rect 13140 17380 13144 17436
rect 13144 17380 13200 17436
rect 13200 17380 13204 17436
rect 13140 17376 13204 17380
rect 24848 17436 24912 17440
rect 24848 17380 24852 17436
rect 24852 17380 24908 17436
rect 24908 17380 24912 17436
rect 24848 17376 24912 17380
rect 24928 17436 24992 17440
rect 24928 17380 24932 17436
rect 24932 17380 24988 17436
rect 24988 17380 24992 17436
rect 24928 17376 24992 17380
rect 25008 17436 25072 17440
rect 25008 17380 25012 17436
rect 25012 17380 25068 17436
rect 25068 17380 25072 17436
rect 25008 17376 25072 17380
rect 25088 17436 25152 17440
rect 25088 17380 25092 17436
rect 25092 17380 25148 17436
rect 25148 17380 25152 17436
rect 25088 17376 25152 17380
rect 36796 17436 36860 17440
rect 36796 17380 36800 17436
rect 36800 17380 36856 17436
rect 36856 17380 36860 17436
rect 36796 17376 36860 17380
rect 36876 17436 36940 17440
rect 36876 17380 36880 17436
rect 36880 17380 36936 17436
rect 36936 17380 36940 17436
rect 36876 17376 36940 17380
rect 36956 17436 37020 17440
rect 36956 17380 36960 17436
rect 36960 17380 37016 17436
rect 37016 17380 37020 17436
rect 36956 17376 37020 17380
rect 37036 17436 37100 17440
rect 37036 17380 37040 17436
rect 37040 17380 37096 17436
rect 37096 17380 37100 17436
rect 37036 17376 37100 17380
rect 6926 16892 6990 16896
rect 6926 16836 6930 16892
rect 6930 16836 6986 16892
rect 6986 16836 6990 16892
rect 6926 16832 6990 16836
rect 7006 16892 7070 16896
rect 7006 16836 7010 16892
rect 7010 16836 7066 16892
rect 7066 16836 7070 16892
rect 7006 16832 7070 16836
rect 7086 16892 7150 16896
rect 7086 16836 7090 16892
rect 7090 16836 7146 16892
rect 7146 16836 7150 16892
rect 7086 16832 7150 16836
rect 7166 16892 7230 16896
rect 7166 16836 7170 16892
rect 7170 16836 7226 16892
rect 7226 16836 7230 16892
rect 7166 16832 7230 16836
rect 18874 16892 18938 16896
rect 18874 16836 18878 16892
rect 18878 16836 18934 16892
rect 18934 16836 18938 16892
rect 18874 16832 18938 16836
rect 18954 16892 19018 16896
rect 18954 16836 18958 16892
rect 18958 16836 19014 16892
rect 19014 16836 19018 16892
rect 18954 16832 19018 16836
rect 19034 16892 19098 16896
rect 19034 16836 19038 16892
rect 19038 16836 19094 16892
rect 19094 16836 19098 16892
rect 19034 16832 19098 16836
rect 19114 16892 19178 16896
rect 19114 16836 19118 16892
rect 19118 16836 19174 16892
rect 19174 16836 19178 16892
rect 19114 16832 19178 16836
rect 30822 16892 30886 16896
rect 30822 16836 30826 16892
rect 30826 16836 30882 16892
rect 30882 16836 30886 16892
rect 30822 16832 30886 16836
rect 30902 16892 30966 16896
rect 30902 16836 30906 16892
rect 30906 16836 30962 16892
rect 30962 16836 30966 16892
rect 30902 16832 30966 16836
rect 30982 16892 31046 16896
rect 30982 16836 30986 16892
rect 30986 16836 31042 16892
rect 31042 16836 31046 16892
rect 30982 16832 31046 16836
rect 31062 16892 31126 16896
rect 31062 16836 31066 16892
rect 31066 16836 31122 16892
rect 31122 16836 31126 16892
rect 31062 16832 31126 16836
rect 42770 16892 42834 16896
rect 42770 16836 42774 16892
rect 42774 16836 42830 16892
rect 42830 16836 42834 16892
rect 42770 16832 42834 16836
rect 42850 16892 42914 16896
rect 42850 16836 42854 16892
rect 42854 16836 42910 16892
rect 42910 16836 42914 16892
rect 42850 16832 42914 16836
rect 42930 16892 42994 16896
rect 42930 16836 42934 16892
rect 42934 16836 42990 16892
rect 42990 16836 42994 16892
rect 42930 16832 42994 16836
rect 43010 16892 43074 16896
rect 43010 16836 43014 16892
rect 43014 16836 43070 16892
rect 43070 16836 43074 16892
rect 43010 16832 43074 16836
rect 12900 16348 12964 16352
rect 12900 16292 12904 16348
rect 12904 16292 12960 16348
rect 12960 16292 12964 16348
rect 12900 16288 12964 16292
rect 12980 16348 13044 16352
rect 12980 16292 12984 16348
rect 12984 16292 13040 16348
rect 13040 16292 13044 16348
rect 12980 16288 13044 16292
rect 13060 16348 13124 16352
rect 13060 16292 13064 16348
rect 13064 16292 13120 16348
rect 13120 16292 13124 16348
rect 13060 16288 13124 16292
rect 13140 16348 13204 16352
rect 13140 16292 13144 16348
rect 13144 16292 13200 16348
rect 13200 16292 13204 16348
rect 13140 16288 13204 16292
rect 24848 16348 24912 16352
rect 24848 16292 24852 16348
rect 24852 16292 24908 16348
rect 24908 16292 24912 16348
rect 24848 16288 24912 16292
rect 24928 16348 24992 16352
rect 24928 16292 24932 16348
rect 24932 16292 24988 16348
rect 24988 16292 24992 16348
rect 24928 16288 24992 16292
rect 25008 16348 25072 16352
rect 25008 16292 25012 16348
rect 25012 16292 25068 16348
rect 25068 16292 25072 16348
rect 25008 16288 25072 16292
rect 25088 16348 25152 16352
rect 25088 16292 25092 16348
rect 25092 16292 25148 16348
rect 25148 16292 25152 16348
rect 25088 16288 25152 16292
rect 36796 16348 36860 16352
rect 36796 16292 36800 16348
rect 36800 16292 36856 16348
rect 36856 16292 36860 16348
rect 36796 16288 36860 16292
rect 36876 16348 36940 16352
rect 36876 16292 36880 16348
rect 36880 16292 36936 16348
rect 36936 16292 36940 16348
rect 36876 16288 36940 16292
rect 36956 16348 37020 16352
rect 36956 16292 36960 16348
rect 36960 16292 37016 16348
rect 37016 16292 37020 16348
rect 36956 16288 37020 16292
rect 37036 16348 37100 16352
rect 37036 16292 37040 16348
rect 37040 16292 37096 16348
rect 37096 16292 37100 16348
rect 37036 16288 37100 16292
rect 6926 15804 6990 15808
rect 6926 15748 6930 15804
rect 6930 15748 6986 15804
rect 6986 15748 6990 15804
rect 6926 15744 6990 15748
rect 7006 15804 7070 15808
rect 7006 15748 7010 15804
rect 7010 15748 7066 15804
rect 7066 15748 7070 15804
rect 7006 15744 7070 15748
rect 7086 15804 7150 15808
rect 7086 15748 7090 15804
rect 7090 15748 7146 15804
rect 7146 15748 7150 15804
rect 7086 15744 7150 15748
rect 7166 15804 7230 15808
rect 7166 15748 7170 15804
rect 7170 15748 7226 15804
rect 7226 15748 7230 15804
rect 7166 15744 7230 15748
rect 18874 15804 18938 15808
rect 18874 15748 18878 15804
rect 18878 15748 18934 15804
rect 18934 15748 18938 15804
rect 18874 15744 18938 15748
rect 18954 15804 19018 15808
rect 18954 15748 18958 15804
rect 18958 15748 19014 15804
rect 19014 15748 19018 15804
rect 18954 15744 19018 15748
rect 19034 15804 19098 15808
rect 19034 15748 19038 15804
rect 19038 15748 19094 15804
rect 19094 15748 19098 15804
rect 19034 15744 19098 15748
rect 19114 15804 19178 15808
rect 19114 15748 19118 15804
rect 19118 15748 19174 15804
rect 19174 15748 19178 15804
rect 19114 15744 19178 15748
rect 30822 15804 30886 15808
rect 30822 15748 30826 15804
rect 30826 15748 30882 15804
rect 30882 15748 30886 15804
rect 30822 15744 30886 15748
rect 30902 15804 30966 15808
rect 30902 15748 30906 15804
rect 30906 15748 30962 15804
rect 30962 15748 30966 15804
rect 30902 15744 30966 15748
rect 30982 15804 31046 15808
rect 30982 15748 30986 15804
rect 30986 15748 31042 15804
rect 31042 15748 31046 15804
rect 30982 15744 31046 15748
rect 31062 15804 31126 15808
rect 31062 15748 31066 15804
rect 31066 15748 31122 15804
rect 31122 15748 31126 15804
rect 31062 15744 31126 15748
rect 42770 15804 42834 15808
rect 42770 15748 42774 15804
rect 42774 15748 42830 15804
rect 42830 15748 42834 15804
rect 42770 15744 42834 15748
rect 42850 15804 42914 15808
rect 42850 15748 42854 15804
rect 42854 15748 42910 15804
rect 42910 15748 42914 15804
rect 42850 15744 42914 15748
rect 42930 15804 42994 15808
rect 42930 15748 42934 15804
rect 42934 15748 42990 15804
rect 42990 15748 42994 15804
rect 42930 15744 42994 15748
rect 43010 15804 43074 15808
rect 43010 15748 43014 15804
rect 43014 15748 43070 15804
rect 43070 15748 43074 15804
rect 43010 15744 43074 15748
rect 12900 15260 12964 15264
rect 12900 15204 12904 15260
rect 12904 15204 12960 15260
rect 12960 15204 12964 15260
rect 12900 15200 12964 15204
rect 12980 15260 13044 15264
rect 12980 15204 12984 15260
rect 12984 15204 13040 15260
rect 13040 15204 13044 15260
rect 12980 15200 13044 15204
rect 13060 15260 13124 15264
rect 13060 15204 13064 15260
rect 13064 15204 13120 15260
rect 13120 15204 13124 15260
rect 13060 15200 13124 15204
rect 13140 15260 13204 15264
rect 13140 15204 13144 15260
rect 13144 15204 13200 15260
rect 13200 15204 13204 15260
rect 13140 15200 13204 15204
rect 24848 15260 24912 15264
rect 24848 15204 24852 15260
rect 24852 15204 24908 15260
rect 24908 15204 24912 15260
rect 24848 15200 24912 15204
rect 24928 15260 24992 15264
rect 24928 15204 24932 15260
rect 24932 15204 24988 15260
rect 24988 15204 24992 15260
rect 24928 15200 24992 15204
rect 25008 15260 25072 15264
rect 25008 15204 25012 15260
rect 25012 15204 25068 15260
rect 25068 15204 25072 15260
rect 25008 15200 25072 15204
rect 25088 15260 25152 15264
rect 25088 15204 25092 15260
rect 25092 15204 25148 15260
rect 25148 15204 25152 15260
rect 25088 15200 25152 15204
rect 36796 15260 36860 15264
rect 36796 15204 36800 15260
rect 36800 15204 36856 15260
rect 36856 15204 36860 15260
rect 36796 15200 36860 15204
rect 36876 15260 36940 15264
rect 36876 15204 36880 15260
rect 36880 15204 36936 15260
rect 36936 15204 36940 15260
rect 36876 15200 36940 15204
rect 36956 15260 37020 15264
rect 36956 15204 36960 15260
rect 36960 15204 37016 15260
rect 37016 15204 37020 15260
rect 36956 15200 37020 15204
rect 37036 15260 37100 15264
rect 37036 15204 37040 15260
rect 37040 15204 37096 15260
rect 37096 15204 37100 15260
rect 37036 15200 37100 15204
rect 6926 14716 6990 14720
rect 6926 14660 6930 14716
rect 6930 14660 6986 14716
rect 6986 14660 6990 14716
rect 6926 14656 6990 14660
rect 7006 14716 7070 14720
rect 7006 14660 7010 14716
rect 7010 14660 7066 14716
rect 7066 14660 7070 14716
rect 7006 14656 7070 14660
rect 7086 14716 7150 14720
rect 7086 14660 7090 14716
rect 7090 14660 7146 14716
rect 7146 14660 7150 14716
rect 7086 14656 7150 14660
rect 7166 14716 7230 14720
rect 7166 14660 7170 14716
rect 7170 14660 7226 14716
rect 7226 14660 7230 14716
rect 7166 14656 7230 14660
rect 18874 14716 18938 14720
rect 18874 14660 18878 14716
rect 18878 14660 18934 14716
rect 18934 14660 18938 14716
rect 18874 14656 18938 14660
rect 18954 14716 19018 14720
rect 18954 14660 18958 14716
rect 18958 14660 19014 14716
rect 19014 14660 19018 14716
rect 18954 14656 19018 14660
rect 19034 14716 19098 14720
rect 19034 14660 19038 14716
rect 19038 14660 19094 14716
rect 19094 14660 19098 14716
rect 19034 14656 19098 14660
rect 19114 14716 19178 14720
rect 19114 14660 19118 14716
rect 19118 14660 19174 14716
rect 19174 14660 19178 14716
rect 19114 14656 19178 14660
rect 30822 14716 30886 14720
rect 30822 14660 30826 14716
rect 30826 14660 30882 14716
rect 30882 14660 30886 14716
rect 30822 14656 30886 14660
rect 30902 14716 30966 14720
rect 30902 14660 30906 14716
rect 30906 14660 30962 14716
rect 30962 14660 30966 14716
rect 30902 14656 30966 14660
rect 30982 14716 31046 14720
rect 30982 14660 30986 14716
rect 30986 14660 31042 14716
rect 31042 14660 31046 14716
rect 30982 14656 31046 14660
rect 31062 14716 31126 14720
rect 31062 14660 31066 14716
rect 31066 14660 31122 14716
rect 31122 14660 31126 14716
rect 31062 14656 31126 14660
rect 42770 14716 42834 14720
rect 42770 14660 42774 14716
rect 42774 14660 42830 14716
rect 42830 14660 42834 14716
rect 42770 14656 42834 14660
rect 42850 14716 42914 14720
rect 42850 14660 42854 14716
rect 42854 14660 42910 14716
rect 42910 14660 42914 14716
rect 42850 14656 42914 14660
rect 42930 14716 42994 14720
rect 42930 14660 42934 14716
rect 42934 14660 42990 14716
rect 42990 14660 42994 14716
rect 42930 14656 42994 14660
rect 43010 14716 43074 14720
rect 43010 14660 43014 14716
rect 43014 14660 43070 14716
rect 43070 14660 43074 14716
rect 43010 14656 43074 14660
rect 12900 14172 12964 14176
rect 12900 14116 12904 14172
rect 12904 14116 12960 14172
rect 12960 14116 12964 14172
rect 12900 14112 12964 14116
rect 12980 14172 13044 14176
rect 12980 14116 12984 14172
rect 12984 14116 13040 14172
rect 13040 14116 13044 14172
rect 12980 14112 13044 14116
rect 13060 14172 13124 14176
rect 13060 14116 13064 14172
rect 13064 14116 13120 14172
rect 13120 14116 13124 14172
rect 13060 14112 13124 14116
rect 13140 14172 13204 14176
rect 13140 14116 13144 14172
rect 13144 14116 13200 14172
rect 13200 14116 13204 14172
rect 13140 14112 13204 14116
rect 24848 14172 24912 14176
rect 24848 14116 24852 14172
rect 24852 14116 24908 14172
rect 24908 14116 24912 14172
rect 24848 14112 24912 14116
rect 24928 14172 24992 14176
rect 24928 14116 24932 14172
rect 24932 14116 24988 14172
rect 24988 14116 24992 14172
rect 24928 14112 24992 14116
rect 25008 14172 25072 14176
rect 25008 14116 25012 14172
rect 25012 14116 25068 14172
rect 25068 14116 25072 14172
rect 25008 14112 25072 14116
rect 25088 14172 25152 14176
rect 25088 14116 25092 14172
rect 25092 14116 25148 14172
rect 25148 14116 25152 14172
rect 25088 14112 25152 14116
rect 36796 14172 36860 14176
rect 36796 14116 36800 14172
rect 36800 14116 36856 14172
rect 36856 14116 36860 14172
rect 36796 14112 36860 14116
rect 36876 14172 36940 14176
rect 36876 14116 36880 14172
rect 36880 14116 36936 14172
rect 36936 14116 36940 14172
rect 36876 14112 36940 14116
rect 36956 14172 37020 14176
rect 36956 14116 36960 14172
rect 36960 14116 37016 14172
rect 37016 14116 37020 14172
rect 36956 14112 37020 14116
rect 37036 14172 37100 14176
rect 37036 14116 37040 14172
rect 37040 14116 37096 14172
rect 37096 14116 37100 14172
rect 37036 14112 37100 14116
rect 6926 13628 6990 13632
rect 6926 13572 6930 13628
rect 6930 13572 6986 13628
rect 6986 13572 6990 13628
rect 6926 13568 6990 13572
rect 7006 13628 7070 13632
rect 7006 13572 7010 13628
rect 7010 13572 7066 13628
rect 7066 13572 7070 13628
rect 7006 13568 7070 13572
rect 7086 13628 7150 13632
rect 7086 13572 7090 13628
rect 7090 13572 7146 13628
rect 7146 13572 7150 13628
rect 7086 13568 7150 13572
rect 7166 13628 7230 13632
rect 7166 13572 7170 13628
rect 7170 13572 7226 13628
rect 7226 13572 7230 13628
rect 7166 13568 7230 13572
rect 18874 13628 18938 13632
rect 18874 13572 18878 13628
rect 18878 13572 18934 13628
rect 18934 13572 18938 13628
rect 18874 13568 18938 13572
rect 18954 13628 19018 13632
rect 18954 13572 18958 13628
rect 18958 13572 19014 13628
rect 19014 13572 19018 13628
rect 18954 13568 19018 13572
rect 19034 13628 19098 13632
rect 19034 13572 19038 13628
rect 19038 13572 19094 13628
rect 19094 13572 19098 13628
rect 19034 13568 19098 13572
rect 19114 13628 19178 13632
rect 19114 13572 19118 13628
rect 19118 13572 19174 13628
rect 19174 13572 19178 13628
rect 19114 13568 19178 13572
rect 30822 13628 30886 13632
rect 30822 13572 30826 13628
rect 30826 13572 30882 13628
rect 30882 13572 30886 13628
rect 30822 13568 30886 13572
rect 30902 13628 30966 13632
rect 30902 13572 30906 13628
rect 30906 13572 30962 13628
rect 30962 13572 30966 13628
rect 30902 13568 30966 13572
rect 30982 13628 31046 13632
rect 30982 13572 30986 13628
rect 30986 13572 31042 13628
rect 31042 13572 31046 13628
rect 30982 13568 31046 13572
rect 31062 13628 31126 13632
rect 31062 13572 31066 13628
rect 31066 13572 31122 13628
rect 31122 13572 31126 13628
rect 31062 13568 31126 13572
rect 42770 13628 42834 13632
rect 42770 13572 42774 13628
rect 42774 13572 42830 13628
rect 42830 13572 42834 13628
rect 42770 13568 42834 13572
rect 42850 13628 42914 13632
rect 42850 13572 42854 13628
rect 42854 13572 42910 13628
rect 42910 13572 42914 13628
rect 42850 13568 42914 13572
rect 42930 13628 42994 13632
rect 42930 13572 42934 13628
rect 42934 13572 42990 13628
rect 42990 13572 42994 13628
rect 42930 13568 42994 13572
rect 43010 13628 43074 13632
rect 43010 13572 43014 13628
rect 43014 13572 43070 13628
rect 43070 13572 43074 13628
rect 43010 13568 43074 13572
rect 12900 13084 12964 13088
rect 12900 13028 12904 13084
rect 12904 13028 12960 13084
rect 12960 13028 12964 13084
rect 12900 13024 12964 13028
rect 12980 13084 13044 13088
rect 12980 13028 12984 13084
rect 12984 13028 13040 13084
rect 13040 13028 13044 13084
rect 12980 13024 13044 13028
rect 13060 13084 13124 13088
rect 13060 13028 13064 13084
rect 13064 13028 13120 13084
rect 13120 13028 13124 13084
rect 13060 13024 13124 13028
rect 13140 13084 13204 13088
rect 13140 13028 13144 13084
rect 13144 13028 13200 13084
rect 13200 13028 13204 13084
rect 13140 13024 13204 13028
rect 24848 13084 24912 13088
rect 24848 13028 24852 13084
rect 24852 13028 24908 13084
rect 24908 13028 24912 13084
rect 24848 13024 24912 13028
rect 24928 13084 24992 13088
rect 24928 13028 24932 13084
rect 24932 13028 24988 13084
rect 24988 13028 24992 13084
rect 24928 13024 24992 13028
rect 25008 13084 25072 13088
rect 25008 13028 25012 13084
rect 25012 13028 25068 13084
rect 25068 13028 25072 13084
rect 25008 13024 25072 13028
rect 25088 13084 25152 13088
rect 25088 13028 25092 13084
rect 25092 13028 25148 13084
rect 25148 13028 25152 13084
rect 25088 13024 25152 13028
rect 36796 13084 36860 13088
rect 36796 13028 36800 13084
rect 36800 13028 36856 13084
rect 36856 13028 36860 13084
rect 36796 13024 36860 13028
rect 36876 13084 36940 13088
rect 36876 13028 36880 13084
rect 36880 13028 36936 13084
rect 36936 13028 36940 13084
rect 36876 13024 36940 13028
rect 36956 13084 37020 13088
rect 36956 13028 36960 13084
rect 36960 13028 37016 13084
rect 37016 13028 37020 13084
rect 36956 13024 37020 13028
rect 37036 13084 37100 13088
rect 37036 13028 37040 13084
rect 37040 13028 37096 13084
rect 37096 13028 37100 13084
rect 37036 13024 37100 13028
rect 6926 12540 6990 12544
rect 6926 12484 6930 12540
rect 6930 12484 6986 12540
rect 6986 12484 6990 12540
rect 6926 12480 6990 12484
rect 7006 12540 7070 12544
rect 7006 12484 7010 12540
rect 7010 12484 7066 12540
rect 7066 12484 7070 12540
rect 7006 12480 7070 12484
rect 7086 12540 7150 12544
rect 7086 12484 7090 12540
rect 7090 12484 7146 12540
rect 7146 12484 7150 12540
rect 7086 12480 7150 12484
rect 7166 12540 7230 12544
rect 7166 12484 7170 12540
rect 7170 12484 7226 12540
rect 7226 12484 7230 12540
rect 7166 12480 7230 12484
rect 18874 12540 18938 12544
rect 18874 12484 18878 12540
rect 18878 12484 18934 12540
rect 18934 12484 18938 12540
rect 18874 12480 18938 12484
rect 18954 12540 19018 12544
rect 18954 12484 18958 12540
rect 18958 12484 19014 12540
rect 19014 12484 19018 12540
rect 18954 12480 19018 12484
rect 19034 12540 19098 12544
rect 19034 12484 19038 12540
rect 19038 12484 19094 12540
rect 19094 12484 19098 12540
rect 19034 12480 19098 12484
rect 19114 12540 19178 12544
rect 19114 12484 19118 12540
rect 19118 12484 19174 12540
rect 19174 12484 19178 12540
rect 19114 12480 19178 12484
rect 30822 12540 30886 12544
rect 30822 12484 30826 12540
rect 30826 12484 30882 12540
rect 30882 12484 30886 12540
rect 30822 12480 30886 12484
rect 30902 12540 30966 12544
rect 30902 12484 30906 12540
rect 30906 12484 30962 12540
rect 30962 12484 30966 12540
rect 30902 12480 30966 12484
rect 30982 12540 31046 12544
rect 30982 12484 30986 12540
rect 30986 12484 31042 12540
rect 31042 12484 31046 12540
rect 30982 12480 31046 12484
rect 31062 12540 31126 12544
rect 31062 12484 31066 12540
rect 31066 12484 31122 12540
rect 31122 12484 31126 12540
rect 31062 12480 31126 12484
rect 42770 12540 42834 12544
rect 42770 12484 42774 12540
rect 42774 12484 42830 12540
rect 42830 12484 42834 12540
rect 42770 12480 42834 12484
rect 42850 12540 42914 12544
rect 42850 12484 42854 12540
rect 42854 12484 42910 12540
rect 42910 12484 42914 12540
rect 42850 12480 42914 12484
rect 42930 12540 42994 12544
rect 42930 12484 42934 12540
rect 42934 12484 42990 12540
rect 42990 12484 42994 12540
rect 42930 12480 42994 12484
rect 43010 12540 43074 12544
rect 43010 12484 43014 12540
rect 43014 12484 43070 12540
rect 43070 12484 43074 12540
rect 43010 12480 43074 12484
rect 12900 11996 12964 12000
rect 12900 11940 12904 11996
rect 12904 11940 12960 11996
rect 12960 11940 12964 11996
rect 12900 11936 12964 11940
rect 12980 11996 13044 12000
rect 12980 11940 12984 11996
rect 12984 11940 13040 11996
rect 13040 11940 13044 11996
rect 12980 11936 13044 11940
rect 13060 11996 13124 12000
rect 13060 11940 13064 11996
rect 13064 11940 13120 11996
rect 13120 11940 13124 11996
rect 13060 11936 13124 11940
rect 13140 11996 13204 12000
rect 13140 11940 13144 11996
rect 13144 11940 13200 11996
rect 13200 11940 13204 11996
rect 13140 11936 13204 11940
rect 24848 11996 24912 12000
rect 24848 11940 24852 11996
rect 24852 11940 24908 11996
rect 24908 11940 24912 11996
rect 24848 11936 24912 11940
rect 24928 11996 24992 12000
rect 24928 11940 24932 11996
rect 24932 11940 24988 11996
rect 24988 11940 24992 11996
rect 24928 11936 24992 11940
rect 25008 11996 25072 12000
rect 25008 11940 25012 11996
rect 25012 11940 25068 11996
rect 25068 11940 25072 11996
rect 25008 11936 25072 11940
rect 25088 11996 25152 12000
rect 25088 11940 25092 11996
rect 25092 11940 25148 11996
rect 25148 11940 25152 11996
rect 25088 11936 25152 11940
rect 36796 11996 36860 12000
rect 36796 11940 36800 11996
rect 36800 11940 36856 11996
rect 36856 11940 36860 11996
rect 36796 11936 36860 11940
rect 36876 11996 36940 12000
rect 36876 11940 36880 11996
rect 36880 11940 36936 11996
rect 36936 11940 36940 11996
rect 36876 11936 36940 11940
rect 36956 11996 37020 12000
rect 36956 11940 36960 11996
rect 36960 11940 37016 11996
rect 37016 11940 37020 11996
rect 36956 11936 37020 11940
rect 37036 11996 37100 12000
rect 37036 11940 37040 11996
rect 37040 11940 37096 11996
rect 37096 11940 37100 11996
rect 37036 11936 37100 11940
rect 6926 11452 6990 11456
rect 6926 11396 6930 11452
rect 6930 11396 6986 11452
rect 6986 11396 6990 11452
rect 6926 11392 6990 11396
rect 7006 11452 7070 11456
rect 7006 11396 7010 11452
rect 7010 11396 7066 11452
rect 7066 11396 7070 11452
rect 7006 11392 7070 11396
rect 7086 11452 7150 11456
rect 7086 11396 7090 11452
rect 7090 11396 7146 11452
rect 7146 11396 7150 11452
rect 7086 11392 7150 11396
rect 7166 11452 7230 11456
rect 7166 11396 7170 11452
rect 7170 11396 7226 11452
rect 7226 11396 7230 11452
rect 7166 11392 7230 11396
rect 18874 11452 18938 11456
rect 18874 11396 18878 11452
rect 18878 11396 18934 11452
rect 18934 11396 18938 11452
rect 18874 11392 18938 11396
rect 18954 11452 19018 11456
rect 18954 11396 18958 11452
rect 18958 11396 19014 11452
rect 19014 11396 19018 11452
rect 18954 11392 19018 11396
rect 19034 11452 19098 11456
rect 19034 11396 19038 11452
rect 19038 11396 19094 11452
rect 19094 11396 19098 11452
rect 19034 11392 19098 11396
rect 19114 11452 19178 11456
rect 19114 11396 19118 11452
rect 19118 11396 19174 11452
rect 19174 11396 19178 11452
rect 19114 11392 19178 11396
rect 30822 11452 30886 11456
rect 30822 11396 30826 11452
rect 30826 11396 30882 11452
rect 30882 11396 30886 11452
rect 30822 11392 30886 11396
rect 30902 11452 30966 11456
rect 30902 11396 30906 11452
rect 30906 11396 30962 11452
rect 30962 11396 30966 11452
rect 30902 11392 30966 11396
rect 30982 11452 31046 11456
rect 30982 11396 30986 11452
rect 30986 11396 31042 11452
rect 31042 11396 31046 11452
rect 30982 11392 31046 11396
rect 31062 11452 31126 11456
rect 31062 11396 31066 11452
rect 31066 11396 31122 11452
rect 31122 11396 31126 11452
rect 31062 11392 31126 11396
rect 42770 11452 42834 11456
rect 42770 11396 42774 11452
rect 42774 11396 42830 11452
rect 42830 11396 42834 11452
rect 42770 11392 42834 11396
rect 42850 11452 42914 11456
rect 42850 11396 42854 11452
rect 42854 11396 42910 11452
rect 42910 11396 42914 11452
rect 42850 11392 42914 11396
rect 42930 11452 42994 11456
rect 42930 11396 42934 11452
rect 42934 11396 42990 11452
rect 42990 11396 42994 11452
rect 42930 11392 42994 11396
rect 43010 11452 43074 11456
rect 43010 11396 43014 11452
rect 43014 11396 43070 11452
rect 43070 11396 43074 11452
rect 43010 11392 43074 11396
rect 12900 10908 12964 10912
rect 12900 10852 12904 10908
rect 12904 10852 12960 10908
rect 12960 10852 12964 10908
rect 12900 10848 12964 10852
rect 12980 10908 13044 10912
rect 12980 10852 12984 10908
rect 12984 10852 13040 10908
rect 13040 10852 13044 10908
rect 12980 10848 13044 10852
rect 13060 10908 13124 10912
rect 13060 10852 13064 10908
rect 13064 10852 13120 10908
rect 13120 10852 13124 10908
rect 13060 10848 13124 10852
rect 13140 10908 13204 10912
rect 13140 10852 13144 10908
rect 13144 10852 13200 10908
rect 13200 10852 13204 10908
rect 13140 10848 13204 10852
rect 24848 10908 24912 10912
rect 24848 10852 24852 10908
rect 24852 10852 24908 10908
rect 24908 10852 24912 10908
rect 24848 10848 24912 10852
rect 24928 10908 24992 10912
rect 24928 10852 24932 10908
rect 24932 10852 24988 10908
rect 24988 10852 24992 10908
rect 24928 10848 24992 10852
rect 25008 10908 25072 10912
rect 25008 10852 25012 10908
rect 25012 10852 25068 10908
rect 25068 10852 25072 10908
rect 25008 10848 25072 10852
rect 25088 10908 25152 10912
rect 25088 10852 25092 10908
rect 25092 10852 25148 10908
rect 25148 10852 25152 10908
rect 25088 10848 25152 10852
rect 36796 10908 36860 10912
rect 36796 10852 36800 10908
rect 36800 10852 36856 10908
rect 36856 10852 36860 10908
rect 36796 10848 36860 10852
rect 36876 10908 36940 10912
rect 36876 10852 36880 10908
rect 36880 10852 36936 10908
rect 36936 10852 36940 10908
rect 36876 10848 36940 10852
rect 36956 10908 37020 10912
rect 36956 10852 36960 10908
rect 36960 10852 37016 10908
rect 37016 10852 37020 10908
rect 36956 10848 37020 10852
rect 37036 10908 37100 10912
rect 37036 10852 37040 10908
rect 37040 10852 37096 10908
rect 37096 10852 37100 10908
rect 37036 10848 37100 10852
rect 6926 10364 6990 10368
rect 6926 10308 6930 10364
rect 6930 10308 6986 10364
rect 6986 10308 6990 10364
rect 6926 10304 6990 10308
rect 7006 10364 7070 10368
rect 7006 10308 7010 10364
rect 7010 10308 7066 10364
rect 7066 10308 7070 10364
rect 7006 10304 7070 10308
rect 7086 10364 7150 10368
rect 7086 10308 7090 10364
rect 7090 10308 7146 10364
rect 7146 10308 7150 10364
rect 7086 10304 7150 10308
rect 7166 10364 7230 10368
rect 7166 10308 7170 10364
rect 7170 10308 7226 10364
rect 7226 10308 7230 10364
rect 7166 10304 7230 10308
rect 18874 10364 18938 10368
rect 18874 10308 18878 10364
rect 18878 10308 18934 10364
rect 18934 10308 18938 10364
rect 18874 10304 18938 10308
rect 18954 10364 19018 10368
rect 18954 10308 18958 10364
rect 18958 10308 19014 10364
rect 19014 10308 19018 10364
rect 18954 10304 19018 10308
rect 19034 10364 19098 10368
rect 19034 10308 19038 10364
rect 19038 10308 19094 10364
rect 19094 10308 19098 10364
rect 19034 10304 19098 10308
rect 19114 10364 19178 10368
rect 19114 10308 19118 10364
rect 19118 10308 19174 10364
rect 19174 10308 19178 10364
rect 19114 10304 19178 10308
rect 30822 10364 30886 10368
rect 30822 10308 30826 10364
rect 30826 10308 30882 10364
rect 30882 10308 30886 10364
rect 30822 10304 30886 10308
rect 30902 10364 30966 10368
rect 30902 10308 30906 10364
rect 30906 10308 30962 10364
rect 30962 10308 30966 10364
rect 30902 10304 30966 10308
rect 30982 10364 31046 10368
rect 30982 10308 30986 10364
rect 30986 10308 31042 10364
rect 31042 10308 31046 10364
rect 30982 10304 31046 10308
rect 31062 10364 31126 10368
rect 31062 10308 31066 10364
rect 31066 10308 31122 10364
rect 31122 10308 31126 10364
rect 31062 10304 31126 10308
rect 42770 10364 42834 10368
rect 42770 10308 42774 10364
rect 42774 10308 42830 10364
rect 42830 10308 42834 10364
rect 42770 10304 42834 10308
rect 42850 10364 42914 10368
rect 42850 10308 42854 10364
rect 42854 10308 42910 10364
rect 42910 10308 42914 10364
rect 42850 10304 42914 10308
rect 42930 10364 42994 10368
rect 42930 10308 42934 10364
rect 42934 10308 42990 10364
rect 42990 10308 42994 10364
rect 42930 10304 42994 10308
rect 43010 10364 43074 10368
rect 43010 10308 43014 10364
rect 43014 10308 43070 10364
rect 43070 10308 43074 10364
rect 43010 10304 43074 10308
rect 12900 9820 12964 9824
rect 12900 9764 12904 9820
rect 12904 9764 12960 9820
rect 12960 9764 12964 9820
rect 12900 9760 12964 9764
rect 12980 9820 13044 9824
rect 12980 9764 12984 9820
rect 12984 9764 13040 9820
rect 13040 9764 13044 9820
rect 12980 9760 13044 9764
rect 13060 9820 13124 9824
rect 13060 9764 13064 9820
rect 13064 9764 13120 9820
rect 13120 9764 13124 9820
rect 13060 9760 13124 9764
rect 13140 9820 13204 9824
rect 13140 9764 13144 9820
rect 13144 9764 13200 9820
rect 13200 9764 13204 9820
rect 13140 9760 13204 9764
rect 24848 9820 24912 9824
rect 24848 9764 24852 9820
rect 24852 9764 24908 9820
rect 24908 9764 24912 9820
rect 24848 9760 24912 9764
rect 24928 9820 24992 9824
rect 24928 9764 24932 9820
rect 24932 9764 24988 9820
rect 24988 9764 24992 9820
rect 24928 9760 24992 9764
rect 25008 9820 25072 9824
rect 25008 9764 25012 9820
rect 25012 9764 25068 9820
rect 25068 9764 25072 9820
rect 25008 9760 25072 9764
rect 25088 9820 25152 9824
rect 25088 9764 25092 9820
rect 25092 9764 25148 9820
rect 25148 9764 25152 9820
rect 25088 9760 25152 9764
rect 36796 9820 36860 9824
rect 36796 9764 36800 9820
rect 36800 9764 36856 9820
rect 36856 9764 36860 9820
rect 36796 9760 36860 9764
rect 36876 9820 36940 9824
rect 36876 9764 36880 9820
rect 36880 9764 36936 9820
rect 36936 9764 36940 9820
rect 36876 9760 36940 9764
rect 36956 9820 37020 9824
rect 36956 9764 36960 9820
rect 36960 9764 37016 9820
rect 37016 9764 37020 9820
rect 36956 9760 37020 9764
rect 37036 9820 37100 9824
rect 37036 9764 37040 9820
rect 37040 9764 37096 9820
rect 37096 9764 37100 9820
rect 37036 9760 37100 9764
rect 6926 9276 6990 9280
rect 6926 9220 6930 9276
rect 6930 9220 6986 9276
rect 6986 9220 6990 9276
rect 6926 9216 6990 9220
rect 7006 9276 7070 9280
rect 7006 9220 7010 9276
rect 7010 9220 7066 9276
rect 7066 9220 7070 9276
rect 7006 9216 7070 9220
rect 7086 9276 7150 9280
rect 7086 9220 7090 9276
rect 7090 9220 7146 9276
rect 7146 9220 7150 9276
rect 7086 9216 7150 9220
rect 7166 9276 7230 9280
rect 7166 9220 7170 9276
rect 7170 9220 7226 9276
rect 7226 9220 7230 9276
rect 7166 9216 7230 9220
rect 18874 9276 18938 9280
rect 18874 9220 18878 9276
rect 18878 9220 18934 9276
rect 18934 9220 18938 9276
rect 18874 9216 18938 9220
rect 18954 9276 19018 9280
rect 18954 9220 18958 9276
rect 18958 9220 19014 9276
rect 19014 9220 19018 9276
rect 18954 9216 19018 9220
rect 19034 9276 19098 9280
rect 19034 9220 19038 9276
rect 19038 9220 19094 9276
rect 19094 9220 19098 9276
rect 19034 9216 19098 9220
rect 19114 9276 19178 9280
rect 19114 9220 19118 9276
rect 19118 9220 19174 9276
rect 19174 9220 19178 9276
rect 19114 9216 19178 9220
rect 30822 9276 30886 9280
rect 30822 9220 30826 9276
rect 30826 9220 30882 9276
rect 30882 9220 30886 9276
rect 30822 9216 30886 9220
rect 30902 9276 30966 9280
rect 30902 9220 30906 9276
rect 30906 9220 30962 9276
rect 30962 9220 30966 9276
rect 30902 9216 30966 9220
rect 30982 9276 31046 9280
rect 30982 9220 30986 9276
rect 30986 9220 31042 9276
rect 31042 9220 31046 9276
rect 30982 9216 31046 9220
rect 31062 9276 31126 9280
rect 31062 9220 31066 9276
rect 31066 9220 31122 9276
rect 31122 9220 31126 9276
rect 31062 9216 31126 9220
rect 42770 9276 42834 9280
rect 42770 9220 42774 9276
rect 42774 9220 42830 9276
rect 42830 9220 42834 9276
rect 42770 9216 42834 9220
rect 42850 9276 42914 9280
rect 42850 9220 42854 9276
rect 42854 9220 42910 9276
rect 42910 9220 42914 9276
rect 42850 9216 42914 9220
rect 42930 9276 42994 9280
rect 42930 9220 42934 9276
rect 42934 9220 42990 9276
rect 42990 9220 42994 9276
rect 42930 9216 42994 9220
rect 43010 9276 43074 9280
rect 43010 9220 43014 9276
rect 43014 9220 43070 9276
rect 43070 9220 43074 9276
rect 43010 9216 43074 9220
rect 12900 8732 12964 8736
rect 12900 8676 12904 8732
rect 12904 8676 12960 8732
rect 12960 8676 12964 8732
rect 12900 8672 12964 8676
rect 12980 8732 13044 8736
rect 12980 8676 12984 8732
rect 12984 8676 13040 8732
rect 13040 8676 13044 8732
rect 12980 8672 13044 8676
rect 13060 8732 13124 8736
rect 13060 8676 13064 8732
rect 13064 8676 13120 8732
rect 13120 8676 13124 8732
rect 13060 8672 13124 8676
rect 13140 8732 13204 8736
rect 13140 8676 13144 8732
rect 13144 8676 13200 8732
rect 13200 8676 13204 8732
rect 13140 8672 13204 8676
rect 24848 8732 24912 8736
rect 24848 8676 24852 8732
rect 24852 8676 24908 8732
rect 24908 8676 24912 8732
rect 24848 8672 24912 8676
rect 24928 8732 24992 8736
rect 24928 8676 24932 8732
rect 24932 8676 24988 8732
rect 24988 8676 24992 8732
rect 24928 8672 24992 8676
rect 25008 8732 25072 8736
rect 25008 8676 25012 8732
rect 25012 8676 25068 8732
rect 25068 8676 25072 8732
rect 25008 8672 25072 8676
rect 25088 8732 25152 8736
rect 25088 8676 25092 8732
rect 25092 8676 25148 8732
rect 25148 8676 25152 8732
rect 25088 8672 25152 8676
rect 36796 8732 36860 8736
rect 36796 8676 36800 8732
rect 36800 8676 36856 8732
rect 36856 8676 36860 8732
rect 36796 8672 36860 8676
rect 36876 8732 36940 8736
rect 36876 8676 36880 8732
rect 36880 8676 36936 8732
rect 36936 8676 36940 8732
rect 36876 8672 36940 8676
rect 36956 8732 37020 8736
rect 36956 8676 36960 8732
rect 36960 8676 37016 8732
rect 37016 8676 37020 8732
rect 36956 8672 37020 8676
rect 37036 8732 37100 8736
rect 37036 8676 37040 8732
rect 37040 8676 37096 8732
rect 37096 8676 37100 8732
rect 37036 8672 37100 8676
rect 6926 8188 6990 8192
rect 6926 8132 6930 8188
rect 6930 8132 6986 8188
rect 6986 8132 6990 8188
rect 6926 8128 6990 8132
rect 7006 8188 7070 8192
rect 7006 8132 7010 8188
rect 7010 8132 7066 8188
rect 7066 8132 7070 8188
rect 7006 8128 7070 8132
rect 7086 8188 7150 8192
rect 7086 8132 7090 8188
rect 7090 8132 7146 8188
rect 7146 8132 7150 8188
rect 7086 8128 7150 8132
rect 7166 8188 7230 8192
rect 7166 8132 7170 8188
rect 7170 8132 7226 8188
rect 7226 8132 7230 8188
rect 7166 8128 7230 8132
rect 18874 8188 18938 8192
rect 18874 8132 18878 8188
rect 18878 8132 18934 8188
rect 18934 8132 18938 8188
rect 18874 8128 18938 8132
rect 18954 8188 19018 8192
rect 18954 8132 18958 8188
rect 18958 8132 19014 8188
rect 19014 8132 19018 8188
rect 18954 8128 19018 8132
rect 19034 8188 19098 8192
rect 19034 8132 19038 8188
rect 19038 8132 19094 8188
rect 19094 8132 19098 8188
rect 19034 8128 19098 8132
rect 19114 8188 19178 8192
rect 19114 8132 19118 8188
rect 19118 8132 19174 8188
rect 19174 8132 19178 8188
rect 19114 8128 19178 8132
rect 30822 8188 30886 8192
rect 30822 8132 30826 8188
rect 30826 8132 30882 8188
rect 30882 8132 30886 8188
rect 30822 8128 30886 8132
rect 30902 8188 30966 8192
rect 30902 8132 30906 8188
rect 30906 8132 30962 8188
rect 30962 8132 30966 8188
rect 30902 8128 30966 8132
rect 30982 8188 31046 8192
rect 30982 8132 30986 8188
rect 30986 8132 31042 8188
rect 31042 8132 31046 8188
rect 30982 8128 31046 8132
rect 31062 8188 31126 8192
rect 31062 8132 31066 8188
rect 31066 8132 31122 8188
rect 31122 8132 31126 8188
rect 31062 8128 31126 8132
rect 42770 8188 42834 8192
rect 42770 8132 42774 8188
rect 42774 8132 42830 8188
rect 42830 8132 42834 8188
rect 42770 8128 42834 8132
rect 42850 8188 42914 8192
rect 42850 8132 42854 8188
rect 42854 8132 42910 8188
rect 42910 8132 42914 8188
rect 42850 8128 42914 8132
rect 42930 8188 42994 8192
rect 42930 8132 42934 8188
rect 42934 8132 42990 8188
rect 42990 8132 42994 8188
rect 42930 8128 42994 8132
rect 43010 8188 43074 8192
rect 43010 8132 43014 8188
rect 43014 8132 43070 8188
rect 43070 8132 43074 8188
rect 43010 8128 43074 8132
rect 12900 7644 12964 7648
rect 12900 7588 12904 7644
rect 12904 7588 12960 7644
rect 12960 7588 12964 7644
rect 12900 7584 12964 7588
rect 12980 7644 13044 7648
rect 12980 7588 12984 7644
rect 12984 7588 13040 7644
rect 13040 7588 13044 7644
rect 12980 7584 13044 7588
rect 13060 7644 13124 7648
rect 13060 7588 13064 7644
rect 13064 7588 13120 7644
rect 13120 7588 13124 7644
rect 13060 7584 13124 7588
rect 13140 7644 13204 7648
rect 13140 7588 13144 7644
rect 13144 7588 13200 7644
rect 13200 7588 13204 7644
rect 13140 7584 13204 7588
rect 24848 7644 24912 7648
rect 24848 7588 24852 7644
rect 24852 7588 24908 7644
rect 24908 7588 24912 7644
rect 24848 7584 24912 7588
rect 24928 7644 24992 7648
rect 24928 7588 24932 7644
rect 24932 7588 24988 7644
rect 24988 7588 24992 7644
rect 24928 7584 24992 7588
rect 25008 7644 25072 7648
rect 25008 7588 25012 7644
rect 25012 7588 25068 7644
rect 25068 7588 25072 7644
rect 25008 7584 25072 7588
rect 25088 7644 25152 7648
rect 25088 7588 25092 7644
rect 25092 7588 25148 7644
rect 25148 7588 25152 7644
rect 25088 7584 25152 7588
rect 36796 7644 36860 7648
rect 36796 7588 36800 7644
rect 36800 7588 36856 7644
rect 36856 7588 36860 7644
rect 36796 7584 36860 7588
rect 36876 7644 36940 7648
rect 36876 7588 36880 7644
rect 36880 7588 36936 7644
rect 36936 7588 36940 7644
rect 36876 7584 36940 7588
rect 36956 7644 37020 7648
rect 36956 7588 36960 7644
rect 36960 7588 37016 7644
rect 37016 7588 37020 7644
rect 36956 7584 37020 7588
rect 37036 7644 37100 7648
rect 37036 7588 37040 7644
rect 37040 7588 37096 7644
rect 37096 7588 37100 7644
rect 37036 7584 37100 7588
rect 6926 7100 6990 7104
rect 6926 7044 6930 7100
rect 6930 7044 6986 7100
rect 6986 7044 6990 7100
rect 6926 7040 6990 7044
rect 7006 7100 7070 7104
rect 7006 7044 7010 7100
rect 7010 7044 7066 7100
rect 7066 7044 7070 7100
rect 7006 7040 7070 7044
rect 7086 7100 7150 7104
rect 7086 7044 7090 7100
rect 7090 7044 7146 7100
rect 7146 7044 7150 7100
rect 7086 7040 7150 7044
rect 7166 7100 7230 7104
rect 7166 7044 7170 7100
rect 7170 7044 7226 7100
rect 7226 7044 7230 7100
rect 7166 7040 7230 7044
rect 18874 7100 18938 7104
rect 18874 7044 18878 7100
rect 18878 7044 18934 7100
rect 18934 7044 18938 7100
rect 18874 7040 18938 7044
rect 18954 7100 19018 7104
rect 18954 7044 18958 7100
rect 18958 7044 19014 7100
rect 19014 7044 19018 7100
rect 18954 7040 19018 7044
rect 19034 7100 19098 7104
rect 19034 7044 19038 7100
rect 19038 7044 19094 7100
rect 19094 7044 19098 7100
rect 19034 7040 19098 7044
rect 19114 7100 19178 7104
rect 19114 7044 19118 7100
rect 19118 7044 19174 7100
rect 19174 7044 19178 7100
rect 19114 7040 19178 7044
rect 30822 7100 30886 7104
rect 30822 7044 30826 7100
rect 30826 7044 30882 7100
rect 30882 7044 30886 7100
rect 30822 7040 30886 7044
rect 30902 7100 30966 7104
rect 30902 7044 30906 7100
rect 30906 7044 30962 7100
rect 30962 7044 30966 7100
rect 30902 7040 30966 7044
rect 30982 7100 31046 7104
rect 30982 7044 30986 7100
rect 30986 7044 31042 7100
rect 31042 7044 31046 7100
rect 30982 7040 31046 7044
rect 31062 7100 31126 7104
rect 31062 7044 31066 7100
rect 31066 7044 31122 7100
rect 31122 7044 31126 7100
rect 31062 7040 31126 7044
rect 42770 7100 42834 7104
rect 42770 7044 42774 7100
rect 42774 7044 42830 7100
rect 42830 7044 42834 7100
rect 42770 7040 42834 7044
rect 42850 7100 42914 7104
rect 42850 7044 42854 7100
rect 42854 7044 42910 7100
rect 42910 7044 42914 7100
rect 42850 7040 42914 7044
rect 42930 7100 42994 7104
rect 42930 7044 42934 7100
rect 42934 7044 42990 7100
rect 42990 7044 42994 7100
rect 42930 7040 42994 7044
rect 43010 7100 43074 7104
rect 43010 7044 43014 7100
rect 43014 7044 43070 7100
rect 43070 7044 43074 7100
rect 43010 7040 43074 7044
rect 12900 6556 12964 6560
rect 12900 6500 12904 6556
rect 12904 6500 12960 6556
rect 12960 6500 12964 6556
rect 12900 6496 12964 6500
rect 12980 6556 13044 6560
rect 12980 6500 12984 6556
rect 12984 6500 13040 6556
rect 13040 6500 13044 6556
rect 12980 6496 13044 6500
rect 13060 6556 13124 6560
rect 13060 6500 13064 6556
rect 13064 6500 13120 6556
rect 13120 6500 13124 6556
rect 13060 6496 13124 6500
rect 13140 6556 13204 6560
rect 13140 6500 13144 6556
rect 13144 6500 13200 6556
rect 13200 6500 13204 6556
rect 13140 6496 13204 6500
rect 24848 6556 24912 6560
rect 24848 6500 24852 6556
rect 24852 6500 24908 6556
rect 24908 6500 24912 6556
rect 24848 6496 24912 6500
rect 24928 6556 24992 6560
rect 24928 6500 24932 6556
rect 24932 6500 24988 6556
rect 24988 6500 24992 6556
rect 24928 6496 24992 6500
rect 25008 6556 25072 6560
rect 25008 6500 25012 6556
rect 25012 6500 25068 6556
rect 25068 6500 25072 6556
rect 25008 6496 25072 6500
rect 25088 6556 25152 6560
rect 25088 6500 25092 6556
rect 25092 6500 25148 6556
rect 25148 6500 25152 6556
rect 25088 6496 25152 6500
rect 36796 6556 36860 6560
rect 36796 6500 36800 6556
rect 36800 6500 36856 6556
rect 36856 6500 36860 6556
rect 36796 6496 36860 6500
rect 36876 6556 36940 6560
rect 36876 6500 36880 6556
rect 36880 6500 36936 6556
rect 36936 6500 36940 6556
rect 36876 6496 36940 6500
rect 36956 6556 37020 6560
rect 36956 6500 36960 6556
rect 36960 6500 37016 6556
rect 37016 6500 37020 6556
rect 36956 6496 37020 6500
rect 37036 6556 37100 6560
rect 37036 6500 37040 6556
rect 37040 6500 37096 6556
rect 37096 6500 37100 6556
rect 37036 6496 37100 6500
rect 6926 6012 6990 6016
rect 6926 5956 6930 6012
rect 6930 5956 6986 6012
rect 6986 5956 6990 6012
rect 6926 5952 6990 5956
rect 7006 6012 7070 6016
rect 7006 5956 7010 6012
rect 7010 5956 7066 6012
rect 7066 5956 7070 6012
rect 7006 5952 7070 5956
rect 7086 6012 7150 6016
rect 7086 5956 7090 6012
rect 7090 5956 7146 6012
rect 7146 5956 7150 6012
rect 7086 5952 7150 5956
rect 7166 6012 7230 6016
rect 7166 5956 7170 6012
rect 7170 5956 7226 6012
rect 7226 5956 7230 6012
rect 7166 5952 7230 5956
rect 18874 6012 18938 6016
rect 18874 5956 18878 6012
rect 18878 5956 18934 6012
rect 18934 5956 18938 6012
rect 18874 5952 18938 5956
rect 18954 6012 19018 6016
rect 18954 5956 18958 6012
rect 18958 5956 19014 6012
rect 19014 5956 19018 6012
rect 18954 5952 19018 5956
rect 19034 6012 19098 6016
rect 19034 5956 19038 6012
rect 19038 5956 19094 6012
rect 19094 5956 19098 6012
rect 19034 5952 19098 5956
rect 19114 6012 19178 6016
rect 19114 5956 19118 6012
rect 19118 5956 19174 6012
rect 19174 5956 19178 6012
rect 19114 5952 19178 5956
rect 30822 6012 30886 6016
rect 30822 5956 30826 6012
rect 30826 5956 30882 6012
rect 30882 5956 30886 6012
rect 30822 5952 30886 5956
rect 30902 6012 30966 6016
rect 30902 5956 30906 6012
rect 30906 5956 30962 6012
rect 30962 5956 30966 6012
rect 30902 5952 30966 5956
rect 30982 6012 31046 6016
rect 30982 5956 30986 6012
rect 30986 5956 31042 6012
rect 31042 5956 31046 6012
rect 30982 5952 31046 5956
rect 31062 6012 31126 6016
rect 31062 5956 31066 6012
rect 31066 5956 31122 6012
rect 31122 5956 31126 6012
rect 31062 5952 31126 5956
rect 42770 6012 42834 6016
rect 42770 5956 42774 6012
rect 42774 5956 42830 6012
rect 42830 5956 42834 6012
rect 42770 5952 42834 5956
rect 42850 6012 42914 6016
rect 42850 5956 42854 6012
rect 42854 5956 42910 6012
rect 42910 5956 42914 6012
rect 42850 5952 42914 5956
rect 42930 6012 42994 6016
rect 42930 5956 42934 6012
rect 42934 5956 42990 6012
rect 42990 5956 42994 6012
rect 42930 5952 42994 5956
rect 43010 6012 43074 6016
rect 43010 5956 43014 6012
rect 43014 5956 43070 6012
rect 43070 5956 43074 6012
rect 43010 5952 43074 5956
rect 12900 5468 12964 5472
rect 12900 5412 12904 5468
rect 12904 5412 12960 5468
rect 12960 5412 12964 5468
rect 12900 5408 12964 5412
rect 12980 5468 13044 5472
rect 12980 5412 12984 5468
rect 12984 5412 13040 5468
rect 13040 5412 13044 5468
rect 12980 5408 13044 5412
rect 13060 5468 13124 5472
rect 13060 5412 13064 5468
rect 13064 5412 13120 5468
rect 13120 5412 13124 5468
rect 13060 5408 13124 5412
rect 13140 5468 13204 5472
rect 13140 5412 13144 5468
rect 13144 5412 13200 5468
rect 13200 5412 13204 5468
rect 13140 5408 13204 5412
rect 24848 5468 24912 5472
rect 24848 5412 24852 5468
rect 24852 5412 24908 5468
rect 24908 5412 24912 5468
rect 24848 5408 24912 5412
rect 24928 5468 24992 5472
rect 24928 5412 24932 5468
rect 24932 5412 24988 5468
rect 24988 5412 24992 5468
rect 24928 5408 24992 5412
rect 25008 5468 25072 5472
rect 25008 5412 25012 5468
rect 25012 5412 25068 5468
rect 25068 5412 25072 5468
rect 25008 5408 25072 5412
rect 25088 5468 25152 5472
rect 25088 5412 25092 5468
rect 25092 5412 25148 5468
rect 25148 5412 25152 5468
rect 25088 5408 25152 5412
rect 36796 5468 36860 5472
rect 36796 5412 36800 5468
rect 36800 5412 36856 5468
rect 36856 5412 36860 5468
rect 36796 5408 36860 5412
rect 36876 5468 36940 5472
rect 36876 5412 36880 5468
rect 36880 5412 36936 5468
rect 36936 5412 36940 5468
rect 36876 5408 36940 5412
rect 36956 5468 37020 5472
rect 36956 5412 36960 5468
rect 36960 5412 37016 5468
rect 37016 5412 37020 5468
rect 36956 5408 37020 5412
rect 37036 5468 37100 5472
rect 37036 5412 37040 5468
rect 37040 5412 37096 5468
rect 37096 5412 37100 5468
rect 37036 5408 37100 5412
rect 6926 4924 6990 4928
rect 6926 4868 6930 4924
rect 6930 4868 6986 4924
rect 6986 4868 6990 4924
rect 6926 4864 6990 4868
rect 7006 4924 7070 4928
rect 7006 4868 7010 4924
rect 7010 4868 7066 4924
rect 7066 4868 7070 4924
rect 7006 4864 7070 4868
rect 7086 4924 7150 4928
rect 7086 4868 7090 4924
rect 7090 4868 7146 4924
rect 7146 4868 7150 4924
rect 7086 4864 7150 4868
rect 7166 4924 7230 4928
rect 7166 4868 7170 4924
rect 7170 4868 7226 4924
rect 7226 4868 7230 4924
rect 7166 4864 7230 4868
rect 18874 4924 18938 4928
rect 18874 4868 18878 4924
rect 18878 4868 18934 4924
rect 18934 4868 18938 4924
rect 18874 4864 18938 4868
rect 18954 4924 19018 4928
rect 18954 4868 18958 4924
rect 18958 4868 19014 4924
rect 19014 4868 19018 4924
rect 18954 4864 19018 4868
rect 19034 4924 19098 4928
rect 19034 4868 19038 4924
rect 19038 4868 19094 4924
rect 19094 4868 19098 4924
rect 19034 4864 19098 4868
rect 19114 4924 19178 4928
rect 19114 4868 19118 4924
rect 19118 4868 19174 4924
rect 19174 4868 19178 4924
rect 19114 4864 19178 4868
rect 30822 4924 30886 4928
rect 30822 4868 30826 4924
rect 30826 4868 30882 4924
rect 30882 4868 30886 4924
rect 30822 4864 30886 4868
rect 30902 4924 30966 4928
rect 30902 4868 30906 4924
rect 30906 4868 30962 4924
rect 30962 4868 30966 4924
rect 30902 4864 30966 4868
rect 30982 4924 31046 4928
rect 30982 4868 30986 4924
rect 30986 4868 31042 4924
rect 31042 4868 31046 4924
rect 30982 4864 31046 4868
rect 31062 4924 31126 4928
rect 31062 4868 31066 4924
rect 31066 4868 31122 4924
rect 31122 4868 31126 4924
rect 31062 4864 31126 4868
rect 42770 4924 42834 4928
rect 42770 4868 42774 4924
rect 42774 4868 42830 4924
rect 42830 4868 42834 4924
rect 42770 4864 42834 4868
rect 42850 4924 42914 4928
rect 42850 4868 42854 4924
rect 42854 4868 42910 4924
rect 42910 4868 42914 4924
rect 42850 4864 42914 4868
rect 42930 4924 42994 4928
rect 42930 4868 42934 4924
rect 42934 4868 42990 4924
rect 42990 4868 42994 4924
rect 42930 4864 42994 4868
rect 43010 4924 43074 4928
rect 43010 4868 43014 4924
rect 43014 4868 43070 4924
rect 43070 4868 43074 4924
rect 43010 4864 43074 4868
rect 12900 4380 12964 4384
rect 12900 4324 12904 4380
rect 12904 4324 12960 4380
rect 12960 4324 12964 4380
rect 12900 4320 12964 4324
rect 12980 4380 13044 4384
rect 12980 4324 12984 4380
rect 12984 4324 13040 4380
rect 13040 4324 13044 4380
rect 12980 4320 13044 4324
rect 13060 4380 13124 4384
rect 13060 4324 13064 4380
rect 13064 4324 13120 4380
rect 13120 4324 13124 4380
rect 13060 4320 13124 4324
rect 13140 4380 13204 4384
rect 13140 4324 13144 4380
rect 13144 4324 13200 4380
rect 13200 4324 13204 4380
rect 13140 4320 13204 4324
rect 24848 4380 24912 4384
rect 24848 4324 24852 4380
rect 24852 4324 24908 4380
rect 24908 4324 24912 4380
rect 24848 4320 24912 4324
rect 24928 4380 24992 4384
rect 24928 4324 24932 4380
rect 24932 4324 24988 4380
rect 24988 4324 24992 4380
rect 24928 4320 24992 4324
rect 25008 4380 25072 4384
rect 25008 4324 25012 4380
rect 25012 4324 25068 4380
rect 25068 4324 25072 4380
rect 25008 4320 25072 4324
rect 25088 4380 25152 4384
rect 25088 4324 25092 4380
rect 25092 4324 25148 4380
rect 25148 4324 25152 4380
rect 25088 4320 25152 4324
rect 36796 4380 36860 4384
rect 36796 4324 36800 4380
rect 36800 4324 36856 4380
rect 36856 4324 36860 4380
rect 36796 4320 36860 4324
rect 36876 4380 36940 4384
rect 36876 4324 36880 4380
rect 36880 4324 36936 4380
rect 36936 4324 36940 4380
rect 36876 4320 36940 4324
rect 36956 4380 37020 4384
rect 36956 4324 36960 4380
rect 36960 4324 37016 4380
rect 37016 4324 37020 4380
rect 36956 4320 37020 4324
rect 37036 4380 37100 4384
rect 37036 4324 37040 4380
rect 37040 4324 37096 4380
rect 37096 4324 37100 4380
rect 37036 4320 37100 4324
rect 6926 3836 6990 3840
rect 6926 3780 6930 3836
rect 6930 3780 6986 3836
rect 6986 3780 6990 3836
rect 6926 3776 6990 3780
rect 7006 3836 7070 3840
rect 7006 3780 7010 3836
rect 7010 3780 7066 3836
rect 7066 3780 7070 3836
rect 7006 3776 7070 3780
rect 7086 3836 7150 3840
rect 7086 3780 7090 3836
rect 7090 3780 7146 3836
rect 7146 3780 7150 3836
rect 7086 3776 7150 3780
rect 7166 3836 7230 3840
rect 7166 3780 7170 3836
rect 7170 3780 7226 3836
rect 7226 3780 7230 3836
rect 7166 3776 7230 3780
rect 18874 3836 18938 3840
rect 18874 3780 18878 3836
rect 18878 3780 18934 3836
rect 18934 3780 18938 3836
rect 18874 3776 18938 3780
rect 18954 3836 19018 3840
rect 18954 3780 18958 3836
rect 18958 3780 19014 3836
rect 19014 3780 19018 3836
rect 18954 3776 19018 3780
rect 19034 3836 19098 3840
rect 19034 3780 19038 3836
rect 19038 3780 19094 3836
rect 19094 3780 19098 3836
rect 19034 3776 19098 3780
rect 19114 3836 19178 3840
rect 19114 3780 19118 3836
rect 19118 3780 19174 3836
rect 19174 3780 19178 3836
rect 19114 3776 19178 3780
rect 30822 3836 30886 3840
rect 30822 3780 30826 3836
rect 30826 3780 30882 3836
rect 30882 3780 30886 3836
rect 30822 3776 30886 3780
rect 30902 3836 30966 3840
rect 30902 3780 30906 3836
rect 30906 3780 30962 3836
rect 30962 3780 30966 3836
rect 30902 3776 30966 3780
rect 30982 3836 31046 3840
rect 30982 3780 30986 3836
rect 30986 3780 31042 3836
rect 31042 3780 31046 3836
rect 30982 3776 31046 3780
rect 31062 3836 31126 3840
rect 31062 3780 31066 3836
rect 31066 3780 31122 3836
rect 31122 3780 31126 3836
rect 31062 3776 31126 3780
rect 42770 3836 42834 3840
rect 42770 3780 42774 3836
rect 42774 3780 42830 3836
rect 42830 3780 42834 3836
rect 42770 3776 42834 3780
rect 42850 3836 42914 3840
rect 42850 3780 42854 3836
rect 42854 3780 42910 3836
rect 42910 3780 42914 3836
rect 42850 3776 42914 3780
rect 42930 3836 42994 3840
rect 42930 3780 42934 3836
rect 42934 3780 42990 3836
rect 42990 3780 42994 3836
rect 42930 3776 42994 3780
rect 43010 3836 43074 3840
rect 43010 3780 43014 3836
rect 43014 3780 43070 3836
rect 43070 3780 43074 3836
rect 43010 3776 43074 3780
rect 12900 3292 12964 3296
rect 12900 3236 12904 3292
rect 12904 3236 12960 3292
rect 12960 3236 12964 3292
rect 12900 3232 12964 3236
rect 12980 3292 13044 3296
rect 12980 3236 12984 3292
rect 12984 3236 13040 3292
rect 13040 3236 13044 3292
rect 12980 3232 13044 3236
rect 13060 3292 13124 3296
rect 13060 3236 13064 3292
rect 13064 3236 13120 3292
rect 13120 3236 13124 3292
rect 13060 3232 13124 3236
rect 13140 3292 13204 3296
rect 13140 3236 13144 3292
rect 13144 3236 13200 3292
rect 13200 3236 13204 3292
rect 13140 3232 13204 3236
rect 24848 3292 24912 3296
rect 24848 3236 24852 3292
rect 24852 3236 24908 3292
rect 24908 3236 24912 3292
rect 24848 3232 24912 3236
rect 24928 3292 24992 3296
rect 24928 3236 24932 3292
rect 24932 3236 24988 3292
rect 24988 3236 24992 3292
rect 24928 3232 24992 3236
rect 25008 3292 25072 3296
rect 25008 3236 25012 3292
rect 25012 3236 25068 3292
rect 25068 3236 25072 3292
rect 25008 3232 25072 3236
rect 25088 3292 25152 3296
rect 25088 3236 25092 3292
rect 25092 3236 25148 3292
rect 25148 3236 25152 3292
rect 25088 3232 25152 3236
rect 36796 3292 36860 3296
rect 36796 3236 36800 3292
rect 36800 3236 36856 3292
rect 36856 3236 36860 3292
rect 36796 3232 36860 3236
rect 36876 3292 36940 3296
rect 36876 3236 36880 3292
rect 36880 3236 36936 3292
rect 36936 3236 36940 3292
rect 36876 3232 36940 3236
rect 36956 3292 37020 3296
rect 36956 3236 36960 3292
rect 36960 3236 37016 3292
rect 37016 3236 37020 3292
rect 36956 3232 37020 3236
rect 37036 3292 37100 3296
rect 37036 3236 37040 3292
rect 37040 3236 37096 3292
rect 37096 3236 37100 3292
rect 37036 3232 37100 3236
rect 6926 2748 6990 2752
rect 6926 2692 6930 2748
rect 6930 2692 6986 2748
rect 6986 2692 6990 2748
rect 6926 2688 6990 2692
rect 7006 2748 7070 2752
rect 7006 2692 7010 2748
rect 7010 2692 7066 2748
rect 7066 2692 7070 2748
rect 7006 2688 7070 2692
rect 7086 2748 7150 2752
rect 7086 2692 7090 2748
rect 7090 2692 7146 2748
rect 7146 2692 7150 2748
rect 7086 2688 7150 2692
rect 7166 2748 7230 2752
rect 7166 2692 7170 2748
rect 7170 2692 7226 2748
rect 7226 2692 7230 2748
rect 7166 2688 7230 2692
rect 18874 2748 18938 2752
rect 18874 2692 18878 2748
rect 18878 2692 18934 2748
rect 18934 2692 18938 2748
rect 18874 2688 18938 2692
rect 18954 2748 19018 2752
rect 18954 2692 18958 2748
rect 18958 2692 19014 2748
rect 19014 2692 19018 2748
rect 18954 2688 19018 2692
rect 19034 2748 19098 2752
rect 19034 2692 19038 2748
rect 19038 2692 19094 2748
rect 19094 2692 19098 2748
rect 19034 2688 19098 2692
rect 19114 2748 19178 2752
rect 19114 2692 19118 2748
rect 19118 2692 19174 2748
rect 19174 2692 19178 2748
rect 19114 2688 19178 2692
rect 30822 2748 30886 2752
rect 30822 2692 30826 2748
rect 30826 2692 30882 2748
rect 30882 2692 30886 2748
rect 30822 2688 30886 2692
rect 30902 2748 30966 2752
rect 30902 2692 30906 2748
rect 30906 2692 30962 2748
rect 30962 2692 30966 2748
rect 30902 2688 30966 2692
rect 30982 2748 31046 2752
rect 30982 2692 30986 2748
rect 30986 2692 31042 2748
rect 31042 2692 31046 2748
rect 30982 2688 31046 2692
rect 31062 2748 31126 2752
rect 31062 2692 31066 2748
rect 31066 2692 31122 2748
rect 31122 2692 31126 2748
rect 31062 2688 31126 2692
rect 42770 2748 42834 2752
rect 42770 2692 42774 2748
rect 42774 2692 42830 2748
rect 42830 2692 42834 2748
rect 42770 2688 42834 2692
rect 42850 2748 42914 2752
rect 42850 2692 42854 2748
rect 42854 2692 42910 2748
rect 42910 2692 42914 2748
rect 42850 2688 42914 2692
rect 42930 2748 42994 2752
rect 42930 2692 42934 2748
rect 42934 2692 42990 2748
rect 42990 2692 42994 2748
rect 42930 2688 42994 2692
rect 43010 2748 43074 2752
rect 43010 2692 43014 2748
rect 43014 2692 43070 2748
rect 43070 2692 43074 2748
rect 43010 2688 43074 2692
rect 12900 2204 12964 2208
rect 12900 2148 12904 2204
rect 12904 2148 12960 2204
rect 12960 2148 12964 2204
rect 12900 2144 12964 2148
rect 12980 2204 13044 2208
rect 12980 2148 12984 2204
rect 12984 2148 13040 2204
rect 13040 2148 13044 2204
rect 12980 2144 13044 2148
rect 13060 2204 13124 2208
rect 13060 2148 13064 2204
rect 13064 2148 13120 2204
rect 13120 2148 13124 2204
rect 13060 2144 13124 2148
rect 13140 2204 13204 2208
rect 13140 2148 13144 2204
rect 13144 2148 13200 2204
rect 13200 2148 13204 2204
rect 13140 2144 13204 2148
rect 24848 2204 24912 2208
rect 24848 2148 24852 2204
rect 24852 2148 24908 2204
rect 24908 2148 24912 2204
rect 24848 2144 24912 2148
rect 24928 2204 24992 2208
rect 24928 2148 24932 2204
rect 24932 2148 24988 2204
rect 24988 2148 24992 2204
rect 24928 2144 24992 2148
rect 25008 2204 25072 2208
rect 25008 2148 25012 2204
rect 25012 2148 25068 2204
rect 25068 2148 25072 2204
rect 25008 2144 25072 2148
rect 25088 2204 25152 2208
rect 25088 2148 25092 2204
rect 25092 2148 25148 2204
rect 25148 2148 25152 2204
rect 25088 2144 25152 2148
rect 36796 2204 36860 2208
rect 36796 2148 36800 2204
rect 36800 2148 36856 2204
rect 36856 2148 36860 2204
rect 36796 2144 36860 2148
rect 36876 2204 36940 2208
rect 36876 2148 36880 2204
rect 36880 2148 36936 2204
rect 36936 2148 36940 2204
rect 36876 2144 36940 2148
rect 36956 2204 37020 2208
rect 36956 2148 36960 2204
rect 36960 2148 37016 2204
rect 37016 2148 37020 2204
rect 36956 2144 37020 2148
rect 37036 2204 37100 2208
rect 37036 2148 37040 2204
rect 37040 2148 37096 2204
rect 37096 2148 37100 2204
rect 37036 2144 37100 2148
<< metal4 >>
rect 6918 27776 7238 27792
rect 6918 27712 6926 27776
rect 6990 27712 7006 27776
rect 7070 27712 7086 27776
rect 7150 27712 7166 27776
rect 7230 27712 7238 27776
rect 6918 26688 7238 27712
rect 6918 26624 6926 26688
rect 6990 26624 7006 26688
rect 7070 26624 7086 26688
rect 7150 26624 7166 26688
rect 7230 26624 7238 26688
rect 6918 25600 7238 26624
rect 6918 25536 6926 25600
rect 6990 25536 7006 25600
rect 7070 25536 7086 25600
rect 7150 25536 7166 25600
rect 7230 25536 7238 25600
rect 6918 24512 7238 25536
rect 6918 24448 6926 24512
rect 6990 24448 7006 24512
rect 7070 24448 7086 24512
rect 7150 24448 7166 24512
rect 7230 24448 7238 24512
rect 6918 23424 7238 24448
rect 6918 23360 6926 23424
rect 6990 23360 7006 23424
rect 7070 23360 7086 23424
rect 7150 23360 7166 23424
rect 7230 23360 7238 23424
rect 6918 22336 7238 23360
rect 6918 22272 6926 22336
rect 6990 22272 7006 22336
rect 7070 22272 7086 22336
rect 7150 22272 7166 22336
rect 7230 22272 7238 22336
rect 6918 21248 7238 22272
rect 6918 21184 6926 21248
rect 6990 21184 7006 21248
rect 7070 21184 7086 21248
rect 7150 21184 7166 21248
rect 7230 21184 7238 21248
rect 6918 20160 7238 21184
rect 6918 20096 6926 20160
rect 6990 20096 7006 20160
rect 7070 20096 7086 20160
rect 7150 20096 7166 20160
rect 7230 20096 7238 20160
rect 6918 19072 7238 20096
rect 6918 19008 6926 19072
rect 6990 19008 7006 19072
rect 7070 19008 7086 19072
rect 7150 19008 7166 19072
rect 7230 19008 7238 19072
rect 6918 17984 7238 19008
rect 6918 17920 6926 17984
rect 6990 17920 7006 17984
rect 7070 17920 7086 17984
rect 7150 17920 7166 17984
rect 7230 17920 7238 17984
rect 6918 16896 7238 17920
rect 6918 16832 6926 16896
rect 6990 16832 7006 16896
rect 7070 16832 7086 16896
rect 7150 16832 7166 16896
rect 7230 16832 7238 16896
rect 6918 15808 7238 16832
rect 6918 15744 6926 15808
rect 6990 15744 7006 15808
rect 7070 15744 7086 15808
rect 7150 15744 7166 15808
rect 7230 15744 7238 15808
rect 6918 14720 7238 15744
rect 6918 14656 6926 14720
rect 6990 14656 7006 14720
rect 7070 14656 7086 14720
rect 7150 14656 7166 14720
rect 7230 14656 7238 14720
rect 6918 13632 7238 14656
rect 6918 13568 6926 13632
rect 6990 13568 7006 13632
rect 7070 13568 7086 13632
rect 7150 13568 7166 13632
rect 7230 13568 7238 13632
rect 6918 12544 7238 13568
rect 6918 12480 6926 12544
rect 6990 12480 7006 12544
rect 7070 12480 7086 12544
rect 7150 12480 7166 12544
rect 7230 12480 7238 12544
rect 6918 11456 7238 12480
rect 6918 11392 6926 11456
rect 6990 11392 7006 11456
rect 7070 11392 7086 11456
rect 7150 11392 7166 11456
rect 7230 11392 7238 11456
rect 6918 10368 7238 11392
rect 6918 10304 6926 10368
rect 6990 10304 7006 10368
rect 7070 10304 7086 10368
rect 7150 10304 7166 10368
rect 7230 10304 7238 10368
rect 6918 9280 7238 10304
rect 6918 9216 6926 9280
rect 6990 9216 7006 9280
rect 7070 9216 7086 9280
rect 7150 9216 7166 9280
rect 7230 9216 7238 9280
rect 6918 8192 7238 9216
rect 6918 8128 6926 8192
rect 6990 8128 7006 8192
rect 7070 8128 7086 8192
rect 7150 8128 7166 8192
rect 7230 8128 7238 8192
rect 6918 7104 7238 8128
rect 6918 7040 6926 7104
rect 6990 7040 7006 7104
rect 7070 7040 7086 7104
rect 7150 7040 7166 7104
rect 7230 7040 7238 7104
rect 6918 6016 7238 7040
rect 6918 5952 6926 6016
rect 6990 5952 7006 6016
rect 7070 5952 7086 6016
rect 7150 5952 7166 6016
rect 7230 5952 7238 6016
rect 6918 4928 7238 5952
rect 6918 4864 6926 4928
rect 6990 4864 7006 4928
rect 7070 4864 7086 4928
rect 7150 4864 7166 4928
rect 7230 4864 7238 4928
rect 6918 3840 7238 4864
rect 6918 3776 6926 3840
rect 6990 3776 7006 3840
rect 7070 3776 7086 3840
rect 7150 3776 7166 3840
rect 7230 3776 7238 3840
rect 6918 2752 7238 3776
rect 6918 2688 6926 2752
rect 6990 2688 7006 2752
rect 7070 2688 7086 2752
rect 7150 2688 7166 2752
rect 7230 2688 7238 2752
rect 6918 2128 7238 2688
rect 12892 27232 13212 27792
rect 12892 27168 12900 27232
rect 12964 27168 12980 27232
rect 13044 27168 13060 27232
rect 13124 27168 13140 27232
rect 13204 27168 13212 27232
rect 12892 26144 13212 27168
rect 12892 26080 12900 26144
rect 12964 26080 12980 26144
rect 13044 26080 13060 26144
rect 13124 26080 13140 26144
rect 13204 26080 13212 26144
rect 12892 25056 13212 26080
rect 12892 24992 12900 25056
rect 12964 24992 12980 25056
rect 13044 24992 13060 25056
rect 13124 24992 13140 25056
rect 13204 24992 13212 25056
rect 12892 23968 13212 24992
rect 12892 23904 12900 23968
rect 12964 23904 12980 23968
rect 13044 23904 13060 23968
rect 13124 23904 13140 23968
rect 13204 23904 13212 23968
rect 12892 22880 13212 23904
rect 12892 22816 12900 22880
rect 12964 22816 12980 22880
rect 13044 22816 13060 22880
rect 13124 22816 13140 22880
rect 13204 22816 13212 22880
rect 12892 21792 13212 22816
rect 12892 21728 12900 21792
rect 12964 21728 12980 21792
rect 13044 21728 13060 21792
rect 13124 21728 13140 21792
rect 13204 21728 13212 21792
rect 12892 20704 13212 21728
rect 12892 20640 12900 20704
rect 12964 20640 12980 20704
rect 13044 20640 13060 20704
rect 13124 20640 13140 20704
rect 13204 20640 13212 20704
rect 12892 19616 13212 20640
rect 12892 19552 12900 19616
rect 12964 19552 12980 19616
rect 13044 19552 13060 19616
rect 13124 19552 13140 19616
rect 13204 19552 13212 19616
rect 12892 18528 13212 19552
rect 12892 18464 12900 18528
rect 12964 18464 12980 18528
rect 13044 18464 13060 18528
rect 13124 18464 13140 18528
rect 13204 18464 13212 18528
rect 12892 17440 13212 18464
rect 12892 17376 12900 17440
rect 12964 17376 12980 17440
rect 13044 17376 13060 17440
rect 13124 17376 13140 17440
rect 13204 17376 13212 17440
rect 12892 16352 13212 17376
rect 12892 16288 12900 16352
rect 12964 16288 12980 16352
rect 13044 16288 13060 16352
rect 13124 16288 13140 16352
rect 13204 16288 13212 16352
rect 12892 15264 13212 16288
rect 12892 15200 12900 15264
rect 12964 15200 12980 15264
rect 13044 15200 13060 15264
rect 13124 15200 13140 15264
rect 13204 15200 13212 15264
rect 12892 14176 13212 15200
rect 12892 14112 12900 14176
rect 12964 14112 12980 14176
rect 13044 14112 13060 14176
rect 13124 14112 13140 14176
rect 13204 14112 13212 14176
rect 12892 13088 13212 14112
rect 12892 13024 12900 13088
rect 12964 13024 12980 13088
rect 13044 13024 13060 13088
rect 13124 13024 13140 13088
rect 13204 13024 13212 13088
rect 12892 12000 13212 13024
rect 12892 11936 12900 12000
rect 12964 11936 12980 12000
rect 13044 11936 13060 12000
rect 13124 11936 13140 12000
rect 13204 11936 13212 12000
rect 12892 10912 13212 11936
rect 12892 10848 12900 10912
rect 12964 10848 12980 10912
rect 13044 10848 13060 10912
rect 13124 10848 13140 10912
rect 13204 10848 13212 10912
rect 12892 9824 13212 10848
rect 12892 9760 12900 9824
rect 12964 9760 12980 9824
rect 13044 9760 13060 9824
rect 13124 9760 13140 9824
rect 13204 9760 13212 9824
rect 12892 8736 13212 9760
rect 12892 8672 12900 8736
rect 12964 8672 12980 8736
rect 13044 8672 13060 8736
rect 13124 8672 13140 8736
rect 13204 8672 13212 8736
rect 12892 7648 13212 8672
rect 12892 7584 12900 7648
rect 12964 7584 12980 7648
rect 13044 7584 13060 7648
rect 13124 7584 13140 7648
rect 13204 7584 13212 7648
rect 12892 6560 13212 7584
rect 12892 6496 12900 6560
rect 12964 6496 12980 6560
rect 13044 6496 13060 6560
rect 13124 6496 13140 6560
rect 13204 6496 13212 6560
rect 12892 5472 13212 6496
rect 12892 5408 12900 5472
rect 12964 5408 12980 5472
rect 13044 5408 13060 5472
rect 13124 5408 13140 5472
rect 13204 5408 13212 5472
rect 12892 4384 13212 5408
rect 12892 4320 12900 4384
rect 12964 4320 12980 4384
rect 13044 4320 13060 4384
rect 13124 4320 13140 4384
rect 13204 4320 13212 4384
rect 12892 3296 13212 4320
rect 12892 3232 12900 3296
rect 12964 3232 12980 3296
rect 13044 3232 13060 3296
rect 13124 3232 13140 3296
rect 13204 3232 13212 3296
rect 12892 2208 13212 3232
rect 12892 2144 12900 2208
rect 12964 2144 12980 2208
rect 13044 2144 13060 2208
rect 13124 2144 13140 2208
rect 13204 2144 13212 2208
rect 12892 2128 13212 2144
rect 18866 27776 19186 27792
rect 18866 27712 18874 27776
rect 18938 27712 18954 27776
rect 19018 27712 19034 27776
rect 19098 27712 19114 27776
rect 19178 27712 19186 27776
rect 18866 26688 19186 27712
rect 18866 26624 18874 26688
rect 18938 26624 18954 26688
rect 19018 26624 19034 26688
rect 19098 26624 19114 26688
rect 19178 26624 19186 26688
rect 18866 25600 19186 26624
rect 18866 25536 18874 25600
rect 18938 25536 18954 25600
rect 19018 25536 19034 25600
rect 19098 25536 19114 25600
rect 19178 25536 19186 25600
rect 18866 24512 19186 25536
rect 18866 24448 18874 24512
rect 18938 24448 18954 24512
rect 19018 24448 19034 24512
rect 19098 24448 19114 24512
rect 19178 24448 19186 24512
rect 18866 23424 19186 24448
rect 18866 23360 18874 23424
rect 18938 23360 18954 23424
rect 19018 23360 19034 23424
rect 19098 23360 19114 23424
rect 19178 23360 19186 23424
rect 18866 22336 19186 23360
rect 18866 22272 18874 22336
rect 18938 22272 18954 22336
rect 19018 22272 19034 22336
rect 19098 22272 19114 22336
rect 19178 22272 19186 22336
rect 18866 21248 19186 22272
rect 18866 21184 18874 21248
rect 18938 21184 18954 21248
rect 19018 21184 19034 21248
rect 19098 21184 19114 21248
rect 19178 21184 19186 21248
rect 18866 20160 19186 21184
rect 18866 20096 18874 20160
rect 18938 20096 18954 20160
rect 19018 20096 19034 20160
rect 19098 20096 19114 20160
rect 19178 20096 19186 20160
rect 18866 19072 19186 20096
rect 18866 19008 18874 19072
rect 18938 19008 18954 19072
rect 19018 19008 19034 19072
rect 19098 19008 19114 19072
rect 19178 19008 19186 19072
rect 18866 17984 19186 19008
rect 18866 17920 18874 17984
rect 18938 17920 18954 17984
rect 19018 17920 19034 17984
rect 19098 17920 19114 17984
rect 19178 17920 19186 17984
rect 18866 16896 19186 17920
rect 18866 16832 18874 16896
rect 18938 16832 18954 16896
rect 19018 16832 19034 16896
rect 19098 16832 19114 16896
rect 19178 16832 19186 16896
rect 18866 15808 19186 16832
rect 18866 15744 18874 15808
rect 18938 15744 18954 15808
rect 19018 15744 19034 15808
rect 19098 15744 19114 15808
rect 19178 15744 19186 15808
rect 18866 14720 19186 15744
rect 18866 14656 18874 14720
rect 18938 14656 18954 14720
rect 19018 14656 19034 14720
rect 19098 14656 19114 14720
rect 19178 14656 19186 14720
rect 18866 13632 19186 14656
rect 18866 13568 18874 13632
rect 18938 13568 18954 13632
rect 19018 13568 19034 13632
rect 19098 13568 19114 13632
rect 19178 13568 19186 13632
rect 18866 12544 19186 13568
rect 18866 12480 18874 12544
rect 18938 12480 18954 12544
rect 19018 12480 19034 12544
rect 19098 12480 19114 12544
rect 19178 12480 19186 12544
rect 18866 11456 19186 12480
rect 18866 11392 18874 11456
rect 18938 11392 18954 11456
rect 19018 11392 19034 11456
rect 19098 11392 19114 11456
rect 19178 11392 19186 11456
rect 18866 10368 19186 11392
rect 18866 10304 18874 10368
rect 18938 10304 18954 10368
rect 19018 10304 19034 10368
rect 19098 10304 19114 10368
rect 19178 10304 19186 10368
rect 18866 9280 19186 10304
rect 18866 9216 18874 9280
rect 18938 9216 18954 9280
rect 19018 9216 19034 9280
rect 19098 9216 19114 9280
rect 19178 9216 19186 9280
rect 18866 8192 19186 9216
rect 18866 8128 18874 8192
rect 18938 8128 18954 8192
rect 19018 8128 19034 8192
rect 19098 8128 19114 8192
rect 19178 8128 19186 8192
rect 18866 7104 19186 8128
rect 18866 7040 18874 7104
rect 18938 7040 18954 7104
rect 19018 7040 19034 7104
rect 19098 7040 19114 7104
rect 19178 7040 19186 7104
rect 18866 6016 19186 7040
rect 18866 5952 18874 6016
rect 18938 5952 18954 6016
rect 19018 5952 19034 6016
rect 19098 5952 19114 6016
rect 19178 5952 19186 6016
rect 18866 4928 19186 5952
rect 18866 4864 18874 4928
rect 18938 4864 18954 4928
rect 19018 4864 19034 4928
rect 19098 4864 19114 4928
rect 19178 4864 19186 4928
rect 18866 3840 19186 4864
rect 18866 3776 18874 3840
rect 18938 3776 18954 3840
rect 19018 3776 19034 3840
rect 19098 3776 19114 3840
rect 19178 3776 19186 3840
rect 18866 2752 19186 3776
rect 18866 2688 18874 2752
rect 18938 2688 18954 2752
rect 19018 2688 19034 2752
rect 19098 2688 19114 2752
rect 19178 2688 19186 2752
rect 18866 2128 19186 2688
rect 24840 27232 25160 27792
rect 24840 27168 24848 27232
rect 24912 27168 24928 27232
rect 24992 27168 25008 27232
rect 25072 27168 25088 27232
rect 25152 27168 25160 27232
rect 24840 26144 25160 27168
rect 24840 26080 24848 26144
rect 24912 26080 24928 26144
rect 24992 26080 25008 26144
rect 25072 26080 25088 26144
rect 25152 26080 25160 26144
rect 24840 25056 25160 26080
rect 24840 24992 24848 25056
rect 24912 24992 24928 25056
rect 24992 24992 25008 25056
rect 25072 24992 25088 25056
rect 25152 24992 25160 25056
rect 24840 23968 25160 24992
rect 24840 23904 24848 23968
rect 24912 23904 24928 23968
rect 24992 23904 25008 23968
rect 25072 23904 25088 23968
rect 25152 23904 25160 23968
rect 24840 22880 25160 23904
rect 24840 22816 24848 22880
rect 24912 22816 24928 22880
rect 24992 22816 25008 22880
rect 25072 22816 25088 22880
rect 25152 22816 25160 22880
rect 24840 21792 25160 22816
rect 24840 21728 24848 21792
rect 24912 21728 24928 21792
rect 24992 21728 25008 21792
rect 25072 21728 25088 21792
rect 25152 21728 25160 21792
rect 24840 20704 25160 21728
rect 24840 20640 24848 20704
rect 24912 20640 24928 20704
rect 24992 20640 25008 20704
rect 25072 20640 25088 20704
rect 25152 20640 25160 20704
rect 24840 19616 25160 20640
rect 24840 19552 24848 19616
rect 24912 19552 24928 19616
rect 24992 19552 25008 19616
rect 25072 19552 25088 19616
rect 25152 19552 25160 19616
rect 24840 18528 25160 19552
rect 24840 18464 24848 18528
rect 24912 18464 24928 18528
rect 24992 18464 25008 18528
rect 25072 18464 25088 18528
rect 25152 18464 25160 18528
rect 24840 17440 25160 18464
rect 24840 17376 24848 17440
rect 24912 17376 24928 17440
rect 24992 17376 25008 17440
rect 25072 17376 25088 17440
rect 25152 17376 25160 17440
rect 24840 16352 25160 17376
rect 24840 16288 24848 16352
rect 24912 16288 24928 16352
rect 24992 16288 25008 16352
rect 25072 16288 25088 16352
rect 25152 16288 25160 16352
rect 24840 15264 25160 16288
rect 24840 15200 24848 15264
rect 24912 15200 24928 15264
rect 24992 15200 25008 15264
rect 25072 15200 25088 15264
rect 25152 15200 25160 15264
rect 24840 14176 25160 15200
rect 24840 14112 24848 14176
rect 24912 14112 24928 14176
rect 24992 14112 25008 14176
rect 25072 14112 25088 14176
rect 25152 14112 25160 14176
rect 24840 13088 25160 14112
rect 24840 13024 24848 13088
rect 24912 13024 24928 13088
rect 24992 13024 25008 13088
rect 25072 13024 25088 13088
rect 25152 13024 25160 13088
rect 24840 12000 25160 13024
rect 24840 11936 24848 12000
rect 24912 11936 24928 12000
rect 24992 11936 25008 12000
rect 25072 11936 25088 12000
rect 25152 11936 25160 12000
rect 24840 10912 25160 11936
rect 24840 10848 24848 10912
rect 24912 10848 24928 10912
rect 24992 10848 25008 10912
rect 25072 10848 25088 10912
rect 25152 10848 25160 10912
rect 24840 9824 25160 10848
rect 24840 9760 24848 9824
rect 24912 9760 24928 9824
rect 24992 9760 25008 9824
rect 25072 9760 25088 9824
rect 25152 9760 25160 9824
rect 24840 8736 25160 9760
rect 24840 8672 24848 8736
rect 24912 8672 24928 8736
rect 24992 8672 25008 8736
rect 25072 8672 25088 8736
rect 25152 8672 25160 8736
rect 24840 7648 25160 8672
rect 24840 7584 24848 7648
rect 24912 7584 24928 7648
rect 24992 7584 25008 7648
rect 25072 7584 25088 7648
rect 25152 7584 25160 7648
rect 24840 6560 25160 7584
rect 24840 6496 24848 6560
rect 24912 6496 24928 6560
rect 24992 6496 25008 6560
rect 25072 6496 25088 6560
rect 25152 6496 25160 6560
rect 24840 5472 25160 6496
rect 24840 5408 24848 5472
rect 24912 5408 24928 5472
rect 24992 5408 25008 5472
rect 25072 5408 25088 5472
rect 25152 5408 25160 5472
rect 24840 4384 25160 5408
rect 24840 4320 24848 4384
rect 24912 4320 24928 4384
rect 24992 4320 25008 4384
rect 25072 4320 25088 4384
rect 25152 4320 25160 4384
rect 24840 3296 25160 4320
rect 24840 3232 24848 3296
rect 24912 3232 24928 3296
rect 24992 3232 25008 3296
rect 25072 3232 25088 3296
rect 25152 3232 25160 3296
rect 24840 2208 25160 3232
rect 24840 2144 24848 2208
rect 24912 2144 24928 2208
rect 24992 2144 25008 2208
rect 25072 2144 25088 2208
rect 25152 2144 25160 2208
rect 24840 2128 25160 2144
rect 30814 27776 31134 27792
rect 30814 27712 30822 27776
rect 30886 27712 30902 27776
rect 30966 27712 30982 27776
rect 31046 27712 31062 27776
rect 31126 27712 31134 27776
rect 30814 26688 31134 27712
rect 30814 26624 30822 26688
rect 30886 26624 30902 26688
rect 30966 26624 30982 26688
rect 31046 26624 31062 26688
rect 31126 26624 31134 26688
rect 30814 25600 31134 26624
rect 30814 25536 30822 25600
rect 30886 25536 30902 25600
rect 30966 25536 30982 25600
rect 31046 25536 31062 25600
rect 31126 25536 31134 25600
rect 30814 24512 31134 25536
rect 30814 24448 30822 24512
rect 30886 24448 30902 24512
rect 30966 24448 30982 24512
rect 31046 24448 31062 24512
rect 31126 24448 31134 24512
rect 30814 23424 31134 24448
rect 30814 23360 30822 23424
rect 30886 23360 30902 23424
rect 30966 23360 30982 23424
rect 31046 23360 31062 23424
rect 31126 23360 31134 23424
rect 30814 22336 31134 23360
rect 30814 22272 30822 22336
rect 30886 22272 30902 22336
rect 30966 22272 30982 22336
rect 31046 22272 31062 22336
rect 31126 22272 31134 22336
rect 30814 21248 31134 22272
rect 30814 21184 30822 21248
rect 30886 21184 30902 21248
rect 30966 21184 30982 21248
rect 31046 21184 31062 21248
rect 31126 21184 31134 21248
rect 30814 20160 31134 21184
rect 30814 20096 30822 20160
rect 30886 20096 30902 20160
rect 30966 20096 30982 20160
rect 31046 20096 31062 20160
rect 31126 20096 31134 20160
rect 30814 19072 31134 20096
rect 30814 19008 30822 19072
rect 30886 19008 30902 19072
rect 30966 19008 30982 19072
rect 31046 19008 31062 19072
rect 31126 19008 31134 19072
rect 30814 17984 31134 19008
rect 30814 17920 30822 17984
rect 30886 17920 30902 17984
rect 30966 17920 30982 17984
rect 31046 17920 31062 17984
rect 31126 17920 31134 17984
rect 30814 16896 31134 17920
rect 30814 16832 30822 16896
rect 30886 16832 30902 16896
rect 30966 16832 30982 16896
rect 31046 16832 31062 16896
rect 31126 16832 31134 16896
rect 30814 15808 31134 16832
rect 30814 15744 30822 15808
rect 30886 15744 30902 15808
rect 30966 15744 30982 15808
rect 31046 15744 31062 15808
rect 31126 15744 31134 15808
rect 30814 14720 31134 15744
rect 30814 14656 30822 14720
rect 30886 14656 30902 14720
rect 30966 14656 30982 14720
rect 31046 14656 31062 14720
rect 31126 14656 31134 14720
rect 30814 13632 31134 14656
rect 30814 13568 30822 13632
rect 30886 13568 30902 13632
rect 30966 13568 30982 13632
rect 31046 13568 31062 13632
rect 31126 13568 31134 13632
rect 30814 12544 31134 13568
rect 30814 12480 30822 12544
rect 30886 12480 30902 12544
rect 30966 12480 30982 12544
rect 31046 12480 31062 12544
rect 31126 12480 31134 12544
rect 30814 11456 31134 12480
rect 30814 11392 30822 11456
rect 30886 11392 30902 11456
rect 30966 11392 30982 11456
rect 31046 11392 31062 11456
rect 31126 11392 31134 11456
rect 30814 10368 31134 11392
rect 30814 10304 30822 10368
rect 30886 10304 30902 10368
rect 30966 10304 30982 10368
rect 31046 10304 31062 10368
rect 31126 10304 31134 10368
rect 30814 9280 31134 10304
rect 30814 9216 30822 9280
rect 30886 9216 30902 9280
rect 30966 9216 30982 9280
rect 31046 9216 31062 9280
rect 31126 9216 31134 9280
rect 30814 8192 31134 9216
rect 30814 8128 30822 8192
rect 30886 8128 30902 8192
rect 30966 8128 30982 8192
rect 31046 8128 31062 8192
rect 31126 8128 31134 8192
rect 30814 7104 31134 8128
rect 30814 7040 30822 7104
rect 30886 7040 30902 7104
rect 30966 7040 30982 7104
rect 31046 7040 31062 7104
rect 31126 7040 31134 7104
rect 30814 6016 31134 7040
rect 30814 5952 30822 6016
rect 30886 5952 30902 6016
rect 30966 5952 30982 6016
rect 31046 5952 31062 6016
rect 31126 5952 31134 6016
rect 30814 4928 31134 5952
rect 30814 4864 30822 4928
rect 30886 4864 30902 4928
rect 30966 4864 30982 4928
rect 31046 4864 31062 4928
rect 31126 4864 31134 4928
rect 30814 3840 31134 4864
rect 30814 3776 30822 3840
rect 30886 3776 30902 3840
rect 30966 3776 30982 3840
rect 31046 3776 31062 3840
rect 31126 3776 31134 3840
rect 30814 2752 31134 3776
rect 30814 2688 30822 2752
rect 30886 2688 30902 2752
rect 30966 2688 30982 2752
rect 31046 2688 31062 2752
rect 31126 2688 31134 2752
rect 30814 2128 31134 2688
rect 36788 27232 37108 27792
rect 36788 27168 36796 27232
rect 36860 27168 36876 27232
rect 36940 27168 36956 27232
rect 37020 27168 37036 27232
rect 37100 27168 37108 27232
rect 36788 26144 37108 27168
rect 36788 26080 36796 26144
rect 36860 26080 36876 26144
rect 36940 26080 36956 26144
rect 37020 26080 37036 26144
rect 37100 26080 37108 26144
rect 36788 25056 37108 26080
rect 36788 24992 36796 25056
rect 36860 24992 36876 25056
rect 36940 24992 36956 25056
rect 37020 24992 37036 25056
rect 37100 24992 37108 25056
rect 36788 23968 37108 24992
rect 36788 23904 36796 23968
rect 36860 23904 36876 23968
rect 36940 23904 36956 23968
rect 37020 23904 37036 23968
rect 37100 23904 37108 23968
rect 36788 22880 37108 23904
rect 36788 22816 36796 22880
rect 36860 22816 36876 22880
rect 36940 22816 36956 22880
rect 37020 22816 37036 22880
rect 37100 22816 37108 22880
rect 36788 21792 37108 22816
rect 36788 21728 36796 21792
rect 36860 21728 36876 21792
rect 36940 21728 36956 21792
rect 37020 21728 37036 21792
rect 37100 21728 37108 21792
rect 36788 20704 37108 21728
rect 36788 20640 36796 20704
rect 36860 20640 36876 20704
rect 36940 20640 36956 20704
rect 37020 20640 37036 20704
rect 37100 20640 37108 20704
rect 36788 19616 37108 20640
rect 36788 19552 36796 19616
rect 36860 19552 36876 19616
rect 36940 19552 36956 19616
rect 37020 19552 37036 19616
rect 37100 19552 37108 19616
rect 36788 18528 37108 19552
rect 36788 18464 36796 18528
rect 36860 18464 36876 18528
rect 36940 18464 36956 18528
rect 37020 18464 37036 18528
rect 37100 18464 37108 18528
rect 36788 17440 37108 18464
rect 36788 17376 36796 17440
rect 36860 17376 36876 17440
rect 36940 17376 36956 17440
rect 37020 17376 37036 17440
rect 37100 17376 37108 17440
rect 36788 16352 37108 17376
rect 36788 16288 36796 16352
rect 36860 16288 36876 16352
rect 36940 16288 36956 16352
rect 37020 16288 37036 16352
rect 37100 16288 37108 16352
rect 36788 15264 37108 16288
rect 36788 15200 36796 15264
rect 36860 15200 36876 15264
rect 36940 15200 36956 15264
rect 37020 15200 37036 15264
rect 37100 15200 37108 15264
rect 36788 14176 37108 15200
rect 36788 14112 36796 14176
rect 36860 14112 36876 14176
rect 36940 14112 36956 14176
rect 37020 14112 37036 14176
rect 37100 14112 37108 14176
rect 36788 13088 37108 14112
rect 36788 13024 36796 13088
rect 36860 13024 36876 13088
rect 36940 13024 36956 13088
rect 37020 13024 37036 13088
rect 37100 13024 37108 13088
rect 36788 12000 37108 13024
rect 36788 11936 36796 12000
rect 36860 11936 36876 12000
rect 36940 11936 36956 12000
rect 37020 11936 37036 12000
rect 37100 11936 37108 12000
rect 36788 10912 37108 11936
rect 36788 10848 36796 10912
rect 36860 10848 36876 10912
rect 36940 10848 36956 10912
rect 37020 10848 37036 10912
rect 37100 10848 37108 10912
rect 36788 9824 37108 10848
rect 36788 9760 36796 9824
rect 36860 9760 36876 9824
rect 36940 9760 36956 9824
rect 37020 9760 37036 9824
rect 37100 9760 37108 9824
rect 36788 8736 37108 9760
rect 36788 8672 36796 8736
rect 36860 8672 36876 8736
rect 36940 8672 36956 8736
rect 37020 8672 37036 8736
rect 37100 8672 37108 8736
rect 36788 7648 37108 8672
rect 36788 7584 36796 7648
rect 36860 7584 36876 7648
rect 36940 7584 36956 7648
rect 37020 7584 37036 7648
rect 37100 7584 37108 7648
rect 36788 6560 37108 7584
rect 36788 6496 36796 6560
rect 36860 6496 36876 6560
rect 36940 6496 36956 6560
rect 37020 6496 37036 6560
rect 37100 6496 37108 6560
rect 36788 5472 37108 6496
rect 36788 5408 36796 5472
rect 36860 5408 36876 5472
rect 36940 5408 36956 5472
rect 37020 5408 37036 5472
rect 37100 5408 37108 5472
rect 36788 4384 37108 5408
rect 36788 4320 36796 4384
rect 36860 4320 36876 4384
rect 36940 4320 36956 4384
rect 37020 4320 37036 4384
rect 37100 4320 37108 4384
rect 36788 3296 37108 4320
rect 36788 3232 36796 3296
rect 36860 3232 36876 3296
rect 36940 3232 36956 3296
rect 37020 3232 37036 3296
rect 37100 3232 37108 3296
rect 36788 2208 37108 3232
rect 36788 2144 36796 2208
rect 36860 2144 36876 2208
rect 36940 2144 36956 2208
rect 37020 2144 37036 2208
rect 37100 2144 37108 2208
rect 36788 2128 37108 2144
rect 42762 27776 43082 27792
rect 42762 27712 42770 27776
rect 42834 27712 42850 27776
rect 42914 27712 42930 27776
rect 42994 27712 43010 27776
rect 43074 27712 43082 27776
rect 42762 26688 43082 27712
rect 42762 26624 42770 26688
rect 42834 26624 42850 26688
rect 42914 26624 42930 26688
rect 42994 26624 43010 26688
rect 43074 26624 43082 26688
rect 42762 25600 43082 26624
rect 42762 25536 42770 25600
rect 42834 25536 42850 25600
rect 42914 25536 42930 25600
rect 42994 25536 43010 25600
rect 43074 25536 43082 25600
rect 42762 24512 43082 25536
rect 42762 24448 42770 24512
rect 42834 24448 42850 24512
rect 42914 24448 42930 24512
rect 42994 24448 43010 24512
rect 43074 24448 43082 24512
rect 42762 23424 43082 24448
rect 42762 23360 42770 23424
rect 42834 23360 42850 23424
rect 42914 23360 42930 23424
rect 42994 23360 43010 23424
rect 43074 23360 43082 23424
rect 42762 22336 43082 23360
rect 42762 22272 42770 22336
rect 42834 22272 42850 22336
rect 42914 22272 42930 22336
rect 42994 22272 43010 22336
rect 43074 22272 43082 22336
rect 42762 21248 43082 22272
rect 42762 21184 42770 21248
rect 42834 21184 42850 21248
rect 42914 21184 42930 21248
rect 42994 21184 43010 21248
rect 43074 21184 43082 21248
rect 42762 20160 43082 21184
rect 42762 20096 42770 20160
rect 42834 20096 42850 20160
rect 42914 20096 42930 20160
rect 42994 20096 43010 20160
rect 43074 20096 43082 20160
rect 42762 19072 43082 20096
rect 42762 19008 42770 19072
rect 42834 19008 42850 19072
rect 42914 19008 42930 19072
rect 42994 19008 43010 19072
rect 43074 19008 43082 19072
rect 42762 17984 43082 19008
rect 42762 17920 42770 17984
rect 42834 17920 42850 17984
rect 42914 17920 42930 17984
rect 42994 17920 43010 17984
rect 43074 17920 43082 17984
rect 42762 16896 43082 17920
rect 42762 16832 42770 16896
rect 42834 16832 42850 16896
rect 42914 16832 42930 16896
rect 42994 16832 43010 16896
rect 43074 16832 43082 16896
rect 42762 15808 43082 16832
rect 42762 15744 42770 15808
rect 42834 15744 42850 15808
rect 42914 15744 42930 15808
rect 42994 15744 43010 15808
rect 43074 15744 43082 15808
rect 42762 14720 43082 15744
rect 42762 14656 42770 14720
rect 42834 14656 42850 14720
rect 42914 14656 42930 14720
rect 42994 14656 43010 14720
rect 43074 14656 43082 14720
rect 42762 13632 43082 14656
rect 42762 13568 42770 13632
rect 42834 13568 42850 13632
rect 42914 13568 42930 13632
rect 42994 13568 43010 13632
rect 43074 13568 43082 13632
rect 42762 12544 43082 13568
rect 42762 12480 42770 12544
rect 42834 12480 42850 12544
rect 42914 12480 42930 12544
rect 42994 12480 43010 12544
rect 43074 12480 43082 12544
rect 42762 11456 43082 12480
rect 42762 11392 42770 11456
rect 42834 11392 42850 11456
rect 42914 11392 42930 11456
rect 42994 11392 43010 11456
rect 43074 11392 43082 11456
rect 42762 10368 43082 11392
rect 42762 10304 42770 10368
rect 42834 10304 42850 10368
rect 42914 10304 42930 10368
rect 42994 10304 43010 10368
rect 43074 10304 43082 10368
rect 42762 9280 43082 10304
rect 42762 9216 42770 9280
rect 42834 9216 42850 9280
rect 42914 9216 42930 9280
rect 42994 9216 43010 9280
rect 43074 9216 43082 9280
rect 42762 8192 43082 9216
rect 42762 8128 42770 8192
rect 42834 8128 42850 8192
rect 42914 8128 42930 8192
rect 42994 8128 43010 8192
rect 43074 8128 43082 8192
rect 42762 7104 43082 8128
rect 42762 7040 42770 7104
rect 42834 7040 42850 7104
rect 42914 7040 42930 7104
rect 42994 7040 43010 7104
rect 43074 7040 43082 7104
rect 42762 6016 43082 7040
rect 42762 5952 42770 6016
rect 42834 5952 42850 6016
rect 42914 5952 42930 6016
rect 42994 5952 43010 6016
rect 43074 5952 43082 6016
rect 42762 4928 43082 5952
rect 42762 4864 42770 4928
rect 42834 4864 42850 4928
rect 42914 4864 42930 4928
rect 42994 4864 43010 4928
rect 43074 4864 43082 4928
rect 42762 3840 43082 4864
rect 42762 3776 42770 3840
rect 42834 3776 42850 3840
rect 42914 3776 42930 3840
rect 42994 3776 43010 3840
rect 43074 3776 43082 3840
rect 42762 2752 43082 3776
rect 42762 2688 42770 2752
rect 42834 2688 42850 2752
rect 42914 2688 42930 2752
rect 42994 2688 43010 2752
rect 43074 2688 43082 2752
rect 42762 2128 43082 2688
use sky130_fd_sc_hd__decap_8  FILLER_0_6 ../openroad/OpenLane/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1659098407
transform 1 0 1656 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17 ../openroad/OpenLane/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1659098407
transform 1 0 2668 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24
timestamp 1659098407
transform 1 0 3312 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29 ../openroad/OpenLane/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1659098407
transform 1 0 3772 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38
timestamp 1659098407
transform 1 0 4600 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_45
timestamp 1659098407
transform 1 0 5244 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_52
timestamp 1659098407
transform 1 0 5888 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_57
timestamp 1659098407
transform 1 0 6348 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_66
timestamp 1659098407
transform 1 0 7176 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_73
timestamp 1659098407
transform 1 0 7820 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_80
timestamp 1659098407
transform 1 0 8464 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_85
timestamp 1659098407
transform 1 0 8924 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_94
timestamp 1659098407
transform 1 0 9752 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_101
timestamp 1659098407
transform 1 0 10396 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_108
timestamp 1659098407
transform 1 0 11040 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_113 ../openroad/OpenLane/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1659098407
transform 1 0 11500 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_118
timestamp 1659098407
transform 1 0 11960 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_125
timestamp 1659098407
transform 1 0 12604 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_132
timestamp 1659098407
transform 1 0 13248 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_144
timestamp 1659098407
transform 1 0 14352 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_153
timestamp 1659098407
transform 1 0 15180 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_164
timestamp 1659098407
transform 1 0 16192 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_169
timestamp 1659098407
transform 1 0 16652 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_178
timestamp 1659098407
transform 1 0 17480 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_185
timestamp 1659098407
transform 1 0 18124 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_192
timestamp 1659098407
transform 1 0 18768 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_197
timestamp 1659098407
transform 1 0 19228 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_206
timestamp 1659098407
transform 1 0 20056 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_213
timestamp 1659098407
transform 1 0 20700 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_220
timestamp 1659098407
transform 1 0 21344 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_225
timestamp 1659098407
transform 1 0 21804 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_230
timestamp 1659098407
transform 1 0 22264 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_238
timestamp 1659098407
transform 1 0 23000 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_244 ../openroad/OpenLane/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1659098407
transform 1 0 23552 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_248
timestamp 1659098407
transform 1 0 23920 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_253
timestamp 1659098407
transform 1 0 24380 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_258
timestamp 1659098407
transform 1 0 24840 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_265
timestamp 1659098407
transform 1 0 25484 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_272
timestamp 1659098407
transform 1 0 26128 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_284
timestamp 1659098407
transform 1 0 27232 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_291
timestamp 1659098407
transform 1 0 27876 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_298
timestamp 1659098407
transform 1 0 28520 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_306
timestamp 1659098407
transform 1 0 29256 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_312
timestamp 1659098407
transform 1 0 29808 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_319
timestamp 1659098407
transform 1 0 30452 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_326
timestamp 1659098407
transform 1 0 31096 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_334
timestamp 1659098407
transform 1 0 31832 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_337
timestamp 1659098407
transform 1 0 32108 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_342
timestamp 1659098407
transform 1 0 32568 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_349
timestamp 1659098407
transform 1 0 33212 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_356
timestamp 1659098407
transform 1 0 33856 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_368
timestamp 1659098407
transform 1 0 34960 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_375
timestamp 1659098407
transform 1 0 35604 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_382
timestamp 1659098407
transform 1 0 36248 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_390
timestamp 1659098407
transform 1 0 36984 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_393
timestamp 1659098407
transform 1 0 37260 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_398
timestamp 1659098407
transform 1 0 37720 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_406 ../openroad/OpenLane/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1659098407
transform 1 0 38456 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_412
timestamp 1659098407
transform 1 0 39008 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_424
timestamp 1659098407
transform 1 0 40112 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_433
timestamp 1659098407
transform 1 0 40940 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_440
timestamp 1659098407
transform 1 0 41584 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_452
timestamp 1659098407
transform 1 0 42688 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_459
timestamp 1659098407
transform 1 0 43332 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_466
timestamp 1659098407
transform 1 0 43976 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_474
timestamp 1659098407
transform 1 0 44712 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_480
timestamp 1659098407
transform 1 0 45264 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_487
timestamp 1659098407
transform 1 0 45908 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_496
timestamp 1659098407
transform 1 0 46736 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_508
timestamp 1659098407
transform 1 0 47840 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_1_6
timestamp 1659098407
transform 1 0 1656 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_13
timestamp 1659098407
transform 1 0 2300 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_20
timestamp 1659098407
transform 1 0 2944 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_1_28
timestamp 1659098407
transform 1 0 3680 0 -1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_1_34 ../openroad/OpenLane/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1659098407
transform 1 0 4232 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_46
timestamp 1659098407
transform 1 0 5336 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_54
timestamp 1659098407
transform 1 0 6072 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_1_57
timestamp 1659098407
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_69
timestamp 1659098407
transform 1 0 7452 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_81
timestamp 1659098407
transform 1 0 8556 0 -1 3264
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_1_90
timestamp 1659098407
transform 1 0 9384 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_102
timestamp 1659098407
transform 1 0 10488 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_110
timestamp 1659098407
transform 1 0 11224 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_1_113
timestamp 1659098407
transform 1 0 11500 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_125
timestamp 1659098407
transform 1 0 12604 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_137
timestamp 1659098407
transform 1 0 13708 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_149
timestamp 1659098407
transform 1 0 14812 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_161
timestamp 1659098407
transform 1 0 15916 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_167
timestamp 1659098407
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_169
timestamp 1659098407
transform 1 0 16652 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_1_174
timestamp 1659098407
transform 1 0 17112 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_186
timestamp 1659098407
transform 1 0 18216 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_198
timestamp 1659098407
transform 1 0 19320 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_202
timestamp 1659098407
transform 1 0 19688 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_214
timestamp 1659098407
transform 1 0 20792 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_222
timestamp 1659098407
transform 1 0 21528 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_1_225
timestamp 1659098407
transform 1 0 21804 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_237
timestamp 1659098407
transform 1 0 22908 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_244
timestamp 1659098407
transform 1 0 23552 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_256
timestamp 1659098407
transform 1 0 24656 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_268
timestamp 1659098407
transform 1 0 25760 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_281
timestamp 1659098407
transform 1 0 26956 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_293
timestamp 1659098407
transform 1 0 28060 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_300
timestamp 1659098407
transform 1 0 28704 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_312
timestamp 1659098407
transform 1 0 29808 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_324
timestamp 1659098407
transform 1 0 30912 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_328
timestamp 1659098407
transform 1 0 31280 0 -1 3264
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_1_337
timestamp 1659098407
transform 1 0 32108 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_349
timestamp 1659098407
transform 1 0 33212 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_361
timestamp 1659098407
transform 1 0 34316 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_373
timestamp 1659098407
transform 1 0 35420 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_1_384
timestamp 1659098407
transform 1 0 36432 0 -1 3264
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_1_393
timestamp 1659098407
transform 1 0 37260 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_405
timestamp 1659098407
transform 1 0 38364 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_417
timestamp 1659098407
transform 1 0 39468 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_429
timestamp 1659098407
transform 1 0 40572 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_441
timestamp 1659098407
transform 1 0 41676 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_447
timestamp 1659098407
transform 1 0 42228 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_449
timestamp 1659098407
transform 1 0 42412 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_461
timestamp 1659098407
transform 1 0 43516 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_468
timestamp 1659098407
transform 1 0 44160 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_1_480
timestamp 1659098407
transform 1 0 45264 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_486
timestamp 1659098407
transform 1 0 45816 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_493
timestamp 1659098407
transform 1 0 46460 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_500
timestamp 1659098407
transform 1 0 47104 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_505
timestamp 1659098407
transform 1 0 47564 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_1_510
timestamp 1659098407
transform 1 0 48024 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_2_6
timestamp 1659098407
transform 1 0 1656 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_13
timestamp 1659098407
transform 1 0 2300 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_20
timestamp 1659098407
transform 1 0 2944 0 1 3264
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_2_29
timestamp 1659098407
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_41
timestamp 1659098407
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_53
timestamp 1659098407
transform 1 0 5980 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_65
timestamp 1659098407
transform 1 0 7084 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_77
timestamp 1659098407
transform 1 0 8188 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_83
timestamp 1659098407
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_85
timestamp 1659098407
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_97
timestamp 1659098407
transform 1 0 10028 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_109
timestamp 1659098407
transform 1 0 11132 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_121
timestamp 1659098407
transform 1 0 12236 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_133
timestamp 1659098407
transform 1 0 13340 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_139
timestamp 1659098407
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_141
timestamp 1659098407
transform 1 0 14076 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_153
timestamp 1659098407
transform 1 0 15180 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_165
timestamp 1659098407
transform 1 0 16284 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_177
timestamp 1659098407
transform 1 0 17388 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_189
timestamp 1659098407
transform 1 0 18492 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_195
timestamp 1659098407
transform 1 0 19044 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_197
timestamp 1659098407
transform 1 0 19228 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_209
timestamp 1659098407
transform 1 0 20332 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_221
timestamp 1659098407
transform 1 0 21436 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_233
timestamp 1659098407
transform 1 0 22540 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_245
timestamp 1659098407
transform 1 0 23644 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_251
timestamp 1659098407
transform 1 0 24196 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_253
timestamp 1659098407
transform 1 0 24380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_265
timestamp 1659098407
transform 1 0 25484 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_277
timestamp 1659098407
transform 1 0 26588 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_289
timestamp 1659098407
transform 1 0 27692 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_301
timestamp 1659098407
transform 1 0 28796 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_307
timestamp 1659098407
transform 1 0 29348 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_309
timestamp 1659098407
transform 1 0 29532 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_321
timestamp 1659098407
transform 1 0 30636 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_333
timestamp 1659098407
transform 1 0 31740 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_345
timestamp 1659098407
transform 1 0 32844 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_357
timestamp 1659098407
transform 1 0 33948 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_363
timestamp 1659098407
transform 1 0 34500 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_365
timestamp 1659098407
transform 1 0 34684 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_377
timestamp 1659098407
transform 1 0 35788 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_389
timestamp 1659098407
transform 1 0 36892 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_401
timestamp 1659098407
transform 1 0 37996 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_413
timestamp 1659098407
transform 1 0 39100 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_419
timestamp 1659098407
transform 1 0 39652 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_421
timestamp 1659098407
transform 1 0 39836 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_433
timestamp 1659098407
transform 1 0 40940 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_445
timestamp 1659098407
transform 1 0 42044 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_457
timestamp 1659098407
transform 1 0 43148 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_469
timestamp 1659098407
transform 1 0 44252 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_475
timestamp 1659098407
transform 1 0 44804 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_477
timestamp 1659098407
transform 1 0 44988 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_489
timestamp 1659098407
transform 1 0 46092 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_2_498
timestamp 1659098407
transform 1 0 46920 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_505
timestamp 1659098407
transform 1 0 47564 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_512
timestamp 1659098407
transform 1 0 48208 0 1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_3_6
timestamp 1659098407
transform 1 0 1656 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_18
timestamp 1659098407
transform 1 0 2760 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_30
timestamp 1659098407
transform 1 0 3864 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_42
timestamp 1659098407
transform 1 0 4968 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_3_54
timestamp 1659098407
transform 1 0 6072 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_3_57
timestamp 1659098407
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_69
timestamp 1659098407
transform 1 0 7452 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_81
timestamp 1659098407
transform 1 0 8556 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_93
timestamp 1659098407
transform 1 0 9660 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_105
timestamp 1659098407
transform 1 0 10764 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_111
timestamp 1659098407
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_113
timestamp 1659098407
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_125
timestamp 1659098407
transform 1 0 12604 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_137
timestamp 1659098407
transform 1 0 13708 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_149
timestamp 1659098407
transform 1 0 14812 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_161
timestamp 1659098407
transform 1 0 15916 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_167
timestamp 1659098407
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_169
timestamp 1659098407
transform 1 0 16652 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_181
timestamp 1659098407
transform 1 0 17756 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_193
timestamp 1659098407
transform 1 0 18860 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_205
timestamp 1659098407
transform 1 0 19964 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_217
timestamp 1659098407
transform 1 0 21068 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_223
timestamp 1659098407
transform 1 0 21620 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_225
timestamp 1659098407
transform 1 0 21804 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_237
timestamp 1659098407
transform 1 0 22908 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_249
timestamp 1659098407
transform 1 0 24012 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_261
timestamp 1659098407
transform 1 0 25116 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_273
timestamp 1659098407
transform 1 0 26220 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_279
timestamp 1659098407
transform 1 0 26772 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_281
timestamp 1659098407
transform 1 0 26956 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_293
timestamp 1659098407
transform 1 0 28060 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_305
timestamp 1659098407
transform 1 0 29164 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_317
timestamp 1659098407
transform 1 0 30268 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_329
timestamp 1659098407
transform 1 0 31372 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_335
timestamp 1659098407
transform 1 0 31924 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_337
timestamp 1659098407
transform 1 0 32108 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_349
timestamp 1659098407
transform 1 0 33212 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_361
timestamp 1659098407
transform 1 0 34316 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_373
timestamp 1659098407
transform 1 0 35420 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_385
timestamp 1659098407
transform 1 0 36524 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_391
timestamp 1659098407
transform 1 0 37076 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_393
timestamp 1659098407
transform 1 0 37260 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_405
timestamp 1659098407
transform 1 0 38364 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_417
timestamp 1659098407
transform 1 0 39468 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_429
timestamp 1659098407
transform 1 0 40572 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_441
timestamp 1659098407
transform 1 0 41676 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_447
timestamp 1659098407
transform 1 0 42228 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_449
timestamp 1659098407
transform 1 0 42412 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_461
timestamp 1659098407
transform 1 0 43516 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_473
timestamp 1659098407
transform 1 0 44620 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_485
timestamp 1659098407
transform 1 0 45724 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_500
timestamp 1659098407
transform 1 0 47104 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_505
timestamp 1659098407
transform 1 0 47564 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_512
timestamp 1659098407
transform 1 0 48208 0 -1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3
timestamp 1659098407
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_15
timestamp 1659098407
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp 1659098407
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_29
timestamp 1659098407
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_41
timestamp 1659098407
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_53
timestamp 1659098407
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_65
timestamp 1659098407
transform 1 0 7084 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_77
timestamp 1659098407
transform 1 0 8188 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_83
timestamp 1659098407
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_85
timestamp 1659098407
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_97
timestamp 1659098407
transform 1 0 10028 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_109
timestamp 1659098407
transform 1 0 11132 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_121
timestamp 1659098407
transform 1 0 12236 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_133
timestamp 1659098407
transform 1 0 13340 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_139
timestamp 1659098407
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_141
timestamp 1659098407
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_153
timestamp 1659098407
transform 1 0 15180 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_165
timestamp 1659098407
transform 1 0 16284 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_177
timestamp 1659098407
transform 1 0 17388 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_189
timestamp 1659098407
transform 1 0 18492 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_195
timestamp 1659098407
transform 1 0 19044 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_197
timestamp 1659098407
transform 1 0 19228 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_209
timestamp 1659098407
transform 1 0 20332 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_221
timestamp 1659098407
transform 1 0 21436 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_233
timestamp 1659098407
transform 1 0 22540 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_245
timestamp 1659098407
transform 1 0 23644 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_251
timestamp 1659098407
transform 1 0 24196 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_253
timestamp 1659098407
transform 1 0 24380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_265
timestamp 1659098407
transform 1 0 25484 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_277
timestamp 1659098407
transform 1 0 26588 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_289
timestamp 1659098407
transform 1 0 27692 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_301
timestamp 1659098407
transform 1 0 28796 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_307
timestamp 1659098407
transform 1 0 29348 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_309
timestamp 1659098407
transform 1 0 29532 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_321
timestamp 1659098407
transform 1 0 30636 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_333
timestamp 1659098407
transform 1 0 31740 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_345
timestamp 1659098407
transform 1 0 32844 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_357
timestamp 1659098407
transform 1 0 33948 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_363
timestamp 1659098407
transform 1 0 34500 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_365
timestamp 1659098407
transform 1 0 34684 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_377
timestamp 1659098407
transform 1 0 35788 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_389
timestamp 1659098407
transform 1 0 36892 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_401
timestamp 1659098407
transform 1 0 37996 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_413
timestamp 1659098407
transform 1 0 39100 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_419
timestamp 1659098407
transform 1 0 39652 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_421
timestamp 1659098407
transform 1 0 39836 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_433
timestamp 1659098407
transform 1 0 40940 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_445
timestamp 1659098407
transform 1 0 42044 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_457
timestamp 1659098407
transform 1 0 43148 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_469
timestamp 1659098407
transform 1 0 44252 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_475
timestamp 1659098407
transform 1 0 44804 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_477
timestamp 1659098407
transform 1 0 44988 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_489
timestamp 1659098407
transform 1 0 46092 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_501
timestamp 1659098407
transform 1 0 47196 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_4_512
timestamp 1659098407
transform 1 0 48208 0 1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_5_6
timestamp 1659098407
transform 1 0 1656 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_18
timestamp 1659098407
transform 1 0 2760 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_30
timestamp 1659098407
transform 1 0 3864 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_42
timestamp 1659098407
transform 1 0 4968 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_5_54
timestamp 1659098407
transform 1 0 6072 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_5_57
timestamp 1659098407
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_69
timestamp 1659098407
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_81
timestamp 1659098407
transform 1 0 8556 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_93
timestamp 1659098407
transform 1 0 9660 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_105
timestamp 1659098407
transform 1 0 10764 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_111
timestamp 1659098407
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_113
timestamp 1659098407
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_125
timestamp 1659098407
transform 1 0 12604 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_137
timestamp 1659098407
transform 1 0 13708 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_149
timestamp 1659098407
transform 1 0 14812 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_161
timestamp 1659098407
transform 1 0 15916 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_167
timestamp 1659098407
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_169
timestamp 1659098407
transform 1 0 16652 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_181
timestamp 1659098407
transform 1 0 17756 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_193
timestamp 1659098407
transform 1 0 18860 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_205
timestamp 1659098407
transform 1 0 19964 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_217
timestamp 1659098407
transform 1 0 21068 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_223
timestamp 1659098407
transform 1 0 21620 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_225
timestamp 1659098407
transform 1 0 21804 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_237
timestamp 1659098407
transform 1 0 22908 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_249
timestamp 1659098407
transform 1 0 24012 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_261
timestamp 1659098407
transform 1 0 25116 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_273
timestamp 1659098407
transform 1 0 26220 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_279
timestamp 1659098407
transform 1 0 26772 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_281
timestamp 1659098407
transform 1 0 26956 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_293
timestamp 1659098407
transform 1 0 28060 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_305
timestamp 1659098407
transform 1 0 29164 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_317
timestamp 1659098407
transform 1 0 30268 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_329
timestamp 1659098407
transform 1 0 31372 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_335
timestamp 1659098407
transform 1 0 31924 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_337
timestamp 1659098407
transform 1 0 32108 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_349
timestamp 1659098407
transform 1 0 33212 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_361
timestamp 1659098407
transform 1 0 34316 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_373
timestamp 1659098407
transform 1 0 35420 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_385
timestamp 1659098407
transform 1 0 36524 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_391
timestamp 1659098407
transform 1 0 37076 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_393
timestamp 1659098407
transform 1 0 37260 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_405
timestamp 1659098407
transform 1 0 38364 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_417
timestamp 1659098407
transform 1 0 39468 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_429
timestamp 1659098407
transform 1 0 40572 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_441
timestamp 1659098407
transform 1 0 41676 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_447
timestamp 1659098407
transform 1 0 42228 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_449
timestamp 1659098407
transform 1 0 42412 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_461
timestamp 1659098407
transform 1 0 43516 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_473
timestamp 1659098407
transform 1 0 44620 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_485
timestamp 1659098407
transform 1 0 45724 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_497
timestamp 1659098407
transform 1 0 46828 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_503
timestamp 1659098407
transform 1 0 47380 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_505
timestamp 1659098407
transform 1 0 47564 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_512
timestamp 1659098407
transform 1 0 48208 0 -1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_6_6
timestamp 1659098407
transform 1 0 1656 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_18
timestamp 1659098407
transform 1 0 2760 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_6_26
timestamp 1659098407
transform 1 0 3496 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_6_29
timestamp 1659098407
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_41
timestamp 1659098407
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_53
timestamp 1659098407
transform 1 0 5980 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_65
timestamp 1659098407
transform 1 0 7084 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_77
timestamp 1659098407
transform 1 0 8188 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_83
timestamp 1659098407
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_85
timestamp 1659098407
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_97
timestamp 1659098407
transform 1 0 10028 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_109
timestamp 1659098407
transform 1 0 11132 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_121
timestamp 1659098407
transform 1 0 12236 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_133
timestamp 1659098407
transform 1 0 13340 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_139
timestamp 1659098407
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_141
timestamp 1659098407
transform 1 0 14076 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_153
timestamp 1659098407
transform 1 0 15180 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_165
timestamp 1659098407
transform 1 0 16284 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_177
timestamp 1659098407
transform 1 0 17388 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_189
timestamp 1659098407
transform 1 0 18492 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_195
timestamp 1659098407
transform 1 0 19044 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_197
timestamp 1659098407
transform 1 0 19228 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_209
timestamp 1659098407
transform 1 0 20332 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_221
timestamp 1659098407
transform 1 0 21436 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_233
timestamp 1659098407
transform 1 0 22540 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_245
timestamp 1659098407
transform 1 0 23644 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_251
timestamp 1659098407
transform 1 0 24196 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_253
timestamp 1659098407
transform 1 0 24380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_265
timestamp 1659098407
transform 1 0 25484 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_277
timestamp 1659098407
transform 1 0 26588 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_289
timestamp 1659098407
transform 1 0 27692 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_301
timestamp 1659098407
transform 1 0 28796 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_307
timestamp 1659098407
transform 1 0 29348 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_309
timestamp 1659098407
transform 1 0 29532 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_321
timestamp 1659098407
transform 1 0 30636 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_333
timestamp 1659098407
transform 1 0 31740 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_345
timestamp 1659098407
transform 1 0 32844 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_357
timestamp 1659098407
transform 1 0 33948 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_363
timestamp 1659098407
transform 1 0 34500 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_365
timestamp 1659098407
transform 1 0 34684 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_377
timestamp 1659098407
transform 1 0 35788 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_389
timestamp 1659098407
transform 1 0 36892 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_401
timestamp 1659098407
transform 1 0 37996 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_413
timestamp 1659098407
transform 1 0 39100 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_419
timestamp 1659098407
transform 1 0 39652 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_421
timestamp 1659098407
transform 1 0 39836 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_433
timestamp 1659098407
transform 1 0 40940 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_445
timestamp 1659098407
transform 1 0 42044 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_457
timestamp 1659098407
transform 1 0 43148 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_469
timestamp 1659098407
transform 1 0 44252 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_475
timestamp 1659098407
transform 1 0 44804 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_477
timestamp 1659098407
transform 1 0 44988 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_489
timestamp 1659098407
transform 1 0 46092 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_501
timestamp 1659098407
transform 1 0 47196 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_6_513
timestamp 1659098407
transform 1 0 48300 0 1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_7_6
timestamp 1659098407
transform 1 0 1656 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_18
timestamp 1659098407
transform 1 0 2760 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_30
timestamp 1659098407
transform 1 0 3864 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_42
timestamp 1659098407
transform 1 0 4968 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_7_54
timestamp 1659098407
transform 1 0 6072 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_7_57
timestamp 1659098407
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_69
timestamp 1659098407
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_81
timestamp 1659098407
transform 1 0 8556 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_93
timestamp 1659098407
transform 1 0 9660 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_105
timestamp 1659098407
transform 1 0 10764 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_111
timestamp 1659098407
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_113
timestamp 1659098407
transform 1 0 11500 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_125
timestamp 1659098407
transform 1 0 12604 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_137
timestamp 1659098407
transform 1 0 13708 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_149
timestamp 1659098407
transform 1 0 14812 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_161
timestamp 1659098407
transform 1 0 15916 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_167
timestamp 1659098407
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_169
timestamp 1659098407
transform 1 0 16652 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_181
timestamp 1659098407
transform 1 0 17756 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_193
timestamp 1659098407
transform 1 0 18860 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_205
timestamp 1659098407
transform 1 0 19964 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_217
timestamp 1659098407
transform 1 0 21068 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_223
timestamp 1659098407
transform 1 0 21620 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_225
timestamp 1659098407
transform 1 0 21804 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_237
timestamp 1659098407
transform 1 0 22908 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_249
timestamp 1659098407
transform 1 0 24012 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_261
timestamp 1659098407
transform 1 0 25116 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_273
timestamp 1659098407
transform 1 0 26220 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_279
timestamp 1659098407
transform 1 0 26772 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_281
timestamp 1659098407
transform 1 0 26956 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_293
timestamp 1659098407
transform 1 0 28060 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_305
timestamp 1659098407
transform 1 0 29164 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_317
timestamp 1659098407
transform 1 0 30268 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_329
timestamp 1659098407
transform 1 0 31372 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_335
timestamp 1659098407
transform 1 0 31924 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_337
timestamp 1659098407
transform 1 0 32108 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_349
timestamp 1659098407
transform 1 0 33212 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_361
timestamp 1659098407
transform 1 0 34316 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_373
timestamp 1659098407
transform 1 0 35420 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_385
timestamp 1659098407
transform 1 0 36524 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_391
timestamp 1659098407
transform 1 0 37076 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_393
timestamp 1659098407
transform 1 0 37260 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_405
timestamp 1659098407
transform 1 0 38364 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_417
timestamp 1659098407
transform 1 0 39468 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_429
timestamp 1659098407
transform 1 0 40572 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_441
timestamp 1659098407
transform 1 0 41676 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_447
timestamp 1659098407
transform 1 0 42228 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_449
timestamp 1659098407
transform 1 0 42412 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_461
timestamp 1659098407
transform 1 0 43516 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_473
timestamp 1659098407
transform 1 0 44620 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_485
timestamp 1659098407
transform 1 0 45724 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_497
timestamp 1659098407
transform 1 0 46828 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_503
timestamp 1659098407
transform 1 0 47380 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_505
timestamp 1659098407
transform 1 0 47564 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_512
timestamp 1659098407
transform 1 0 48208 0 -1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3
timestamp 1659098407
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_15
timestamp 1659098407
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp 1659098407
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_29
timestamp 1659098407
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_41
timestamp 1659098407
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_53
timestamp 1659098407
transform 1 0 5980 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_65
timestamp 1659098407
transform 1 0 7084 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_77
timestamp 1659098407
transform 1 0 8188 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_83
timestamp 1659098407
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_85
timestamp 1659098407
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_97
timestamp 1659098407
transform 1 0 10028 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_109
timestamp 1659098407
transform 1 0 11132 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_121
timestamp 1659098407
transform 1 0 12236 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_133
timestamp 1659098407
transform 1 0 13340 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_139
timestamp 1659098407
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_141
timestamp 1659098407
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_153
timestamp 1659098407
transform 1 0 15180 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_165
timestamp 1659098407
transform 1 0 16284 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_177
timestamp 1659098407
transform 1 0 17388 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_189
timestamp 1659098407
transform 1 0 18492 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_195
timestamp 1659098407
transform 1 0 19044 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_197
timestamp 1659098407
transform 1 0 19228 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_209
timestamp 1659098407
transform 1 0 20332 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_221
timestamp 1659098407
transform 1 0 21436 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_233
timestamp 1659098407
transform 1 0 22540 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_245
timestamp 1659098407
transform 1 0 23644 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_251
timestamp 1659098407
transform 1 0 24196 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_253
timestamp 1659098407
transform 1 0 24380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_265
timestamp 1659098407
transform 1 0 25484 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_277
timestamp 1659098407
transform 1 0 26588 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_289
timestamp 1659098407
transform 1 0 27692 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_301
timestamp 1659098407
transform 1 0 28796 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_307
timestamp 1659098407
transform 1 0 29348 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_309
timestamp 1659098407
transform 1 0 29532 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_321
timestamp 1659098407
transform 1 0 30636 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_333
timestamp 1659098407
transform 1 0 31740 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_345
timestamp 1659098407
transform 1 0 32844 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_357
timestamp 1659098407
transform 1 0 33948 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_363
timestamp 1659098407
transform 1 0 34500 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_365
timestamp 1659098407
transform 1 0 34684 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_377
timestamp 1659098407
transform 1 0 35788 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_389
timestamp 1659098407
transform 1 0 36892 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_401
timestamp 1659098407
transform 1 0 37996 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_413
timestamp 1659098407
transform 1 0 39100 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_419
timestamp 1659098407
transform 1 0 39652 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_421
timestamp 1659098407
transform 1 0 39836 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_433
timestamp 1659098407
transform 1 0 40940 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_445
timestamp 1659098407
transform 1 0 42044 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_457
timestamp 1659098407
transform 1 0 43148 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_469
timestamp 1659098407
transform 1 0 44252 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_475
timestamp 1659098407
transform 1 0 44804 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_477
timestamp 1659098407
transform 1 0 44988 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_489
timestamp 1659098407
transform 1 0 46092 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_501
timestamp 1659098407
transform 1 0 47196 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_8_513
timestamp 1659098407
transform 1 0 48300 0 1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_6
timestamp 1659098407
transform 1 0 1656 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_18
timestamp 1659098407
transform 1 0 2760 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_30
timestamp 1659098407
transform 1 0 3864 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_42
timestamp 1659098407
transform 1 0 4968 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_9_54
timestamp 1659098407
transform 1 0 6072 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_57
timestamp 1659098407
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_69
timestamp 1659098407
transform 1 0 7452 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_81
timestamp 1659098407
transform 1 0 8556 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_93
timestamp 1659098407
transform 1 0 9660 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_105
timestamp 1659098407
transform 1 0 10764 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_111
timestamp 1659098407
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_113
timestamp 1659098407
transform 1 0 11500 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_125
timestamp 1659098407
transform 1 0 12604 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_137
timestamp 1659098407
transform 1 0 13708 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_149
timestamp 1659098407
transform 1 0 14812 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_161
timestamp 1659098407
transform 1 0 15916 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_167
timestamp 1659098407
transform 1 0 16468 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_169
timestamp 1659098407
transform 1 0 16652 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_181
timestamp 1659098407
transform 1 0 17756 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_193
timestamp 1659098407
transform 1 0 18860 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_205
timestamp 1659098407
transform 1 0 19964 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_217
timestamp 1659098407
transform 1 0 21068 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_223
timestamp 1659098407
transform 1 0 21620 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_225
timestamp 1659098407
transform 1 0 21804 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_237
timestamp 1659098407
transform 1 0 22908 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_249
timestamp 1659098407
transform 1 0 24012 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_261
timestamp 1659098407
transform 1 0 25116 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_273
timestamp 1659098407
transform 1 0 26220 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_279
timestamp 1659098407
transform 1 0 26772 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_281
timestamp 1659098407
transform 1 0 26956 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_293
timestamp 1659098407
transform 1 0 28060 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_305
timestamp 1659098407
transform 1 0 29164 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_317
timestamp 1659098407
transform 1 0 30268 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_329
timestamp 1659098407
transform 1 0 31372 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_335
timestamp 1659098407
transform 1 0 31924 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_337
timestamp 1659098407
transform 1 0 32108 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_349
timestamp 1659098407
transform 1 0 33212 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_361
timestamp 1659098407
transform 1 0 34316 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_373
timestamp 1659098407
transform 1 0 35420 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_385
timestamp 1659098407
transform 1 0 36524 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_391
timestamp 1659098407
transform 1 0 37076 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_393
timestamp 1659098407
transform 1 0 37260 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_405
timestamp 1659098407
transform 1 0 38364 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_417
timestamp 1659098407
transform 1 0 39468 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_429
timestamp 1659098407
transform 1 0 40572 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_441
timestamp 1659098407
transform 1 0 41676 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_447
timestamp 1659098407
transform 1 0 42228 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_449
timestamp 1659098407
transform 1 0 42412 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_461
timestamp 1659098407
transform 1 0 43516 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_473
timestamp 1659098407
transform 1 0 44620 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_485
timestamp 1659098407
transform 1 0 45724 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_497
timestamp 1659098407
transform 1 0 46828 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_503
timestamp 1659098407
transform 1 0 47380 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_505
timestamp 1659098407
transform 1 0 47564 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_512
timestamp 1659098407
transform 1 0 48208 0 -1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_10_6
timestamp 1659098407
transform 1 0 1656 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_18
timestamp 1659098407
transform 1 0 2760 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_26
timestamp 1659098407
transform 1 0 3496 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_10_29
timestamp 1659098407
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_41
timestamp 1659098407
transform 1 0 4876 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_53
timestamp 1659098407
transform 1 0 5980 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_65
timestamp 1659098407
transform 1 0 7084 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_77
timestamp 1659098407
transform 1 0 8188 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_83
timestamp 1659098407
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_85
timestamp 1659098407
transform 1 0 8924 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_97
timestamp 1659098407
transform 1 0 10028 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_109
timestamp 1659098407
transform 1 0 11132 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_121
timestamp 1659098407
transform 1 0 12236 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_133
timestamp 1659098407
transform 1 0 13340 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_139
timestamp 1659098407
transform 1 0 13892 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_141
timestamp 1659098407
transform 1 0 14076 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_153
timestamp 1659098407
transform 1 0 15180 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_165
timestamp 1659098407
transform 1 0 16284 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_177
timestamp 1659098407
transform 1 0 17388 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_189
timestamp 1659098407
transform 1 0 18492 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_195
timestamp 1659098407
transform 1 0 19044 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_197
timestamp 1659098407
transform 1 0 19228 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_209
timestamp 1659098407
transform 1 0 20332 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_221
timestamp 1659098407
transform 1 0 21436 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_233
timestamp 1659098407
transform 1 0 22540 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_245
timestamp 1659098407
transform 1 0 23644 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_251
timestamp 1659098407
transform 1 0 24196 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_253
timestamp 1659098407
transform 1 0 24380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_265
timestamp 1659098407
transform 1 0 25484 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_277
timestamp 1659098407
transform 1 0 26588 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_289
timestamp 1659098407
transform 1 0 27692 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_301
timestamp 1659098407
transform 1 0 28796 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_307
timestamp 1659098407
transform 1 0 29348 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_309
timestamp 1659098407
transform 1 0 29532 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_321
timestamp 1659098407
transform 1 0 30636 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_333
timestamp 1659098407
transform 1 0 31740 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_345
timestamp 1659098407
transform 1 0 32844 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_357
timestamp 1659098407
transform 1 0 33948 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_363
timestamp 1659098407
transform 1 0 34500 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_365
timestamp 1659098407
transform 1 0 34684 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_377
timestamp 1659098407
transform 1 0 35788 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_389
timestamp 1659098407
transform 1 0 36892 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_401
timestamp 1659098407
transform 1 0 37996 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_413
timestamp 1659098407
transform 1 0 39100 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_419
timestamp 1659098407
transform 1 0 39652 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_421
timestamp 1659098407
transform 1 0 39836 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_433
timestamp 1659098407
transform 1 0 40940 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_445
timestamp 1659098407
transform 1 0 42044 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_457
timestamp 1659098407
transform 1 0 43148 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_469
timestamp 1659098407
transform 1 0 44252 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_475
timestamp 1659098407
transform 1 0 44804 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_477
timestamp 1659098407
transform 1 0 44988 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_489
timestamp 1659098407
transform 1 0 46092 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_501
timestamp 1659098407
transform 1 0 47196 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_10_512
timestamp 1659098407
transform 1 0 48208 0 1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_11_6
timestamp 1659098407
transform 1 0 1656 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_18
timestamp 1659098407
transform 1 0 2760 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_30
timestamp 1659098407
transform 1 0 3864 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_42
timestamp 1659098407
transform 1 0 4968 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_11_54
timestamp 1659098407
transform 1 0 6072 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_11_57
timestamp 1659098407
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_69
timestamp 1659098407
transform 1 0 7452 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_81
timestamp 1659098407
transform 1 0 8556 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_93
timestamp 1659098407
transform 1 0 9660 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_105
timestamp 1659098407
transform 1 0 10764 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_111
timestamp 1659098407
transform 1 0 11316 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_113
timestamp 1659098407
transform 1 0 11500 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_125
timestamp 1659098407
transform 1 0 12604 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_137
timestamp 1659098407
transform 1 0 13708 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_149
timestamp 1659098407
transform 1 0 14812 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_161
timestamp 1659098407
transform 1 0 15916 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_167
timestamp 1659098407
transform 1 0 16468 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_169
timestamp 1659098407
transform 1 0 16652 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_181
timestamp 1659098407
transform 1 0 17756 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_193
timestamp 1659098407
transform 1 0 18860 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_205
timestamp 1659098407
transform 1 0 19964 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_217
timestamp 1659098407
transform 1 0 21068 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_223
timestamp 1659098407
transform 1 0 21620 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_225
timestamp 1659098407
transform 1 0 21804 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_237
timestamp 1659098407
transform 1 0 22908 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_249
timestamp 1659098407
transform 1 0 24012 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_261
timestamp 1659098407
transform 1 0 25116 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_273
timestamp 1659098407
transform 1 0 26220 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_279
timestamp 1659098407
transform 1 0 26772 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_281
timestamp 1659098407
transform 1 0 26956 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_293
timestamp 1659098407
transform 1 0 28060 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_305
timestamp 1659098407
transform 1 0 29164 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_317
timestamp 1659098407
transform 1 0 30268 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_329
timestamp 1659098407
transform 1 0 31372 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_335
timestamp 1659098407
transform 1 0 31924 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_337
timestamp 1659098407
transform 1 0 32108 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_349
timestamp 1659098407
transform 1 0 33212 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_361
timestamp 1659098407
transform 1 0 34316 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_373
timestamp 1659098407
transform 1 0 35420 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_385
timestamp 1659098407
transform 1 0 36524 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_391
timestamp 1659098407
transform 1 0 37076 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_393
timestamp 1659098407
transform 1 0 37260 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_405
timestamp 1659098407
transform 1 0 38364 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_417
timestamp 1659098407
transform 1 0 39468 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_429
timestamp 1659098407
transform 1 0 40572 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_441
timestamp 1659098407
transform 1 0 41676 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_447
timestamp 1659098407
transform 1 0 42228 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_449
timestamp 1659098407
transform 1 0 42412 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_461
timestamp 1659098407
transform 1 0 43516 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_473
timestamp 1659098407
transform 1 0 44620 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_485
timestamp 1659098407
transform 1 0 45724 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_497
timestamp 1659098407
transform 1 0 46828 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_503
timestamp 1659098407
transform 1 0 47380 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_505
timestamp 1659098407
transform 1 0 47564 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_11_513
timestamp 1659098407
transform 1 0 48300 0 -1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_12_6
timestamp 1659098407
transform 1 0 1656 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_18
timestamp 1659098407
transform 1 0 2760 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_12_26
timestamp 1659098407
transform 1 0 3496 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_12_29
timestamp 1659098407
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_41
timestamp 1659098407
transform 1 0 4876 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_53
timestamp 1659098407
transform 1 0 5980 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_65
timestamp 1659098407
transform 1 0 7084 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_77
timestamp 1659098407
transform 1 0 8188 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_83
timestamp 1659098407
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_85
timestamp 1659098407
transform 1 0 8924 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_97
timestamp 1659098407
transform 1 0 10028 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_109
timestamp 1659098407
transform 1 0 11132 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_121
timestamp 1659098407
transform 1 0 12236 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_133
timestamp 1659098407
transform 1 0 13340 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_139
timestamp 1659098407
transform 1 0 13892 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_141
timestamp 1659098407
transform 1 0 14076 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_153
timestamp 1659098407
transform 1 0 15180 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_165
timestamp 1659098407
transform 1 0 16284 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_177
timestamp 1659098407
transform 1 0 17388 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_189
timestamp 1659098407
transform 1 0 18492 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_195
timestamp 1659098407
transform 1 0 19044 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_197
timestamp 1659098407
transform 1 0 19228 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_209
timestamp 1659098407
transform 1 0 20332 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_221
timestamp 1659098407
transform 1 0 21436 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_233
timestamp 1659098407
transform 1 0 22540 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_245
timestamp 1659098407
transform 1 0 23644 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_251
timestamp 1659098407
transform 1 0 24196 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_253
timestamp 1659098407
transform 1 0 24380 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_265
timestamp 1659098407
transform 1 0 25484 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_277
timestamp 1659098407
transform 1 0 26588 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_289
timestamp 1659098407
transform 1 0 27692 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_301
timestamp 1659098407
transform 1 0 28796 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_307
timestamp 1659098407
transform 1 0 29348 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_309
timestamp 1659098407
transform 1 0 29532 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_321
timestamp 1659098407
transform 1 0 30636 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_333
timestamp 1659098407
transform 1 0 31740 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_345
timestamp 1659098407
transform 1 0 32844 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_357
timestamp 1659098407
transform 1 0 33948 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_363
timestamp 1659098407
transform 1 0 34500 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_365
timestamp 1659098407
transform 1 0 34684 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_377
timestamp 1659098407
transform 1 0 35788 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_389
timestamp 1659098407
transform 1 0 36892 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_401
timestamp 1659098407
transform 1 0 37996 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_413
timestamp 1659098407
transform 1 0 39100 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_419
timestamp 1659098407
transform 1 0 39652 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_421
timestamp 1659098407
transform 1 0 39836 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_433
timestamp 1659098407
transform 1 0 40940 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_445
timestamp 1659098407
transform 1 0 42044 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_457
timestamp 1659098407
transform 1 0 43148 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_469
timestamp 1659098407
transform 1 0 44252 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_475
timestamp 1659098407
transform 1 0 44804 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_477
timestamp 1659098407
transform 1 0 44988 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_489
timestamp 1659098407
transform 1 0 46092 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_501
timestamp 1659098407
transform 1 0 47196 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_12_512
timestamp 1659098407
transform 1 0 48208 0 1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_13_3
timestamp 1659098407
transform 1 0 1380 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_15
timestamp 1659098407
transform 1 0 2484 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_27
timestamp 1659098407
transform 1 0 3588 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_39
timestamp 1659098407
transform 1 0 4692 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_51
timestamp 1659098407
transform 1 0 5796 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_55
timestamp 1659098407
transform 1 0 6164 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_57
timestamp 1659098407
transform 1 0 6348 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_69
timestamp 1659098407
transform 1 0 7452 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_81
timestamp 1659098407
transform 1 0 8556 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_93
timestamp 1659098407
transform 1 0 9660 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_105
timestamp 1659098407
transform 1 0 10764 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_111
timestamp 1659098407
transform 1 0 11316 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_113
timestamp 1659098407
transform 1 0 11500 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_125
timestamp 1659098407
transform 1 0 12604 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_137
timestamp 1659098407
transform 1 0 13708 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_149
timestamp 1659098407
transform 1 0 14812 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_161
timestamp 1659098407
transform 1 0 15916 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_167
timestamp 1659098407
transform 1 0 16468 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_169
timestamp 1659098407
transform 1 0 16652 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_181
timestamp 1659098407
transform 1 0 17756 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_193
timestamp 1659098407
transform 1 0 18860 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_205
timestamp 1659098407
transform 1 0 19964 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_217
timestamp 1659098407
transform 1 0 21068 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_223
timestamp 1659098407
transform 1 0 21620 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_225
timestamp 1659098407
transform 1 0 21804 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_237
timestamp 1659098407
transform 1 0 22908 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_249
timestamp 1659098407
transform 1 0 24012 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_261
timestamp 1659098407
transform 1 0 25116 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_273
timestamp 1659098407
transform 1 0 26220 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_279
timestamp 1659098407
transform 1 0 26772 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_281
timestamp 1659098407
transform 1 0 26956 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_293
timestamp 1659098407
transform 1 0 28060 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_305
timestamp 1659098407
transform 1 0 29164 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_317
timestamp 1659098407
transform 1 0 30268 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_329
timestamp 1659098407
transform 1 0 31372 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_335
timestamp 1659098407
transform 1 0 31924 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_337
timestamp 1659098407
transform 1 0 32108 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_349
timestamp 1659098407
transform 1 0 33212 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_361
timestamp 1659098407
transform 1 0 34316 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_373
timestamp 1659098407
transform 1 0 35420 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_385
timestamp 1659098407
transform 1 0 36524 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_391
timestamp 1659098407
transform 1 0 37076 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_393
timestamp 1659098407
transform 1 0 37260 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_405
timestamp 1659098407
transform 1 0 38364 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_417
timestamp 1659098407
transform 1 0 39468 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_429
timestamp 1659098407
transform 1 0 40572 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_441
timestamp 1659098407
transform 1 0 41676 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_447
timestamp 1659098407
transform 1 0 42228 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_449
timestamp 1659098407
transform 1 0 42412 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_461
timestamp 1659098407
transform 1 0 43516 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_473
timestamp 1659098407
transform 1 0 44620 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_485
timestamp 1659098407
transform 1 0 45724 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_13_492
timestamp 1659098407
transform 1 0 46368 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_505
timestamp 1659098407
transform 1 0 47564 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_13_513
timestamp 1659098407
transform 1 0 48300 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_14_3
timestamp 1659098407
transform 1 0 1380 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_15
timestamp 1659098407
transform 1 0 2484 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_27
timestamp 1659098407
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_29
timestamp 1659098407
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_41
timestamp 1659098407
transform 1 0 4876 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_53
timestamp 1659098407
transform 1 0 5980 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_65
timestamp 1659098407
transform 1 0 7084 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_77
timestamp 1659098407
transform 1 0 8188 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_83
timestamp 1659098407
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_85
timestamp 1659098407
transform 1 0 8924 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_97
timestamp 1659098407
transform 1 0 10028 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_109
timestamp 1659098407
transform 1 0 11132 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_121
timestamp 1659098407
transform 1 0 12236 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_133
timestamp 1659098407
transform 1 0 13340 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_139
timestamp 1659098407
transform 1 0 13892 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_141
timestamp 1659098407
transform 1 0 14076 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_153
timestamp 1659098407
transform 1 0 15180 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_165
timestamp 1659098407
transform 1 0 16284 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_177
timestamp 1659098407
transform 1 0 17388 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_189
timestamp 1659098407
transform 1 0 18492 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_195
timestamp 1659098407
transform 1 0 19044 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_197
timestamp 1659098407
transform 1 0 19228 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_209
timestamp 1659098407
transform 1 0 20332 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_221
timestamp 1659098407
transform 1 0 21436 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_233
timestamp 1659098407
transform 1 0 22540 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_245
timestamp 1659098407
transform 1 0 23644 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_251
timestamp 1659098407
transform 1 0 24196 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_253
timestamp 1659098407
transform 1 0 24380 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_265
timestamp 1659098407
transform 1 0 25484 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_277
timestamp 1659098407
transform 1 0 26588 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_289
timestamp 1659098407
transform 1 0 27692 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_301
timestamp 1659098407
transform 1 0 28796 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_307
timestamp 1659098407
transform 1 0 29348 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_309
timestamp 1659098407
transform 1 0 29532 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_321
timestamp 1659098407
transform 1 0 30636 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_333
timestamp 1659098407
transform 1 0 31740 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_345
timestamp 1659098407
transform 1 0 32844 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_357
timestamp 1659098407
transform 1 0 33948 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_363
timestamp 1659098407
transform 1 0 34500 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_365
timestamp 1659098407
transform 1 0 34684 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_377
timestamp 1659098407
transform 1 0 35788 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_389
timestamp 1659098407
transform 1 0 36892 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_401
timestamp 1659098407
transform 1 0 37996 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_413
timestamp 1659098407
transform 1 0 39100 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_419
timestamp 1659098407
transform 1 0 39652 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_421
timestamp 1659098407
transform 1 0 39836 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_433
timestamp 1659098407
transform 1 0 40940 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_445
timestamp 1659098407
transform 1 0 42044 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_457
timestamp 1659098407
transform 1 0 43148 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_469
timestamp 1659098407
transform 1 0 44252 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_475
timestamp 1659098407
transform 1 0 44804 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_477
timestamp 1659098407
transform 1 0 44988 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_489
timestamp 1659098407
transform 1 0 46092 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_501
timestamp 1659098407
transform 1 0 47196 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_14_512
timestamp 1659098407
transform 1 0 48208 0 1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_15_3
timestamp 1659098407
transform 1 0 1380 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_15
timestamp 1659098407
transform 1 0 2484 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_27
timestamp 1659098407
transform 1 0 3588 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_39
timestamp 1659098407
transform 1 0 4692 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_51
timestamp 1659098407
transform 1 0 5796 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_55
timestamp 1659098407
transform 1 0 6164 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_57
timestamp 1659098407
transform 1 0 6348 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_69
timestamp 1659098407
transform 1 0 7452 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_81
timestamp 1659098407
transform 1 0 8556 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_93
timestamp 1659098407
transform 1 0 9660 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_105
timestamp 1659098407
transform 1 0 10764 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_111
timestamp 1659098407
transform 1 0 11316 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_113
timestamp 1659098407
transform 1 0 11500 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_125
timestamp 1659098407
transform 1 0 12604 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_137
timestamp 1659098407
transform 1 0 13708 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_149
timestamp 1659098407
transform 1 0 14812 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_161
timestamp 1659098407
transform 1 0 15916 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_167
timestamp 1659098407
transform 1 0 16468 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_169
timestamp 1659098407
transform 1 0 16652 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_181
timestamp 1659098407
transform 1 0 17756 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_193
timestamp 1659098407
transform 1 0 18860 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_205
timestamp 1659098407
transform 1 0 19964 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_217
timestamp 1659098407
transform 1 0 21068 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_223
timestamp 1659098407
transform 1 0 21620 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_225
timestamp 1659098407
transform 1 0 21804 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_237
timestamp 1659098407
transform 1 0 22908 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_249
timestamp 1659098407
transform 1 0 24012 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_261
timestamp 1659098407
transform 1 0 25116 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_273
timestamp 1659098407
transform 1 0 26220 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_279
timestamp 1659098407
transform 1 0 26772 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_281
timestamp 1659098407
transform 1 0 26956 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_293
timestamp 1659098407
transform 1 0 28060 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_305
timestamp 1659098407
transform 1 0 29164 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_317
timestamp 1659098407
transform 1 0 30268 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_329
timestamp 1659098407
transform 1 0 31372 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_335
timestamp 1659098407
transform 1 0 31924 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_337
timestamp 1659098407
transform 1 0 32108 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_349
timestamp 1659098407
transform 1 0 33212 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_361
timestamp 1659098407
transform 1 0 34316 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_373
timestamp 1659098407
transform 1 0 35420 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_385
timestamp 1659098407
transform 1 0 36524 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_391
timestamp 1659098407
transform 1 0 37076 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_393
timestamp 1659098407
transform 1 0 37260 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_405
timestamp 1659098407
transform 1 0 38364 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_417
timestamp 1659098407
transform 1 0 39468 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_429
timestamp 1659098407
transform 1 0 40572 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_441
timestamp 1659098407
transform 1 0 41676 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_447
timestamp 1659098407
transform 1 0 42228 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_449
timestamp 1659098407
transform 1 0 42412 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_461
timestamp 1659098407
transform 1 0 43516 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_473
timestamp 1659098407
transform 1 0 44620 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_485
timestamp 1659098407
transform 1 0 45724 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_497
timestamp 1659098407
transform 1 0 46828 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_503
timestamp 1659098407
transform 1 0 47380 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_508
timestamp 1659098407
transform 1 0 47840 0 -1 10880
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_16_6
timestamp 1659098407
transform 1 0 1656 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_18
timestamp 1659098407
transform 1 0 2760 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_26
timestamp 1659098407
transform 1 0 3496 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_16_29
timestamp 1659098407
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_41
timestamp 1659098407
transform 1 0 4876 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_53
timestamp 1659098407
transform 1 0 5980 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_65
timestamp 1659098407
transform 1 0 7084 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_77
timestamp 1659098407
transform 1 0 8188 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_83
timestamp 1659098407
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_85
timestamp 1659098407
transform 1 0 8924 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_97
timestamp 1659098407
transform 1 0 10028 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_109
timestamp 1659098407
transform 1 0 11132 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_121
timestamp 1659098407
transform 1 0 12236 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_133
timestamp 1659098407
transform 1 0 13340 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_139
timestamp 1659098407
transform 1 0 13892 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_141
timestamp 1659098407
transform 1 0 14076 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_153
timestamp 1659098407
transform 1 0 15180 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_165
timestamp 1659098407
transform 1 0 16284 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_177
timestamp 1659098407
transform 1 0 17388 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_189
timestamp 1659098407
transform 1 0 18492 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_195
timestamp 1659098407
transform 1 0 19044 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_197
timestamp 1659098407
transform 1 0 19228 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_209
timestamp 1659098407
transform 1 0 20332 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_221
timestamp 1659098407
transform 1 0 21436 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_233
timestamp 1659098407
transform 1 0 22540 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_245
timestamp 1659098407
transform 1 0 23644 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_251
timestamp 1659098407
transform 1 0 24196 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_253
timestamp 1659098407
transform 1 0 24380 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_265
timestamp 1659098407
transform 1 0 25484 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_277
timestamp 1659098407
transform 1 0 26588 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_289
timestamp 1659098407
transform 1 0 27692 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_301
timestamp 1659098407
transform 1 0 28796 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_307
timestamp 1659098407
transform 1 0 29348 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_309
timestamp 1659098407
transform 1 0 29532 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_321
timestamp 1659098407
transform 1 0 30636 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_333
timestamp 1659098407
transform 1 0 31740 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_345
timestamp 1659098407
transform 1 0 32844 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_357
timestamp 1659098407
transform 1 0 33948 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_363
timestamp 1659098407
transform 1 0 34500 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_365
timestamp 1659098407
transform 1 0 34684 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_377
timestamp 1659098407
transform 1 0 35788 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_389
timestamp 1659098407
transform 1 0 36892 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_401
timestamp 1659098407
transform 1 0 37996 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_413
timestamp 1659098407
transform 1 0 39100 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_419
timestamp 1659098407
transform 1 0 39652 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_421
timestamp 1659098407
transform 1 0 39836 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_433
timestamp 1659098407
transform 1 0 40940 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_445
timestamp 1659098407
transform 1 0 42044 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_457
timestamp 1659098407
transform 1 0 43148 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_469
timestamp 1659098407
transform 1 0 44252 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_475
timestamp 1659098407
transform 1 0 44804 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_477
timestamp 1659098407
transform 1 0 44988 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_489
timestamp 1659098407
transform 1 0 46092 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_497
timestamp 1659098407
transform 1 0 46828 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_504
timestamp 1659098407
transform 1 0 47472 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_6
timestamp 1659098407
transform 1 0 1656 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_18
timestamp 1659098407
transform 1 0 2760 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_30
timestamp 1659098407
transform 1 0 3864 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_42
timestamp 1659098407
transform 1 0 4968 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_17_54
timestamp 1659098407
transform 1 0 6072 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_17_57
timestamp 1659098407
transform 1 0 6348 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_69
timestamp 1659098407
transform 1 0 7452 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_81
timestamp 1659098407
transform 1 0 8556 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_93
timestamp 1659098407
transform 1 0 9660 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_105
timestamp 1659098407
transform 1 0 10764 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_111
timestamp 1659098407
transform 1 0 11316 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_113
timestamp 1659098407
transform 1 0 11500 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_125
timestamp 1659098407
transform 1 0 12604 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_137
timestamp 1659098407
transform 1 0 13708 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_149
timestamp 1659098407
transform 1 0 14812 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_161
timestamp 1659098407
transform 1 0 15916 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_167
timestamp 1659098407
transform 1 0 16468 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_169
timestamp 1659098407
transform 1 0 16652 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_181
timestamp 1659098407
transform 1 0 17756 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_193
timestamp 1659098407
transform 1 0 18860 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_205
timestamp 1659098407
transform 1 0 19964 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_217
timestamp 1659098407
transform 1 0 21068 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_223
timestamp 1659098407
transform 1 0 21620 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_225
timestamp 1659098407
transform 1 0 21804 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_237
timestamp 1659098407
transform 1 0 22908 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_249
timestamp 1659098407
transform 1 0 24012 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_261
timestamp 1659098407
transform 1 0 25116 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_273
timestamp 1659098407
transform 1 0 26220 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_279
timestamp 1659098407
transform 1 0 26772 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_281
timestamp 1659098407
transform 1 0 26956 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_293
timestamp 1659098407
transform 1 0 28060 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_305
timestamp 1659098407
transform 1 0 29164 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_317
timestamp 1659098407
transform 1 0 30268 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_329
timestamp 1659098407
transform 1 0 31372 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_335
timestamp 1659098407
transform 1 0 31924 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_337
timestamp 1659098407
transform 1 0 32108 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_349
timestamp 1659098407
transform 1 0 33212 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_361
timestamp 1659098407
transform 1 0 34316 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_373
timestamp 1659098407
transform 1 0 35420 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_385
timestamp 1659098407
transform 1 0 36524 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_391
timestamp 1659098407
transform 1 0 37076 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_393
timestamp 1659098407
transform 1 0 37260 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_405
timestamp 1659098407
transform 1 0 38364 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_417
timestamp 1659098407
transform 1 0 39468 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_429
timestamp 1659098407
transform 1 0 40572 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_441
timestamp 1659098407
transform 1 0 41676 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_447
timestamp 1659098407
transform 1 0 42228 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_449
timestamp 1659098407
transform 1 0 42412 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_461
timestamp 1659098407
transform 1 0 43516 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_473
timestamp 1659098407
transform 1 0 44620 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_485
timestamp 1659098407
transform 1 0 45724 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_497
timestamp 1659098407
transform 1 0 46828 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_503
timestamp 1659098407
transform 1 0 47380 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_505
timestamp 1659098407
transform 1 0 47564 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_512
timestamp 1659098407
transform 1 0 48208 0 -1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_18_3
timestamp 1659098407
transform 1 0 1380 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_15
timestamp 1659098407
transform 1 0 2484 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_27
timestamp 1659098407
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_29
timestamp 1659098407
transform 1 0 3772 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_41
timestamp 1659098407
transform 1 0 4876 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_53
timestamp 1659098407
transform 1 0 5980 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_65
timestamp 1659098407
transform 1 0 7084 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_77
timestamp 1659098407
transform 1 0 8188 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_83
timestamp 1659098407
transform 1 0 8740 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_85
timestamp 1659098407
transform 1 0 8924 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_97
timestamp 1659098407
transform 1 0 10028 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_109
timestamp 1659098407
transform 1 0 11132 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_121
timestamp 1659098407
transform 1 0 12236 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_133
timestamp 1659098407
transform 1 0 13340 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_139
timestamp 1659098407
transform 1 0 13892 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_141
timestamp 1659098407
transform 1 0 14076 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_153
timestamp 1659098407
transform 1 0 15180 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_165
timestamp 1659098407
transform 1 0 16284 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_177
timestamp 1659098407
transform 1 0 17388 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_189
timestamp 1659098407
transform 1 0 18492 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_195
timestamp 1659098407
transform 1 0 19044 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_197
timestamp 1659098407
transform 1 0 19228 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_209
timestamp 1659098407
transform 1 0 20332 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_221
timestamp 1659098407
transform 1 0 21436 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_233
timestamp 1659098407
transform 1 0 22540 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_245
timestamp 1659098407
transform 1 0 23644 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_251
timestamp 1659098407
transform 1 0 24196 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_253
timestamp 1659098407
transform 1 0 24380 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_265
timestamp 1659098407
transform 1 0 25484 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_277
timestamp 1659098407
transform 1 0 26588 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_289
timestamp 1659098407
transform 1 0 27692 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_301
timestamp 1659098407
transform 1 0 28796 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_307
timestamp 1659098407
transform 1 0 29348 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_309
timestamp 1659098407
transform 1 0 29532 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_321
timestamp 1659098407
transform 1 0 30636 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_333
timestamp 1659098407
transform 1 0 31740 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_345
timestamp 1659098407
transform 1 0 32844 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_357
timestamp 1659098407
transform 1 0 33948 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_363
timestamp 1659098407
transform 1 0 34500 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_365
timestamp 1659098407
transform 1 0 34684 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_377
timestamp 1659098407
transform 1 0 35788 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_389
timestamp 1659098407
transform 1 0 36892 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_401
timestamp 1659098407
transform 1 0 37996 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_413
timestamp 1659098407
transform 1 0 39100 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_419
timestamp 1659098407
transform 1 0 39652 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_421
timestamp 1659098407
transform 1 0 39836 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_433
timestamp 1659098407
transform 1 0 40940 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_445
timestamp 1659098407
transform 1 0 42044 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_457
timestamp 1659098407
transform 1 0 43148 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_469
timestamp 1659098407
transform 1 0 44252 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_475
timestamp 1659098407
transform 1 0 44804 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_477
timestamp 1659098407
transform 1 0 44988 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_489
timestamp 1659098407
transform 1 0 46092 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_501
timestamp 1659098407
transform 1 0 47196 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_18_512
timestamp 1659098407
transform 1 0 48208 0 1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_19_6
timestamp 1659098407
transform 1 0 1656 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_18
timestamp 1659098407
transform 1 0 2760 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_30
timestamp 1659098407
transform 1 0 3864 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_42
timestamp 1659098407
transform 1 0 4968 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_19_54
timestamp 1659098407
transform 1 0 6072 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_19_57
timestamp 1659098407
transform 1 0 6348 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_69
timestamp 1659098407
transform 1 0 7452 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_81
timestamp 1659098407
transform 1 0 8556 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_93
timestamp 1659098407
transform 1 0 9660 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_105
timestamp 1659098407
transform 1 0 10764 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_111
timestamp 1659098407
transform 1 0 11316 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_113
timestamp 1659098407
transform 1 0 11500 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_125
timestamp 1659098407
transform 1 0 12604 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_137
timestamp 1659098407
transform 1 0 13708 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_149
timestamp 1659098407
transform 1 0 14812 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_161
timestamp 1659098407
transform 1 0 15916 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_167
timestamp 1659098407
transform 1 0 16468 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_169
timestamp 1659098407
transform 1 0 16652 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_181
timestamp 1659098407
transform 1 0 17756 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_193
timestamp 1659098407
transform 1 0 18860 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_205
timestamp 1659098407
transform 1 0 19964 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_217
timestamp 1659098407
transform 1 0 21068 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_223
timestamp 1659098407
transform 1 0 21620 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_225
timestamp 1659098407
transform 1 0 21804 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_237
timestamp 1659098407
transform 1 0 22908 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_249
timestamp 1659098407
transform 1 0 24012 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_261
timestamp 1659098407
transform 1 0 25116 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_273
timestamp 1659098407
transform 1 0 26220 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_279
timestamp 1659098407
transform 1 0 26772 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_281
timestamp 1659098407
transform 1 0 26956 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_293
timestamp 1659098407
transform 1 0 28060 0 -1 13056
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_19_319
timestamp 1659098407
transform 1 0 30452 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_331
timestamp 1659098407
transform 1 0 31556 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_335
timestamp 1659098407
transform 1 0 31924 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_337
timestamp 1659098407
transform 1 0 32108 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_349
timestamp 1659098407
transform 1 0 33212 0 -1 13056
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_19_375
timestamp 1659098407
transform 1 0 35604 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_387
timestamp 1659098407
transform 1 0 36708 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_391
timestamp 1659098407
transform 1 0 37076 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_393
timestamp 1659098407
transform 1 0 37260 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_405
timestamp 1659098407
transform 1 0 38364 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_417
timestamp 1659098407
transform 1 0 39468 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_19_429
timestamp 1659098407
transform 1 0 40572 0 -1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_19_435
timestamp 1659098407
transform 1 0 41124 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_19_447
timestamp 1659098407
transform 1 0 42228 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_449
timestamp 1659098407
transform 1 0 42412 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_461
timestamp 1659098407
transform 1 0 43516 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_473
timestamp 1659098407
transform 1 0 44620 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_480
timestamp 1659098407
transform 1 0 45264 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_487
timestamp 1659098407
transform 1 0 45908 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_19_494
timestamp 1659098407
transform 1 0 46552 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_502
timestamp 1659098407
transform 1 0 47288 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_19_508
timestamp 1659098407
transform 1 0 47840 0 -1 13056
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_20_3
timestamp 1659098407
transform 1 0 1380 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_15
timestamp 1659098407
transform 1 0 2484 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_27
timestamp 1659098407
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_29
timestamp 1659098407
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_41
timestamp 1659098407
transform 1 0 4876 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_53
timestamp 1659098407
transform 1 0 5980 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_65
timestamp 1659098407
transform 1 0 7084 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_77
timestamp 1659098407
transform 1 0 8188 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_83
timestamp 1659098407
transform 1 0 8740 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_85
timestamp 1659098407
transform 1 0 8924 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_97
timestamp 1659098407
transform 1 0 10028 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_109
timestamp 1659098407
transform 1 0 11132 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_121
timestamp 1659098407
transform 1 0 12236 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_133
timestamp 1659098407
transform 1 0 13340 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_139
timestamp 1659098407
transform 1 0 13892 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_141
timestamp 1659098407
transform 1 0 14076 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_153
timestamp 1659098407
transform 1 0 15180 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_165
timestamp 1659098407
transform 1 0 16284 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_177
timestamp 1659098407
transform 1 0 17388 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_189
timestamp 1659098407
transform 1 0 18492 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_195
timestamp 1659098407
transform 1 0 19044 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_197
timestamp 1659098407
transform 1 0 19228 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_209
timestamp 1659098407
transform 1 0 20332 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_221
timestamp 1659098407
transform 1 0 21436 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_229
timestamp 1659098407
transform 1 0 22172 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_20_235
timestamp 1659098407
transform 1 0 22724 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_247
timestamp 1659098407
transform 1 0 23828 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_251
timestamp 1659098407
transform 1 0 24196 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_253
timestamp 1659098407
transform 1 0 24380 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_265
timestamp 1659098407
transform 1 0 25484 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_277
timestamp 1659098407
transform 1 0 26588 0 1 13056
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_20_293
timestamp 1659098407
transform 1 0 28060 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_20_305
timestamp 1659098407
transform 1 0 29164 0 1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_20_309
timestamp 1659098407
transform 1 0 29532 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_321
timestamp 1659098407
transform 1 0 30636 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_333
timestamp 1659098407
transform 1 0 31740 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_339
timestamp 1659098407
transform 1 0 32292 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_348
timestamp 1659098407
transform 1 0 33120 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_360
timestamp 1659098407
transform 1 0 34224 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_365
timestamp 1659098407
transform 1 0 34684 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_20_387
timestamp 1659098407
transform 1 0 36708 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_399
timestamp 1659098407
transform 1 0 37812 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_411
timestamp 1659098407
transform 1 0 38916 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_419
timestamp 1659098407
transform 1 0 39652 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_421
timestamp 1659098407
transform 1 0 39836 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_433
timestamp 1659098407
transform 1 0 40940 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_445
timestamp 1659098407
transform 1 0 42044 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_457
timestamp 1659098407
transform 1 0 43148 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_469
timestamp 1659098407
transform 1 0 44252 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_475
timestamp 1659098407
transform 1 0 44804 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_477
timestamp 1659098407
transform 1 0 44988 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_489
timestamp 1659098407
transform 1 0 46092 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_501
timestamp 1659098407
transform 1 0 47196 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_20_512
timestamp 1659098407
transform 1 0 48208 0 1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_21_6
timestamp 1659098407
transform 1 0 1656 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_18
timestamp 1659098407
transform 1 0 2760 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_30
timestamp 1659098407
transform 1 0 3864 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_42
timestamp 1659098407
transform 1 0 4968 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_21_54
timestamp 1659098407
transform 1 0 6072 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_21_57
timestamp 1659098407
transform 1 0 6348 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_69
timestamp 1659098407
transform 1 0 7452 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_81
timestamp 1659098407
transform 1 0 8556 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_93
timestamp 1659098407
transform 1 0 9660 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_105
timestamp 1659098407
transform 1 0 10764 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_111
timestamp 1659098407
transform 1 0 11316 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_113
timestamp 1659098407
transform 1 0 11500 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_125
timestamp 1659098407
transform 1 0 12604 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_137
timestamp 1659098407
transform 1 0 13708 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_149
timestamp 1659098407
transform 1 0 14812 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_161
timestamp 1659098407
transform 1 0 15916 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_167
timestamp 1659098407
transform 1 0 16468 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_169
timestamp 1659098407
transform 1 0 16652 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_181
timestamp 1659098407
transform 1 0 17756 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_193
timestamp 1659098407
transform 1 0 18860 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_205
timestamp 1659098407
transform 1 0 19964 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_217
timestamp 1659098407
transform 1 0 21068 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_223
timestamp 1659098407
transform 1 0 21620 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_225
timestamp 1659098407
transform 1 0 21804 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_237
timestamp 1659098407
transform 1 0 22908 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_249
timestamp 1659098407
transform 1 0 24012 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_255
timestamp 1659098407
transform 1 0 24564 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_276
timestamp 1659098407
transform 1 0 26496 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_21_281
timestamp 1659098407
transform 1 0 26956 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_289
timestamp 1659098407
transform 1 0 27692 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_21_311
timestamp 1659098407
transform 1 0 29716 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_323
timestamp 1659098407
transform 1 0 30820 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_21_335
timestamp 1659098407
transform 1 0 31924 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_337
timestamp 1659098407
transform 1 0 32108 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_345
timestamp 1659098407
transform 1 0 32844 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_21_367
timestamp 1659098407
transform 1 0 34868 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_379
timestamp 1659098407
transform 1 0 35972 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_21_391
timestamp 1659098407
transform 1 0 37076 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_393
timestamp 1659098407
transform 1 0 37260 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_405
timestamp 1659098407
transform 1 0 38364 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_417
timestamp 1659098407
transform 1 0 39468 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_429
timestamp 1659098407
transform 1 0 40572 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_441
timestamp 1659098407
transform 1 0 41676 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_447
timestamp 1659098407
transform 1 0 42228 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_449
timestamp 1659098407
transform 1 0 42412 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_457
timestamp 1659098407
transform 1 0 43148 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_478
timestamp 1659098407
transform 1 0 45080 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_490
timestamp 1659098407
transform 1 0 46184 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_21_502
timestamp 1659098407
transform 1 0 47288 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_505
timestamp 1659098407
transform 1 0 47564 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_512
timestamp 1659098407
transform 1 0 48208 0 -1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_22_6
timestamp 1659098407
transform 1 0 1656 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_18
timestamp 1659098407
transform 1 0 2760 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_26
timestamp 1659098407
transform 1 0 3496 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_22_29
timestamp 1659098407
transform 1 0 3772 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_41
timestamp 1659098407
transform 1 0 4876 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_53
timestamp 1659098407
transform 1 0 5980 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_65
timestamp 1659098407
transform 1 0 7084 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_77
timestamp 1659098407
transform 1 0 8188 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_83
timestamp 1659098407
transform 1 0 8740 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_85
timestamp 1659098407
transform 1 0 8924 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_97
timestamp 1659098407
transform 1 0 10028 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_109
timestamp 1659098407
transform 1 0 11132 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_121
timestamp 1659098407
transform 1 0 12236 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_133
timestamp 1659098407
transform 1 0 13340 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_139
timestamp 1659098407
transform 1 0 13892 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_141
timestamp 1659098407
transform 1 0 14076 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_153
timestamp 1659098407
transform 1 0 15180 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_165
timestamp 1659098407
transform 1 0 16284 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_177
timestamp 1659098407
transform 1 0 17388 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_189
timestamp 1659098407
transform 1 0 18492 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_195
timestamp 1659098407
transform 1 0 19044 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_197
timestamp 1659098407
transform 1 0 19228 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_209
timestamp 1659098407
transform 1 0 20332 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_221
timestamp 1659098407
transform 1 0 21436 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_233
timestamp 1659098407
transform 1 0 22540 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_245
timestamp 1659098407
transform 1 0 23644 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_251
timestamp 1659098407
transform 1 0 24196 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_253
timestamp 1659098407
transform 1 0 24380 0 1 14144
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_22_264
timestamp 1659098407
transform 1 0 25392 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_276
timestamp 1659098407
transform 1 0 26496 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_288
timestamp 1659098407
transform 1 0 27600 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_300
timestamp 1659098407
transform 1 0 28704 0 1 14144
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_22_309
timestamp 1659098407
transform 1 0 29532 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_321
timestamp 1659098407
transform 1 0 30636 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_333
timestamp 1659098407
transform 1 0 31740 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_345
timestamp 1659098407
transform 1 0 32844 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_357
timestamp 1659098407
transform 1 0 33948 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_363
timestamp 1659098407
transform 1 0 34500 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_365
timestamp 1659098407
transform 1 0 34684 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_377
timestamp 1659098407
transform 1 0 35788 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_389
timestamp 1659098407
transform 1 0 36892 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_401
timestamp 1659098407
transform 1 0 37996 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_22_413
timestamp 1659098407
transform 1 0 39100 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_419
timestamp 1659098407
transform 1 0 39652 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_441
timestamp 1659098407
transform 1 0 41676 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_449
timestamp 1659098407
transform 1 0 42412 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_22_459
timestamp 1659098407
transform 1 0 43332 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_471
timestamp 1659098407
transform 1 0 44436 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_475
timestamp 1659098407
transform 1 0 44804 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_477
timestamp 1659098407
transform 1 0 44988 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_489
timestamp 1659098407
transform 1 0 46092 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_501
timestamp 1659098407
transform 1 0 47196 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_22_512
timestamp 1659098407
transform 1 0 48208 0 1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_23_3
timestamp 1659098407
transform 1 0 1380 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_15
timestamp 1659098407
transform 1 0 2484 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_27
timestamp 1659098407
transform 1 0 3588 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_39
timestamp 1659098407
transform 1 0 4692 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_51
timestamp 1659098407
transform 1 0 5796 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_55
timestamp 1659098407
transform 1 0 6164 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_57
timestamp 1659098407
transform 1 0 6348 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_69
timestamp 1659098407
transform 1 0 7452 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_81
timestamp 1659098407
transform 1 0 8556 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_93
timestamp 1659098407
transform 1 0 9660 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_105
timestamp 1659098407
transform 1 0 10764 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_111
timestamp 1659098407
transform 1 0 11316 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_113
timestamp 1659098407
transform 1 0 11500 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_125
timestamp 1659098407
transform 1 0 12604 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_137
timestamp 1659098407
transform 1 0 13708 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_149
timestamp 1659098407
transform 1 0 14812 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_161
timestamp 1659098407
transform 1 0 15916 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_167
timestamp 1659098407
transform 1 0 16468 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_169
timestamp 1659098407
transform 1 0 16652 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_181
timestamp 1659098407
transform 1 0 17756 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_193
timestamp 1659098407
transform 1 0 18860 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_205
timestamp 1659098407
transform 1 0 19964 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_217
timestamp 1659098407
transform 1 0 21068 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_223
timestamp 1659098407
transform 1 0 21620 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_225
timestamp 1659098407
transform 1 0 21804 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_233
timestamp 1659098407
transform 1 0 22540 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_23_238
timestamp 1659098407
transform 1 0 23000 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_250
timestamp 1659098407
transform 1 0 24104 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_262
timestamp 1659098407
transform 1 0 25208 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_274
timestamp 1659098407
transform 1 0 26312 0 -1 15232
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_23_281
timestamp 1659098407
transform 1 0 26956 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_293
timestamp 1659098407
transform 1 0 28060 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_305
timestamp 1659098407
transform 1 0 29164 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_317
timestamp 1659098407
transform 1 0 30268 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_329
timestamp 1659098407
transform 1 0 31372 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_335
timestamp 1659098407
transform 1 0 31924 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_337
timestamp 1659098407
transform 1 0 32108 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_349
timestamp 1659098407
transform 1 0 33212 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_361
timestamp 1659098407
transform 1 0 34316 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_373
timestamp 1659098407
transform 1 0 35420 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_385
timestamp 1659098407
transform 1 0 36524 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_391
timestamp 1659098407
transform 1 0 37076 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_393
timestamp 1659098407
transform 1 0 37260 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_405
timestamp 1659098407
transform 1 0 38364 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_417
timestamp 1659098407
transform 1 0 39468 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_429
timestamp 1659098407
transform 1 0 40572 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_441
timestamp 1659098407
transform 1 0 41676 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_447
timestamp 1659098407
transform 1 0 42228 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_449
timestamp 1659098407
transform 1 0 42412 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_461
timestamp 1659098407
transform 1 0 43516 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_473
timestamp 1659098407
transform 1 0 44620 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_485
timestamp 1659098407
transform 1 0 45724 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_497
timestamp 1659098407
transform 1 0 46828 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_503
timestamp 1659098407
transform 1 0 47380 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_505
timestamp 1659098407
transform 1 0 47564 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_23_513
timestamp 1659098407
transform 1 0 48300 0 -1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_24_6
timestamp 1659098407
transform 1 0 1656 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_18
timestamp 1659098407
transform 1 0 2760 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_26
timestamp 1659098407
transform 1 0 3496 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_24_29
timestamp 1659098407
transform 1 0 3772 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_41
timestamp 1659098407
transform 1 0 4876 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_53
timestamp 1659098407
transform 1 0 5980 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_65
timestamp 1659098407
transform 1 0 7084 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_77
timestamp 1659098407
transform 1 0 8188 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_83
timestamp 1659098407
transform 1 0 8740 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_85
timestamp 1659098407
transform 1 0 8924 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_97
timestamp 1659098407
transform 1 0 10028 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_109
timestamp 1659098407
transform 1 0 11132 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_121
timestamp 1659098407
transform 1 0 12236 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_133
timestamp 1659098407
transform 1 0 13340 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_139
timestamp 1659098407
transform 1 0 13892 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_141
timestamp 1659098407
transform 1 0 14076 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_153
timestamp 1659098407
transform 1 0 15180 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_165
timestamp 1659098407
transform 1 0 16284 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_177
timestamp 1659098407
transform 1 0 17388 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_189
timestamp 1659098407
transform 1 0 18492 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_195
timestamp 1659098407
transform 1 0 19044 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_197
timestamp 1659098407
transform 1 0 19228 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_209
timestamp 1659098407
transform 1 0 20332 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_221
timestamp 1659098407
transform 1 0 21436 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_233
timestamp 1659098407
transform 1 0 22540 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_245
timestamp 1659098407
transform 1 0 23644 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_251
timestamp 1659098407
transform 1 0 24196 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_253
timestamp 1659098407
transform 1 0 24380 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_265
timestamp 1659098407
transform 1 0 25484 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_277
timestamp 1659098407
transform 1 0 26588 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_289
timestamp 1659098407
transform 1 0 27692 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_301
timestamp 1659098407
transform 1 0 28796 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_307
timestamp 1659098407
transform 1 0 29348 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_309
timestamp 1659098407
transform 1 0 29532 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_321
timestamp 1659098407
transform 1 0 30636 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_333
timestamp 1659098407
transform 1 0 31740 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_345
timestamp 1659098407
transform 1 0 32844 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_357
timestamp 1659098407
transform 1 0 33948 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_363
timestamp 1659098407
transform 1 0 34500 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_365
timestamp 1659098407
transform 1 0 34684 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_377
timestamp 1659098407
transform 1 0 35788 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_389
timestamp 1659098407
transform 1 0 36892 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_401
timestamp 1659098407
transform 1 0 37996 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_413
timestamp 1659098407
transform 1 0 39100 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_419
timestamp 1659098407
transform 1 0 39652 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_421
timestamp 1659098407
transform 1 0 39836 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_433
timestamp 1659098407
transform 1 0 40940 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_445
timestamp 1659098407
transform 1 0 42044 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_457
timestamp 1659098407
transform 1 0 43148 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_469
timestamp 1659098407
transform 1 0 44252 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_475
timestamp 1659098407
transform 1 0 44804 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_477
timestamp 1659098407
transform 1 0 44988 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_489
timestamp 1659098407
transform 1 0 46092 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_501
timestamp 1659098407
transform 1 0 47196 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_24_513
timestamp 1659098407
transform 1 0 48300 0 1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_25_6
timestamp 1659098407
transform 1 0 1656 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_18
timestamp 1659098407
transform 1 0 2760 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_30
timestamp 1659098407
transform 1 0 3864 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_42
timestamp 1659098407
transform 1 0 4968 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_25_54
timestamp 1659098407
transform 1 0 6072 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_25_57
timestamp 1659098407
transform 1 0 6348 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_69
timestamp 1659098407
transform 1 0 7452 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_81
timestamp 1659098407
transform 1 0 8556 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_93
timestamp 1659098407
transform 1 0 9660 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_105
timestamp 1659098407
transform 1 0 10764 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_111
timestamp 1659098407
transform 1 0 11316 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_113
timestamp 1659098407
transform 1 0 11500 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_125
timestamp 1659098407
transform 1 0 12604 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_137
timestamp 1659098407
transform 1 0 13708 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_149
timestamp 1659098407
transform 1 0 14812 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_161
timestamp 1659098407
transform 1 0 15916 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_167
timestamp 1659098407
transform 1 0 16468 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_169
timestamp 1659098407
transform 1 0 16652 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_181
timestamp 1659098407
transform 1 0 17756 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_193
timestamp 1659098407
transform 1 0 18860 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_205
timestamp 1659098407
transform 1 0 19964 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_217
timestamp 1659098407
transform 1 0 21068 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_223
timestamp 1659098407
transform 1 0 21620 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_225
timestamp 1659098407
transform 1 0 21804 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_237
timestamp 1659098407
transform 1 0 22908 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_249
timestamp 1659098407
transform 1 0 24012 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_261
timestamp 1659098407
transform 1 0 25116 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_273
timestamp 1659098407
transform 1 0 26220 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_279
timestamp 1659098407
transform 1 0 26772 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_281
timestamp 1659098407
transform 1 0 26956 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_293
timestamp 1659098407
transform 1 0 28060 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_305
timestamp 1659098407
transform 1 0 29164 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_317
timestamp 1659098407
transform 1 0 30268 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_329
timestamp 1659098407
transform 1 0 31372 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_335
timestamp 1659098407
transform 1 0 31924 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_337
timestamp 1659098407
transform 1 0 32108 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_349
timestamp 1659098407
transform 1 0 33212 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_361
timestamp 1659098407
transform 1 0 34316 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_373
timestamp 1659098407
transform 1 0 35420 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_385
timestamp 1659098407
transform 1 0 36524 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_391
timestamp 1659098407
transform 1 0 37076 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_393
timestamp 1659098407
transform 1 0 37260 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_405
timestamp 1659098407
transform 1 0 38364 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_417
timestamp 1659098407
transform 1 0 39468 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_429
timestamp 1659098407
transform 1 0 40572 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_441
timestamp 1659098407
transform 1 0 41676 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_447
timestamp 1659098407
transform 1 0 42228 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_449
timestamp 1659098407
transform 1 0 42412 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_461
timestamp 1659098407
transform 1 0 43516 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_473
timestamp 1659098407
transform 1 0 44620 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_485
timestamp 1659098407
transform 1 0 45724 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_497
timestamp 1659098407
transform 1 0 46828 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_503
timestamp 1659098407
transform 1 0 47380 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_505
timestamp 1659098407
transform 1 0 47564 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_512
timestamp 1659098407
transform 1 0 48208 0 -1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_26_3
timestamp 1659098407
transform 1 0 1380 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_15
timestamp 1659098407
transform 1 0 2484 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_27
timestamp 1659098407
transform 1 0 3588 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_29
timestamp 1659098407
transform 1 0 3772 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_41
timestamp 1659098407
transform 1 0 4876 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_53
timestamp 1659098407
transform 1 0 5980 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_65
timestamp 1659098407
transform 1 0 7084 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_77
timestamp 1659098407
transform 1 0 8188 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_83
timestamp 1659098407
transform 1 0 8740 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_85
timestamp 1659098407
transform 1 0 8924 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_97
timestamp 1659098407
transform 1 0 10028 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_109
timestamp 1659098407
transform 1 0 11132 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_121
timestamp 1659098407
transform 1 0 12236 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_133
timestamp 1659098407
transform 1 0 13340 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_139
timestamp 1659098407
transform 1 0 13892 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_141
timestamp 1659098407
transform 1 0 14076 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_153
timestamp 1659098407
transform 1 0 15180 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_165
timestamp 1659098407
transform 1 0 16284 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_177
timestamp 1659098407
transform 1 0 17388 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_189
timestamp 1659098407
transform 1 0 18492 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_195
timestamp 1659098407
transform 1 0 19044 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_197
timestamp 1659098407
transform 1 0 19228 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_209
timestamp 1659098407
transform 1 0 20332 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_221
timestamp 1659098407
transform 1 0 21436 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_233
timestamp 1659098407
transform 1 0 22540 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_245
timestamp 1659098407
transform 1 0 23644 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_251
timestamp 1659098407
transform 1 0 24196 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_253
timestamp 1659098407
transform 1 0 24380 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_265
timestamp 1659098407
transform 1 0 25484 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_277
timestamp 1659098407
transform 1 0 26588 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_289
timestamp 1659098407
transform 1 0 27692 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_301
timestamp 1659098407
transform 1 0 28796 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_307
timestamp 1659098407
transform 1 0 29348 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_309
timestamp 1659098407
transform 1 0 29532 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_321
timestamp 1659098407
transform 1 0 30636 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_333
timestamp 1659098407
transform 1 0 31740 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_345
timestamp 1659098407
transform 1 0 32844 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_357
timestamp 1659098407
transform 1 0 33948 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_363
timestamp 1659098407
transform 1 0 34500 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_365
timestamp 1659098407
transform 1 0 34684 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_377
timestamp 1659098407
transform 1 0 35788 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_389
timestamp 1659098407
transform 1 0 36892 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_401
timestamp 1659098407
transform 1 0 37996 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_413
timestamp 1659098407
transform 1 0 39100 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_419
timestamp 1659098407
transform 1 0 39652 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_421
timestamp 1659098407
transform 1 0 39836 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_433
timestamp 1659098407
transform 1 0 40940 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_445
timestamp 1659098407
transform 1 0 42044 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_457
timestamp 1659098407
transform 1 0 43148 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_469
timestamp 1659098407
transform 1 0 44252 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_475
timestamp 1659098407
transform 1 0 44804 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_477
timestamp 1659098407
transform 1 0 44988 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_489
timestamp 1659098407
transform 1 0 46092 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_501
timestamp 1659098407
transform 1 0 47196 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_26_512
timestamp 1659098407
transform 1 0 48208 0 1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_27_3
timestamp 1659098407
transform 1 0 1380 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_15
timestamp 1659098407
transform 1 0 2484 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_27
timestamp 1659098407
transform 1 0 3588 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_39
timestamp 1659098407
transform 1 0 4692 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_51
timestamp 1659098407
transform 1 0 5796 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_55
timestamp 1659098407
transform 1 0 6164 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_57
timestamp 1659098407
transform 1 0 6348 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_69
timestamp 1659098407
transform 1 0 7452 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_81
timestamp 1659098407
transform 1 0 8556 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_93
timestamp 1659098407
transform 1 0 9660 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_105
timestamp 1659098407
transform 1 0 10764 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_111
timestamp 1659098407
transform 1 0 11316 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_113
timestamp 1659098407
transform 1 0 11500 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_125
timestamp 1659098407
transform 1 0 12604 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_137
timestamp 1659098407
transform 1 0 13708 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_149
timestamp 1659098407
transform 1 0 14812 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_161
timestamp 1659098407
transform 1 0 15916 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_167
timestamp 1659098407
transform 1 0 16468 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_169
timestamp 1659098407
transform 1 0 16652 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_181
timestamp 1659098407
transform 1 0 17756 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_193
timestamp 1659098407
transform 1 0 18860 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_205
timestamp 1659098407
transform 1 0 19964 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_217
timestamp 1659098407
transform 1 0 21068 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_223
timestamp 1659098407
transform 1 0 21620 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_225
timestamp 1659098407
transform 1 0 21804 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_237
timestamp 1659098407
transform 1 0 22908 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_249
timestamp 1659098407
transform 1 0 24012 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_261
timestamp 1659098407
transform 1 0 25116 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_273
timestamp 1659098407
transform 1 0 26220 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_279
timestamp 1659098407
transform 1 0 26772 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_281
timestamp 1659098407
transform 1 0 26956 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_293
timestamp 1659098407
transform 1 0 28060 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_305
timestamp 1659098407
transform 1 0 29164 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_317
timestamp 1659098407
transform 1 0 30268 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_329
timestamp 1659098407
transform 1 0 31372 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_335
timestamp 1659098407
transform 1 0 31924 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_337
timestamp 1659098407
transform 1 0 32108 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_349
timestamp 1659098407
transform 1 0 33212 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_361
timestamp 1659098407
transform 1 0 34316 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_373
timestamp 1659098407
transform 1 0 35420 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_385
timestamp 1659098407
transform 1 0 36524 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_391
timestamp 1659098407
transform 1 0 37076 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_393
timestamp 1659098407
transform 1 0 37260 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_405
timestamp 1659098407
transform 1 0 38364 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_417
timestamp 1659098407
transform 1 0 39468 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_429
timestamp 1659098407
transform 1 0 40572 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_441
timestamp 1659098407
transform 1 0 41676 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_447
timestamp 1659098407
transform 1 0 42228 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_449
timestamp 1659098407
transform 1 0 42412 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_461
timestamp 1659098407
transform 1 0 43516 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_473
timestamp 1659098407
transform 1 0 44620 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_485
timestamp 1659098407
transform 1 0 45724 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_497
timestamp 1659098407
transform 1 0 46828 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_503
timestamp 1659098407
transform 1 0 47380 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_505
timestamp 1659098407
transform 1 0 47564 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_512
timestamp 1659098407
transform 1 0 48208 0 -1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_28_3
timestamp 1659098407
transform 1 0 1380 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_15
timestamp 1659098407
transform 1 0 2484 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_27
timestamp 1659098407
transform 1 0 3588 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_29
timestamp 1659098407
transform 1 0 3772 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_41
timestamp 1659098407
transform 1 0 4876 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_53
timestamp 1659098407
transform 1 0 5980 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_65
timestamp 1659098407
transform 1 0 7084 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_77
timestamp 1659098407
transform 1 0 8188 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_83
timestamp 1659098407
transform 1 0 8740 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_85
timestamp 1659098407
transform 1 0 8924 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_97
timestamp 1659098407
transform 1 0 10028 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_109
timestamp 1659098407
transform 1 0 11132 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_121
timestamp 1659098407
transform 1 0 12236 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_133
timestamp 1659098407
transform 1 0 13340 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_139
timestamp 1659098407
transform 1 0 13892 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_141
timestamp 1659098407
transform 1 0 14076 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_153
timestamp 1659098407
transform 1 0 15180 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_165
timestamp 1659098407
transform 1 0 16284 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_177
timestamp 1659098407
transform 1 0 17388 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_189
timestamp 1659098407
transform 1 0 18492 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_195
timestamp 1659098407
transform 1 0 19044 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_197
timestamp 1659098407
transform 1 0 19228 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_209
timestamp 1659098407
transform 1 0 20332 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_221
timestamp 1659098407
transform 1 0 21436 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_233
timestamp 1659098407
transform 1 0 22540 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_245
timestamp 1659098407
transform 1 0 23644 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_251
timestamp 1659098407
transform 1 0 24196 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_253
timestamp 1659098407
transform 1 0 24380 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_265
timestamp 1659098407
transform 1 0 25484 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_277
timestamp 1659098407
transform 1 0 26588 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_289
timestamp 1659098407
transform 1 0 27692 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_301
timestamp 1659098407
transform 1 0 28796 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_307
timestamp 1659098407
transform 1 0 29348 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_309
timestamp 1659098407
transform 1 0 29532 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_321
timestamp 1659098407
transform 1 0 30636 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_333
timestamp 1659098407
transform 1 0 31740 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_345
timestamp 1659098407
transform 1 0 32844 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_357
timestamp 1659098407
transform 1 0 33948 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_363
timestamp 1659098407
transform 1 0 34500 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_365
timestamp 1659098407
transform 1 0 34684 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_377
timestamp 1659098407
transform 1 0 35788 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_389
timestamp 1659098407
transform 1 0 36892 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_401
timestamp 1659098407
transform 1 0 37996 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_413
timestamp 1659098407
transform 1 0 39100 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_419
timestamp 1659098407
transform 1 0 39652 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_421
timestamp 1659098407
transform 1 0 39836 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_433
timestamp 1659098407
transform 1 0 40940 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_445
timestamp 1659098407
transform 1 0 42044 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_457
timestamp 1659098407
transform 1 0 43148 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_469
timestamp 1659098407
transform 1 0 44252 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_475
timestamp 1659098407
transform 1 0 44804 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_477
timestamp 1659098407
transform 1 0 44988 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_489
timestamp 1659098407
transform 1 0 46092 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_501
timestamp 1659098407
transform 1 0 47196 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_28_513
timestamp 1659098407
transform 1 0 48300 0 1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_29_3
timestamp 1659098407
transform 1 0 1380 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_15
timestamp 1659098407
transform 1 0 2484 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_27
timestamp 1659098407
transform 1 0 3588 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_39
timestamp 1659098407
transform 1 0 4692 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_51
timestamp 1659098407
transform 1 0 5796 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_55
timestamp 1659098407
transform 1 0 6164 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_57
timestamp 1659098407
transform 1 0 6348 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_69
timestamp 1659098407
transform 1 0 7452 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_81
timestamp 1659098407
transform 1 0 8556 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_93
timestamp 1659098407
transform 1 0 9660 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_105
timestamp 1659098407
transform 1 0 10764 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_111
timestamp 1659098407
transform 1 0 11316 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_113
timestamp 1659098407
transform 1 0 11500 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_125
timestamp 1659098407
transform 1 0 12604 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_137
timestamp 1659098407
transform 1 0 13708 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_149
timestamp 1659098407
transform 1 0 14812 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_161
timestamp 1659098407
transform 1 0 15916 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_167
timestamp 1659098407
transform 1 0 16468 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_169
timestamp 1659098407
transform 1 0 16652 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_181
timestamp 1659098407
transform 1 0 17756 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_193
timestamp 1659098407
transform 1 0 18860 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_205
timestamp 1659098407
transform 1 0 19964 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_217
timestamp 1659098407
transform 1 0 21068 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_223
timestamp 1659098407
transform 1 0 21620 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_225
timestamp 1659098407
transform 1 0 21804 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_237
timestamp 1659098407
transform 1 0 22908 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_249
timestamp 1659098407
transform 1 0 24012 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_261
timestamp 1659098407
transform 1 0 25116 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_273
timestamp 1659098407
transform 1 0 26220 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_279
timestamp 1659098407
transform 1 0 26772 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_281
timestamp 1659098407
transform 1 0 26956 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_293
timestamp 1659098407
transform 1 0 28060 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_305
timestamp 1659098407
transform 1 0 29164 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_317
timestamp 1659098407
transform 1 0 30268 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_329
timestamp 1659098407
transform 1 0 31372 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_335
timestamp 1659098407
transform 1 0 31924 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_337
timestamp 1659098407
transform 1 0 32108 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_349
timestamp 1659098407
transform 1 0 33212 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_361
timestamp 1659098407
transform 1 0 34316 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_373
timestamp 1659098407
transform 1 0 35420 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_385
timestamp 1659098407
transform 1 0 36524 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_391
timestamp 1659098407
transform 1 0 37076 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_393
timestamp 1659098407
transform 1 0 37260 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_405
timestamp 1659098407
transform 1 0 38364 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_417
timestamp 1659098407
transform 1 0 39468 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_429
timestamp 1659098407
transform 1 0 40572 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_441
timestamp 1659098407
transform 1 0 41676 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_447
timestamp 1659098407
transform 1 0 42228 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_449
timestamp 1659098407
transform 1 0 42412 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_461
timestamp 1659098407
transform 1 0 43516 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_473
timestamp 1659098407
transform 1 0 44620 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_485
timestamp 1659098407
transform 1 0 45724 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_497
timestamp 1659098407
transform 1 0 46828 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_503
timestamp 1659098407
transform 1 0 47380 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_505
timestamp 1659098407
transform 1 0 47564 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_512
timestamp 1659098407
transform 1 0 48208 0 -1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_30_6
timestamp 1659098407
transform 1 0 1656 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_18
timestamp 1659098407
transform 1 0 2760 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_30_26
timestamp 1659098407
transform 1 0 3496 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_30_29
timestamp 1659098407
transform 1 0 3772 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_41
timestamp 1659098407
transform 1 0 4876 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_53
timestamp 1659098407
transform 1 0 5980 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_65
timestamp 1659098407
transform 1 0 7084 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_77
timestamp 1659098407
transform 1 0 8188 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_83
timestamp 1659098407
transform 1 0 8740 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_85
timestamp 1659098407
transform 1 0 8924 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_97
timestamp 1659098407
transform 1 0 10028 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_109
timestamp 1659098407
transform 1 0 11132 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_121
timestamp 1659098407
transform 1 0 12236 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_133
timestamp 1659098407
transform 1 0 13340 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_139
timestamp 1659098407
transform 1 0 13892 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_141
timestamp 1659098407
transform 1 0 14076 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_153
timestamp 1659098407
transform 1 0 15180 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_165
timestamp 1659098407
transform 1 0 16284 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_177
timestamp 1659098407
transform 1 0 17388 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_189
timestamp 1659098407
transform 1 0 18492 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_195
timestamp 1659098407
transform 1 0 19044 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_197
timestamp 1659098407
transform 1 0 19228 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_209
timestamp 1659098407
transform 1 0 20332 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_221
timestamp 1659098407
transform 1 0 21436 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_233
timestamp 1659098407
transform 1 0 22540 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_245
timestamp 1659098407
transform 1 0 23644 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_251
timestamp 1659098407
transform 1 0 24196 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_253
timestamp 1659098407
transform 1 0 24380 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_265
timestamp 1659098407
transform 1 0 25484 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_277
timestamp 1659098407
transform 1 0 26588 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_289
timestamp 1659098407
transform 1 0 27692 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_301
timestamp 1659098407
transform 1 0 28796 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_307
timestamp 1659098407
transform 1 0 29348 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_309
timestamp 1659098407
transform 1 0 29532 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_321
timestamp 1659098407
transform 1 0 30636 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_333
timestamp 1659098407
transform 1 0 31740 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_345
timestamp 1659098407
transform 1 0 32844 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_357
timestamp 1659098407
transform 1 0 33948 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_363
timestamp 1659098407
transform 1 0 34500 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_365
timestamp 1659098407
transform 1 0 34684 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_377
timestamp 1659098407
transform 1 0 35788 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_389
timestamp 1659098407
transform 1 0 36892 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_401
timestamp 1659098407
transform 1 0 37996 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_413
timestamp 1659098407
transform 1 0 39100 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_419
timestamp 1659098407
transform 1 0 39652 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_421
timestamp 1659098407
transform 1 0 39836 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_433
timestamp 1659098407
transform 1 0 40940 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_445
timestamp 1659098407
transform 1 0 42044 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_457
timestamp 1659098407
transform 1 0 43148 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_469
timestamp 1659098407
transform 1 0 44252 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_475
timestamp 1659098407
transform 1 0 44804 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_477
timestamp 1659098407
transform 1 0 44988 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_489
timestamp 1659098407
transform 1 0 46092 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_501
timestamp 1659098407
transform 1 0 47196 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_30_512
timestamp 1659098407
transform 1 0 48208 0 1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_31_6
timestamp 1659098407
transform 1 0 1656 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_18
timestamp 1659098407
transform 1 0 2760 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_30
timestamp 1659098407
transform 1 0 3864 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_42
timestamp 1659098407
transform 1 0 4968 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_31_54
timestamp 1659098407
transform 1 0 6072 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_31_57
timestamp 1659098407
transform 1 0 6348 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_69
timestamp 1659098407
transform 1 0 7452 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_81
timestamp 1659098407
transform 1 0 8556 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_93
timestamp 1659098407
transform 1 0 9660 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_105
timestamp 1659098407
transform 1 0 10764 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_111
timestamp 1659098407
transform 1 0 11316 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_113
timestamp 1659098407
transform 1 0 11500 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_125
timestamp 1659098407
transform 1 0 12604 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_137
timestamp 1659098407
transform 1 0 13708 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_149
timestamp 1659098407
transform 1 0 14812 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_161
timestamp 1659098407
transform 1 0 15916 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_167
timestamp 1659098407
transform 1 0 16468 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_169
timestamp 1659098407
transform 1 0 16652 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_181
timestamp 1659098407
transform 1 0 17756 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_193
timestamp 1659098407
transform 1 0 18860 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_205
timestamp 1659098407
transform 1 0 19964 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_217
timestamp 1659098407
transform 1 0 21068 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_223
timestamp 1659098407
transform 1 0 21620 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_225
timestamp 1659098407
transform 1 0 21804 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_237
timestamp 1659098407
transform 1 0 22908 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_249
timestamp 1659098407
transform 1 0 24012 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_261
timestamp 1659098407
transform 1 0 25116 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_273
timestamp 1659098407
transform 1 0 26220 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_279
timestamp 1659098407
transform 1 0 26772 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_281
timestamp 1659098407
transform 1 0 26956 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_293
timestamp 1659098407
transform 1 0 28060 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_305
timestamp 1659098407
transform 1 0 29164 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_317
timestamp 1659098407
transform 1 0 30268 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_329
timestamp 1659098407
transform 1 0 31372 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_335
timestamp 1659098407
transform 1 0 31924 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_337
timestamp 1659098407
transform 1 0 32108 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_349
timestamp 1659098407
transform 1 0 33212 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_361
timestamp 1659098407
transform 1 0 34316 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_373
timestamp 1659098407
transform 1 0 35420 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_385
timestamp 1659098407
transform 1 0 36524 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_391
timestamp 1659098407
transform 1 0 37076 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_393
timestamp 1659098407
transform 1 0 37260 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_405
timestamp 1659098407
transform 1 0 38364 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_417
timestamp 1659098407
transform 1 0 39468 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_429
timestamp 1659098407
transform 1 0 40572 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_441
timestamp 1659098407
transform 1 0 41676 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_447
timestamp 1659098407
transform 1 0 42228 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_449
timestamp 1659098407
transform 1 0 42412 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_461
timestamp 1659098407
transform 1 0 43516 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_473
timestamp 1659098407
transform 1 0 44620 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_485
timestamp 1659098407
transform 1 0 45724 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_497
timestamp 1659098407
transform 1 0 46828 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_503
timestamp 1659098407
transform 1 0 47380 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_505
timestamp 1659098407
transform 1 0 47564 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_512
timestamp 1659098407
transform 1 0 48208 0 -1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_32_6
timestamp 1659098407
transform 1 0 1656 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_18
timestamp 1659098407
transform 1 0 2760 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_32_26
timestamp 1659098407
transform 1 0 3496 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_32_29
timestamp 1659098407
transform 1 0 3772 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_41
timestamp 1659098407
transform 1 0 4876 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_53
timestamp 1659098407
transform 1 0 5980 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_65
timestamp 1659098407
transform 1 0 7084 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_77
timestamp 1659098407
transform 1 0 8188 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_83
timestamp 1659098407
transform 1 0 8740 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_85
timestamp 1659098407
transform 1 0 8924 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_97
timestamp 1659098407
transform 1 0 10028 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_109
timestamp 1659098407
transform 1 0 11132 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_121
timestamp 1659098407
transform 1 0 12236 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_133
timestamp 1659098407
transform 1 0 13340 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_139
timestamp 1659098407
transform 1 0 13892 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_141
timestamp 1659098407
transform 1 0 14076 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_153
timestamp 1659098407
transform 1 0 15180 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_165
timestamp 1659098407
transform 1 0 16284 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_177
timestamp 1659098407
transform 1 0 17388 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_189
timestamp 1659098407
transform 1 0 18492 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_195
timestamp 1659098407
transform 1 0 19044 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_197
timestamp 1659098407
transform 1 0 19228 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_209
timestamp 1659098407
transform 1 0 20332 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_221
timestamp 1659098407
transform 1 0 21436 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_233
timestamp 1659098407
transform 1 0 22540 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_245
timestamp 1659098407
transform 1 0 23644 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_251
timestamp 1659098407
transform 1 0 24196 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_253
timestamp 1659098407
transform 1 0 24380 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_265
timestamp 1659098407
transform 1 0 25484 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_277
timestamp 1659098407
transform 1 0 26588 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_289
timestamp 1659098407
transform 1 0 27692 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_301
timestamp 1659098407
transform 1 0 28796 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_307
timestamp 1659098407
transform 1 0 29348 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_309
timestamp 1659098407
transform 1 0 29532 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_321
timestamp 1659098407
transform 1 0 30636 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_333
timestamp 1659098407
transform 1 0 31740 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_345
timestamp 1659098407
transform 1 0 32844 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_357
timestamp 1659098407
transform 1 0 33948 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_363
timestamp 1659098407
transform 1 0 34500 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_365
timestamp 1659098407
transform 1 0 34684 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_377
timestamp 1659098407
transform 1 0 35788 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_389
timestamp 1659098407
transform 1 0 36892 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_401
timestamp 1659098407
transform 1 0 37996 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_413
timestamp 1659098407
transform 1 0 39100 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_419
timestamp 1659098407
transform 1 0 39652 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_421
timestamp 1659098407
transform 1 0 39836 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_433
timestamp 1659098407
transform 1 0 40940 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_445
timestamp 1659098407
transform 1 0 42044 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_457
timestamp 1659098407
transform 1 0 43148 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_469
timestamp 1659098407
transform 1 0 44252 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_475
timestamp 1659098407
transform 1 0 44804 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_477
timestamp 1659098407
transform 1 0 44988 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_489
timestamp 1659098407
transform 1 0 46092 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_501
timestamp 1659098407
transform 1 0 47196 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_32_513
timestamp 1659098407
transform 1 0 48300 0 1 19584
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_33_3
timestamp 1659098407
transform 1 0 1380 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_15
timestamp 1659098407
transform 1 0 2484 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_27
timestamp 1659098407
transform 1 0 3588 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_39
timestamp 1659098407
transform 1 0 4692 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_51
timestamp 1659098407
transform 1 0 5796 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_55
timestamp 1659098407
transform 1 0 6164 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_57
timestamp 1659098407
transform 1 0 6348 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_69
timestamp 1659098407
transform 1 0 7452 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_81
timestamp 1659098407
transform 1 0 8556 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_93
timestamp 1659098407
transform 1 0 9660 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_105
timestamp 1659098407
transform 1 0 10764 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_111
timestamp 1659098407
transform 1 0 11316 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_113
timestamp 1659098407
transform 1 0 11500 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_125
timestamp 1659098407
transform 1 0 12604 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_137
timestamp 1659098407
transform 1 0 13708 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_149
timestamp 1659098407
transform 1 0 14812 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_161
timestamp 1659098407
transform 1 0 15916 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_167
timestamp 1659098407
transform 1 0 16468 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_169
timestamp 1659098407
transform 1 0 16652 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_181
timestamp 1659098407
transform 1 0 17756 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_193
timestamp 1659098407
transform 1 0 18860 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_205
timestamp 1659098407
transform 1 0 19964 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_217
timestamp 1659098407
transform 1 0 21068 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_223
timestamp 1659098407
transform 1 0 21620 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_225
timestamp 1659098407
transform 1 0 21804 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_237
timestamp 1659098407
transform 1 0 22908 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_249
timestamp 1659098407
transform 1 0 24012 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_261
timestamp 1659098407
transform 1 0 25116 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_273
timestamp 1659098407
transform 1 0 26220 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_279
timestamp 1659098407
transform 1 0 26772 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_281
timestamp 1659098407
transform 1 0 26956 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_293
timestamp 1659098407
transform 1 0 28060 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_305
timestamp 1659098407
transform 1 0 29164 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_317
timestamp 1659098407
transform 1 0 30268 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_329
timestamp 1659098407
transform 1 0 31372 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_335
timestamp 1659098407
transform 1 0 31924 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_337
timestamp 1659098407
transform 1 0 32108 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_349
timestamp 1659098407
transform 1 0 33212 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_361
timestamp 1659098407
transform 1 0 34316 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_373
timestamp 1659098407
transform 1 0 35420 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_385
timestamp 1659098407
transform 1 0 36524 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_391
timestamp 1659098407
transform 1 0 37076 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_393
timestamp 1659098407
transform 1 0 37260 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_405
timestamp 1659098407
transform 1 0 38364 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_417
timestamp 1659098407
transform 1 0 39468 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_429
timestamp 1659098407
transform 1 0 40572 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_441
timestamp 1659098407
transform 1 0 41676 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_447
timestamp 1659098407
transform 1 0 42228 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_449
timestamp 1659098407
transform 1 0 42412 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_461
timestamp 1659098407
transform 1 0 43516 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_473
timestamp 1659098407
transform 1 0 44620 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_485
timestamp 1659098407
transform 1 0 45724 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_497
timestamp 1659098407
transform 1 0 46828 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_503
timestamp 1659098407
transform 1 0 47380 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_505
timestamp 1659098407
transform 1 0 47564 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_33_513
timestamp 1659098407
transform 1 0 48300 0 -1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_34_6
timestamp 1659098407
transform 1 0 1656 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_18
timestamp 1659098407
transform 1 0 2760 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_34_26
timestamp 1659098407
transform 1 0 3496 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_34_29
timestamp 1659098407
transform 1 0 3772 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_41
timestamp 1659098407
transform 1 0 4876 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_53
timestamp 1659098407
transform 1 0 5980 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_65
timestamp 1659098407
transform 1 0 7084 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_77
timestamp 1659098407
transform 1 0 8188 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_83
timestamp 1659098407
transform 1 0 8740 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_85
timestamp 1659098407
transform 1 0 8924 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_97
timestamp 1659098407
transform 1 0 10028 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_109
timestamp 1659098407
transform 1 0 11132 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_121
timestamp 1659098407
transform 1 0 12236 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_133
timestamp 1659098407
transform 1 0 13340 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_139
timestamp 1659098407
transform 1 0 13892 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_141
timestamp 1659098407
transform 1 0 14076 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_153
timestamp 1659098407
transform 1 0 15180 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_165
timestamp 1659098407
transform 1 0 16284 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_177
timestamp 1659098407
transform 1 0 17388 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_189
timestamp 1659098407
transform 1 0 18492 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_195
timestamp 1659098407
transform 1 0 19044 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_197
timestamp 1659098407
transform 1 0 19228 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_209
timestamp 1659098407
transform 1 0 20332 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_221
timestamp 1659098407
transform 1 0 21436 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_233
timestamp 1659098407
transform 1 0 22540 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_245
timestamp 1659098407
transform 1 0 23644 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_251
timestamp 1659098407
transform 1 0 24196 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_253
timestamp 1659098407
transform 1 0 24380 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_265
timestamp 1659098407
transform 1 0 25484 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_277
timestamp 1659098407
transform 1 0 26588 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_289
timestamp 1659098407
transform 1 0 27692 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_301
timestamp 1659098407
transform 1 0 28796 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_307
timestamp 1659098407
transform 1 0 29348 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_309
timestamp 1659098407
transform 1 0 29532 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_321
timestamp 1659098407
transform 1 0 30636 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_333
timestamp 1659098407
transform 1 0 31740 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_345
timestamp 1659098407
transform 1 0 32844 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_357
timestamp 1659098407
transform 1 0 33948 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_363
timestamp 1659098407
transform 1 0 34500 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_365
timestamp 1659098407
transform 1 0 34684 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_377
timestamp 1659098407
transform 1 0 35788 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_389
timestamp 1659098407
transform 1 0 36892 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_401
timestamp 1659098407
transform 1 0 37996 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_413
timestamp 1659098407
transform 1 0 39100 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_419
timestamp 1659098407
transform 1 0 39652 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_421
timestamp 1659098407
transform 1 0 39836 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_433
timestamp 1659098407
transform 1 0 40940 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_445
timestamp 1659098407
transform 1 0 42044 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_457
timestamp 1659098407
transform 1 0 43148 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_469
timestamp 1659098407
transform 1 0 44252 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_475
timestamp 1659098407
transform 1 0 44804 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_477
timestamp 1659098407
transform 1 0 44988 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_489
timestamp 1659098407
transform 1 0 46092 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_501
timestamp 1659098407
transform 1 0 47196 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_34_512
timestamp 1659098407
transform 1 0 48208 0 1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_35_6
timestamp 1659098407
transform 1 0 1656 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_18
timestamp 1659098407
transform 1 0 2760 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_30
timestamp 1659098407
transform 1 0 3864 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_42
timestamp 1659098407
transform 1 0 4968 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_35_54
timestamp 1659098407
transform 1 0 6072 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_35_57
timestamp 1659098407
transform 1 0 6348 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_69
timestamp 1659098407
transform 1 0 7452 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_81
timestamp 1659098407
transform 1 0 8556 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_93
timestamp 1659098407
transform 1 0 9660 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_105
timestamp 1659098407
transform 1 0 10764 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_111
timestamp 1659098407
transform 1 0 11316 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_113
timestamp 1659098407
transform 1 0 11500 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_125
timestamp 1659098407
transform 1 0 12604 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_137
timestamp 1659098407
transform 1 0 13708 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_149
timestamp 1659098407
transform 1 0 14812 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_161
timestamp 1659098407
transform 1 0 15916 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_167
timestamp 1659098407
transform 1 0 16468 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_169
timestamp 1659098407
transform 1 0 16652 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_181
timestamp 1659098407
transform 1 0 17756 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_193
timestamp 1659098407
transform 1 0 18860 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_205
timestamp 1659098407
transform 1 0 19964 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_217
timestamp 1659098407
transform 1 0 21068 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_223
timestamp 1659098407
transform 1 0 21620 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_225
timestamp 1659098407
transform 1 0 21804 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_237
timestamp 1659098407
transform 1 0 22908 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_249
timestamp 1659098407
transform 1 0 24012 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_261
timestamp 1659098407
transform 1 0 25116 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_273
timestamp 1659098407
transform 1 0 26220 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_279
timestamp 1659098407
transform 1 0 26772 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_281
timestamp 1659098407
transform 1 0 26956 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_293
timestamp 1659098407
transform 1 0 28060 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_305
timestamp 1659098407
transform 1 0 29164 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_317
timestamp 1659098407
transform 1 0 30268 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_329
timestamp 1659098407
transform 1 0 31372 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_335
timestamp 1659098407
transform 1 0 31924 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_337
timestamp 1659098407
transform 1 0 32108 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_349
timestamp 1659098407
transform 1 0 33212 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_361
timestamp 1659098407
transform 1 0 34316 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_373
timestamp 1659098407
transform 1 0 35420 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_385
timestamp 1659098407
transform 1 0 36524 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_391
timestamp 1659098407
transform 1 0 37076 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_393
timestamp 1659098407
transform 1 0 37260 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_405
timestamp 1659098407
transform 1 0 38364 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_417
timestamp 1659098407
transform 1 0 39468 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_429
timestamp 1659098407
transform 1 0 40572 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_441
timestamp 1659098407
transform 1 0 41676 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_447
timestamp 1659098407
transform 1 0 42228 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_449
timestamp 1659098407
transform 1 0 42412 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_461
timestamp 1659098407
transform 1 0 43516 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_473
timestamp 1659098407
transform 1 0 44620 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_485
timestamp 1659098407
transform 1 0 45724 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_497
timestamp 1659098407
transform 1 0 46828 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_503
timestamp 1659098407
transform 1 0 47380 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_35_505
timestamp 1659098407
transform 1 0 47564 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_35_513
timestamp 1659098407
transform 1 0 48300 0 -1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_36_6
timestamp 1659098407
transform 1 0 1656 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_36_18
timestamp 1659098407
transform 1 0 2760 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_36_26
timestamp 1659098407
transform 1 0 3496 0 1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_36_29
timestamp 1659098407
transform 1 0 3772 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_41
timestamp 1659098407
transform 1 0 4876 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_53
timestamp 1659098407
transform 1 0 5980 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_65
timestamp 1659098407
transform 1 0 7084 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_77
timestamp 1659098407
transform 1 0 8188 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_83
timestamp 1659098407
transform 1 0 8740 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_85
timestamp 1659098407
transform 1 0 8924 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_97
timestamp 1659098407
transform 1 0 10028 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_109
timestamp 1659098407
transform 1 0 11132 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_121
timestamp 1659098407
transform 1 0 12236 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_133
timestamp 1659098407
transform 1 0 13340 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_139
timestamp 1659098407
transform 1 0 13892 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_141
timestamp 1659098407
transform 1 0 14076 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_153
timestamp 1659098407
transform 1 0 15180 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_165
timestamp 1659098407
transform 1 0 16284 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_177
timestamp 1659098407
transform 1 0 17388 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_189
timestamp 1659098407
transform 1 0 18492 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_195
timestamp 1659098407
transform 1 0 19044 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_197
timestamp 1659098407
transform 1 0 19228 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_209
timestamp 1659098407
transform 1 0 20332 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_221
timestamp 1659098407
transform 1 0 21436 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_233
timestamp 1659098407
transform 1 0 22540 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_245
timestamp 1659098407
transform 1 0 23644 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_251
timestamp 1659098407
transform 1 0 24196 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_253
timestamp 1659098407
transform 1 0 24380 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_265
timestamp 1659098407
transform 1 0 25484 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_277
timestamp 1659098407
transform 1 0 26588 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_289
timestamp 1659098407
transform 1 0 27692 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_301
timestamp 1659098407
transform 1 0 28796 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_307
timestamp 1659098407
transform 1 0 29348 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_309
timestamp 1659098407
transform 1 0 29532 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_321
timestamp 1659098407
transform 1 0 30636 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_333
timestamp 1659098407
transform 1 0 31740 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_345
timestamp 1659098407
transform 1 0 32844 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_357
timestamp 1659098407
transform 1 0 33948 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_363
timestamp 1659098407
transform 1 0 34500 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_365
timestamp 1659098407
transform 1 0 34684 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_377
timestamp 1659098407
transform 1 0 35788 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_389
timestamp 1659098407
transform 1 0 36892 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_401
timestamp 1659098407
transform 1 0 37996 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_413
timestamp 1659098407
transform 1 0 39100 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_419
timestamp 1659098407
transform 1 0 39652 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_421
timestamp 1659098407
transform 1 0 39836 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_433
timestamp 1659098407
transform 1 0 40940 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_445
timestamp 1659098407
transform 1 0 42044 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_457
timestamp 1659098407
transform 1 0 43148 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_469
timestamp 1659098407
transform 1 0 44252 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_475
timestamp 1659098407
transform 1 0 44804 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_477
timestamp 1659098407
transform 1 0 44988 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_489
timestamp 1659098407
transform 1 0 46092 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_36_501
timestamp 1659098407
transform 1 0 47196 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_36_512
timestamp 1659098407
transform 1 0 48208 0 1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_37_3
timestamp 1659098407
transform 1 0 1380 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_15
timestamp 1659098407
transform 1 0 2484 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_27
timestamp 1659098407
transform 1 0 3588 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_39
timestamp 1659098407
transform 1 0 4692 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_51
timestamp 1659098407
transform 1 0 5796 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_55
timestamp 1659098407
transform 1 0 6164 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_57
timestamp 1659098407
transform 1 0 6348 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_69
timestamp 1659098407
transform 1 0 7452 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_81
timestamp 1659098407
transform 1 0 8556 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_93
timestamp 1659098407
transform 1 0 9660 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_105
timestamp 1659098407
transform 1 0 10764 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_111
timestamp 1659098407
transform 1 0 11316 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_113
timestamp 1659098407
transform 1 0 11500 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_125
timestamp 1659098407
transform 1 0 12604 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_137
timestamp 1659098407
transform 1 0 13708 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_149
timestamp 1659098407
transform 1 0 14812 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_161
timestamp 1659098407
transform 1 0 15916 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_167
timestamp 1659098407
transform 1 0 16468 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_169
timestamp 1659098407
transform 1 0 16652 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_181
timestamp 1659098407
transform 1 0 17756 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_193
timestamp 1659098407
transform 1 0 18860 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_205
timestamp 1659098407
transform 1 0 19964 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_217
timestamp 1659098407
transform 1 0 21068 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_223
timestamp 1659098407
transform 1 0 21620 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_225
timestamp 1659098407
transform 1 0 21804 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_237
timestamp 1659098407
transform 1 0 22908 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_249
timestamp 1659098407
transform 1 0 24012 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_261
timestamp 1659098407
transform 1 0 25116 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_273
timestamp 1659098407
transform 1 0 26220 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_279
timestamp 1659098407
transform 1 0 26772 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_281
timestamp 1659098407
transform 1 0 26956 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_293
timestamp 1659098407
transform 1 0 28060 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_305
timestamp 1659098407
transform 1 0 29164 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_317
timestamp 1659098407
transform 1 0 30268 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_329
timestamp 1659098407
transform 1 0 31372 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_335
timestamp 1659098407
transform 1 0 31924 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_337
timestamp 1659098407
transform 1 0 32108 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_349
timestamp 1659098407
transform 1 0 33212 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_361
timestamp 1659098407
transform 1 0 34316 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_373
timestamp 1659098407
transform 1 0 35420 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_385
timestamp 1659098407
transform 1 0 36524 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_391
timestamp 1659098407
transform 1 0 37076 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_393
timestamp 1659098407
transform 1 0 37260 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_405
timestamp 1659098407
transform 1 0 38364 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_417
timestamp 1659098407
transform 1 0 39468 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_429
timestamp 1659098407
transform 1 0 40572 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_441
timestamp 1659098407
transform 1 0 41676 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_447
timestamp 1659098407
transform 1 0 42228 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_449
timestamp 1659098407
transform 1 0 42412 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_461
timestamp 1659098407
transform 1 0 43516 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_473
timestamp 1659098407
transform 1 0 44620 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_485
timestamp 1659098407
transform 1 0 45724 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_497
timestamp 1659098407
transform 1 0 46828 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_503
timestamp 1659098407
transform 1 0 47380 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_505
timestamp 1659098407
transform 1 0 47564 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_512
timestamp 1659098407
transform 1 0 48208 0 -1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_38_3
timestamp 1659098407
transform 1 0 1380 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_15
timestamp 1659098407
transform 1 0 2484 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_38_27
timestamp 1659098407
transform 1 0 3588 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_29
timestamp 1659098407
transform 1 0 3772 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_41
timestamp 1659098407
transform 1 0 4876 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_53
timestamp 1659098407
transform 1 0 5980 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_65
timestamp 1659098407
transform 1 0 7084 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_77
timestamp 1659098407
transform 1 0 8188 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_83
timestamp 1659098407
transform 1 0 8740 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_85
timestamp 1659098407
transform 1 0 8924 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_97
timestamp 1659098407
transform 1 0 10028 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_109
timestamp 1659098407
transform 1 0 11132 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_121
timestamp 1659098407
transform 1 0 12236 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_133
timestamp 1659098407
transform 1 0 13340 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_139
timestamp 1659098407
transform 1 0 13892 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_141
timestamp 1659098407
transform 1 0 14076 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_153
timestamp 1659098407
transform 1 0 15180 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_165
timestamp 1659098407
transform 1 0 16284 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_177
timestamp 1659098407
transform 1 0 17388 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_189
timestamp 1659098407
transform 1 0 18492 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_195
timestamp 1659098407
transform 1 0 19044 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_197
timestamp 1659098407
transform 1 0 19228 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_209
timestamp 1659098407
transform 1 0 20332 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_221
timestamp 1659098407
transform 1 0 21436 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_233
timestamp 1659098407
transform 1 0 22540 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_245
timestamp 1659098407
transform 1 0 23644 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_251
timestamp 1659098407
transform 1 0 24196 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_253
timestamp 1659098407
transform 1 0 24380 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_265
timestamp 1659098407
transform 1 0 25484 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_277
timestamp 1659098407
transform 1 0 26588 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_289
timestamp 1659098407
transform 1 0 27692 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_301
timestamp 1659098407
transform 1 0 28796 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_307
timestamp 1659098407
transform 1 0 29348 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_309
timestamp 1659098407
transform 1 0 29532 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_321
timestamp 1659098407
transform 1 0 30636 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_333
timestamp 1659098407
transform 1 0 31740 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_345
timestamp 1659098407
transform 1 0 32844 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_357
timestamp 1659098407
transform 1 0 33948 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_363
timestamp 1659098407
transform 1 0 34500 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_365
timestamp 1659098407
transform 1 0 34684 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_377
timestamp 1659098407
transform 1 0 35788 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_389
timestamp 1659098407
transform 1 0 36892 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_401
timestamp 1659098407
transform 1 0 37996 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_413
timestamp 1659098407
transform 1 0 39100 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_419
timestamp 1659098407
transform 1 0 39652 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_421
timestamp 1659098407
transform 1 0 39836 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_433
timestamp 1659098407
transform 1 0 40940 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_445
timestamp 1659098407
transform 1 0 42044 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_457
timestamp 1659098407
transform 1 0 43148 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_469
timestamp 1659098407
transform 1 0 44252 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_475
timestamp 1659098407
transform 1 0 44804 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_477
timestamp 1659098407
transform 1 0 44988 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_489
timestamp 1659098407
transform 1 0 46092 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_501
timestamp 1659098407
transform 1 0 47196 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_38_513
timestamp 1659098407
transform 1 0 48300 0 1 22848
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_39_6
timestamp 1659098407
transform 1 0 1656 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_18
timestamp 1659098407
transform 1 0 2760 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_30
timestamp 1659098407
transform 1 0 3864 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_42
timestamp 1659098407
transform 1 0 4968 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_39_54
timestamp 1659098407
transform 1 0 6072 0 -1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_39_57
timestamp 1659098407
transform 1 0 6348 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_69
timestamp 1659098407
transform 1 0 7452 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_81
timestamp 1659098407
transform 1 0 8556 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_93
timestamp 1659098407
transform 1 0 9660 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_105
timestamp 1659098407
transform 1 0 10764 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_111
timestamp 1659098407
transform 1 0 11316 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_113
timestamp 1659098407
transform 1 0 11500 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_125
timestamp 1659098407
transform 1 0 12604 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_137
timestamp 1659098407
transform 1 0 13708 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_149
timestamp 1659098407
transform 1 0 14812 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_161
timestamp 1659098407
transform 1 0 15916 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_167
timestamp 1659098407
transform 1 0 16468 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_169
timestamp 1659098407
transform 1 0 16652 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_181
timestamp 1659098407
transform 1 0 17756 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_193
timestamp 1659098407
transform 1 0 18860 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_205
timestamp 1659098407
transform 1 0 19964 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_217
timestamp 1659098407
transform 1 0 21068 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_223
timestamp 1659098407
transform 1 0 21620 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_225
timestamp 1659098407
transform 1 0 21804 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_237
timestamp 1659098407
transform 1 0 22908 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_249
timestamp 1659098407
transform 1 0 24012 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_261
timestamp 1659098407
transform 1 0 25116 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_273
timestamp 1659098407
transform 1 0 26220 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_279
timestamp 1659098407
transform 1 0 26772 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_281
timestamp 1659098407
transform 1 0 26956 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_293
timestamp 1659098407
transform 1 0 28060 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_305
timestamp 1659098407
transform 1 0 29164 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_317
timestamp 1659098407
transform 1 0 30268 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_329
timestamp 1659098407
transform 1 0 31372 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_335
timestamp 1659098407
transform 1 0 31924 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_337
timestamp 1659098407
transform 1 0 32108 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_349
timestamp 1659098407
transform 1 0 33212 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_361
timestamp 1659098407
transform 1 0 34316 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_373
timestamp 1659098407
transform 1 0 35420 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_385
timestamp 1659098407
transform 1 0 36524 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_391
timestamp 1659098407
transform 1 0 37076 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_393
timestamp 1659098407
transform 1 0 37260 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_405
timestamp 1659098407
transform 1 0 38364 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_417
timestamp 1659098407
transform 1 0 39468 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_429
timestamp 1659098407
transform 1 0 40572 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_441
timestamp 1659098407
transform 1 0 41676 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_447
timestamp 1659098407
transform 1 0 42228 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_449
timestamp 1659098407
transform 1 0 42412 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_461
timestamp 1659098407
transform 1 0 43516 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_473
timestamp 1659098407
transform 1 0 44620 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_485
timestamp 1659098407
transform 1 0 45724 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_497
timestamp 1659098407
transform 1 0 46828 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_503
timestamp 1659098407
transform 1 0 47380 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_505
timestamp 1659098407
transform 1 0 47564 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_512
timestamp 1659098407
transform 1 0 48208 0 -1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_40_6
timestamp 1659098407
transform 1 0 1656 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_18
timestamp 1659098407
transform 1 0 2760 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_40_26
timestamp 1659098407
transform 1 0 3496 0 1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_40_29
timestamp 1659098407
transform 1 0 3772 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_41
timestamp 1659098407
transform 1 0 4876 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_53
timestamp 1659098407
transform 1 0 5980 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_65
timestamp 1659098407
transform 1 0 7084 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_77
timestamp 1659098407
transform 1 0 8188 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_83
timestamp 1659098407
transform 1 0 8740 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_85
timestamp 1659098407
transform 1 0 8924 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_97
timestamp 1659098407
transform 1 0 10028 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_109
timestamp 1659098407
transform 1 0 11132 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_121
timestamp 1659098407
transform 1 0 12236 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_133
timestamp 1659098407
transform 1 0 13340 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_139
timestamp 1659098407
transform 1 0 13892 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_141
timestamp 1659098407
transform 1 0 14076 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_153
timestamp 1659098407
transform 1 0 15180 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_165
timestamp 1659098407
transform 1 0 16284 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_177
timestamp 1659098407
transform 1 0 17388 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_189
timestamp 1659098407
transform 1 0 18492 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_195
timestamp 1659098407
transform 1 0 19044 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_197
timestamp 1659098407
transform 1 0 19228 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_209
timestamp 1659098407
transform 1 0 20332 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_221
timestamp 1659098407
transform 1 0 21436 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_233
timestamp 1659098407
transform 1 0 22540 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_245
timestamp 1659098407
transform 1 0 23644 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_251
timestamp 1659098407
transform 1 0 24196 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_253
timestamp 1659098407
transform 1 0 24380 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_265
timestamp 1659098407
transform 1 0 25484 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_277
timestamp 1659098407
transform 1 0 26588 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_289
timestamp 1659098407
transform 1 0 27692 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_301
timestamp 1659098407
transform 1 0 28796 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_307
timestamp 1659098407
transform 1 0 29348 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_309
timestamp 1659098407
transform 1 0 29532 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_321
timestamp 1659098407
transform 1 0 30636 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_333
timestamp 1659098407
transform 1 0 31740 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_345
timestamp 1659098407
transform 1 0 32844 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_357
timestamp 1659098407
transform 1 0 33948 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_363
timestamp 1659098407
transform 1 0 34500 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_365
timestamp 1659098407
transform 1 0 34684 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_377
timestamp 1659098407
transform 1 0 35788 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_389
timestamp 1659098407
transform 1 0 36892 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_401
timestamp 1659098407
transform 1 0 37996 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_413
timestamp 1659098407
transform 1 0 39100 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_419
timestamp 1659098407
transform 1 0 39652 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_421
timestamp 1659098407
transform 1 0 39836 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_433
timestamp 1659098407
transform 1 0 40940 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_445
timestamp 1659098407
transform 1 0 42044 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_457
timestamp 1659098407
transform 1 0 43148 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_469
timestamp 1659098407
transform 1 0 44252 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_475
timestamp 1659098407
transform 1 0 44804 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_477
timestamp 1659098407
transform 1 0 44988 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_489
timestamp 1659098407
transform 1 0 46092 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_501
timestamp 1659098407
transform 1 0 47196 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_40_512
timestamp 1659098407
transform 1 0 48208 0 1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_41_6
timestamp 1659098407
transform 1 0 1656 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_18
timestamp 1659098407
transform 1 0 2760 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_30
timestamp 1659098407
transform 1 0 3864 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_42
timestamp 1659098407
transform 1 0 4968 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_41_54
timestamp 1659098407
transform 1 0 6072 0 -1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_41_57
timestamp 1659098407
transform 1 0 6348 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_69
timestamp 1659098407
transform 1 0 7452 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_81
timestamp 1659098407
transform 1 0 8556 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_93
timestamp 1659098407
transform 1 0 9660 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_105
timestamp 1659098407
transform 1 0 10764 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_111
timestamp 1659098407
transform 1 0 11316 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_113
timestamp 1659098407
transform 1 0 11500 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_125
timestamp 1659098407
transform 1 0 12604 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_137
timestamp 1659098407
transform 1 0 13708 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_149
timestamp 1659098407
transform 1 0 14812 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_161
timestamp 1659098407
transform 1 0 15916 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_167
timestamp 1659098407
transform 1 0 16468 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_169
timestamp 1659098407
transform 1 0 16652 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_181
timestamp 1659098407
transform 1 0 17756 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_193
timestamp 1659098407
transform 1 0 18860 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_205
timestamp 1659098407
transform 1 0 19964 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_217
timestamp 1659098407
transform 1 0 21068 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_223
timestamp 1659098407
transform 1 0 21620 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_225
timestamp 1659098407
transform 1 0 21804 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_237
timestamp 1659098407
transform 1 0 22908 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_249
timestamp 1659098407
transform 1 0 24012 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_261
timestamp 1659098407
transform 1 0 25116 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_273
timestamp 1659098407
transform 1 0 26220 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_279
timestamp 1659098407
transform 1 0 26772 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_281
timestamp 1659098407
transform 1 0 26956 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_293
timestamp 1659098407
transform 1 0 28060 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_305
timestamp 1659098407
transform 1 0 29164 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_317
timestamp 1659098407
transform 1 0 30268 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_329
timestamp 1659098407
transform 1 0 31372 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_335
timestamp 1659098407
transform 1 0 31924 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_337
timestamp 1659098407
transform 1 0 32108 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_349
timestamp 1659098407
transform 1 0 33212 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_361
timestamp 1659098407
transform 1 0 34316 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_373
timestamp 1659098407
transform 1 0 35420 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_385
timestamp 1659098407
transform 1 0 36524 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_391
timestamp 1659098407
transform 1 0 37076 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_393
timestamp 1659098407
transform 1 0 37260 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_405
timestamp 1659098407
transform 1 0 38364 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_417
timestamp 1659098407
transform 1 0 39468 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_429
timestamp 1659098407
transform 1 0 40572 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_441
timestamp 1659098407
transform 1 0 41676 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_447
timestamp 1659098407
transform 1 0 42228 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_449
timestamp 1659098407
transform 1 0 42412 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_461
timestamp 1659098407
transform 1 0 43516 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_473
timestamp 1659098407
transform 1 0 44620 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_485
timestamp 1659098407
transform 1 0 45724 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_497
timestamp 1659098407
transform 1 0 46828 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_503
timestamp 1659098407
transform 1 0 47380 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_505
timestamp 1659098407
transform 1 0 47564 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_512
timestamp 1659098407
transform 1 0 48208 0 -1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_42_6
timestamp 1659098407
transform 1 0 1656 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_42_18
timestamp 1659098407
transform 1 0 2760 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_42_26
timestamp 1659098407
transform 1 0 3496 0 1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_42_29
timestamp 1659098407
transform 1 0 3772 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_41
timestamp 1659098407
transform 1 0 4876 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_53
timestamp 1659098407
transform 1 0 5980 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_65
timestamp 1659098407
transform 1 0 7084 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_77
timestamp 1659098407
transform 1 0 8188 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_83
timestamp 1659098407
transform 1 0 8740 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_85
timestamp 1659098407
transform 1 0 8924 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_97
timestamp 1659098407
transform 1 0 10028 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_109
timestamp 1659098407
transform 1 0 11132 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_121
timestamp 1659098407
transform 1 0 12236 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_133
timestamp 1659098407
transform 1 0 13340 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_139
timestamp 1659098407
transform 1 0 13892 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_141
timestamp 1659098407
transform 1 0 14076 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_153
timestamp 1659098407
transform 1 0 15180 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_165
timestamp 1659098407
transform 1 0 16284 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_177
timestamp 1659098407
transform 1 0 17388 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_189
timestamp 1659098407
transform 1 0 18492 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_195
timestamp 1659098407
transform 1 0 19044 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_197
timestamp 1659098407
transform 1 0 19228 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_209
timestamp 1659098407
transform 1 0 20332 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_221
timestamp 1659098407
transform 1 0 21436 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_233
timestamp 1659098407
transform 1 0 22540 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_245
timestamp 1659098407
transform 1 0 23644 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_251
timestamp 1659098407
transform 1 0 24196 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_253
timestamp 1659098407
transform 1 0 24380 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_265
timestamp 1659098407
transform 1 0 25484 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_277
timestamp 1659098407
transform 1 0 26588 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_289
timestamp 1659098407
transform 1 0 27692 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_301
timestamp 1659098407
transform 1 0 28796 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_307
timestamp 1659098407
transform 1 0 29348 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_309
timestamp 1659098407
transform 1 0 29532 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_321
timestamp 1659098407
transform 1 0 30636 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_333
timestamp 1659098407
transform 1 0 31740 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_345
timestamp 1659098407
transform 1 0 32844 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_357
timestamp 1659098407
transform 1 0 33948 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_363
timestamp 1659098407
transform 1 0 34500 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_365
timestamp 1659098407
transform 1 0 34684 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_377
timestamp 1659098407
transform 1 0 35788 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_389
timestamp 1659098407
transform 1 0 36892 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_401
timestamp 1659098407
transform 1 0 37996 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_413
timestamp 1659098407
transform 1 0 39100 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_419
timestamp 1659098407
transform 1 0 39652 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_421
timestamp 1659098407
transform 1 0 39836 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_433
timestamp 1659098407
transform 1 0 40940 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_445
timestamp 1659098407
transform 1 0 42044 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_457
timestamp 1659098407
transform 1 0 43148 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_469
timestamp 1659098407
transform 1 0 44252 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_475
timestamp 1659098407
transform 1 0 44804 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_477
timestamp 1659098407
transform 1 0 44988 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_489
timestamp 1659098407
transform 1 0 46092 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_42_501
timestamp 1659098407
transform 1 0 47196 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_42_512
timestamp 1659098407
transform 1 0 48208 0 1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_43_6
timestamp 1659098407
transform 1 0 1656 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_18
timestamp 1659098407
transform 1 0 2760 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_30
timestamp 1659098407
transform 1 0 3864 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_42
timestamp 1659098407
transform 1 0 4968 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_43_54
timestamp 1659098407
transform 1 0 6072 0 -1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_43_57
timestamp 1659098407
transform 1 0 6348 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_69
timestamp 1659098407
transform 1 0 7452 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_81
timestamp 1659098407
transform 1 0 8556 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_93
timestamp 1659098407
transform 1 0 9660 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_105
timestamp 1659098407
transform 1 0 10764 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_111
timestamp 1659098407
transform 1 0 11316 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_113
timestamp 1659098407
transform 1 0 11500 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_125
timestamp 1659098407
transform 1 0 12604 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_137
timestamp 1659098407
transform 1 0 13708 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_149
timestamp 1659098407
transform 1 0 14812 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_161
timestamp 1659098407
transform 1 0 15916 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_167
timestamp 1659098407
transform 1 0 16468 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_169
timestamp 1659098407
transform 1 0 16652 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_181
timestamp 1659098407
transform 1 0 17756 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_193
timestamp 1659098407
transform 1 0 18860 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_205
timestamp 1659098407
transform 1 0 19964 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_217
timestamp 1659098407
transform 1 0 21068 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_223
timestamp 1659098407
transform 1 0 21620 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_225
timestamp 1659098407
transform 1 0 21804 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_237
timestamp 1659098407
transform 1 0 22908 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_249
timestamp 1659098407
transform 1 0 24012 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_261
timestamp 1659098407
transform 1 0 25116 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_273
timestamp 1659098407
transform 1 0 26220 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_279
timestamp 1659098407
transform 1 0 26772 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_281
timestamp 1659098407
transform 1 0 26956 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_293
timestamp 1659098407
transform 1 0 28060 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_305
timestamp 1659098407
transform 1 0 29164 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_317
timestamp 1659098407
transform 1 0 30268 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_329
timestamp 1659098407
transform 1 0 31372 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_335
timestamp 1659098407
transform 1 0 31924 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_337
timestamp 1659098407
transform 1 0 32108 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_349
timestamp 1659098407
transform 1 0 33212 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_361
timestamp 1659098407
transform 1 0 34316 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_373
timestamp 1659098407
transform 1 0 35420 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_385
timestamp 1659098407
transform 1 0 36524 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_391
timestamp 1659098407
transform 1 0 37076 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_393
timestamp 1659098407
transform 1 0 37260 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_405
timestamp 1659098407
transform 1 0 38364 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_417
timestamp 1659098407
transform 1 0 39468 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_429
timestamp 1659098407
transform 1 0 40572 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_441
timestamp 1659098407
transform 1 0 41676 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_447
timestamp 1659098407
transform 1 0 42228 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_449
timestamp 1659098407
transform 1 0 42412 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_461
timestamp 1659098407
transform 1 0 43516 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_473
timestamp 1659098407
transform 1 0 44620 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_485
timestamp 1659098407
transform 1 0 45724 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_500
timestamp 1659098407
transform 1 0 47104 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_505
timestamp 1659098407
transform 1 0 47564 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_512
timestamp 1659098407
transform 1 0 48208 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_6
timestamp 1659098407
transform 1 0 1656 0 1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_44_13
timestamp 1659098407
transform 1 0 2300 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_44_25
timestamp 1659098407
transform 1 0 3404 0 1 26112
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_44_29
timestamp 1659098407
transform 1 0 3772 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_41
timestamp 1659098407
transform 1 0 4876 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_53
timestamp 1659098407
transform 1 0 5980 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_65
timestamp 1659098407
transform 1 0 7084 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_77
timestamp 1659098407
transform 1 0 8188 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_83
timestamp 1659098407
transform 1 0 8740 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_85
timestamp 1659098407
transform 1 0 8924 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_97
timestamp 1659098407
transform 1 0 10028 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_109
timestamp 1659098407
transform 1 0 11132 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_121
timestamp 1659098407
transform 1 0 12236 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_133
timestamp 1659098407
transform 1 0 13340 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_139
timestamp 1659098407
transform 1 0 13892 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_141
timestamp 1659098407
transform 1 0 14076 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_153
timestamp 1659098407
transform 1 0 15180 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_165
timestamp 1659098407
transform 1 0 16284 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_177
timestamp 1659098407
transform 1 0 17388 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_189
timestamp 1659098407
transform 1 0 18492 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_195
timestamp 1659098407
transform 1 0 19044 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_197
timestamp 1659098407
transform 1 0 19228 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_209
timestamp 1659098407
transform 1 0 20332 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_221
timestamp 1659098407
transform 1 0 21436 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_233
timestamp 1659098407
transform 1 0 22540 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_245
timestamp 1659098407
transform 1 0 23644 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_251
timestamp 1659098407
transform 1 0 24196 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_253
timestamp 1659098407
transform 1 0 24380 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_265
timestamp 1659098407
transform 1 0 25484 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_277
timestamp 1659098407
transform 1 0 26588 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_289
timestamp 1659098407
transform 1 0 27692 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_301
timestamp 1659098407
transform 1 0 28796 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_307
timestamp 1659098407
transform 1 0 29348 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_309
timestamp 1659098407
transform 1 0 29532 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_321
timestamp 1659098407
transform 1 0 30636 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_333
timestamp 1659098407
transform 1 0 31740 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_345
timestamp 1659098407
transform 1 0 32844 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_357
timestamp 1659098407
transform 1 0 33948 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_363
timestamp 1659098407
transform 1 0 34500 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_365
timestamp 1659098407
transform 1 0 34684 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_377
timestamp 1659098407
transform 1 0 35788 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_389
timestamp 1659098407
transform 1 0 36892 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_401
timestamp 1659098407
transform 1 0 37996 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_413
timestamp 1659098407
transform 1 0 39100 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_419
timestamp 1659098407
transform 1 0 39652 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_421
timestamp 1659098407
transform 1 0 39836 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_433
timestamp 1659098407
transform 1 0 40940 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_445
timestamp 1659098407
transform 1 0 42044 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_457
timestamp 1659098407
transform 1 0 43148 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_469
timestamp 1659098407
transform 1 0 44252 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_475
timestamp 1659098407
transform 1 0 44804 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_477
timestamp 1659098407
transform 1 0 44988 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_489
timestamp 1659098407
transform 1 0 46092 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_44_498
timestamp 1659098407
transform 1 0 46920 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_505
timestamp 1659098407
transform 1 0 47564 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_512
timestamp 1659098407
transform 1 0 48208 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_6
timestamp 1659098407
transform 1 0 1656 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_13
timestamp 1659098407
transform 1 0 2300 0 -1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_45_20
timestamp 1659098407
transform 1 0 2944 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_32
timestamp 1659098407
transform 1 0 4048 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_44
timestamp 1659098407
transform 1 0 5152 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_45_57
timestamp 1659098407
transform 1 0 6348 0 -1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_45_62
timestamp 1659098407
transform 1 0 6808 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_74
timestamp 1659098407
transform 1 0 7912 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_45_86
timestamp 1659098407
transform 1 0 9016 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_90
timestamp 1659098407
transform 1 0 9384 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_45_102
timestamp 1659098407
transform 1 0 10488 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_45_110
timestamp 1659098407
transform 1 0 11224 0 -1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_45_113
timestamp 1659098407
transform 1 0 11500 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_125
timestamp 1659098407
transform 1 0 12604 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_137
timestamp 1659098407
transform 1 0 13708 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_149
timestamp 1659098407
transform 1 0 14812 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_161
timestamp 1659098407
transform 1 0 15916 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_167
timestamp 1659098407
transform 1 0 16468 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_169
timestamp 1659098407
transform 1 0 16652 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_181
timestamp 1659098407
transform 1 0 17756 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_193
timestamp 1659098407
transform 1 0 18860 0 -1 27200
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_45_202
timestamp 1659098407
transform 1 0 19688 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_45_214
timestamp 1659098407
transform 1 0 20792 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_45_222
timestamp 1659098407
transform 1 0 21528 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_225
timestamp 1659098407
transform 1 0 21804 0 -1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_45_230
timestamp 1659098407
transform 1 0 22264 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_242
timestamp 1659098407
transform 1 0 23368 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_254
timestamp 1659098407
transform 1 0 24472 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_266
timestamp 1659098407
transform 1 0 25576 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_45_278
timestamp 1659098407
transform 1 0 26680 0 -1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_45_281
timestamp 1659098407
transform 1 0 26956 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_293
timestamp 1659098407
transform 1 0 28060 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_305
timestamp 1659098407
transform 1 0 29164 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_317
timestamp 1659098407
transform 1 0 30268 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_329
timestamp 1659098407
transform 1 0 31372 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_335
timestamp 1659098407
transform 1 0 31924 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_337
timestamp 1659098407
transform 1 0 32108 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_349
timestamp 1659098407
transform 1 0 33212 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_361
timestamp 1659098407
transform 1 0 34316 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_45_373
timestamp 1659098407
transform 1 0 35420 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_45_384
timestamp 1659098407
transform 1 0 36432 0 -1 27200
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_45_393
timestamp 1659098407
transform 1 0 37260 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_405
timestamp 1659098407
transform 1 0 38364 0 -1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_45_412
timestamp 1659098407
transform 1 0 39008 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_424
timestamp 1659098407
transform 1 0 40112 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_436
timestamp 1659098407
transform 1 0 41216 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_452
timestamp 1659098407
transform 1 0 42688 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_45_464
timestamp 1659098407
transform 1 0 43792 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_468
timestamp 1659098407
transform 1 0 44160 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_45_480
timestamp 1659098407
transform 1 0 45264 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_45_486
timestamp 1659098407
transform 1 0 45816 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_493
timestamp 1659098407
transform 1 0 46460 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_500
timestamp 1659098407
transform 1 0 47104 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_45_508
timestamp 1659098407
transform 1 0 47840 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_46_6
timestamp 1659098407
transform 1 0 1656 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_13
timestamp 1659098407
transform 1 0 2300 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_46_20
timestamp 1659098407
transform 1 0 2944 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_46_29
timestamp 1659098407
transform 1 0 3772 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_46_34
timestamp 1659098407
transform 1 0 4232 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_46_45
timestamp 1659098407
transform 1 0 5244 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_52
timestamp 1659098407
transform 1 0 5888 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_46_57
timestamp 1659098407
transform 1 0 6348 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_46_66
timestamp 1659098407
transform 1 0 7176 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_73
timestamp 1659098407
transform 1 0 7820 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_80
timestamp 1659098407
transform 1 0 8464 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_46_85
timestamp 1659098407
transform 1 0 8924 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_46_94
timestamp 1659098407
transform 1 0 9752 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_101
timestamp 1659098407
transform 1 0 10396 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_108
timestamp 1659098407
transform 1 0 11040 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_46_113
timestamp 1659098407
transform 1 0 11500 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_118
timestamp 1659098407
transform 1 0 11960 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_125
timestamp 1659098407
transform 1 0 12604 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_46_132
timestamp 1659098407
transform 1 0 13248 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_46_144
timestamp 1659098407
transform 1 0 14352 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_46_153
timestamp 1659098407
transform 1 0 15180 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_46_160
timestamp 1659098407
transform 1 0 15824 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_46_172
timestamp 1659098407
transform 1 0 16928 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_46_180
timestamp 1659098407
transform 1 0 17664 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_185
timestamp 1659098407
transform 1 0 18124 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_192
timestamp 1659098407
transform 1 0 18768 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_46_197
timestamp 1659098407
transform 1 0 19228 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_46_206
timestamp 1659098407
transform 1 0 20056 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_213
timestamp 1659098407
transform 1 0 20700 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_220
timestamp 1659098407
transform 1 0 21344 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_46_225
timestamp 1659098407
transform 1 0 21804 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_46_234
timestamp 1659098407
transform 1 0 22632 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_241
timestamp 1659098407
transform 1 0 23276 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_248
timestamp 1659098407
transform 1 0 23920 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_46_253
timestamp 1659098407
transform 1 0 24380 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_258
timestamp 1659098407
transform 1 0 24840 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_265
timestamp 1659098407
transform 1 0 25484 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_46_272
timestamp 1659098407
transform 1 0 26128 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_46_284
timestamp 1659098407
transform 1 0 27232 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_46_293
timestamp 1659098407
transform 1 0 28060 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_46_300
timestamp 1659098407
transform 1 0 28704 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_46_312
timestamp 1659098407
transform 1 0 29808 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_46_321
timestamp 1659098407
transform 1 0 30636 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_46_328
timestamp 1659098407
transform 1 0 31280 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_46_337
timestamp 1659098407
transform 1 0 32108 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_46_342
timestamp 1659098407
transform 1 0 32568 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_46_350
timestamp 1659098407
transform 1 0 33304 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_46_356
timestamp 1659098407
transform 1 0 33856 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_46_368
timestamp 1659098407
transform 1 0 34960 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_375
timestamp 1659098407
transform 1 0 35604 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_46_382
timestamp 1659098407
transform 1 0 36248 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_46_390
timestamp 1659098407
transform 1 0 36984 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_396
timestamp 1659098407
transform 1 0 37536 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_403
timestamp 1659098407
transform 1 0 38180 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_46_410
timestamp 1659098407
transform 1 0 38824 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_46_418
timestamp 1659098407
transform 1 0 39560 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_46_421
timestamp 1659098407
transform 1 0 39836 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_426
timestamp 1659098407
transform 1 0 40296 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_433
timestamp 1659098407
transform 1 0 40940 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_46_440
timestamp 1659098407
transform 1 0 41584 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_46_449
timestamp 1659098407
transform 1 0 42412 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_461
timestamp 1659098407
transform 1 0 43516 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_46_468
timestamp 1659098407
transform 1 0 44160 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_46_477
timestamp 1659098407
transform 1 0 44988 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_482
timestamp 1659098407
transform 1 0 45448 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_489
timestamp 1659098407
transform 1 0 46092 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_46_496
timestamp 1659098407
transform 1 0 46736 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_46_505
timestamp 1659098407
transform 1 0 47564 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_46_512
timestamp 1659098407
transform 1 0 48208 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1659098407
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1659098407
transform -1 0 48852 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1659098407
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1659098407
transform -1 0 48852 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1659098407
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1659098407
transform -1 0 48852 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1659098407
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1659098407
transform -1 0 48852 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1659098407
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1659098407
transform -1 0 48852 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1659098407
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1659098407
transform -1 0 48852 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1659098407
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1659098407
transform -1 0 48852 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1659098407
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1659098407
transform -1 0 48852 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1659098407
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1659098407
transform -1 0 48852 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1659098407
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1659098407
transform -1 0 48852 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1659098407
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1659098407
transform -1 0 48852 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1659098407
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1659098407
transform -1 0 48852 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1659098407
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1659098407
transform -1 0 48852 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1659098407
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1659098407
transform -1 0 48852 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1659098407
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1659098407
transform -1 0 48852 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1659098407
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1659098407
transform -1 0 48852 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1659098407
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1659098407
transform -1 0 48852 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1659098407
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1659098407
transform -1 0 48852 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1659098407
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1659098407
transform -1 0 48852 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1659098407
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1659098407
transform -1 0 48852 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1659098407
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1659098407
transform -1 0 48852 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1659098407
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1659098407
transform -1 0 48852 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1659098407
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1659098407
transform -1 0 48852 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1659098407
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1659098407
transform -1 0 48852 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1659098407
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1659098407
transform -1 0 48852 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1659098407
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1659098407
transform -1 0 48852 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1659098407
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1659098407
transform -1 0 48852 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1659098407
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1659098407
transform -1 0 48852 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1659098407
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1659098407
transform -1 0 48852 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1659098407
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1659098407
transform -1 0 48852 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1659098407
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1659098407
transform -1 0 48852 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1659098407
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1659098407
transform -1 0 48852 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1659098407
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1659098407
transform -1 0 48852 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1659098407
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1659098407
transform -1 0 48852 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1659098407
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1659098407
transform -1 0 48852 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1659098407
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1659098407
transform -1 0 48852 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1659098407
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1659098407
transform -1 0 48852 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1659098407
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1659098407
transform -1 0 48852 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1659098407
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1659098407
transform -1 0 48852 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1659098407
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1659098407
transform -1 0 48852 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1659098407
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1659098407
transform -1 0 48852 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1659098407
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1659098407
transform -1 0 48852 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1659098407
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1659098407
transform -1 0 48852 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1659098407
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1659098407
transform -1 0 48852 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1659098407
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1659098407
transform -1 0 48852 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1659098407
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1659098407
transform -1 0 48852 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1659098407
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1659098407
transform -1 0 48852 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_94 ../openroad/OpenLane/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1659098407
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_95
timestamp 1659098407
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_96
timestamp 1659098407
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_97
timestamp 1659098407
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_98
timestamp 1659098407
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_99
timestamp 1659098407
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_100
timestamp 1659098407
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_101
timestamp 1659098407
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_102
timestamp 1659098407
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_103
timestamp 1659098407
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_104
timestamp 1659098407
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_105
timestamp 1659098407
transform 1 0 32016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_106
timestamp 1659098407
transform 1 0 34592 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_107
timestamp 1659098407
transform 1 0 37168 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_108
timestamp 1659098407
transform 1 0 39744 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_109
timestamp 1659098407
transform 1 0 42320 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_110
timestamp 1659098407
transform 1 0 44896 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_111
timestamp 1659098407
transform 1 0 47472 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_112
timestamp 1659098407
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_113
timestamp 1659098407
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_114
timestamp 1659098407
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_115
timestamp 1659098407
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_116
timestamp 1659098407
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_117
timestamp 1659098407
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_118
timestamp 1659098407
transform 1 0 37168 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_119
timestamp 1659098407
transform 1 0 42320 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_120
timestamp 1659098407
transform 1 0 47472 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_121
timestamp 1659098407
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_122
timestamp 1659098407
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_123
timestamp 1659098407
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_124
timestamp 1659098407
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_125
timestamp 1659098407
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_126
timestamp 1659098407
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_127
timestamp 1659098407
transform 1 0 34592 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_128
timestamp 1659098407
transform 1 0 39744 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_129
timestamp 1659098407
transform 1 0 44896 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_130
timestamp 1659098407
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_131
timestamp 1659098407
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_132
timestamp 1659098407
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_133
timestamp 1659098407
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_134
timestamp 1659098407
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_135
timestamp 1659098407
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_136
timestamp 1659098407
transform 1 0 37168 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_137
timestamp 1659098407
transform 1 0 42320 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_138
timestamp 1659098407
transform 1 0 47472 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_139
timestamp 1659098407
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_140
timestamp 1659098407
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_141
timestamp 1659098407
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_142
timestamp 1659098407
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_143
timestamp 1659098407
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_144
timestamp 1659098407
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_145
timestamp 1659098407
transform 1 0 34592 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_146
timestamp 1659098407
transform 1 0 39744 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_147
timestamp 1659098407
transform 1 0 44896 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_148
timestamp 1659098407
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_149
timestamp 1659098407
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_150
timestamp 1659098407
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_151
timestamp 1659098407
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_152
timestamp 1659098407
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_153
timestamp 1659098407
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_154
timestamp 1659098407
transform 1 0 37168 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_155
timestamp 1659098407
transform 1 0 42320 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_156
timestamp 1659098407
transform 1 0 47472 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_157
timestamp 1659098407
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_158
timestamp 1659098407
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_159
timestamp 1659098407
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160
timestamp 1659098407
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 1659098407
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 1659098407
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 1659098407
transform 1 0 34592 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_164
timestamp 1659098407
transform 1 0 39744 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_165
timestamp 1659098407
transform 1 0 44896 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166
timestamp 1659098407
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1659098407
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1659098407
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1659098407
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1659098407
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1659098407
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1659098407
transform 1 0 37168 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1659098407
transform 1 0 42320 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1659098407
transform 1 0 47472 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1659098407
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1659098407
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1659098407
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1659098407
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1659098407
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1659098407
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1659098407
transform 1 0 34592 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1659098407
transform 1 0 39744 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1659098407
transform 1 0 44896 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1659098407
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1659098407
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1659098407
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1659098407
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1659098407
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1659098407
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1659098407
transform 1 0 37168 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1659098407
transform 1 0 42320 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1659098407
transform 1 0 47472 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1659098407
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1659098407
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1659098407
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1659098407
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1659098407
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1659098407
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1659098407
transform 1 0 34592 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1659098407
transform 1 0 39744 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1659098407
transform 1 0 44896 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1659098407
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1659098407
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1659098407
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1659098407
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1659098407
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1659098407
transform 1 0 32016 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1659098407
transform 1 0 37168 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1659098407
transform 1 0 42320 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1659098407
transform 1 0 47472 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1659098407
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1659098407
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1659098407
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1659098407
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1659098407
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1659098407
transform 1 0 29440 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1659098407
transform 1 0 34592 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1659098407
transform 1 0 39744 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1659098407
transform 1 0 44896 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1659098407
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1659098407
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1659098407
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1659098407
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1659098407
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1659098407
transform 1 0 32016 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1659098407
transform 1 0 37168 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1659098407
transform 1 0 42320 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1659098407
transform 1 0 47472 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1659098407
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1659098407
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1659098407
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1659098407
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1659098407
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1659098407
transform 1 0 29440 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1659098407
transform 1 0 34592 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1659098407
transform 1 0 39744 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1659098407
transform 1 0 44896 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1659098407
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1659098407
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1659098407
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1659098407
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1659098407
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1659098407
transform 1 0 32016 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1659098407
transform 1 0 37168 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1659098407
transform 1 0 42320 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1659098407
transform 1 0 47472 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1659098407
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1659098407
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1659098407
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1659098407
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1659098407
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1659098407
transform 1 0 29440 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1659098407
transform 1 0 34592 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1659098407
transform 1 0 39744 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1659098407
transform 1 0 44896 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1659098407
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1659098407
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1659098407
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1659098407
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1659098407
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1659098407
transform 1 0 32016 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1659098407
transform 1 0 37168 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1659098407
transform 1 0 42320 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1659098407
transform 1 0 47472 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1659098407
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1659098407
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1659098407
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1659098407
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1659098407
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1659098407
transform 1 0 29440 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1659098407
transform 1 0 34592 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1659098407
transform 1 0 39744 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1659098407
transform 1 0 44896 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1659098407
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1659098407
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1659098407
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1659098407
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1659098407
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1659098407
transform 1 0 32016 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1659098407
transform 1 0 37168 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1659098407
transform 1 0 42320 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1659098407
transform 1 0 47472 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1659098407
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1659098407
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1659098407
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1659098407
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1659098407
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1659098407
transform 1 0 29440 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1659098407
transform 1 0 34592 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1659098407
transform 1 0 39744 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1659098407
transform 1 0 44896 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1659098407
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1659098407
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1659098407
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1659098407
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1659098407
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1659098407
transform 1 0 32016 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1659098407
transform 1 0 37168 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1659098407
transform 1 0 42320 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1659098407
transform 1 0 47472 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1659098407
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1659098407
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1659098407
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1659098407
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1659098407
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1659098407
transform 1 0 29440 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1659098407
transform 1 0 34592 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1659098407
transform 1 0 39744 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1659098407
transform 1 0 44896 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1659098407
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1659098407
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1659098407
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1659098407
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1659098407
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1659098407
transform 1 0 32016 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1659098407
transform 1 0 37168 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1659098407
transform 1 0 42320 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1659098407
transform 1 0 47472 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1659098407
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1659098407
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1659098407
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1659098407
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1659098407
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1659098407
transform 1 0 29440 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1659098407
transform 1 0 34592 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1659098407
transform 1 0 39744 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1659098407
transform 1 0 44896 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1659098407
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1659098407
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1659098407
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1659098407
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1659098407
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1659098407
transform 1 0 32016 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1659098407
transform 1 0 37168 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1659098407
transform 1 0 42320 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1659098407
transform 1 0 47472 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1659098407
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1659098407
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1659098407
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1659098407
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1659098407
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1659098407
transform 1 0 29440 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1659098407
transform 1 0 34592 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1659098407
transform 1 0 39744 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1659098407
transform 1 0 44896 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1659098407
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1659098407
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1659098407
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1659098407
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1659098407
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1659098407
transform 1 0 32016 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1659098407
transform 1 0 37168 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1659098407
transform 1 0 42320 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1659098407
transform 1 0 47472 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1659098407
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 1659098407
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 1659098407
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 1659098407
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 1659098407
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 1659098407
transform 1 0 29440 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 1659098407
transform 1 0 34592 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 1659098407
transform 1 0 39744 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 1659098407
transform 1 0 44896 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 1659098407
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 1659098407
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 1659098407
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 1659098407
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 1659098407
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 1659098407
transform 1 0 32016 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 1659098407
transform 1 0 37168 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 1659098407
transform 1 0 42320 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 1659098407
transform 1 0 47472 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 1659098407
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_374
timestamp 1659098407
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_375
timestamp 1659098407
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_376
timestamp 1659098407
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_377
timestamp 1659098407
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_378
timestamp 1659098407
transform 1 0 29440 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_379
timestamp 1659098407
transform 1 0 34592 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_380
timestamp 1659098407
transform 1 0 39744 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_381
timestamp 1659098407
transform 1 0 44896 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_382
timestamp 1659098407
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_383
timestamp 1659098407
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_384
timestamp 1659098407
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_385
timestamp 1659098407
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_386
timestamp 1659098407
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_387
timestamp 1659098407
transform 1 0 32016 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_388
timestamp 1659098407
transform 1 0 37168 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_389
timestamp 1659098407
transform 1 0 42320 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_390
timestamp 1659098407
transform 1 0 47472 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_391
timestamp 1659098407
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_392
timestamp 1659098407
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_393
timestamp 1659098407
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_394
timestamp 1659098407
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_395
timestamp 1659098407
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_396
timestamp 1659098407
transform 1 0 29440 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_397
timestamp 1659098407
transform 1 0 34592 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_398
timestamp 1659098407
transform 1 0 39744 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_399
timestamp 1659098407
transform 1 0 44896 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_400
timestamp 1659098407
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_401
timestamp 1659098407
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_402
timestamp 1659098407
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_403
timestamp 1659098407
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_404
timestamp 1659098407
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_405
timestamp 1659098407
transform 1 0 32016 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_406
timestamp 1659098407
transform 1 0 37168 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_407
timestamp 1659098407
transform 1 0 42320 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_408
timestamp 1659098407
transform 1 0 47472 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_409
timestamp 1659098407
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_410
timestamp 1659098407
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_411
timestamp 1659098407
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_412
timestamp 1659098407
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_413
timestamp 1659098407
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_414
timestamp 1659098407
transform 1 0 29440 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_415
timestamp 1659098407
transform 1 0 34592 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_416
timestamp 1659098407
transform 1 0 39744 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_417
timestamp 1659098407
transform 1 0 44896 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_418
timestamp 1659098407
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_419
timestamp 1659098407
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_420
timestamp 1659098407
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_421
timestamp 1659098407
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_422
timestamp 1659098407
transform 1 0 26864 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_423
timestamp 1659098407
transform 1 0 32016 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_424
timestamp 1659098407
transform 1 0 37168 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_425
timestamp 1659098407
transform 1 0 42320 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_426
timestamp 1659098407
transform 1 0 47472 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_427
timestamp 1659098407
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_428
timestamp 1659098407
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_429
timestamp 1659098407
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_430
timestamp 1659098407
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_431
timestamp 1659098407
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_432
timestamp 1659098407
transform 1 0 29440 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_433
timestamp 1659098407
transform 1 0 34592 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_434
timestamp 1659098407
transform 1 0 39744 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_435
timestamp 1659098407
transform 1 0 44896 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_436
timestamp 1659098407
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_437
timestamp 1659098407
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_438
timestamp 1659098407
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_439
timestamp 1659098407
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_440
timestamp 1659098407
transform 1 0 26864 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_441
timestamp 1659098407
transform 1 0 32016 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_442
timestamp 1659098407
transform 1 0 37168 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_443
timestamp 1659098407
transform 1 0 42320 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_444
timestamp 1659098407
transform 1 0 47472 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_445
timestamp 1659098407
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_446
timestamp 1659098407
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_447
timestamp 1659098407
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_448
timestamp 1659098407
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_449
timestamp 1659098407
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_450
timestamp 1659098407
transform 1 0 29440 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_451
timestamp 1659098407
transform 1 0 34592 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_452
timestamp 1659098407
transform 1 0 39744 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_453
timestamp 1659098407
transform 1 0 44896 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_454
timestamp 1659098407
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_455
timestamp 1659098407
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_456
timestamp 1659098407
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_457
timestamp 1659098407
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_458
timestamp 1659098407
transform 1 0 26864 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_459
timestamp 1659098407
transform 1 0 32016 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_460
timestamp 1659098407
transform 1 0 37168 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_461
timestamp 1659098407
transform 1 0 42320 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_462
timestamp 1659098407
transform 1 0 47472 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_463
timestamp 1659098407
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_464
timestamp 1659098407
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_465
timestamp 1659098407
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_466
timestamp 1659098407
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_467
timestamp 1659098407
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_468
timestamp 1659098407
transform 1 0 29440 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_469
timestamp 1659098407
transform 1 0 34592 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_470
timestamp 1659098407
transform 1 0 39744 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_471
timestamp 1659098407
transform 1 0 44896 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_472
timestamp 1659098407
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_473
timestamp 1659098407
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_474
timestamp 1659098407
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_475
timestamp 1659098407
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_476
timestamp 1659098407
transform 1 0 26864 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_477
timestamp 1659098407
transform 1 0 32016 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_478
timestamp 1659098407
transform 1 0 37168 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_479
timestamp 1659098407
transform 1 0 42320 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_480
timestamp 1659098407
transform 1 0 47472 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_481
timestamp 1659098407
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_482
timestamp 1659098407
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_483
timestamp 1659098407
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_484
timestamp 1659098407
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_485
timestamp 1659098407
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_486
timestamp 1659098407
transform 1 0 29440 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_487
timestamp 1659098407
transform 1 0 34592 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_488
timestamp 1659098407
transform 1 0 39744 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_489
timestamp 1659098407
transform 1 0 44896 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_490
timestamp 1659098407
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_491
timestamp 1659098407
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_492
timestamp 1659098407
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_493
timestamp 1659098407
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_494
timestamp 1659098407
transform 1 0 26864 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_495
timestamp 1659098407
transform 1 0 32016 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_496
timestamp 1659098407
transform 1 0 37168 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_497
timestamp 1659098407
transform 1 0 42320 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_498
timestamp 1659098407
transform 1 0 47472 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_499
timestamp 1659098407
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_500
timestamp 1659098407
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_501
timestamp 1659098407
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_502
timestamp 1659098407
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_503
timestamp 1659098407
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_504
timestamp 1659098407
transform 1 0 29440 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_505
timestamp 1659098407
transform 1 0 34592 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_506
timestamp 1659098407
transform 1 0 39744 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_507
timestamp 1659098407
transform 1 0 44896 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_508
timestamp 1659098407
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_509
timestamp 1659098407
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_510
timestamp 1659098407
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_511
timestamp 1659098407
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_512
timestamp 1659098407
transform 1 0 26864 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_513
timestamp 1659098407
transform 1 0 32016 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_514
timestamp 1659098407
transform 1 0 37168 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_515
timestamp 1659098407
transform 1 0 42320 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_516
timestamp 1659098407
transform 1 0 47472 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_517
timestamp 1659098407
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_518
timestamp 1659098407
transform 1 0 6256 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_519
timestamp 1659098407
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_520
timestamp 1659098407
transform 1 0 11408 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_521
timestamp 1659098407
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_522
timestamp 1659098407
transform 1 0 16560 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_523
timestamp 1659098407
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_524
timestamp 1659098407
transform 1 0 21712 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_525
timestamp 1659098407
transform 1 0 24288 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_526
timestamp 1659098407
transform 1 0 26864 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_527
timestamp 1659098407
transform 1 0 29440 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_528
timestamp 1659098407
transform 1 0 32016 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_529
timestamp 1659098407
transform 1 0 34592 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_530
timestamp 1659098407
transform 1 0 37168 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_531
timestamp 1659098407
transform 1 0 39744 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_532
timestamp 1659098407
transform 1 0 42320 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_533
timestamp 1659098407
transform 1 0 44896 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_534
timestamp 1659098407
transform 1 0 47472 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__nand2_1  _008_ ../openroad/OpenLane/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1659098407
transform -1 0 47840 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _009_ ../openroad/OpenLane/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1659098407
transform -1 0 47472 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _010_ ../openroad/OpenLane/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1659098407
transform -1 0 46368 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _011_ ../openroad/OpenLane/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1659098407
transform 1 0 47564 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _012_
timestamp 1659098407
transform -1 0 45264 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _013_
timestamp 1659098407
transform -1 0 46552 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _014_
timestamp 1659098407
transform -1 0 45908 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _015_
timestamp 1659098407
transform -1 0 41124 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  _016_ ../openroad/OpenLane/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1659098407
transform 1 0 43240 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _017_
timestamp 1659098407
transform 1 0 39836 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _018_
timestamp 1659098407
transform 1 0 34868 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _019_
timestamp 1659098407
transform 1 0 27876 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__conb_1  _020__153 ../openroad/OpenLane/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1659098407
transform 1 0 25116 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  _020_
timestamp 1659098407
transform 1 0 24656 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__buf_2  _220_
timestamp 1659098407
transform -1 0 22724 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _221_ ../openroad/OpenLane/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1659098407
transform 1 0 22724 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  clk_rst_gen_7
timestamp 1659098407
transform -1 0 1656 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  clk_rst_gen_8
timestamp 1659098407
transform 1 0 47932 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  clk_rst_gen_9
timestamp 1659098407
transform -1 0 27232 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  clk_rst_gen_10
timestamp 1659098407
transform 1 0 47932 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  clk_rst_gen_11
timestamp 1659098407
transform -1 0 1656 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  clk_rst_gen_12
timestamp 1659098407
transform 1 0 23644 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  clk_rst_gen_13
timestamp 1659098407
transform -1 0 39008 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  clk_rst_gen_14
timestamp 1659098407
transform 1 0 47932 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  clk_rst_gen_15
timestamp 1659098407
transform 1 0 10764 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  clk_rst_gen_16
timestamp 1659098407
transform -1 0 27232 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  clk_rst_gen_17
timestamp 1659098407
transform 1 0 17848 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  clk_rst_gen_18
timestamp 1659098407
transform -1 0 34960 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  clk_rst_gen_19
timestamp 1659098407
transform 1 0 4968 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  clk_rst_gen_20
timestamp 1659098407
transform -1 0 31280 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  clk_rst_gen_21
timestamp 1659098407
transform 1 0 47932 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  clk_rst_gen_22
timestamp 1659098407
transform 1 0 47932 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  clk_rst_gen_23
timestamp 1659098407
transform 1 0 47932 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  clk_rst_gen_24
timestamp 1659098407
transform -1 0 1656 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  clk_rst_gen_25
timestamp 1659098407
transform -1 0 46736 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  clk_rst_gen_26
timestamp 1659098407
transform -1 0 14352 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  clk_rst_gen_27
timestamp 1659098407
transform 1 0 47932 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  clk_rst_gen_28
timestamp 1659098407
transform 1 0 18492 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  clk_rst_gen_29
timestamp 1659098407
transform -1 0 6808 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  clk_rst_gen_30
timestamp 1659098407
transform -1 0 9384 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  clk_rst_gen_31
timestamp 1659098407
transform -1 0 44160 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  clk_rst_gen_32
timestamp 1659098407
transform -1 0 1656 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  clk_rst_gen_33
timestamp 1659098407
transform -1 0 1656 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  clk_rst_gen_34
timestamp 1659098407
transform 1 0 47932 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  clk_rst_gen_35
timestamp 1659098407
transform -1 0 2300 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  clk_rst_gen_36
timestamp 1659098407
transform -1 0 41584 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  clk_rst_gen_37
timestamp 1659098407
transform 1 0 20424 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  clk_rst_gen_38
timestamp 1659098407
transform -1 0 32568 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  clk_rst_gen_39
timestamp 1659098407
transform 1 0 47932 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  clk_rst_gen_40
timestamp 1659098407
transform -1 0 22264 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  clk_rst_gen_41
timestamp 1659098407
transform -1 0 44160 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  clk_rst_gen_42
timestamp 1659098407
transform 1 0 47932 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  clk_rst_gen_43
timestamp 1659098407
transform -1 0 46092 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  clk_rst_gen_44
timestamp 1659098407
transform 1 0 46184 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  clk_rst_gen_45
timestamp 1659098407
transform -1 0 1656 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  clk_rst_gen_46
timestamp 1659098407
transform -1 0 1656 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  clk_rst_gen_47
timestamp 1659098407
transform 1 0 18492 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  clk_rst_gen_48
timestamp 1659098407
transform 1 0 23000 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  clk_rst_gen_49
timestamp 1659098407
transform 1 0 46828 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  clk_rst_gen_50
timestamp 1659098407
transform -1 0 33856 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  clk_rst_gen_51
timestamp 1659098407
transform -1 0 2300 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  clk_rst_gen_52
timestamp 1659098407
transform -1 0 35604 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  clk_rst_gen_53
timestamp 1659098407
transform 1 0 46644 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  clk_rst_gen_54
timestamp 1659098407
transform -1 0 42688 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  clk_rst_gen_55
timestamp 1659098407
transform -1 0 33856 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  clk_rst_gen_56
timestamp 1659098407
transform -1 0 1656 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  clk_rst_gen_57
timestamp 1659098407
transform -1 0 30636 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  clk_rst_gen_58
timestamp 1659098407
transform -1 0 2944 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  clk_rst_gen_59
timestamp 1659098407
transform -1 0 37720 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  clk_rst_gen_60
timestamp 1659098407
transform 1 0 5612 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  clk_rst_gen_61
timestamp 1659098407
transform 1 0 17848 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  clk_rst_gen_62
timestamp 1659098407
transform -1 0 1656 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  clk_rst_gen_63
timestamp 1659098407
transform -1 0 40940 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  clk_rst_gen_64
timestamp 1659098407
transform -1 0 1656 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  clk_rst_gen_65
timestamp 1659098407
transform 1 0 45540 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  clk_rst_gen_66
timestamp 1659098407
transform -1 0 39008 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  clk_rst_gen_67
timestamp 1659098407
transform -1 0 1656 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  clk_rst_gen_68
timestamp 1659098407
transform -1 0 17112 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  clk_rst_gen_69
timestamp 1659098407
transform 1 0 47932 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  clk_rst_gen_70
timestamp 1659098407
transform -1 0 24840 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  clk_rst_gen_71
timestamp 1659098407
transform -1 0 19688 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  clk_rst_gen_72
timestamp 1659098407
transform -1 0 1656 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  clk_rst_gen_73
timestamp 1659098407
transform -1 0 31096 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  clk_rst_gen_74
timestamp 1659098407
transform 1 0 47932 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  clk_rst_gen_75
timestamp 1659098407
transform 1 0 47932 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  clk_rst_gen_76
timestamp 1659098407
transform -1 0 2300 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  clk_rst_gen_77
timestamp 1659098407
transform -1 0 15180 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  clk_rst_gen_78
timestamp 1659098407
transform -1 0 40112 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  clk_rst_gen_79
timestamp 1659098407
transform -1 0 36432 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  clk_rst_gen_80
timestamp 1659098407
transform 1 0 17204 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  clk_rst_gen_81
timestamp 1659098407
transform 1 0 3036 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  clk_rst_gen_82
timestamp 1659098407
transform 1 0 46828 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  clk_rst_gen_83
timestamp 1659098407
transform 1 0 47932 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  clk_rst_gen_84
timestamp 1659098407
transform -1 0 13248 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  clk_rst_gen_85
timestamp 1659098407
transform 1 0 47932 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  clk_rst_gen_86
timestamp 1659098407
transform 1 0 5612 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  clk_rst_gen_87
timestamp 1659098407
transform -1 0 26128 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  clk_rst_gen_88
timestamp 1659098407
transform 1 0 47932 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  clk_rst_gen_89
timestamp 1659098407
transform -1 0 1656 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  clk_rst_gen_90
timestamp 1659098407
transform 1 0 10120 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  clk_rst_gen_91
timestamp 1659098407
transform -1 0 14352 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  clk_rst_gen_92
timestamp 1659098407
transform -1 0 43332 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  clk_rst_gen_93
timestamp 1659098407
transform -1 0 38824 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  clk_rst_gen_94
timestamp 1659098407
transform 1 0 47932 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  clk_rst_gen_95
timestamp 1659098407
transform -1 0 19688 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  clk_rst_gen_96
timestamp 1659098407
transform 1 0 21068 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  clk_rst_gen_97
timestamp 1659098407
transform 1 0 19780 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  clk_rst_gen_98
timestamp 1659098407
transform -1 0 1656 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  clk_rst_gen_99
timestamp 1659098407
transform 1 0 6900 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  clk_rst_gen_100
timestamp 1659098407
transform -1 0 1656 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  clk_rst_gen_101
timestamp 1659098407
transform 1 0 19780 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  clk_rst_gen_102
timestamp 1659098407
transform 1 0 7544 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  clk_rst_gen_103
timestamp 1659098407
transform -1 0 1656 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  clk_rst_gen_104
timestamp 1659098407
transform 1 0 4968 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  clk_rst_gen_105
timestamp 1659098407
transform 1 0 47932 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  clk_rst_gen_106
timestamp 1659098407
transform 1 0 47932 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  clk_rst_gen_107
timestamp 1659098407
transform -1 0 9384 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  clk_rst_gen_108
timestamp 1659098407
transform 1 0 47932 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  clk_rst_gen_109
timestamp 1659098407
transform -1 0 47840 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  clk_rst_gen_110
timestamp 1659098407
transform -1 0 24840 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  clk_rst_gen_111
timestamp 1659098407
transform 1 0 47288 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  clk_rst_gen_112
timestamp 1659098407
transform 1 0 10764 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  clk_rst_gen_113
timestamp 1659098407
transform -1 0 1656 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  clk_rst_gen_114
timestamp 1659098407
transform -1 0 29808 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  clk_rst_gen_115
timestamp 1659098407
transform -1 0 46736 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  clk_rst_gen_116
timestamp 1659098407
transform -1 0 1656 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  clk_rst_gen_117
timestamp 1659098407
transform -1 0 1656 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  clk_rst_gen_118
timestamp 1659098407
transform 1 0 47932 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  clk_rst_gen_119
timestamp 1659098407
transform -1 0 45448 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  clk_rst_gen_120
timestamp 1659098407
transform -1 0 41584 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  clk_rst_gen_121
timestamp 1659098407
transform -1 0 44160 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  clk_rst_gen_122
timestamp 1659098407
transform 1 0 2392 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  clk_rst_gen_123
timestamp 1659098407
transform 1 0 47932 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  clk_rst_gen_124
timestamp 1659098407
transform -1 0 37536 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  clk_rst_gen_125
timestamp 1659098407
transform 1 0 8188 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  clk_rst_gen_126
timestamp 1659098407
transform -1 0 15824 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  clk_rst_gen_127
timestamp 1659098407
transform -1 0 28704 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  clk_rst_gen_128
timestamp 1659098407
transform -1 0 1656 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  clk_rst_gen_129
timestamp 1659098407
transform -1 0 4232 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  clk_rst_gen_130
timestamp 1659098407
transform 1 0 47932 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  clk_rst_gen_131
timestamp 1659098407
transform -1 0 1656 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  clk_rst_gen_132
timestamp 1659098407
transform -1 0 1656 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  clk_rst_gen_133
timestamp 1659098407
transform -1 0 25484 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  clk_rst_gen_134
timestamp 1659098407
transform -1 0 2300 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  clk_rst_gen_135
timestamp 1659098407
transform -1 0 30452 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  clk_rst_gen_136
timestamp 1659098407
transform -1 0 1656 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  clk_rst_gen_137
timestamp 1659098407
transform 1 0 10120 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  clk_rst_gen_138
timestamp 1659098407
transform -1 0 26128 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  clk_rst_gen_139
timestamp 1659098407
transform -1 0 1656 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  clk_rst_gen_140
timestamp 1659098407
transform 1 0 7544 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  clk_rst_gen_141
timestamp 1659098407
transform -1 0 34960 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  clk_rst_gen_142
timestamp 1659098407
transform -1 0 25484 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  clk_rst_gen_143
timestamp 1659098407
transform 1 0 20424 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  clk_rst_gen_144
timestamp 1659098407
transform -1 0 40296 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  clk_rst_gen_145
timestamp 1659098407
transform 1 0 47932 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  clk_rst_gen_146
timestamp 1659098407
transform -1 0 2944 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  clk_rst_gen_147
timestamp 1659098407
transform 1 0 47932 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  clk_rst_gen_148
timestamp 1659098407
transform 1 0 8188 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  clk_rst_gen_149
timestamp 1659098407
transform -1 0 15180 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  clk_rst_gen_150
timestamp 1659098407
transform -1 0 1656 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  clk_rst_gen_151
timestamp 1659098407
transform -1 0 23552 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  clk_rst_gen_152
timestamp 1659098407
transform -1 0 38180 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  clk_rst_gen_154
timestamp 1659098407
transform 1 0 32292 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  clk_rst_gen_155
timestamp 1659098407
transform 1 0 2024 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  clk_rst_gen_156
timestamp 1659098407
transform 1 0 12328 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  clk_rst_gen_157
timestamp 1659098407
transform 1 0 1380 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  clk_rst_gen_158
timestamp 1659098407
transform 1 0 1380 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  clk_rst_gen_159
timestamp 1659098407
transform -1 0 7176 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  clk_rst_gen_160
timestamp 1659098407
transform 1 0 11684 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  clk_rst_gen_161
timestamp 1659098407
transform -1 0 48208 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  clk_rst_gen_162
timestamp 1659098407
transform 1 0 2668 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  clk_rst_gen_163
timestamp 1659098407
transform -1 0 9752 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  clk_rst_gen_164
timestamp 1659098407
transform 1 0 1380 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  clk_rst_gen_165
timestamp 1659098407
transform 1 0 29532 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  clk_rst_gen_166
timestamp 1659098407
transform 1 0 35972 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  clk_rst_gen_167
timestamp 1659098407
transform -1 0 4600 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  clk_rst_gen_168
timestamp 1659098407
transform 1 0 35328 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  clk_rst_gen_169
timestamp 1659098407
transform 1 0 1380 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  clk_rst_gen_170
timestamp 1659098407
transform 1 0 32936 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  clk_rst_gen_171
timestamp 1659098407
transform 1 0 40664 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  clk_rst_gen_172
timestamp 1659098407
transform 1 0 1380 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  clk_rst_gen_173
timestamp 1659098407
transform -1 0 47564 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  clk_rst_gen_174
timestamp 1659098407
transform 1 0 36156 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  clk_rst_gen_175
timestamp 1659098407
transform -1 0 48208 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  clk_rst_gen_176
timestamp 1659098407
transform -1 0 47104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  clk_rst_gen_177
timestamp 1659098407
transform 1 0 3956 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  clk_rst_gen_178
timestamp 1659098407
transform 1 0 35972 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  clk_rst_gen_179
timestamp 1659098407
transform 1 0 45632 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  clk_rst_gen_180
timestamp 1659098407
transform 1 0 11684 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  clk_rst_gen_181
timestamp 1659098407
transform 1 0 31004 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  clk_rst_gen_182
timestamp 1659098407
transform 1 0 47748 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  clk_rst_gen_183
timestamp 1659098407
transform 1 0 12972 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  clk_rst_gen_184
timestamp 1659098407
transform 1 0 28244 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  clk_rst_gen_185
timestamp 1659098407
transform 1 0 1380 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  clk_rst_gen_186
timestamp 1659098407
transform 1 0 16652 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  clk_rst_gen_187
timestamp 1659098407
transform 1 0 12328 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  clk_rst_gen_188
timestamp 1659098407
transform 1 0 47564 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  clk_rst_gen_189
timestamp 1659098407
transform -1 0 46460 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  clk_rst_gen_190
timestamp 1659098407
transform 1 0 27784 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  clk_rst_gen_191
timestamp 1659098407
transform -1 0 46920 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  clk_rst_gen_192
timestamp 1659098407
transform 1 0 1380 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  clk_rst_gen_193
timestamp 1659098407
transform -1 0 22632 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  clk_rst_gen_194
timestamp 1659098407
transform 1 0 27600 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  clk_rst_gen_195
timestamp 1659098407
transform 1 0 44988 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  clk_rst_gen_196
timestamp 1659098407
transform -1 0 23920 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  clk_rst_gen_197
timestamp 1659098407
transform 1 0 42412 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  clk_rst_gen_198
timestamp 1659098407
transform -1 0 21344 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  clk_rst_gen_199
timestamp 1659098407
transform 1 0 2668 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  clk_rst_gen_200
timestamp 1659098407
transform -1 0 48208 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  clk_rst_gen_201
timestamp 1659098407
transform 1 0 28428 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  clk_rst_gen_202
timestamp 1659098407
transform -1 0 47104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  clk_rst_gen_203
timestamp 1659098407
transform -1 0 9752 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  clk_rst_gen_204
timestamp 1659098407
transform 1 0 43700 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  clk_rst_gen_205
timestamp 1659098407
transform -1 0 16192 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk_i ../openroad/OpenLane/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1659098407
transform -1 0 34868 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_clk_i
timestamp 1659098407
transform -1 0 30452 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_clk_i
timestamp 1659098407
transform 1 0 33764 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold1 ../openroad/OpenLane/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1659098407
transform 1 0 27324 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold2
timestamp 1659098407
transform 1 0 32384 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold3
timestamp 1659098407
transform 1 0 42596 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold4
timestamp 1659098407
transform 1 0 38364 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input1 ../openroad/OpenLane/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1659098407
transform 1 0 42596 0 1 27200
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 1659098407
transform -1 0 45816 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1659098407
transform 1 0 47932 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output4
timestamp 1659098407
transform 1 0 21988 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output5
timestamp 1659098407
transform -1 0 23000 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output6
timestamp 1659098407
transform 1 0 47840 0 1 27200
box -38 -48 406 592
<< labels >>
flabel metal3 s 49200 14968 50000 15088 0 FreeSans 480 0 0 0 clk_i
port 0 nsew signal input
flabel metal2 s 21914 0 21970 800 0 FreeSans 224 90 0 0 clk_o
port 1 nsew signal tristate
flabel metal2 s 4526 29200 4582 30000 0 FreeSans 224 90 0 0 clk_sel_i
port 2 nsew signal input
flabel metal3 s 0 4088 800 4208 0 FreeSans 480 0 0 0 clk_standalone_i
port 3 nsew signal input
flabel metal2 s 22558 0 22614 800 0 FreeSans 224 90 0 0 fll_ack_o
port 4 nsew signal tristate
flabel metal3 s 49200 29248 50000 29368 0 FreeSans 480 0 0 0 fll_add_i[0]
port 5 nsew signal input
flabel metal2 s 48318 0 48374 800 0 FreeSans 224 90 0 0 fll_add_i[1]
port 6 nsew signal input
flabel metal2 s 16762 29200 16818 30000 0 FreeSans 224 90 0 0 fll_data_i[0]
port 7 nsew signal input
flabel metal3 s 0 9528 800 9648 0 FreeSans 480 0 0 0 fll_data_i[10]
port 8 nsew signal input
flabel metal2 s 3238 29200 3294 30000 0 FreeSans 224 90 0 0 fll_data_i[11]
port 9 nsew signal input
flabel metal3 s 49200 21088 50000 21208 0 FreeSans 480 0 0 0 fll_data_i[12]
port 10 nsew signal input
flabel metal2 s 39946 0 40002 800 0 FreeSans 224 90 0 0 fll_data_i[13]
port 11 nsew signal input
flabel metal2 s 32862 29200 32918 30000 0 FreeSans 224 90 0 0 fll_data_i[14]
port 12 nsew signal input
flabel metal2 s 14186 29200 14242 30000 0 FreeSans 224 90 0 0 fll_data_i[15]
port 13 nsew signal input
flabel metal3 s 49200 8168 50000 8288 0 FreeSans 480 0 0 0 fll_data_i[16]
port 14 nsew signal input
flabel metal2 s 6458 0 6514 800 0 FreeSans 224 90 0 0 fll_data_i[17]
port 15 nsew signal input
flabel metal3 s 0 10208 800 10328 0 FreeSans 480 0 0 0 fll_data_i[18]
port 16 nsew signal input
flabel metal2 s 31574 29200 31630 30000 0 FreeSans 224 90 0 0 fll_data_i[19]
port 17 nsew signal input
flabel metal2 s 27066 29200 27122 30000 0 FreeSans 224 90 0 0 fll_data_i[1]
port 18 nsew signal input
flabel metal3 s 0 17688 800 17808 0 FreeSans 480 0 0 0 fll_data_i[20]
port 19 nsew signal input
flabel metal3 s 49200 10208 50000 10328 0 FreeSans 480 0 0 0 fll_data_i[21]
port 20 nsew signal input
flabel metal2 s 1950 0 2006 800 0 FreeSans 224 90 0 0 fll_data_i[22]
port 21 nsew signal input
flabel metal3 s 0 16328 800 16448 0 FreeSans 480 0 0 0 fll_data_i[23]
port 22 nsew signal input
flabel metal3 s 49200 10888 50000 11008 0 FreeSans 480 0 0 0 fll_data_i[24]
port 23 nsew signal input
flabel metal2 s 39302 29200 39358 30000 0 FreeSans 224 90 0 0 fll_data_i[25]
port 24 nsew signal input
flabel metal2 s 45742 0 45798 800 0 FreeSans 224 90 0 0 fll_data_i[26]
port 25 nsew signal input
flabel metal2 s 44454 29200 44510 30000 0 FreeSans 224 90 0 0 fll_data_i[27]
port 26 nsew signal input
flabel metal2 s 2594 29200 2650 30000 0 FreeSans 224 90 0 0 fll_data_i[28]
port 27 nsew signal input
flabel metal3 s 0 12928 800 13048 0 FreeSans 480 0 0 0 fll_data_i[29]
port 28 nsew signal input
flabel metal2 s 14186 0 14242 800 0 FreeSans 224 90 0 0 fll_data_i[2]
port 29 nsew signal input
flabel metal3 s 0 2728 800 2848 0 FreeSans 480 0 0 0 fll_data_i[30]
port 30 nsew signal input
flabel metal3 s 49200 5448 50000 5568 0 FreeSans 480 0 0 0 fll_data_i[31]
port 31 nsew signal input
flabel metal2 s 17406 29200 17462 30000 0 FreeSans 224 90 0 0 fll_data_i[3]
port 32 nsew signal input
flabel metal3 s 0 26528 800 26648 0 FreeSans 480 0 0 0 fll_data_i[4]
port 33 nsew signal input
flabel metal3 s 0 17008 800 17128 0 FreeSans 480 0 0 0 fll_data_i[5]
port 34 nsew signal input
flabel metal2 s 36726 0 36782 800 0 FreeSans 224 90 0 0 fll_data_i[6]
port 35 nsew signal input
flabel metal3 s 0 22448 800 22568 0 FreeSans 480 0 0 0 fll_data_i[7]
port 36 nsew signal input
flabel metal2 s 29642 29200 29698 30000 0 FreeSans 224 90 0 0 fll_data_i[8]
port 37 nsew signal input
flabel metal2 s 31574 0 31630 800 0 FreeSans 224 90 0 0 fll_data_i[9]
port 38 nsew signal input
flabel metal3 s 0 14288 800 14408 0 FreeSans 480 0 0 0 fll_lock_o
port 39 nsew signal tristate
flabel metal3 s 49200 12248 50000 12368 0 FreeSans 480 0 0 0 fll_r_data_o[0]
port 40 nsew signal tristate
flabel metal2 s 34150 0 34206 800 0 FreeSans 224 90 0 0 fll_r_data_o[10]
port 41 nsew signal tristate
flabel metal2 s 5170 29200 5226 30000 0 FreeSans 224 90 0 0 fll_r_data_o[11]
port 42 nsew signal tristate
flabel metal2 s 30930 29200 30986 30000 0 FreeSans 224 90 0 0 fll_r_data_o[12]
port 43 nsew signal tristate
flabel metal3 s 49200 4768 50000 4888 0 FreeSans 480 0 0 0 fll_r_data_o[13]
port 44 nsew signal tristate
flabel metal3 s 49200 4088 50000 4208 0 FreeSans 480 0 0 0 fll_r_data_o[14]
port 45 nsew signal tristate
flabel metal3 s 49200 15648 50000 15768 0 FreeSans 480 0 0 0 fll_r_data_o[15]
port 46 nsew signal tristate
flabel metal3 s 0 12248 800 12368 0 FreeSans 480 0 0 0 fll_r_data_o[16]
port 47 nsew signal tristate
flabel metal2 s 46386 29200 46442 30000 0 FreeSans 224 90 0 0 fll_r_data_o[17]
port 48 nsew signal tristate
flabel metal2 s 13542 0 13598 800 0 FreeSans 224 90 0 0 fll_r_data_o[18]
port 49 nsew signal tristate
flabel metal3 s 49200 17008 50000 17128 0 FreeSans 480 0 0 0 fll_r_data_o[19]
port 50 nsew signal tristate
flabel metal2 s 26422 29200 26478 30000 0 FreeSans 224 90 0 0 fll_r_data_o[1]
port 51 nsew signal tristate
flabel metal2 s 18694 29200 18750 30000 0 FreeSans 224 90 0 0 fll_r_data_o[20]
port 52 nsew signal tristate
flabel metal2 s 6458 29200 6514 30000 0 FreeSans 224 90 0 0 fll_r_data_o[21]
port 53 nsew signal tristate
flabel metal2 s 9034 0 9090 800 0 FreeSans 224 90 0 0 fll_r_data_o[22]
port 54 nsew signal tristate
flabel metal2 s 43166 29200 43222 30000 0 FreeSans 224 90 0 0 fll_r_data_o[23]
port 55 nsew signal tristate
flabel metal3 s 0 8168 800 8288 0 FreeSans 480 0 0 0 fll_r_data_o[24]
port 56 nsew signal tristate
flabel metal3 s 0 4768 800 4888 0 FreeSans 480 0 0 0 fll_r_data_o[25]
port 57 nsew signal tristate
flabel metal3 s 49200 26528 50000 26648 0 FreeSans 480 0 0 0 fll_r_data_o[26]
port 58 nsew signal tristate
flabel metal2 s 1950 29200 2006 30000 0 FreeSans 224 90 0 0 fll_r_data_o[27]
port 59 nsew signal tristate
flabel metal2 s 41234 29200 41290 30000 0 FreeSans 224 90 0 0 fll_r_data_o[28]
port 60 nsew signal tristate
flabel metal2 s 20626 29200 20682 30000 0 FreeSans 224 90 0 0 fll_r_data_o[29]
port 61 nsew signal tristate
flabel metal3 s 49200 23808 50000 23928 0 FreeSans 480 0 0 0 fll_r_data_o[2]
port 62 nsew signal tristate
flabel metal2 s 32218 29200 32274 30000 0 FreeSans 224 90 0 0 fll_r_data_o[30]
port 63 nsew signal tristate
flabel metal3 s 49200 9528 50000 9648 0 FreeSans 480 0 0 0 fll_r_data_o[31]
port 64 nsew signal tristate
flabel metal3 s 0 3408 800 3528 0 FreeSans 480 0 0 0 fll_r_data_o[3]
port 65 nsew signal tristate
flabel metal2 s 23846 0 23902 800 0 FreeSans 224 90 0 0 fll_r_data_o[4]
port 66 nsew signal tristate
flabel metal2 s 38658 0 38714 800 0 FreeSans 224 90 0 0 fll_r_data_o[5]
port 67 nsew signal tristate
flabel metal3 s 49200 20408 50000 20528 0 FreeSans 480 0 0 0 fll_r_data_o[6]
port 68 nsew signal tristate
flabel metal2 s 10966 29200 11022 30000 0 FreeSans 224 90 0 0 fll_r_data_o[7]
port 69 nsew signal tristate
flabel metal2 s 26422 0 26478 800 0 FreeSans 224 90 0 0 fll_r_data_o[8]
port 70 nsew signal tristate
flabel metal2 s 18050 29200 18106 30000 0 FreeSans 224 90 0 0 fll_r_data_o[9]
port 71 nsew signal tristate
flabel metal2 s 42522 29200 42578 30000 0 FreeSans 224 90 0 0 fll_req_i
port 72 nsew signal input
flabel metal2 s 15474 0 15530 800 0 FreeSans 224 90 0 0 fll_wrn_i
port 73 nsew signal input
flabel metal2 s 32218 0 32274 800 0 FreeSans 224 90 0 0 io_oeb[0]
port 74 nsew signal tristate
flabel metal3 s 0 7488 800 7608 0 FreeSans 480 0 0 0 io_oeb[10]
port 75 nsew signal tristate
flabel metal2 s 28998 29200 29054 30000 0 FreeSans 224 90 0 0 io_oeb[11]
port 76 nsew signal tristate
flabel metal2 s 35438 29200 35494 30000 0 FreeSans 224 90 0 0 io_oeb[12]
port 77 nsew signal tristate
flabel metal2 s 4526 0 4582 800 0 FreeSans 224 90 0 0 io_oeb[13]
port 78 nsew signal tristate
flabel metal2 s 34794 29200 34850 30000 0 FreeSans 224 90 0 0 io_oeb[14]
port 79 nsew signal tristate
flabel metal3 s 0 6808 800 6928 0 FreeSans 480 0 0 0 io_oeb[15]
port 80 nsew signal tristate
flabel metal2 s 32862 0 32918 800 0 FreeSans 224 90 0 0 io_oeb[16]
port 81 nsew signal tristate
flabel metal2 s 40590 29200 40646 30000 0 FreeSans 224 90 0 0 io_oeb[17]
port 82 nsew signal tristate
flabel metal2 s 1306 29200 1362 30000 0 FreeSans 224 90 0 0 io_oeb[18]
port 83 nsew signal tristate
flabel metal2 s 49606 0 49662 800 0 FreeSans 224 90 0 0 io_oeb[19]
port 84 nsew signal tristate
flabel metal3 s 0 29248 800 29368 0 FreeSans 480 0 0 0 io_oeb[1]
port 85 nsew signal tristate
flabel metal2 s 36082 0 36138 800 0 FreeSans 224 90 0 0 io_oeb[20]
port 86 nsew signal tristate
flabel metal3 s 49200 25848 50000 25968 0 FreeSans 480 0 0 0 io_oeb[21]
port 87 nsew signal tristate
flabel metal3 s 49200 2728 50000 2848 0 FreeSans 480 0 0 0 io_oeb[22]
port 88 nsew signal tristate
flabel metal2 s 3882 0 3938 800 0 FreeSans 224 90 0 0 io_oeb[23]
port 89 nsew signal tristate
flabel metal2 s 35438 0 35494 800 0 FreeSans 224 90 0 0 io_oeb[24]
port 90 nsew signal tristate
flabel metal2 s 45098 0 45154 800 0 FreeSans 224 90 0 0 io_oeb[25]
port 91 nsew signal tristate
flabel metal2 s 21914 29200 21970 30000 0 FreeSans 224 90 0 0 io_oeb[26]
port 92 nsew signal tristate
flabel metal2 s 43810 0 43866 800 0 FreeSans 224 90 0 0 io_oeb[27]
port 93 nsew signal tristate
flabel metal3 s 49200 11568 50000 11688 0 FreeSans 480 0 0 0 io_oeb[28]
port 94 nsew signal tristate
flabel metal2 s 45742 29200 45798 30000 0 FreeSans 224 90 0 0 io_oeb[29]
port 95 nsew signal tristate
flabel metal2 s 12254 0 12310 800 0 FreeSans 224 90 0 0 io_oeb[2]
port 96 nsew signal tristate
flabel metal3 s 49200 688 50000 808 0 FreeSans 480 0 0 0 io_oeb[30]
port 97 nsew signal tristate
flabel metal3 s 0 1368 800 1488 0 FreeSans 480 0 0 0 io_oeb[31]
port 98 nsew signal tristate
flabel metal3 s 0 18368 800 18488 0 FreeSans 480 0 0 0 io_oeb[32]
port 99 nsew signal tristate
flabel metal2 s 18694 0 18750 800 0 FreeSans 224 90 0 0 io_oeb[33]
port 100 nsew signal tristate
flabel metal2 s 23202 29200 23258 30000 0 FreeSans 224 90 0 0 io_oeb[34]
port 101 nsew signal tristate
flabel metal2 s 47674 29200 47730 30000 0 FreeSans 224 90 0 0 io_oeb[35]
port 102 nsew signal tristate
flabel metal2 s 33506 29200 33562 30000 0 FreeSans 224 90 0 0 io_oeb[36]
port 103 nsew signal tristate
flabel metal3 s 0 2048 800 2168 0 FreeSans 480 0 0 0 io_oeb[37]
port 104 nsew signal tristate
flabel metal3 s 0 6128 800 6248 0 FreeSans 480 0 0 0 io_oeb[3]
port 105 nsew signal tristate
flabel metal3 s 0 23808 800 23928 0 FreeSans 480 0 0 0 io_oeb[4]
port 106 nsew signal tristate
flabel metal2 s 7102 29200 7158 30000 0 FreeSans 224 90 0 0 io_oeb[5]
port 107 nsew signal tristate
flabel metal2 s 11610 0 11666 800 0 FreeSans 224 90 0 0 io_oeb[6]
port 108 nsew signal tristate
flabel metal3 s 49200 6808 50000 6928 0 FreeSans 480 0 0 0 io_oeb[7]
port 109 nsew signal tristate
flabel metal2 s 662 29200 718 30000 0 FreeSans 224 90 0 0 io_oeb[8]
port 110 nsew signal tristate
flabel metal2 s 9678 0 9734 800 0 FreeSans 224 90 0 0 io_oeb[9]
port 111 nsew signal tristate
flabel metal2 s 11610 29200 11666 30000 0 FreeSans 224 90 0 0 io_out[0]
port 112 nsew signal tristate
flabel metal2 s 27710 29200 27766 30000 0 FreeSans 224 90 0 0 io_out[10]
port 113 nsew signal tristate
flabel metal3 s 49200 27208 50000 27328 0 FreeSans 480 0 0 0 io_out[11]
port 114 nsew signal tristate
flabel metal3 s 0 11568 800 11688 0 FreeSans 480 0 0 0 io_out[12]
port 115 nsew signal tristate
flabel metal2 s 22558 29200 22614 30000 0 FreeSans 224 90 0 0 io_out[13]
port 116 nsew signal tristate
flabel metal2 s 27066 0 27122 800 0 FreeSans 224 90 0 0 io_out[14]
port 117 nsew signal tristate
flabel metal2 s 44454 0 44510 800 0 FreeSans 224 90 0 0 io_out[15]
port 118 nsew signal tristate
flabel metal2 s 23846 29200 23902 30000 0 FreeSans 224 90 0 0 io_out[16]
port 119 nsew signal tristate
flabel metal2 s 41878 0 41934 800 0 FreeSans 224 90 0 0 io_out[17]
port 120 nsew signal tristate
flabel metal2 s 21270 0 21326 800 0 FreeSans 224 90 0 0 io_out[18]
port 121 nsew signal tristate
flabel metal3 s 0 8 800 128 0 FreeSans 480 0 0 0 io_out[19]
port 122 nsew signal tristate
flabel metal2 s 30930 0 30986 800 0 FreeSans 224 90 0 0 io_out[1]
port 123 nsew signal tristate
flabel metal3 s 49200 18368 50000 18488 0 FreeSans 480 0 0 0 io_out[20]
port 124 nsew signal tristate
flabel metal2 s 28354 29200 28410 30000 0 FreeSans 224 90 0 0 io_out[21]
port 125 nsew signal tristate
flabel metal2 s 49606 29200 49662 30000 0 FreeSans 224 90 0 0 io_out[22]
port 126 nsew signal tristate
flabel metal2 s 9678 29200 9734 30000 0 FreeSans 224 90 0 0 io_out[23]
port 127 nsew signal tristate
flabel metal2 s 43166 0 43222 800 0 FreeSans 224 90 0 0 io_out[24]
port 128 nsew signal tristate
flabel metal2 s 16118 0 16174 800 0 FreeSans 224 90 0 0 io_out[25]
port 129 nsew signal tristate
flabel metal2 s 47674 0 47730 800 0 FreeSans 224 90 0 0 io_out[2]
port 130 nsew signal tristate
flabel metal2 s 12898 29200 12954 30000 0 FreeSans 224 90 0 0 io_out[3]
port 131 nsew signal tristate
flabel metal2 s 27710 0 27766 800 0 FreeSans 224 90 0 0 io_out[4]
port 132 nsew signal tristate
flabel metal3 s 0 10888 800 11008 0 FreeSans 480 0 0 0 io_out[5]
port 133 nsew signal tristate
flabel metal2 s 16118 29200 16174 30000 0 FreeSans 224 90 0 0 io_out[6]
port 134 nsew signal tristate
flabel metal2 s 12254 29200 12310 30000 0 FreeSans 224 90 0 0 io_out[7]
port 135 nsew signal tristate
flabel metal2 s 47030 29200 47086 30000 0 FreeSans 224 90 0 0 io_out[8]
port 136 nsew signal tristate
flabel metal2 s 48962 29200 49018 30000 0 FreeSans 224 90 0 0 io_out[9]
port 137 nsew signal tristate
flabel metal2 s 34794 0 34850 800 0 FreeSans 224 90 0 0 la_data_out[0]
port 138 nsew signal tristate
flabel metal3 s 0 21088 800 21208 0 FreeSans 480 0 0 0 la_data_out[10]
port 139 nsew signal tristate
flabel metal2 s 40590 0 40646 800 0 FreeSans 224 90 0 0 la_data_out[11]
port 140 nsew signal tristate
flabel metal3 s 0 23128 800 23248 0 FreeSans 480 0 0 0 la_data_out[12]
port 141 nsew signal tristate
flabel metal3 s 49200 28568 50000 28688 0 FreeSans 480 0 0 0 la_data_out[13]
port 142 nsew signal tristate
flabel metal2 s 38658 29200 38714 30000 0 FreeSans 224 90 0 0 la_data_out[14]
port 143 nsew signal tristate
flabel metal3 s 0 25168 800 25288 0 FreeSans 480 0 0 0 la_data_out[15]
port 144 nsew signal tristate
flabel metal2 s 16762 0 16818 800 0 FreeSans 224 90 0 0 la_data_out[16]
port 145 nsew signal tristate
flabel metal3 s 49200 3408 50000 3528 0 FreeSans 480 0 0 0 la_data_out[17]
port 146 nsew signal tristate
flabel metal2 s 24490 29200 24546 30000 0 FreeSans 224 90 0 0 la_data_out[18]
port 147 nsew signal tristate
flabel metal2 s 19338 0 19394 800 0 FreeSans 224 90 0 0 la_data_out[19]
port 148 nsew signal tristate
flabel metal3 s 49200 8 50000 128 0 FreeSans 480 0 0 0 la_data_out[1]
port 149 nsew signal tristate
flabel metal3 s 0 21768 800 21888 0 FreeSans 480 0 0 0 la_data_out[20]
port 150 nsew signal tristate
flabel metal2 s 30286 0 30342 800 0 FreeSans 224 90 0 0 la_data_out[21]
port 151 nsew signal tristate
flabel metal3 s 49200 25168 50000 25288 0 FreeSans 480 0 0 0 la_data_out[22]
port 152 nsew signal tristate
flabel metal3 s 49200 16328 50000 16448 0 FreeSans 480 0 0 0 la_data_out[23]
port 153 nsew signal tristate
flabel metal3 s 0 28568 800 28688 0 FreeSans 480 0 0 0 la_data_out[24]
port 154 nsew signal tristate
flabel metal2 s 14830 29200 14886 30000 0 FreeSans 224 90 0 0 la_data_out[25]
port 155 nsew signal tristate
flabel metal2 s 39302 0 39358 800 0 FreeSans 224 90 0 0 la_data_out[26]
port 156 nsew signal tristate
flabel metal2 s 36082 29200 36138 30000 0 FreeSans 224 90 0 0 la_data_out[27]
port 157 nsew signal tristate
flabel metal2 s 17406 0 17462 800 0 FreeSans 224 90 0 0 la_data_out[28]
port 158 nsew signal tristate
flabel metal2 s 3238 0 3294 800 0 FreeSans 224 90 0 0 la_data_out[29]
port 159 nsew signal tristate
flabel metal2 s 41878 29200 41934 30000 0 FreeSans 224 90 0 0 la_data_out[2]
port 160 nsew signal tristate
flabel metal3 s 49200 1368 50000 1488 0 FreeSans 480 0 0 0 la_data_out[30]
port 161 nsew signal tristate
flabel metal3 s 49200 14288 50000 14408 0 FreeSans 480 0 0 0 la_data_out[31]
port 162 nsew signal tristate
flabel metal2 s 12898 0 12954 800 0 FreeSans 224 90 0 0 la_data_out[32]
port 163 nsew signal tristate
flabel metal3 s 49200 23128 50000 23248 0 FreeSans 480 0 0 0 la_data_out[33]
port 164 nsew signal tristate
flabel metal2 s 5814 29200 5870 30000 0 FreeSans 224 90 0 0 la_data_out[34]
port 165 nsew signal tristate
flabel metal2 s 25778 0 25834 800 0 FreeSans 224 90 0 0 la_data_out[35]
port 166 nsew signal tristate
flabel metal3 s 49200 24488 50000 24608 0 FreeSans 480 0 0 0 la_data_out[36]
port 167 nsew signal tristate
flabel metal3 s 0 19728 800 19848 0 FreeSans 480 0 0 0 la_data_out[37]
port 168 nsew signal tristate
flabel metal2 s 10322 0 10378 800 0 FreeSans 224 90 0 0 la_data_out[38]
port 169 nsew signal tristate
flabel metal2 s 13542 29200 13598 30000 0 FreeSans 224 90 0 0 la_data_out[39]
port 170 nsew signal tristate
flabel metal2 s 33506 0 33562 800 0 FreeSans 224 90 0 0 la_data_out[3]
port 171 nsew signal tristate
flabel metal2 s 42522 0 42578 800 0 FreeSans 224 90 0 0 la_data_out[40]
port 172 nsew signal tristate
flabel metal2 s 38014 29200 38070 30000 0 FreeSans 224 90 0 0 la_data_out[41]
port 173 nsew signal tristate
flabel metal3 s 49200 13608 50000 13728 0 FreeSans 480 0 0 0 la_data_out[42]
port 174 nsew signal tristate
flabel metal2 s 19338 29200 19394 30000 0 FreeSans 224 90 0 0 la_data_out[43]
port 175 nsew signal tristate
flabel metal2 s 21270 29200 21326 30000 0 FreeSans 224 90 0 0 la_data_out[44]
port 176 nsew signal tristate
flabel metal2 s 19982 29200 20038 30000 0 FreeSans 224 90 0 0 la_data_out[45]
port 177 nsew signal tristate
flabel metal2 s 1306 0 1362 800 0 FreeSans 224 90 0 0 la_data_out[46]
port 178 nsew signal tristate
flabel metal2 s 7102 0 7158 800 0 FreeSans 224 90 0 0 la_data_out[47]
port 179 nsew signal tristate
flabel metal3 s 0 27888 800 28008 0 FreeSans 480 0 0 0 la_data_out[48]
port 180 nsew signal tristate
flabel metal2 s 19982 0 20038 800 0 FreeSans 224 90 0 0 la_data_out[49]
port 181 nsew signal tristate
flabel metal3 s 0 27208 800 27328 0 FreeSans 480 0 0 0 la_data_out[4]
port 182 nsew signal tristate
flabel metal2 s 7746 29200 7802 30000 0 FreeSans 224 90 0 0 la_data_out[50]
port 183 nsew signal tristate
flabel metal3 s 0 15648 800 15768 0 FreeSans 480 0 0 0 la_data_out[51]
port 184 nsew signal tristate
flabel metal2 s 5170 0 5226 800 0 FreeSans 224 90 0 0 la_data_out[52]
port 185 nsew signal tristate
flabel metal3 s 49200 6128 50000 6248 0 FreeSans 480 0 0 0 la_data_out[53]
port 186 nsew signal tristate
flabel metal3 s 49200 22448 50000 22568 0 FreeSans 480 0 0 0 la_data_out[54]
port 187 nsew signal tristate
flabel metal2 s 9034 29200 9090 30000 0 FreeSans 224 90 0 0 la_data_out[55]
port 188 nsew signal tristate
flabel metal3 s 49200 12928 50000 13048 0 FreeSans 480 0 0 0 la_data_out[56]
port 189 nsew signal tristate
flabel metal2 s 47030 0 47086 800 0 FreeSans 224 90 0 0 la_data_out[57]
port 190 nsew signal tristate
flabel metal2 s 24490 0 24546 800 0 FreeSans 224 90 0 0 la_data_out[58]
port 191 nsew signal tristate
flabel metal3 s 49200 27888 50000 28008 0 FreeSans 480 0 0 0 la_data_out[59]
port 192 nsew signal tristate
flabel metal2 s 30286 29200 30342 30000 0 FreeSans 224 90 0 0 la_data_out[5]
port 193 nsew signal tristate
flabel metal2 s 10966 0 11022 800 0 FreeSans 224 90 0 0 la_data_out[60]
port 194 nsew signal tristate
flabel metal3 s 0 24488 800 24608 0 FreeSans 480 0 0 0 la_data_out[61]
port 195 nsew signal tristate
flabel metal2 s 28998 0 29054 800 0 FreeSans 224 90 0 0 la_data_out[62]
port 196 nsew signal tristate
flabel metal2 s 46386 0 46442 800 0 FreeSans 224 90 0 0 la_data_out[63]
port 197 nsew signal tristate
flabel metal3 s 0 688 800 808 0 FreeSans 480 0 0 0 la_data_out[6]
port 198 nsew signal tristate
flabel metal2 s 37370 0 37426 800 0 FreeSans 224 90 0 0 la_data_out[7]
port 199 nsew signal tristate
flabel metal2 s 5814 0 5870 800 0 FreeSans 224 90 0 0 la_data_out[8]
port 200 nsew signal tristate
flabel metal2 s 18050 0 18106 800 0 FreeSans 224 90 0 0 la_data_out[9]
port 201 nsew signal tristate
flabel metal3 s 49200 2048 50000 2168 0 FreeSans 480 0 0 0 rstn_i
port 202 nsew signal input
flabel metal2 s 48318 29200 48374 30000 0 FreeSans 224 90 0 0 rstn_o
port 203 nsew signal tristate
flabel metal3 s 49200 19728 50000 19848 0 FreeSans 480 0 0 0 scan_en_i
port 204 nsew signal input
flabel metal2 s 38014 0 38070 800 0 FreeSans 224 90 0 0 scan_i
port 205 nsew signal input
flabel metal3 s 0 13608 800 13728 0 FreeSans 480 0 0 0 scan_o
port 206 nsew signal tristate
flabel metal3 s 49200 7488 50000 7608 0 FreeSans 480 0 0 0 testmode_i
port 207 nsew signal input
flabel metal2 s 662 0 718 800 0 FreeSans 224 90 0 0 user_irq[0]
port 208 nsew signal tristate
flabel metal3 s 49200 21768 50000 21888 0 FreeSans 480 0 0 0 user_irq[1]
port 209 nsew signal tristate
flabel metal2 s 45098 29200 45154 30000 0 FreeSans 224 90 0 0 user_irq[2]
port 210 nsew signal tristate
flabel metal4 s 6918 2128 7238 27792 0 FreeSans 1920 90 0 0 vccd1
port 211 nsew power bidirectional
flabel metal4 s 18866 2128 19186 27792 0 FreeSans 1920 90 0 0 vccd1
port 211 nsew power bidirectional
flabel metal4 s 30814 2128 31134 27792 0 FreeSans 1920 90 0 0 vccd1
port 211 nsew power bidirectional
flabel metal4 s 42762 2128 43082 27792 0 FreeSans 1920 90 0 0 vccd1
port 211 nsew power bidirectional
flabel metal4 s 12892 2128 13212 27792 0 FreeSans 1920 90 0 0 vssd1
port 212 nsew ground bidirectional
flabel metal4 s 24840 2128 25160 27792 0 FreeSans 1920 90 0 0 vssd1
port 212 nsew ground bidirectional
flabel metal4 s 36788 2128 37108 27792 0 FreeSans 1920 90 0 0 vssd1
port 212 nsew ground bidirectional
flabel metal2 s 41234 0 41290 800 0 FreeSans 224 90 0 0 wbs_ack_o
port 213 nsew signal tristate
flabel metal2 s 43810 29200 43866 30000 0 FreeSans 224 90 0 0 wbs_dat_o[0]
port 214 nsew signal tristate
flabel metal3 s 0 14968 800 15088 0 FreeSans 480 0 0 0 wbs_dat_o[10]
port 215 nsew signal tristate
flabel metal3 s 0 20408 800 20528 0 FreeSans 480 0 0 0 wbs_dat_o[11]
port 216 nsew signal tristate
flabel metal2 s 25134 0 25190 800 0 FreeSans 224 90 0 0 wbs_dat_o[12]
port 217 nsew signal tristate
flabel metal2 s 18 0 74 800 0 FreeSans 224 90 0 0 wbs_dat_o[13]
port 218 nsew signal tristate
flabel metal2 s 29642 0 29698 800 0 FreeSans 224 90 0 0 wbs_dat_o[14]
port 219 nsew signal tristate
flabel metal3 s 0 25848 800 25968 0 FreeSans 480 0 0 0 wbs_dat_o[15]
port 220 nsew signal tristate
flabel metal2 s 10322 29200 10378 30000 0 FreeSans 224 90 0 0 wbs_dat_o[16]
port 221 nsew signal tristate
flabel metal2 s 25778 29200 25834 30000 0 FreeSans 224 90 0 0 wbs_dat_o[17]
port 222 nsew signal tristate
flabel metal3 s 0 19048 800 19168 0 FreeSans 480 0 0 0 wbs_dat_o[18]
port 223 nsew signal tristate
flabel metal2 s 7746 0 7802 800 0 FreeSans 224 90 0 0 wbs_dat_o[19]
port 224 nsew signal tristate
flabel metal2 s 2594 0 2650 800 0 FreeSans 224 90 0 0 wbs_dat_o[1]
port 225 nsew signal tristate
flabel metal2 s 34150 29200 34206 30000 0 FreeSans 224 90 0 0 wbs_dat_o[20]
port 226 nsew signal tristate
flabel metal2 s 25134 29200 25190 30000 0 FreeSans 224 90 0 0 wbs_dat_o[21]
port 227 nsew signal tristate
flabel metal2 s 20626 0 20682 800 0 FreeSans 224 90 0 0 wbs_dat_o[22]
port 228 nsew signal tristate
flabel metal2 s 39946 29200 40002 30000 0 FreeSans 224 90 0 0 wbs_dat_o[23]
port 229 nsew signal tristate
flabel metal2 s 48962 0 49018 800 0 FreeSans 224 90 0 0 wbs_dat_o[24]
port 230 nsew signal tristate
flabel metal2 s 18 29200 74 30000 0 FreeSans 224 90 0 0 wbs_dat_o[25]
port 231 nsew signal tristate
flabel metal3 s 49200 19048 50000 19168 0 FreeSans 480 0 0 0 wbs_dat_o[26]
port 232 nsew signal tristate
flabel metal2 s 8390 0 8446 800 0 FreeSans 224 90 0 0 wbs_dat_o[27]
port 233 nsew signal tristate
flabel metal2 s 14830 0 14886 800 0 FreeSans 224 90 0 0 wbs_dat_o[28]
port 234 nsew signal tristate
flabel metal3 s 0 5448 800 5568 0 FreeSans 480 0 0 0 wbs_dat_o[29]
port 235 nsew signal tristate
flabel metal3 s 49200 17688 50000 17808 0 FreeSans 480 0 0 0 wbs_dat_o[2]
port 236 nsew signal tristate
flabel metal2 s 23202 0 23258 800 0 FreeSans 224 90 0 0 wbs_dat_o[30]
port 237 nsew signal tristate
flabel metal2 s 37370 29200 37426 30000 0 FreeSans 224 90 0 0 wbs_dat_o[31]
port 238 nsew signal tristate
flabel metal2 s 36726 29200 36782 30000 0 FreeSans 224 90 0 0 wbs_dat_o[3]
port 239 nsew signal tristate
flabel metal2 s 8390 29200 8446 30000 0 FreeSans 224 90 0 0 wbs_dat_o[4]
port 240 nsew signal tristate
flabel metal2 s 15474 29200 15530 30000 0 FreeSans 224 90 0 0 wbs_dat_o[5]
port 241 nsew signal tristate
flabel metal2 s 28354 0 28410 800 0 FreeSans 224 90 0 0 wbs_dat_o[6]
port 242 nsew signal tristate
flabel metal3 s 0 8848 800 8968 0 FreeSans 480 0 0 0 wbs_dat_o[7]
port 243 nsew signal tristate
flabel metal2 s 3882 29200 3938 30000 0 FreeSans 224 90 0 0 wbs_dat_o[8]
port 244 nsew signal tristate
flabel metal3 s 49200 8848 50000 8968 0 FreeSans 480 0 0 0 wbs_dat_o[9]
port 245 nsew signal tristate
<< properties >>
string FIXED_BBOX 0 0 50000 30000
<< end >>
