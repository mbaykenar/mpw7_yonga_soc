magic
tech sky130A
magscale 1 2
timestamp 1649977179
<< nwell >>
rect -66 377 834 897
<< pwell >>
rect 13 43 764 283
rect -26 -43 794 43
<< mvnmos >>
rect 101 173 201 257
rect 243 173 343 257
rect 385 173 485 257
rect 585 107 685 257
<< mvpmos >>
rect 87 517 187 601
rect 243 517 343 601
rect 399 517 499 601
rect 578 443 678 743
<< mvndiff >>
rect 39 232 101 257
rect 39 198 51 232
rect 85 198 101 232
rect 39 173 101 198
rect 201 173 243 257
rect 343 173 385 257
rect 485 249 585 257
rect 485 215 540 249
rect 574 215 585 249
rect 485 173 585 215
rect 528 149 585 173
rect 528 115 540 149
rect 574 115 585 149
rect 528 107 585 115
rect 685 245 738 257
rect 685 211 696 245
rect 730 211 738 245
rect 685 153 738 211
rect 685 119 696 153
rect 730 119 738 153
rect 685 107 738 119
<< mvpdiff >>
rect 521 735 578 743
rect 521 701 533 735
rect 567 701 578 735
rect 521 652 578 701
rect 521 618 533 652
rect 567 618 578 652
rect 521 601 578 618
rect 30 576 87 601
rect 30 542 42 576
rect 76 542 87 576
rect 30 517 87 542
rect 187 580 243 601
rect 187 546 198 580
rect 232 546 243 580
rect 187 517 243 546
rect 343 576 399 601
rect 343 542 354 576
rect 388 542 399 576
rect 343 517 399 542
rect 499 568 578 601
rect 499 534 533 568
rect 567 534 578 568
rect 499 517 578 534
rect 521 485 578 517
rect 521 451 533 485
rect 567 451 578 485
rect 521 443 578 451
rect 678 735 735 743
rect 678 701 689 735
rect 723 701 735 735
rect 678 652 735 701
rect 678 618 689 652
rect 723 618 735 652
rect 678 568 735 618
rect 678 534 689 568
rect 723 534 735 568
rect 678 485 735 534
rect 678 451 689 485
rect 723 451 735 485
rect 678 443 735 451
<< mvndiffc >>
rect 51 198 85 232
rect 540 215 574 249
rect 540 115 574 149
rect 696 211 730 245
rect 696 119 730 153
<< mvpdiffc >>
rect 533 701 567 735
rect 533 618 567 652
rect 42 542 76 576
rect 198 546 232 580
rect 354 542 388 576
rect 533 534 567 568
rect 533 451 567 485
rect 689 701 723 735
rect 689 618 723 652
rect 689 534 723 568
rect 689 451 723 485
<< mvpsubdiff >>
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 768 17
<< mvnsubdiff >>
rect 0 797 31 831
rect 65 797 127 831
rect 161 797 223 831
rect 257 797 319 831
rect 353 797 415 831
rect 449 797 511 831
rect 545 797 607 831
rect 641 797 703 831
rect 737 797 768 831
<< mvpsubdiffcont >>
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
<< mvnsubdiffcont >>
rect 31 797 65 831
rect 127 797 161 831
rect 223 797 257 831
rect 319 797 353 831
rect 415 797 449 831
rect 511 797 545 831
rect 607 797 641 831
rect 703 797 737 831
<< poly >>
rect 578 743 678 769
rect 87 601 187 627
rect 243 601 343 627
rect 399 601 499 627
rect 87 379 187 517
rect 243 469 343 517
rect 243 435 263 469
rect 297 435 343 469
rect 87 329 201 379
rect 87 295 137 329
rect 171 295 201 329
rect 87 279 201 295
rect 101 257 201 279
rect 243 257 343 435
rect 399 379 499 517
rect 385 329 499 379
rect 385 295 401 329
rect 435 295 499 329
rect 385 279 499 295
rect 578 417 678 443
rect 578 383 685 417
rect 578 349 598 383
rect 632 349 685 383
rect 578 283 685 349
rect 385 257 485 279
rect 585 257 685 283
rect 101 147 201 173
rect 243 147 343 173
rect 385 147 485 173
rect 585 81 685 107
<< polycont >>
rect 263 435 297 469
rect 137 295 171 329
rect 401 295 435 329
rect 598 349 632 383
<< locali >>
rect 0 797 31 831
rect 65 797 127 831
rect 161 797 223 831
rect 257 797 319 831
rect 353 797 415 831
rect 449 797 511 831
rect 545 797 607 831
rect 641 797 703 831
rect 737 797 768 831
rect 112 735 302 741
rect 112 701 118 735
rect 152 701 190 735
rect 224 701 262 735
rect 296 701 302 735
rect 26 576 76 609
rect 26 542 42 576
rect 26 399 76 542
rect 112 580 302 701
rect 440 735 630 751
rect 440 701 446 735
rect 480 701 518 735
rect 567 701 590 735
rect 624 701 630 735
rect 440 652 630 701
rect 440 618 533 652
rect 567 618 630 652
rect 112 546 198 580
rect 232 546 302 580
rect 112 534 302 546
rect 354 576 404 609
rect 388 542 404 576
rect 121 469 313 498
rect 121 435 263 469
rect 297 435 313 469
rect 354 399 404 542
rect 440 568 630 618
rect 440 534 533 568
rect 567 534 630 568
rect 440 485 630 534
rect 440 451 533 485
rect 567 451 630 485
rect 440 435 630 451
rect 673 735 743 751
rect 673 701 689 735
rect 723 701 743 735
rect 673 652 743 701
rect 673 618 689 652
rect 723 618 743 652
rect 673 568 743 618
rect 673 534 689 568
rect 723 534 743 568
rect 673 485 743 534
rect 673 451 689 485
rect 723 451 743 485
rect 673 435 743 451
rect 26 383 648 399
rect 26 365 598 383
rect 26 232 85 365
rect 582 349 598 365
rect 632 349 648 383
rect 582 333 648 349
rect 26 198 51 232
rect 26 165 85 198
rect 121 295 137 329
rect 171 295 187 329
rect 121 162 187 295
rect 223 295 401 329
rect 435 295 451 329
rect 223 162 451 295
rect 487 249 648 265
rect 487 215 540 249
rect 574 215 648 249
rect 487 149 648 215
rect 487 115 540 149
rect 574 115 648 149
rect 487 113 648 115
rect 487 79 497 113
rect 531 79 603 113
rect 637 79 648 113
rect 682 245 743 435
rect 682 211 696 245
rect 730 211 743 245
rect 682 153 743 211
rect 682 119 696 153
rect 730 119 743 153
rect 682 99 743 119
rect 487 73 648 79
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 768 17
<< viali >>
rect 31 797 65 831
rect 127 797 161 831
rect 223 797 257 831
rect 319 797 353 831
rect 415 797 449 831
rect 511 797 545 831
rect 607 797 641 831
rect 703 797 737 831
rect 118 701 152 735
rect 190 701 224 735
rect 262 701 296 735
rect 446 701 480 735
rect 518 701 533 735
rect 533 701 552 735
rect 590 701 624 735
rect 497 79 531 113
rect 603 79 637 113
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
<< metal1 >>
rect 0 831 768 837
rect 0 797 31 831
rect 65 797 127 831
rect 161 797 223 831
rect 257 797 319 831
rect 353 797 415 831
rect 449 797 511 831
rect 545 797 607 831
rect 641 797 703 831
rect 737 797 768 831
rect 0 791 768 797
rect 0 735 768 763
rect 0 701 118 735
rect 152 701 190 735
rect 224 701 262 735
rect 296 701 446 735
rect 480 701 518 735
rect 552 701 590 735
rect 624 701 768 735
rect 0 689 768 701
rect 0 113 768 125
rect 0 79 497 113
rect 531 79 603 113
rect 637 79 768 113
rect 0 51 768 79
rect 0 17 768 23
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 768 17
rect 0 -23 768 -17
<< labels >>
rlabel comment s 0 0 0 0 4 and3_1
flabel metal1 s 0 51 768 125 0 FreeSans 340 0 0 0 VGND
port 4 nsew ground bidirectional
flabel metal1 s 0 0 768 23 0 FreeSans 340 0 0 0 VNB
port 5 nsew ground bidirectional
flabel metal1 s 0 689 768 763 0 FreeSans 340 0 0 0 VPWR
port 7 nsew power bidirectional
flabel metal1 s 0 791 768 814 0 FreeSans 340 0 0 0 VPB
port 6 nsew power bidirectional
flabel locali s 127 168 161 202 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 127 242 161 276 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 127 464 161 498 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 223 464 257 498 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 223 168 257 202 0 FreeSans 340 0 0 0 C
port 3 nsew signal input
flabel locali s 223 242 257 276 0 FreeSans 340 0 0 0 C
port 3 nsew signal input
flabel locali s 319 168 353 202 0 FreeSans 340 0 0 0 C
port 3 nsew signal input
flabel locali s 319 242 353 276 0 FreeSans 340 0 0 0 C
port 3 nsew signal input
flabel locali s 415 168 449 202 0 FreeSans 340 0 0 0 C
port 3 nsew signal input
flabel locali s 415 242 449 276 0 FreeSans 340 0 0 0 C
port 3 nsew signal input
flabel locali s 703 168 737 202 0 FreeSans 340 0 0 0 X
port 8 nsew signal output
flabel locali s 703 242 737 276 0 FreeSans 340 0 0 0 X
port 8 nsew signal output
flabel locali s 703 316 737 350 0 FreeSans 340 0 0 0 X
port 8 nsew signal output
flabel locali s 703 390 737 424 0 FreeSans 340 0 0 0 X
port 8 nsew signal output
flabel locali s 703 464 737 498 0 FreeSans 340 0 0 0 X
port 8 nsew signal output
flabel locali s 703 538 737 572 0 FreeSans 340 0 0 0 X
port 8 nsew signal output
flabel locali s 703 612 737 646 0 FreeSans 340 0 0 0 X
port 8 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 768 814
string GDS_END 813630
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hvl/gds/sky130_fd_sc_hvl.gds
string GDS_START 803460
string LEFclass CORE
string LEFsite unithv
string LEFsymmetry X Y
<< end >>
