magic
tech sky130B
magscale 1 2
timestamp 1649977179
<< dnwell >>
rect -2476 -1400 2776 7401
<< nwell >>
rect -10 0 310 6000
<< pwell >>
rect -1102 -26 -374 6026
rect 674 -26 1402 6026
<< obsactive >>
rect -2676 -1600 2976 7601
<< locali >>
rect -1068 5969 -934 5991
rect -1068 31 -1054 5969
rect -948 31 -934 5969
rect -1068 9 -934 31
rect -830 5969 -696 5991
rect -830 31 -816 5969
rect -710 31 -696 5969
rect 996 5969 1130 5991
rect 15 5933 285 5957
rect 15 67 25 5933
rect 275 67 285 5933
rect 15 43 285 67
rect -830 9 -696 31
rect 996 31 1010 5969
rect 1116 31 1130 5969
rect 996 9 1130 31
rect 1234 5969 1368 5991
rect 1234 31 1248 5969
rect 1354 31 1368 5969
rect 1234 9 1368 31
rect -209 -459 555 -443
rect -209 -493 -180 -459
rect -146 -493 -106 -459
rect -72 -493 -32 -459
rect 2 -493 42 -459
rect 76 -493 116 -459
rect 150 -493 190 -459
rect 224 -493 264 -459
rect 298 -493 338 -459
rect 372 -493 412 -459
rect 446 -493 486 -459
rect 520 -493 555 -459
rect -209 -533 555 -493
rect -209 -567 -180 -533
rect -146 -567 -106 -533
rect -72 -567 -32 -533
rect 2 -567 42 -533
rect 76 -567 116 -533
rect 150 -567 190 -533
rect 224 -567 264 -533
rect 298 -567 338 -533
rect 372 -567 412 -533
rect 446 -567 486 -533
rect 520 -567 555 -533
rect -209 -607 555 -567
rect -209 -641 -180 -607
rect -146 -641 -106 -607
rect -72 -641 -32 -607
rect 2 -641 42 -607
rect 76 -641 116 -607
rect 150 -641 190 -607
rect 224 -641 264 -607
rect 298 -641 338 -607
rect 372 -641 412 -607
rect 446 -641 486 -607
rect 520 -641 555 -607
rect -209 -657 555 -641
<< viali >>
rect -1054 31 -948 5969
rect -816 31 -710 5969
rect 25 67 275 5933
rect 1010 31 1116 5969
rect 1248 31 1354 5969
rect -180 -493 -146 -459
rect -106 -493 -72 -459
rect -32 -493 2 -459
rect 42 -493 76 -459
rect 116 -493 150 -459
rect 190 -493 224 -459
rect 264 -493 298 -459
rect 338 -493 372 -459
rect 412 -493 446 -459
rect 486 -493 520 -459
rect -180 -567 -146 -533
rect -106 -567 -72 -533
rect -32 -567 2 -533
rect 42 -567 76 -533
rect 116 -567 150 -533
rect 190 -567 224 -533
rect 264 -567 298 -533
rect 338 -567 372 -533
rect 412 -567 446 -533
rect 486 -567 520 -533
rect -180 -641 -146 -607
rect -106 -641 -72 -607
rect -32 -641 2 -607
rect 42 -641 76 -607
rect 116 -641 150 -607
rect 190 -641 224 -607
rect 264 -641 298 -607
rect 338 -641 372 -607
rect 412 -641 446 -607
rect 486 -641 520 -607
<< metal1 >>
rect -1066 5969 -936 5981
rect -1066 31 -1054 5969
rect -948 31 -936 5969
rect -1066 19 -936 31
rect -828 5969 -698 5981
rect -828 31 -816 5969
rect -710 31 -698 5969
rect 998 5969 1128 5981
rect 13 5939 287 5945
rect 13 5933 28 5939
rect 272 5933 287 5939
rect 13 67 25 5933
rect 275 67 287 5933
rect 13 63 28 67
rect 272 63 287 67
rect 13 55 287 63
rect -828 19 -698 31
rect 998 31 1010 5969
rect 1116 31 1128 5969
rect 998 19 1128 31
rect 1236 5969 1366 5981
rect 1236 31 1248 5969
rect 1354 31 1366 5969
rect 1236 19 1366 31
rect -209 -450 555 -443
rect -209 -502 -189 -450
rect -137 -502 -115 -450
rect -63 -502 -41 -450
rect 11 -502 33 -450
rect 85 -502 107 -450
rect 159 -502 181 -450
rect 233 -502 255 -450
rect 307 -502 329 -450
rect 381 -502 403 -450
rect 455 -502 477 -450
rect 529 -502 555 -450
rect -209 -524 555 -502
rect -209 -576 -189 -524
rect -137 -576 -115 -524
rect -63 -576 -41 -524
rect 11 -576 33 -524
rect 85 -576 107 -524
rect 159 -576 181 -524
rect 233 -576 255 -524
rect 307 -576 329 -524
rect 381 -576 403 -524
rect 455 -576 477 -524
rect 529 -576 555 -524
rect -209 -598 555 -576
rect -209 -650 -189 -598
rect -137 -650 -115 -598
rect -63 -650 -41 -598
rect 11 -650 33 -598
rect 85 -650 107 -598
rect 159 -650 181 -598
rect 233 -650 255 -598
rect 307 -650 329 -598
rect 381 -650 403 -598
rect 455 -650 477 -598
rect 529 -650 555 -598
rect -209 -657 555 -650
<< via1 >>
rect 28 5933 272 5939
rect 28 67 272 5933
rect 28 63 272 67
rect -189 -459 -137 -450
rect -189 -493 -180 -459
rect -180 -493 -146 -459
rect -146 -493 -137 -459
rect -189 -502 -137 -493
rect -115 -459 -63 -450
rect -115 -493 -106 -459
rect -106 -493 -72 -459
rect -72 -493 -63 -459
rect -115 -502 -63 -493
rect -41 -459 11 -450
rect -41 -493 -32 -459
rect -32 -493 2 -459
rect 2 -493 11 -459
rect -41 -502 11 -493
rect 33 -459 85 -450
rect 33 -493 42 -459
rect 42 -493 76 -459
rect 76 -493 85 -459
rect 33 -502 85 -493
rect 107 -459 159 -450
rect 107 -493 116 -459
rect 116 -493 150 -459
rect 150 -493 159 -459
rect 107 -502 159 -493
rect 181 -459 233 -450
rect 181 -493 190 -459
rect 190 -493 224 -459
rect 224 -493 233 -459
rect 181 -502 233 -493
rect 255 -459 307 -450
rect 255 -493 264 -459
rect 264 -493 298 -459
rect 298 -493 307 -459
rect 255 -502 307 -493
rect 329 -459 381 -450
rect 329 -493 338 -459
rect 338 -493 372 -459
rect 372 -493 381 -459
rect 329 -502 381 -493
rect 403 -459 455 -450
rect 403 -493 412 -459
rect 412 -493 446 -459
rect 446 -493 455 -459
rect 403 -502 455 -493
rect 477 -459 529 -450
rect 477 -493 486 -459
rect 486 -493 520 -459
rect 520 -493 529 -459
rect 477 -502 529 -493
rect -189 -533 -137 -524
rect -189 -567 -180 -533
rect -180 -567 -146 -533
rect -146 -567 -137 -533
rect -189 -576 -137 -567
rect -115 -533 -63 -524
rect -115 -567 -106 -533
rect -106 -567 -72 -533
rect -72 -567 -63 -533
rect -115 -576 -63 -567
rect -41 -533 11 -524
rect -41 -567 -32 -533
rect -32 -567 2 -533
rect 2 -567 11 -533
rect -41 -576 11 -567
rect 33 -533 85 -524
rect 33 -567 42 -533
rect 42 -567 76 -533
rect 76 -567 85 -533
rect 33 -576 85 -567
rect 107 -533 159 -524
rect 107 -567 116 -533
rect 116 -567 150 -533
rect 150 -567 159 -533
rect 107 -576 159 -567
rect 181 -533 233 -524
rect 181 -567 190 -533
rect 190 -567 224 -533
rect 224 -567 233 -533
rect 181 -576 233 -567
rect 255 -533 307 -524
rect 255 -567 264 -533
rect 264 -567 298 -533
rect 298 -567 307 -533
rect 255 -576 307 -567
rect 329 -533 381 -524
rect 329 -567 338 -533
rect 338 -567 372 -533
rect 372 -567 381 -533
rect 329 -576 381 -567
rect 403 -533 455 -524
rect 403 -567 412 -533
rect 412 -567 446 -533
rect 446 -567 455 -533
rect 403 -576 455 -567
rect 477 -533 529 -524
rect 477 -567 486 -533
rect 486 -567 520 -533
rect 520 -567 529 -533
rect 477 -576 529 -567
rect -189 -607 -137 -598
rect -189 -641 -180 -607
rect -180 -641 -146 -607
rect -146 -641 -137 -607
rect -189 -650 -137 -641
rect -115 -607 -63 -598
rect -115 -641 -106 -607
rect -106 -641 -72 -607
rect -72 -641 -63 -607
rect -115 -650 -63 -641
rect -41 -607 11 -598
rect -41 -641 -32 -607
rect -32 -641 2 -607
rect 2 -641 11 -607
rect -41 -650 11 -641
rect 33 -607 85 -598
rect 33 -641 42 -607
rect 42 -641 76 -607
rect 76 -641 85 -607
rect 33 -650 85 -641
rect 107 -607 159 -598
rect 107 -641 116 -607
rect 116 -641 150 -607
rect 150 -641 159 -607
rect 107 -650 159 -641
rect 181 -607 233 -598
rect 181 -641 190 -607
rect 190 -641 224 -607
rect 224 -641 233 -607
rect 181 -650 233 -641
rect 255 -607 307 -598
rect 255 -641 264 -607
rect 264 -641 298 -607
rect 298 -641 307 -607
rect 255 -650 307 -641
rect 329 -607 381 -598
rect 329 -641 338 -607
rect 338 -641 372 -607
rect 372 -641 381 -607
rect 329 -650 381 -641
rect 403 -607 455 -598
rect 403 -641 412 -607
rect 412 -641 446 -607
rect 446 -641 455 -607
rect 403 -650 455 -641
rect 477 -607 529 -598
rect 477 -641 486 -607
rect 486 -641 520 -607
rect 520 -641 529 -607
rect 477 -650 529 -641
<< metal2 >>
rect 22 5939 278 5945
rect 22 63 28 5939
rect 272 63 278 5939
rect 22 57 278 63
rect -209 -450 555 -443
rect -209 -502 -189 -450
rect -137 -502 -115 -450
rect -63 -502 -41 -450
rect 11 -502 33 -450
rect 85 -502 107 -450
rect 159 -502 181 -450
rect 233 -502 255 -450
rect 307 -502 329 -450
rect 381 -502 403 -450
rect 455 -502 477 -450
rect 529 -502 555 -450
rect -209 -524 555 -502
rect -209 -576 -189 -524
rect -137 -576 -115 -524
rect -63 -576 -41 -524
rect 11 -576 33 -524
rect 85 -576 107 -524
rect 159 -576 181 -524
rect 233 -576 255 -524
rect 307 -576 329 -524
rect 381 -576 403 -524
rect 455 -576 477 -524
rect 529 -576 555 -524
rect -209 -598 555 -576
rect -209 -650 -189 -598
rect -137 -650 -115 -598
rect -63 -650 -41 -598
rect 11 -650 33 -598
rect 85 -650 107 -598
rect 159 -650 181 -598
rect 233 -650 255 -598
rect 307 -650 329 -598
rect 381 -650 403 -598
rect 455 -650 477 -598
rect 529 -650 555 -598
rect -209 -657 555 -650
<< properties >>
string GDS_END 8388676
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_pr/gds/sky130_fd_pr.gds
string GDS_START 8207760
<< end >>
