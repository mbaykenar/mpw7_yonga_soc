magic
tech sky130B
magscale 12 1
timestamp 1598776399
<< metal5 >>
rect 0 75 30 105
rect 0 45 30 60
rect 15 -15 30 45
rect 0 -25 30 -15
rect 0 -30 25 -25
<< properties >>
string FIXED_BBOX 0 -30 45 105
<< end >>
