magic
tech sky130B
magscale 12 1
timestamp 1598786533
<< metal5 >>
rect 30 90 45 105
rect 20 80 55 90
rect 5 65 70 80
rect 20 55 55 65
rect 30 40 45 55
<< properties >>
string FIXED_BBOX 0 -30 90 105
<< end >>
