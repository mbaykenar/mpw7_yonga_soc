magic
tech sky130A
magscale 1 2
timestamp 1649977179
<< labels >>
rlabel poly s 75 74 75 74 4 G
port 1 nsew
rlabel mvpsubdiff s 25 74 25 74 4 S
rlabel mvpsubdiff s 125 74 125 74 4 D
<< properties >>
string GDS_END 106906
string GDS_FILE $PDKPATH/libs.ref/sky130_sram_macros/gds/sky130_sram_2kbyte_1rw1r_32x512_8.gds
string GDS_START 106258
<< end >>
