magic
tech sky130B
magscale 1 2
timestamp 1649977179
<< metal4 >>
rect 0 39976 254 40000
rect 15746 39976 16000 40000
rect 0 39965 16000 39976
rect 0 39729 162 39965
rect 398 39729 483 39965
rect 719 39729 804 39965
rect 1040 39729 1125 39965
rect 1361 39729 1446 39965
rect 1682 39729 1767 39965
rect 2003 39729 2088 39965
rect 2324 39729 2409 39965
rect 2645 39729 2730 39965
rect 2966 39729 3051 39965
rect 3287 39729 3372 39965
rect 3608 39729 3693 39965
rect 3929 39729 4014 39965
rect 4250 39729 4335 39965
rect 4571 39729 4656 39965
rect 4892 39729 4977 39965
rect 5213 39729 5298 39965
rect 5534 39729 5619 39965
rect 5855 39729 5940 39965
rect 6176 39729 6261 39965
rect 6497 39729 6582 39965
rect 6818 39729 6903 39965
rect 7139 39729 7224 39965
rect 7460 39729 7545 39965
rect 7781 39729 7866 39965
rect 8102 39729 8187 39965
rect 8423 39729 8508 39965
rect 8744 39729 8829 39965
rect 9065 39729 9150 39965
rect 9386 39729 9471 39965
rect 9707 39729 9792 39965
rect 10028 39729 10113 39965
rect 10349 39729 10434 39965
rect 10670 39729 10755 39965
rect 10991 39729 11076 39965
rect 11312 39729 11397 39965
rect 11633 39729 11718 39965
rect 11954 39729 12038 39965
rect 12274 39729 12358 39965
rect 12594 39729 12678 39965
rect 12914 39729 12998 39965
rect 13234 39729 13318 39965
rect 13554 39729 13638 39965
rect 13874 39729 13958 39965
rect 14194 39729 14278 39965
rect 14514 39729 14598 39965
rect 14834 39729 14918 39965
rect 15154 39729 15238 39965
rect 15474 39729 15558 39965
rect 15794 39729 16000 39965
rect 0 39641 16000 39729
rect 0 39405 162 39641
rect 398 39405 483 39641
rect 719 39405 804 39641
rect 1040 39405 1125 39641
rect 1361 39405 1446 39641
rect 1682 39405 1767 39641
rect 2003 39405 2088 39641
rect 2324 39405 2409 39641
rect 2645 39405 2730 39641
rect 2966 39405 3051 39641
rect 3287 39405 3372 39641
rect 3608 39405 3693 39641
rect 3929 39405 4014 39641
rect 4250 39405 4335 39641
rect 4571 39405 4656 39641
rect 4892 39405 4977 39641
rect 5213 39405 5298 39641
rect 5534 39405 5619 39641
rect 5855 39405 5940 39641
rect 6176 39405 6261 39641
rect 6497 39405 6582 39641
rect 6818 39405 6903 39641
rect 7139 39405 7224 39641
rect 7460 39405 7545 39641
rect 7781 39405 7866 39641
rect 8102 39405 8187 39641
rect 8423 39405 8508 39641
rect 8744 39405 8829 39641
rect 9065 39405 9150 39641
rect 9386 39405 9471 39641
rect 9707 39405 9792 39641
rect 10028 39405 10113 39641
rect 10349 39405 10434 39641
rect 10670 39405 10755 39641
rect 10991 39405 11076 39641
rect 11312 39405 11397 39641
rect 11633 39405 11718 39641
rect 11954 39405 12038 39641
rect 12274 39405 12358 39641
rect 12594 39405 12678 39641
rect 12914 39405 12998 39641
rect 13234 39405 13318 39641
rect 13554 39405 13638 39641
rect 13874 39405 13958 39641
rect 14194 39405 14278 39641
rect 14514 39405 14598 39641
rect 14834 39405 14918 39641
rect 15154 39405 15238 39641
rect 15474 39405 15558 39641
rect 15794 39405 16000 39641
rect 0 39317 16000 39405
rect 0 39081 162 39317
rect 398 39081 483 39317
rect 719 39081 804 39317
rect 1040 39081 1125 39317
rect 1361 39081 1446 39317
rect 1682 39081 1767 39317
rect 2003 39081 2088 39317
rect 2324 39081 2409 39317
rect 2645 39081 2730 39317
rect 2966 39081 3051 39317
rect 3287 39081 3372 39317
rect 3608 39081 3693 39317
rect 3929 39081 4014 39317
rect 4250 39081 4335 39317
rect 4571 39081 4656 39317
rect 4892 39081 4977 39317
rect 5213 39081 5298 39317
rect 5534 39081 5619 39317
rect 5855 39081 5940 39317
rect 6176 39081 6261 39317
rect 6497 39081 6582 39317
rect 6818 39081 6903 39317
rect 7139 39081 7224 39317
rect 7460 39081 7545 39317
rect 7781 39081 7866 39317
rect 8102 39081 8187 39317
rect 8423 39081 8508 39317
rect 8744 39081 8829 39317
rect 9065 39081 9150 39317
rect 9386 39081 9471 39317
rect 9707 39081 9792 39317
rect 10028 39081 10113 39317
rect 10349 39081 10434 39317
rect 10670 39081 10755 39317
rect 10991 39081 11076 39317
rect 11312 39081 11397 39317
rect 11633 39081 11718 39317
rect 11954 39081 12038 39317
rect 12274 39081 12358 39317
rect 12594 39081 12678 39317
rect 12914 39081 12998 39317
rect 13234 39081 13318 39317
rect 13554 39081 13638 39317
rect 13874 39081 13958 39317
rect 14194 39081 14278 39317
rect 14514 39081 14598 39317
rect 14834 39081 14918 39317
rect 15154 39081 15238 39317
rect 15474 39081 15558 39317
rect 15794 39081 16000 39317
rect 0 38993 16000 39081
rect 0 38757 162 38993
rect 398 38757 483 38993
rect 719 38757 804 38993
rect 1040 38757 1125 38993
rect 1361 38757 1446 38993
rect 1682 38757 1767 38993
rect 2003 38757 2088 38993
rect 2324 38757 2409 38993
rect 2645 38757 2730 38993
rect 2966 38757 3051 38993
rect 3287 38757 3372 38993
rect 3608 38757 3693 38993
rect 3929 38757 4014 38993
rect 4250 38757 4335 38993
rect 4571 38757 4656 38993
rect 4892 38757 4977 38993
rect 5213 38757 5298 38993
rect 5534 38757 5619 38993
rect 5855 38757 5940 38993
rect 6176 38757 6261 38993
rect 6497 38757 6582 38993
rect 6818 38757 6903 38993
rect 7139 38757 7224 38993
rect 7460 38757 7545 38993
rect 7781 38757 7866 38993
rect 8102 38757 8187 38993
rect 8423 38757 8508 38993
rect 8744 38757 8829 38993
rect 9065 38757 9150 38993
rect 9386 38757 9471 38993
rect 9707 38757 9792 38993
rect 10028 38757 10113 38993
rect 10349 38757 10434 38993
rect 10670 38757 10755 38993
rect 10991 38757 11076 38993
rect 11312 38757 11397 38993
rect 11633 38757 11718 38993
rect 11954 38757 12038 38993
rect 12274 38757 12358 38993
rect 12594 38757 12678 38993
rect 12914 38757 12998 38993
rect 13234 38757 13318 38993
rect 13554 38757 13638 38993
rect 13874 38757 13958 38993
rect 14194 38757 14278 38993
rect 14514 38757 14598 38993
rect 14834 38757 14918 38993
rect 15154 38757 15238 38993
rect 15474 38757 15558 38993
rect 15794 38757 16000 38993
rect 0 38669 16000 38757
rect 0 38433 162 38669
rect 398 38433 483 38669
rect 719 38433 804 38669
rect 1040 38433 1125 38669
rect 1361 38433 1446 38669
rect 1682 38433 1767 38669
rect 2003 38433 2088 38669
rect 2324 38433 2409 38669
rect 2645 38433 2730 38669
rect 2966 38433 3051 38669
rect 3287 38433 3372 38669
rect 3608 38433 3693 38669
rect 3929 38433 4014 38669
rect 4250 38433 4335 38669
rect 4571 38433 4656 38669
rect 4892 38433 4977 38669
rect 5213 38433 5298 38669
rect 5534 38433 5619 38669
rect 5855 38433 5940 38669
rect 6176 38433 6261 38669
rect 6497 38433 6582 38669
rect 6818 38433 6903 38669
rect 7139 38433 7224 38669
rect 7460 38433 7545 38669
rect 7781 38433 7866 38669
rect 8102 38433 8187 38669
rect 8423 38433 8508 38669
rect 8744 38433 8829 38669
rect 9065 38433 9150 38669
rect 9386 38433 9471 38669
rect 9707 38433 9792 38669
rect 10028 38433 10113 38669
rect 10349 38433 10434 38669
rect 10670 38433 10755 38669
rect 10991 38433 11076 38669
rect 11312 38433 11397 38669
rect 11633 38433 11718 38669
rect 11954 38433 12038 38669
rect 12274 38433 12358 38669
rect 12594 38433 12678 38669
rect 12914 38433 12998 38669
rect 13234 38433 13318 38669
rect 13554 38433 13638 38669
rect 13874 38433 13958 38669
rect 14194 38433 14278 38669
rect 14514 38433 14598 38669
rect 14834 38433 14918 38669
rect 15154 38433 15238 38669
rect 15474 38433 15558 38669
rect 15794 38433 16000 38669
rect 0 38345 16000 38433
rect 0 38109 162 38345
rect 398 38109 483 38345
rect 719 38109 804 38345
rect 1040 38109 1125 38345
rect 1361 38109 1446 38345
rect 1682 38109 1767 38345
rect 2003 38109 2088 38345
rect 2324 38109 2409 38345
rect 2645 38109 2730 38345
rect 2966 38109 3051 38345
rect 3287 38109 3372 38345
rect 3608 38109 3693 38345
rect 3929 38109 4014 38345
rect 4250 38109 4335 38345
rect 4571 38109 4656 38345
rect 4892 38109 4977 38345
rect 5213 38109 5298 38345
rect 5534 38109 5619 38345
rect 5855 38109 5940 38345
rect 6176 38109 6261 38345
rect 6497 38109 6582 38345
rect 6818 38109 6903 38345
rect 7139 38109 7224 38345
rect 7460 38109 7545 38345
rect 7781 38109 7866 38345
rect 8102 38109 8187 38345
rect 8423 38109 8508 38345
rect 8744 38109 8829 38345
rect 9065 38109 9150 38345
rect 9386 38109 9471 38345
rect 9707 38109 9792 38345
rect 10028 38109 10113 38345
rect 10349 38109 10434 38345
rect 10670 38109 10755 38345
rect 10991 38109 11076 38345
rect 11312 38109 11397 38345
rect 11633 38109 11718 38345
rect 11954 38109 12038 38345
rect 12274 38109 12358 38345
rect 12594 38109 12678 38345
rect 12914 38109 12998 38345
rect 13234 38109 13318 38345
rect 13554 38109 13638 38345
rect 13874 38109 13958 38345
rect 14194 38109 14278 38345
rect 14514 38109 14598 38345
rect 14834 38109 14918 38345
rect 15154 38109 15238 38345
rect 15474 38109 15558 38345
rect 15794 38109 16000 38345
rect 0 38021 16000 38109
rect 0 37785 162 38021
rect 398 37785 483 38021
rect 719 37785 804 38021
rect 1040 37785 1125 38021
rect 1361 37785 1446 38021
rect 1682 37785 1767 38021
rect 2003 37785 2088 38021
rect 2324 37785 2409 38021
rect 2645 37785 2730 38021
rect 2966 37785 3051 38021
rect 3287 37785 3372 38021
rect 3608 37785 3693 38021
rect 3929 37785 4014 38021
rect 4250 37785 4335 38021
rect 4571 37785 4656 38021
rect 4892 37785 4977 38021
rect 5213 37785 5298 38021
rect 5534 37785 5619 38021
rect 5855 37785 5940 38021
rect 6176 37785 6261 38021
rect 6497 37785 6582 38021
rect 6818 37785 6903 38021
rect 7139 37785 7224 38021
rect 7460 37785 7545 38021
rect 7781 37785 7866 38021
rect 8102 37785 8187 38021
rect 8423 37785 8508 38021
rect 8744 37785 8829 38021
rect 9065 37785 9150 38021
rect 9386 37785 9471 38021
rect 9707 37785 9792 38021
rect 10028 37785 10113 38021
rect 10349 37785 10434 38021
rect 10670 37785 10755 38021
rect 10991 37785 11076 38021
rect 11312 37785 11397 38021
rect 11633 37785 11718 38021
rect 11954 37785 12038 38021
rect 12274 37785 12358 38021
rect 12594 37785 12678 38021
rect 12914 37785 12998 38021
rect 13234 37785 13318 38021
rect 13554 37785 13638 38021
rect 13874 37785 13958 38021
rect 14194 37785 14278 38021
rect 14514 37785 14598 38021
rect 14834 37785 14918 38021
rect 15154 37785 15238 38021
rect 15474 37785 15558 38021
rect 15794 37785 16000 38021
rect 0 37697 16000 37785
rect 0 37461 162 37697
rect 398 37461 483 37697
rect 719 37461 804 37697
rect 1040 37461 1125 37697
rect 1361 37461 1446 37697
rect 1682 37461 1767 37697
rect 2003 37461 2088 37697
rect 2324 37461 2409 37697
rect 2645 37461 2730 37697
rect 2966 37461 3051 37697
rect 3287 37461 3372 37697
rect 3608 37461 3693 37697
rect 3929 37461 4014 37697
rect 4250 37461 4335 37697
rect 4571 37461 4656 37697
rect 4892 37461 4977 37697
rect 5213 37461 5298 37697
rect 5534 37461 5619 37697
rect 5855 37461 5940 37697
rect 6176 37461 6261 37697
rect 6497 37461 6582 37697
rect 6818 37461 6903 37697
rect 7139 37461 7224 37697
rect 7460 37461 7545 37697
rect 7781 37461 7866 37697
rect 8102 37461 8187 37697
rect 8423 37461 8508 37697
rect 8744 37461 8829 37697
rect 9065 37461 9150 37697
rect 9386 37461 9471 37697
rect 9707 37461 9792 37697
rect 10028 37461 10113 37697
rect 10349 37461 10434 37697
rect 10670 37461 10755 37697
rect 10991 37461 11076 37697
rect 11312 37461 11397 37697
rect 11633 37461 11718 37697
rect 11954 37461 12038 37697
rect 12274 37461 12358 37697
rect 12594 37461 12678 37697
rect 12914 37461 12998 37697
rect 13234 37461 13318 37697
rect 13554 37461 13638 37697
rect 13874 37461 13958 37697
rect 14194 37461 14278 37697
rect 14514 37461 14598 37697
rect 14834 37461 14918 37697
rect 15154 37461 15238 37697
rect 15474 37461 15558 37697
rect 15794 37461 16000 37697
rect 0 37373 16000 37461
rect 0 37137 162 37373
rect 398 37137 483 37373
rect 719 37137 804 37373
rect 1040 37137 1125 37373
rect 1361 37137 1446 37373
rect 1682 37137 1767 37373
rect 2003 37137 2088 37373
rect 2324 37137 2409 37373
rect 2645 37137 2730 37373
rect 2966 37137 3051 37373
rect 3287 37137 3372 37373
rect 3608 37137 3693 37373
rect 3929 37137 4014 37373
rect 4250 37137 4335 37373
rect 4571 37137 4656 37373
rect 4892 37137 4977 37373
rect 5213 37137 5298 37373
rect 5534 37137 5619 37373
rect 5855 37137 5940 37373
rect 6176 37137 6261 37373
rect 6497 37137 6582 37373
rect 6818 37137 6903 37373
rect 7139 37137 7224 37373
rect 7460 37137 7545 37373
rect 7781 37137 7866 37373
rect 8102 37137 8187 37373
rect 8423 37137 8508 37373
rect 8744 37137 8829 37373
rect 9065 37137 9150 37373
rect 9386 37137 9471 37373
rect 9707 37137 9792 37373
rect 10028 37137 10113 37373
rect 10349 37137 10434 37373
rect 10670 37137 10755 37373
rect 10991 37137 11076 37373
rect 11312 37137 11397 37373
rect 11633 37137 11718 37373
rect 11954 37137 12038 37373
rect 12274 37137 12358 37373
rect 12594 37137 12678 37373
rect 12914 37137 12998 37373
rect 13234 37137 13318 37373
rect 13554 37137 13638 37373
rect 13874 37137 13958 37373
rect 14194 37137 14278 37373
rect 14514 37137 14598 37373
rect 14834 37137 14918 37373
rect 15154 37137 15238 37373
rect 15474 37137 15558 37373
rect 15794 37137 16000 37373
rect 0 37049 16000 37137
rect 0 36813 162 37049
rect 398 36813 483 37049
rect 719 36813 804 37049
rect 1040 36813 1125 37049
rect 1361 36813 1446 37049
rect 1682 36813 1767 37049
rect 2003 36813 2088 37049
rect 2324 36813 2409 37049
rect 2645 36813 2730 37049
rect 2966 36813 3051 37049
rect 3287 36813 3372 37049
rect 3608 36813 3693 37049
rect 3929 36813 4014 37049
rect 4250 36813 4335 37049
rect 4571 36813 4656 37049
rect 4892 36813 4977 37049
rect 5213 36813 5298 37049
rect 5534 36813 5619 37049
rect 5855 36813 5940 37049
rect 6176 36813 6261 37049
rect 6497 36813 6582 37049
rect 6818 36813 6903 37049
rect 7139 36813 7224 37049
rect 7460 36813 7545 37049
rect 7781 36813 7866 37049
rect 8102 36813 8187 37049
rect 8423 36813 8508 37049
rect 8744 36813 8829 37049
rect 9065 36813 9150 37049
rect 9386 36813 9471 37049
rect 9707 36813 9792 37049
rect 10028 36813 10113 37049
rect 10349 36813 10434 37049
rect 10670 36813 10755 37049
rect 10991 36813 11076 37049
rect 11312 36813 11397 37049
rect 11633 36813 11718 37049
rect 11954 36813 12038 37049
rect 12274 36813 12358 37049
rect 12594 36813 12678 37049
rect 12914 36813 12998 37049
rect 13234 36813 13318 37049
rect 13554 36813 13638 37049
rect 13874 36813 13958 37049
rect 14194 36813 14278 37049
rect 14514 36813 14598 37049
rect 14834 36813 14918 37049
rect 15154 36813 15238 37049
rect 15474 36813 15558 37049
rect 15794 36813 16000 37049
rect 0 36725 16000 36813
rect 0 36489 162 36725
rect 398 36489 483 36725
rect 719 36489 804 36725
rect 1040 36489 1125 36725
rect 1361 36489 1446 36725
rect 1682 36489 1767 36725
rect 2003 36489 2088 36725
rect 2324 36489 2409 36725
rect 2645 36489 2730 36725
rect 2966 36489 3051 36725
rect 3287 36489 3372 36725
rect 3608 36489 3693 36725
rect 3929 36489 4014 36725
rect 4250 36489 4335 36725
rect 4571 36489 4656 36725
rect 4892 36489 4977 36725
rect 5213 36489 5298 36725
rect 5534 36489 5619 36725
rect 5855 36489 5940 36725
rect 6176 36489 6261 36725
rect 6497 36489 6582 36725
rect 6818 36489 6903 36725
rect 7139 36489 7224 36725
rect 7460 36489 7545 36725
rect 7781 36489 7866 36725
rect 8102 36489 8187 36725
rect 8423 36489 8508 36725
rect 8744 36489 8829 36725
rect 9065 36489 9150 36725
rect 9386 36489 9471 36725
rect 9707 36489 9792 36725
rect 10028 36489 10113 36725
rect 10349 36489 10434 36725
rect 10670 36489 10755 36725
rect 10991 36489 11076 36725
rect 11312 36489 11397 36725
rect 11633 36489 11718 36725
rect 11954 36489 12038 36725
rect 12274 36489 12358 36725
rect 12594 36489 12678 36725
rect 12914 36489 12998 36725
rect 13234 36489 13318 36725
rect 13554 36489 13638 36725
rect 13874 36489 13958 36725
rect 14194 36489 14278 36725
rect 14514 36489 14598 36725
rect 14834 36489 14918 36725
rect 15154 36489 15238 36725
rect 15474 36489 15558 36725
rect 15794 36489 16000 36725
rect 0 36401 16000 36489
rect 0 36165 162 36401
rect 398 36165 483 36401
rect 719 36165 804 36401
rect 1040 36165 1125 36401
rect 1361 36165 1446 36401
rect 1682 36165 1767 36401
rect 2003 36165 2088 36401
rect 2324 36165 2409 36401
rect 2645 36165 2730 36401
rect 2966 36165 3051 36401
rect 3287 36165 3372 36401
rect 3608 36165 3693 36401
rect 3929 36165 4014 36401
rect 4250 36165 4335 36401
rect 4571 36165 4656 36401
rect 4892 36165 4977 36401
rect 5213 36165 5298 36401
rect 5534 36165 5619 36401
rect 5855 36165 5940 36401
rect 6176 36165 6261 36401
rect 6497 36165 6582 36401
rect 6818 36165 6903 36401
rect 7139 36165 7224 36401
rect 7460 36165 7545 36401
rect 7781 36165 7866 36401
rect 8102 36165 8187 36401
rect 8423 36165 8508 36401
rect 8744 36165 8829 36401
rect 9065 36165 9150 36401
rect 9386 36165 9471 36401
rect 9707 36165 9792 36401
rect 10028 36165 10113 36401
rect 10349 36165 10434 36401
rect 10670 36165 10755 36401
rect 10991 36165 11076 36401
rect 11312 36165 11397 36401
rect 11633 36165 11718 36401
rect 11954 36165 12038 36401
rect 12274 36165 12358 36401
rect 12594 36165 12678 36401
rect 12914 36165 12998 36401
rect 13234 36165 13318 36401
rect 13554 36165 13638 36401
rect 13874 36165 13958 36401
rect 14194 36165 14278 36401
rect 14514 36165 14598 36401
rect 14834 36165 14918 36401
rect 15154 36165 15238 36401
rect 15474 36165 15558 36401
rect 15794 36165 16000 36401
rect 0 36077 16000 36165
rect 0 35841 162 36077
rect 398 35841 483 36077
rect 719 35841 804 36077
rect 1040 35841 1125 36077
rect 1361 35841 1446 36077
rect 1682 35841 1767 36077
rect 2003 35841 2088 36077
rect 2324 35841 2409 36077
rect 2645 35841 2730 36077
rect 2966 35841 3051 36077
rect 3287 35841 3372 36077
rect 3608 35841 3693 36077
rect 3929 35841 4014 36077
rect 4250 35841 4335 36077
rect 4571 35841 4656 36077
rect 4892 35841 4977 36077
rect 5213 35841 5298 36077
rect 5534 35841 5619 36077
rect 5855 35841 5940 36077
rect 6176 35841 6261 36077
rect 6497 35841 6582 36077
rect 6818 35841 6903 36077
rect 7139 35841 7224 36077
rect 7460 35841 7545 36077
rect 7781 35841 7866 36077
rect 8102 35841 8187 36077
rect 8423 35841 8508 36077
rect 8744 35841 8829 36077
rect 9065 35841 9150 36077
rect 9386 35841 9471 36077
rect 9707 35841 9792 36077
rect 10028 35841 10113 36077
rect 10349 35841 10434 36077
rect 10670 35841 10755 36077
rect 10991 35841 11076 36077
rect 11312 35841 11397 36077
rect 11633 35841 11718 36077
rect 11954 35841 12038 36077
rect 12274 35841 12358 36077
rect 12594 35841 12678 36077
rect 12914 35841 12998 36077
rect 13234 35841 13318 36077
rect 13554 35841 13638 36077
rect 13874 35841 13958 36077
rect 14194 35841 14278 36077
rect 14514 35841 14598 36077
rect 14834 35841 14918 36077
rect 15154 35841 15238 36077
rect 15474 35841 15558 36077
rect 15794 35841 16000 36077
rect 0 35753 16000 35841
rect 0 35517 162 35753
rect 398 35517 483 35753
rect 719 35517 804 35753
rect 1040 35517 1125 35753
rect 1361 35517 1446 35753
rect 1682 35517 1767 35753
rect 2003 35517 2088 35753
rect 2324 35517 2409 35753
rect 2645 35517 2730 35753
rect 2966 35517 3051 35753
rect 3287 35517 3372 35753
rect 3608 35517 3693 35753
rect 3929 35517 4014 35753
rect 4250 35517 4335 35753
rect 4571 35517 4656 35753
rect 4892 35517 4977 35753
rect 5213 35517 5298 35753
rect 5534 35517 5619 35753
rect 5855 35517 5940 35753
rect 6176 35517 6261 35753
rect 6497 35517 6582 35753
rect 6818 35517 6903 35753
rect 7139 35517 7224 35753
rect 7460 35517 7545 35753
rect 7781 35517 7866 35753
rect 8102 35517 8187 35753
rect 8423 35517 8508 35753
rect 8744 35517 8829 35753
rect 9065 35517 9150 35753
rect 9386 35517 9471 35753
rect 9707 35517 9792 35753
rect 10028 35517 10113 35753
rect 10349 35517 10434 35753
rect 10670 35517 10755 35753
rect 10991 35517 11076 35753
rect 11312 35517 11397 35753
rect 11633 35517 11718 35753
rect 11954 35517 12038 35753
rect 12274 35517 12358 35753
rect 12594 35517 12678 35753
rect 12914 35517 12998 35753
rect 13234 35517 13318 35753
rect 13554 35517 13638 35753
rect 13874 35517 13958 35753
rect 14194 35517 14278 35753
rect 14514 35517 14598 35753
rect 14834 35517 14918 35753
rect 15154 35517 15238 35753
rect 15474 35517 15558 35753
rect 15794 35517 16000 35753
rect 0 35429 16000 35517
rect 0 35193 162 35429
rect 398 35193 483 35429
rect 719 35193 804 35429
rect 1040 35193 1125 35429
rect 1361 35193 1446 35429
rect 1682 35193 1767 35429
rect 2003 35193 2088 35429
rect 2324 35193 2409 35429
rect 2645 35193 2730 35429
rect 2966 35193 3051 35429
rect 3287 35193 3372 35429
rect 3608 35193 3693 35429
rect 3929 35193 4014 35429
rect 4250 35193 4335 35429
rect 4571 35193 4656 35429
rect 4892 35193 4977 35429
rect 5213 35193 5298 35429
rect 5534 35193 5619 35429
rect 5855 35193 5940 35429
rect 6176 35193 6261 35429
rect 6497 35193 6582 35429
rect 6818 35193 6903 35429
rect 7139 35193 7224 35429
rect 7460 35193 7545 35429
rect 7781 35193 7866 35429
rect 8102 35193 8187 35429
rect 8423 35193 8508 35429
rect 8744 35193 8829 35429
rect 9065 35193 9150 35429
rect 9386 35193 9471 35429
rect 9707 35193 9792 35429
rect 10028 35193 10113 35429
rect 10349 35193 10434 35429
rect 10670 35193 10755 35429
rect 10991 35193 11076 35429
rect 11312 35193 11397 35429
rect 11633 35193 11718 35429
rect 11954 35193 12038 35429
rect 12274 35193 12358 35429
rect 12594 35193 12678 35429
rect 12914 35193 12998 35429
rect 13234 35193 13318 35429
rect 13554 35193 13638 35429
rect 13874 35193 13958 35429
rect 14194 35193 14278 35429
rect 14514 35193 14598 35429
rect 14834 35193 14918 35429
rect 15154 35193 15238 35429
rect 15474 35193 15558 35429
rect 15794 35193 16000 35429
rect 0 35182 16000 35193
rect 0 35157 254 35182
rect 15746 35157 16000 35182
rect 0 18973 254 19000
rect 15746 18973 16000 19000
rect 0 18972 16000 18973
rect 0 18736 162 18972
rect 398 18736 483 18972
rect 719 18736 804 18972
rect 1040 18736 1125 18972
rect 1361 18736 1446 18972
rect 1682 18736 1767 18972
rect 2003 18736 2088 18972
rect 2324 18736 2409 18972
rect 2645 18736 2730 18972
rect 2966 18736 3051 18972
rect 3287 18736 3372 18972
rect 3608 18736 3693 18972
rect 3929 18736 4014 18972
rect 4250 18736 4335 18972
rect 4571 18736 4656 18972
rect 4892 18736 4977 18972
rect 5213 18736 5298 18972
rect 5534 18736 5619 18972
rect 5855 18736 5940 18972
rect 6176 18736 6261 18972
rect 6497 18736 6582 18972
rect 6818 18736 6903 18972
rect 7139 18736 7224 18972
rect 7460 18736 7545 18972
rect 7781 18736 7866 18972
rect 8102 18736 8187 18972
rect 8423 18736 8508 18972
rect 8744 18736 8829 18972
rect 9065 18736 9150 18972
rect 9386 18736 9471 18972
rect 9707 18736 9792 18972
rect 10028 18736 10113 18972
rect 10349 18736 10434 18972
rect 10670 18736 10755 18972
rect 10991 18736 11076 18972
rect 11312 18736 11397 18972
rect 11633 18736 11718 18972
rect 11954 18736 12038 18972
rect 12274 18736 12358 18972
rect 12594 18736 12678 18972
rect 12914 18736 12998 18972
rect 13234 18736 13318 18972
rect 13554 18736 13638 18972
rect 13874 18736 13958 18972
rect 14194 18736 14278 18972
rect 14514 18736 14598 18972
rect 14834 18736 14918 18972
rect 15154 18736 15238 18972
rect 15474 18736 15558 18972
rect 15794 18736 16000 18972
rect 0 18636 16000 18736
rect 0 18400 162 18636
rect 398 18400 483 18636
rect 719 18400 804 18636
rect 1040 18400 1125 18636
rect 1361 18400 1446 18636
rect 1682 18400 1767 18636
rect 2003 18400 2088 18636
rect 2324 18400 2409 18636
rect 2645 18400 2730 18636
rect 2966 18400 3051 18636
rect 3287 18400 3372 18636
rect 3608 18400 3693 18636
rect 3929 18400 4014 18636
rect 4250 18400 4335 18636
rect 4571 18400 4656 18636
rect 4892 18400 4977 18636
rect 5213 18400 5298 18636
rect 5534 18400 5619 18636
rect 5855 18400 5940 18636
rect 6176 18400 6261 18636
rect 6497 18400 6582 18636
rect 6818 18400 6903 18636
rect 7139 18400 7224 18636
rect 7460 18400 7545 18636
rect 7781 18400 7866 18636
rect 8102 18400 8187 18636
rect 8423 18400 8508 18636
rect 8744 18400 8829 18636
rect 9065 18400 9150 18636
rect 9386 18400 9471 18636
rect 9707 18400 9792 18636
rect 10028 18400 10113 18636
rect 10349 18400 10434 18636
rect 10670 18400 10755 18636
rect 10991 18400 11076 18636
rect 11312 18400 11397 18636
rect 11633 18400 11718 18636
rect 11954 18400 12038 18636
rect 12274 18400 12358 18636
rect 12594 18400 12678 18636
rect 12914 18400 12998 18636
rect 13234 18400 13318 18636
rect 13554 18400 13638 18636
rect 13874 18400 13958 18636
rect 14194 18400 14278 18636
rect 14514 18400 14598 18636
rect 14834 18400 14918 18636
rect 15154 18400 15238 18636
rect 15474 18400 15558 18636
rect 15794 18400 16000 18636
rect 0 18300 16000 18400
rect 0 18064 162 18300
rect 398 18064 483 18300
rect 719 18064 804 18300
rect 1040 18064 1125 18300
rect 1361 18064 1446 18300
rect 1682 18064 1767 18300
rect 2003 18064 2088 18300
rect 2324 18064 2409 18300
rect 2645 18064 2730 18300
rect 2966 18064 3051 18300
rect 3287 18064 3372 18300
rect 3608 18064 3693 18300
rect 3929 18064 4014 18300
rect 4250 18064 4335 18300
rect 4571 18064 4656 18300
rect 4892 18064 4977 18300
rect 5213 18064 5298 18300
rect 5534 18064 5619 18300
rect 5855 18064 5940 18300
rect 6176 18064 6261 18300
rect 6497 18064 6582 18300
rect 6818 18064 6903 18300
rect 7139 18064 7224 18300
rect 7460 18064 7545 18300
rect 7781 18064 7866 18300
rect 8102 18064 8187 18300
rect 8423 18064 8508 18300
rect 8744 18064 8829 18300
rect 9065 18064 9150 18300
rect 9386 18064 9471 18300
rect 9707 18064 9792 18300
rect 10028 18064 10113 18300
rect 10349 18064 10434 18300
rect 10670 18064 10755 18300
rect 10991 18064 11076 18300
rect 11312 18064 11397 18300
rect 11633 18064 11718 18300
rect 11954 18064 12038 18300
rect 12274 18064 12358 18300
rect 12594 18064 12678 18300
rect 12914 18064 12998 18300
rect 13234 18064 13318 18300
rect 13554 18064 13638 18300
rect 13874 18064 13958 18300
rect 14194 18064 14278 18300
rect 14514 18064 14598 18300
rect 14834 18064 14918 18300
rect 15154 18064 15238 18300
rect 15474 18064 15558 18300
rect 15794 18064 16000 18300
rect 0 17964 16000 18064
rect 0 17728 162 17964
rect 398 17728 483 17964
rect 719 17728 804 17964
rect 1040 17728 1125 17964
rect 1361 17728 1446 17964
rect 1682 17728 1767 17964
rect 2003 17728 2088 17964
rect 2324 17728 2409 17964
rect 2645 17728 2730 17964
rect 2966 17728 3051 17964
rect 3287 17728 3372 17964
rect 3608 17728 3693 17964
rect 3929 17728 4014 17964
rect 4250 17728 4335 17964
rect 4571 17728 4656 17964
rect 4892 17728 4977 17964
rect 5213 17728 5298 17964
rect 5534 17728 5619 17964
rect 5855 17728 5940 17964
rect 6176 17728 6261 17964
rect 6497 17728 6582 17964
rect 6818 17728 6903 17964
rect 7139 17728 7224 17964
rect 7460 17728 7545 17964
rect 7781 17728 7866 17964
rect 8102 17728 8187 17964
rect 8423 17728 8508 17964
rect 8744 17728 8829 17964
rect 9065 17728 9150 17964
rect 9386 17728 9471 17964
rect 9707 17728 9792 17964
rect 10028 17728 10113 17964
rect 10349 17728 10434 17964
rect 10670 17728 10755 17964
rect 10991 17728 11076 17964
rect 11312 17728 11397 17964
rect 11633 17728 11718 17964
rect 11954 17728 12038 17964
rect 12274 17728 12358 17964
rect 12594 17728 12678 17964
rect 12914 17728 12998 17964
rect 13234 17728 13318 17964
rect 13554 17728 13638 17964
rect 13874 17728 13958 17964
rect 14194 17728 14278 17964
rect 14514 17728 14598 17964
rect 14834 17728 14918 17964
rect 15154 17728 15238 17964
rect 15474 17728 15558 17964
rect 15794 17728 16000 17964
rect 0 17628 16000 17728
rect 0 17392 162 17628
rect 398 17392 483 17628
rect 719 17392 804 17628
rect 1040 17392 1125 17628
rect 1361 17392 1446 17628
rect 1682 17392 1767 17628
rect 2003 17392 2088 17628
rect 2324 17392 2409 17628
rect 2645 17392 2730 17628
rect 2966 17392 3051 17628
rect 3287 17392 3372 17628
rect 3608 17392 3693 17628
rect 3929 17392 4014 17628
rect 4250 17392 4335 17628
rect 4571 17392 4656 17628
rect 4892 17392 4977 17628
rect 5213 17392 5298 17628
rect 5534 17392 5619 17628
rect 5855 17392 5940 17628
rect 6176 17392 6261 17628
rect 6497 17392 6582 17628
rect 6818 17392 6903 17628
rect 7139 17392 7224 17628
rect 7460 17392 7545 17628
rect 7781 17392 7866 17628
rect 8102 17392 8187 17628
rect 8423 17392 8508 17628
rect 8744 17392 8829 17628
rect 9065 17392 9150 17628
rect 9386 17392 9471 17628
rect 9707 17392 9792 17628
rect 10028 17392 10113 17628
rect 10349 17392 10434 17628
rect 10670 17392 10755 17628
rect 10991 17392 11076 17628
rect 11312 17392 11397 17628
rect 11633 17392 11718 17628
rect 11954 17392 12038 17628
rect 12274 17392 12358 17628
rect 12594 17392 12678 17628
rect 12914 17392 12998 17628
rect 13234 17392 13318 17628
rect 13554 17392 13638 17628
rect 13874 17392 13958 17628
rect 14194 17392 14278 17628
rect 14514 17392 14598 17628
rect 14834 17392 14918 17628
rect 15154 17392 15238 17628
rect 15474 17392 15558 17628
rect 15794 17392 16000 17628
rect 0 17292 16000 17392
rect 0 17056 162 17292
rect 398 17056 483 17292
rect 719 17056 804 17292
rect 1040 17056 1125 17292
rect 1361 17056 1446 17292
rect 1682 17056 1767 17292
rect 2003 17056 2088 17292
rect 2324 17056 2409 17292
rect 2645 17056 2730 17292
rect 2966 17056 3051 17292
rect 3287 17056 3372 17292
rect 3608 17056 3693 17292
rect 3929 17056 4014 17292
rect 4250 17056 4335 17292
rect 4571 17056 4656 17292
rect 4892 17056 4977 17292
rect 5213 17056 5298 17292
rect 5534 17056 5619 17292
rect 5855 17056 5940 17292
rect 6176 17056 6261 17292
rect 6497 17056 6582 17292
rect 6818 17056 6903 17292
rect 7139 17056 7224 17292
rect 7460 17056 7545 17292
rect 7781 17056 7866 17292
rect 8102 17056 8187 17292
rect 8423 17056 8508 17292
rect 8744 17056 8829 17292
rect 9065 17056 9150 17292
rect 9386 17056 9471 17292
rect 9707 17056 9792 17292
rect 10028 17056 10113 17292
rect 10349 17056 10434 17292
rect 10670 17056 10755 17292
rect 10991 17056 11076 17292
rect 11312 17056 11397 17292
rect 11633 17056 11718 17292
rect 11954 17056 12038 17292
rect 12274 17056 12358 17292
rect 12594 17056 12678 17292
rect 12914 17056 12998 17292
rect 13234 17056 13318 17292
rect 13554 17056 13638 17292
rect 13874 17056 13958 17292
rect 14194 17056 14278 17292
rect 14514 17056 14598 17292
rect 14834 17056 14918 17292
rect 15154 17056 15238 17292
rect 15474 17056 15558 17292
rect 15794 17056 16000 17292
rect 0 16956 16000 17056
rect 0 16720 162 16956
rect 398 16720 483 16956
rect 719 16720 804 16956
rect 1040 16720 1125 16956
rect 1361 16720 1446 16956
rect 1682 16720 1767 16956
rect 2003 16720 2088 16956
rect 2324 16720 2409 16956
rect 2645 16720 2730 16956
rect 2966 16720 3051 16956
rect 3287 16720 3372 16956
rect 3608 16720 3693 16956
rect 3929 16720 4014 16956
rect 4250 16720 4335 16956
rect 4571 16720 4656 16956
rect 4892 16720 4977 16956
rect 5213 16720 5298 16956
rect 5534 16720 5619 16956
rect 5855 16720 5940 16956
rect 6176 16720 6261 16956
rect 6497 16720 6582 16956
rect 6818 16720 6903 16956
rect 7139 16720 7224 16956
rect 7460 16720 7545 16956
rect 7781 16720 7866 16956
rect 8102 16720 8187 16956
rect 8423 16720 8508 16956
rect 8744 16720 8829 16956
rect 9065 16720 9150 16956
rect 9386 16720 9471 16956
rect 9707 16720 9792 16956
rect 10028 16720 10113 16956
rect 10349 16720 10434 16956
rect 10670 16720 10755 16956
rect 10991 16720 11076 16956
rect 11312 16720 11397 16956
rect 11633 16720 11718 16956
rect 11954 16720 12038 16956
rect 12274 16720 12358 16956
rect 12594 16720 12678 16956
rect 12914 16720 12998 16956
rect 13234 16720 13318 16956
rect 13554 16720 13638 16956
rect 13874 16720 13958 16956
rect 14194 16720 14278 16956
rect 14514 16720 14598 16956
rect 14834 16720 14918 16956
rect 15154 16720 15238 16956
rect 15474 16720 15558 16956
rect 15794 16720 16000 16956
rect 0 16620 16000 16720
rect 0 16384 162 16620
rect 398 16384 483 16620
rect 719 16384 804 16620
rect 1040 16384 1125 16620
rect 1361 16384 1446 16620
rect 1682 16384 1767 16620
rect 2003 16384 2088 16620
rect 2324 16384 2409 16620
rect 2645 16384 2730 16620
rect 2966 16384 3051 16620
rect 3287 16384 3372 16620
rect 3608 16384 3693 16620
rect 3929 16384 4014 16620
rect 4250 16384 4335 16620
rect 4571 16384 4656 16620
rect 4892 16384 4977 16620
rect 5213 16384 5298 16620
rect 5534 16384 5619 16620
rect 5855 16384 5940 16620
rect 6176 16384 6261 16620
rect 6497 16384 6582 16620
rect 6818 16384 6903 16620
rect 7139 16384 7224 16620
rect 7460 16384 7545 16620
rect 7781 16384 7866 16620
rect 8102 16384 8187 16620
rect 8423 16384 8508 16620
rect 8744 16384 8829 16620
rect 9065 16384 9150 16620
rect 9386 16384 9471 16620
rect 9707 16384 9792 16620
rect 10028 16384 10113 16620
rect 10349 16384 10434 16620
rect 10670 16384 10755 16620
rect 10991 16384 11076 16620
rect 11312 16384 11397 16620
rect 11633 16384 11718 16620
rect 11954 16384 12038 16620
rect 12274 16384 12358 16620
rect 12594 16384 12678 16620
rect 12914 16384 12998 16620
rect 13234 16384 13318 16620
rect 13554 16384 13638 16620
rect 13874 16384 13958 16620
rect 14194 16384 14278 16620
rect 14514 16384 14598 16620
rect 14834 16384 14918 16620
rect 15154 16384 15238 16620
rect 15474 16384 15558 16620
rect 15794 16384 16000 16620
rect 0 16284 16000 16384
rect 0 16048 162 16284
rect 398 16048 483 16284
rect 719 16048 804 16284
rect 1040 16048 1125 16284
rect 1361 16048 1446 16284
rect 1682 16048 1767 16284
rect 2003 16048 2088 16284
rect 2324 16048 2409 16284
rect 2645 16048 2730 16284
rect 2966 16048 3051 16284
rect 3287 16048 3372 16284
rect 3608 16048 3693 16284
rect 3929 16048 4014 16284
rect 4250 16048 4335 16284
rect 4571 16048 4656 16284
rect 4892 16048 4977 16284
rect 5213 16048 5298 16284
rect 5534 16048 5619 16284
rect 5855 16048 5940 16284
rect 6176 16048 6261 16284
rect 6497 16048 6582 16284
rect 6818 16048 6903 16284
rect 7139 16048 7224 16284
rect 7460 16048 7545 16284
rect 7781 16048 7866 16284
rect 8102 16048 8187 16284
rect 8423 16048 8508 16284
rect 8744 16048 8829 16284
rect 9065 16048 9150 16284
rect 9386 16048 9471 16284
rect 9707 16048 9792 16284
rect 10028 16048 10113 16284
rect 10349 16048 10434 16284
rect 10670 16048 10755 16284
rect 10991 16048 11076 16284
rect 11312 16048 11397 16284
rect 11633 16048 11718 16284
rect 11954 16048 12038 16284
rect 12274 16048 12358 16284
rect 12594 16048 12678 16284
rect 12914 16048 12998 16284
rect 13234 16048 13318 16284
rect 13554 16048 13638 16284
rect 13874 16048 13958 16284
rect 14194 16048 14278 16284
rect 14514 16048 14598 16284
rect 14834 16048 14918 16284
rect 15154 16048 15238 16284
rect 15474 16048 15558 16284
rect 15794 16048 16000 16284
rect 0 15948 16000 16048
rect 0 15712 162 15948
rect 398 15712 483 15948
rect 719 15712 804 15948
rect 1040 15712 1125 15948
rect 1361 15712 1446 15948
rect 1682 15712 1767 15948
rect 2003 15712 2088 15948
rect 2324 15712 2409 15948
rect 2645 15712 2730 15948
rect 2966 15712 3051 15948
rect 3287 15712 3372 15948
rect 3608 15712 3693 15948
rect 3929 15712 4014 15948
rect 4250 15712 4335 15948
rect 4571 15712 4656 15948
rect 4892 15712 4977 15948
rect 5213 15712 5298 15948
rect 5534 15712 5619 15948
rect 5855 15712 5940 15948
rect 6176 15712 6261 15948
rect 6497 15712 6582 15948
rect 6818 15712 6903 15948
rect 7139 15712 7224 15948
rect 7460 15712 7545 15948
rect 7781 15712 7866 15948
rect 8102 15712 8187 15948
rect 8423 15712 8508 15948
rect 8744 15712 8829 15948
rect 9065 15712 9150 15948
rect 9386 15712 9471 15948
rect 9707 15712 9792 15948
rect 10028 15712 10113 15948
rect 10349 15712 10434 15948
rect 10670 15712 10755 15948
rect 10991 15712 11076 15948
rect 11312 15712 11397 15948
rect 11633 15712 11718 15948
rect 11954 15712 12038 15948
rect 12274 15712 12358 15948
rect 12594 15712 12678 15948
rect 12914 15712 12998 15948
rect 13234 15712 13318 15948
rect 13554 15712 13638 15948
rect 13874 15712 13958 15948
rect 14194 15712 14278 15948
rect 14514 15712 14598 15948
rect 14834 15712 14918 15948
rect 15154 15712 15238 15948
rect 15474 15712 15558 15948
rect 15794 15712 16000 15948
rect 0 15612 16000 15712
rect 0 15376 162 15612
rect 398 15376 483 15612
rect 719 15376 804 15612
rect 1040 15376 1125 15612
rect 1361 15376 1446 15612
rect 1682 15376 1767 15612
rect 2003 15376 2088 15612
rect 2324 15376 2409 15612
rect 2645 15376 2730 15612
rect 2966 15376 3051 15612
rect 3287 15376 3372 15612
rect 3608 15376 3693 15612
rect 3929 15376 4014 15612
rect 4250 15376 4335 15612
rect 4571 15376 4656 15612
rect 4892 15376 4977 15612
rect 5213 15376 5298 15612
rect 5534 15376 5619 15612
rect 5855 15376 5940 15612
rect 6176 15376 6261 15612
rect 6497 15376 6582 15612
rect 6818 15376 6903 15612
rect 7139 15376 7224 15612
rect 7460 15376 7545 15612
rect 7781 15376 7866 15612
rect 8102 15376 8187 15612
rect 8423 15376 8508 15612
rect 8744 15376 8829 15612
rect 9065 15376 9150 15612
rect 9386 15376 9471 15612
rect 9707 15376 9792 15612
rect 10028 15376 10113 15612
rect 10349 15376 10434 15612
rect 10670 15376 10755 15612
rect 10991 15376 11076 15612
rect 11312 15376 11397 15612
rect 11633 15376 11718 15612
rect 11954 15376 12038 15612
rect 12274 15376 12358 15612
rect 12594 15376 12678 15612
rect 12914 15376 12998 15612
rect 13234 15376 13318 15612
rect 13554 15376 13638 15612
rect 13874 15376 13958 15612
rect 14194 15376 14278 15612
rect 14514 15376 14598 15612
rect 14834 15376 14918 15612
rect 15154 15376 15238 15612
rect 15474 15376 15558 15612
rect 15794 15376 16000 15612
rect 0 15276 16000 15376
rect 0 15040 162 15276
rect 398 15040 483 15276
rect 719 15040 804 15276
rect 1040 15040 1125 15276
rect 1361 15040 1446 15276
rect 1682 15040 1767 15276
rect 2003 15040 2088 15276
rect 2324 15040 2409 15276
rect 2645 15040 2730 15276
rect 2966 15040 3051 15276
rect 3287 15040 3372 15276
rect 3608 15040 3693 15276
rect 3929 15040 4014 15276
rect 4250 15040 4335 15276
rect 4571 15040 4656 15276
rect 4892 15040 4977 15276
rect 5213 15040 5298 15276
rect 5534 15040 5619 15276
rect 5855 15040 5940 15276
rect 6176 15040 6261 15276
rect 6497 15040 6582 15276
rect 6818 15040 6903 15276
rect 7139 15040 7224 15276
rect 7460 15040 7545 15276
rect 7781 15040 7866 15276
rect 8102 15040 8187 15276
rect 8423 15040 8508 15276
rect 8744 15040 8829 15276
rect 9065 15040 9150 15276
rect 9386 15040 9471 15276
rect 9707 15040 9792 15276
rect 10028 15040 10113 15276
rect 10349 15040 10434 15276
rect 10670 15040 10755 15276
rect 10991 15040 11076 15276
rect 11312 15040 11397 15276
rect 11633 15040 11718 15276
rect 11954 15040 12038 15276
rect 12274 15040 12358 15276
rect 12594 15040 12678 15276
rect 12914 15040 12998 15276
rect 13234 15040 13318 15276
rect 13554 15040 13638 15276
rect 13874 15040 13958 15276
rect 14194 15040 14278 15276
rect 14514 15040 14598 15276
rect 14834 15040 14918 15276
rect 15154 15040 15238 15276
rect 15474 15040 15558 15276
rect 15794 15040 16000 15276
rect 0 14940 16000 15040
rect 0 14704 162 14940
rect 398 14704 483 14940
rect 719 14704 804 14940
rect 1040 14704 1125 14940
rect 1361 14704 1446 14940
rect 1682 14704 1767 14940
rect 2003 14704 2088 14940
rect 2324 14704 2409 14940
rect 2645 14704 2730 14940
rect 2966 14704 3051 14940
rect 3287 14704 3372 14940
rect 3608 14704 3693 14940
rect 3929 14704 4014 14940
rect 4250 14704 4335 14940
rect 4571 14704 4656 14940
rect 4892 14704 4977 14940
rect 5213 14704 5298 14940
rect 5534 14704 5619 14940
rect 5855 14704 5940 14940
rect 6176 14704 6261 14940
rect 6497 14704 6582 14940
rect 6818 14704 6903 14940
rect 7139 14704 7224 14940
rect 7460 14704 7545 14940
rect 7781 14704 7866 14940
rect 8102 14704 8187 14940
rect 8423 14704 8508 14940
rect 8744 14704 8829 14940
rect 9065 14704 9150 14940
rect 9386 14704 9471 14940
rect 9707 14704 9792 14940
rect 10028 14704 10113 14940
rect 10349 14704 10434 14940
rect 10670 14704 10755 14940
rect 10991 14704 11076 14940
rect 11312 14704 11397 14940
rect 11633 14704 11718 14940
rect 11954 14704 12038 14940
rect 12274 14704 12358 14940
rect 12594 14704 12678 14940
rect 12914 14704 12998 14940
rect 13234 14704 13318 14940
rect 13554 14704 13638 14940
rect 13874 14704 13958 14940
rect 14194 14704 14278 14940
rect 14514 14704 14598 14940
rect 14834 14704 14918 14940
rect 15154 14704 15238 14940
rect 15474 14704 15558 14940
rect 15794 14704 16000 14940
rect 0 14604 16000 14704
rect 0 14368 162 14604
rect 398 14368 483 14604
rect 719 14368 804 14604
rect 1040 14368 1125 14604
rect 1361 14368 1446 14604
rect 1682 14368 1767 14604
rect 2003 14368 2088 14604
rect 2324 14368 2409 14604
rect 2645 14368 2730 14604
rect 2966 14368 3051 14604
rect 3287 14368 3372 14604
rect 3608 14368 3693 14604
rect 3929 14368 4014 14604
rect 4250 14368 4335 14604
rect 4571 14368 4656 14604
rect 4892 14368 4977 14604
rect 5213 14368 5298 14604
rect 5534 14368 5619 14604
rect 5855 14368 5940 14604
rect 6176 14368 6261 14604
rect 6497 14368 6582 14604
rect 6818 14368 6903 14604
rect 7139 14368 7224 14604
rect 7460 14368 7545 14604
rect 7781 14368 7866 14604
rect 8102 14368 8187 14604
rect 8423 14368 8508 14604
rect 8744 14368 8829 14604
rect 9065 14368 9150 14604
rect 9386 14368 9471 14604
rect 9707 14368 9792 14604
rect 10028 14368 10113 14604
rect 10349 14368 10434 14604
rect 10670 14368 10755 14604
rect 10991 14368 11076 14604
rect 11312 14368 11397 14604
rect 11633 14368 11718 14604
rect 11954 14368 12038 14604
rect 12274 14368 12358 14604
rect 12594 14368 12678 14604
rect 12914 14368 12998 14604
rect 13234 14368 13318 14604
rect 13554 14368 13638 14604
rect 13874 14368 13958 14604
rect 14194 14368 14278 14604
rect 14514 14368 14598 14604
rect 14834 14368 14918 14604
rect 15154 14368 15238 14604
rect 15474 14368 15558 14604
rect 15794 14368 16000 14604
rect 0 14268 16000 14368
rect 0 14032 162 14268
rect 398 14032 483 14268
rect 719 14032 804 14268
rect 1040 14032 1125 14268
rect 1361 14032 1446 14268
rect 1682 14032 1767 14268
rect 2003 14032 2088 14268
rect 2324 14032 2409 14268
rect 2645 14032 2730 14268
rect 2966 14032 3051 14268
rect 3287 14032 3372 14268
rect 3608 14032 3693 14268
rect 3929 14032 4014 14268
rect 4250 14032 4335 14268
rect 4571 14032 4656 14268
rect 4892 14032 4977 14268
rect 5213 14032 5298 14268
rect 5534 14032 5619 14268
rect 5855 14032 5940 14268
rect 6176 14032 6261 14268
rect 6497 14032 6582 14268
rect 6818 14032 6903 14268
rect 7139 14032 7224 14268
rect 7460 14032 7545 14268
rect 7781 14032 7866 14268
rect 8102 14032 8187 14268
rect 8423 14032 8508 14268
rect 8744 14032 8829 14268
rect 9065 14032 9150 14268
rect 9386 14032 9471 14268
rect 9707 14032 9792 14268
rect 10028 14032 10113 14268
rect 10349 14032 10434 14268
rect 10670 14032 10755 14268
rect 10991 14032 11076 14268
rect 11312 14032 11397 14268
rect 11633 14032 11718 14268
rect 11954 14032 12038 14268
rect 12274 14032 12358 14268
rect 12594 14032 12678 14268
rect 12914 14032 12998 14268
rect 13234 14032 13318 14268
rect 13554 14032 13638 14268
rect 13874 14032 13958 14268
rect 14194 14032 14278 14268
rect 14514 14032 14598 14268
rect 14834 14032 14918 14268
rect 15154 14032 15238 14268
rect 15474 14032 15558 14268
rect 15794 14032 16000 14268
rect 0 14031 16000 14032
rect 0 14007 254 14031
rect 15746 14007 16000 14031
rect 0 13663 254 13707
rect 15746 13663 16000 13707
rect 0 13427 162 13663
rect 398 13427 483 13663
rect 719 13427 804 13663
rect 1040 13427 1125 13663
rect 1361 13427 1446 13663
rect 1682 13427 1767 13663
rect 2003 13427 2088 13663
rect 2324 13427 2409 13663
rect 2645 13427 2730 13663
rect 2966 13427 3051 13663
rect 3287 13427 3372 13663
rect 3608 13427 3693 13663
rect 3929 13427 4014 13663
rect 4250 13427 4335 13663
rect 4571 13427 4656 13663
rect 4892 13427 4977 13663
rect 5213 13427 5298 13663
rect 5534 13427 5619 13663
rect 5855 13427 5940 13663
rect 6176 13427 6261 13663
rect 6497 13427 6582 13663
rect 6818 13427 6903 13663
rect 7139 13427 7224 13663
rect 7460 13427 7545 13663
rect 7781 13427 7866 13663
rect 8102 13427 8187 13663
rect 8423 13427 8508 13663
rect 8744 13427 8829 13663
rect 9065 13427 9150 13663
rect 9386 13427 9471 13663
rect 9707 13427 9792 13663
rect 10028 13427 10113 13663
rect 10349 13427 10434 13663
rect 10670 13427 10755 13663
rect 10991 13427 11076 13663
rect 11312 13427 11397 13663
rect 11633 13427 11718 13663
rect 11954 13427 12038 13663
rect 12274 13427 12358 13663
rect 12594 13427 12678 13663
rect 12914 13427 12998 13663
rect 13234 13427 13318 13663
rect 13554 13427 13638 13663
rect 13874 13427 13958 13663
rect 14194 13427 14278 13663
rect 14514 13427 14598 13663
rect 14834 13427 14918 13663
rect 15154 13427 15238 13663
rect 15474 13427 15558 13663
rect 15794 13427 16000 13663
rect 0 13097 16000 13427
rect 0 12861 162 13097
rect 398 12861 483 13097
rect 719 12861 804 13097
rect 1040 12861 1125 13097
rect 1361 12861 1446 13097
rect 1682 12861 1767 13097
rect 2003 12861 2088 13097
rect 2324 12861 2409 13097
rect 2645 12861 2730 13097
rect 2966 12861 3051 13097
rect 3287 12861 3372 13097
rect 3608 12861 3693 13097
rect 3929 12861 4014 13097
rect 4250 12861 4335 13097
rect 4571 12861 4656 13097
rect 4892 12861 4977 13097
rect 5213 12861 5298 13097
rect 5534 12861 5619 13097
rect 5855 12861 5940 13097
rect 6176 12861 6261 13097
rect 6497 12861 6582 13097
rect 6818 12861 6903 13097
rect 7139 12861 7224 13097
rect 7460 12861 7545 13097
rect 7781 12861 7866 13097
rect 8102 12861 8187 13097
rect 8423 12861 8508 13097
rect 8744 12861 8829 13097
rect 9065 12861 9150 13097
rect 9386 12861 9471 13097
rect 9707 12861 9792 13097
rect 10028 12861 10113 13097
rect 10349 12861 10434 13097
rect 10670 12861 10755 13097
rect 10991 12861 11076 13097
rect 11312 12861 11397 13097
rect 11633 12861 11718 13097
rect 11954 12861 12038 13097
rect 12274 12861 12358 13097
rect 12594 12861 12678 13097
rect 12914 12861 12998 13097
rect 13234 12861 13318 13097
rect 13554 12861 13638 13097
rect 13874 12861 13958 13097
rect 14194 12861 14278 13097
rect 14514 12861 14598 13097
rect 14834 12861 14918 13097
rect 15154 12861 15238 13097
rect 15474 12861 15558 13097
rect 15794 12861 16000 13097
rect 0 12817 254 12861
rect 15746 12817 16000 12861
rect 0 12493 254 12537
rect 15746 12493 16000 12537
rect 0 12257 162 12493
rect 398 12257 483 12493
rect 719 12257 804 12493
rect 1040 12257 1125 12493
rect 1361 12257 1446 12493
rect 1682 12257 1767 12493
rect 2003 12257 2088 12493
rect 2324 12257 2409 12493
rect 2645 12257 2730 12493
rect 2966 12257 3051 12493
rect 3287 12257 3372 12493
rect 3608 12257 3693 12493
rect 3929 12257 4014 12493
rect 4250 12257 4335 12493
rect 4571 12257 4656 12493
rect 4892 12257 4977 12493
rect 5213 12257 5298 12493
rect 5534 12257 5619 12493
rect 5855 12257 5940 12493
rect 6176 12257 6261 12493
rect 6497 12257 6582 12493
rect 6818 12257 6903 12493
rect 7139 12257 7224 12493
rect 7460 12257 7545 12493
rect 7781 12257 7866 12493
rect 8102 12257 8187 12493
rect 8423 12257 8508 12493
rect 8744 12257 8829 12493
rect 9065 12257 9150 12493
rect 9386 12257 9471 12493
rect 9707 12257 9792 12493
rect 10028 12257 10113 12493
rect 10349 12257 10434 12493
rect 10670 12257 10755 12493
rect 10991 12257 11076 12493
rect 11312 12257 11397 12493
rect 11633 12257 11718 12493
rect 11954 12257 12039 12493
rect 12275 12257 12359 12493
rect 12595 12257 12679 12493
rect 12915 12257 12999 12493
rect 13235 12257 13319 12493
rect 13555 12257 13639 12493
rect 13875 12257 13959 12493
rect 14195 12257 14279 12493
rect 14515 12257 14599 12493
rect 14835 12257 14919 12493
rect 15155 12257 15239 12493
rect 15475 12257 15559 12493
rect 15795 12257 16000 12493
rect 0 11927 16000 12257
rect 0 11691 162 11927
rect 398 11691 483 11927
rect 719 11691 804 11927
rect 1040 11691 1125 11927
rect 1361 11691 1446 11927
rect 1682 11691 1767 11927
rect 2003 11691 2088 11927
rect 2324 11691 2409 11927
rect 2645 11691 2730 11927
rect 2966 11691 3051 11927
rect 3287 11691 3372 11927
rect 3608 11691 3693 11927
rect 3929 11691 4014 11927
rect 4250 11691 4335 11927
rect 4571 11691 4656 11927
rect 4892 11691 4977 11927
rect 5213 11691 5298 11927
rect 5534 11691 5619 11927
rect 5855 11691 5940 11927
rect 6176 11691 6261 11927
rect 6497 11691 6582 11927
rect 6818 11691 6903 11927
rect 7139 11691 7224 11927
rect 7460 11691 7545 11927
rect 7781 11691 7866 11927
rect 8102 11691 8187 11927
rect 8423 11691 8508 11927
rect 8744 11691 8829 11927
rect 9065 11691 9150 11927
rect 9386 11691 9471 11927
rect 9707 11691 9792 11927
rect 10028 11691 10113 11927
rect 10349 11691 10434 11927
rect 10670 11691 10755 11927
rect 10991 11691 11076 11927
rect 11312 11691 11397 11927
rect 11633 11691 11718 11927
rect 11954 11691 12039 11927
rect 12275 11691 12359 11927
rect 12595 11691 12679 11927
rect 12915 11691 12999 11927
rect 13235 11691 13319 11927
rect 13555 11691 13639 11927
rect 13875 11691 13959 11927
rect 14195 11691 14279 11927
rect 14515 11691 14599 11927
rect 14835 11691 14919 11927
rect 15155 11691 15239 11927
rect 15475 11691 15559 11927
rect 15795 11691 16000 11927
rect 0 11647 254 11691
rect 15746 11647 16000 11691
rect 0 11281 254 11347
rect 15746 11281 16000 11347
rect 0 10625 254 11221
rect 15746 10625 16000 11221
rect 0 10329 162 10565
rect 398 10329 483 10565
rect 719 10329 804 10565
rect 1040 10329 1125 10565
rect 1361 10329 1446 10565
rect 1682 10329 1767 10565
rect 2003 10329 2088 10565
rect 2324 10329 2409 10565
rect 2645 10329 2730 10565
rect 2966 10329 3051 10565
rect 3287 10329 3372 10565
rect 3608 10329 3693 10565
rect 3929 10329 4014 10565
rect 4250 10329 4335 10565
rect 4571 10329 4656 10565
rect 4892 10329 4977 10565
rect 5213 10329 5298 10565
rect 5534 10329 5619 10565
rect 5855 10329 5940 10565
rect 6176 10329 6261 10565
rect 6497 10329 6582 10565
rect 6818 10329 6903 10565
rect 7139 10329 7224 10565
rect 7460 10329 7545 10565
rect 7781 10329 7866 10565
rect 8102 10329 8187 10565
rect 8423 10329 8508 10565
rect 8744 10329 8829 10565
rect 9065 10329 9150 10565
rect 9386 10329 9471 10565
rect 9707 10329 9792 10565
rect 10028 10329 10113 10565
rect 10349 10329 10434 10565
rect 10670 10329 10755 10565
rect 10991 10329 11076 10565
rect 11312 10329 11397 10565
rect 11633 10329 11718 10565
rect 11954 10329 12038 10565
rect 12274 10329 12358 10565
rect 12594 10329 12678 10565
rect 12914 10329 12998 10565
rect 13234 10329 13318 10565
rect 13554 10329 13638 10565
rect 13874 10329 13958 10565
rect 14194 10329 14278 10565
rect 14514 10329 14598 10565
rect 14834 10329 14918 10565
rect 15154 10329 15238 10565
rect 15474 10329 15558 10565
rect 15794 10329 16000 10565
rect 0 9673 254 10269
rect 15746 9673 16000 10269
rect 0 9547 254 9613
rect 15746 9547 16000 9613
rect 0 9203 254 9247
rect 15746 9203 16000 9247
rect 0 8967 162 9203
rect 398 8967 483 9203
rect 719 8967 804 9203
rect 1040 8967 1125 9203
rect 1361 8967 1446 9203
rect 1682 8967 1767 9203
rect 2003 8967 2088 9203
rect 2324 8967 2409 9203
rect 2645 8967 2730 9203
rect 2966 8967 3051 9203
rect 3287 8967 3372 9203
rect 3608 8967 3693 9203
rect 3929 8967 4014 9203
rect 4250 8967 4335 9203
rect 4571 8967 4656 9203
rect 4892 8967 4977 9203
rect 5213 8967 5298 9203
rect 5534 8967 5619 9203
rect 5855 8967 5940 9203
rect 6176 8967 6261 9203
rect 6497 8967 6582 9203
rect 6818 8967 6903 9203
rect 7139 8967 7224 9203
rect 7460 8967 7545 9203
rect 7781 8967 7866 9203
rect 8102 8967 8187 9203
rect 8423 8967 8508 9203
rect 8744 8967 8829 9203
rect 9065 8967 9150 9203
rect 9386 8967 9471 9203
rect 9707 8967 9792 9203
rect 10028 8967 10113 9203
rect 10349 8967 10434 9203
rect 10670 8967 10755 9203
rect 10991 8967 11076 9203
rect 11312 8967 11397 9203
rect 11633 8967 11717 9203
rect 11953 8967 12037 9203
rect 12273 8967 12357 9203
rect 12593 8967 12677 9203
rect 12913 8967 12997 9203
rect 13233 8967 13317 9203
rect 13553 8967 13637 9203
rect 13873 8967 13957 9203
rect 14193 8967 14277 9203
rect 14513 8967 14597 9203
rect 14833 8967 14917 9203
rect 15153 8967 15237 9203
rect 15473 8967 15557 9203
rect 15793 8967 16000 9203
rect 0 8597 16000 8967
rect 0 8361 162 8597
rect 398 8361 483 8597
rect 719 8361 804 8597
rect 1040 8361 1125 8597
rect 1361 8361 1446 8597
rect 1682 8361 1767 8597
rect 2003 8361 2088 8597
rect 2324 8361 2409 8597
rect 2645 8361 2730 8597
rect 2966 8361 3051 8597
rect 3287 8361 3372 8597
rect 3608 8361 3693 8597
rect 3929 8361 4014 8597
rect 4250 8361 4335 8597
rect 4571 8361 4656 8597
rect 4892 8361 4977 8597
rect 5213 8361 5298 8597
rect 5534 8361 5619 8597
rect 5855 8361 5940 8597
rect 6176 8361 6261 8597
rect 6497 8361 6582 8597
rect 6818 8361 6903 8597
rect 7139 8361 7224 8597
rect 7460 8361 7545 8597
rect 7781 8361 7866 8597
rect 8102 8361 8187 8597
rect 8423 8361 8508 8597
rect 8744 8361 8829 8597
rect 9065 8361 9150 8597
rect 9386 8361 9471 8597
rect 9707 8361 9792 8597
rect 10028 8361 10113 8597
rect 10349 8361 10434 8597
rect 10670 8361 10755 8597
rect 10991 8361 11076 8597
rect 11312 8361 11397 8597
rect 11633 8361 11717 8597
rect 11953 8361 12037 8597
rect 12273 8361 12357 8597
rect 12593 8361 12677 8597
rect 12913 8361 12997 8597
rect 13233 8361 13317 8597
rect 13553 8361 13637 8597
rect 13873 8361 13957 8597
rect 14193 8361 14277 8597
rect 14513 8361 14597 8597
rect 14833 8361 14917 8597
rect 15153 8361 15237 8597
rect 15473 8361 15557 8597
rect 15793 8361 16000 8597
rect 0 8317 254 8361
rect 15746 8317 16000 8361
rect 0 7993 254 8037
rect 15746 7993 16000 8037
rect 0 7757 162 7993
rect 398 7757 483 7993
rect 719 7757 804 7993
rect 1040 7757 1125 7993
rect 1361 7757 1446 7993
rect 1682 7757 1767 7993
rect 2003 7757 2088 7993
rect 2324 7757 2409 7993
rect 2645 7757 2730 7993
rect 2966 7757 3051 7993
rect 3287 7757 3372 7993
rect 3608 7757 3693 7993
rect 3929 7757 4014 7993
rect 4250 7757 4335 7993
rect 4571 7757 4656 7993
rect 4892 7757 4977 7993
rect 5213 7757 5298 7993
rect 5534 7757 5619 7993
rect 5855 7757 5940 7993
rect 6176 7757 6261 7993
rect 6497 7757 6582 7993
rect 6818 7757 6903 7993
rect 7139 7757 7224 7993
rect 7460 7757 7545 7993
rect 7781 7757 7866 7993
rect 8102 7757 8187 7993
rect 8423 7757 8508 7993
rect 8744 7757 8829 7993
rect 9065 7757 9150 7993
rect 9386 7757 9471 7993
rect 9707 7757 9792 7993
rect 10028 7757 10113 7993
rect 10349 7757 10434 7993
rect 10670 7757 10755 7993
rect 10991 7757 11076 7993
rect 11312 7757 11397 7993
rect 11633 7757 11718 7993
rect 11954 7757 12039 7993
rect 12275 7757 12359 7993
rect 12595 7757 12679 7993
rect 12915 7757 12999 7993
rect 13235 7757 13319 7993
rect 13555 7757 13639 7993
rect 13875 7757 13959 7993
rect 14195 7757 14279 7993
rect 14515 7757 14599 7993
rect 14835 7757 14919 7993
rect 15155 7757 15239 7993
rect 15475 7757 15559 7993
rect 15795 7757 16000 7993
rect 0 7627 16000 7757
rect 0 7391 162 7627
rect 398 7391 483 7627
rect 719 7391 804 7627
rect 1040 7391 1125 7627
rect 1361 7391 1446 7627
rect 1682 7391 1767 7627
rect 2003 7391 2088 7627
rect 2324 7391 2409 7627
rect 2645 7391 2730 7627
rect 2966 7391 3051 7627
rect 3287 7391 3372 7627
rect 3608 7391 3693 7627
rect 3929 7391 4014 7627
rect 4250 7391 4335 7627
rect 4571 7391 4656 7627
rect 4892 7391 4977 7627
rect 5213 7391 5298 7627
rect 5534 7391 5619 7627
rect 5855 7391 5940 7627
rect 6176 7391 6261 7627
rect 6497 7391 6582 7627
rect 6818 7391 6903 7627
rect 7139 7391 7224 7627
rect 7460 7391 7545 7627
rect 7781 7391 7866 7627
rect 8102 7391 8187 7627
rect 8423 7391 8508 7627
rect 8744 7391 8829 7627
rect 9065 7391 9150 7627
rect 9386 7391 9471 7627
rect 9707 7391 9792 7627
rect 10028 7391 10113 7627
rect 10349 7391 10434 7627
rect 10670 7391 10755 7627
rect 10991 7391 11076 7627
rect 11312 7391 11397 7627
rect 11633 7391 11718 7627
rect 11954 7391 12039 7627
rect 12275 7391 12359 7627
rect 12595 7391 12679 7627
rect 12915 7391 12999 7627
rect 13235 7391 13319 7627
rect 13555 7391 13639 7627
rect 13875 7391 13959 7627
rect 14195 7391 14279 7627
rect 14515 7391 14599 7627
rect 14835 7391 14919 7627
rect 15155 7391 15239 7627
rect 15475 7391 15559 7627
rect 15795 7391 16000 7627
rect 0 7347 254 7391
rect 15746 7347 16000 7391
rect 0 7023 254 7067
rect 15746 7023 16000 7067
rect 0 6787 162 7023
rect 398 6787 483 7023
rect 719 6787 804 7023
rect 1040 6787 1125 7023
rect 1361 6787 1446 7023
rect 1682 6787 1767 7023
rect 2003 6787 2088 7023
rect 2324 6787 2409 7023
rect 2645 6787 2730 7023
rect 2966 6787 3051 7023
rect 3287 6787 3372 7023
rect 3608 6787 3693 7023
rect 3929 6787 4014 7023
rect 4250 6787 4335 7023
rect 4571 6787 4656 7023
rect 4892 6787 4977 7023
rect 5213 6787 5298 7023
rect 5534 6787 5619 7023
rect 5855 6787 5940 7023
rect 6176 6787 6261 7023
rect 6497 6787 6582 7023
rect 6818 6787 6903 7023
rect 7139 6787 7224 7023
rect 7460 6787 7545 7023
rect 7781 6787 7866 7023
rect 8102 6787 8187 7023
rect 8423 6787 8508 7023
rect 8744 6787 8829 7023
rect 9065 6787 9150 7023
rect 9386 6787 9471 7023
rect 9707 6787 9792 7023
rect 10028 6787 10113 7023
rect 10349 6787 10434 7023
rect 10670 6787 10755 7023
rect 10991 6787 11076 7023
rect 11312 6787 11397 7023
rect 11633 6787 11718 7023
rect 11954 6787 12038 7023
rect 12274 6787 12358 7023
rect 12594 6787 12678 7023
rect 12914 6787 12998 7023
rect 13234 6787 13318 7023
rect 13554 6787 13638 7023
rect 13874 6787 13958 7023
rect 14194 6787 14278 7023
rect 14514 6787 14598 7023
rect 14834 6787 14918 7023
rect 15154 6787 15238 7023
rect 15474 6787 15558 7023
rect 15794 6787 16000 7023
rect 0 6657 16000 6787
rect 0 6421 162 6657
rect 398 6421 483 6657
rect 719 6421 804 6657
rect 1040 6421 1125 6657
rect 1361 6421 1446 6657
rect 1682 6421 1767 6657
rect 2003 6421 2088 6657
rect 2324 6421 2409 6657
rect 2645 6421 2730 6657
rect 2966 6421 3051 6657
rect 3287 6421 3372 6657
rect 3608 6421 3693 6657
rect 3929 6421 4014 6657
rect 4250 6421 4335 6657
rect 4571 6421 4656 6657
rect 4892 6421 4977 6657
rect 5213 6421 5298 6657
rect 5534 6421 5619 6657
rect 5855 6421 5940 6657
rect 6176 6421 6261 6657
rect 6497 6421 6582 6657
rect 6818 6421 6903 6657
rect 7139 6421 7224 6657
rect 7460 6421 7545 6657
rect 7781 6421 7866 6657
rect 8102 6421 8187 6657
rect 8423 6421 8508 6657
rect 8744 6421 8829 6657
rect 9065 6421 9150 6657
rect 9386 6421 9471 6657
rect 9707 6421 9792 6657
rect 10028 6421 10113 6657
rect 10349 6421 10434 6657
rect 10670 6421 10755 6657
rect 10991 6421 11076 6657
rect 11312 6421 11397 6657
rect 11633 6421 11718 6657
rect 11954 6421 12038 6657
rect 12274 6421 12358 6657
rect 12594 6421 12678 6657
rect 12914 6421 12998 6657
rect 13234 6421 13318 6657
rect 13554 6421 13638 6657
rect 13874 6421 13958 6657
rect 14194 6421 14278 6657
rect 14514 6421 14598 6657
rect 14834 6421 14918 6657
rect 15154 6421 15238 6657
rect 15474 6421 15558 6657
rect 15794 6421 16000 6657
rect 0 6377 254 6421
rect 15746 6377 16000 6421
rect 0 6053 254 6097
rect 15746 6053 16000 6097
rect 0 5817 161 6053
rect 397 5817 482 6053
rect 718 5817 803 6053
rect 1039 5817 1124 6053
rect 1360 5817 1445 6053
rect 1681 5817 1766 6053
rect 2002 5817 2087 6053
rect 2323 5817 2408 6053
rect 2644 5817 2729 6053
rect 2965 5817 3050 6053
rect 3286 5817 3371 6053
rect 3607 5817 3692 6053
rect 3928 5817 4013 6053
rect 4249 5817 4334 6053
rect 4570 5817 4655 6053
rect 4891 5817 4976 6053
rect 5212 5817 5297 6053
rect 5533 5817 5618 6053
rect 5854 5817 5939 6053
rect 6175 5817 6260 6053
rect 6496 5817 6581 6053
rect 6817 5817 6902 6053
rect 7138 5817 7223 6053
rect 7459 5817 7544 6053
rect 7780 5817 7865 6053
rect 8101 5817 8186 6053
rect 8422 5817 8507 6053
rect 8743 5817 8828 6053
rect 9064 5817 9149 6053
rect 9385 5817 9470 6053
rect 9706 5817 9791 6053
rect 10027 5817 10112 6053
rect 10348 5817 10433 6053
rect 10669 5817 10754 6053
rect 10990 5817 11075 6053
rect 11311 5817 11396 6053
rect 11632 5817 11717 6053
rect 11953 5817 12038 6053
rect 12274 5817 12358 6053
rect 12594 5817 12678 6053
rect 12914 5817 12998 6053
rect 13234 5817 13318 6053
rect 13554 5817 13638 6053
rect 13874 5817 13958 6053
rect 14194 5817 14278 6053
rect 14514 5817 14598 6053
rect 14834 5817 14918 6053
rect 15154 5817 15238 6053
rect 15474 5817 15558 6053
rect 15794 5817 16000 6053
rect 0 5447 16000 5817
rect 0 5211 161 5447
rect 397 5211 482 5447
rect 718 5211 803 5447
rect 1039 5211 1124 5447
rect 1360 5211 1445 5447
rect 1681 5211 1766 5447
rect 2002 5211 2087 5447
rect 2323 5211 2408 5447
rect 2644 5211 2729 5447
rect 2965 5211 3050 5447
rect 3286 5211 3371 5447
rect 3607 5211 3692 5447
rect 3928 5211 4013 5447
rect 4249 5211 4334 5447
rect 4570 5211 4655 5447
rect 4891 5211 4976 5447
rect 5212 5211 5297 5447
rect 5533 5211 5618 5447
rect 5854 5211 5939 5447
rect 6175 5211 6260 5447
rect 6496 5211 6581 5447
rect 6817 5211 6902 5447
rect 7138 5211 7223 5447
rect 7459 5211 7544 5447
rect 7780 5211 7865 5447
rect 8101 5211 8186 5447
rect 8422 5211 8507 5447
rect 8743 5211 8828 5447
rect 9064 5211 9149 5447
rect 9385 5211 9470 5447
rect 9706 5211 9791 5447
rect 10027 5211 10112 5447
rect 10348 5211 10433 5447
rect 10669 5211 10754 5447
rect 10990 5211 11075 5447
rect 11311 5211 11396 5447
rect 11632 5211 11717 5447
rect 11953 5211 12038 5447
rect 12274 5211 12358 5447
rect 12594 5211 12678 5447
rect 12914 5211 12998 5447
rect 13234 5211 13318 5447
rect 13554 5211 13638 5447
rect 13874 5211 13958 5447
rect 14194 5211 14278 5447
rect 14514 5211 14598 5447
rect 14834 5211 14918 5447
rect 15154 5211 15238 5447
rect 15474 5211 15558 5447
rect 15794 5211 16000 5447
rect 0 5167 254 5211
rect 15746 5167 16000 5211
rect 0 4843 254 4887
rect 15746 4843 16000 4887
rect 0 4607 161 4843
rect 397 4607 482 4843
rect 718 4607 803 4843
rect 1039 4607 1124 4843
rect 1360 4607 1445 4843
rect 1681 4607 1766 4843
rect 2002 4607 2087 4843
rect 2323 4607 2408 4843
rect 2644 4607 2729 4843
rect 2965 4607 3050 4843
rect 3286 4607 3371 4843
rect 3607 4607 3692 4843
rect 3928 4607 4013 4843
rect 4249 4607 4334 4843
rect 4570 4607 4655 4843
rect 4891 4607 4976 4843
rect 5212 4607 5297 4843
rect 5533 4607 5618 4843
rect 5854 4607 5939 4843
rect 6175 4607 6260 4843
rect 6496 4607 6581 4843
rect 6817 4607 6902 4843
rect 7138 4607 7223 4843
rect 7459 4607 7544 4843
rect 7780 4607 7865 4843
rect 8101 4607 8186 4843
rect 8422 4607 8507 4843
rect 8743 4607 8828 4843
rect 9064 4607 9149 4843
rect 9385 4607 9470 4843
rect 9706 4607 9791 4843
rect 10027 4607 10112 4843
rect 10348 4607 10433 4843
rect 10669 4607 10754 4843
rect 10990 4607 11075 4843
rect 11311 4607 11396 4843
rect 11632 4607 11717 4843
rect 11953 4607 12037 4843
rect 12273 4607 12357 4843
rect 12593 4607 12677 4843
rect 12913 4607 12997 4843
rect 13233 4607 13317 4843
rect 13553 4607 13637 4843
rect 13873 4607 13957 4843
rect 14193 4607 14277 4843
rect 14513 4607 14597 4843
rect 14833 4607 14917 4843
rect 15153 4607 15237 4843
rect 15473 4607 15557 4843
rect 15793 4607 16000 4843
rect 0 4237 16000 4607
rect 0 4001 161 4237
rect 397 4001 482 4237
rect 718 4001 803 4237
rect 1039 4001 1124 4237
rect 1360 4001 1445 4237
rect 1681 4001 1766 4237
rect 2002 4001 2087 4237
rect 2323 4001 2408 4237
rect 2644 4001 2729 4237
rect 2965 4001 3050 4237
rect 3286 4001 3371 4237
rect 3607 4001 3692 4237
rect 3928 4001 4013 4237
rect 4249 4001 4334 4237
rect 4570 4001 4655 4237
rect 4891 4001 4976 4237
rect 5212 4001 5297 4237
rect 5533 4001 5618 4237
rect 5854 4001 5939 4237
rect 6175 4001 6260 4237
rect 6496 4001 6581 4237
rect 6817 4001 6902 4237
rect 7138 4001 7223 4237
rect 7459 4001 7544 4237
rect 7780 4001 7865 4237
rect 8101 4001 8186 4237
rect 8422 4001 8507 4237
rect 8743 4001 8828 4237
rect 9064 4001 9149 4237
rect 9385 4001 9470 4237
rect 9706 4001 9791 4237
rect 10027 4001 10112 4237
rect 10348 4001 10433 4237
rect 10669 4001 10754 4237
rect 10990 4001 11075 4237
rect 11311 4001 11396 4237
rect 11632 4001 11717 4237
rect 11953 4001 12037 4237
rect 12273 4001 12357 4237
rect 12593 4001 12677 4237
rect 12913 4001 12997 4237
rect 13233 4001 13317 4237
rect 13553 4001 13637 4237
rect 13873 4001 13957 4237
rect 14193 4001 14277 4237
rect 14513 4001 14597 4237
rect 14833 4001 14917 4237
rect 15153 4001 15237 4237
rect 15473 4001 15557 4237
rect 15793 4001 16000 4237
rect 0 3957 254 4001
rect 15746 3957 16000 4001
rect 0 3633 193 3677
rect 0 3397 162 3633
rect 398 3397 483 3633
rect 719 3397 804 3633
rect 1040 3397 1125 3633
rect 1361 3397 1446 3633
rect 1682 3397 1767 3633
rect 2003 3397 2088 3633
rect 2324 3397 2409 3633
rect 2645 3397 2730 3633
rect 2966 3397 3051 3633
rect 3287 3397 3372 3633
rect 3608 3397 3693 3633
rect 3929 3397 4014 3633
rect 4250 3397 4335 3633
rect 4571 3397 4656 3633
rect 4892 3397 4977 3633
rect 5213 3397 5298 3633
rect 5534 3397 5619 3633
rect 5855 3397 5940 3633
rect 6176 3397 6261 3633
rect 6497 3397 6582 3633
rect 6818 3397 6903 3633
rect 7139 3397 7224 3633
rect 7460 3397 7545 3633
rect 7781 3397 7866 3633
rect 8102 3397 8187 3633
rect 8423 3397 8508 3633
rect 8744 3397 8829 3633
rect 9065 3397 9150 3633
rect 9386 3397 9471 3633
rect 9707 3397 9792 3633
rect 10028 3397 10113 3633
rect 10349 3397 10434 3633
rect 10670 3397 10755 3633
rect 10991 3397 11076 3633
rect 11312 3397 11397 3633
rect 11633 3397 11718 3633
rect 11954 3397 12038 3633
rect 12274 3397 12358 3633
rect 12594 3397 12678 3633
rect 12914 3397 12998 3633
rect 13234 3397 13318 3633
rect 13554 3397 13638 3633
rect 13874 3397 13958 3633
rect 14194 3397 14278 3633
rect 14514 3397 14598 3633
rect 14834 3397 14918 3633
rect 15154 3397 15238 3633
rect 15474 3397 15558 3633
rect 0 3267 15794 3397
rect 0 3031 162 3267
rect 398 3031 483 3267
rect 719 3031 804 3267
rect 1040 3031 1125 3267
rect 1361 3031 1446 3267
rect 1682 3031 1767 3267
rect 2003 3031 2088 3267
rect 2324 3031 2409 3267
rect 2645 3031 2730 3267
rect 2966 3031 3051 3267
rect 3287 3031 3372 3267
rect 3608 3031 3693 3267
rect 3929 3031 4014 3267
rect 4250 3031 4335 3267
rect 4571 3031 4656 3267
rect 4892 3031 4977 3267
rect 5213 3031 5298 3267
rect 5534 3031 5619 3267
rect 5855 3031 5940 3267
rect 6176 3031 6261 3267
rect 6497 3031 6582 3267
rect 6818 3031 6903 3267
rect 7139 3031 7224 3267
rect 7460 3031 7545 3267
rect 7781 3031 7866 3267
rect 8102 3031 8187 3267
rect 8423 3031 8508 3267
rect 8744 3031 8829 3267
rect 9065 3031 9150 3267
rect 9386 3031 9471 3267
rect 9707 3031 9792 3267
rect 10028 3031 10113 3267
rect 10349 3031 10434 3267
rect 10670 3031 10755 3267
rect 10991 3031 11076 3267
rect 11312 3031 11397 3267
rect 11633 3031 11718 3267
rect 11954 3031 12038 3267
rect 12274 3031 12358 3267
rect 12594 3031 12678 3267
rect 12914 3031 12998 3267
rect 13234 3031 13318 3267
rect 13554 3031 13638 3267
rect 13874 3031 13958 3267
rect 14194 3031 14278 3267
rect 14514 3031 14598 3267
rect 14834 3031 14918 3267
rect 15154 3031 15238 3267
rect 15474 3031 15558 3267
rect 0 2987 193 3031
rect 15807 2987 16000 3677
rect 0 2663 254 2707
rect 15746 2663 16000 2707
rect 0 2427 163 2663
rect 399 2427 484 2663
rect 720 2427 805 2663
rect 1041 2427 1126 2663
rect 1362 2427 1447 2663
rect 1683 2427 1768 2663
rect 2004 2427 2089 2663
rect 2325 2427 2410 2663
rect 2646 2427 2731 2663
rect 2967 2427 3052 2663
rect 3288 2427 3373 2663
rect 3609 2427 3694 2663
rect 3930 2427 4015 2663
rect 4251 2427 4336 2663
rect 4572 2427 4657 2663
rect 4893 2427 4978 2663
rect 5214 2427 5299 2663
rect 5535 2427 5620 2663
rect 5856 2427 5941 2663
rect 6177 2427 6262 2663
rect 6498 2427 6583 2663
rect 6819 2427 6904 2663
rect 7140 2427 7225 2663
rect 7461 2427 7546 2663
rect 7782 2427 7867 2663
rect 8103 2427 8188 2663
rect 8424 2427 8509 2663
rect 8745 2427 8830 2663
rect 9066 2427 9151 2663
rect 9387 2427 9472 2663
rect 9708 2427 9793 2663
rect 10029 2427 10114 2663
rect 10350 2427 10435 2663
rect 10671 2427 10756 2663
rect 10992 2427 11077 2663
rect 11313 2427 11397 2663
rect 11633 2427 11717 2663
rect 11953 2427 12037 2663
rect 12273 2427 12357 2663
rect 12593 2427 12677 2663
rect 12913 2427 12997 2663
rect 13233 2427 13317 2663
rect 13553 2427 13637 2663
rect 13873 2427 13957 2663
rect 14193 2427 14277 2663
rect 14513 2427 14597 2663
rect 14833 2427 14917 2663
rect 15153 2427 15237 2663
rect 15473 2427 15557 2663
rect 15793 2427 16000 2663
rect 0 2057 16000 2427
rect 0 1821 163 2057
rect 399 1821 484 2057
rect 720 1821 805 2057
rect 1041 1821 1126 2057
rect 1362 1821 1447 2057
rect 1683 1821 1768 2057
rect 2004 1821 2089 2057
rect 2325 1821 2410 2057
rect 2646 1821 2731 2057
rect 2967 1821 3052 2057
rect 3288 1821 3373 2057
rect 3609 1821 3694 2057
rect 3930 1821 4015 2057
rect 4251 1821 4336 2057
rect 4572 1821 4657 2057
rect 4893 1821 4978 2057
rect 5214 1821 5299 2057
rect 5535 1821 5620 2057
rect 5856 1821 5941 2057
rect 6177 1821 6262 2057
rect 6498 1821 6583 2057
rect 6819 1821 6904 2057
rect 7140 1821 7225 2057
rect 7461 1821 7546 2057
rect 7782 1821 7867 2057
rect 8103 1821 8188 2057
rect 8424 1821 8509 2057
rect 8745 1821 8830 2057
rect 9066 1821 9151 2057
rect 9387 1821 9472 2057
rect 9708 1821 9793 2057
rect 10029 1821 10114 2057
rect 10350 1821 10435 2057
rect 10671 1821 10756 2057
rect 10992 1821 11077 2057
rect 11313 1821 11397 2057
rect 11633 1821 11717 2057
rect 11953 1821 12037 2057
rect 12273 1821 12357 2057
rect 12593 1821 12677 2057
rect 12913 1821 12997 2057
rect 13233 1821 13317 2057
rect 13553 1821 13637 2057
rect 13873 1821 13957 2057
rect 14193 1821 14277 2057
rect 14513 1821 14597 2057
rect 14833 1821 14917 2057
rect 15153 1821 15237 2057
rect 15473 1821 15557 2057
rect 15793 1821 16000 2057
rect 0 1777 254 1821
rect 15746 1777 16000 1821
rect 0 1453 254 1497
rect 15746 1453 16000 1497
rect 0 1452 16000 1453
rect 0 1216 162 1452
rect 398 1216 483 1452
rect 719 1216 804 1452
rect 1040 1216 1125 1452
rect 1361 1216 1446 1452
rect 1682 1216 1767 1452
rect 2003 1216 2088 1452
rect 2324 1216 2409 1452
rect 2645 1216 2730 1452
rect 2966 1216 3051 1452
rect 3287 1216 3372 1452
rect 3608 1216 3693 1452
rect 3929 1216 4014 1452
rect 4250 1216 4335 1452
rect 4571 1216 4656 1452
rect 4892 1216 4977 1452
rect 5213 1216 5298 1452
rect 5534 1216 5619 1452
rect 5855 1216 5940 1452
rect 6176 1216 6261 1452
rect 6497 1216 6582 1452
rect 6818 1216 6903 1452
rect 7139 1216 7224 1452
rect 7460 1216 7545 1452
rect 7781 1216 7866 1452
rect 8102 1216 8187 1452
rect 8423 1216 8508 1452
rect 8744 1216 8829 1452
rect 9065 1216 9150 1452
rect 9386 1216 9471 1452
rect 9707 1216 9792 1452
rect 10028 1216 10113 1452
rect 10349 1216 10434 1452
rect 10670 1216 10755 1452
rect 10991 1216 11076 1452
rect 11312 1216 11397 1452
rect 11633 1216 11718 1452
rect 11954 1216 12038 1452
rect 12274 1216 12358 1452
rect 12594 1216 12678 1452
rect 12914 1216 12998 1452
rect 13234 1216 13318 1452
rect 13554 1216 13638 1452
rect 13874 1216 13958 1452
rect 14194 1216 14278 1452
rect 14514 1216 14598 1452
rect 14834 1216 14918 1452
rect 15154 1216 15238 1452
rect 15474 1216 15558 1452
rect 15794 1216 16000 1452
rect 0 1070 16000 1216
rect 0 834 162 1070
rect 398 834 483 1070
rect 719 834 804 1070
rect 1040 834 1125 1070
rect 1361 834 1446 1070
rect 1682 834 1767 1070
rect 2003 834 2088 1070
rect 2324 834 2409 1070
rect 2645 834 2730 1070
rect 2966 834 3051 1070
rect 3287 834 3372 1070
rect 3608 834 3693 1070
rect 3929 834 4014 1070
rect 4250 834 4335 1070
rect 4571 834 4656 1070
rect 4892 834 4977 1070
rect 5213 834 5298 1070
rect 5534 834 5619 1070
rect 5855 834 5940 1070
rect 6176 834 6261 1070
rect 6497 834 6582 1070
rect 6818 834 6903 1070
rect 7139 834 7224 1070
rect 7460 834 7545 1070
rect 7781 834 7866 1070
rect 8102 834 8187 1070
rect 8423 834 8508 1070
rect 8744 834 8829 1070
rect 9065 834 9150 1070
rect 9386 834 9471 1070
rect 9707 834 9792 1070
rect 10028 834 10113 1070
rect 10349 834 10434 1070
rect 10670 834 10755 1070
rect 10991 834 11076 1070
rect 11312 834 11397 1070
rect 11633 834 11718 1070
rect 11954 834 12038 1070
rect 12274 834 12358 1070
rect 12594 834 12678 1070
rect 12914 834 12998 1070
rect 13234 834 13318 1070
rect 13554 834 13638 1070
rect 13874 834 13958 1070
rect 14194 834 14278 1070
rect 14514 834 14598 1070
rect 14834 834 14918 1070
rect 15154 834 15238 1070
rect 15474 834 15558 1070
rect 15794 834 16000 1070
rect 0 688 16000 834
rect 0 452 162 688
rect 398 452 483 688
rect 719 452 804 688
rect 1040 452 1125 688
rect 1361 452 1446 688
rect 1682 452 1767 688
rect 2003 452 2088 688
rect 2324 452 2409 688
rect 2645 452 2730 688
rect 2966 452 3051 688
rect 3287 452 3372 688
rect 3608 452 3693 688
rect 3929 452 4014 688
rect 4250 452 4335 688
rect 4571 452 4656 688
rect 4892 452 4977 688
rect 5213 452 5298 688
rect 5534 452 5619 688
rect 5855 452 5940 688
rect 6176 452 6261 688
rect 6497 452 6582 688
rect 6818 452 6903 688
rect 7139 452 7224 688
rect 7460 452 7545 688
rect 7781 452 7866 688
rect 8102 452 8187 688
rect 8423 452 8508 688
rect 8744 452 8829 688
rect 9065 452 9150 688
rect 9386 452 9471 688
rect 9707 452 9792 688
rect 10028 452 10113 688
rect 10349 452 10434 688
rect 10670 452 10755 688
rect 10991 452 11076 688
rect 11312 452 11397 688
rect 11633 452 11718 688
rect 11954 452 12038 688
rect 12274 452 12358 688
rect 12594 452 12678 688
rect 12914 452 12998 688
rect 13234 452 13318 688
rect 13554 452 13638 688
rect 13874 452 13958 688
rect 14194 452 14278 688
rect 14514 452 14598 688
rect 14834 452 14918 688
rect 15154 452 15238 688
rect 15474 452 15558 688
rect 15794 452 16000 688
rect 0 451 16000 452
rect 0 407 254 451
rect 15746 407 16000 451
<< via4 >>
rect 162 39729 398 39965
rect 483 39729 719 39965
rect 804 39729 1040 39965
rect 1125 39729 1361 39965
rect 1446 39729 1682 39965
rect 1767 39729 2003 39965
rect 2088 39729 2324 39965
rect 2409 39729 2645 39965
rect 2730 39729 2966 39965
rect 3051 39729 3287 39965
rect 3372 39729 3608 39965
rect 3693 39729 3929 39965
rect 4014 39729 4250 39965
rect 4335 39729 4571 39965
rect 4656 39729 4892 39965
rect 4977 39729 5213 39965
rect 5298 39729 5534 39965
rect 5619 39729 5855 39965
rect 5940 39729 6176 39965
rect 6261 39729 6497 39965
rect 6582 39729 6818 39965
rect 6903 39729 7139 39965
rect 7224 39729 7460 39965
rect 7545 39729 7781 39965
rect 7866 39729 8102 39965
rect 8187 39729 8423 39965
rect 8508 39729 8744 39965
rect 8829 39729 9065 39965
rect 9150 39729 9386 39965
rect 9471 39729 9707 39965
rect 9792 39729 10028 39965
rect 10113 39729 10349 39965
rect 10434 39729 10670 39965
rect 10755 39729 10991 39965
rect 11076 39729 11312 39965
rect 11397 39729 11633 39965
rect 11718 39729 11954 39965
rect 12038 39729 12274 39965
rect 12358 39729 12594 39965
rect 12678 39729 12914 39965
rect 12998 39729 13234 39965
rect 13318 39729 13554 39965
rect 13638 39729 13874 39965
rect 13958 39729 14194 39965
rect 14278 39729 14514 39965
rect 14598 39729 14834 39965
rect 14918 39729 15154 39965
rect 15238 39729 15474 39965
rect 15558 39729 15794 39965
rect 162 39405 398 39641
rect 483 39405 719 39641
rect 804 39405 1040 39641
rect 1125 39405 1361 39641
rect 1446 39405 1682 39641
rect 1767 39405 2003 39641
rect 2088 39405 2324 39641
rect 2409 39405 2645 39641
rect 2730 39405 2966 39641
rect 3051 39405 3287 39641
rect 3372 39405 3608 39641
rect 3693 39405 3929 39641
rect 4014 39405 4250 39641
rect 4335 39405 4571 39641
rect 4656 39405 4892 39641
rect 4977 39405 5213 39641
rect 5298 39405 5534 39641
rect 5619 39405 5855 39641
rect 5940 39405 6176 39641
rect 6261 39405 6497 39641
rect 6582 39405 6818 39641
rect 6903 39405 7139 39641
rect 7224 39405 7460 39641
rect 7545 39405 7781 39641
rect 7866 39405 8102 39641
rect 8187 39405 8423 39641
rect 8508 39405 8744 39641
rect 8829 39405 9065 39641
rect 9150 39405 9386 39641
rect 9471 39405 9707 39641
rect 9792 39405 10028 39641
rect 10113 39405 10349 39641
rect 10434 39405 10670 39641
rect 10755 39405 10991 39641
rect 11076 39405 11312 39641
rect 11397 39405 11633 39641
rect 11718 39405 11954 39641
rect 12038 39405 12274 39641
rect 12358 39405 12594 39641
rect 12678 39405 12914 39641
rect 12998 39405 13234 39641
rect 13318 39405 13554 39641
rect 13638 39405 13874 39641
rect 13958 39405 14194 39641
rect 14278 39405 14514 39641
rect 14598 39405 14834 39641
rect 14918 39405 15154 39641
rect 15238 39405 15474 39641
rect 15558 39405 15794 39641
rect 162 39081 398 39317
rect 483 39081 719 39317
rect 804 39081 1040 39317
rect 1125 39081 1361 39317
rect 1446 39081 1682 39317
rect 1767 39081 2003 39317
rect 2088 39081 2324 39317
rect 2409 39081 2645 39317
rect 2730 39081 2966 39317
rect 3051 39081 3287 39317
rect 3372 39081 3608 39317
rect 3693 39081 3929 39317
rect 4014 39081 4250 39317
rect 4335 39081 4571 39317
rect 4656 39081 4892 39317
rect 4977 39081 5213 39317
rect 5298 39081 5534 39317
rect 5619 39081 5855 39317
rect 5940 39081 6176 39317
rect 6261 39081 6497 39317
rect 6582 39081 6818 39317
rect 6903 39081 7139 39317
rect 7224 39081 7460 39317
rect 7545 39081 7781 39317
rect 7866 39081 8102 39317
rect 8187 39081 8423 39317
rect 8508 39081 8744 39317
rect 8829 39081 9065 39317
rect 9150 39081 9386 39317
rect 9471 39081 9707 39317
rect 9792 39081 10028 39317
rect 10113 39081 10349 39317
rect 10434 39081 10670 39317
rect 10755 39081 10991 39317
rect 11076 39081 11312 39317
rect 11397 39081 11633 39317
rect 11718 39081 11954 39317
rect 12038 39081 12274 39317
rect 12358 39081 12594 39317
rect 12678 39081 12914 39317
rect 12998 39081 13234 39317
rect 13318 39081 13554 39317
rect 13638 39081 13874 39317
rect 13958 39081 14194 39317
rect 14278 39081 14514 39317
rect 14598 39081 14834 39317
rect 14918 39081 15154 39317
rect 15238 39081 15474 39317
rect 15558 39081 15794 39317
rect 162 38757 398 38993
rect 483 38757 719 38993
rect 804 38757 1040 38993
rect 1125 38757 1361 38993
rect 1446 38757 1682 38993
rect 1767 38757 2003 38993
rect 2088 38757 2324 38993
rect 2409 38757 2645 38993
rect 2730 38757 2966 38993
rect 3051 38757 3287 38993
rect 3372 38757 3608 38993
rect 3693 38757 3929 38993
rect 4014 38757 4250 38993
rect 4335 38757 4571 38993
rect 4656 38757 4892 38993
rect 4977 38757 5213 38993
rect 5298 38757 5534 38993
rect 5619 38757 5855 38993
rect 5940 38757 6176 38993
rect 6261 38757 6497 38993
rect 6582 38757 6818 38993
rect 6903 38757 7139 38993
rect 7224 38757 7460 38993
rect 7545 38757 7781 38993
rect 7866 38757 8102 38993
rect 8187 38757 8423 38993
rect 8508 38757 8744 38993
rect 8829 38757 9065 38993
rect 9150 38757 9386 38993
rect 9471 38757 9707 38993
rect 9792 38757 10028 38993
rect 10113 38757 10349 38993
rect 10434 38757 10670 38993
rect 10755 38757 10991 38993
rect 11076 38757 11312 38993
rect 11397 38757 11633 38993
rect 11718 38757 11954 38993
rect 12038 38757 12274 38993
rect 12358 38757 12594 38993
rect 12678 38757 12914 38993
rect 12998 38757 13234 38993
rect 13318 38757 13554 38993
rect 13638 38757 13874 38993
rect 13958 38757 14194 38993
rect 14278 38757 14514 38993
rect 14598 38757 14834 38993
rect 14918 38757 15154 38993
rect 15238 38757 15474 38993
rect 15558 38757 15794 38993
rect 162 38433 398 38669
rect 483 38433 719 38669
rect 804 38433 1040 38669
rect 1125 38433 1361 38669
rect 1446 38433 1682 38669
rect 1767 38433 2003 38669
rect 2088 38433 2324 38669
rect 2409 38433 2645 38669
rect 2730 38433 2966 38669
rect 3051 38433 3287 38669
rect 3372 38433 3608 38669
rect 3693 38433 3929 38669
rect 4014 38433 4250 38669
rect 4335 38433 4571 38669
rect 4656 38433 4892 38669
rect 4977 38433 5213 38669
rect 5298 38433 5534 38669
rect 5619 38433 5855 38669
rect 5940 38433 6176 38669
rect 6261 38433 6497 38669
rect 6582 38433 6818 38669
rect 6903 38433 7139 38669
rect 7224 38433 7460 38669
rect 7545 38433 7781 38669
rect 7866 38433 8102 38669
rect 8187 38433 8423 38669
rect 8508 38433 8744 38669
rect 8829 38433 9065 38669
rect 9150 38433 9386 38669
rect 9471 38433 9707 38669
rect 9792 38433 10028 38669
rect 10113 38433 10349 38669
rect 10434 38433 10670 38669
rect 10755 38433 10991 38669
rect 11076 38433 11312 38669
rect 11397 38433 11633 38669
rect 11718 38433 11954 38669
rect 12038 38433 12274 38669
rect 12358 38433 12594 38669
rect 12678 38433 12914 38669
rect 12998 38433 13234 38669
rect 13318 38433 13554 38669
rect 13638 38433 13874 38669
rect 13958 38433 14194 38669
rect 14278 38433 14514 38669
rect 14598 38433 14834 38669
rect 14918 38433 15154 38669
rect 15238 38433 15474 38669
rect 15558 38433 15794 38669
rect 162 38109 398 38345
rect 483 38109 719 38345
rect 804 38109 1040 38345
rect 1125 38109 1361 38345
rect 1446 38109 1682 38345
rect 1767 38109 2003 38345
rect 2088 38109 2324 38345
rect 2409 38109 2645 38345
rect 2730 38109 2966 38345
rect 3051 38109 3287 38345
rect 3372 38109 3608 38345
rect 3693 38109 3929 38345
rect 4014 38109 4250 38345
rect 4335 38109 4571 38345
rect 4656 38109 4892 38345
rect 4977 38109 5213 38345
rect 5298 38109 5534 38345
rect 5619 38109 5855 38345
rect 5940 38109 6176 38345
rect 6261 38109 6497 38345
rect 6582 38109 6818 38345
rect 6903 38109 7139 38345
rect 7224 38109 7460 38345
rect 7545 38109 7781 38345
rect 7866 38109 8102 38345
rect 8187 38109 8423 38345
rect 8508 38109 8744 38345
rect 8829 38109 9065 38345
rect 9150 38109 9386 38345
rect 9471 38109 9707 38345
rect 9792 38109 10028 38345
rect 10113 38109 10349 38345
rect 10434 38109 10670 38345
rect 10755 38109 10991 38345
rect 11076 38109 11312 38345
rect 11397 38109 11633 38345
rect 11718 38109 11954 38345
rect 12038 38109 12274 38345
rect 12358 38109 12594 38345
rect 12678 38109 12914 38345
rect 12998 38109 13234 38345
rect 13318 38109 13554 38345
rect 13638 38109 13874 38345
rect 13958 38109 14194 38345
rect 14278 38109 14514 38345
rect 14598 38109 14834 38345
rect 14918 38109 15154 38345
rect 15238 38109 15474 38345
rect 15558 38109 15794 38345
rect 162 37785 398 38021
rect 483 37785 719 38021
rect 804 37785 1040 38021
rect 1125 37785 1361 38021
rect 1446 37785 1682 38021
rect 1767 37785 2003 38021
rect 2088 37785 2324 38021
rect 2409 37785 2645 38021
rect 2730 37785 2966 38021
rect 3051 37785 3287 38021
rect 3372 37785 3608 38021
rect 3693 37785 3929 38021
rect 4014 37785 4250 38021
rect 4335 37785 4571 38021
rect 4656 37785 4892 38021
rect 4977 37785 5213 38021
rect 5298 37785 5534 38021
rect 5619 37785 5855 38021
rect 5940 37785 6176 38021
rect 6261 37785 6497 38021
rect 6582 37785 6818 38021
rect 6903 37785 7139 38021
rect 7224 37785 7460 38021
rect 7545 37785 7781 38021
rect 7866 37785 8102 38021
rect 8187 37785 8423 38021
rect 8508 37785 8744 38021
rect 8829 37785 9065 38021
rect 9150 37785 9386 38021
rect 9471 37785 9707 38021
rect 9792 37785 10028 38021
rect 10113 37785 10349 38021
rect 10434 37785 10670 38021
rect 10755 37785 10991 38021
rect 11076 37785 11312 38021
rect 11397 37785 11633 38021
rect 11718 37785 11954 38021
rect 12038 37785 12274 38021
rect 12358 37785 12594 38021
rect 12678 37785 12914 38021
rect 12998 37785 13234 38021
rect 13318 37785 13554 38021
rect 13638 37785 13874 38021
rect 13958 37785 14194 38021
rect 14278 37785 14514 38021
rect 14598 37785 14834 38021
rect 14918 37785 15154 38021
rect 15238 37785 15474 38021
rect 15558 37785 15794 38021
rect 162 37461 398 37697
rect 483 37461 719 37697
rect 804 37461 1040 37697
rect 1125 37461 1361 37697
rect 1446 37461 1682 37697
rect 1767 37461 2003 37697
rect 2088 37461 2324 37697
rect 2409 37461 2645 37697
rect 2730 37461 2966 37697
rect 3051 37461 3287 37697
rect 3372 37461 3608 37697
rect 3693 37461 3929 37697
rect 4014 37461 4250 37697
rect 4335 37461 4571 37697
rect 4656 37461 4892 37697
rect 4977 37461 5213 37697
rect 5298 37461 5534 37697
rect 5619 37461 5855 37697
rect 5940 37461 6176 37697
rect 6261 37461 6497 37697
rect 6582 37461 6818 37697
rect 6903 37461 7139 37697
rect 7224 37461 7460 37697
rect 7545 37461 7781 37697
rect 7866 37461 8102 37697
rect 8187 37461 8423 37697
rect 8508 37461 8744 37697
rect 8829 37461 9065 37697
rect 9150 37461 9386 37697
rect 9471 37461 9707 37697
rect 9792 37461 10028 37697
rect 10113 37461 10349 37697
rect 10434 37461 10670 37697
rect 10755 37461 10991 37697
rect 11076 37461 11312 37697
rect 11397 37461 11633 37697
rect 11718 37461 11954 37697
rect 12038 37461 12274 37697
rect 12358 37461 12594 37697
rect 12678 37461 12914 37697
rect 12998 37461 13234 37697
rect 13318 37461 13554 37697
rect 13638 37461 13874 37697
rect 13958 37461 14194 37697
rect 14278 37461 14514 37697
rect 14598 37461 14834 37697
rect 14918 37461 15154 37697
rect 15238 37461 15474 37697
rect 15558 37461 15794 37697
rect 162 37137 398 37373
rect 483 37137 719 37373
rect 804 37137 1040 37373
rect 1125 37137 1361 37373
rect 1446 37137 1682 37373
rect 1767 37137 2003 37373
rect 2088 37137 2324 37373
rect 2409 37137 2645 37373
rect 2730 37137 2966 37373
rect 3051 37137 3287 37373
rect 3372 37137 3608 37373
rect 3693 37137 3929 37373
rect 4014 37137 4250 37373
rect 4335 37137 4571 37373
rect 4656 37137 4892 37373
rect 4977 37137 5213 37373
rect 5298 37137 5534 37373
rect 5619 37137 5855 37373
rect 5940 37137 6176 37373
rect 6261 37137 6497 37373
rect 6582 37137 6818 37373
rect 6903 37137 7139 37373
rect 7224 37137 7460 37373
rect 7545 37137 7781 37373
rect 7866 37137 8102 37373
rect 8187 37137 8423 37373
rect 8508 37137 8744 37373
rect 8829 37137 9065 37373
rect 9150 37137 9386 37373
rect 9471 37137 9707 37373
rect 9792 37137 10028 37373
rect 10113 37137 10349 37373
rect 10434 37137 10670 37373
rect 10755 37137 10991 37373
rect 11076 37137 11312 37373
rect 11397 37137 11633 37373
rect 11718 37137 11954 37373
rect 12038 37137 12274 37373
rect 12358 37137 12594 37373
rect 12678 37137 12914 37373
rect 12998 37137 13234 37373
rect 13318 37137 13554 37373
rect 13638 37137 13874 37373
rect 13958 37137 14194 37373
rect 14278 37137 14514 37373
rect 14598 37137 14834 37373
rect 14918 37137 15154 37373
rect 15238 37137 15474 37373
rect 15558 37137 15794 37373
rect 162 36813 398 37049
rect 483 36813 719 37049
rect 804 36813 1040 37049
rect 1125 36813 1361 37049
rect 1446 36813 1682 37049
rect 1767 36813 2003 37049
rect 2088 36813 2324 37049
rect 2409 36813 2645 37049
rect 2730 36813 2966 37049
rect 3051 36813 3287 37049
rect 3372 36813 3608 37049
rect 3693 36813 3929 37049
rect 4014 36813 4250 37049
rect 4335 36813 4571 37049
rect 4656 36813 4892 37049
rect 4977 36813 5213 37049
rect 5298 36813 5534 37049
rect 5619 36813 5855 37049
rect 5940 36813 6176 37049
rect 6261 36813 6497 37049
rect 6582 36813 6818 37049
rect 6903 36813 7139 37049
rect 7224 36813 7460 37049
rect 7545 36813 7781 37049
rect 7866 36813 8102 37049
rect 8187 36813 8423 37049
rect 8508 36813 8744 37049
rect 8829 36813 9065 37049
rect 9150 36813 9386 37049
rect 9471 36813 9707 37049
rect 9792 36813 10028 37049
rect 10113 36813 10349 37049
rect 10434 36813 10670 37049
rect 10755 36813 10991 37049
rect 11076 36813 11312 37049
rect 11397 36813 11633 37049
rect 11718 36813 11954 37049
rect 12038 36813 12274 37049
rect 12358 36813 12594 37049
rect 12678 36813 12914 37049
rect 12998 36813 13234 37049
rect 13318 36813 13554 37049
rect 13638 36813 13874 37049
rect 13958 36813 14194 37049
rect 14278 36813 14514 37049
rect 14598 36813 14834 37049
rect 14918 36813 15154 37049
rect 15238 36813 15474 37049
rect 15558 36813 15794 37049
rect 162 36489 398 36725
rect 483 36489 719 36725
rect 804 36489 1040 36725
rect 1125 36489 1361 36725
rect 1446 36489 1682 36725
rect 1767 36489 2003 36725
rect 2088 36489 2324 36725
rect 2409 36489 2645 36725
rect 2730 36489 2966 36725
rect 3051 36489 3287 36725
rect 3372 36489 3608 36725
rect 3693 36489 3929 36725
rect 4014 36489 4250 36725
rect 4335 36489 4571 36725
rect 4656 36489 4892 36725
rect 4977 36489 5213 36725
rect 5298 36489 5534 36725
rect 5619 36489 5855 36725
rect 5940 36489 6176 36725
rect 6261 36489 6497 36725
rect 6582 36489 6818 36725
rect 6903 36489 7139 36725
rect 7224 36489 7460 36725
rect 7545 36489 7781 36725
rect 7866 36489 8102 36725
rect 8187 36489 8423 36725
rect 8508 36489 8744 36725
rect 8829 36489 9065 36725
rect 9150 36489 9386 36725
rect 9471 36489 9707 36725
rect 9792 36489 10028 36725
rect 10113 36489 10349 36725
rect 10434 36489 10670 36725
rect 10755 36489 10991 36725
rect 11076 36489 11312 36725
rect 11397 36489 11633 36725
rect 11718 36489 11954 36725
rect 12038 36489 12274 36725
rect 12358 36489 12594 36725
rect 12678 36489 12914 36725
rect 12998 36489 13234 36725
rect 13318 36489 13554 36725
rect 13638 36489 13874 36725
rect 13958 36489 14194 36725
rect 14278 36489 14514 36725
rect 14598 36489 14834 36725
rect 14918 36489 15154 36725
rect 15238 36489 15474 36725
rect 15558 36489 15794 36725
rect 162 36165 398 36401
rect 483 36165 719 36401
rect 804 36165 1040 36401
rect 1125 36165 1361 36401
rect 1446 36165 1682 36401
rect 1767 36165 2003 36401
rect 2088 36165 2324 36401
rect 2409 36165 2645 36401
rect 2730 36165 2966 36401
rect 3051 36165 3287 36401
rect 3372 36165 3608 36401
rect 3693 36165 3929 36401
rect 4014 36165 4250 36401
rect 4335 36165 4571 36401
rect 4656 36165 4892 36401
rect 4977 36165 5213 36401
rect 5298 36165 5534 36401
rect 5619 36165 5855 36401
rect 5940 36165 6176 36401
rect 6261 36165 6497 36401
rect 6582 36165 6818 36401
rect 6903 36165 7139 36401
rect 7224 36165 7460 36401
rect 7545 36165 7781 36401
rect 7866 36165 8102 36401
rect 8187 36165 8423 36401
rect 8508 36165 8744 36401
rect 8829 36165 9065 36401
rect 9150 36165 9386 36401
rect 9471 36165 9707 36401
rect 9792 36165 10028 36401
rect 10113 36165 10349 36401
rect 10434 36165 10670 36401
rect 10755 36165 10991 36401
rect 11076 36165 11312 36401
rect 11397 36165 11633 36401
rect 11718 36165 11954 36401
rect 12038 36165 12274 36401
rect 12358 36165 12594 36401
rect 12678 36165 12914 36401
rect 12998 36165 13234 36401
rect 13318 36165 13554 36401
rect 13638 36165 13874 36401
rect 13958 36165 14194 36401
rect 14278 36165 14514 36401
rect 14598 36165 14834 36401
rect 14918 36165 15154 36401
rect 15238 36165 15474 36401
rect 15558 36165 15794 36401
rect 162 35841 398 36077
rect 483 35841 719 36077
rect 804 35841 1040 36077
rect 1125 35841 1361 36077
rect 1446 35841 1682 36077
rect 1767 35841 2003 36077
rect 2088 35841 2324 36077
rect 2409 35841 2645 36077
rect 2730 35841 2966 36077
rect 3051 35841 3287 36077
rect 3372 35841 3608 36077
rect 3693 35841 3929 36077
rect 4014 35841 4250 36077
rect 4335 35841 4571 36077
rect 4656 35841 4892 36077
rect 4977 35841 5213 36077
rect 5298 35841 5534 36077
rect 5619 35841 5855 36077
rect 5940 35841 6176 36077
rect 6261 35841 6497 36077
rect 6582 35841 6818 36077
rect 6903 35841 7139 36077
rect 7224 35841 7460 36077
rect 7545 35841 7781 36077
rect 7866 35841 8102 36077
rect 8187 35841 8423 36077
rect 8508 35841 8744 36077
rect 8829 35841 9065 36077
rect 9150 35841 9386 36077
rect 9471 35841 9707 36077
rect 9792 35841 10028 36077
rect 10113 35841 10349 36077
rect 10434 35841 10670 36077
rect 10755 35841 10991 36077
rect 11076 35841 11312 36077
rect 11397 35841 11633 36077
rect 11718 35841 11954 36077
rect 12038 35841 12274 36077
rect 12358 35841 12594 36077
rect 12678 35841 12914 36077
rect 12998 35841 13234 36077
rect 13318 35841 13554 36077
rect 13638 35841 13874 36077
rect 13958 35841 14194 36077
rect 14278 35841 14514 36077
rect 14598 35841 14834 36077
rect 14918 35841 15154 36077
rect 15238 35841 15474 36077
rect 15558 35841 15794 36077
rect 162 35517 398 35753
rect 483 35517 719 35753
rect 804 35517 1040 35753
rect 1125 35517 1361 35753
rect 1446 35517 1682 35753
rect 1767 35517 2003 35753
rect 2088 35517 2324 35753
rect 2409 35517 2645 35753
rect 2730 35517 2966 35753
rect 3051 35517 3287 35753
rect 3372 35517 3608 35753
rect 3693 35517 3929 35753
rect 4014 35517 4250 35753
rect 4335 35517 4571 35753
rect 4656 35517 4892 35753
rect 4977 35517 5213 35753
rect 5298 35517 5534 35753
rect 5619 35517 5855 35753
rect 5940 35517 6176 35753
rect 6261 35517 6497 35753
rect 6582 35517 6818 35753
rect 6903 35517 7139 35753
rect 7224 35517 7460 35753
rect 7545 35517 7781 35753
rect 7866 35517 8102 35753
rect 8187 35517 8423 35753
rect 8508 35517 8744 35753
rect 8829 35517 9065 35753
rect 9150 35517 9386 35753
rect 9471 35517 9707 35753
rect 9792 35517 10028 35753
rect 10113 35517 10349 35753
rect 10434 35517 10670 35753
rect 10755 35517 10991 35753
rect 11076 35517 11312 35753
rect 11397 35517 11633 35753
rect 11718 35517 11954 35753
rect 12038 35517 12274 35753
rect 12358 35517 12594 35753
rect 12678 35517 12914 35753
rect 12998 35517 13234 35753
rect 13318 35517 13554 35753
rect 13638 35517 13874 35753
rect 13958 35517 14194 35753
rect 14278 35517 14514 35753
rect 14598 35517 14834 35753
rect 14918 35517 15154 35753
rect 15238 35517 15474 35753
rect 15558 35517 15794 35753
rect 162 35193 398 35429
rect 483 35193 719 35429
rect 804 35193 1040 35429
rect 1125 35193 1361 35429
rect 1446 35193 1682 35429
rect 1767 35193 2003 35429
rect 2088 35193 2324 35429
rect 2409 35193 2645 35429
rect 2730 35193 2966 35429
rect 3051 35193 3287 35429
rect 3372 35193 3608 35429
rect 3693 35193 3929 35429
rect 4014 35193 4250 35429
rect 4335 35193 4571 35429
rect 4656 35193 4892 35429
rect 4977 35193 5213 35429
rect 5298 35193 5534 35429
rect 5619 35193 5855 35429
rect 5940 35193 6176 35429
rect 6261 35193 6497 35429
rect 6582 35193 6818 35429
rect 6903 35193 7139 35429
rect 7224 35193 7460 35429
rect 7545 35193 7781 35429
rect 7866 35193 8102 35429
rect 8187 35193 8423 35429
rect 8508 35193 8744 35429
rect 8829 35193 9065 35429
rect 9150 35193 9386 35429
rect 9471 35193 9707 35429
rect 9792 35193 10028 35429
rect 10113 35193 10349 35429
rect 10434 35193 10670 35429
rect 10755 35193 10991 35429
rect 11076 35193 11312 35429
rect 11397 35193 11633 35429
rect 11718 35193 11954 35429
rect 12038 35193 12274 35429
rect 12358 35193 12594 35429
rect 12678 35193 12914 35429
rect 12998 35193 13234 35429
rect 13318 35193 13554 35429
rect 13638 35193 13874 35429
rect 13958 35193 14194 35429
rect 14278 35193 14514 35429
rect 14598 35193 14834 35429
rect 14918 35193 15154 35429
rect 15238 35193 15474 35429
rect 15558 35193 15794 35429
rect 162 18736 398 18972
rect 483 18736 719 18972
rect 804 18736 1040 18972
rect 1125 18736 1361 18972
rect 1446 18736 1682 18972
rect 1767 18736 2003 18972
rect 2088 18736 2324 18972
rect 2409 18736 2645 18972
rect 2730 18736 2966 18972
rect 3051 18736 3287 18972
rect 3372 18736 3608 18972
rect 3693 18736 3929 18972
rect 4014 18736 4250 18972
rect 4335 18736 4571 18972
rect 4656 18736 4892 18972
rect 4977 18736 5213 18972
rect 5298 18736 5534 18972
rect 5619 18736 5855 18972
rect 5940 18736 6176 18972
rect 6261 18736 6497 18972
rect 6582 18736 6818 18972
rect 6903 18736 7139 18972
rect 7224 18736 7460 18972
rect 7545 18736 7781 18972
rect 7866 18736 8102 18972
rect 8187 18736 8423 18972
rect 8508 18736 8744 18972
rect 8829 18736 9065 18972
rect 9150 18736 9386 18972
rect 9471 18736 9707 18972
rect 9792 18736 10028 18972
rect 10113 18736 10349 18972
rect 10434 18736 10670 18972
rect 10755 18736 10991 18972
rect 11076 18736 11312 18972
rect 11397 18736 11633 18972
rect 11718 18736 11954 18972
rect 12038 18736 12274 18972
rect 12358 18736 12594 18972
rect 12678 18736 12914 18972
rect 12998 18736 13234 18972
rect 13318 18736 13554 18972
rect 13638 18736 13874 18972
rect 13958 18736 14194 18972
rect 14278 18736 14514 18972
rect 14598 18736 14834 18972
rect 14918 18736 15154 18972
rect 15238 18736 15474 18972
rect 15558 18736 15794 18972
rect 162 18400 398 18636
rect 483 18400 719 18636
rect 804 18400 1040 18636
rect 1125 18400 1361 18636
rect 1446 18400 1682 18636
rect 1767 18400 2003 18636
rect 2088 18400 2324 18636
rect 2409 18400 2645 18636
rect 2730 18400 2966 18636
rect 3051 18400 3287 18636
rect 3372 18400 3608 18636
rect 3693 18400 3929 18636
rect 4014 18400 4250 18636
rect 4335 18400 4571 18636
rect 4656 18400 4892 18636
rect 4977 18400 5213 18636
rect 5298 18400 5534 18636
rect 5619 18400 5855 18636
rect 5940 18400 6176 18636
rect 6261 18400 6497 18636
rect 6582 18400 6818 18636
rect 6903 18400 7139 18636
rect 7224 18400 7460 18636
rect 7545 18400 7781 18636
rect 7866 18400 8102 18636
rect 8187 18400 8423 18636
rect 8508 18400 8744 18636
rect 8829 18400 9065 18636
rect 9150 18400 9386 18636
rect 9471 18400 9707 18636
rect 9792 18400 10028 18636
rect 10113 18400 10349 18636
rect 10434 18400 10670 18636
rect 10755 18400 10991 18636
rect 11076 18400 11312 18636
rect 11397 18400 11633 18636
rect 11718 18400 11954 18636
rect 12038 18400 12274 18636
rect 12358 18400 12594 18636
rect 12678 18400 12914 18636
rect 12998 18400 13234 18636
rect 13318 18400 13554 18636
rect 13638 18400 13874 18636
rect 13958 18400 14194 18636
rect 14278 18400 14514 18636
rect 14598 18400 14834 18636
rect 14918 18400 15154 18636
rect 15238 18400 15474 18636
rect 15558 18400 15794 18636
rect 162 18064 398 18300
rect 483 18064 719 18300
rect 804 18064 1040 18300
rect 1125 18064 1361 18300
rect 1446 18064 1682 18300
rect 1767 18064 2003 18300
rect 2088 18064 2324 18300
rect 2409 18064 2645 18300
rect 2730 18064 2966 18300
rect 3051 18064 3287 18300
rect 3372 18064 3608 18300
rect 3693 18064 3929 18300
rect 4014 18064 4250 18300
rect 4335 18064 4571 18300
rect 4656 18064 4892 18300
rect 4977 18064 5213 18300
rect 5298 18064 5534 18300
rect 5619 18064 5855 18300
rect 5940 18064 6176 18300
rect 6261 18064 6497 18300
rect 6582 18064 6818 18300
rect 6903 18064 7139 18300
rect 7224 18064 7460 18300
rect 7545 18064 7781 18300
rect 7866 18064 8102 18300
rect 8187 18064 8423 18300
rect 8508 18064 8744 18300
rect 8829 18064 9065 18300
rect 9150 18064 9386 18300
rect 9471 18064 9707 18300
rect 9792 18064 10028 18300
rect 10113 18064 10349 18300
rect 10434 18064 10670 18300
rect 10755 18064 10991 18300
rect 11076 18064 11312 18300
rect 11397 18064 11633 18300
rect 11718 18064 11954 18300
rect 12038 18064 12274 18300
rect 12358 18064 12594 18300
rect 12678 18064 12914 18300
rect 12998 18064 13234 18300
rect 13318 18064 13554 18300
rect 13638 18064 13874 18300
rect 13958 18064 14194 18300
rect 14278 18064 14514 18300
rect 14598 18064 14834 18300
rect 14918 18064 15154 18300
rect 15238 18064 15474 18300
rect 15558 18064 15794 18300
rect 162 17728 398 17964
rect 483 17728 719 17964
rect 804 17728 1040 17964
rect 1125 17728 1361 17964
rect 1446 17728 1682 17964
rect 1767 17728 2003 17964
rect 2088 17728 2324 17964
rect 2409 17728 2645 17964
rect 2730 17728 2966 17964
rect 3051 17728 3287 17964
rect 3372 17728 3608 17964
rect 3693 17728 3929 17964
rect 4014 17728 4250 17964
rect 4335 17728 4571 17964
rect 4656 17728 4892 17964
rect 4977 17728 5213 17964
rect 5298 17728 5534 17964
rect 5619 17728 5855 17964
rect 5940 17728 6176 17964
rect 6261 17728 6497 17964
rect 6582 17728 6818 17964
rect 6903 17728 7139 17964
rect 7224 17728 7460 17964
rect 7545 17728 7781 17964
rect 7866 17728 8102 17964
rect 8187 17728 8423 17964
rect 8508 17728 8744 17964
rect 8829 17728 9065 17964
rect 9150 17728 9386 17964
rect 9471 17728 9707 17964
rect 9792 17728 10028 17964
rect 10113 17728 10349 17964
rect 10434 17728 10670 17964
rect 10755 17728 10991 17964
rect 11076 17728 11312 17964
rect 11397 17728 11633 17964
rect 11718 17728 11954 17964
rect 12038 17728 12274 17964
rect 12358 17728 12594 17964
rect 12678 17728 12914 17964
rect 12998 17728 13234 17964
rect 13318 17728 13554 17964
rect 13638 17728 13874 17964
rect 13958 17728 14194 17964
rect 14278 17728 14514 17964
rect 14598 17728 14834 17964
rect 14918 17728 15154 17964
rect 15238 17728 15474 17964
rect 15558 17728 15794 17964
rect 162 17392 398 17628
rect 483 17392 719 17628
rect 804 17392 1040 17628
rect 1125 17392 1361 17628
rect 1446 17392 1682 17628
rect 1767 17392 2003 17628
rect 2088 17392 2324 17628
rect 2409 17392 2645 17628
rect 2730 17392 2966 17628
rect 3051 17392 3287 17628
rect 3372 17392 3608 17628
rect 3693 17392 3929 17628
rect 4014 17392 4250 17628
rect 4335 17392 4571 17628
rect 4656 17392 4892 17628
rect 4977 17392 5213 17628
rect 5298 17392 5534 17628
rect 5619 17392 5855 17628
rect 5940 17392 6176 17628
rect 6261 17392 6497 17628
rect 6582 17392 6818 17628
rect 6903 17392 7139 17628
rect 7224 17392 7460 17628
rect 7545 17392 7781 17628
rect 7866 17392 8102 17628
rect 8187 17392 8423 17628
rect 8508 17392 8744 17628
rect 8829 17392 9065 17628
rect 9150 17392 9386 17628
rect 9471 17392 9707 17628
rect 9792 17392 10028 17628
rect 10113 17392 10349 17628
rect 10434 17392 10670 17628
rect 10755 17392 10991 17628
rect 11076 17392 11312 17628
rect 11397 17392 11633 17628
rect 11718 17392 11954 17628
rect 12038 17392 12274 17628
rect 12358 17392 12594 17628
rect 12678 17392 12914 17628
rect 12998 17392 13234 17628
rect 13318 17392 13554 17628
rect 13638 17392 13874 17628
rect 13958 17392 14194 17628
rect 14278 17392 14514 17628
rect 14598 17392 14834 17628
rect 14918 17392 15154 17628
rect 15238 17392 15474 17628
rect 15558 17392 15794 17628
rect 162 17056 398 17292
rect 483 17056 719 17292
rect 804 17056 1040 17292
rect 1125 17056 1361 17292
rect 1446 17056 1682 17292
rect 1767 17056 2003 17292
rect 2088 17056 2324 17292
rect 2409 17056 2645 17292
rect 2730 17056 2966 17292
rect 3051 17056 3287 17292
rect 3372 17056 3608 17292
rect 3693 17056 3929 17292
rect 4014 17056 4250 17292
rect 4335 17056 4571 17292
rect 4656 17056 4892 17292
rect 4977 17056 5213 17292
rect 5298 17056 5534 17292
rect 5619 17056 5855 17292
rect 5940 17056 6176 17292
rect 6261 17056 6497 17292
rect 6582 17056 6818 17292
rect 6903 17056 7139 17292
rect 7224 17056 7460 17292
rect 7545 17056 7781 17292
rect 7866 17056 8102 17292
rect 8187 17056 8423 17292
rect 8508 17056 8744 17292
rect 8829 17056 9065 17292
rect 9150 17056 9386 17292
rect 9471 17056 9707 17292
rect 9792 17056 10028 17292
rect 10113 17056 10349 17292
rect 10434 17056 10670 17292
rect 10755 17056 10991 17292
rect 11076 17056 11312 17292
rect 11397 17056 11633 17292
rect 11718 17056 11954 17292
rect 12038 17056 12274 17292
rect 12358 17056 12594 17292
rect 12678 17056 12914 17292
rect 12998 17056 13234 17292
rect 13318 17056 13554 17292
rect 13638 17056 13874 17292
rect 13958 17056 14194 17292
rect 14278 17056 14514 17292
rect 14598 17056 14834 17292
rect 14918 17056 15154 17292
rect 15238 17056 15474 17292
rect 15558 17056 15794 17292
rect 162 16720 398 16956
rect 483 16720 719 16956
rect 804 16720 1040 16956
rect 1125 16720 1361 16956
rect 1446 16720 1682 16956
rect 1767 16720 2003 16956
rect 2088 16720 2324 16956
rect 2409 16720 2645 16956
rect 2730 16720 2966 16956
rect 3051 16720 3287 16956
rect 3372 16720 3608 16956
rect 3693 16720 3929 16956
rect 4014 16720 4250 16956
rect 4335 16720 4571 16956
rect 4656 16720 4892 16956
rect 4977 16720 5213 16956
rect 5298 16720 5534 16956
rect 5619 16720 5855 16956
rect 5940 16720 6176 16956
rect 6261 16720 6497 16956
rect 6582 16720 6818 16956
rect 6903 16720 7139 16956
rect 7224 16720 7460 16956
rect 7545 16720 7781 16956
rect 7866 16720 8102 16956
rect 8187 16720 8423 16956
rect 8508 16720 8744 16956
rect 8829 16720 9065 16956
rect 9150 16720 9386 16956
rect 9471 16720 9707 16956
rect 9792 16720 10028 16956
rect 10113 16720 10349 16956
rect 10434 16720 10670 16956
rect 10755 16720 10991 16956
rect 11076 16720 11312 16956
rect 11397 16720 11633 16956
rect 11718 16720 11954 16956
rect 12038 16720 12274 16956
rect 12358 16720 12594 16956
rect 12678 16720 12914 16956
rect 12998 16720 13234 16956
rect 13318 16720 13554 16956
rect 13638 16720 13874 16956
rect 13958 16720 14194 16956
rect 14278 16720 14514 16956
rect 14598 16720 14834 16956
rect 14918 16720 15154 16956
rect 15238 16720 15474 16956
rect 15558 16720 15794 16956
rect 162 16384 398 16620
rect 483 16384 719 16620
rect 804 16384 1040 16620
rect 1125 16384 1361 16620
rect 1446 16384 1682 16620
rect 1767 16384 2003 16620
rect 2088 16384 2324 16620
rect 2409 16384 2645 16620
rect 2730 16384 2966 16620
rect 3051 16384 3287 16620
rect 3372 16384 3608 16620
rect 3693 16384 3929 16620
rect 4014 16384 4250 16620
rect 4335 16384 4571 16620
rect 4656 16384 4892 16620
rect 4977 16384 5213 16620
rect 5298 16384 5534 16620
rect 5619 16384 5855 16620
rect 5940 16384 6176 16620
rect 6261 16384 6497 16620
rect 6582 16384 6818 16620
rect 6903 16384 7139 16620
rect 7224 16384 7460 16620
rect 7545 16384 7781 16620
rect 7866 16384 8102 16620
rect 8187 16384 8423 16620
rect 8508 16384 8744 16620
rect 8829 16384 9065 16620
rect 9150 16384 9386 16620
rect 9471 16384 9707 16620
rect 9792 16384 10028 16620
rect 10113 16384 10349 16620
rect 10434 16384 10670 16620
rect 10755 16384 10991 16620
rect 11076 16384 11312 16620
rect 11397 16384 11633 16620
rect 11718 16384 11954 16620
rect 12038 16384 12274 16620
rect 12358 16384 12594 16620
rect 12678 16384 12914 16620
rect 12998 16384 13234 16620
rect 13318 16384 13554 16620
rect 13638 16384 13874 16620
rect 13958 16384 14194 16620
rect 14278 16384 14514 16620
rect 14598 16384 14834 16620
rect 14918 16384 15154 16620
rect 15238 16384 15474 16620
rect 15558 16384 15794 16620
rect 162 16048 398 16284
rect 483 16048 719 16284
rect 804 16048 1040 16284
rect 1125 16048 1361 16284
rect 1446 16048 1682 16284
rect 1767 16048 2003 16284
rect 2088 16048 2324 16284
rect 2409 16048 2645 16284
rect 2730 16048 2966 16284
rect 3051 16048 3287 16284
rect 3372 16048 3608 16284
rect 3693 16048 3929 16284
rect 4014 16048 4250 16284
rect 4335 16048 4571 16284
rect 4656 16048 4892 16284
rect 4977 16048 5213 16284
rect 5298 16048 5534 16284
rect 5619 16048 5855 16284
rect 5940 16048 6176 16284
rect 6261 16048 6497 16284
rect 6582 16048 6818 16284
rect 6903 16048 7139 16284
rect 7224 16048 7460 16284
rect 7545 16048 7781 16284
rect 7866 16048 8102 16284
rect 8187 16048 8423 16284
rect 8508 16048 8744 16284
rect 8829 16048 9065 16284
rect 9150 16048 9386 16284
rect 9471 16048 9707 16284
rect 9792 16048 10028 16284
rect 10113 16048 10349 16284
rect 10434 16048 10670 16284
rect 10755 16048 10991 16284
rect 11076 16048 11312 16284
rect 11397 16048 11633 16284
rect 11718 16048 11954 16284
rect 12038 16048 12274 16284
rect 12358 16048 12594 16284
rect 12678 16048 12914 16284
rect 12998 16048 13234 16284
rect 13318 16048 13554 16284
rect 13638 16048 13874 16284
rect 13958 16048 14194 16284
rect 14278 16048 14514 16284
rect 14598 16048 14834 16284
rect 14918 16048 15154 16284
rect 15238 16048 15474 16284
rect 15558 16048 15794 16284
rect 162 15712 398 15948
rect 483 15712 719 15948
rect 804 15712 1040 15948
rect 1125 15712 1361 15948
rect 1446 15712 1682 15948
rect 1767 15712 2003 15948
rect 2088 15712 2324 15948
rect 2409 15712 2645 15948
rect 2730 15712 2966 15948
rect 3051 15712 3287 15948
rect 3372 15712 3608 15948
rect 3693 15712 3929 15948
rect 4014 15712 4250 15948
rect 4335 15712 4571 15948
rect 4656 15712 4892 15948
rect 4977 15712 5213 15948
rect 5298 15712 5534 15948
rect 5619 15712 5855 15948
rect 5940 15712 6176 15948
rect 6261 15712 6497 15948
rect 6582 15712 6818 15948
rect 6903 15712 7139 15948
rect 7224 15712 7460 15948
rect 7545 15712 7781 15948
rect 7866 15712 8102 15948
rect 8187 15712 8423 15948
rect 8508 15712 8744 15948
rect 8829 15712 9065 15948
rect 9150 15712 9386 15948
rect 9471 15712 9707 15948
rect 9792 15712 10028 15948
rect 10113 15712 10349 15948
rect 10434 15712 10670 15948
rect 10755 15712 10991 15948
rect 11076 15712 11312 15948
rect 11397 15712 11633 15948
rect 11718 15712 11954 15948
rect 12038 15712 12274 15948
rect 12358 15712 12594 15948
rect 12678 15712 12914 15948
rect 12998 15712 13234 15948
rect 13318 15712 13554 15948
rect 13638 15712 13874 15948
rect 13958 15712 14194 15948
rect 14278 15712 14514 15948
rect 14598 15712 14834 15948
rect 14918 15712 15154 15948
rect 15238 15712 15474 15948
rect 15558 15712 15794 15948
rect 162 15376 398 15612
rect 483 15376 719 15612
rect 804 15376 1040 15612
rect 1125 15376 1361 15612
rect 1446 15376 1682 15612
rect 1767 15376 2003 15612
rect 2088 15376 2324 15612
rect 2409 15376 2645 15612
rect 2730 15376 2966 15612
rect 3051 15376 3287 15612
rect 3372 15376 3608 15612
rect 3693 15376 3929 15612
rect 4014 15376 4250 15612
rect 4335 15376 4571 15612
rect 4656 15376 4892 15612
rect 4977 15376 5213 15612
rect 5298 15376 5534 15612
rect 5619 15376 5855 15612
rect 5940 15376 6176 15612
rect 6261 15376 6497 15612
rect 6582 15376 6818 15612
rect 6903 15376 7139 15612
rect 7224 15376 7460 15612
rect 7545 15376 7781 15612
rect 7866 15376 8102 15612
rect 8187 15376 8423 15612
rect 8508 15376 8744 15612
rect 8829 15376 9065 15612
rect 9150 15376 9386 15612
rect 9471 15376 9707 15612
rect 9792 15376 10028 15612
rect 10113 15376 10349 15612
rect 10434 15376 10670 15612
rect 10755 15376 10991 15612
rect 11076 15376 11312 15612
rect 11397 15376 11633 15612
rect 11718 15376 11954 15612
rect 12038 15376 12274 15612
rect 12358 15376 12594 15612
rect 12678 15376 12914 15612
rect 12998 15376 13234 15612
rect 13318 15376 13554 15612
rect 13638 15376 13874 15612
rect 13958 15376 14194 15612
rect 14278 15376 14514 15612
rect 14598 15376 14834 15612
rect 14918 15376 15154 15612
rect 15238 15376 15474 15612
rect 15558 15376 15794 15612
rect 162 15040 398 15276
rect 483 15040 719 15276
rect 804 15040 1040 15276
rect 1125 15040 1361 15276
rect 1446 15040 1682 15276
rect 1767 15040 2003 15276
rect 2088 15040 2324 15276
rect 2409 15040 2645 15276
rect 2730 15040 2966 15276
rect 3051 15040 3287 15276
rect 3372 15040 3608 15276
rect 3693 15040 3929 15276
rect 4014 15040 4250 15276
rect 4335 15040 4571 15276
rect 4656 15040 4892 15276
rect 4977 15040 5213 15276
rect 5298 15040 5534 15276
rect 5619 15040 5855 15276
rect 5940 15040 6176 15276
rect 6261 15040 6497 15276
rect 6582 15040 6818 15276
rect 6903 15040 7139 15276
rect 7224 15040 7460 15276
rect 7545 15040 7781 15276
rect 7866 15040 8102 15276
rect 8187 15040 8423 15276
rect 8508 15040 8744 15276
rect 8829 15040 9065 15276
rect 9150 15040 9386 15276
rect 9471 15040 9707 15276
rect 9792 15040 10028 15276
rect 10113 15040 10349 15276
rect 10434 15040 10670 15276
rect 10755 15040 10991 15276
rect 11076 15040 11312 15276
rect 11397 15040 11633 15276
rect 11718 15040 11954 15276
rect 12038 15040 12274 15276
rect 12358 15040 12594 15276
rect 12678 15040 12914 15276
rect 12998 15040 13234 15276
rect 13318 15040 13554 15276
rect 13638 15040 13874 15276
rect 13958 15040 14194 15276
rect 14278 15040 14514 15276
rect 14598 15040 14834 15276
rect 14918 15040 15154 15276
rect 15238 15040 15474 15276
rect 15558 15040 15794 15276
rect 162 14704 398 14940
rect 483 14704 719 14940
rect 804 14704 1040 14940
rect 1125 14704 1361 14940
rect 1446 14704 1682 14940
rect 1767 14704 2003 14940
rect 2088 14704 2324 14940
rect 2409 14704 2645 14940
rect 2730 14704 2966 14940
rect 3051 14704 3287 14940
rect 3372 14704 3608 14940
rect 3693 14704 3929 14940
rect 4014 14704 4250 14940
rect 4335 14704 4571 14940
rect 4656 14704 4892 14940
rect 4977 14704 5213 14940
rect 5298 14704 5534 14940
rect 5619 14704 5855 14940
rect 5940 14704 6176 14940
rect 6261 14704 6497 14940
rect 6582 14704 6818 14940
rect 6903 14704 7139 14940
rect 7224 14704 7460 14940
rect 7545 14704 7781 14940
rect 7866 14704 8102 14940
rect 8187 14704 8423 14940
rect 8508 14704 8744 14940
rect 8829 14704 9065 14940
rect 9150 14704 9386 14940
rect 9471 14704 9707 14940
rect 9792 14704 10028 14940
rect 10113 14704 10349 14940
rect 10434 14704 10670 14940
rect 10755 14704 10991 14940
rect 11076 14704 11312 14940
rect 11397 14704 11633 14940
rect 11718 14704 11954 14940
rect 12038 14704 12274 14940
rect 12358 14704 12594 14940
rect 12678 14704 12914 14940
rect 12998 14704 13234 14940
rect 13318 14704 13554 14940
rect 13638 14704 13874 14940
rect 13958 14704 14194 14940
rect 14278 14704 14514 14940
rect 14598 14704 14834 14940
rect 14918 14704 15154 14940
rect 15238 14704 15474 14940
rect 15558 14704 15794 14940
rect 162 14368 398 14604
rect 483 14368 719 14604
rect 804 14368 1040 14604
rect 1125 14368 1361 14604
rect 1446 14368 1682 14604
rect 1767 14368 2003 14604
rect 2088 14368 2324 14604
rect 2409 14368 2645 14604
rect 2730 14368 2966 14604
rect 3051 14368 3287 14604
rect 3372 14368 3608 14604
rect 3693 14368 3929 14604
rect 4014 14368 4250 14604
rect 4335 14368 4571 14604
rect 4656 14368 4892 14604
rect 4977 14368 5213 14604
rect 5298 14368 5534 14604
rect 5619 14368 5855 14604
rect 5940 14368 6176 14604
rect 6261 14368 6497 14604
rect 6582 14368 6818 14604
rect 6903 14368 7139 14604
rect 7224 14368 7460 14604
rect 7545 14368 7781 14604
rect 7866 14368 8102 14604
rect 8187 14368 8423 14604
rect 8508 14368 8744 14604
rect 8829 14368 9065 14604
rect 9150 14368 9386 14604
rect 9471 14368 9707 14604
rect 9792 14368 10028 14604
rect 10113 14368 10349 14604
rect 10434 14368 10670 14604
rect 10755 14368 10991 14604
rect 11076 14368 11312 14604
rect 11397 14368 11633 14604
rect 11718 14368 11954 14604
rect 12038 14368 12274 14604
rect 12358 14368 12594 14604
rect 12678 14368 12914 14604
rect 12998 14368 13234 14604
rect 13318 14368 13554 14604
rect 13638 14368 13874 14604
rect 13958 14368 14194 14604
rect 14278 14368 14514 14604
rect 14598 14368 14834 14604
rect 14918 14368 15154 14604
rect 15238 14368 15474 14604
rect 15558 14368 15794 14604
rect 162 14032 398 14268
rect 483 14032 719 14268
rect 804 14032 1040 14268
rect 1125 14032 1361 14268
rect 1446 14032 1682 14268
rect 1767 14032 2003 14268
rect 2088 14032 2324 14268
rect 2409 14032 2645 14268
rect 2730 14032 2966 14268
rect 3051 14032 3287 14268
rect 3372 14032 3608 14268
rect 3693 14032 3929 14268
rect 4014 14032 4250 14268
rect 4335 14032 4571 14268
rect 4656 14032 4892 14268
rect 4977 14032 5213 14268
rect 5298 14032 5534 14268
rect 5619 14032 5855 14268
rect 5940 14032 6176 14268
rect 6261 14032 6497 14268
rect 6582 14032 6818 14268
rect 6903 14032 7139 14268
rect 7224 14032 7460 14268
rect 7545 14032 7781 14268
rect 7866 14032 8102 14268
rect 8187 14032 8423 14268
rect 8508 14032 8744 14268
rect 8829 14032 9065 14268
rect 9150 14032 9386 14268
rect 9471 14032 9707 14268
rect 9792 14032 10028 14268
rect 10113 14032 10349 14268
rect 10434 14032 10670 14268
rect 10755 14032 10991 14268
rect 11076 14032 11312 14268
rect 11397 14032 11633 14268
rect 11718 14032 11954 14268
rect 12038 14032 12274 14268
rect 12358 14032 12594 14268
rect 12678 14032 12914 14268
rect 12998 14032 13234 14268
rect 13318 14032 13554 14268
rect 13638 14032 13874 14268
rect 13958 14032 14194 14268
rect 14278 14032 14514 14268
rect 14598 14032 14834 14268
rect 14918 14032 15154 14268
rect 15238 14032 15474 14268
rect 15558 14032 15794 14268
rect 162 13427 398 13663
rect 483 13427 719 13663
rect 804 13427 1040 13663
rect 1125 13427 1361 13663
rect 1446 13427 1682 13663
rect 1767 13427 2003 13663
rect 2088 13427 2324 13663
rect 2409 13427 2645 13663
rect 2730 13427 2966 13663
rect 3051 13427 3287 13663
rect 3372 13427 3608 13663
rect 3693 13427 3929 13663
rect 4014 13427 4250 13663
rect 4335 13427 4571 13663
rect 4656 13427 4892 13663
rect 4977 13427 5213 13663
rect 5298 13427 5534 13663
rect 5619 13427 5855 13663
rect 5940 13427 6176 13663
rect 6261 13427 6497 13663
rect 6582 13427 6818 13663
rect 6903 13427 7139 13663
rect 7224 13427 7460 13663
rect 7545 13427 7781 13663
rect 7866 13427 8102 13663
rect 8187 13427 8423 13663
rect 8508 13427 8744 13663
rect 8829 13427 9065 13663
rect 9150 13427 9386 13663
rect 9471 13427 9707 13663
rect 9792 13427 10028 13663
rect 10113 13427 10349 13663
rect 10434 13427 10670 13663
rect 10755 13427 10991 13663
rect 11076 13427 11312 13663
rect 11397 13427 11633 13663
rect 11718 13427 11954 13663
rect 12038 13427 12274 13663
rect 12358 13427 12594 13663
rect 12678 13427 12914 13663
rect 12998 13427 13234 13663
rect 13318 13427 13554 13663
rect 13638 13427 13874 13663
rect 13958 13427 14194 13663
rect 14278 13427 14514 13663
rect 14598 13427 14834 13663
rect 14918 13427 15154 13663
rect 15238 13427 15474 13663
rect 15558 13427 15794 13663
rect 162 12861 398 13097
rect 483 12861 719 13097
rect 804 12861 1040 13097
rect 1125 12861 1361 13097
rect 1446 12861 1682 13097
rect 1767 12861 2003 13097
rect 2088 12861 2324 13097
rect 2409 12861 2645 13097
rect 2730 12861 2966 13097
rect 3051 12861 3287 13097
rect 3372 12861 3608 13097
rect 3693 12861 3929 13097
rect 4014 12861 4250 13097
rect 4335 12861 4571 13097
rect 4656 12861 4892 13097
rect 4977 12861 5213 13097
rect 5298 12861 5534 13097
rect 5619 12861 5855 13097
rect 5940 12861 6176 13097
rect 6261 12861 6497 13097
rect 6582 12861 6818 13097
rect 6903 12861 7139 13097
rect 7224 12861 7460 13097
rect 7545 12861 7781 13097
rect 7866 12861 8102 13097
rect 8187 12861 8423 13097
rect 8508 12861 8744 13097
rect 8829 12861 9065 13097
rect 9150 12861 9386 13097
rect 9471 12861 9707 13097
rect 9792 12861 10028 13097
rect 10113 12861 10349 13097
rect 10434 12861 10670 13097
rect 10755 12861 10991 13097
rect 11076 12861 11312 13097
rect 11397 12861 11633 13097
rect 11718 12861 11954 13097
rect 12038 12861 12274 13097
rect 12358 12861 12594 13097
rect 12678 12861 12914 13097
rect 12998 12861 13234 13097
rect 13318 12861 13554 13097
rect 13638 12861 13874 13097
rect 13958 12861 14194 13097
rect 14278 12861 14514 13097
rect 14598 12861 14834 13097
rect 14918 12861 15154 13097
rect 15238 12861 15474 13097
rect 15558 12861 15794 13097
rect 162 12257 398 12493
rect 483 12257 719 12493
rect 804 12257 1040 12493
rect 1125 12257 1361 12493
rect 1446 12257 1682 12493
rect 1767 12257 2003 12493
rect 2088 12257 2324 12493
rect 2409 12257 2645 12493
rect 2730 12257 2966 12493
rect 3051 12257 3287 12493
rect 3372 12257 3608 12493
rect 3693 12257 3929 12493
rect 4014 12257 4250 12493
rect 4335 12257 4571 12493
rect 4656 12257 4892 12493
rect 4977 12257 5213 12493
rect 5298 12257 5534 12493
rect 5619 12257 5855 12493
rect 5940 12257 6176 12493
rect 6261 12257 6497 12493
rect 6582 12257 6818 12493
rect 6903 12257 7139 12493
rect 7224 12257 7460 12493
rect 7545 12257 7781 12493
rect 7866 12257 8102 12493
rect 8187 12257 8423 12493
rect 8508 12257 8744 12493
rect 8829 12257 9065 12493
rect 9150 12257 9386 12493
rect 9471 12257 9707 12493
rect 9792 12257 10028 12493
rect 10113 12257 10349 12493
rect 10434 12257 10670 12493
rect 10755 12257 10991 12493
rect 11076 12257 11312 12493
rect 11397 12257 11633 12493
rect 11718 12257 11954 12493
rect 12039 12257 12275 12493
rect 12359 12257 12595 12493
rect 12679 12257 12915 12493
rect 12999 12257 13235 12493
rect 13319 12257 13555 12493
rect 13639 12257 13875 12493
rect 13959 12257 14195 12493
rect 14279 12257 14515 12493
rect 14599 12257 14835 12493
rect 14919 12257 15155 12493
rect 15239 12257 15475 12493
rect 15559 12257 15795 12493
rect 162 11691 398 11927
rect 483 11691 719 11927
rect 804 11691 1040 11927
rect 1125 11691 1361 11927
rect 1446 11691 1682 11927
rect 1767 11691 2003 11927
rect 2088 11691 2324 11927
rect 2409 11691 2645 11927
rect 2730 11691 2966 11927
rect 3051 11691 3287 11927
rect 3372 11691 3608 11927
rect 3693 11691 3929 11927
rect 4014 11691 4250 11927
rect 4335 11691 4571 11927
rect 4656 11691 4892 11927
rect 4977 11691 5213 11927
rect 5298 11691 5534 11927
rect 5619 11691 5855 11927
rect 5940 11691 6176 11927
rect 6261 11691 6497 11927
rect 6582 11691 6818 11927
rect 6903 11691 7139 11927
rect 7224 11691 7460 11927
rect 7545 11691 7781 11927
rect 7866 11691 8102 11927
rect 8187 11691 8423 11927
rect 8508 11691 8744 11927
rect 8829 11691 9065 11927
rect 9150 11691 9386 11927
rect 9471 11691 9707 11927
rect 9792 11691 10028 11927
rect 10113 11691 10349 11927
rect 10434 11691 10670 11927
rect 10755 11691 10991 11927
rect 11076 11691 11312 11927
rect 11397 11691 11633 11927
rect 11718 11691 11954 11927
rect 12039 11691 12275 11927
rect 12359 11691 12595 11927
rect 12679 11691 12915 11927
rect 12999 11691 13235 11927
rect 13319 11691 13555 11927
rect 13639 11691 13875 11927
rect 13959 11691 14195 11927
rect 14279 11691 14515 11927
rect 14599 11691 14835 11927
rect 14919 11691 15155 11927
rect 15239 11691 15475 11927
rect 15559 11691 15795 11927
rect 162 10329 398 10565
rect 483 10329 719 10565
rect 804 10329 1040 10565
rect 1125 10329 1361 10565
rect 1446 10329 1682 10565
rect 1767 10329 2003 10565
rect 2088 10329 2324 10565
rect 2409 10329 2645 10565
rect 2730 10329 2966 10565
rect 3051 10329 3287 10565
rect 3372 10329 3608 10565
rect 3693 10329 3929 10565
rect 4014 10329 4250 10565
rect 4335 10329 4571 10565
rect 4656 10329 4892 10565
rect 4977 10329 5213 10565
rect 5298 10329 5534 10565
rect 5619 10329 5855 10565
rect 5940 10329 6176 10565
rect 6261 10329 6497 10565
rect 6582 10329 6818 10565
rect 6903 10329 7139 10565
rect 7224 10329 7460 10565
rect 7545 10329 7781 10565
rect 7866 10329 8102 10565
rect 8187 10329 8423 10565
rect 8508 10329 8744 10565
rect 8829 10329 9065 10565
rect 9150 10329 9386 10565
rect 9471 10329 9707 10565
rect 9792 10329 10028 10565
rect 10113 10329 10349 10565
rect 10434 10329 10670 10565
rect 10755 10329 10991 10565
rect 11076 10329 11312 10565
rect 11397 10329 11633 10565
rect 11718 10329 11954 10565
rect 12038 10329 12274 10565
rect 12358 10329 12594 10565
rect 12678 10329 12914 10565
rect 12998 10329 13234 10565
rect 13318 10329 13554 10565
rect 13638 10329 13874 10565
rect 13958 10329 14194 10565
rect 14278 10329 14514 10565
rect 14598 10329 14834 10565
rect 14918 10329 15154 10565
rect 15238 10329 15474 10565
rect 15558 10329 15794 10565
rect 162 8967 398 9203
rect 483 8967 719 9203
rect 804 8967 1040 9203
rect 1125 8967 1361 9203
rect 1446 8967 1682 9203
rect 1767 8967 2003 9203
rect 2088 8967 2324 9203
rect 2409 8967 2645 9203
rect 2730 8967 2966 9203
rect 3051 8967 3287 9203
rect 3372 8967 3608 9203
rect 3693 8967 3929 9203
rect 4014 8967 4250 9203
rect 4335 8967 4571 9203
rect 4656 8967 4892 9203
rect 4977 8967 5213 9203
rect 5298 8967 5534 9203
rect 5619 8967 5855 9203
rect 5940 8967 6176 9203
rect 6261 8967 6497 9203
rect 6582 8967 6818 9203
rect 6903 8967 7139 9203
rect 7224 8967 7460 9203
rect 7545 8967 7781 9203
rect 7866 8967 8102 9203
rect 8187 8967 8423 9203
rect 8508 8967 8744 9203
rect 8829 8967 9065 9203
rect 9150 8967 9386 9203
rect 9471 8967 9707 9203
rect 9792 8967 10028 9203
rect 10113 8967 10349 9203
rect 10434 8967 10670 9203
rect 10755 8967 10991 9203
rect 11076 8967 11312 9203
rect 11397 8967 11633 9203
rect 11717 8967 11953 9203
rect 12037 8967 12273 9203
rect 12357 8967 12593 9203
rect 12677 8967 12913 9203
rect 12997 8967 13233 9203
rect 13317 8967 13553 9203
rect 13637 8967 13873 9203
rect 13957 8967 14193 9203
rect 14277 8967 14513 9203
rect 14597 8967 14833 9203
rect 14917 8967 15153 9203
rect 15237 8967 15473 9203
rect 15557 8967 15793 9203
rect 162 8361 398 8597
rect 483 8361 719 8597
rect 804 8361 1040 8597
rect 1125 8361 1361 8597
rect 1446 8361 1682 8597
rect 1767 8361 2003 8597
rect 2088 8361 2324 8597
rect 2409 8361 2645 8597
rect 2730 8361 2966 8597
rect 3051 8361 3287 8597
rect 3372 8361 3608 8597
rect 3693 8361 3929 8597
rect 4014 8361 4250 8597
rect 4335 8361 4571 8597
rect 4656 8361 4892 8597
rect 4977 8361 5213 8597
rect 5298 8361 5534 8597
rect 5619 8361 5855 8597
rect 5940 8361 6176 8597
rect 6261 8361 6497 8597
rect 6582 8361 6818 8597
rect 6903 8361 7139 8597
rect 7224 8361 7460 8597
rect 7545 8361 7781 8597
rect 7866 8361 8102 8597
rect 8187 8361 8423 8597
rect 8508 8361 8744 8597
rect 8829 8361 9065 8597
rect 9150 8361 9386 8597
rect 9471 8361 9707 8597
rect 9792 8361 10028 8597
rect 10113 8361 10349 8597
rect 10434 8361 10670 8597
rect 10755 8361 10991 8597
rect 11076 8361 11312 8597
rect 11397 8361 11633 8597
rect 11717 8361 11953 8597
rect 12037 8361 12273 8597
rect 12357 8361 12593 8597
rect 12677 8361 12913 8597
rect 12997 8361 13233 8597
rect 13317 8361 13553 8597
rect 13637 8361 13873 8597
rect 13957 8361 14193 8597
rect 14277 8361 14513 8597
rect 14597 8361 14833 8597
rect 14917 8361 15153 8597
rect 15237 8361 15473 8597
rect 15557 8361 15793 8597
rect 162 7757 398 7993
rect 483 7757 719 7993
rect 804 7757 1040 7993
rect 1125 7757 1361 7993
rect 1446 7757 1682 7993
rect 1767 7757 2003 7993
rect 2088 7757 2324 7993
rect 2409 7757 2645 7993
rect 2730 7757 2966 7993
rect 3051 7757 3287 7993
rect 3372 7757 3608 7993
rect 3693 7757 3929 7993
rect 4014 7757 4250 7993
rect 4335 7757 4571 7993
rect 4656 7757 4892 7993
rect 4977 7757 5213 7993
rect 5298 7757 5534 7993
rect 5619 7757 5855 7993
rect 5940 7757 6176 7993
rect 6261 7757 6497 7993
rect 6582 7757 6818 7993
rect 6903 7757 7139 7993
rect 7224 7757 7460 7993
rect 7545 7757 7781 7993
rect 7866 7757 8102 7993
rect 8187 7757 8423 7993
rect 8508 7757 8744 7993
rect 8829 7757 9065 7993
rect 9150 7757 9386 7993
rect 9471 7757 9707 7993
rect 9792 7757 10028 7993
rect 10113 7757 10349 7993
rect 10434 7757 10670 7993
rect 10755 7757 10991 7993
rect 11076 7757 11312 7993
rect 11397 7757 11633 7993
rect 11718 7757 11954 7993
rect 12039 7757 12275 7993
rect 12359 7757 12595 7993
rect 12679 7757 12915 7993
rect 12999 7757 13235 7993
rect 13319 7757 13555 7993
rect 13639 7757 13875 7993
rect 13959 7757 14195 7993
rect 14279 7757 14515 7993
rect 14599 7757 14835 7993
rect 14919 7757 15155 7993
rect 15239 7757 15475 7993
rect 15559 7757 15795 7993
rect 162 7391 398 7627
rect 483 7391 719 7627
rect 804 7391 1040 7627
rect 1125 7391 1361 7627
rect 1446 7391 1682 7627
rect 1767 7391 2003 7627
rect 2088 7391 2324 7627
rect 2409 7391 2645 7627
rect 2730 7391 2966 7627
rect 3051 7391 3287 7627
rect 3372 7391 3608 7627
rect 3693 7391 3929 7627
rect 4014 7391 4250 7627
rect 4335 7391 4571 7627
rect 4656 7391 4892 7627
rect 4977 7391 5213 7627
rect 5298 7391 5534 7627
rect 5619 7391 5855 7627
rect 5940 7391 6176 7627
rect 6261 7391 6497 7627
rect 6582 7391 6818 7627
rect 6903 7391 7139 7627
rect 7224 7391 7460 7627
rect 7545 7391 7781 7627
rect 7866 7391 8102 7627
rect 8187 7391 8423 7627
rect 8508 7391 8744 7627
rect 8829 7391 9065 7627
rect 9150 7391 9386 7627
rect 9471 7391 9707 7627
rect 9792 7391 10028 7627
rect 10113 7391 10349 7627
rect 10434 7391 10670 7627
rect 10755 7391 10991 7627
rect 11076 7391 11312 7627
rect 11397 7391 11633 7627
rect 11718 7391 11954 7627
rect 12039 7391 12275 7627
rect 12359 7391 12595 7627
rect 12679 7391 12915 7627
rect 12999 7391 13235 7627
rect 13319 7391 13555 7627
rect 13639 7391 13875 7627
rect 13959 7391 14195 7627
rect 14279 7391 14515 7627
rect 14599 7391 14835 7627
rect 14919 7391 15155 7627
rect 15239 7391 15475 7627
rect 15559 7391 15795 7627
rect 162 6787 398 7023
rect 483 6787 719 7023
rect 804 6787 1040 7023
rect 1125 6787 1361 7023
rect 1446 6787 1682 7023
rect 1767 6787 2003 7023
rect 2088 6787 2324 7023
rect 2409 6787 2645 7023
rect 2730 6787 2966 7023
rect 3051 6787 3287 7023
rect 3372 6787 3608 7023
rect 3693 6787 3929 7023
rect 4014 6787 4250 7023
rect 4335 6787 4571 7023
rect 4656 6787 4892 7023
rect 4977 6787 5213 7023
rect 5298 6787 5534 7023
rect 5619 6787 5855 7023
rect 5940 6787 6176 7023
rect 6261 6787 6497 7023
rect 6582 6787 6818 7023
rect 6903 6787 7139 7023
rect 7224 6787 7460 7023
rect 7545 6787 7781 7023
rect 7866 6787 8102 7023
rect 8187 6787 8423 7023
rect 8508 6787 8744 7023
rect 8829 6787 9065 7023
rect 9150 6787 9386 7023
rect 9471 6787 9707 7023
rect 9792 6787 10028 7023
rect 10113 6787 10349 7023
rect 10434 6787 10670 7023
rect 10755 6787 10991 7023
rect 11076 6787 11312 7023
rect 11397 6787 11633 7023
rect 11718 6787 11954 7023
rect 12038 6787 12274 7023
rect 12358 6787 12594 7023
rect 12678 6787 12914 7023
rect 12998 6787 13234 7023
rect 13318 6787 13554 7023
rect 13638 6787 13874 7023
rect 13958 6787 14194 7023
rect 14278 6787 14514 7023
rect 14598 6787 14834 7023
rect 14918 6787 15154 7023
rect 15238 6787 15474 7023
rect 15558 6787 15794 7023
rect 162 6421 398 6657
rect 483 6421 719 6657
rect 804 6421 1040 6657
rect 1125 6421 1361 6657
rect 1446 6421 1682 6657
rect 1767 6421 2003 6657
rect 2088 6421 2324 6657
rect 2409 6421 2645 6657
rect 2730 6421 2966 6657
rect 3051 6421 3287 6657
rect 3372 6421 3608 6657
rect 3693 6421 3929 6657
rect 4014 6421 4250 6657
rect 4335 6421 4571 6657
rect 4656 6421 4892 6657
rect 4977 6421 5213 6657
rect 5298 6421 5534 6657
rect 5619 6421 5855 6657
rect 5940 6421 6176 6657
rect 6261 6421 6497 6657
rect 6582 6421 6818 6657
rect 6903 6421 7139 6657
rect 7224 6421 7460 6657
rect 7545 6421 7781 6657
rect 7866 6421 8102 6657
rect 8187 6421 8423 6657
rect 8508 6421 8744 6657
rect 8829 6421 9065 6657
rect 9150 6421 9386 6657
rect 9471 6421 9707 6657
rect 9792 6421 10028 6657
rect 10113 6421 10349 6657
rect 10434 6421 10670 6657
rect 10755 6421 10991 6657
rect 11076 6421 11312 6657
rect 11397 6421 11633 6657
rect 11718 6421 11954 6657
rect 12038 6421 12274 6657
rect 12358 6421 12594 6657
rect 12678 6421 12914 6657
rect 12998 6421 13234 6657
rect 13318 6421 13554 6657
rect 13638 6421 13874 6657
rect 13958 6421 14194 6657
rect 14278 6421 14514 6657
rect 14598 6421 14834 6657
rect 14918 6421 15154 6657
rect 15238 6421 15474 6657
rect 15558 6421 15794 6657
rect 161 5817 397 6053
rect 482 5817 718 6053
rect 803 5817 1039 6053
rect 1124 5817 1360 6053
rect 1445 5817 1681 6053
rect 1766 5817 2002 6053
rect 2087 5817 2323 6053
rect 2408 5817 2644 6053
rect 2729 5817 2965 6053
rect 3050 5817 3286 6053
rect 3371 5817 3607 6053
rect 3692 5817 3928 6053
rect 4013 5817 4249 6053
rect 4334 5817 4570 6053
rect 4655 5817 4891 6053
rect 4976 5817 5212 6053
rect 5297 5817 5533 6053
rect 5618 5817 5854 6053
rect 5939 5817 6175 6053
rect 6260 5817 6496 6053
rect 6581 5817 6817 6053
rect 6902 5817 7138 6053
rect 7223 5817 7459 6053
rect 7544 5817 7780 6053
rect 7865 5817 8101 6053
rect 8186 5817 8422 6053
rect 8507 5817 8743 6053
rect 8828 5817 9064 6053
rect 9149 5817 9385 6053
rect 9470 5817 9706 6053
rect 9791 5817 10027 6053
rect 10112 5817 10348 6053
rect 10433 5817 10669 6053
rect 10754 5817 10990 6053
rect 11075 5817 11311 6053
rect 11396 5817 11632 6053
rect 11717 5817 11953 6053
rect 12038 5817 12274 6053
rect 12358 5817 12594 6053
rect 12678 5817 12914 6053
rect 12998 5817 13234 6053
rect 13318 5817 13554 6053
rect 13638 5817 13874 6053
rect 13958 5817 14194 6053
rect 14278 5817 14514 6053
rect 14598 5817 14834 6053
rect 14918 5817 15154 6053
rect 15238 5817 15474 6053
rect 15558 5817 15794 6053
rect 161 5211 397 5447
rect 482 5211 718 5447
rect 803 5211 1039 5447
rect 1124 5211 1360 5447
rect 1445 5211 1681 5447
rect 1766 5211 2002 5447
rect 2087 5211 2323 5447
rect 2408 5211 2644 5447
rect 2729 5211 2965 5447
rect 3050 5211 3286 5447
rect 3371 5211 3607 5447
rect 3692 5211 3928 5447
rect 4013 5211 4249 5447
rect 4334 5211 4570 5447
rect 4655 5211 4891 5447
rect 4976 5211 5212 5447
rect 5297 5211 5533 5447
rect 5618 5211 5854 5447
rect 5939 5211 6175 5447
rect 6260 5211 6496 5447
rect 6581 5211 6817 5447
rect 6902 5211 7138 5447
rect 7223 5211 7459 5447
rect 7544 5211 7780 5447
rect 7865 5211 8101 5447
rect 8186 5211 8422 5447
rect 8507 5211 8743 5447
rect 8828 5211 9064 5447
rect 9149 5211 9385 5447
rect 9470 5211 9706 5447
rect 9791 5211 10027 5447
rect 10112 5211 10348 5447
rect 10433 5211 10669 5447
rect 10754 5211 10990 5447
rect 11075 5211 11311 5447
rect 11396 5211 11632 5447
rect 11717 5211 11953 5447
rect 12038 5211 12274 5447
rect 12358 5211 12594 5447
rect 12678 5211 12914 5447
rect 12998 5211 13234 5447
rect 13318 5211 13554 5447
rect 13638 5211 13874 5447
rect 13958 5211 14194 5447
rect 14278 5211 14514 5447
rect 14598 5211 14834 5447
rect 14918 5211 15154 5447
rect 15238 5211 15474 5447
rect 15558 5211 15794 5447
rect 161 4607 397 4843
rect 482 4607 718 4843
rect 803 4607 1039 4843
rect 1124 4607 1360 4843
rect 1445 4607 1681 4843
rect 1766 4607 2002 4843
rect 2087 4607 2323 4843
rect 2408 4607 2644 4843
rect 2729 4607 2965 4843
rect 3050 4607 3286 4843
rect 3371 4607 3607 4843
rect 3692 4607 3928 4843
rect 4013 4607 4249 4843
rect 4334 4607 4570 4843
rect 4655 4607 4891 4843
rect 4976 4607 5212 4843
rect 5297 4607 5533 4843
rect 5618 4607 5854 4843
rect 5939 4607 6175 4843
rect 6260 4607 6496 4843
rect 6581 4607 6817 4843
rect 6902 4607 7138 4843
rect 7223 4607 7459 4843
rect 7544 4607 7780 4843
rect 7865 4607 8101 4843
rect 8186 4607 8422 4843
rect 8507 4607 8743 4843
rect 8828 4607 9064 4843
rect 9149 4607 9385 4843
rect 9470 4607 9706 4843
rect 9791 4607 10027 4843
rect 10112 4607 10348 4843
rect 10433 4607 10669 4843
rect 10754 4607 10990 4843
rect 11075 4607 11311 4843
rect 11396 4607 11632 4843
rect 11717 4607 11953 4843
rect 12037 4607 12273 4843
rect 12357 4607 12593 4843
rect 12677 4607 12913 4843
rect 12997 4607 13233 4843
rect 13317 4607 13553 4843
rect 13637 4607 13873 4843
rect 13957 4607 14193 4843
rect 14277 4607 14513 4843
rect 14597 4607 14833 4843
rect 14917 4607 15153 4843
rect 15237 4607 15473 4843
rect 15557 4607 15793 4843
rect 161 4001 397 4237
rect 482 4001 718 4237
rect 803 4001 1039 4237
rect 1124 4001 1360 4237
rect 1445 4001 1681 4237
rect 1766 4001 2002 4237
rect 2087 4001 2323 4237
rect 2408 4001 2644 4237
rect 2729 4001 2965 4237
rect 3050 4001 3286 4237
rect 3371 4001 3607 4237
rect 3692 4001 3928 4237
rect 4013 4001 4249 4237
rect 4334 4001 4570 4237
rect 4655 4001 4891 4237
rect 4976 4001 5212 4237
rect 5297 4001 5533 4237
rect 5618 4001 5854 4237
rect 5939 4001 6175 4237
rect 6260 4001 6496 4237
rect 6581 4001 6817 4237
rect 6902 4001 7138 4237
rect 7223 4001 7459 4237
rect 7544 4001 7780 4237
rect 7865 4001 8101 4237
rect 8186 4001 8422 4237
rect 8507 4001 8743 4237
rect 8828 4001 9064 4237
rect 9149 4001 9385 4237
rect 9470 4001 9706 4237
rect 9791 4001 10027 4237
rect 10112 4001 10348 4237
rect 10433 4001 10669 4237
rect 10754 4001 10990 4237
rect 11075 4001 11311 4237
rect 11396 4001 11632 4237
rect 11717 4001 11953 4237
rect 12037 4001 12273 4237
rect 12357 4001 12593 4237
rect 12677 4001 12913 4237
rect 12997 4001 13233 4237
rect 13317 4001 13553 4237
rect 13637 4001 13873 4237
rect 13957 4001 14193 4237
rect 14277 4001 14513 4237
rect 14597 4001 14833 4237
rect 14917 4001 15153 4237
rect 15237 4001 15473 4237
rect 15557 4001 15793 4237
rect 162 3397 398 3633
rect 483 3397 719 3633
rect 804 3397 1040 3633
rect 1125 3397 1361 3633
rect 1446 3397 1682 3633
rect 1767 3397 2003 3633
rect 2088 3397 2324 3633
rect 2409 3397 2645 3633
rect 2730 3397 2966 3633
rect 3051 3397 3287 3633
rect 3372 3397 3608 3633
rect 3693 3397 3929 3633
rect 4014 3397 4250 3633
rect 4335 3397 4571 3633
rect 4656 3397 4892 3633
rect 4977 3397 5213 3633
rect 5298 3397 5534 3633
rect 5619 3397 5855 3633
rect 5940 3397 6176 3633
rect 6261 3397 6497 3633
rect 6582 3397 6818 3633
rect 6903 3397 7139 3633
rect 7224 3397 7460 3633
rect 7545 3397 7781 3633
rect 7866 3397 8102 3633
rect 8187 3397 8423 3633
rect 8508 3397 8744 3633
rect 8829 3397 9065 3633
rect 9150 3397 9386 3633
rect 9471 3397 9707 3633
rect 9792 3397 10028 3633
rect 10113 3397 10349 3633
rect 10434 3397 10670 3633
rect 10755 3397 10991 3633
rect 11076 3397 11312 3633
rect 11397 3397 11633 3633
rect 11718 3397 11954 3633
rect 12038 3397 12274 3633
rect 12358 3397 12594 3633
rect 12678 3397 12914 3633
rect 12998 3397 13234 3633
rect 13318 3397 13554 3633
rect 13638 3397 13874 3633
rect 13958 3397 14194 3633
rect 14278 3397 14514 3633
rect 14598 3397 14834 3633
rect 14918 3397 15154 3633
rect 15238 3397 15474 3633
rect 15558 3397 15794 3633
rect 162 3031 398 3267
rect 483 3031 719 3267
rect 804 3031 1040 3267
rect 1125 3031 1361 3267
rect 1446 3031 1682 3267
rect 1767 3031 2003 3267
rect 2088 3031 2324 3267
rect 2409 3031 2645 3267
rect 2730 3031 2966 3267
rect 3051 3031 3287 3267
rect 3372 3031 3608 3267
rect 3693 3031 3929 3267
rect 4014 3031 4250 3267
rect 4335 3031 4571 3267
rect 4656 3031 4892 3267
rect 4977 3031 5213 3267
rect 5298 3031 5534 3267
rect 5619 3031 5855 3267
rect 5940 3031 6176 3267
rect 6261 3031 6497 3267
rect 6582 3031 6818 3267
rect 6903 3031 7139 3267
rect 7224 3031 7460 3267
rect 7545 3031 7781 3267
rect 7866 3031 8102 3267
rect 8187 3031 8423 3267
rect 8508 3031 8744 3267
rect 8829 3031 9065 3267
rect 9150 3031 9386 3267
rect 9471 3031 9707 3267
rect 9792 3031 10028 3267
rect 10113 3031 10349 3267
rect 10434 3031 10670 3267
rect 10755 3031 10991 3267
rect 11076 3031 11312 3267
rect 11397 3031 11633 3267
rect 11718 3031 11954 3267
rect 12038 3031 12274 3267
rect 12358 3031 12594 3267
rect 12678 3031 12914 3267
rect 12998 3031 13234 3267
rect 13318 3031 13554 3267
rect 13638 3031 13874 3267
rect 13958 3031 14194 3267
rect 14278 3031 14514 3267
rect 14598 3031 14834 3267
rect 14918 3031 15154 3267
rect 15238 3031 15474 3267
rect 15558 3031 15794 3267
rect 163 2427 399 2663
rect 484 2427 720 2663
rect 805 2427 1041 2663
rect 1126 2427 1362 2663
rect 1447 2427 1683 2663
rect 1768 2427 2004 2663
rect 2089 2427 2325 2663
rect 2410 2427 2646 2663
rect 2731 2427 2967 2663
rect 3052 2427 3288 2663
rect 3373 2427 3609 2663
rect 3694 2427 3930 2663
rect 4015 2427 4251 2663
rect 4336 2427 4572 2663
rect 4657 2427 4893 2663
rect 4978 2427 5214 2663
rect 5299 2427 5535 2663
rect 5620 2427 5856 2663
rect 5941 2427 6177 2663
rect 6262 2427 6498 2663
rect 6583 2427 6819 2663
rect 6904 2427 7140 2663
rect 7225 2427 7461 2663
rect 7546 2427 7782 2663
rect 7867 2427 8103 2663
rect 8188 2427 8424 2663
rect 8509 2427 8745 2663
rect 8830 2427 9066 2663
rect 9151 2427 9387 2663
rect 9472 2427 9708 2663
rect 9793 2427 10029 2663
rect 10114 2427 10350 2663
rect 10435 2427 10671 2663
rect 10756 2427 10992 2663
rect 11077 2427 11313 2663
rect 11397 2427 11633 2663
rect 11717 2427 11953 2663
rect 12037 2427 12273 2663
rect 12357 2427 12593 2663
rect 12677 2427 12913 2663
rect 12997 2427 13233 2663
rect 13317 2427 13553 2663
rect 13637 2427 13873 2663
rect 13957 2427 14193 2663
rect 14277 2427 14513 2663
rect 14597 2427 14833 2663
rect 14917 2427 15153 2663
rect 15237 2427 15473 2663
rect 15557 2427 15793 2663
rect 163 1821 399 2057
rect 484 1821 720 2057
rect 805 1821 1041 2057
rect 1126 1821 1362 2057
rect 1447 1821 1683 2057
rect 1768 1821 2004 2057
rect 2089 1821 2325 2057
rect 2410 1821 2646 2057
rect 2731 1821 2967 2057
rect 3052 1821 3288 2057
rect 3373 1821 3609 2057
rect 3694 1821 3930 2057
rect 4015 1821 4251 2057
rect 4336 1821 4572 2057
rect 4657 1821 4893 2057
rect 4978 1821 5214 2057
rect 5299 1821 5535 2057
rect 5620 1821 5856 2057
rect 5941 1821 6177 2057
rect 6262 1821 6498 2057
rect 6583 1821 6819 2057
rect 6904 1821 7140 2057
rect 7225 1821 7461 2057
rect 7546 1821 7782 2057
rect 7867 1821 8103 2057
rect 8188 1821 8424 2057
rect 8509 1821 8745 2057
rect 8830 1821 9066 2057
rect 9151 1821 9387 2057
rect 9472 1821 9708 2057
rect 9793 1821 10029 2057
rect 10114 1821 10350 2057
rect 10435 1821 10671 2057
rect 10756 1821 10992 2057
rect 11077 1821 11313 2057
rect 11397 1821 11633 2057
rect 11717 1821 11953 2057
rect 12037 1821 12273 2057
rect 12357 1821 12593 2057
rect 12677 1821 12913 2057
rect 12997 1821 13233 2057
rect 13317 1821 13553 2057
rect 13637 1821 13873 2057
rect 13957 1821 14193 2057
rect 14277 1821 14513 2057
rect 14597 1821 14833 2057
rect 14917 1821 15153 2057
rect 15237 1821 15473 2057
rect 15557 1821 15793 2057
rect 162 1216 398 1452
rect 483 1216 719 1452
rect 804 1216 1040 1452
rect 1125 1216 1361 1452
rect 1446 1216 1682 1452
rect 1767 1216 2003 1452
rect 2088 1216 2324 1452
rect 2409 1216 2645 1452
rect 2730 1216 2966 1452
rect 3051 1216 3287 1452
rect 3372 1216 3608 1452
rect 3693 1216 3929 1452
rect 4014 1216 4250 1452
rect 4335 1216 4571 1452
rect 4656 1216 4892 1452
rect 4977 1216 5213 1452
rect 5298 1216 5534 1452
rect 5619 1216 5855 1452
rect 5940 1216 6176 1452
rect 6261 1216 6497 1452
rect 6582 1216 6818 1452
rect 6903 1216 7139 1452
rect 7224 1216 7460 1452
rect 7545 1216 7781 1452
rect 7866 1216 8102 1452
rect 8187 1216 8423 1452
rect 8508 1216 8744 1452
rect 8829 1216 9065 1452
rect 9150 1216 9386 1452
rect 9471 1216 9707 1452
rect 9792 1216 10028 1452
rect 10113 1216 10349 1452
rect 10434 1216 10670 1452
rect 10755 1216 10991 1452
rect 11076 1216 11312 1452
rect 11397 1216 11633 1452
rect 11718 1216 11954 1452
rect 12038 1216 12274 1452
rect 12358 1216 12594 1452
rect 12678 1216 12914 1452
rect 12998 1216 13234 1452
rect 13318 1216 13554 1452
rect 13638 1216 13874 1452
rect 13958 1216 14194 1452
rect 14278 1216 14514 1452
rect 14598 1216 14834 1452
rect 14918 1216 15154 1452
rect 15238 1216 15474 1452
rect 15558 1216 15794 1452
rect 162 834 398 1070
rect 483 834 719 1070
rect 804 834 1040 1070
rect 1125 834 1361 1070
rect 1446 834 1682 1070
rect 1767 834 2003 1070
rect 2088 834 2324 1070
rect 2409 834 2645 1070
rect 2730 834 2966 1070
rect 3051 834 3287 1070
rect 3372 834 3608 1070
rect 3693 834 3929 1070
rect 4014 834 4250 1070
rect 4335 834 4571 1070
rect 4656 834 4892 1070
rect 4977 834 5213 1070
rect 5298 834 5534 1070
rect 5619 834 5855 1070
rect 5940 834 6176 1070
rect 6261 834 6497 1070
rect 6582 834 6818 1070
rect 6903 834 7139 1070
rect 7224 834 7460 1070
rect 7545 834 7781 1070
rect 7866 834 8102 1070
rect 8187 834 8423 1070
rect 8508 834 8744 1070
rect 8829 834 9065 1070
rect 9150 834 9386 1070
rect 9471 834 9707 1070
rect 9792 834 10028 1070
rect 10113 834 10349 1070
rect 10434 834 10670 1070
rect 10755 834 10991 1070
rect 11076 834 11312 1070
rect 11397 834 11633 1070
rect 11718 834 11954 1070
rect 12038 834 12274 1070
rect 12358 834 12594 1070
rect 12678 834 12914 1070
rect 12998 834 13234 1070
rect 13318 834 13554 1070
rect 13638 834 13874 1070
rect 13958 834 14194 1070
rect 14278 834 14514 1070
rect 14598 834 14834 1070
rect 14918 834 15154 1070
rect 15238 834 15474 1070
rect 15558 834 15794 1070
rect 162 452 398 688
rect 483 452 719 688
rect 804 452 1040 688
rect 1125 452 1361 688
rect 1446 452 1682 688
rect 1767 452 2003 688
rect 2088 452 2324 688
rect 2409 452 2645 688
rect 2730 452 2966 688
rect 3051 452 3287 688
rect 3372 452 3608 688
rect 3693 452 3929 688
rect 4014 452 4250 688
rect 4335 452 4571 688
rect 4656 452 4892 688
rect 4977 452 5213 688
rect 5298 452 5534 688
rect 5619 452 5855 688
rect 5940 452 6176 688
rect 6261 452 6497 688
rect 6582 452 6818 688
rect 6903 452 7139 688
rect 7224 452 7460 688
rect 7545 452 7781 688
rect 7866 452 8102 688
rect 8187 452 8423 688
rect 8508 452 8744 688
rect 8829 452 9065 688
rect 9150 452 9386 688
rect 9471 452 9707 688
rect 9792 452 10028 688
rect 10113 452 10349 688
rect 10434 452 10670 688
rect 10755 452 10991 688
rect 11076 452 11312 688
rect 11397 452 11633 688
rect 11718 452 11954 688
rect 12038 452 12274 688
rect 12358 452 12594 688
rect 12678 452 12914 688
rect 12998 452 13234 688
rect 13318 452 13554 688
rect 13638 452 13874 688
rect 13958 452 14194 688
rect 14278 452 14514 688
rect 14598 452 14834 688
rect 14918 452 15154 688
rect 15238 452 15474 688
rect 15558 452 15794 688
<< metal5 >>
rect 0 39965 16000 40000
rect 0 39729 162 39965
rect 398 39729 483 39965
rect 719 39729 804 39965
rect 1040 39729 1125 39965
rect 1361 39729 1446 39965
rect 1682 39729 1767 39965
rect 2003 39729 2088 39965
rect 2324 39729 2409 39965
rect 2645 39729 2730 39965
rect 2966 39729 3051 39965
rect 3287 39729 3372 39965
rect 3608 39729 3693 39965
rect 3929 39729 4014 39965
rect 4250 39729 4335 39965
rect 4571 39729 4656 39965
rect 4892 39729 4977 39965
rect 5213 39729 5298 39965
rect 5534 39729 5619 39965
rect 5855 39729 5940 39965
rect 6176 39729 6261 39965
rect 6497 39729 6582 39965
rect 6818 39729 6903 39965
rect 7139 39729 7224 39965
rect 7460 39729 7545 39965
rect 7781 39729 7866 39965
rect 8102 39729 8187 39965
rect 8423 39729 8508 39965
rect 8744 39729 8829 39965
rect 9065 39729 9150 39965
rect 9386 39729 9471 39965
rect 9707 39729 9792 39965
rect 10028 39729 10113 39965
rect 10349 39729 10434 39965
rect 10670 39729 10755 39965
rect 10991 39729 11076 39965
rect 11312 39729 11397 39965
rect 11633 39729 11718 39965
rect 11954 39729 12038 39965
rect 12274 39729 12358 39965
rect 12594 39729 12678 39965
rect 12914 39729 12998 39965
rect 13234 39729 13318 39965
rect 13554 39729 13638 39965
rect 13874 39729 13958 39965
rect 14194 39729 14278 39965
rect 14514 39729 14598 39965
rect 14834 39729 14918 39965
rect 15154 39729 15238 39965
rect 15474 39729 15558 39965
rect 15794 39729 16000 39965
rect 0 39641 16000 39729
rect 0 39405 162 39641
rect 398 39405 483 39641
rect 719 39405 804 39641
rect 1040 39405 1125 39641
rect 1361 39405 1446 39641
rect 1682 39405 1767 39641
rect 2003 39405 2088 39641
rect 2324 39405 2409 39641
rect 2645 39405 2730 39641
rect 2966 39405 3051 39641
rect 3287 39405 3372 39641
rect 3608 39405 3693 39641
rect 3929 39405 4014 39641
rect 4250 39405 4335 39641
rect 4571 39405 4656 39641
rect 4892 39405 4977 39641
rect 5213 39405 5298 39641
rect 5534 39405 5619 39641
rect 5855 39405 5940 39641
rect 6176 39405 6261 39641
rect 6497 39405 6582 39641
rect 6818 39405 6903 39641
rect 7139 39405 7224 39641
rect 7460 39405 7545 39641
rect 7781 39405 7866 39641
rect 8102 39405 8187 39641
rect 8423 39405 8508 39641
rect 8744 39405 8829 39641
rect 9065 39405 9150 39641
rect 9386 39405 9471 39641
rect 9707 39405 9792 39641
rect 10028 39405 10113 39641
rect 10349 39405 10434 39641
rect 10670 39405 10755 39641
rect 10991 39405 11076 39641
rect 11312 39405 11397 39641
rect 11633 39405 11718 39641
rect 11954 39405 12038 39641
rect 12274 39405 12358 39641
rect 12594 39405 12678 39641
rect 12914 39405 12998 39641
rect 13234 39405 13318 39641
rect 13554 39405 13638 39641
rect 13874 39405 13958 39641
rect 14194 39405 14278 39641
rect 14514 39405 14598 39641
rect 14834 39405 14918 39641
rect 15154 39405 15238 39641
rect 15474 39405 15558 39641
rect 15794 39405 16000 39641
rect 0 39317 16000 39405
rect 0 39081 162 39317
rect 398 39081 483 39317
rect 719 39081 804 39317
rect 1040 39081 1125 39317
rect 1361 39081 1446 39317
rect 1682 39081 1767 39317
rect 2003 39081 2088 39317
rect 2324 39081 2409 39317
rect 2645 39081 2730 39317
rect 2966 39081 3051 39317
rect 3287 39081 3372 39317
rect 3608 39081 3693 39317
rect 3929 39081 4014 39317
rect 4250 39081 4335 39317
rect 4571 39081 4656 39317
rect 4892 39081 4977 39317
rect 5213 39081 5298 39317
rect 5534 39081 5619 39317
rect 5855 39081 5940 39317
rect 6176 39081 6261 39317
rect 6497 39081 6582 39317
rect 6818 39081 6903 39317
rect 7139 39081 7224 39317
rect 7460 39081 7545 39317
rect 7781 39081 7866 39317
rect 8102 39081 8187 39317
rect 8423 39081 8508 39317
rect 8744 39081 8829 39317
rect 9065 39081 9150 39317
rect 9386 39081 9471 39317
rect 9707 39081 9792 39317
rect 10028 39081 10113 39317
rect 10349 39081 10434 39317
rect 10670 39081 10755 39317
rect 10991 39081 11076 39317
rect 11312 39081 11397 39317
rect 11633 39081 11718 39317
rect 11954 39081 12038 39317
rect 12274 39081 12358 39317
rect 12594 39081 12678 39317
rect 12914 39081 12998 39317
rect 13234 39081 13318 39317
rect 13554 39081 13638 39317
rect 13874 39081 13958 39317
rect 14194 39081 14278 39317
rect 14514 39081 14598 39317
rect 14834 39081 14918 39317
rect 15154 39081 15238 39317
rect 15474 39081 15558 39317
rect 15794 39081 16000 39317
rect 0 38993 16000 39081
rect 0 38757 162 38993
rect 398 38757 483 38993
rect 719 38757 804 38993
rect 1040 38757 1125 38993
rect 1361 38757 1446 38993
rect 1682 38757 1767 38993
rect 2003 38757 2088 38993
rect 2324 38757 2409 38993
rect 2645 38757 2730 38993
rect 2966 38757 3051 38993
rect 3287 38757 3372 38993
rect 3608 38757 3693 38993
rect 3929 38757 4014 38993
rect 4250 38757 4335 38993
rect 4571 38757 4656 38993
rect 4892 38757 4977 38993
rect 5213 38757 5298 38993
rect 5534 38757 5619 38993
rect 5855 38757 5940 38993
rect 6176 38757 6261 38993
rect 6497 38757 6582 38993
rect 6818 38757 6903 38993
rect 7139 38757 7224 38993
rect 7460 38757 7545 38993
rect 7781 38757 7866 38993
rect 8102 38757 8187 38993
rect 8423 38757 8508 38993
rect 8744 38757 8829 38993
rect 9065 38757 9150 38993
rect 9386 38757 9471 38993
rect 9707 38757 9792 38993
rect 10028 38757 10113 38993
rect 10349 38757 10434 38993
rect 10670 38757 10755 38993
rect 10991 38757 11076 38993
rect 11312 38757 11397 38993
rect 11633 38757 11718 38993
rect 11954 38757 12038 38993
rect 12274 38757 12358 38993
rect 12594 38757 12678 38993
rect 12914 38757 12998 38993
rect 13234 38757 13318 38993
rect 13554 38757 13638 38993
rect 13874 38757 13958 38993
rect 14194 38757 14278 38993
rect 14514 38757 14598 38993
rect 14834 38757 14918 38993
rect 15154 38757 15238 38993
rect 15474 38757 15558 38993
rect 15794 38757 16000 38993
rect 0 38669 16000 38757
rect 0 38433 162 38669
rect 398 38433 483 38669
rect 719 38433 804 38669
rect 1040 38433 1125 38669
rect 1361 38433 1446 38669
rect 1682 38433 1767 38669
rect 2003 38433 2088 38669
rect 2324 38433 2409 38669
rect 2645 38433 2730 38669
rect 2966 38433 3051 38669
rect 3287 38433 3372 38669
rect 3608 38433 3693 38669
rect 3929 38433 4014 38669
rect 4250 38433 4335 38669
rect 4571 38433 4656 38669
rect 4892 38433 4977 38669
rect 5213 38433 5298 38669
rect 5534 38433 5619 38669
rect 5855 38433 5940 38669
rect 6176 38433 6261 38669
rect 6497 38433 6582 38669
rect 6818 38433 6903 38669
rect 7139 38433 7224 38669
rect 7460 38433 7545 38669
rect 7781 38433 7866 38669
rect 8102 38433 8187 38669
rect 8423 38433 8508 38669
rect 8744 38433 8829 38669
rect 9065 38433 9150 38669
rect 9386 38433 9471 38669
rect 9707 38433 9792 38669
rect 10028 38433 10113 38669
rect 10349 38433 10434 38669
rect 10670 38433 10755 38669
rect 10991 38433 11076 38669
rect 11312 38433 11397 38669
rect 11633 38433 11718 38669
rect 11954 38433 12038 38669
rect 12274 38433 12358 38669
rect 12594 38433 12678 38669
rect 12914 38433 12998 38669
rect 13234 38433 13318 38669
rect 13554 38433 13638 38669
rect 13874 38433 13958 38669
rect 14194 38433 14278 38669
rect 14514 38433 14598 38669
rect 14834 38433 14918 38669
rect 15154 38433 15238 38669
rect 15474 38433 15558 38669
rect 15794 38433 16000 38669
rect 0 38345 16000 38433
rect 0 38109 162 38345
rect 398 38109 483 38345
rect 719 38109 804 38345
rect 1040 38109 1125 38345
rect 1361 38109 1446 38345
rect 1682 38109 1767 38345
rect 2003 38109 2088 38345
rect 2324 38109 2409 38345
rect 2645 38109 2730 38345
rect 2966 38109 3051 38345
rect 3287 38109 3372 38345
rect 3608 38109 3693 38345
rect 3929 38109 4014 38345
rect 4250 38109 4335 38345
rect 4571 38109 4656 38345
rect 4892 38109 4977 38345
rect 5213 38109 5298 38345
rect 5534 38109 5619 38345
rect 5855 38109 5940 38345
rect 6176 38109 6261 38345
rect 6497 38109 6582 38345
rect 6818 38109 6903 38345
rect 7139 38109 7224 38345
rect 7460 38109 7545 38345
rect 7781 38109 7866 38345
rect 8102 38109 8187 38345
rect 8423 38109 8508 38345
rect 8744 38109 8829 38345
rect 9065 38109 9150 38345
rect 9386 38109 9471 38345
rect 9707 38109 9792 38345
rect 10028 38109 10113 38345
rect 10349 38109 10434 38345
rect 10670 38109 10755 38345
rect 10991 38109 11076 38345
rect 11312 38109 11397 38345
rect 11633 38109 11718 38345
rect 11954 38109 12038 38345
rect 12274 38109 12358 38345
rect 12594 38109 12678 38345
rect 12914 38109 12998 38345
rect 13234 38109 13318 38345
rect 13554 38109 13638 38345
rect 13874 38109 13958 38345
rect 14194 38109 14278 38345
rect 14514 38109 14598 38345
rect 14834 38109 14918 38345
rect 15154 38109 15238 38345
rect 15474 38109 15558 38345
rect 15794 38109 16000 38345
rect 0 38021 16000 38109
rect 0 37785 162 38021
rect 398 37785 483 38021
rect 719 37785 804 38021
rect 1040 37785 1125 38021
rect 1361 37785 1446 38021
rect 1682 37785 1767 38021
rect 2003 37785 2088 38021
rect 2324 37785 2409 38021
rect 2645 37785 2730 38021
rect 2966 37785 3051 38021
rect 3287 37785 3372 38021
rect 3608 37785 3693 38021
rect 3929 37785 4014 38021
rect 4250 37785 4335 38021
rect 4571 37785 4656 38021
rect 4892 37785 4977 38021
rect 5213 37785 5298 38021
rect 5534 37785 5619 38021
rect 5855 37785 5940 38021
rect 6176 37785 6261 38021
rect 6497 37785 6582 38021
rect 6818 37785 6903 38021
rect 7139 37785 7224 38021
rect 7460 37785 7545 38021
rect 7781 37785 7866 38021
rect 8102 37785 8187 38021
rect 8423 37785 8508 38021
rect 8744 37785 8829 38021
rect 9065 37785 9150 38021
rect 9386 37785 9471 38021
rect 9707 37785 9792 38021
rect 10028 37785 10113 38021
rect 10349 37785 10434 38021
rect 10670 37785 10755 38021
rect 10991 37785 11076 38021
rect 11312 37785 11397 38021
rect 11633 37785 11718 38021
rect 11954 37785 12038 38021
rect 12274 37785 12358 38021
rect 12594 37785 12678 38021
rect 12914 37785 12998 38021
rect 13234 37785 13318 38021
rect 13554 37785 13638 38021
rect 13874 37785 13958 38021
rect 14194 37785 14278 38021
rect 14514 37785 14598 38021
rect 14834 37785 14918 38021
rect 15154 37785 15238 38021
rect 15474 37785 15558 38021
rect 15794 37785 16000 38021
rect 0 37697 16000 37785
rect 0 37461 162 37697
rect 398 37461 483 37697
rect 719 37461 804 37697
rect 1040 37461 1125 37697
rect 1361 37461 1446 37697
rect 1682 37461 1767 37697
rect 2003 37461 2088 37697
rect 2324 37461 2409 37697
rect 2645 37461 2730 37697
rect 2966 37461 3051 37697
rect 3287 37461 3372 37697
rect 3608 37461 3693 37697
rect 3929 37461 4014 37697
rect 4250 37461 4335 37697
rect 4571 37461 4656 37697
rect 4892 37461 4977 37697
rect 5213 37461 5298 37697
rect 5534 37461 5619 37697
rect 5855 37461 5940 37697
rect 6176 37461 6261 37697
rect 6497 37461 6582 37697
rect 6818 37461 6903 37697
rect 7139 37461 7224 37697
rect 7460 37461 7545 37697
rect 7781 37461 7866 37697
rect 8102 37461 8187 37697
rect 8423 37461 8508 37697
rect 8744 37461 8829 37697
rect 9065 37461 9150 37697
rect 9386 37461 9471 37697
rect 9707 37461 9792 37697
rect 10028 37461 10113 37697
rect 10349 37461 10434 37697
rect 10670 37461 10755 37697
rect 10991 37461 11076 37697
rect 11312 37461 11397 37697
rect 11633 37461 11718 37697
rect 11954 37461 12038 37697
rect 12274 37461 12358 37697
rect 12594 37461 12678 37697
rect 12914 37461 12998 37697
rect 13234 37461 13318 37697
rect 13554 37461 13638 37697
rect 13874 37461 13958 37697
rect 14194 37461 14278 37697
rect 14514 37461 14598 37697
rect 14834 37461 14918 37697
rect 15154 37461 15238 37697
rect 15474 37461 15558 37697
rect 15794 37461 16000 37697
rect 0 37373 16000 37461
rect 0 37137 162 37373
rect 398 37137 483 37373
rect 719 37137 804 37373
rect 1040 37137 1125 37373
rect 1361 37137 1446 37373
rect 1682 37137 1767 37373
rect 2003 37137 2088 37373
rect 2324 37137 2409 37373
rect 2645 37137 2730 37373
rect 2966 37137 3051 37373
rect 3287 37137 3372 37373
rect 3608 37137 3693 37373
rect 3929 37137 4014 37373
rect 4250 37137 4335 37373
rect 4571 37137 4656 37373
rect 4892 37137 4977 37373
rect 5213 37137 5298 37373
rect 5534 37137 5619 37373
rect 5855 37137 5940 37373
rect 6176 37137 6261 37373
rect 6497 37137 6582 37373
rect 6818 37137 6903 37373
rect 7139 37137 7224 37373
rect 7460 37137 7545 37373
rect 7781 37137 7866 37373
rect 8102 37137 8187 37373
rect 8423 37137 8508 37373
rect 8744 37137 8829 37373
rect 9065 37137 9150 37373
rect 9386 37137 9471 37373
rect 9707 37137 9792 37373
rect 10028 37137 10113 37373
rect 10349 37137 10434 37373
rect 10670 37137 10755 37373
rect 10991 37137 11076 37373
rect 11312 37137 11397 37373
rect 11633 37137 11718 37373
rect 11954 37137 12038 37373
rect 12274 37137 12358 37373
rect 12594 37137 12678 37373
rect 12914 37137 12998 37373
rect 13234 37137 13318 37373
rect 13554 37137 13638 37373
rect 13874 37137 13958 37373
rect 14194 37137 14278 37373
rect 14514 37137 14598 37373
rect 14834 37137 14918 37373
rect 15154 37137 15238 37373
rect 15474 37137 15558 37373
rect 15794 37137 16000 37373
rect 0 37049 16000 37137
rect 0 36813 162 37049
rect 398 36813 483 37049
rect 719 36813 804 37049
rect 1040 36813 1125 37049
rect 1361 36813 1446 37049
rect 1682 36813 1767 37049
rect 2003 36813 2088 37049
rect 2324 36813 2409 37049
rect 2645 36813 2730 37049
rect 2966 36813 3051 37049
rect 3287 36813 3372 37049
rect 3608 36813 3693 37049
rect 3929 36813 4014 37049
rect 4250 36813 4335 37049
rect 4571 36813 4656 37049
rect 4892 36813 4977 37049
rect 5213 36813 5298 37049
rect 5534 36813 5619 37049
rect 5855 36813 5940 37049
rect 6176 36813 6261 37049
rect 6497 36813 6582 37049
rect 6818 36813 6903 37049
rect 7139 36813 7224 37049
rect 7460 36813 7545 37049
rect 7781 36813 7866 37049
rect 8102 36813 8187 37049
rect 8423 36813 8508 37049
rect 8744 36813 8829 37049
rect 9065 36813 9150 37049
rect 9386 36813 9471 37049
rect 9707 36813 9792 37049
rect 10028 36813 10113 37049
rect 10349 36813 10434 37049
rect 10670 36813 10755 37049
rect 10991 36813 11076 37049
rect 11312 36813 11397 37049
rect 11633 36813 11718 37049
rect 11954 36813 12038 37049
rect 12274 36813 12358 37049
rect 12594 36813 12678 37049
rect 12914 36813 12998 37049
rect 13234 36813 13318 37049
rect 13554 36813 13638 37049
rect 13874 36813 13958 37049
rect 14194 36813 14278 37049
rect 14514 36813 14598 37049
rect 14834 36813 14918 37049
rect 15154 36813 15238 37049
rect 15474 36813 15558 37049
rect 15794 36813 16000 37049
rect 0 36725 16000 36813
rect 0 36489 162 36725
rect 398 36489 483 36725
rect 719 36489 804 36725
rect 1040 36489 1125 36725
rect 1361 36489 1446 36725
rect 1682 36489 1767 36725
rect 2003 36489 2088 36725
rect 2324 36489 2409 36725
rect 2645 36489 2730 36725
rect 2966 36489 3051 36725
rect 3287 36489 3372 36725
rect 3608 36489 3693 36725
rect 3929 36489 4014 36725
rect 4250 36489 4335 36725
rect 4571 36489 4656 36725
rect 4892 36489 4977 36725
rect 5213 36489 5298 36725
rect 5534 36489 5619 36725
rect 5855 36489 5940 36725
rect 6176 36489 6261 36725
rect 6497 36489 6582 36725
rect 6818 36489 6903 36725
rect 7139 36489 7224 36725
rect 7460 36489 7545 36725
rect 7781 36489 7866 36725
rect 8102 36489 8187 36725
rect 8423 36489 8508 36725
rect 8744 36489 8829 36725
rect 9065 36489 9150 36725
rect 9386 36489 9471 36725
rect 9707 36489 9792 36725
rect 10028 36489 10113 36725
rect 10349 36489 10434 36725
rect 10670 36489 10755 36725
rect 10991 36489 11076 36725
rect 11312 36489 11397 36725
rect 11633 36489 11718 36725
rect 11954 36489 12038 36725
rect 12274 36489 12358 36725
rect 12594 36489 12678 36725
rect 12914 36489 12998 36725
rect 13234 36489 13318 36725
rect 13554 36489 13638 36725
rect 13874 36489 13958 36725
rect 14194 36489 14278 36725
rect 14514 36489 14598 36725
rect 14834 36489 14918 36725
rect 15154 36489 15238 36725
rect 15474 36489 15558 36725
rect 15794 36489 16000 36725
rect 0 36401 16000 36489
rect 0 36165 162 36401
rect 398 36165 483 36401
rect 719 36165 804 36401
rect 1040 36165 1125 36401
rect 1361 36165 1446 36401
rect 1682 36165 1767 36401
rect 2003 36165 2088 36401
rect 2324 36165 2409 36401
rect 2645 36165 2730 36401
rect 2966 36165 3051 36401
rect 3287 36165 3372 36401
rect 3608 36165 3693 36401
rect 3929 36165 4014 36401
rect 4250 36165 4335 36401
rect 4571 36165 4656 36401
rect 4892 36165 4977 36401
rect 5213 36165 5298 36401
rect 5534 36165 5619 36401
rect 5855 36165 5940 36401
rect 6176 36165 6261 36401
rect 6497 36165 6582 36401
rect 6818 36165 6903 36401
rect 7139 36165 7224 36401
rect 7460 36165 7545 36401
rect 7781 36165 7866 36401
rect 8102 36165 8187 36401
rect 8423 36165 8508 36401
rect 8744 36165 8829 36401
rect 9065 36165 9150 36401
rect 9386 36165 9471 36401
rect 9707 36165 9792 36401
rect 10028 36165 10113 36401
rect 10349 36165 10434 36401
rect 10670 36165 10755 36401
rect 10991 36165 11076 36401
rect 11312 36165 11397 36401
rect 11633 36165 11718 36401
rect 11954 36165 12038 36401
rect 12274 36165 12358 36401
rect 12594 36165 12678 36401
rect 12914 36165 12998 36401
rect 13234 36165 13318 36401
rect 13554 36165 13638 36401
rect 13874 36165 13958 36401
rect 14194 36165 14278 36401
rect 14514 36165 14598 36401
rect 14834 36165 14918 36401
rect 15154 36165 15238 36401
rect 15474 36165 15558 36401
rect 15794 36165 16000 36401
rect 0 36077 16000 36165
rect 0 35841 162 36077
rect 398 35841 483 36077
rect 719 35841 804 36077
rect 1040 35841 1125 36077
rect 1361 35841 1446 36077
rect 1682 35841 1767 36077
rect 2003 35841 2088 36077
rect 2324 35841 2409 36077
rect 2645 35841 2730 36077
rect 2966 35841 3051 36077
rect 3287 35841 3372 36077
rect 3608 35841 3693 36077
rect 3929 35841 4014 36077
rect 4250 35841 4335 36077
rect 4571 35841 4656 36077
rect 4892 35841 4977 36077
rect 5213 35841 5298 36077
rect 5534 35841 5619 36077
rect 5855 35841 5940 36077
rect 6176 35841 6261 36077
rect 6497 35841 6582 36077
rect 6818 35841 6903 36077
rect 7139 35841 7224 36077
rect 7460 35841 7545 36077
rect 7781 35841 7866 36077
rect 8102 35841 8187 36077
rect 8423 35841 8508 36077
rect 8744 35841 8829 36077
rect 9065 35841 9150 36077
rect 9386 35841 9471 36077
rect 9707 35841 9792 36077
rect 10028 35841 10113 36077
rect 10349 35841 10434 36077
rect 10670 35841 10755 36077
rect 10991 35841 11076 36077
rect 11312 35841 11397 36077
rect 11633 35841 11718 36077
rect 11954 35841 12038 36077
rect 12274 35841 12358 36077
rect 12594 35841 12678 36077
rect 12914 35841 12998 36077
rect 13234 35841 13318 36077
rect 13554 35841 13638 36077
rect 13874 35841 13958 36077
rect 14194 35841 14278 36077
rect 14514 35841 14598 36077
rect 14834 35841 14918 36077
rect 15154 35841 15238 36077
rect 15474 35841 15558 36077
rect 15794 35841 16000 36077
rect 0 35753 16000 35841
rect 0 35517 162 35753
rect 398 35517 483 35753
rect 719 35517 804 35753
rect 1040 35517 1125 35753
rect 1361 35517 1446 35753
rect 1682 35517 1767 35753
rect 2003 35517 2088 35753
rect 2324 35517 2409 35753
rect 2645 35517 2730 35753
rect 2966 35517 3051 35753
rect 3287 35517 3372 35753
rect 3608 35517 3693 35753
rect 3929 35517 4014 35753
rect 4250 35517 4335 35753
rect 4571 35517 4656 35753
rect 4892 35517 4977 35753
rect 5213 35517 5298 35753
rect 5534 35517 5619 35753
rect 5855 35517 5940 35753
rect 6176 35517 6261 35753
rect 6497 35517 6582 35753
rect 6818 35517 6903 35753
rect 7139 35517 7224 35753
rect 7460 35517 7545 35753
rect 7781 35517 7866 35753
rect 8102 35517 8187 35753
rect 8423 35517 8508 35753
rect 8744 35517 8829 35753
rect 9065 35517 9150 35753
rect 9386 35517 9471 35753
rect 9707 35517 9792 35753
rect 10028 35517 10113 35753
rect 10349 35517 10434 35753
rect 10670 35517 10755 35753
rect 10991 35517 11076 35753
rect 11312 35517 11397 35753
rect 11633 35517 11718 35753
rect 11954 35517 12038 35753
rect 12274 35517 12358 35753
rect 12594 35517 12678 35753
rect 12914 35517 12998 35753
rect 13234 35517 13318 35753
rect 13554 35517 13638 35753
rect 13874 35517 13958 35753
rect 14194 35517 14278 35753
rect 14514 35517 14598 35753
rect 14834 35517 14918 35753
rect 15154 35517 15238 35753
rect 15474 35517 15558 35753
rect 15794 35517 16000 35753
rect 0 35429 16000 35517
rect 0 35193 162 35429
rect 398 35193 483 35429
rect 719 35193 804 35429
rect 1040 35193 1125 35429
rect 1361 35193 1446 35429
rect 1682 35193 1767 35429
rect 2003 35193 2088 35429
rect 2324 35193 2409 35429
rect 2645 35193 2730 35429
rect 2966 35193 3051 35429
rect 3287 35193 3372 35429
rect 3608 35193 3693 35429
rect 3929 35193 4014 35429
rect 4250 35193 4335 35429
rect 4571 35193 4656 35429
rect 4892 35193 4977 35429
rect 5213 35193 5298 35429
rect 5534 35193 5619 35429
rect 5855 35193 5940 35429
rect 6176 35193 6261 35429
rect 6497 35193 6582 35429
rect 6818 35193 6903 35429
rect 7139 35193 7224 35429
rect 7460 35193 7545 35429
rect 7781 35193 7866 35429
rect 8102 35193 8187 35429
rect 8423 35193 8508 35429
rect 8744 35193 8829 35429
rect 9065 35193 9150 35429
rect 9386 35193 9471 35429
rect 9707 35193 9792 35429
rect 10028 35193 10113 35429
rect 10349 35193 10434 35429
rect 10670 35193 10755 35429
rect 10991 35193 11076 35429
rect 11312 35193 11397 35429
rect 11633 35193 11718 35429
rect 11954 35193 12038 35429
rect 12274 35193 12358 35429
rect 12594 35193 12678 35429
rect 12914 35193 12998 35429
rect 13234 35193 13318 35429
rect 13554 35193 13638 35429
rect 13874 35193 13958 35429
rect 14194 35193 14278 35429
rect 14514 35193 14598 35429
rect 14834 35193 14918 35429
rect 15154 35193 15238 35429
rect 15474 35193 15558 35429
rect 15794 35193 16000 35429
rect 0 35157 16000 35193
rect 6374 25521 10682 29830
rect 0 18972 16000 18997
rect 0 18736 162 18972
rect 398 18736 483 18972
rect 719 18736 804 18972
rect 1040 18736 1125 18972
rect 1361 18736 1446 18972
rect 1682 18736 1767 18972
rect 2003 18736 2088 18972
rect 2324 18736 2409 18972
rect 2645 18736 2730 18972
rect 2966 18736 3051 18972
rect 3287 18736 3372 18972
rect 3608 18736 3693 18972
rect 3929 18736 4014 18972
rect 4250 18736 4335 18972
rect 4571 18736 4656 18972
rect 4892 18736 4977 18972
rect 5213 18736 5298 18972
rect 5534 18736 5619 18972
rect 5855 18736 5940 18972
rect 6176 18736 6261 18972
rect 6497 18736 6582 18972
rect 6818 18736 6903 18972
rect 7139 18736 7224 18972
rect 7460 18736 7545 18972
rect 7781 18736 7866 18972
rect 8102 18736 8187 18972
rect 8423 18736 8508 18972
rect 8744 18736 8829 18972
rect 9065 18736 9150 18972
rect 9386 18736 9471 18972
rect 9707 18736 9792 18972
rect 10028 18736 10113 18972
rect 10349 18736 10434 18972
rect 10670 18736 10755 18972
rect 10991 18736 11076 18972
rect 11312 18736 11397 18972
rect 11633 18736 11718 18972
rect 11954 18736 12038 18972
rect 12274 18736 12358 18972
rect 12594 18736 12678 18972
rect 12914 18736 12998 18972
rect 13234 18736 13318 18972
rect 13554 18736 13638 18972
rect 13874 18736 13958 18972
rect 14194 18736 14278 18972
rect 14514 18736 14598 18972
rect 14834 18736 14918 18972
rect 15154 18736 15238 18972
rect 15474 18736 15558 18972
rect 15794 18736 16000 18972
rect 0 18636 16000 18736
rect 0 18400 162 18636
rect 398 18400 483 18636
rect 719 18400 804 18636
rect 1040 18400 1125 18636
rect 1361 18400 1446 18636
rect 1682 18400 1767 18636
rect 2003 18400 2088 18636
rect 2324 18400 2409 18636
rect 2645 18400 2730 18636
rect 2966 18400 3051 18636
rect 3287 18400 3372 18636
rect 3608 18400 3693 18636
rect 3929 18400 4014 18636
rect 4250 18400 4335 18636
rect 4571 18400 4656 18636
rect 4892 18400 4977 18636
rect 5213 18400 5298 18636
rect 5534 18400 5619 18636
rect 5855 18400 5940 18636
rect 6176 18400 6261 18636
rect 6497 18400 6582 18636
rect 6818 18400 6903 18636
rect 7139 18400 7224 18636
rect 7460 18400 7545 18636
rect 7781 18400 7866 18636
rect 8102 18400 8187 18636
rect 8423 18400 8508 18636
rect 8744 18400 8829 18636
rect 9065 18400 9150 18636
rect 9386 18400 9471 18636
rect 9707 18400 9792 18636
rect 10028 18400 10113 18636
rect 10349 18400 10434 18636
rect 10670 18400 10755 18636
rect 10991 18400 11076 18636
rect 11312 18400 11397 18636
rect 11633 18400 11718 18636
rect 11954 18400 12038 18636
rect 12274 18400 12358 18636
rect 12594 18400 12678 18636
rect 12914 18400 12998 18636
rect 13234 18400 13318 18636
rect 13554 18400 13638 18636
rect 13874 18400 13958 18636
rect 14194 18400 14278 18636
rect 14514 18400 14598 18636
rect 14834 18400 14918 18636
rect 15154 18400 15238 18636
rect 15474 18400 15558 18636
rect 15794 18400 16000 18636
rect 0 18300 16000 18400
rect 0 18064 162 18300
rect 398 18064 483 18300
rect 719 18064 804 18300
rect 1040 18064 1125 18300
rect 1361 18064 1446 18300
rect 1682 18064 1767 18300
rect 2003 18064 2088 18300
rect 2324 18064 2409 18300
rect 2645 18064 2730 18300
rect 2966 18064 3051 18300
rect 3287 18064 3372 18300
rect 3608 18064 3693 18300
rect 3929 18064 4014 18300
rect 4250 18064 4335 18300
rect 4571 18064 4656 18300
rect 4892 18064 4977 18300
rect 5213 18064 5298 18300
rect 5534 18064 5619 18300
rect 5855 18064 5940 18300
rect 6176 18064 6261 18300
rect 6497 18064 6582 18300
rect 6818 18064 6903 18300
rect 7139 18064 7224 18300
rect 7460 18064 7545 18300
rect 7781 18064 7866 18300
rect 8102 18064 8187 18300
rect 8423 18064 8508 18300
rect 8744 18064 8829 18300
rect 9065 18064 9150 18300
rect 9386 18064 9471 18300
rect 9707 18064 9792 18300
rect 10028 18064 10113 18300
rect 10349 18064 10434 18300
rect 10670 18064 10755 18300
rect 10991 18064 11076 18300
rect 11312 18064 11397 18300
rect 11633 18064 11718 18300
rect 11954 18064 12038 18300
rect 12274 18064 12358 18300
rect 12594 18064 12678 18300
rect 12914 18064 12998 18300
rect 13234 18064 13318 18300
rect 13554 18064 13638 18300
rect 13874 18064 13958 18300
rect 14194 18064 14278 18300
rect 14514 18064 14598 18300
rect 14834 18064 14918 18300
rect 15154 18064 15238 18300
rect 15474 18064 15558 18300
rect 15794 18064 16000 18300
rect 0 17964 16000 18064
rect 0 17728 162 17964
rect 398 17728 483 17964
rect 719 17728 804 17964
rect 1040 17728 1125 17964
rect 1361 17728 1446 17964
rect 1682 17728 1767 17964
rect 2003 17728 2088 17964
rect 2324 17728 2409 17964
rect 2645 17728 2730 17964
rect 2966 17728 3051 17964
rect 3287 17728 3372 17964
rect 3608 17728 3693 17964
rect 3929 17728 4014 17964
rect 4250 17728 4335 17964
rect 4571 17728 4656 17964
rect 4892 17728 4977 17964
rect 5213 17728 5298 17964
rect 5534 17728 5619 17964
rect 5855 17728 5940 17964
rect 6176 17728 6261 17964
rect 6497 17728 6582 17964
rect 6818 17728 6903 17964
rect 7139 17728 7224 17964
rect 7460 17728 7545 17964
rect 7781 17728 7866 17964
rect 8102 17728 8187 17964
rect 8423 17728 8508 17964
rect 8744 17728 8829 17964
rect 9065 17728 9150 17964
rect 9386 17728 9471 17964
rect 9707 17728 9792 17964
rect 10028 17728 10113 17964
rect 10349 17728 10434 17964
rect 10670 17728 10755 17964
rect 10991 17728 11076 17964
rect 11312 17728 11397 17964
rect 11633 17728 11718 17964
rect 11954 17728 12038 17964
rect 12274 17728 12358 17964
rect 12594 17728 12678 17964
rect 12914 17728 12998 17964
rect 13234 17728 13318 17964
rect 13554 17728 13638 17964
rect 13874 17728 13958 17964
rect 14194 17728 14278 17964
rect 14514 17728 14598 17964
rect 14834 17728 14918 17964
rect 15154 17728 15238 17964
rect 15474 17728 15558 17964
rect 15794 17728 16000 17964
rect 0 17628 16000 17728
rect 0 17392 162 17628
rect 398 17392 483 17628
rect 719 17392 804 17628
rect 1040 17392 1125 17628
rect 1361 17392 1446 17628
rect 1682 17392 1767 17628
rect 2003 17392 2088 17628
rect 2324 17392 2409 17628
rect 2645 17392 2730 17628
rect 2966 17392 3051 17628
rect 3287 17392 3372 17628
rect 3608 17392 3693 17628
rect 3929 17392 4014 17628
rect 4250 17392 4335 17628
rect 4571 17392 4656 17628
rect 4892 17392 4977 17628
rect 5213 17392 5298 17628
rect 5534 17392 5619 17628
rect 5855 17392 5940 17628
rect 6176 17392 6261 17628
rect 6497 17392 6582 17628
rect 6818 17392 6903 17628
rect 7139 17392 7224 17628
rect 7460 17392 7545 17628
rect 7781 17392 7866 17628
rect 8102 17392 8187 17628
rect 8423 17392 8508 17628
rect 8744 17392 8829 17628
rect 9065 17392 9150 17628
rect 9386 17392 9471 17628
rect 9707 17392 9792 17628
rect 10028 17392 10113 17628
rect 10349 17392 10434 17628
rect 10670 17392 10755 17628
rect 10991 17392 11076 17628
rect 11312 17392 11397 17628
rect 11633 17392 11718 17628
rect 11954 17392 12038 17628
rect 12274 17392 12358 17628
rect 12594 17392 12678 17628
rect 12914 17392 12998 17628
rect 13234 17392 13318 17628
rect 13554 17392 13638 17628
rect 13874 17392 13958 17628
rect 14194 17392 14278 17628
rect 14514 17392 14598 17628
rect 14834 17392 14918 17628
rect 15154 17392 15238 17628
rect 15474 17392 15558 17628
rect 15794 17392 16000 17628
rect 0 17292 16000 17392
rect 0 17056 162 17292
rect 398 17056 483 17292
rect 719 17056 804 17292
rect 1040 17056 1125 17292
rect 1361 17056 1446 17292
rect 1682 17056 1767 17292
rect 2003 17056 2088 17292
rect 2324 17056 2409 17292
rect 2645 17056 2730 17292
rect 2966 17056 3051 17292
rect 3287 17056 3372 17292
rect 3608 17056 3693 17292
rect 3929 17056 4014 17292
rect 4250 17056 4335 17292
rect 4571 17056 4656 17292
rect 4892 17056 4977 17292
rect 5213 17056 5298 17292
rect 5534 17056 5619 17292
rect 5855 17056 5940 17292
rect 6176 17056 6261 17292
rect 6497 17056 6582 17292
rect 6818 17056 6903 17292
rect 7139 17056 7224 17292
rect 7460 17056 7545 17292
rect 7781 17056 7866 17292
rect 8102 17056 8187 17292
rect 8423 17056 8508 17292
rect 8744 17056 8829 17292
rect 9065 17056 9150 17292
rect 9386 17056 9471 17292
rect 9707 17056 9792 17292
rect 10028 17056 10113 17292
rect 10349 17056 10434 17292
rect 10670 17056 10755 17292
rect 10991 17056 11076 17292
rect 11312 17056 11397 17292
rect 11633 17056 11718 17292
rect 11954 17056 12038 17292
rect 12274 17056 12358 17292
rect 12594 17056 12678 17292
rect 12914 17056 12998 17292
rect 13234 17056 13318 17292
rect 13554 17056 13638 17292
rect 13874 17056 13958 17292
rect 14194 17056 14278 17292
rect 14514 17056 14598 17292
rect 14834 17056 14918 17292
rect 15154 17056 15238 17292
rect 15474 17056 15558 17292
rect 15794 17056 16000 17292
rect 0 16956 16000 17056
rect 0 16720 162 16956
rect 398 16720 483 16956
rect 719 16720 804 16956
rect 1040 16720 1125 16956
rect 1361 16720 1446 16956
rect 1682 16720 1767 16956
rect 2003 16720 2088 16956
rect 2324 16720 2409 16956
rect 2645 16720 2730 16956
rect 2966 16720 3051 16956
rect 3287 16720 3372 16956
rect 3608 16720 3693 16956
rect 3929 16720 4014 16956
rect 4250 16720 4335 16956
rect 4571 16720 4656 16956
rect 4892 16720 4977 16956
rect 5213 16720 5298 16956
rect 5534 16720 5619 16956
rect 5855 16720 5940 16956
rect 6176 16720 6261 16956
rect 6497 16720 6582 16956
rect 6818 16720 6903 16956
rect 7139 16720 7224 16956
rect 7460 16720 7545 16956
rect 7781 16720 7866 16956
rect 8102 16720 8187 16956
rect 8423 16720 8508 16956
rect 8744 16720 8829 16956
rect 9065 16720 9150 16956
rect 9386 16720 9471 16956
rect 9707 16720 9792 16956
rect 10028 16720 10113 16956
rect 10349 16720 10434 16956
rect 10670 16720 10755 16956
rect 10991 16720 11076 16956
rect 11312 16720 11397 16956
rect 11633 16720 11718 16956
rect 11954 16720 12038 16956
rect 12274 16720 12358 16956
rect 12594 16720 12678 16956
rect 12914 16720 12998 16956
rect 13234 16720 13318 16956
rect 13554 16720 13638 16956
rect 13874 16720 13958 16956
rect 14194 16720 14278 16956
rect 14514 16720 14598 16956
rect 14834 16720 14918 16956
rect 15154 16720 15238 16956
rect 15474 16720 15558 16956
rect 15794 16720 16000 16956
rect 0 16620 16000 16720
rect 0 16384 162 16620
rect 398 16384 483 16620
rect 719 16384 804 16620
rect 1040 16384 1125 16620
rect 1361 16384 1446 16620
rect 1682 16384 1767 16620
rect 2003 16384 2088 16620
rect 2324 16384 2409 16620
rect 2645 16384 2730 16620
rect 2966 16384 3051 16620
rect 3287 16384 3372 16620
rect 3608 16384 3693 16620
rect 3929 16384 4014 16620
rect 4250 16384 4335 16620
rect 4571 16384 4656 16620
rect 4892 16384 4977 16620
rect 5213 16384 5298 16620
rect 5534 16384 5619 16620
rect 5855 16384 5940 16620
rect 6176 16384 6261 16620
rect 6497 16384 6582 16620
rect 6818 16384 6903 16620
rect 7139 16384 7224 16620
rect 7460 16384 7545 16620
rect 7781 16384 7866 16620
rect 8102 16384 8187 16620
rect 8423 16384 8508 16620
rect 8744 16384 8829 16620
rect 9065 16384 9150 16620
rect 9386 16384 9471 16620
rect 9707 16384 9792 16620
rect 10028 16384 10113 16620
rect 10349 16384 10434 16620
rect 10670 16384 10755 16620
rect 10991 16384 11076 16620
rect 11312 16384 11397 16620
rect 11633 16384 11718 16620
rect 11954 16384 12038 16620
rect 12274 16384 12358 16620
rect 12594 16384 12678 16620
rect 12914 16384 12998 16620
rect 13234 16384 13318 16620
rect 13554 16384 13638 16620
rect 13874 16384 13958 16620
rect 14194 16384 14278 16620
rect 14514 16384 14598 16620
rect 14834 16384 14918 16620
rect 15154 16384 15238 16620
rect 15474 16384 15558 16620
rect 15794 16384 16000 16620
rect 0 16284 16000 16384
rect 0 16048 162 16284
rect 398 16048 483 16284
rect 719 16048 804 16284
rect 1040 16048 1125 16284
rect 1361 16048 1446 16284
rect 1682 16048 1767 16284
rect 2003 16048 2088 16284
rect 2324 16048 2409 16284
rect 2645 16048 2730 16284
rect 2966 16048 3051 16284
rect 3287 16048 3372 16284
rect 3608 16048 3693 16284
rect 3929 16048 4014 16284
rect 4250 16048 4335 16284
rect 4571 16048 4656 16284
rect 4892 16048 4977 16284
rect 5213 16048 5298 16284
rect 5534 16048 5619 16284
rect 5855 16048 5940 16284
rect 6176 16048 6261 16284
rect 6497 16048 6582 16284
rect 6818 16048 6903 16284
rect 7139 16048 7224 16284
rect 7460 16048 7545 16284
rect 7781 16048 7866 16284
rect 8102 16048 8187 16284
rect 8423 16048 8508 16284
rect 8744 16048 8829 16284
rect 9065 16048 9150 16284
rect 9386 16048 9471 16284
rect 9707 16048 9792 16284
rect 10028 16048 10113 16284
rect 10349 16048 10434 16284
rect 10670 16048 10755 16284
rect 10991 16048 11076 16284
rect 11312 16048 11397 16284
rect 11633 16048 11718 16284
rect 11954 16048 12038 16284
rect 12274 16048 12358 16284
rect 12594 16048 12678 16284
rect 12914 16048 12998 16284
rect 13234 16048 13318 16284
rect 13554 16048 13638 16284
rect 13874 16048 13958 16284
rect 14194 16048 14278 16284
rect 14514 16048 14598 16284
rect 14834 16048 14918 16284
rect 15154 16048 15238 16284
rect 15474 16048 15558 16284
rect 15794 16048 16000 16284
rect 0 15948 16000 16048
rect 0 15712 162 15948
rect 398 15712 483 15948
rect 719 15712 804 15948
rect 1040 15712 1125 15948
rect 1361 15712 1446 15948
rect 1682 15712 1767 15948
rect 2003 15712 2088 15948
rect 2324 15712 2409 15948
rect 2645 15712 2730 15948
rect 2966 15712 3051 15948
rect 3287 15712 3372 15948
rect 3608 15712 3693 15948
rect 3929 15712 4014 15948
rect 4250 15712 4335 15948
rect 4571 15712 4656 15948
rect 4892 15712 4977 15948
rect 5213 15712 5298 15948
rect 5534 15712 5619 15948
rect 5855 15712 5940 15948
rect 6176 15712 6261 15948
rect 6497 15712 6582 15948
rect 6818 15712 6903 15948
rect 7139 15712 7224 15948
rect 7460 15712 7545 15948
rect 7781 15712 7866 15948
rect 8102 15712 8187 15948
rect 8423 15712 8508 15948
rect 8744 15712 8829 15948
rect 9065 15712 9150 15948
rect 9386 15712 9471 15948
rect 9707 15712 9792 15948
rect 10028 15712 10113 15948
rect 10349 15712 10434 15948
rect 10670 15712 10755 15948
rect 10991 15712 11076 15948
rect 11312 15712 11397 15948
rect 11633 15712 11718 15948
rect 11954 15712 12038 15948
rect 12274 15712 12358 15948
rect 12594 15712 12678 15948
rect 12914 15712 12998 15948
rect 13234 15712 13318 15948
rect 13554 15712 13638 15948
rect 13874 15712 13958 15948
rect 14194 15712 14278 15948
rect 14514 15712 14598 15948
rect 14834 15712 14918 15948
rect 15154 15712 15238 15948
rect 15474 15712 15558 15948
rect 15794 15712 16000 15948
rect 0 15612 16000 15712
rect 0 15376 162 15612
rect 398 15376 483 15612
rect 719 15376 804 15612
rect 1040 15376 1125 15612
rect 1361 15376 1446 15612
rect 1682 15376 1767 15612
rect 2003 15376 2088 15612
rect 2324 15376 2409 15612
rect 2645 15376 2730 15612
rect 2966 15376 3051 15612
rect 3287 15376 3372 15612
rect 3608 15376 3693 15612
rect 3929 15376 4014 15612
rect 4250 15376 4335 15612
rect 4571 15376 4656 15612
rect 4892 15376 4977 15612
rect 5213 15376 5298 15612
rect 5534 15376 5619 15612
rect 5855 15376 5940 15612
rect 6176 15376 6261 15612
rect 6497 15376 6582 15612
rect 6818 15376 6903 15612
rect 7139 15376 7224 15612
rect 7460 15376 7545 15612
rect 7781 15376 7866 15612
rect 8102 15376 8187 15612
rect 8423 15376 8508 15612
rect 8744 15376 8829 15612
rect 9065 15376 9150 15612
rect 9386 15376 9471 15612
rect 9707 15376 9792 15612
rect 10028 15376 10113 15612
rect 10349 15376 10434 15612
rect 10670 15376 10755 15612
rect 10991 15376 11076 15612
rect 11312 15376 11397 15612
rect 11633 15376 11718 15612
rect 11954 15376 12038 15612
rect 12274 15376 12358 15612
rect 12594 15376 12678 15612
rect 12914 15376 12998 15612
rect 13234 15376 13318 15612
rect 13554 15376 13638 15612
rect 13874 15376 13958 15612
rect 14194 15376 14278 15612
rect 14514 15376 14598 15612
rect 14834 15376 14918 15612
rect 15154 15376 15238 15612
rect 15474 15376 15558 15612
rect 15794 15376 16000 15612
rect 0 15276 16000 15376
rect 0 15040 162 15276
rect 398 15040 483 15276
rect 719 15040 804 15276
rect 1040 15040 1125 15276
rect 1361 15040 1446 15276
rect 1682 15040 1767 15276
rect 2003 15040 2088 15276
rect 2324 15040 2409 15276
rect 2645 15040 2730 15276
rect 2966 15040 3051 15276
rect 3287 15040 3372 15276
rect 3608 15040 3693 15276
rect 3929 15040 4014 15276
rect 4250 15040 4335 15276
rect 4571 15040 4656 15276
rect 4892 15040 4977 15276
rect 5213 15040 5298 15276
rect 5534 15040 5619 15276
rect 5855 15040 5940 15276
rect 6176 15040 6261 15276
rect 6497 15040 6582 15276
rect 6818 15040 6903 15276
rect 7139 15040 7224 15276
rect 7460 15040 7545 15276
rect 7781 15040 7866 15276
rect 8102 15040 8187 15276
rect 8423 15040 8508 15276
rect 8744 15040 8829 15276
rect 9065 15040 9150 15276
rect 9386 15040 9471 15276
rect 9707 15040 9792 15276
rect 10028 15040 10113 15276
rect 10349 15040 10434 15276
rect 10670 15040 10755 15276
rect 10991 15040 11076 15276
rect 11312 15040 11397 15276
rect 11633 15040 11718 15276
rect 11954 15040 12038 15276
rect 12274 15040 12358 15276
rect 12594 15040 12678 15276
rect 12914 15040 12998 15276
rect 13234 15040 13318 15276
rect 13554 15040 13638 15276
rect 13874 15040 13958 15276
rect 14194 15040 14278 15276
rect 14514 15040 14598 15276
rect 14834 15040 14918 15276
rect 15154 15040 15238 15276
rect 15474 15040 15558 15276
rect 15794 15040 16000 15276
rect 0 14940 16000 15040
rect 0 14704 162 14940
rect 398 14704 483 14940
rect 719 14704 804 14940
rect 1040 14704 1125 14940
rect 1361 14704 1446 14940
rect 1682 14704 1767 14940
rect 2003 14704 2088 14940
rect 2324 14704 2409 14940
rect 2645 14704 2730 14940
rect 2966 14704 3051 14940
rect 3287 14704 3372 14940
rect 3608 14704 3693 14940
rect 3929 14704 4014 14940
rect 4250 14704 4335 14940
rect 4571 14704 4656 14940
rect 4892 14704 4977 14940
rect 5213 14704 5298 14940
rect 5534 14704 5619 14940
rect 5855 14704 5940 14940
rect 6176 14704 6261 14940
rect 6497 14704 6582 14940
rect 6818 14704 6903 14940
rect 7139 14704 7224 14940
rect 7460 14704 7545 14940
rect 7781 14704 7866 14940
rect 8102 14704 8187 14940
rect 8423 14704 8508 14940
rect 8744 14704 8829 14940
rect 9065 14704 9150 14940
rect 9386 14704 9471 14940
rect 9707 14704 9792 14940
rect 10028 14704 10113 14940
rect 10349 14704 10434 14940
rect 10670 14704 10755 14940
rect 10991 14704 11076 14940
rect 11312 14704 11397 14940
rect 11633 14704 11718 14940
rect 11954 14704 12038 14940
rect 12274 14704 12358 14940
rect 12594 14704 12678 14940
rect 12914 14704 12998 14940
rect 13234 14704 13318 14940
rect 13554 14704 13638 14940
rect 13874 14704 13958 14940
rect 14194 14704 14278 14940
rect 14514 14704 14598 14940
rect 14834 14704 14918 14940
rect 15154 14704 15238 14940
rect 15474 14704 15558 14940
rect 15794 14704 16000 14940
rect 0 14604 16000 14704
rect 0 14368 162 14604
rect 398 14368 483 14604
rect 719 14368 804 14604
rect 1040 14368 1125 14604
rect 1361 14368 1446 14604
rect 1682 14368 1767 14604
rect 2003 14368 2088 14604
rect 2324 14368 2409 14604
rect 2645 14368 2730 14604
rect 2966 14368 3051 14604
rect 3287 14368 3372 14604
rect 3608 14368 3693 14604
rect 3929 14368 4014 14604
rect 4250 14368 4335 14604
rect 4571 14368 4656 14604
rect 4892 14368 4977 14604
rect 5213 14368 5298 14604
rect 5534 14368 5619 14604
rect 5855 14368 5940 14604
rect 6176 14368 6261 14604
rect 6497 14368 6582 14604
rect 6818 14368 6903 14604
rect 7139 14368 7224 14604
rect 7460 14368 7545 14604
rect 7781 14368 7866 14604
rect 8102 14368 8187 14604
rect 8423 14368 8508 14604
rect 8744 14368 8829 14604
rect 9065 14368 9150 14604
rect 9386 14368 9471 14604
rect 9707 14368 9792 14604
rect 10028 14368 10113 14604
rect 10349 14368 10434 14604
rect 10670 14368 10755 14604
rect 10991 14368 11076 14604
rect 11312 14368 11397 14604
rect 11633 14368 11718 14604
rect 11954 14368 12038 14604
rect 12274 14368 12358 14604
rect 12594 14368 12678 14604
rect 12914 14368 12998 14604
rect 13234 14368 13318 14604
rect 13554 14368 13638 14604
rect 13874 14368 13958 14604
rect 14194 14368 14278 14604
rect 14514 14368 14598 14604
rect 14834 14368 14918 14604
rect 15154 14368 15238 14604
rect 15474 14368 15558 14604
rect 15794 14368 16000 14604
rect 0 14268 16000 14368
rect 0 14032 162 14268
rect 398 14032 483 14268
rect 719 14032 804 14268
rect 1040 14032 1125 14268
rect 1361 14032 1446 14268
rect 1682 14032 1767 14268
rect 2003 14032 2088 14268
rect 2324 14032 2409 14268
rect 2645 14032 2730 14268
rect 2966 14032 3051 14268
rect 3287 14032 3372 14268
rect 3608 14032 3693 14268
rect 3929 14032 4014 14268
rect 4250 14032 4335 14268
rect 4571 14032 4656 14268
rect 4892 14032 4977 14268
rect 5213 14032 5298 14268
rect 5534 14032 5619 14268
rect 5855 14032 5940 14268
rect 6176 14032 6261 14268
rect 6497 14032 6582 14268
rect 6818 14032 6903 14268
rect 7139 14032 7224 14268
rect 7460 14032 7545 14268
rect 7781 14032 7866 14268
rect 8102 14032 8187 14268
rect 8423 14032 8508 14268
rect 8744 14032 8829 14268
rect 9065 14032 9150 14268
rect 9386 14032 9471 14268
rect 9707 14032 9792 14268
rect 10028 14032 10113 14268
rect 10349 14032 10434 14268
rect 10670 14032 10755 14268
rect 10991 14032 11076 14268
rect 11312 14032 11397 14268
rect 11633 14032 11718 14268
rect 11954 14032 12038 14268
rect 12274 14032 12358 14268
rect 12594 14032 12678 14268
rect 12914 14032 12998 14268
rect 13234 14032 13318 14268
rect 13554 14032 13638 14268
rect 13874 14032 13958 14268
rect 14194 14032 14278 14268
rect 14514 14032 14598 14268
rect 14834 14032 14918 14268
rect 15154 14032 15238 14268
rect 15474 14032 15558 14268
rect 15794 14032 16000 14268
rect 0 14007 16000 14032
rect 0 13663 16000 13687
rect 0 13427 162 13663
rect 398 13427 483 13663
rect 719 13427 804 13663
rect 1040 13427 1125 13663
rect 1361 13427 1446 13663
rect 1682 13427 1767 13663
rect 2003 13427 2088 13663
rect 2324 13427 2409 13663
rect 2645 13427 2730 13663
rect 2966 13427 3051 13663
rect 3287 13427 3372 13663
rect 3608 13427 3693 13663
rect 3929 13427 4014 13663
rect 4250 13427 4335 13663
rect 4571 13427 4656 13663
rect 4892 13427 4977 13663
rect 5213 13427 5298 13663
rect 5534 13427 5619 13663
rect 5855 13427 5940 13663
rect 6176 13427 6261 13663
rect 6497 13427 6582 13663
rect 6818 13427 6903 13663
rect 7139 13427 7224 13663
rect 7460 13427 7545 13663
rect 7781 13427 7866 13663
rect 8102 13427 8187 13663
rect 8423 13427 8508 13663
rect 8744 13427 8829 13663
rect 9065 13427 9150 13663
rect 9386 13427 9471 13663
rect 9707 13427 9792 13663
rect 10028 13427 10113 13663
rect 10349 13427 10434 13663
rect 10670 13427 10755 13663
rect 10991 13427 11076 13663
rect 11312 13427 11397 13663
rect 11633 13427 11718 13663
rect 11954 13427 12038 13663
rect 12274 13427 12358 13663
rect 12594 13427 12678 13663
rect 12914 13427 12998 13663
rect 13234 13427 13318 13663
rect 13554 13427 13638 13663
rect 13874 13427 13958 13663
rect 14194 13427 14278 13663
rect 14514 13427 14598 13663
rect 14834 13427 14918 13663
rect 15154 13427 15238 13663
rect 15474 13427 15558 13663
rect 15794 13427 16000 13663
rect 0 13097 16000 13427
rect 0 12861 162 13097
rect 398 12861 483 13097
rect 719 12861 804 13097
rect 1040 12861 1125 13097
rect 1361 12861 1446 13097
rect 1682 12861 1767 13097
rect 2003 12861 2088 13097
rect 2324 12861 2409 13097
rect 2645 12861 2730 13097
rect 2966 12861 3051 13097
rect 3287 12861 3372 13097
rect 3608 12861 3693 13097
rect 3929 12861 4014 13097
rect 4250 12861 4335 13097
rect 4571 12861 4656 13097
rect 4892 12861 4977 13097
rect 5213 12861 5298 13097
rect 5534 12861 5619 13097
rect 5855 12861 5940 13097
rect 6176 12861 6261 13097
rect 6497 12861 6582 13097
rect 6818 12861 6903 13097
rect 7139 12861 7224 13097
rect 7460 12861 7545 13097
rect 7781 12861 7866 13097
rect 8102 12861 8187 13097
rect 8423 12861 8508 13097
rect 8744 12861 8829 13097
rect 9065 12861 9150 13097
rect 9386 12861 9471 13097
rect 9707 12861 9792 13097
rect 10028 12861 10113 13097
rect 10349 12861 10434 13097
rect 10670 12861 10755 13097
rect 10991 12861 11076 13097
rect 11312 12861 11397 13097
rect 11633 12861 11718 13097
rect 11954 12861 12038 13097
rect 12274 12861 12358 13097
rect 12594 12861 12678 13097
rect 12914 12861 12998 13097
rect 13234 12861 13318 13097
rect 13554 12861 13638 13097
rect 13874 12861 13958 13097
rect 14194 12861 14278 13097
rect 14514 12861 14598 13097
rect 14834 12861 14918 13097
rect 15154 12861 15238 13097
rect 15474 12861 15558 13097
rect 15794 12861 16000 13097
rect 0 12837 16000 12861
rect 0 12493 16000 12517
rect 0 12257 162 12493
rect 398 12257 483 12493
rect 719 12257 804 12493
rect 1040 12257 1125 12493
rect 1361 12257 1446 12493
rect 1682 12257 1767 12493
rect 2003 12257 2088 12493
rect 2324 12257 2409 12493
rect 2645 12257 2730 12493
rect 2966 12257 3051 12493
rect 3287 12257 3372 12493
rect 3608 12257 3693 12493
rect 3929 12257 4014 12493
rect 4250 12257 4335 12493
rect 4571 12257 4656 12493
rect 4892 12257 4977 12493
rect 5213 12257 5298 12493
rect 5534 12257 5619 12493
rect 5855 12257 5940 12493
rect 6176 12257 6261 12493
rect 6497 12257 6582 12493
rect 6818 12257 6903 12493
rect 7139 12257 7224 12493
rect 7460 12257 7545 12493
rect 7781 12257 7866 12493
rect 8102 12257 8187 12493
rect 8423 12257 8508 12493
rect 8744 12257 8829 12493
rect 9065 12257 9150 12493
rect 9386 12257 9471 12493
rect 9707 12257 9792 12493
rect 10028 12257 10113 12493
rect 10349 12257 10434 12493
rect 10670 12257 10755 12493
rect 10991 12257 11076 12493
rect 11312 12257 11397 12493
rect 11633 12257 11718 12493
rect 11954 12257 12039 12493
rect 12275 12257 12359 12493
rect 12595 12257 12679 12493
rect 12915 12257 12999 12493
rect 13235 12257 13319 12493
rect 13555 12257 13639 12493
rect 13875 12257 13959 12493
rect 14195 12257 14279 12493
rect 14515 12257 14599 12493
rect 14835 12257 14919 12493
rect 15155 12257 15239 12493
rect 15475 12257 15559 12493
rect 15795 12257 16000 12493
rect 0 11927 16000 12257
rect 0 11691 162 11927
rect 398 11691 483 11927
rect 719 11691 804 11927
rect 1040 11691 1125 11927
rect 1361 11691 1446 11927
rect 1682 11691 1767 11927
rect 2003 11691 2088 11927
rect 2324 11691 2409 11927
rect 2645 11691 2730 11927
rect 2966 11691 3051 11927
rect 3287 11691 3372 11927
rect 3608 11691 3693 11927
rect 3929 11691 4014 11927
rect 4250 11691 4335 11927
rect 4571 11691 4656 11927
rect 4892 11691 4977 11927
rect 5213 11691 5298 11927
rect 5534 11691 5619 11927
rect 5855 11691 5940 11927
rect 6176 11691 6261 11927
rect 6497 11691 6582 11927
rect 6818 11691 6903 11927
rect 7139 11691 7224 11927
rect 7460 11691 7545 11927
rect 7781 11691 7866 11927
rect 8102 11691 8187 11927
rect 8423 11691 8508 11927
rect 8744 11691 8829 11927
rect 9065 11691 9150 11927
rect 9386 11691 9471 11927
rect 9707 11691 9792 11927
rect 10028 11691 10113 11927
rect 10349 11691 10434 11927
rect 10670 11691 10755 11927
rect 10991 11691 11076 11927
rect 11312 11691 11397 11927
rect 11633 11691 11718 11927
rect 11954 11691 12039 11927
rect 12275 11691 12359 11927
rect 12595 11691 12679 11927
rect 12915 11691 12999 11927
rect 13235 11691 13319 11927
rect 13555 11691 13639 11927
rect 13875 11691 13959 11927
rect 14195 11691 14279 11927
rect 14515 11691 14599 11927
rect 14835 11691 14919 11927
rect 15155 11691 15239 11927
rect 15475 11691 15559 11927
rect 15795 11691 16000 11927
rect 0 11667 16000 11691
rect 0 10565 16000 11347
rect 0 10329 162 10565
rect 398 10329 483 10565
rect 719 10329 804 10565
rect 1040 10329 1125 10565
rect 1361 10329 1446 10565
rect 1682 10329 1767 10565
rect 2003 10329 2088 10565
rect 2324 10329 2409 10565
rect 2645 10329 2730 10565
rect 2966 10329 3051 10565
rect 3287 10329 3372 10565
rect 3608 10329 3693 10565
rect 3929 10329 4014 10565
rect 4250 10329 4335 10565
rect 4571 10329 4656 10565
rect 4892 10329 4977 10565
rect 5213 10329 5298 10565
rect 5534 10329 5619 10565
rect 5855 10329 5940 10565
rect 6176 10329 6261 10565
rect 6497 10329 6582 10565
rect 6818 10329 6903 10565
rect 7139 10329 7224 10565
rect 7460 10329 7545 10565
rect 7781 10329 7866 10565
rect 8102 10329 8187 10565
rect 8423 10329 8508 10565
rect 8744 10329 8829 10565
rect 9065 10329 9150 10565
rect 9386 10329 9471 10565
rect 9707 10329 9792 10565
rect 10028 10329 10113 10565
rect 10349 10329 10434 10565
rect 10670 10329 10755 10565
rect 10991 10329 11076 10565
rect 11312 10329 11397 10565
rect 11633 10329 11718 10565
rect 11954 10329 12038 10565
rect 12274 10329 12358 10565
rect 12594 10329 12678 10565
rect 12914 10329 12998 10565
rect 13234 10329 13318 10565
rect 13554 10329 13638 10565
rect 13874 10329 13958 10565
rect 14194 10329 14278 10565
rect 14514 10329 14598 10565
rect 14834 10329 14918 10565
rect 15154 10329 15238 10565
rect 15474 10329 15558 10565
rect 15794 10329 16000 10565
rect 0 9547 16000 10329
rect 0 9203 16000 9227
rect 0 8967 162 9203
rect 398 8967 483 9203
rect 719 8967 804 9203
rect 1040 8967 1125 9203
rect 1361 8967 1446 9203
rect 1682 8967 1767 9203
rect 2003 8967 2088 9203
rect 2324 8967 2409 9203
rect 2645 8967 2730 9203
rect 2966 8967 3051 9203
rect 3287 8967 3372 9203
rect 3608 8967 3693 9203
rect 3929 8967 4014 9203
rect 4250 8967 4335 9203
rect 4571 8967 4656 9203
rect 4892 8967 4977 9203
rect 5213 8967 5298 9203
rect 5534 8967 5619 9203
rect 5855 8967 5940 9203
rect 6176 8967 6261 9203
rect 6497 8967 6582 9203
rect 6818 8967 6903 9203
rect 7139 8967 7224 9203
rect 7460 8967 7545 9203
rect 7781 8967 7866 9203
rect 8102 8967 8187 9203
rect 8423 8967 8508 9203
rect 8744 8967 8829 9203
rect 9065 8967 9150 9203
rect 9386 8967 9471 9203
rect 9707 8967 9792 9203
rect 10028 8967 10113 9203
rect 10349 8967 10434 9203
rect 10670 8967 10755 9203
rect 10991 8967 11076 9203
rect 11312 8967 11397 9203
rect 11633 8967 11717 9203
rect 11953 8967 12037 9203
rect 12273 8967 12357 9203
rect 12593 8967 12677 9203
rect 12913 8967 12997 9203
rect 13233 8967 13317 9203
rect 13553 8967 13637 9203
rect 13873 8967 13957 9203
rect 14193 8967 14277 9203
rect 14513 8967 14597 9203
rect 14833 8967 14917 9203
rect 15153 8967 15237 9203
rect 15473 8967 15557 9203
rect 15793 8967 16000 9203
rect 0 8597 16000 8967
rect 0 8361 162 8597
rect 398 8361 483 8597
rect 719 8361 804 8597
rect 1040 8361 1125 8597
rect 1361 8361 1446 8597
rect 1682 8361 1767 8597
rect 2003 8361 2088 8597
rect 2324 8361 2409 8597
rect 2645 8361 2730 8597
rect 2966 8361 3051 8597
rect 3287 8361 3372 8597
rect 3608 8361 3693 8597
rect 3929 8361 4014 8597
rect 4250 8361 4335 8597
rect 4571 8361 4656 8597
rect 4892 8361 4977 8597
rect 5213 8361 5298 8597
rect 5534 8361 5619 8597
rect 5855 8361 5940 8597
rect 6176 8361 6261 8597
rect 6497 8361 6582 8597
rect 6818 8361 6903 8597
rect 7139 8361 7224 8597
rect 7460 8361 7545 8597
rect 7781 8361 7866 8597
rect 8102 8361 8187 8597
rect 8423 8361 8508 8597
rect 8744 8361 8829 8597
rect 9065 8361 9150 8597
rect 9386 8361 9471 8597
rect 9707 8361 9792 8597
rect 10028 8361 10113 8597
rect 10349 8361 10434 8597
rect 10670 8361 10755 8597
rect 10991 8361 11076 8597
rect 11312 8361 11397 8597
rect 11633 8361 11717 8597
rect 11953 8361 12037 8597
rect 12273 8361 12357 8597
rect 12593 8361 12677 8597
rect 12913 8361 12997 8597
rect 13233 8361 13317 8597
rect 13553 8361 13637 8597
rect 13873 8361 13957 8597
rect 14193 8361 14277 8597
rect 14513 8361 14597 8597
rect 14833 8361 14917 8597
rect 15153 8361 15237 8597
rect 15473 8361 15557 8597
rect 15793 8361 16000 8597
rect 0 8337 16000 8361
rect 0 7993 16000 8017
rect 0 7757 162 7993
rect 398 7757 483 7993
rect 719 7757 804 7993
rect 1040 7757 1125 7993
rect 1361 7757 1446 7993
rect 1682 7757 1767 7993
rect 2003 7757 2088 7993
rect 2324 7757 2409 7993
rect 2645 7757 2730 7993
rect 2966 7757 3051 7993
rect 3287 7757 3372 7993
rect 3608 7757 3693 7993
rect 3929 7757 4014 7993
rect 4250 7757 4335 7993
rect 4571 7757 4656 7993
rect 4892 7757 4977 7993
rect 5213 7757 5298 7993
rect 5534 7757 5619 7993
rect 5855 7757 5940 7993
rect 6176 7757 6261 7993
rect 6497 7757 6582 7993
rect 6818 7757 6903 7993
rect 7139 7757 7224 7993
rect 7460 7757 7545 7993
rect 7781 7757 7866 7993
rect 8102 7757 8187 7993
rect 8423 7757 8508 7993
rect 8744 7757 8829 7993
rect 9065 7757 9150 7993
rect 9386 7757 9471 7993
rect 9707 7757 9792 7993
rect 10028 7757 10113 7993
rect 10349 7757 10434 7993
rect 10670 7757 10755 7993
rect 10991 7757 11076 7993
rect 11312 7757 11397 7993
rect 11633 7757 11718 7993
rect 11954 7757 12039 7993
rect 12275 7757 12359 7993
rect 12595 7757 12679 7993
rect 12915 7757 12999 7993
rect 13235 7757 13319 7993
rect 13555 7757 13639 7993
rect 13875 7757 13959 7993
rect 14195 7757 14279 7993
rect 14515 7757 14599 7993
rect 14835 7757 14919 7993
rect 15155 7757 15239 7993
rect 15475 7757 15559 7993
rect 15795 7757 16000 7993
rect 0 7627 16000 7757
rect 0 7391 162 7627
rect 398 7391 483 7627
rect 719 7391 804 7627
rect 1040 7391 1125 7627
rect 1361 7391 1446 7627
rect 1682 7391 1767 7627
rect 2003 7391 2088 7627
rect 2324 7391 2409 7627
rect 2645 7391 2730 7627
rect 2966 7391 3051 7627
rect 3287 7391 3372 7627
rect 3608 7391 3693 7627
rect 3929 7391 4014 7627
rect 4250 7391 4335 7627
rect 4571 7391 4656 7627
rect 4892 7391 4977 7627
rect 5213 7391 5298 7627
rect 5534 7391 5619 7627
rect 5855 7391 5940 7627
rect 6176 7391 6261 7627
rect 6497 7391 6582 7627
rect 6818 7391 6903 7627
rect 7139 7391 7224 7627
rect 7460 7391 7545 7627
rect 7781 7391 7866 7627
rect 8102 7391 8187 7627
rect 8423 7391 8508 7627
rect 8744 7391 8829 7627
rect 9065 7391 9150 7627
rect 9386 7391 9471 7627
rect 9707 7391 9792 7627
rect 10028 7391 10113 7627
rect 10349 7391 10434 7627
rect 10670 7391 10755 7627
rect 10991 7391 11076 7627
rect 11312 7391 11397 7627
rect 11633 7391 11718 7627
rect 11954 7391 12039 7627
rect 12275 7391 12359 7627
rect 12595 7391 12679 7627
rect 12915 7391 12999 7627
rect 13235 7391 13319 7627
rect 13555 7391 13639 7627
rect 13875 7391 13959 7627
rect 14195 7391 14279 7627
rect 14515 7391 14599 7627
rect 14835 7391 14919 7627
rect 15155 7391 15239 7627
rect 15475 7391 15559 7627
rect 15795 7391 16000 7627
rect 0 7367 16000 7391
rect 0 7023 16000 7047
rect 0 6787 162 7023
rect 398 6787 483 7023
rect 719 6787 804 7023
rect 1040 6787 1125 7023
rect 1361 6787 1446 7023
rect 1682 6787 1767 7023
rect 2003 6787 2088 7023
rect 2324 6787 2409 7023
rect 2645 6787 2730 7023
rect 2966 6787 3051 7023
rect 3287 6787 3372 7023
rect 3608 6787 3693 7023
rect 3929 6787 4014 7023
rect 4250 6787 4335 7023
rect 4571 6787 4656 7023
rect 4892 6787 4977 7023
rect 5213 6787 5298 7023
rect 5534 6787 5619 7023
rect 5855 6787 5940 7023
rect 6176 6787 6261 7023
rect 6497 6787 6582 7023
rect 6818 6787 6903 7023
rect 7139 6787 7224 7023
rect 7460 6787 7545 7023
rect 7781 6787 7866 7023
rect 8102 6787 8187 7023
rect 8423 6787 8508 7023
rect 8744 6787 8829 7023
rect 9065 6787 9150 7023
rect 9386 6787 9471 7023
rect 9707 6787 9792 7023
rect 10028 6787 10113 7023
rect 10349 6787 10434 7023
rect 10670 6787 10755 7023
rect 10991 6787 11076 7023
rect 11312 6787 11397 7023
rect 11633 6787 11718 7023
rect 11954 6787 12038 7023
rect 12274 6787 12358 7023
rect 12594 6787 12678 7023
rect 12914 6787 12998 7023
rect 13234 6787 13318 7023
rect 13554 6787 13638 7023
rect 13874 6787 13958 7023
rect 14194 6787 14278 7023
rect 14514 6787 14598 7023
rect 14834 6787 14918 7023
rect 15154 6787 15238 7023
rect 15474 6787 15558 7023
rect 15794 6787 16000 7023
rect 0 6657 16000 6787
rect 0 6421 162 6657
rect 398 6421 483 6657
rect 719 6421 804 6657
rect 1040 6421 1125 6657
rect 1361 6421 1446 6657
rect 1682 6421 1767 6657
rect 2003 6421 2088 6657
rect 2324 6421 2409 6657
rect 2645 6421 2730 6657
rect 2966 6421 3051 6657
rect 3287 6421 3372 6657
rect 3608 6421 3693 6657
rect 3929 6421 4014 6657
rect 4250 6421 4335 6657
rect 4571 6421 4656 6657
rect 4892 6421 4977 6657
rect 5213 6421 5298 6657
rect 5534 6421 5619 6657
rect 5855 6421 5940 6657
rect 6176 6421 6261 6657
rect 6497 6421 6582 6657
rect 6818 6421 6903 6657
rect 7139 6421 7224 6657
rect 7460 6421 7545 6657
rect 7781 6421 7866 6657
rect 8102 6421 8187 6657
rect 8423 6421 8508 6657
rect 8744 6421 8829 6657
rect 9065 6421 9150 6657
rect 9386 6421 9471 6657
rect 9707 6421 9792 6657
rect 10028 6421 10113 6657
rect 10349 6421 10434 6657
rect 10670 6421 10755 6657
rect 10991 6421 11076 6657
rect 11312 6421 11397 6657
rect 11633 6421 11718 6657
rect 11954 6421 12038 6657
rect 12274 6421 12358 6657
rect 12594 6421 12678 6657
rect 12914 6421 12998 6657
rect 13234 6421 13318 6657
rect 13554 6421 13638 6657
rect 13874 6421 13958 6657
rect 14194 6421 14278 6657
rect 14514 6421 14598 6657
rect 14834 6421 14918 6657
rect 15154 6421 15238 6657
rect 15474 6421 15558 6657
rect 15794 6421 16000 6657
rect 0 6397 16000 6421
rect 0 6053 16000 6077
rect 0 5817 161 6053
rect 397 5817 482 6053
rect 718 5817 803 6053
rect 1039 5817 1124 6053
rect 1360 5817 1445 6053
rect 1681 5817 1766 6053
rect 2002 5817 2087 6053
rect 2323 5817 2408 6053
rect 2644 5817 2729 6053
rect 2965 5817 3050 6053
rect 3286 5817 3371 6053
rect 3607 5817 3692 6053
rect 3928 5817 4013 6053
rect 4249 5817 4334 6053
rect 4570 5817 4655 6053
rect 4891 5817 4976 6053
rect 5212 5817 5297 6053
rect 5533 5817 5618 6053
rect 5854 5817 5939 6053
rect 6175 5817 6260 6053
rect 6496 5817 6581 6053
rect 6817 5817 6902 6053
rect 7138 5817 7223 6053
rect 7459 5817 7544 6053
rect 7780 5817 7865 6053
rect 8101 5817 8186 6053
rect 8422 5817 8507 6053
rect 8743 5817 8828 6053
rect 9064 5817 9149 6053
rect 9385 5817 9470 6053
rect 9706 5817 9791 6053
rect 10027 5817 10112 6053
rect 10348 5817 10433 6053
rect 10669 5817 10754 6053
rect 10990 5817 11075 6053
rect 11311 5817 11396 6053
rect 11632 5817 11717 6053
rect 11953 5817 12038 6053
rect 12274 5817 12358 6053
rect 12594 5817 12678 6053
rect 12914 5817 12998 6053
rect 13234 5817 13318 6053
rect 13554 5817 13638 6053
rect 13874 5817 13958 6053
rect 14194 5817 14278 6053
rect 14514 5817 14598 6053
rect 14834 5817 14918 6053
rect 15154 5817 15238 6053
rect 15474 5817 15558 6053
rect 15794 5817 16000 6053
rect 0 5447 16000 5817
rect 0 5211 161 5447
rect 397 5211 482 5447
rect 718 5211 803 5447
rect 1039 5211 1124 5447
rect 1360 5211 1445 5447
rect 1681 5211 1766 5447
rect 2002 5211 2087 5447
rect 2323 5211 2408 5447
rect 2644 5211 2729 5447
rect 2965 5211 3050 5447
rect 3286 5211 3371 5447
rect 3607 5211 3692 5447
rect 3928 5211 4013 5447
rect 4249 5211 4334 5447
rect 4570 5211 4655 5447
rect 4891 5211 4976 5447
rect 5212 5211 5297 5447
rect 5533 5211 5618 5447
rect 5854 5211 5939 5447
rect 6175 5211 6260 5447
rect 6496 5211 6581 5447
rect 6817 5211 6902 5447
rect 7138 5211 7223 5447
rect 7459 5211 7544 5447
rect 7780 5211 7865 5447
rect 8101 5211 8186 5447
rect 8422 5211 8507 5447
rect 8743 5211 8828 5447
rect 9064 5211 9149 5447
rect 9385 5211 9470 5447
rect 9706 5211 9791 5447
rect 10027 5211 10112 5447
rect 10348 5211 10433 5447
rect 10669 5211 10754 5447
rect 10990 5211 11075 5447
rect 11311 5211 11396 5447
rect 11632 5211 11717 5447
rect 11953 5211 12038 5447
rect 12274 5211 12358 5447
rect 12594 5211 12678 5447
rect 12914 5211 12998 5447
rect 13234 5211 13318 5447
rect 13554 5211 13638 5447
rect 13874 5211 13958 5447
rect 14194 5211 14278 5447
rect 14514 5211 14598 5447
rect 14834 5211 14918 5447
rect 15154 5211 15238 5447
rect 15474 5211 15558 5447
rect 15794 5211 16000 5447
rect 0 5187 16000 5211
rect 0 4843 16000 4867
rect 0 4607 161 4843
rect 397 4607 482 4843
rect 718 4607 803 4843
rect 1039 4607 1124 4843
rect 1360 4607 1445 4843
rect 1681 4607 1766 4843
rect 2002 4607 2087 4843
rect 2323 4607 2408 4843
rect 2644 4607 2729 4843
rect 2965 4607 3050 4843
rect 3286 4607 3371 4843
rect 3607 4607 3692 4843
rect 3928 4607 4013 4843
rect 4249 4607 4334 4843
rect 4570 4607 4655 4843
rect 4891 4607 4976 4843
rect 5212 4607 5297 4843
rect 5533 4607 5618 4843
rect 5854 4607 5939 4843
rect 6175 4607 6260 4843
rect 6496 4607 6581 4843
rect 6817 4607 6902 4843
rect 7138 4607 7223 4843
rect 7459 4607 7544 4843
rect 7780 4607 7865 4843
rect 8101 4607 8186 4843
rect 8422 4607 8507 4843
rect 8743 4607 8828 4843
rect 9064 4607 9149 4843
rect 9385 4607 9470 4843
rect 9706 4607 9791 4843
rect 10027 4607 10112 4843
rect 10348 4607 10433 4843
rect 10669 4607 10754 4843
rect 10990 4607 11075 4843
rect 11311 4607 11396 4843
rect 11632 4607 11717 4843
rect 11953 4607 12037 4843
rect 12273 4607 12357 4843
rect 12593 4607 12677 4843
rect 12913 4607 12997 4843
rect 13233 4607 13317 4843
rect 13553 4607 13637 4843
rect 13873 4607 13957 4843
rect 14193 4607 14277 4843
rect 14513 4607 14597 4843
rect 14833 4607 14917 4843
rect 15153 4607 15237 4843
rect 15473 4607 15557 4843
rect 15793 4607 16000 4843
rect 0 4237 16000 4607
rect 0 4001 161 4237
rect 397 4001 482 4237
rect 718 4001 803 4237
rect 1039 4001 1124 4237
rect 1360 4001 1445 4237
rect 1681 4001 1766 4237
rect 2002 4001 2087 4237
rect 2323 4001 2408 4237
rect 2644 4001 2729 4237
rect 2965 4001 3050 4237
rect 3286 4001 3371 4237
rect 3607 4001 3692 4237
rect 3928 4001 4013 4237
rect 4249 4001 4334 4237
rect 4570 4001 4655 4237
rect 4891 4001 4976 4237
rect 5212 4001 5297 4237
rect 5533 4001 5618 4237
rect 5854 4001 5939 4237
rect 6175 4001 6260 4237
rect 6496 4001 6581 4237
rect 6817 4001 6902 4237
rect 7138 4001 7223 4237
rect 7459 4001 7544 4237
rect 7780 4001 7865 4237
rect 8101 4001 8186 4237
rect 8422 4001 8507 4237
rect 8743 4001 8828 4237
rect 9064 4001 9149 4237
rect 9385 4001 9470 4237
rect 9706 4001 9791 4237
rect 10027 4001 10112 4237
rect 10348 4001 10433 4237
rect 10669 4001 10754 4237
rect 10990 4001 11075 4237
rect 11311 4001 11396 4237
rect 11632 4001 11717 4237
rect 11953 4001 12037 4237
rect 12273 4001 12357 4237
rect 12593 4001 12677 4237
rect 12913 4001 12997 4237
rect 13233 4001 13317 4237
rect 13553 4001 13637 4237
rect 13873 4001 13957 4237
rect 14193 4001 14277 4237
rect 14513 4001 14597 4237
rect 14833 4001 14917 4237
rect 15153 4001 15237 4237
rect 15473 4001 15557 4237
rect 15793 4001 16000 4237
rect 0 3977 16000 4001
rect 0 3633 16000 3657
rect 0 3397 162 3633
rect 398 3397 483 3633
rect 719 3397 804 3633
rect 1040 3397 1125 3633
rect 1361 3397 1446 3633
rect 1682 3397 1767 3633
rect 2003 3397 2088 3633
rect 2324 3397 2409 3633
rect 2645 3397 2730 3633
rect 2966 3397 3051 3633
rect 3287 3397 3372 3633
rect 3608 3397 3693 3633
rect 3929 3397 4014 3633
rect 4250 3397 4335 3633
rect 4571 3397 4656 3633
rect 4892 3397 4977 3633
rect 5213 3397 5298 3633
rect 5534 3397 5619 3633
rect 5855 3397 5940 3633
rect 6176 3397 6261 3633
rect 6497 3397 6582 3633
rect 6818 3397 6903 3633
rect 7139 3397 7224 3633
rect 7460 3397 7545 3633
rect 7781 3397 7866 3633
rect 8102 3397 8187 3633
rect 8423 3397 8508 3633
rect 8744 3397 8829 3633
rect 9065 3397 9150 3633
rect 9386 3397 9471 3633
rect 9707 3397 9792 3633
rect 10028 3397 10113 3633
rect 10349 3397 10434 3633
rect 10670 3397 10755 3633
rect 10991 3397 11076 3633
rect 11312 3397 11397 3633
rect 11633 3397 11718 3633
rect 11954 3397 12038 3633
rect 12274 3397 12358 3633
rect 12594 3397 12678 3633
rect 12914 3397 12998 3633
rect 13234 3397 13318 3633
rect 13554 3397 13638 3633
rect 13874 3397 13958 3633
rect 14194 3397 14278 3633
rect 14514 3397 14598 3633
rect 14834 3397 14918 3633
rect 15154 3397 15238 3633
rect 15474 3397 15558 3633
rect 15794 3397 16000 3633
rect 0 3267 16000 3397
rect 0 3031 162 3267
rect 398 3031 483 3267
rect 719 3031 804 3267
rect 1040 3031 1125 3267
rect 1361 3031 1446 3267
rect 1682 3031 1767 3267
rect 2003 3031 2088 3267
rect 2324 3031 2409 3267
rect 2645 3031 2730 3267
rect 2966 3031 3051 3267
rect 3287 3031 3372 3267
rect 3608 3031 3693 3267
rect 3929 3031 4014 3267
rect 4250 3031 4335 3267
rect 4571 3031 4656 3267
rect 4892 3031 4977 3267
rect 5213 3031 5298 3267
rect 5534 3031 5619 3267
rect 5855 3031 5940 3267
rect 6176 3031 6261 3267
rect 6497 3031 6582 3267
rect 6818 3031 6903 3267
rect 7139 3031 7224 3267
rect 7460 3031 7545 3267
rect 7781 3031 7866 3267
rect 8102 3031 8187 3267
rect 8423 3031 8508 3267
rect 8744 3031 8829 3267
rect 9065 3031 9150 3267
rect 9386 3031 9471 3267
rect 9707 3031 9792 3267
rect 10028 3031 10113 3267
rect 10349 3031 10434 3267
rect 10670 3031 10755 3267
rect 10991 3031 11076 3267
rect 11312 3031 11397 3267
rect 11633 3031 11718 3267
rect 11954 3031 12038 3267
rect 12274 3031 12358 3267
rect 12594 3031 12678 3267
rect 12914 3031 12998 3267
rect 13234 3031 13318 3267
rect 13554 3031 13638 3267
rect 13874 3031 13958 3267
rect 14194 3031 14278 3267
rect 14514 3031 14598 3267
rect 14834 3031 14918 3267
rect 15154 3031 15238 3267
rect 15474 3031 15558 3267
rect 15794 3031 16000 3267
rect 0 3007 16000 3031
rect 0 2663 16000 2687
rect 0 2427 163 2663
rect 399 2427 484 2663
rect 720 2427 805 2663
rect 1041 2427 1126 2663
rect 1362 2427 1447 2663
rect 1683 2427 1768 2663
rect 2004 2427 2089 2663
rect 2325 2427 2410 2663
rect 2646 2427 2731 2663
rect 2967 2427 3052 2663
rect 3288 2427 3373 2663
rect 3609 2427 3694 2663
rect 3930 2427 4015 2663
rect 4251 2427 4336 2663
rect 4572 2427 4657 2663
rect 4893 2427 4978 2663
rect 5214 2427 5299 2663
rect 5535 2427 5620 2663
rect 5856 2427 5941 2663
rect 6177 2427 6262 2663
rect 6498 2427 6583 2663
rect 6819 2427 6904 2663
rect 7140 2427 7225 2663
rect 7461 2427 7546 2663
rect 7782 2427 7867 2663
rect 8103 2427 8188 2663
rect 8424 2427 8509 2663
rect 8745 2427 8830 2663
rect 9066 2427 9151 2663
rect 9387 2427 9472 2663
rect 9708 2427 9793 2663
rect 10029 2427 10114 2663
rect 10350 2427 10435 2663
rect 10671 2427 10756 2663
rect 10992 2427 11077 2663
rect 11313 2427 11397 2663
rect 11633 2427 11717 2663
rect 11953 2427 12037 2663
rect 12273 2427 12357 2663
rect 12593 2427 12677 2663
rect 12913 2427 12997 2663
rect 13233 2427 13317 2663
rect 13553 2427 13637 2663
rect 13873 2427 13957 2663
rect 14193 2427 14277 2663
rect 14513 2427 14597 2663
rect 14833 2427 14917 2663
rect 15153 2427 15237 2663
rect 15473 2427 15557 2663
rect 15793 2427 16000 2663
rect 0 2057 16000 2427
rect 0 1821 163 2057
rect 399 1821 484 2057
rect 720 1821 805 2057
rect 1041 1821 1126 2057
rect 1362 1821 1447 2057
rect 1683 1821 1768 2057
rect 2004 1821 2089 2057
rect 2325 1821 2410 2057
rect 2646 1821 2731 2057
rect 2967 1821 3052 2057
rect 3288 1821 3373 2057
rect 3609 1821 3694 2057
rect 3930 1821 4015 2057
rect 4251 1821 4336 2057
rect 4572 1821 4657 2057
rect 4893 1821 4978 2057
rect 5214 1821 5299 2057
rect 5535 1821 5620 2057
rect 5856 1821 5941 2057
rect 6177 1821 6262 2057
rect 6498 1821 6583 2057
rect 6819 1821 6904 2057
rect 7140 1821 7225 2057
rect 7461 1821 7546 2057
rect 7782 1821 7867 2057
rect 8103 1821 8188 2057
rect 8424 1821 8509 2057
rect 8745 1821 8830 2057
rect 9066 1821 9151 2057
rect 9387 1821 9472 2057
rect 9708 1821 9793 2057
rect 10029 1821 10114 2057
rect 10350 1821 10435 2057
rect 10671 1821 10756 2057
rect 10992 1821 11077 2057
rect 11313 1821 11397 2057
rect 11633 1821 11717 2057
rect 11953 1821 12037 2057
rect 12273 1821 12357 2057
rect 12593 1821 12677 2057
rect 12913 1821 12997 2057
rect 13233 1821 13317 2057
rect 13553 1821 13637 2057
rect 13873 1821 13957 2057
rect 14193 1821 14277 2057
rect 14513 1821 14597 2057
rect 14833 1821 14917 2057
rect 15153 1821 15237 2057
rect 15473 1821 15557 2057
rect 15793 1821 16000 2057
rect 0 1797 16000 1821
rect 0 1452 16000 1477
rect 0 1216 162 1452
rect 398 1216 483 1452
rect 719 1216 804 1452
rect 1040 1216 1125 1452
rect 1361 1216 1446 1452
rect 1682 1216 1767 1452
rect 2003 1216 2088 1452
rect 2324 1216 2409 1452
rect 2645 1216 2730 1452
rect 2966 1216 3051 1452
rect 3287 1216 3372 1452
rect 3608 1216 3693 1452
rect 3929 1216 4014 1452
rect 4250 1216 4335 1452
rect 4571 1216 4656 1452
rect 4892 1216 4977 1452
rect 5213 1216 5298 1452
rect 5534 1216 5619 1452
rect 5855 1216 5940 1452
rect 6176 1216 6261 1452
rect 6497 1216 6582 1452
rect 6818 1216 6903 1452
rect 7139 1216 7224 1452
rect 7460 1216 7545 1452
rect 7781 1216 7866 1452
rect 8102 1216 8187 1452
rect 8423 1216 8508 1452
rect 8744 1216 8829 1452
rect 9065 1216 9150 1452
rect 9386 1216 9471 1452
rect 9707 1216 9792 1452
rect 10028 1216 10113 1452
rect 10349 1216 10434 1452
rect 10670 1216 10755 1452
rect 10991 1216 11076 1452
rect 11312 1216 11397 1452
rect 11633 1216 11718 1452
rect 11954 1216 12038 1452
rect 12274 1216 12358 1452
rect 12594 1216 12678 1452
rect 12914 1216 12998 1452
rect 13234 1216 13318 1452
rect 13554 1216 13638 1452
rect 13874 1216 13958 1452
rect 14194 1216 14278 1452
rect 14514 1216 14598 1452
rect 14834 1216 14918 1452
rect 15154 1216 15238 1452
rect 15474 1216 15558 1452
rect 15794 1216 16000 1452
rect 0 1070 16000 1216
rect 0 834 162 1070
rect 398 834 483 1070
rect 719 834 804 1070
rect 1040 834 1125 1070
rect 1361 834 1446 1070
rect 1682 834 1767 1070
rect 2003 834 2088 1070
rect 2324 834 2409 1070
rect 2645 834 2730 1070
rect 2966 834 3051 1070
rect 3287 834 3372 1070
rect 3608 834 3693 1070
rect 3929 834 4014 1070
rect 4250 834 4335 1070
rect 4571 834 4656 1070
rect 4892 834 4977 1070
rect 5213 834 5298 1070
rect 5534 834 5619 1070
rect 5855 834 5940 1070
rect 6176 834 6261 1070
rect 6497 834 6582 1070
rect 6818 834 6903 1070
rect 7139 834 7224 1070
rect 7460 834 7545 1070
rect 7781 834 7866 1070
rect 8102 834 8187 1070
rect 8423 834 8508 1070
rect 8744 834 8829 1070
rect 9065 834 9150 1070
rect 9386 834 9471 1070
rect 9707 834 9792 1070
rect 10028 834 10113 1070
rect 10349 834 10434 1070
rect 10670 834 10755 1070
rect 10991 834 11076 1070
rect 11312 834 11397 1070
rect 11633 834 11718 1070
rect 11954 834 12038 1070
rect 12274 834 12358 1070
rect 12594 834 12678 1070
rect 12914 834 12998 1070
rect 13234 834 13318 1070
rect 13554 834 13638 1070
rect 13874 834 13958 1070
rect 14194 834 14278 1070
rect 14514 834 14598 1070
rect 14834 834 14918 1070
rect 15154 834 15238 1070
rect 15474 834 15558 1070
rect 15794 834 16000 1070
rect 0 688 16000 834
rect 0 452 162 688
rect 398 452 483 688
rect 719 452 804 688
rect 1040 452 1125 688
rect 1361 452 1446 688
rect 1682 452 1767 688
rect 2003 452 2088 688
rect 2324 452 2409 688
rect 2645 452 2730 688
rect 2966 452 3051 688
rect 3287 452 3372 688
rect 3608 452 3693 688
rect 3929 452 4014 688
rect 4250 452 4335 688
rect 4571 452 4656 688
rect 4892 452 4977 688
rect 5213 452 5298 688
rect 5534 452 5619 688
rect 5855 452 5940 688
rect 6176 452 6261 688
rect 6497 452 6582 688
rect 6818 452 6903 688
rect 7139 452 7224 688
rect 7460 452 7545 688
rect 7781 452 7866 688
rect 8102 452 8187 688
rect 8423 452 8508 688
rect 8744 452 8829 688
rect 9065 452 9150 688
rect 9386 452 9471 688
rect 9707 452 9792 688
rect 10028 452 10113 688
rect 10349 452 10434 688
rect 10670 452 10755 688
rect 10991 452 11076 688
rect 11312 452 11397 688
rect 11633 452 11718 688
rect 11954 452 12038 688
rect 12274 452 12358 688
rect 12594 452 12678 688
rect 12914 452 12998 688
rect 13234 452 13318 688
rect 13554 452 13638 688
rect 13874 452 13958 688
rect 14194 452 14278 688
rect 14514 452 14598 688
rect 14834 452 14918 688
rect 15154 452 15238 688
rect 15474 452 15558 688
rect 15794 452 16000 688
rect 0 427 16000 452
use sky130_fd_io__overlay_gpiov2_m4  sky130_fd_io__overlay_gpiov2_m4_0
timestamp 1649977179
transform 1 0 0 0 1 0
box 0 407 16000 40000
<< labels >>
flabel metal5 s 6374 25521 10682 29830 3 FreeSans 2000 0 0 0 PAD
port 1 nsew signal default
flabel metal5 s 0 35157 254 40000 3 FreeSans 520 0 0 0 VSSIO
port 2 nsew ground bidirectional
flabel metal5 s 15746 35157 16000 40000 3 FreeSans 520 180 0 0 VSSIO
port 2 nsew ground bidirectional
flabel metal5 s 15746 3977 16000 4867 3 FreeSans 520 180 0 0 VDDIO
port 3 nsew power bidirectional
flabel metal5 s 15746 427 16000 1477 3 FreeSans 520 180 0 0 VCCHIB
port 4 nsew power bidirectional
flabel metal5 s 15746 14007 16000 18997 3 FreeSans 520 180 0 0 VDDIO
port 3 nsew power bidirectional
flabel metal5 s 15746 12837 16000 13687 3 FreeSans 520 180 0 0 VDDIO_Q
port 5 nsew power bidirectional
flabel metal5 s 15746 1797 16000 2687 3 FreeSans 520 180 0 0 VCCD
port 6 nsew power bidirectional
flabel metal5 s 15746 7368 16000 8017 3 FreeSans 520 180 0 0 VSSA
port 7 nsew ground bidirectional
flabel metal5 s 15746 6397 16000 7047 3 FreeSans 520 180 0 0 VSWITCH
port 8 nsew power bidirectional
flabel metal5 s 15746 5187 16000 6077 3 FreeSans 520 180 0 0 VSSIO
port 2 nsew ground bidirectional
flabel metal5 s 15746 11667 16000 12517 3 FreeSans 520 180 0 0 VSSIO_Q
port 9 nsew ground bidirectional
flabel metal5 s 15746 8337 16000 9227 3 FreeSans 520 180 0 0 VSSD
port 10 nsew ground bidirectional
flabel metal5 s 15807 3007 16000 3657 3 FreeSans 520 180 0 0 VDDA
port 11 nsew power bidirectional
flabel metal5 s 15746 9547 16000 11347 3 FreeSans 520 180 0 0 VSSA
port 7 nsew ground bidirectional
flabel metal5 s 0 427 254 1477 3 FreeSans 520 0 0 0 VCCHIB
port 4 nsew power bidirectional
flabel metal5 s 0 7368 254 8017 3 FreeSans 520 0 0 0 VSSA
port 7 nsew ground bidirectional
flabel metal5 s 0 9547 254 11347 3 FreeSans 520 0 0 0 VSSA
port 7 nsew ground bidirectional
flabel metal5 s 0 12837 254 13687 3 FreeSans 520 0 0 0 VDDIO_Q
port 5 nsew power bidirectional
flabel metal5 s 0 1797 254 2687 3 FreeSans 520 0 0 0 VCCD
port 6 nsew power bidirectional
flabel metal5 s 0 3977 254 4867 3 FreeSans 520 0 0 0 VDDIO
port 3 nsew power bidirectional
flabel metal5 s 0 3007 193 3657 3 FreeSans 520 0 0 0 VDDA
port 11 nsew power bidirectional
flabel metal5 s 0 5187 254 6077 3 FreeSans 520 0 0 0 VSSIO
port 2 nsew ground bidirectional
flabel metal5 s 0 6397 254 7047 3 FreeSans 520 0 0 0 VSWITCH
port 8 nsew power bidirectional
flabel metal5 s 0 11667 254 12517 3 FreeSans 520 0 0 0 VSSIO_Q
port 9 nsew ground bidirectional
flabel metal5 s 0 8337 254 9227 3 FreeSans 520 0 0 0 VSSD
port 10 nsew ground bidirectional
flabel metal5 s 0 14007 254 18997 3 FreeSans 520 0 0 0 VDDIO
port 3 nsew power bidirectional
flabel metal4 s 0 6377 254 7067 3 FreeSans 520 0 0 0 VSWITCH
port 8 nsew power bidirectional
flabel metal4 s 15746 6377 16000 7067 3 FreeSans 520 180 0 0 VSWITCH
port 8 nsew power bidirectional
flabel metal4 s 0 11647 254 12537 3 FreeSans 520 0 0 0 VSSIO_Q
port 9 nsew ground bidirectional
flabel metal4 s 15746 11647 16000 12537 3 FreeSans 520 180 0 0 VSSIO_Q
port 9 nsew ground bidirectional
flabel metal4 s 0 5167 254 6097 3 FreeSans 520 0 0 0 VSSIO
port 2 nsew ground bidirectional
flabel metal4 s 0 35157 254 40000 3 FreeSans 520 0 0 0 VSSIO
port 2 nsew ground bidirectional
flabel metal4 s 15746 5167 16000 6097 3 FreeSans 520 180 0 0 VSSIO
port 2 nsew ground bidirectional
flabel metal4 s 15746 35157 16000 40000 3 FreeSans 520 180 0 0 VSSIO
port 2 nsew ground bidirectional
flabel metal4 s 0 8317 254 9247 3 FreeSans 520 0 0 0 VSSD
port 10 nsew ground bidirectional
flabel metal4 s 15746 8317 16000 9247 3 FreeSans 520 180 0 0 VSSD
port 10 nsew ground bidirectional
flabel metal4 s 0 7347 254 8037 3 FreeSans 520 0 0 0 VSSA
port 7 nsew ground bidirectional
flabel metal4 s 0 11281 254 11347 3 FreeSans 520 0 0 0 VSSA
port 7 nsew ground bidirectional
flabel metal4 s 0 10329 254 10565 3 FreeSans 520 0 0 0 VSSA
port 7 nsew ground bidirectional
flabel metal4 s 0 9547 254 9613 3 FreeSans 520 0 0 0 VSSA
port 7 nsew ground bidirectional
flabel metal4 s 15746 7347 16000 8037 3 FreeSans 520 180 0 0 VSSA
port 7 nsew ground bidirectional
flabel metal4 s 15746 9547 16000 9613 3 FreeSans 520 180 0 0 VSSA
port 7 nsew ground bidirectional
flabel metal4 s 15746 11281 16000 11347 3 FreeSans 520 180 0 0 VSSA
port 7 nsew ground bidirectional
flabel metal4 s 15746 10329 16000 10565 3 FreeSans 520 180 0 0 VSSA
port 7 nsew ground bidirectional
flabel metal4 s 0 12817 254 13707 3 FreeSans 520 0 0 0 VDDIO_Q
port 5 nsew power bidirectional
flabel metal4 s 15746 12817 16000 13707 3 FreeSans 520 180 0 0 VDDIO_Q
port 5 nsew power bidirectional
flabel metal4 s 0 14007 254 19000 3 FreeSans 520 0 0 0 VDDIO
port 3 nsew power bidirectional
flabel metal4 s 0 3957 254 4887 3 FreeSans 520 0 0 0 VDDIO
port 3 nsew power bidirectional
flabel metal4 s 15746 14007 16000 19000 3 FreeSans 520 180 0 0 VDDIO
port 3 nsew power bidirectional
flabel metal4 s 15746 3957 16000 4887 3 FreeSans 520 180 0 0 VDDIO
port 3 nsew power bidirectional
flabel metal4 s 0 2987 193 3677 3 FreeSans 520 0 0 0 VDDA
port 11 nsew power bidirectional
flabel metal4 s 15807 2987 16000 3677 3 FreeSans 520 180 0 0 VDDA
port 11 nsew power bidirectional
flabel metal4 s 0 407 254 1497 3 FreeSans 520 0 0 0 VCCHIB
port 4 nsew power bidirectional
flabel metal4 s 15746 407 16000 1497 3 FreeSans 520 180 0 0 VCCHIB
port 4 nsew power bidirectional
flabel metal4 s 15746 10625 16000 11221 3 FreeSans 520 180 0 0 AMUXBUS_A
port 12 nsew signal default
flabel metal4 s 0 10625 254 11221 3 FreeSans 520 0 0 0 AMUXBUS_A
port 12 nsew signal default
flabel metal4 s 15746 9673 16000 10269 3 FreeSans 520 180 0 0 AMUXBUS_B
port 13 nsew signal default
flabel metal4 s 0 9673 254 10269 3 FreeSans 520 0 0 0 AMUXBUS_B
port 13 nsew signal default
flabel metal4 s 15746 1777 16000 2707 3 FreeSans 520 180 0 0 VCCD
port 6 nsew power bidirectional
flabel metal4 s 0 1777 254 2707 3 FreeSans 520 0 0 0 VCCD
port 6 nsew power bidirectional
rlabel metal4 s 15746 10625 16000 11221 1 AMUXBUS_A
port 12 nsew signal default
rlabel metal4 s 15746 9673 16000 10269 1 AMUXBUS_B
port 13 nsew signal default
rlabel metal5 s 0 1797 16000 2687 1 VCCD
port 6 nsew power bidirectional
rlabel metal5 s 0 427 16000 1477 1 VCCHIB
port 4 nsew power bidirectional
rlabel metal4 s 15807 2987 16000 3677 1 VDDA
port 11 nsew power bidirectional
rlabel metal5 s 0 3007 16000 3657 1 VDDA
port 11 nsew power bidirectional
rlabel metal4 s 15746 18973 16000 19000 1 VDDIO
port 3 nsew power bidirectional
rlabel metal4 s 15746 14007 16000 14031 1 VDDIO
port 3 nsew power bidirectional
rlabel metal4 s 0 18973 254 19000 1 VDDIO
port 3 nsew power bidirectional
rlabel metal4 s 0 14031 16000 18973 1 VDDIO
port 3 nsew power bidirectional
rlabel metal4 s 0 14007 254 14031 1 VDDIO
port 3 nsew power bidirectional
rlabel metal5 s 0 3977 16000 4867 1 VDDIO
port 3 nsew power bidirectional
rlabel metal5 s 0 14007 16000 18997 1 VDDIO
port 3 nsew power bidirectional
rlabel metal5 s 0 12837 16000 13687 1 VDDIO_Q
port 5 nsew power bidirectional
rlabel metal4 s 0 9547 254 9613 1 VSSA
port 7 nsew ground bidirectional
rlabel metal4 s 0 10329 16000 10565 1 VSSA
port 7 nsew ground bidirectional
rlabel metal4 s 0 11281 254 11347 1 VSSA
port 7 nsew ground bidirectional
rlabel metal4 s 15746 9547 16000 9613 1 VSSA
port 7 nsew ground bidirectional
rlabel metal4 s 15746 11281 16000 11347 1 VSSA
port 7 nsew ground bidirectional
rlabel metal5 s 0 7367 16000 8017 1 VSSA
port 7 nsew ground bidirectional
rlabel metal5 s 0 9547 16000 11347 1 VSSA
port 7 nsew ground bidirectional
rlabel metal5 s 0 8337 16000 9227 1 VSSD
port 10 nsew ground bidirectional
rlabel metal4 s 15746 6053 16000 6097 1 VSSIO
port 2 nsew ground bidirectional
rlabel metal4 s 15746 5167 16000 5211 1 VSSIO
port 2 nsew ground bidirectional
rlabel metal4 s 0 6053 254 6097 1 VSSIO
port 2 nsew ground bidirectional
rlabel metal4 s 0 5211 16000 6053 1 VSSIO
port 2 nsew ground bidirectional
rlabel metal4 s 0 5167 254 5211 1 VSSIO
port 2 nsew ground bidirectional
rlabel metal5 s 0 35157 16000 40000 1 VSSIO
port 2 nsew ground bidirectional
rlabel metal5 s 0 5187 16000 6077 1 VSSIO
port 2 nsew ground bidirectional
rlabel metal5 s 0 11667 16000 12517 1 VSSIO_Q
port 9 nsew ground bidirectional
rlabel metal5 s 0 6397 16000 7047 1 VSWITCH
port 8 nsew power bidirectional
<< properties >>
string FIXED_BBOX 0 0 16000 40000
string GDS_END 192116
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 18226
string LEFclass PAD
string LEFsymmetry X Y R90
<< end >>
