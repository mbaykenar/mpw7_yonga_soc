magic
tech sky130B
magscale 1 2
timestamp 1649977179
<< pwell >>
rect 15 163 867 817
<< nmoslvt >>
rect 171 189 201 791
rect 257 189 307 791
rect 363 189 413 791
rect 469 189 519 791
rect 575 189 625 791
rect 681 189 711 791
<< ndiff >>
rect 111 779 171 791
rect 111 745 126 779
rect 160 745 171 779
rect 111 711 171 745
rect 111 677 126 711
rect 160 677 171 711
rect 111 643 171 677
rect 111 609 126 643
rect 160 609 171 643
rect 111 575 171 609
rect 111 541 126 575
rect 160 541 171 575
rect 111 507 171 541
rect 111 473 126 507
rect 160 473 171 507
rect 111 439 171 473
rect 111 405 126 439
rect 160 405 171 439
rect 111 371 171 405
rect 111 337 126 371
rect 160 337 171 371
rect 111 303 171 337
rect 111 269 126 303
rect 160 269 171 303
rect 111 235 171 269
rect 111 201 126 235
rect 160 201 171 235
rect 111 189 171 201
rect 201 779 257 791
rect 201 745 212 779
rect 246 745 257 779
rect 201 711 257 745
rect 201 677 212 711
rect 246 677 257 711
rect 201 643 257 677
rect 201 609 212 643
rect 246 609 257 643
rect 201 575 257 609
rect 201 541 212 575
rect 246 541 257 575
rect 201 507 257 541
rect 201 473 212 507
rect 246 473 257 507
rect 201 439 257 473
rect 201 405 212 439
rect 246 405 257 439
rect 201 371 257 405
rect 201 337 212 371
rect 246 337 257 371
rect 201 303 257 337
rect 201 269 212 303
rect 246 269 257 303
rect 201 235 257 269
rect 201 201 212 235
rect 246 201 257 235
rect 201 189 257 201
rect 307 779 363 791
rect 307 745 318 779
rect 352 745 363 779
rect 307 711 363 745
rect 307 677 318 711
rect 352 677 363 711
rect 307 643 363 677
rect 307 609 318 643
rect 352 609 363 643
rect 307 575 363 609
rect 307 541 318 575
rect 352 541 363 575
rect 307 507 363 541
rect 307 473 318 507
rect 352 473 363 507
rect 307 439 363 473
rect 307 405 318 439
rect 352 405 363 439
rect 307 371 363 405
rect 307 337 318 371
rect 352 337 363 371
rect 307 303 363 337
rect 307 269 318 303
rect 352 269 363 303
rect 307 235 363 269
rect 307 201 318 235
rect 352 201 363 235
rect 307 189 363 201
rect 413 779 469 791
rect 413 745 424 779
rect 458 745 469 779
rect 413 711 469 745
rect 413 677 424 711
rect 458 677 469 711
rect 413 643 469 677
rect 413 609 424 643
rect 458 609 469 643
rect 413 575 469 609
rect 413 541 424 575
rect 458 541 469 575
rect 413 507 469 541
rect 413 473 424 507
rect 458 473 469 507
rect 413 439 469 473
rect 413 405 424 439
rect 458 405 469 439
rect 413 371 469 405
rect 413 337 424 371
rect 458 337 469 371
rect 413 303 469 337
rect 413 269 424 303
rect 458 269 469 303
rect 413 235 469 269
rect 413 201 424 235
rect 458 201 469 235
rect 413 189 469 201
rect 519 779 575 791
rect 519 745 530 779
rect 564 745 575 779
rect 519 711 575 745
rect 519 677 530 711
rect 564 677 575 711
rect 519 643 575 677
rect 519 609 530 643
rect 564 609 575 643
rect 519 575 575 609
rect 519 541 530 575
rect 564 541 575 575
rect 519 507 575 541
rect 519 473 530 507
rect 564 473 575 507
rect 519 439 575 473
rect 519 405 530 439
rect 564 405 575 439
rect 519 371 575 405
rect 519 337 530 371
rect 564 337 575 371
rect 519 303 575 337
rect 519 269 530 303
rect 564 269 575 303
rect 519 235 575 269
rect 519 201 530 235
rect 564 201 575 235
rect 519 189 575 201
rect 625 779 681 791
rect 625 745 636 779
rect 670 745 681 779
rect 625 711 681 745
rect 625 677 636 711
rect 670 677 681 711
rect 625 643 681 677
rect 625 609 636 643
rect 670 609 681 643
rect 625 575 681 609
rect 625 541 636 575
rect 670 541 681 575
rect 625 507 681 541
rect 625 473 636 507
rect 670 473 681 507
rect 625 439 681 473
rect 625 405 636 439
rect 670 405 681 439
rect 625 371 681 405
rect 625 337 636 371
rect 670 337 681 371
rect 625 303 681 337
rect 625 269 636 303
rect 670 269 681 303
rect 625 235 681 269
rect 625 201 636 235
rect 670 201 681 235
rect 625 189 681 201
rect 711 779 771 791
rect 711 745 722 779
rect 756 745 771 779
rect 711 711 771 745
rect 711 677 722 711
rect 756 677 771 711
rect 711 643 771 677
rect 711 609 722 643
rect 756 609 771 643
rect 711 575 771 609
rect 711 541 722 575
rect 756 541 771 575
rect 711 507 771 541
rect 711 473 722 507
rect 756 473 771 507
rect 711 439 771 473
rect 711 405 722 439
rect 756 405 771 439
rect 711 371 771 405
rect 711 337 722 371
rect 756 337 771 371
rect 711 303 771 337
rect 711 269 722 303
rect 756 269 771 303
rect 711 235 771 269
rect 711 201 722 235
rect 756 201 771 235
rect 711 189 771 201
<< ndiffc >>
rect 126 745 160 779
rect 126 677 160 711
rect 126 609 160 643
rect 126 541 160 575
rect 126 473 160 507
rect 126 405 160 439
rect 126 337 160 371
rect 126 269 160 303
rect 126 201 160 235
rect 212 745 246 779
rect 212 677 246 711
rect 212 609 246 643
rect 212 541 246 575
rect 212 473 246 507
rect 212 405 246 439
rect 212 337 246 371
rect 212 269 246 303
rect 212 201 246 235
rect 318 745 352 779
rect 318 677 352 711
rect 318 609 352 643
rect 318 541 352 575
rect 318 473 352 507
rect 318 405 352 439
rect 318 337 352 371
rect 318 269 352 303
rect 318 201 352 235
rect 424 745 458 779
rect 424 677 458 711
rect 424 609 458 643
rect 424 541 458 575
rect 424 473 458 507
rect 424 405 458 439
rect 424 337 458 371
rect 424 269 458 303
rect 424 201 458 235
rect 530 745 564 779
rect 530 677 564 711
rect 530 609 564 643
rect 530 541 564 575
rect 530 473 564 507
rect 530 405 564 439
rect 530 337 564 371
rect 530 269 564 303
rect 530 201 564 235
rect 636 745 670 779
rect 636 677 670 711
rect 636 609 670 643
rect 636 541 670 575
rect 636 473 670 507
rect 636 405 670 439
rect 636 337 670 371
rect 636 269 670 303
rect 636 201 670 235
rect 722 745 756 779
rect 722 677 756 711
rect 722 609 756 643
rect 722 541 756 575
rect 722 473 756 507
rect 722 405 756 439
rect 722 337 756 371
rect 722 269 756 303
rect 722 201 756 235
<< psubdiff >>
rect 41 779 111 791
rect 41 745 58 779
rect 92 745 111 779
rect 41 711 111 745
rect 41 677 58 711
rect 92 677 111 711
rect 41 643 111 677
rect 41 609 58 643
rect 92 609 111 643
rect 41 575 111 609
rect 41 541 58 575
rect 92 541 111 575
rect 41 507 111 541
rect 41 473 58 507
rect 92 473 111 507
rect 41 439 111 473
rect 41 405 58 439
rect 92 405 111 439
rect 41 371 111 405
rect 41 337 58 371
rect 92 337 111 371
rect 41 303 111 337
rect 41 269 58 303
rect 92 269 111 303
rect 41 235 111 269
rect 41 201 58 235
rect 92 201 111 235
rect 41 189 111 201
rect 771 779 841 791
rect 771 745 790 779
rect 824 745 841 779
rect 771 711 841 745
rect 771 677 790 711
rect 824 677 841 711
rect 771 643 841 677
rect 771 609 790 643
rect 824 609 841 643
rect 771 575 841 609
rect 771 541 790 575
rect 824 541 841 575
rect 771 507 841 541
rect 771 473 790 507
rect 824 473 841 507
rect 771 439 841 473
rect 771 405 790 439
rect 824 405 841 439
rect 771 371 841 405
rect 771 337 790 371
rect 824 337 841 371
rect 771 303 841 337
rect 771 269 790 303
rect 824 269 841 303
rect 771 235 841 269
rect 771 201 790 235
rect 824 201 841 235
rect 771 189 841 201
<< psubdiffcont >>
rect 58 745 92 779
rect 58 677 92 711
rect 58 609 92 643
rect 58 541 92 575
rect 58 473 92 507
rect 58 405 92 439
rect 58 337 92 371
rect 58 269 92 303
rect 58 201 92 235
rect 790 745 824 779
rect 790 677 824 711
rect 790 609 824 643
rect 790 541 824 575
rect 790 473 824 507
rect 790 405 824 439
rect 790 337 824 371
rect 790 269 824 303
rect 790 201 824 235
<< poly >>
rect 243 959 639 980
rect 120 867 201 883
rect 120 833 136 867
rect 170 833 201 867
rect 243 857 288 959
rect 594 857 639 959
rect 243 841 639 857
rect 681 867 762 883
rect 120 817 201 833
rect 171 791 201 817
rect 257 791 307 841
rect 363 791 413 841
rect 469 791 519 841
rect 575 791 625 841
rect 681 833 712 867
rect 746 833 762 867
rect 681 817 762 833
rect 681 791 711 817
rect 171 163 201 189
rect 120 147 201 163
rect 120 113 136 147
rect 170 113 201 147
rect 257 139 307 189
rect 363 139 413 189
rect 469 139 519 189
rect 575 139 625 189
rect 681 163 711 189
rect 681 147 762 163
rect 120 97 201 113
rect 243 123 639 139
rect 243 21 288 123
rect 594 21 639 123
rect 681 113 712 147
rect 746 113 762 147
rect 681 97 762 113
rect 243 0 639 21
<< polycont >>
rect 136 833 170 867
rect 288 857 594 959
rect 712 833 746 867
rect 136 113 170 147
rect 288 21 594 123
rect 712 113 746 147
<< locali >>
rect 266 961 616 980
rect 120 867 186 883
rect 120 833 136 867
rect 170 833 186 867
rect 266 855 280 961
rect 602 855 616 961
rect 266 841 616 855
rect 696 867 762 883
rect 120 817 186 833
rect 696 833 712 867
rect 746 833 762 867
rect 696 817 762 833
rect 120 795 160 817
rect 722 795 762 817
rect 41 779 160 795
rect 41 745 58 779
rect 92 759 126 779
rect 94 745 126 759
rect 41 725 60 745
rect 94 725 160 745
rect 41 711 160 725
rect 41 677 58 711
rect 92 687 126 711
rect 94 677 126 687
rect 41 653 60 677
rect 94 653 160 677
rect 41 643 160 653
rect 41 609 58 643
rect 92 615 126 643
rect 94 609 126 615
rect 41 581 60 609
rect 94 581 160 609
rect 41 575 160 581
rect 41 541 58 575
rect 92 543 126 575
rect 94 541 126 543
rect 41 509 60 541
rect 94 509 160 541
rect 41 507 160 509
rect 41 473 58 507
rect 92 473 126 507
rect 41 471 160 473
rect 41 439 60 471
rect 94 439 160 471
rect 41 405 58 439
rect 94 437 126 439
rect 92 405 126 437
rect 41 399 160 405
rect 41 371 60 399
rect 94 371 160 399
rect 41 337 58 371
rect 94 365 126 371
rect 92 337 126 365
rect 41 327 160 337
rect 41 303 60 327
rect 94 303 160 327
rect 41 269 58 303
rect 94 293 126 303
rect 92 269 126 293
rect 41 255 160 269
rect 41 235 60 255
rect 94 235 160 255
rect 41 201 58 235
rect 94 221 126 235
rect 92 201 126 221
rect 41 185 160 201
rect 212 779 246 795
rect 212 711 246 725
rect 212 643 246 653
rect 212 575 246 581
rect 212 507 246 509
rect 212 471 246 473
rect 212 399 246 405
rect 212 327 246 337
rect 212 255 246 269
rect 212 185 246 201
rect 318 779 352 795
rect 318 711 352 725
rect 318 643 352 653
rect 318 575 352 581
rect 318 507 352 509
rect 318 471 352 473
rect 318 399 352 405
rect 318 327 352 337
rect 318 255 352 269
rect 318 185 352 201
rect 424 779 458 795
rect 424 711 458 725
rect 424 643 458 653
rect 424 575 458 581
rect 424 507 458 509
rect 424 471 458 473
rect 424 399 458 405
rect 424 327 458 337
rect 424 255 458 269
rect 424 185 458 201
rect 530 779 564 795
rect 530 711 564 725
rect 530 643 564 653
rect 530 575 564 581
rect 530 507 564 509
rect 530 471 564 473
rect 530 399 564 405
rect 530 327 564 337
rect 530 255 564 269
rect 530 185 564 201
rect 636 779 670 795
rect 636 711 670 725
rect 636 643 670 653
rect 636 575 670 581
rect 636 507 670 509
rect 636 471 670 473
rect 636 399 670 405
rect 636 327 670 337
rect 636 255 670 269
rect 636 185 670 201
rect 722 779 841 795
rect 756 759 790 779
rect 756 745 788 759
rect 824 745 841 779
rect 722 725 788 745
rect 822 725 841 745
rect 722 711 841 725
rect 756 687 790 711
rect 756 677 788 687
rect 824 677 841 711
rect 722 653 788 677
rect 822 653 841 677
rect 722 643 841 653
rect 756 615 790 643
rect 756 609 788 615
rect 824 609 841 643
rect 722 581 788 609
rect 822 581 841 609
rect 722 575 841 581
rect 756 543 790 575
rect 756 541 788 543
rect 824 541 841 575
rect 722 509 788 541
rect 822 509 841 541
rect 722 507 841 509
rect 756 473 790 507
rect 824 473 841 507
rect 722 471 841 473
rect 722 439 788 471
rect 822 439 841 471
rect 756 437 788 439
rect 756 405 790 437
rect 824 405 841 439
rect 722 399 841 405
rect 722 371 788 399
rect 822 371 841 399
rect 756 365 788 371
rect 756 337 790 365
rect 824 337 841 371
rect 722 327 841 337
rect 722 303 788 327
rect 822 303 841 327
rect 756 293 788 303
rect 756 269 790 293
rect 824 269 841 303
rect 722 255 841 269
rect 722 235 788 255
rect 822 235 841 255
rect 756 221 788 235
rect 756 201 790 221
rect 824 201 841 235
rect 722 185 841 201
rect 120 163 160 185
rect 722 163 762 185
rect 120 147 186 163
rect 120 113 136 147
rect 170 113 186 147
rect 696 147 762 163
rect 120 97 186 113
rect 266 125 616 139
rect 266 19 280 125
rect 602 19 616 125
rect 696 113 712 147
rect 746 113 762 147
rect 696 97 762 113
rect 266 0 616 19
<< viali >>
rect 280 959 602 961
rect 280 857 288 959
rect 288 857 594 959
rect 594 857 602 959
rect 280 855 602 857
rect 60 745 92 759
rect 92 745 94 759
rect 60 725 94 745
rect 60 677 92 687
rect 92 677 94 687
rect 60 653 94 677
rect 60 609 92 615
rect 92 609 94 615
rect 60 581 94 609
rect 60 541 92 543
rect 92 541 94 543
rect 60 509 94 541
rect 60 439 94 471
rect 60 437 92 439
rect 92 437 94 439
rect 60 371 94 399
rect 60 365 92 371
rect 92 365 94 371
rect 60 303 94 327
rect 60 293 92 303
rect 92 293 94 303
rect 60 235 94 255
rect 60 221 92 235
rect 92 221 94 235
rect 212 745 246 759
rect 212 725 246 745
rect 212 677 246 687
rect 212 653 246 677
rect 212 609 246 615
rect 212 581 246 609
rect 212 541 246 543
rect 212 509 246 541
rect 212 439 246 471
rect 212 437 246 439
rect 212 371 246 399
rect 212 365 246 371
rect 212 303 246 327
rect 212 293 246 303
rect 212 235 246 255
rect 212 221 246 235
rect 318 745 352 759
rect 318 725 352 745
rect 318 677 352 687
rect 318 653 352 677
rect 318 609 352 615
rect 318 581 352 609
rect 318 541 352 543
rect 318 509 352 541
rect 318 439 352 471
rect 318 437 352 439
rect 318 371 352 399
rect 318 365 352 371
rect 318 303 352 327
rect 318 293 352 303
rect 318 235 352 255
rect 318 221 352 235
rect 424 745 458 759
rect 424 725 458 745
rect 424 677 458 687
rect 424 653 458 677
rect 424 609 458 615
rect 424 581 458 609
rect 424 541 458 543
rect 424 509 458 541
rect 424 439 458 471
rect 424 437 458 439
rect 424 371 458 399
rect 424 365 458 371
rect 424 303 458 327
rect 424 293 458 303
rect 424 235 458 255
rect 424 221 458 235
rect 530 745 564 759
rect 530 725 564 745
rect 530 677 564 687
rect 530 653 564 677
rect 530 609 564 615
rect 530 581 564 609
rect 530 541 564 543
rect 530 509 564 541
rect 530 439 564 471
rect 530 437 564 439
rect 530 371 564 399
rect 530 365 564 371
rect 530 303 564 327
rect 530 293 564 303
rect 530 235 564 255
rect 530 221 564 235
rect 636 745 670 759
rect 636 725 670 745
rect 636 677 670 687
rect 636 653 670 677
rect 636 609 670 615
rect 636 581 670 609
rect 636 541 670 543
rect 636 509 670 541
rect 636 439 670 471
rect 636 437 670 439
rect 636 371 670 399
rect 636 365 670 371
rect 636 303 670 327
rect 636 293 670 303
rect 636 235 670 255
rect 636 221 670 235
rect 788 745 790 759
rect 790 745 822 759
rect 788 725 822 745
rect 788 677 790 687
rect 790 677 822 687
rect 788 653 822 677
rect 788 609 790 615
rect 790 609 822 615
rect 788 581 822 609
rect 788 541 790 543
rect 790 541 822 543
rect 788 509 822 541
rect 788 439 822 471
rect 788 437 790 439
rect 790 437 822 439
rect 788 371 822 399
rect 788 365 790 371
rect 790 365 822 371
rect 788 303 822 327
rect 788 293 790 303
rect 790 293 822 303
rect 788 235 822 255
rect 788 221 790 235
rect 790 221 822 235
rect 280 123 602 125
rect 280 21 288 123
rect 288 21 594 123
rect 594 21 602 123
rect 280 19 602 21
<< metal1 >>
rect 264 961 618 980
rect 264 855 280 961
rect 602 855 618 961
rect 264 843 618 855
rect 41 759 100 771
rect 41 725 60 759
rect 94 725 100 759
rect 41 687 100 725
rect 41 653 60 687
rect 94 653 100 687
rect 41 615 100 653
rect 41 581 60 615
rect 94 581 100 615
rect 41 543 100 581
rect 41 509 60 543
rect 94 509 100 543
rect 41 471 100 509
rect 41 437 60 471
rect 94 437 100 471
rect 41 399 100 437
rect 41 365 60 399
rect 94 365 100 399
rect 41 327 100 365
rect 41 293 60 327
rect 94 293 100 327
rect 41 255 100 293
rect 41 221 60 255
rect 94 221 100 255
rect 41 209 100 221
rect 203 759 255 771
rect 203 725 212 759
rect 246 725 255 759
rect 203 687 255 725
rect 203 653 212 687
rect 246 653 255 687
rect 203 615 255 653
rect 203 581 212 615
rect 246 581 255 615
rect 203 543 255 581
rect 203 509 212 543
rect 246 509 255 543
rect 203 471 255 509
rect 203 459 212 471
rect 246 459 255 471
rect 203 399 255 407
rect 203 395 212 399
rect 246 395 255 399
rect 203 331 255 343
rect 203 267 255 279
rect 203 209 255 215
rect 309 765 361 771
rect 309 701 361 713
rect 309 637 361 649
rect 309 581 318 585
rect 352 581 361 585
rect 309 573 361 581
rect 309 509 318 521
rect 352 509 361 521
rect 309 471 361 509
rect 309 437 318 471
rect 352 437 361 471
rect 309 399 361 437
rect 309 365 318 399
rect 352 365 361 399
rect 309 327 361 365
rect 309 293 318 327
rect 352 293 361 327
rect 309 255 361 293
rect 309 221 318 255
rect 352 221 361 255
rect 309 209 361 221
rect 415 759 467 771
rect 415 725 424 759
rect 458 725 467 759
rect 415 687 467 725
rect 415 653 424 687
rect 458 653 467 687
rect 415 615 467 653
rect 415 581 424 615
rect 458 581 467 615
rect 415 543 467 581
rect 415 509 424 543
rect 458 509 467 543
rect 415 471 467 509
rect 415 459 424 471
rect 458 459 467 471
rect 415 399 467 407
rect 415 395 424 399
rect 458 395 467 399
rect 415 331 467 343
rect 415 267 467 279
rect 415 209 467 215
rect 521 765 573 771
rect 521 701 573 713
rect 521 637 573 649
rect 521 581 530 585
rect 564 581 573 585
rect 521 573 573 581
rect 521 509 530 521
rect 564 509 573 521
rect 521 471 573 509
rect 521 437 530 471
rect 564 437 573 471
rect 521 399 573 437
rect 521 365 530 399
rect 564 365 573 399
rect 521 327 573 365
rect 521 293 530 327
rect 564 293 573 327
rect 521 255 573 293
rect 521 221 530 255
rect 564 221 573 255
rect 521 209 573 221
rect 627 759 679 771
rect 627 725 636 759
rect 670 725 679 759
rect 627 687 679 725
rect 627 653 636 687
rect 670 653 679 687
rect 627 615 679 653
rect 627 581 636 615
rect 670 581 679 615
rect 627 543 679 581
rect 627 509 636 543
rect 670 509 679 543
rect 627 471 679 509
rect 627 459 636 471
rect 670 459 679 471
rect 627 399 679 407
rect 627 395 636 399
rect 670 395 679 399
rect 627 331 679 343
rect 627 267 679 279
rect 627 209 679 215
rect 782 759 841 771
rect 782 725 788 759
rect 822 725 841 759
rect 782 687 841 725
rect 782 653 788 687
rect 822 653 841 687
rect 782 615 841 653
rect 782 581 788 615
rect 822 581 841 615
rect 782 543 841 581
rect 782 509 788 543
rect 822 509 841 543
rect 782 471 841 509
rect 782 437 788 471
rect 822 437 841 471
rect 782 399 841 437
rect 782 365 788 399
rect 822 365 841 399
rect 782 327 841 365
rect 782 293 788 327
rect 822 293 841 327
rect 782 255 841 293
rect 782 221 788 255
rect 822 221 841 255
rect 782 209 841 221
rect 264 125 618 137
rect 264 19 280 125
rect 602 19 618 125
rect 264 0 618 19
<< via1 >>
rect 203 437 212 459
rect 212 437 246 459
rect 246 437 255 459
rect 203 407 255 437
rect 203 365 212 395
rect 212 365 246 395
rect 246 365 255 395
rect 203 343 255 365
rect 203 327 255 331
rect 203 293 212 327
rect 212 293 246 327
rect 246 293 255 327
rect 203 279 255 293
rect 203 255 255 267
rect 203 221 212 255
rect 212 221 246 255
rect 246 221 255 255
rect 203 215 255 221
rect 309 759 361 765
rect 309 725 318 759
rect 318 725 352 759
rect 352 725 361 759
rect 309 713 361 725
rect 309 687 361 701
rect 309 653 318 687
rect 318 653 352 687
rect 352 653 361 687
rect 309 649 361 653
rect 309 615 361 637
rect 309 585 318 615
rect 318 585 352 615
rect 352 585 361 615
rect 309 543 361 573
rect 309 521 318 543
rect 318 521 352 543
rect 352 521 361 543
rect 415 437 424 459
rect 424 437 458 459
rect 458 437 467 459
rect 415 407 467 437
rect 415 365 424 395
rect 424 365 458 395
rect 458 365 467 395
rect 415 343 467 365
rect 415 327 467 331
rect 415 293 424 327
rect 424 293 458 327
rect 458 293 467 327
rect 415 279 467 293
rect 415 255 467 267
rect 415 221 424 255
rect 424 221 458 255
rect 458 221 467 255
rect 415 215 467 221
rect 521 759 573 765
rect 521 725 530 759
rect 530 725 564 759
rect 564 725 573 759
rect 521 713 573 725
rect 521 687 573 701
rect 521 653 530 687
rect 530 653 564 687
rect 564 653 573 687
rect 521 649 573 653
rect 521 615 573 637
rect 521 585 530 615
rect 530 585 564 615
rect 564 585 573 615
rect 521 543 573 573
rect 521 521 530 543
rect 530 521 564 543
rect 564 521 573 543
rect 627 437 636 459
rect 636 437 670 459
rect 670 437 679 459
rect 627 407 679 437
rect 627 365 636 395
rect 636 365 670 395
rect 670 365 679 395
rect 627 343 679 365
rect 627 327 679 331
rect 627 293 636 327
rect 636 293 670 327
rect 670 293 679 327
rect 627 279 679 293
rect 627 255 679 267
rect 627 221 636 255
rect 636 221 670 255
rect 670 221 679 255
rect 627 215 679 221
<< metal2 >>
rect 14 765 868 771
rect 14 713 309 765
rect 361 713 521 765
rect 573 713 868 765
rect 14 701 868 713
rect 14 649 309 701
rect 361 649 521 701
rect 573 649 868 701
rect 14 637 868 649
rect 14 585 309 637
rect 361 585 521 637
rect 573 585 868 637
rect 14 573 868 585
rect 14 521 309 573
rect 361 521 521 573
rect 573 521 868 573
rect 14 515 868 521
rect 14 459 868 465
rect 14 407 203 459
rect 255 407 415 459
rect 467 407 627 459
rect 679 407 868 459
rect 14 395 868 407
rect 14 343 203 395
rect 255 343 415 395
rect 467 343 627 395
rect 679 343 868 395
rect 14 331 868 343
rect 14 279 203 331
rect 255 279 415 331
rect 467 279 627 331
rect 679 279 868 331
rect 14 267 868 279
rect 14 215 203 267
rect 255 215 415 267
rect 467 215 627 267
rect 679 215 868 267
rect 14 209 868 215
<< labels >>
flabel metal1 s 321 42 571 92 0 FreeSans 200 0 0 0 GATE
port 2 nsew
flabel metal1 s 321 878 571 928 0 FreeSans 200 0 0 0 GATE
port 2 nsew
flabel metal1 s 41 466 100 496 0 FreeSans 200 90 0 0 SUBSTRATE
port 4 nsew
flabel metal1 s 782 469 841 499 0 FreeSans 200 90 0 0 SUBSTRATE
port 4 nsew
flabel comment s 693 502 693 502 0 FreeSans 180 90 0 0 dummy_poly
flabel comment s 182 502 182 502 0 FreeSans 180 90 0 0 dummy_poly
flabel comment s 269 490 269 490 0 FreeSans 300 0 0 0 S
flabel comment s 355 490 355 490 0 FreeSans 300 0 0 0 S
flabel comment s 441 490 441 490 0 FreeSans 300 0 0 0 S
flabel comment s 527 490 527 490 0 FreeSans 300 0 0 0 S
flabel comment s 269 490 269 490 0 FreeSans 300 0 0 0 S
flabel comment s 355 490 355 490 0 FreeSans 300 0 0 0 D
flabel comment s 441 490 441 490 0 FreeSans 300 0 0 0 S
flabel comment s 527 490 527 490 0 FreeSans 300 0 0 0 D
flabel comment s 613 490 613 490 0 FreeSans 300 0 0 0 S
flabel metal2 s 14 280 35 408 7 FreeSans 300 180 0 0 SOURCE
port 3 nsew
flabel metal2 s 14 589 35 717 7 FreeSans 300 180 0 0 DRAIN
port 1 nsew
<< properties >>
string GDS_END 6467638
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_pr/gds/sky130_fd_pr.gds
string GDS_START 6446684
<< end >>
