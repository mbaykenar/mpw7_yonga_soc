magic
tech sky130B
magscale 12 1
timestamp 1598765253
<< metal5 >>
rect 0 90 45 105
rect 0 60 15 90
rect 0 45 30 60
rect 0 0 15 45
<< properties >>
string FIXED_BBOX 0 -30 60 105
<< end >>
