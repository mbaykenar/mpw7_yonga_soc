magic
tech sky130A
magscale 1 2
timestamp 1649977179
<< nwell >>
rect -38 261 2890 582
<< pwell >>
rect 37 157 1011 203
rect 37 21 2834 157
rect 37 17 64 21
rect 30 -17 64 17
rect 1041 -17 1075 21
<< locali >>
rect 17 215 123 264
rect 1475 347 1520 492
rect 1640 347 1692 492
rect 1812 347 1864 492
rect 1984 347 2036 492
rect 2153 347 2205 492
rect 2325 347 2377 492
rect 2497 347 2549 492
rect 1475 344 2549 347
rect 2671 344 2729 492
rect 1475 299 2817 344
rect 652 215 940 255
rect 2584 181 2817 299
rect 1468 147 2817 181
rect 1468 56 1520 147
rect 1640 56 1692 147
rect 1812 56 1864 147
rect 1981 56 2036 147
rect 2153 56 2205 147
rect 2325 56 2377 147
rect 2497 56 2549 147
rect 2671 56 2723 147
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2053 561
rect 2087 527 2145 561
rect 2179 527 2237 561
rect 2271 527 2329 561
rect 2363 527 2421 561
rect 2455 527 2513 561
rect 2547 527 2605 561
rect 2639 527 2697 561
rect 2731 527 2789 561
rect 2823 527 2852 561
rect 26 299 107 527
rect 141 315 207 493
rect 241 459 653 493
rect 241 315 317 459
rect 351 349 385 425
rect 419 387 485 459
rect 519 349 553 425
rect 157 255 207 315
rect 351 289 553 349
rect 587 333 653 459
rect 687 367 737 527
rect 771 333 805 493
rect 839 367 905 527
rect 939 333 995 493
rect 587 291 995 333
rect 1031 459 1097 493
rect 1031 425 1047 459
rect 1081 425 1097 459
rect 1031 299 1097 425
rect 157 215 453 255
rect 49 17 107 181
rect 157 163 207 215
rect 487 193 553 289
rect 1131 265 1169 493
rect 1203 459 1269 493
rect 1203 425 1219 459
rect 1253 425 1269 459
rect 1203 299 1269 425
rect 1303 265 1341 492
rect 1375 459 1441 493
rect 1375 425 1390 459
rect 1424 425 1441 459
rect 1375 299 1441 425
rect 1554 459 1606 493
rect 1554 425 1560 459
rect 1594 425 1606 459
rect 1554 381 1606 425
rect 1726 459 1778 493
rect 1726 425 1736 459
rect 1770 425 1778 459
rect 1726 381 1778 425
rect 1898 459 1950 493
rect 1898 425 1908 459
rect 1942 425 1950 459
rect 1898 381 1950 425
rect 2070 459 2119 493
rect 2070 425 2079 459
rect 2113 425 2119 459
rect 2070 381 2119 425
rect 2242 459 2291 493
rect 2242 425 2251 459
rect 2285 425 2291 459
rect 2242 381 2291 425
rect 2414 459 2463 493
rect 2414 425 2422 459
rect 2456 425 2463 459
rect 2414 381 2463 425
rect 2586 459 2637 493
rect 2586 425 2592 459
rect 2626 425 2637 459
rect 2586 381 2637 425
rect 2763 459 2817 493
rect 2763 425 2768 459
rect 2802 425 2817 459
rect 2763 378 2817 425
rect 487 181 619 193
rect 141 51 207 163
rect 243 17 301 181
rect 335 145 905 181
rect 335 51 401 145
rect 435 17 469 111
rect 503 51 569 145
rect 603 17 637 111
rect 671 51 737 145
rect 771 17 805 111
rect 839 51 905 145
rect 939 113 995 181
rect 1029 147 1092 265
rect 1131 215 2550 265
rect 939 17 1090 113
rect 1131 53 1176 215
rect 1210 17 1262 122
rect 1298 53 1348 215
rect 1382 17 1434 129
rect 1554 17 1606 113
rect 1726 17 1778 113
rect 1898 17 1947 113
rect 2070 17 2119 113
rect 2241 17 2291 113
rect 2413 17 2463 113
rect 2585 17 2637 113
rect 2757 17 2817 113
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2053 17
rect 2087 -17 2145 17
rect 2179 -17 2237 17
rect 2271 -17 2329 17
rect 2363 -17 2421 17
rect 2455 -17 2513 17
rect 2547 -17 2605 17
rect 2639 -17 2697 17
rect 2731 -17 2789 17
rect 2823 -17 2852 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 1593 527 1627 561
rect 1685 527 1719 561
rect 1777 527 1811 561
rect 1869 527 1903 561
rect 1961 527 1995 561
rect 2053 527 2087 561
rect 2145 527 2179 561
rect 2237 527 2271 561
rect 2329 527 2363 561
rect 2421 527 2455 561
rect 2513 527 2547 561
rect 2605 527 2639 561
rect 2697 527 2731 561
rect 2789 527 2823 561
rect 1047 425 1081 459
rect 1219 425 1253 459
rect 1390 425 1424 459
rect 1560 425 1594 459
rect 1736 425 1770 459
rect 1908 425 1942 459
rect 2079 425 2113 459
rect 2251 425 2285 459
rect 2422 425 2456 459
rect 2592 425 2626 459
rect 2768 425 2802 459
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1593 -17 1627 17
rect 1685 -17 1719 17
rect 1777 -17 1811 17
rect 1869 -17 1903 17
rect 1961 -17 1995 17
rect 2053 -17 2087 17
rect 2145 -17 2179 17
rect 2237 -17 2271 17
rect 2329 -17 2363 17
rect 2421 -17 2455 17
rect 2513 -17 2547 17
rect 2605 -17 2639 17
rect 2697 -17 2731 17
rect 2789 -17 2823 17
<< metal1 >>
rect 0 561 2852 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2053 561
rect 2087 527 2145 561
rect 2179 527 2237 561
rect 2271 527 2329 561
rect 2363 527 2421 561
rect 2455 527 2513 561
rect 2547 527 2605 561
rect 2639 527 2697 561
rect 2731 527 2789 561
rect 2823 527 2852 561
rect 0 496 2852 527
rect 14 459 2838 468
rect 14 428 1047 459
rect 1035 425 1047 428
rect 1081 428 1219 459
rect 1081 425 1093 428
rect 1035 416 1093 425
rect 1207 425 1219 428
rect 1253 428 1390 459
rect 1253 425 1265 428
rect 1207 416 1265 425
rect 1378 425 1390 428
rect 1424 428 1560 459
rect 1424 425 1436 428
rect 1378 416 1436 425
rect 1548 425 1560 428
rect 1594 428 1736 459
rect 1594 425 1606 428
rect 1548 416 1606 425
rect 1724 425 1736 428
rect 1770 428 1908 459
rect 1770 425 1782 428
rect 1724 416 1782 425
rect 1896 425 1908 428
rect 1942 428 2079 459
rect 1942 425 1954 428
rect 1896 416 1954 425
rect 2067 425 2079 428
rect 2113 428 2251 459
rect 2113 425 2125 428
rect 2067 416 2125 425
rect 2239 425 2251 428
rect 2285 428 2422 459
rect 2285 425 2297 428
rect 2239 416 2297 425
rect 2410 425 2422 428
rect 2456 428 2592 459
rect 2456 425 2468 428
rect 2410 416 2468 425
rect 2580 425 2592 428
rect 2626 428 2768 459
rect 2626 425 2638 428
rect 2580 416 2638 425
rect 2756 425 2768 428
rect 2802 428 2838 459
rect 2802 425 2814 428
rect 2756 416 2814 425
rect 0 17 2852 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2053 17
rect 2087 -17 2145 17
rect 2179 -17 2237 17
rect 2271 -17 2329 17
rect 2363 -17 2421 17
rect 2455 -17 2513 17
rect 2547 -17 2605 17
rect 2639 -17 2697 17
rect 2731 -17 2789 17
rect 2823 -17 2852 17
rect 0 -48 2852 -17
<< obsm1 >>
rect 493 184 623 193
rect 1030 184 1088 193
rect 493 156 1088 184
rect 493 147 623 156
rect 1030 147 1088 156
<< labels >>
rlabel locali s 17 215 123 264 6 A
port 1 nsew signal input
rlabel locali s 652 215 940 255 6 SLEEP
port 2 nsew signal input
rlabel metal1 s 2756 416 2814 428 6 KAPWR
port 3 nsew power bidirectional abutment
rlabel metal1 s 2580 416 2638 428 6 KAPWR
port 3 nsew power bidirectional abutment
rlabel metal1 s 2410 416 2468 428 6 KAPWR
port 3 nsew power bidirectional abutment
rlabel metal1 s 2239 416 2297 428 6 KAPWR
port 3 nsew power bidirectional abutment
rlabel metal1 s 2067 416 2125 428 6 KAPWR
port 3 nsew power bidirectional abutment
rlabel metal1 s 1896 416 1954 428 6 KAPWR
port 3 nsew power bidirectional abutment
rlabel metal1 s 1724 416 1782 428 6 KAPWR
port 3 nsew power bidirectional abutment
rlabel metal1 s 1548 416 1606 428 6 KAPWR
port 3 nsew power bidirectional abutment
rlabel metal1 s 1378 416 1436 428 6 KAPWR
port 3 nsew power bidirectional abutment
rlabel metal1 s 1207 416 1265 428 6 KAPWR
port 3 nsew power bidirectional abutment
rlabel metal1 s 1035 416 1093 428 6 KAPWR
port 3 nsew power bidirectional abutment
rlabel metal1 s 14 428 2838 468 6 KAPWR
port 3 nsew power bidirectional abutment
rlabel metal1 s 0 -48 2852 48 8 VGND
port 4 nsew ground bidirectional abutment
rlabel pwell s 1041 -17 1075 21 6 VNB
port 5 nsew ground bidirectional
rlabel pwell s 30 -17 64 17 8 VNB
port 5 nsew ground bidirectional
rlabel pwell s 37 17 64 21 6 VNB
port 5 nsew ground bidirectional
rlabel pwell s 37 21 2834 157 6 VNB
port 5 nsew ground bidirectional
rlabel pwell s 37 157 1011 203 6 VNB
port 5 nsew ground bidirectional
rlabel nwell s -38 261 2890 582 6 VPB
port 6 nsew power bidirectional
rlabel metal1 s 0 496 2852 592 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 2671 56 2723 147 6 X
port 8 nsew signal output
rlabel locali s 2497 56 2549 147 6 X
port 8 nsew signal output
rlabel locali s 2325 56 2377 147 6 X
port 8 nsew signal output
rlabel locali s 2153 56 2205 147 6 X
port 8 nsew signal output
rlabel locali s 1981 56 2036 147 6 X
port 8 nsew signal output
rlabel locali s 1812 56 1864 147 6 X
port 8 nsew signal output
rlabel locali s 1640 56 1692 147 6 X
port 8 nsew signal output
rlabel locali s 1468 56 1520 147 6 X
port 8 nsew signal output
rlabel locali s 1468 147 2817 181 6 X
port 8 nsew signal output
rlabel locali s 2584 181 2817 299 6 X
port 8 nsew signal output
rlabel locali s 1475 299 2817 344 6 X
port 8 nsew signal output
rlabel locali s 2671 344 2729 492 6 X
port 8 nsew signal output
rlabel locali s 1475 344 2549 347 6 X
port 8 nsew signal output
rlabel locali s 2497 347 2549 492 6 X
port 8 nsew signal output
rlabel locali s 2325 347 2377 492 6 X
port 8 nsew signal output
rlabel locali s 2153 347 2205 492 6 X
port 8 nsew signal output
rlabel locali s 1984 347 2036 492 6 X
port 8 nsew signal output
rlabel locali s 1812 347 1864 492 6 X
port 8 nsew signal output
rlabel locali s 1640 347 1692 492 6 X
port 8 nsew signal output
rlabel locali s 1475 347 1520 492 6 X
port 8 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 2852 544
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_END 2444532
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 2422616
<< end >>
