magic
tech sky130B
magscale 12 1
timestamp 1598769216
<< metal5 >>
rect 0 55 15 105
rect 30 55 45 105
rect 60 55 75 105
rect 0 45 75 55
rect 5 30 70 45
rect 10 15 65 30
rect 15 0 30 15
rect 45 0 60 15
<< properties >>
string FIXED_BBOX 0 -30 90 105
<< end >>
