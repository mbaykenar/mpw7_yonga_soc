magic
tech sky130B
timestamp 1649977179
<< properties >>
string GDS_END 3201280
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 3200636
<< end >>
