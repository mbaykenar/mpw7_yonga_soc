magic
tech sky130B
magscale 1 2
timestamp 1649977179
<< dnwell >>
rect 1822 1724 134872 81473
<< nwell >>
rect 1738 81389 134956 81557
rect 1738 1808 1906 81389
rect 134788 1808 134956 81389
rect 1738 1640 134956 1808
<< nsubdiff >>
rect 2133 81490 2183 81514
rect 2133 81456 2141 81490
rect 2175 81456 2183 81490
rect 2133 81432 2183 81456
rect 2469 81490 2519 81514
rect 2469 81456 2477 81490
rect 2511 81456 2519 81490
rect 2469 81432 2519 81456
rect 2805 81490 2855 81514
rect 2805 81456 2813 81490
rect 2847 81456 2855 81490
rect 2805 81432 2855 81456
rect 3141 81490 3191 81514
rect 3141 81456 3149 81490
rect 3183 81456 3191 81490
rect 3141 81432 3191 81456
rect 3477 81490 3527 81514
rect 3477 81456 3485 81490
rect 3519 81456 3527 81490
rect 3477 81432 3527 81456
rect 3813 81490 3863 81514
rect 3813 81456 3821 81490
rect 3855 81456 3863 81490
rect 3813 81432 3863 81456
rect 4149 81490 4199 81514
rect 4149 81456 4157 81490
rect 4191 81456 4199 81490
rect 4149 81432 4199 81456
rect 4485 81490 4535 81514
rect 4485 81456 4493 81490
rect 4527 81456 4535 81490
rect 4485 81432 4535 81456
rect 4821 81490 4871 81514
rect 4821 81456 4829 81490
rect 4863 81456 4871 81490
rect 4821 81432 4871 81456
rect 5157 81490 5207 81514
rect 5157 81456 5165 81490
rect 5199 81456 5207 81490
rect 5157 81432 5207 81456
rect 5493 81490 5543 81514
rect 5493 81456 5501 81490
rect 5535 81456 5543 81490
rect 5493 81432 5543 81456
rect 5829 81490 5879 81514
rect 5829 81456 5837 81490
rect 5871 81456 5879 81490
rect 5829 81432 5879 81456
rect 6165 81490 6215 81514
rect 6165 81456 6173 81490
rect 6207 81456 6215 81490
rect 6165 81432 6215 81456
rect 6501 81490 6551 81514
rect 6501 81456 6509 81490
rect 6543 81456 6551 81490
rect 6501 81432 6551 81456
rect 6837 81490 6887 81514
rect 6837 81456 6845 81490
rect 6879 81456 6887 81490
rect 6837 81432 6887 81456
rect 7173 81490 7223 81514
rect 7173 81456 7181 81490
rect 7215 81456 7223 81490
rect 7173 81432 7223 81456
rect 7509 81490 7559 81514
rect 7509 81456 7517 81490
rect 7551 81456 7559 81490
rect 7509 81432 7559 81456
rect 7845 81490 7895 81514
rect 7845 81456 7853 81490
rect 7887 81456 7895 81490
rect 7845 81432 7895 81456
rect 8181 81490 8231 81514
rect 8181 81456 8189 81490
rect 8223 81456 8231 81490
rect 8181 81432 8231 81456
rect 8517 81490 8567 81514
rect 8517 81456 8525 81490
rect 8559 81456 8567 81490
rect 8517 81432 8567 81456
rect 8853 81490 8903 81514
rect 8853 81456 8861 81490
rect 8895 81456 8903 81490
rect 8853 81432 8903 81456
rect 9189 81490 9239 81514
rect 9189 81456 9197 81490
rect 9231 81456 9239 81490
rect 9189 81432 9239 81456
rect 9525 81490 9575 81514
rect 9525 81456 9533 81490
rect 9567 81456 9575 81490
rect 9525 81432 9575 81456
rect 9861 81490 9911 81514
rect 9861 81456 9869 81490
rect 9903 81456 9911 81490
rect 9861 81432 9911 81456
rect 10197 81490 10247 81514
rect 10197 81456 10205 81490
rect 10239 81456 10247 81490
rect 10197 81432 10247 81456
rect 10533 81490 10583 81514
rect 10533 81456 10541 81490
rect 10575 81456 10583 81490
rect 10533 81432 10583 81456
rect 10869 81490 10919 81514
rect 10869 81456 10877 81490
rect 10911 81456 10919 81490
rect 10869 81432 10919 81456
rect 11205 81490 11255 81514
rect 11205 81456 11213 81490
rect 11247 81456 11255 81490
rect 11205 81432 11255 81456
rect 11541 81490 11591 81514
rect 11541 81456 11549 81490
rect 11583 81456 11591 81490
rect 11541 81432 11591 81456
rect 11877 81490 11927 81514
rect 11877 81456 11885 81490
rect 11919 81456 11927 81490
rect 11877 81432 11927 81456
rect 12213 81490 12263 81514
rect 12213 81456 12221 81490
rect 12255 81456 12263 81490
rect 12213 81432 12263 81456
rect 12549 81490 12599 81514
rect 12549 81456 12557 81490
rect 12591 81456 12599 81490
rect 12549 81432 12599 81456
rect 12885 81490 12935 81514
rect 12885 81456 12893 81490
rect 12927 81456 12935 81490
rect 12885 81432 12935 81456
rect 13221 81490 13271 81514
rect 13221 81456 13229 81490
rect 13263 81456 13271 81490
rect 13221 81432 13271 81456
rect 13557 81490 13607 81514
rect 13557 81456 13565 81490
rect 13599 81456 13607 81490
rect 13557 81432 13607 81456
rect 13893 81490 13943 81514
rect 13893 81456 13901 81490
rect 13935 81456 13943 81490
rect 13893 81432 13943 81456
rect 14229 81490 14279 81514
rect 14229 81456 14237 81490
rect 14271 81456 14279 81490
rect 14229 81432 14279 81456
rect 14565 81490 14615 81514
rect 14565 81456 14573 81490
rect 14607 81456 14615 81490
rect 14565 81432 14615 81456
rect 14901 81490 14951 81514
rect 14901 81456 14909 81490
rect 14943 81456 14951 81490
rect 14901 81432 14951 81456
rect 15237 81490 15287 81514
rect 15237 81456 15245 81490
rect 15279 81456 15287 81490
rect 15237 81432 15287 81456
rect 15573 81490 15623 81514
rect 15573 81456 15581 81490
rect 15615 81456 15623 81490
rect 15573 81432 15623 81456
rect 15909 81490 15959 81514
rect 15909 81456 15917 81490
rect 15951 81456 15959 81490
rect 15909 81432 15959 81456
rect 16245 81490 16295 81514
rect 16245 81456 16253 81490
rect 16287 81456 16295 81490
rect 16245 81432 16295 81456
rect 16581 81490 16631 81514
rect 16581 81456 16589 81490
rect 16623 81456 16631 81490
rect 16581 81432 16631 81456
rect 16917 81490 16967 81514
rect 16917 81456 16925 81490
rect 16959 81456 16967 81490
rect 16917 81432 16967 81456
rect 17253 81490 17303 81514
rect 17253 81456 17261 81490
rect 17295 81456 17303 81490
rect 17253 81432 17303 81456
rect 17589 81490 17639 81514
rect 17589 81456 17597 81490
rect 17631 81456 17639 81490
rect 17589 81432 17639 81456
rect 17925 81490 17975 81514
rect 17925 81456 17933 81490
rect 17967 81456 17975 81490
rect 17925 81432 17975 81456
rect 18261 81490 18311 81514
rect 18261 81456 18269 81490
rect 18303 81456 18311 81490
rect 18261 81432 18311 81456
rect 18597 81490 18647 81514
rect 18597 81456 18605 81490
rect 18639 81456 18647 81490
rect 18597 81432 18647 81456
rect 18933 81490 18983 81514
rect 18933 81456 18941 81490
rect 18975 81456 18983 81490
rect 18933 81432 18983 81456
rect 19269 81490 19319 81514
rect 19269 81456 19277 81490
rect 19311 81456 19319 81490
rect 19269 81432 19319 81456
rect 19605 81490 19655 81514
rect 19605 81456 19613 81490
rect 19647 81456 19655 81490
rect 19605 81432 19655 81456
rect 19941 81490 19991 81514
rect 19941 81456 19949 81490
rect 19983 81456 19991 81490
rect 19941 81432 19991 81456
rect 20277 81490 20327 81514
rect 20277 81456 20285 81490
rect 20319 81456 20327 81490
rect 20277 81432 20327 81456
rect 20613 81490 20663 81514
rect 20613 81456 20621 81490
rect 20655 81456 20663 81490
rect 20613 81432 20663 81456
rect 20949 81490 20999 81514
rect 20949 81456 20957 81490
rect 20991 81456 20999 81490
rect 20949 81432 20999 81456
rect 21285 81490 21335 81514
rect 21285 81456 21293 81490
rect 21327 81456 21335 81490
rect 21285 81432 21335 81456
rect 21621 81490 21671 81514
rect 21621 81456 21629 81490
rect 21663 81456 21671 81490
rect 21621 81432 21671 81456
rect 21957 81490 22007 81514
rect 21957 81456 21965 81490
rect 21999 81456 22007 81490
rect 21957 81432 22007 81456
rect 22293 81490 22343 81514
rect 22293 81456 22301 81490
rect 22335 81456 22343 81490
rect 22293 81432 22343 81456
rect 22629 81490 22679 81514
rect 22629 81456 22637 81490
rect 22671 81456 22679 81490
rect 22629 81432 22679 81456
rect 22965 81490 23015 81514
rect 22965 81456 22973 81490
rect 23007 81456 23015 81490
rect 22965 81432 23015 81456
rect 23301 81490 23351 81514
rect 23301 81456 23309 81490
rect 23343 81456 23351 81490
rect 23301 81432 23351 81456
rect 23637 81490 23687 81514
rect 23637 81456 23645 81490
rect 23679 81456 23687 81490
rect 23637 81432 23687 81456
rect 23973 81490 24023 81514
rect 23973 81456 23981 81490
rect 24015 81456 24023 81490
rect 23973 81432 24023 81456
rect 24309 81490 24359 81514
rect 24309 81456 24317 81490
rect 24351 81456 24359 81490
rect 24309 81432 24359 81456
rect 24645 81490 24695 81514
rect 24645 81456 24653 81490
rect 24687 81456 24695 81490
rect 24645 81432 24695 81456
rect 24981 81490 25031 81514
rect 24981 81456 24989 81490
rect 25023 81456 25031 81490
rect 24981 81432 25031 81456
rect 25317 81490 25367 81514
rect 25317 81456 25325 81490
rect 25359 81456 25367 81490
rect 25317 81432 25367 81456
rect 25653 81490 25703 81514
rect 25653 81456 25661 81490
rect 25695 81456 25703 81490
rect 25653 81432 25703 81456
rect 25989 81490 26039 81514
rect 25989 81456 25997 81490
rect 26031 81456 26039 81490
rect 25989 81432 26039 81456
rect 26325 81490 26375 81514
rect 26325 81456 26333 81490
rect 26367 81456 26375 81490
rect 26325 81432 26375 81456
rect 26661 81490 26711 81514
rect 26661 81456 26669 81490
rect 26703 81456 26711 81490
rect 26661 81432 26711 81456
rect 26997 81490 27047 81514
rect 26997 81456 27005 81490
rect 27039 81456 27047 81490
rect 26997 81432 27047 81456
rect 27333 81490 27383 81514
rect 27333 81456 27341 81490
rect 27375 81456 27383 81490
rect 27333 81432 27383 81456
rect 27669 81490 27719 81514
rect 27669 81456 27677 81490
rect 27711 81456 27719 81490
rect 27669 81432 27719 81456
rect 28005 81490 28055 81514
rect 28005 81456 28013 81490
rect 28047 81456 28055 81490
rect 28005 81432 28055 81456
rect 28341 81490 28391 81514
rect 28341 81456 28349 81490
rect 28383 81456 28391 81490
rect 28341 81432 28391 81456
rect 28677 81490 28727 81514
rect 28677 81456 28685 81490
rect 28719 81456 28727 81490
rect 28677 81432 28727 81456
rect 29013 81490 29063 81514
rect 29013 81456 29021 81490
rect 29055 81456 29063 81490
rect 29013 81432 29063 81456
rect 29349 81490 29399 81514
rect 29349 81456 29357 81490
rect 29391 81456 29399 81490
rect 29349 81432 29399 81456
rect 29685 81490 29735 81514
rect 29685 81456 29693 81490
rect 29727 81456 29735 81490
rect 29685 81432 29735 81456
rect 30021 81490 30071 81514
rect 30021 81456 30029 81490
rect 30063 81456 30071 81490
rect 30021 81432 30071 81456
rect 30357 81490 30407 81514
rect 30357 81456 30365 81490
rect 30399 81456 30407 81490
rect 30357 81432 30407 81456
rect 30693 81490 30743 81514
rect 30693 81456 30701 81490
rect 30735 81456 30743 81490
rect 30693 81432 30743 81456
rect 31029 81490 31079 81514
rect 31029 81456 31037 81490
rect 31071 81456 31079 81490
rect 31029 81432 31079 81456
rect 31365 81490 31415 81514
rect 31365 81456 31373 81490
rect 31407 81456 31415 81490
rect 31365 81432 31415 81456
rect 31701 81490 31751 81514
rect 31701 81456 31709 81490
rect 31743 81456 31751 81490
rect 31701 81432 31751 81456
rect 32037 81490 32087 81514
rect 32037 81456 32045 81490
rect 32079 81456 32087 81490
rect 32037 81432 32087 81456
rect 32373 81490 32423 81514
rect 32373 81456 32381 81490
rect 32415 81456 32423 81490
rect 32373 81432 32423 81456
rect 32709 81490 32759 81514
rect 32709 81456 32717 81490
rect 32751 81456 32759 81490
rect 32709 81432 32759 81456
rect 33045 81490 33095 81514
rect 33045 81456 33053 81490
rect 33087 81456 33095 81490
rect 33045 81432 33095 81456
rect 33381 81490 33431 81514
rect 33381 81456 33389 81490
rect 33423 81456 33431 81490
rect 33381 81432 33431 81456
rect 33717 81490 33767 81514
rect 33717 81456 33725 81490
rect 33759 81456 33767 81490
rect 33717 81432 33767 81456
rect 34053 81490 34103 81514
rect 34053 81456 34061 81490
rect 34095 81456 34103 81490
rect 34053 81432 34103 81456
rect 34389 81490 34439 81514
rect 34389 81456 34397 81490
rect 34431 81456 34439 81490
rect 34389 81432 34439 81456
rect 34725 81490 34775 81514
rect 34725 81456 34733 81490
rect 34767 81456 34775 81490
rect 34725 81432 34775 81456
rect 35061 81490 35111 81514
rect 35061 81456 35069 81490
rect 35103 81456 35111 81490
rect 35061 81432 35111 81456
rect 35397 81490 35447 81514
rect 35397 81456 35405 81490
rect 35439 81456 35447 81490
rect 35397 81432 35447 81456
rect 35733 81490 35783 81514
rect 35733 81456 35741 81490
rect 35775 81456 35783 81490
rect 35733 81432 35783 81456
rect 36069 81490 36119 81514
rect 36069 81456 36077 81490
rect 36111 81456 36119 81490
rect 36069 81432 36119 81456
rect 36405 81490 36455 81514
rect 36405 81456 36413 81490
rect 36447 81456 36455 81490
rect 36405 81432 36455 81456
rect 36741 81490 36791 81514
rect 36741 81456 36749 81490
rect 36783 81456 36791 81490
rect 36741 81432 36791 81456
rect 37077 81490 37127 81514
rect 37077 81456 37085 81490
rect 37119 81456 37127 81490
rect 37077 81432 37127 81456
rect 37413 81490 37463 81514
rect 37413 81456 37421 81490
rect 37455 81456 37463 81490
rect 37413 81432 37463 81456
rect 37749 81490 37799 81514
rect 37749 81456 37757 81490
rect 37791 81456 37799 81490
rect 37749 81432 37799 81456
rect 38085 81490 38135 81514
rect 38085 81456 38093 81490
rect 38127 81456 38135 81490
rect 38085 81432 38135 81456
rect 38421 81490 38471 81514
rect 38421 81456 38429 81490
rect 38463 81456 38471 81490
rect 38421 81432 38471 81456
rect 38757 81490 38807 81514
rect 38757 81456 38765 81490
rect 38799 81456 38807 81490
rect 38757 81432 38807 81456
rect 39093 81490 39143 81514
rect 39093 81456 39101 81490
rect 39135 81456 39143 81490
rect 39093 81432 39143 81456
rect 39429 81490 39479 81514
rect 39429 81456 39437 81490
rect 39471 81456 39479 81490
rect 39429 81432 39479 81456
rect 39765 81490 39815 81514
rect 39765 81456 39773 81490
rect 39807 81456 39815 81490
rect 39765 81432 39815 81456
rect 40101 81490 40151 81514
rect 40101 81456 40109 81490
rect 40143 81456 40151 81490
rect 40101 81432 40151 81456
rect 40437 81490 40487 81514
rect 40437 81456 40445 81490
rect 40479 81456 40487 81490
rect 40437 81432 40487 81456
rect 40773 81490 40823 81514
rect 40773 81456 40781 81490
rect 40815 81456 40823 81490
rect 40773 81432 40823 81456
rect 41109 81490 41159 81514
rect 41109 81456 41117 81490
rect 41151 81456 41159 81490
rect 41109 81432 41159 81456
rect 41445 81490 41495 81514
rect 41445 81456 41453 81490
rect 41487 81456 41495 81490
rect 41445 81432 41495 81456
rect 41781 81490 41831 81514
rect 41781 81456 41789 81490
rect 41823 81456 41831 81490
rect 41781 81432 41831 81456
rect 42117 81490 42167 81514
rect 42117 81456 42125 81490
rect 42159 81456 42167 81490
rect 42117 81432 42167 81456
rect 42453 81490 42503 81514
rect 42453 81456 42461 81490
rect 42495 81456 42503 81490
rect 42453 81432 42503 81456
rect 42789 81490 42839 81514
rect 42789 81456 42797 81490
rect 42831 81456 42839 81490
rect 42789 81432 42839 81456
rect 43125 81490 43175 81514
rect 43125 81456 43133 81490
rect 43167 81456 43175 81490
rect 43125 81432 43175 81456
rect 43461 81490 43511 81514
rect 43461 81456 43469 81490
rect 43503 81456 43511 81490
rect 43461 81432 43511 81456
rect 43797 81490 43847 81514
rect 43797 81456 43805 81490
rect 43839 81456 43847 81490
rect 43797 81432 43847 81456
rect 44133 81490 44183 81514
rect 44133 81456 44141 81490
rect 44175 81456 44183 81490
rect 44133 81432 44183 81456
rect 44469 81490 44519 81514
rect 44469 81456 44477 81490
rect 44511 81456 44519 81490
rect 44469 81432 44519 81456
rect 44805 81490 44855 81514
rect 44805 81456 44813 81490
rect 44847 81456 44855 81490
rect 44805 81432 44855 81456
rect 45141 81490 45191 81514
rect 45141 81456 45149 81490
rect 45183 81456 45191 81490
rect 45141 81432 45191 81456
rect 45477 81490 45527 81514
rect 45477 81456 45485 81490
rect 45519 81456 45527 81490
rect 45477 81432 45527 81456
rect 45813 81490 45863 81514
rect 45813 81456 45821 81490
rect 45855 81456 45863 81490
rect 45813 81432 45863 81456
rect 46149 81490 46199 81514
rect 46149 81456 46157 81490
rect 46191 81456 46199 81490
rect 46149 81432 46199 81456
rect 46485 81490 46535 81514
rect 46485 81456 46493 81490
rect 46527 81456 46535 81490
rect 46485 81432 46535 81456
rect 46821 81490 46871 81514
rect 46821 81456 46829 81490
rect 46863 81456 46871 81490
rect 46821 81432 46871 81456
rect 47157 81490 47207 81514
rect 47157 81456 47165 81490
rect 47199 81456 47207 81490
rect 47157 81432 47207 81456
rect 47493 81490 47543 81514
rect 47493 81456 47501 81490
rect 47535 81456 47543 81490
rect 47493 81432 47543 81456
rect 47829 81490 47879 81514
rect 47829 81456 47837 81490
rect 47871 81456 47879 81490
rect 47829 81432 47879 81456
rect 48165 81490 48215 81514
rect 48165 81456 48173 81490
rect 48207 81456 48215 81490
rect 48165 81432 48215 81456
rect 48501 81490 48551 81514
rect 48501 81456 48509 81490
rect 48543 81456 48551 81490
rect 48501 81432 48551 81456
rect 48837 81490 48887 81514
rect 48837 81456 48845 81490
rect 48879 81456 48887 81490
rect 48837 81432 48887 81456
rect 49173 81490 49223 81514
rect 49173 81456 49181 81490
rect 49215 81456 49223 81490
rect 49173 81432 49223 81456
rect 49509 81490 49559 81514
rect 49509 81456 49517 81490
rect 49551 81456 49559 81490
rect 49509 81432 49559 81456
rect 49845 81490 49895 81514
rect 49845 81456 49853 81490
rect 49887 81456 49895 81490
rect 49845 81432 49895 81456
rect 50181 81490 50231 81514
rect 50181 81456 50189 81490
rect 50223 81456 50231 81490
rect 50181 81432 50231 81456
rect 50517 81490 50567 81514
rect 50517 81456 50525 81490
rect 50559 81456 50567 81490
rect 50517 81432 50567 81456
rect 50853 81490 50903 81514
rect 50853 81456 50861 81490
rect 50895 81456 50903 81490
rect 50853 81432 50903 81456
rect 51189 81490 51239 81514
rect 51189 81456 51197 81490
rect 51231 81456 51239 81490
rect 51189 81432 51239 81456
rect 51525 81490 51575 81514
rect 51525 81456 51533 81490
rect 51567 81456 51575 81490
rect 51525 81432 51575 81456
rect 51861 81490 51911 81514
rect 51861 81456 51869 81490
rect 51903 81456 51911 81490
rect 51861 81432 51911 81456
rect 52197 81490 52247 81514
rect 52197 81456 52205 81490
rect 52239 81456 52247 81490
rect 52197 81432 52247 81456
rect 52533 81490 52583 81514
rect 52533 81456 52541 81490
rect 52575 81456 52583 81490
rect 52533 81432 52583 81456
rect 52869 81490 52919 81514
rect 52869 81456 52877 81490
rect 52911 81456 52919 81490
rect 52869 81432 52919 81456
rect 53205 81490 53255 81514
rect 53205 81456 53213 81490
rect 53247 81456 53255 81490
rect 53205 81432 53255 81456
rect 53541 81490 53591 81514
rect 53541 81456 53549 81490
rect 53583 81456 53591 81490
rect 53541 81432 53591 81456
rect 53877 81490 53927 81514
rect 53877 81456 53885 81490
rect 53919 81456 53927 81490
rect 53877 81432 53927 81456
rect 54213 81490 54263 81514
rect 54213 81456 54221 81490
rect 54255 81456 54263 81490
rect 54213 81432 54263 81456
rect 54549 81490 54599 81514
rect 54549 81456 54557 81490
rect 54591 81456 54599 81490
rect 54549 81432 54599 81456
rect 54885 81490 54935 81514
rect 54885 81456 54893 81490
rect 54927 81456 54935 81490
rect 54885 81432 54935 81456
rect 55221 81490 55271 81514
rect 55221 81456 55229 81490
rect 55263 81456 55271 81490
rect 55221 81432 55271 81456
rect 55557 81490 55607 81514
rect 55557 81456 55565 81490
rect 55599 81456 55607 81490
rect 55557 81432 55607 81456
rect 55893 81490 55943 81514
rect 55893 81456 55901 81490
rect 55935 81456 55943 81490
rect 55893 81432 55943 81456
rect 56229 81490 56279 81514
rect 56229 81456 56237 81490
rect 56271 81456 56279 81490
rect 56229 81432 56279 81456
rect 56565 81490 56615 81514
rect 56565 81456 56573 81490
rect 56607 81456 56615 81490
rect 56565 81432 56615 81456
rect 56901 81490 56951 81514
rect 56901 81456 56909 81490
rect 56943 81456 56951 81490
rect 56901 81432 56951 81456
rect 57237 81490 57287 81514
rect 57237 81456 57245 81490
rect 57279 81456 57287 81490
rect 57237 81432 57287 81456
rect 57573 81490 57623 81514
rect 57573 81456 57581 81490
rect 57615 81456 57623 81490
rect 57573 81432 57623 81456
rect 57909 81490 57959 81514
rect 57909 81456 57917 81490
rect 57951 81456 57959 81490
rect 57909 81432 57959 81456
rect 58245 81490 58295 81514
rect 58245 81456 58253 81490
rect 58287 81456 58295 81490
rect 58245 81432 58295 81456
rect 58581 81490 58631 81514
rect 58581 81456 58589 81490
rect 58623 81456 58631 81490
rect 58581 81432 58631 81456
rect 58917 81490 58967 81514
rect 58917 81456 58925 81490
rect 58959 81456 58967 81490
rect 58917 81432 58967 81456
rect 59253 81490 59303 81514
rect 59253 81456 59261 81490
rect 59295 81456 59303 81490
rect 59253 81432 59303 81456
rect 59589 81490 59639 81514
rect 59589 81456 59597 81490
rect 59631 81456 59639 81490
rect 59589 81432 59639 81456
rect 59925 81490 59975 81514
rect 59925 81456 59933 81490
rect 59967 81456 59975 81490
rect 59925 81432 59975 81456
rect 60261 81490 60311 81514
rect 60261 81456 60269 81490
rect 60303 81456 60311 81490
rect 60261 81432 60311 81456
rect 60597 81490 60647 81514
rect 60597 81456 60605 81490
rect 60639 81456 60647 81490
rect 60597 81432 60647 81456
rect 60933 81490 60983 81514
rect 60933 81456 60941 81490
rect 60975 81456 60983 81490
rect 60933 81432 60983 81456
rect 61269 81490 61319 81514
rect 61269 81456 61277 81490
rect 61311 81456 61319 81490
rect 61269 81432 61319 81456
rect 61605 81490 61655 81514
rect 61605 81456 61613 81490
rect 61647 81456 61655 81490
rect 61605 81432 61655 81456
rect 61941 81490 61991 81514
rect 61941 81456 61949 81490
rect 61983 81456 61991 81490
rect 61941 81432 61991 81456
rect 62277 81490 62327 81514
rect 62277 81456 62285 81490
rect 62319 81456 62327 81490
rect 62277 81432 62327 81456
rect 62613 81490 62663 81514
rect 62613 81456 62621 81490
rect 62655 81456 62663 81490
rect 62613 81432 62663 81456
rect 62949 81490 62999 81514
rect 62949 81456 62957 81490
rect 62991 81456 62999 81490
rect 62949 81432 62999 81456
rect 63285 81490 63335 81514
rect 63285 81456 63293 81490
rect 63327 81456 63335 81490
rect 63285 81432 63335 81456
rect 63621 81490 63671 81514
rect 63621 81456 63629 81490
rect 63663 81456 63671 81490
rect 63621 81432 63671 81456
rect 63957 81490 64007 81514
rect 63957 81456 63965 81490
rect 63999 81456 64007 81490
rect 63957 81432 64007 81456
rect 64293 81490 64343 81514
rect 64293 81456 64301 81490
rect 64335 81456 64343 81490
rect 64293 81432 64343 81456
rect 64629 81490 64679 81514
rect 64629 81456 64637 81490
rect 64671 81456 64679 81490
rect 64629 81432 64679 81456
rect 64965 81490 65015 81514
rect 64965 81456 64973 81490
rect 65007 81456 65015 81490
rect 64965 81432 65015 81456
rect 65301 81490 65351 81514
rect 65301 81456 65309 81490
rect 65343 81456 65351 81490
rect 65301 81432 65351 81456
rect 65637 81490 65687 81514
rect 65637 81456 65645 81490
rect 65679 81456 65687 81490
rect 65637 81432 65687 81456
rect 65973 81490 66023 81514
rect 65973 81456 65981 81490
rect 66015 81456 66023 81490
rect 65973 81432 66023 81456
rect 66309 81490 66359 81514
rect 66309 81456 66317 81490
rect 66351 81456 66359 81490
rect 66309 81432 66359 81456
rect 66645 81490 66695 81514
rect 66645 81456 66653 81490
rect 66687 81456 66695 81490
rect 66645 81432 66695 81456
rect 66981 81490 67031 81514
rect 66981 81456 66989 81490
rect 67023 81456 67031 81490
rect 66981 81432 67031 81456
rect 67317 81490 67367 81514
rect 67317 81456 67325 81490
rect 67359 81456 67367 81490
rect 67317 81432 67367 81456
rect 67653 81490 67703 81514
rect 67653 81456 67661 81490
rect 67695 81456 67703 81490
rect 67653 81432 67703 81456
rect 67989 81490 68039 81514
rect 67989 81456 67997 81490
rect 68031 81456 68039 81490
rect 67989 81432 68039 81456
rect 68325 81490 68375 81514
rect 68325 81456 68333 81490
rect 68367 81456 68375 81490
rect 68325 81432 68375 81456
rect 68661 81490 68711 81514
rect 68661 81456 68669 81490
rect 68703 81456 68711 81490
rect 68661 81432 68711 81456
rect 68997 81490 69047 81514
rect 68997 81456 69005 81490
rect 69039 81456 69047 81490
rect 68997 81432 69047 81456
rect 69333 81490 69383 81514
rect 69333 81456 69341 81490
rect 69375 81456 69383 81490
rect 69333 81432 69383 81456
rect 69669 81490 69719 81514
rect 69669 81456 69677 81490
rect 69711 81456 69719 81490
rect 69669 81432 69719 81456
rect 70005 81490 70055 81514
rect 70005 81456 70013 81490
rect 70047 81456 70055 81490
rect 70005 81432 70055 81456
rect 70341 81490 70391 81514
rect 70341 81456 70349 81490
rect 70383 81456 70391 81490
rect 70341 81432 70391 81456
rect 70677 81490 70727 81514
rect 70677 81456 70685 81490
rect 70719 81456 70727 81490
rect 70677 81432 70727 81456
rect 71013 81490 71063 81514
rect 71013 81456 71021 81490
rect 71055 81456 71063 81490
rect 71013 81432 71063 81456
rect 71349 81490 71399 81514
rect 71349 81456 71357 81490
rect 71391 81456 71399 81490
rect 71349 81432 71399 81456
rect 71685 81490 71735 81514
rect 71685 81456 71693 81490
rect 71727 81456 71735 81490
rect 71685 81432 71735 81456
rect 72021 81490 72071 81514
rect 72021 81456 72029 81490
rect 72063 81456 72071 81490
rect 72021 81432 72071 81456
rect 72357 81490 72407 81514
rect 72357 81456 72365 81490
rect 72399 81456 72407 81490
rect 72357 81432 72407 81456
rect 72693 81490 72743 81514
rect 72693 81456 72701 81490
rect 72735 81456 72743 81490
rect 72693 81432 72743 81456
rect 73029 81490 73079 81514
rect 73029 81456 73037 81490
rect 73071 81456 73079 81490
rect 73029 81432 73079 81456
rect 73365 81490 73415 81514
rect 73365 81456 73373 81490
rect 73407 81456 73415 81490
rect 73365 81432 73415 81456
rect 73701 81490 73751 81514
rect 73701 81456 73709 81490
rect 73743 81456 73751 81490
rect 73701 81432 73751 81456
rect 74037 81490 74087 81514
rect 74037 81456 74045 81490
rect 74079 81456 74087 81490
rect 74037 81432 74087 81456
rect 74373 81490 74423 81514
rect 74373 81456 74381 81490
rect 74415 81456 74423 81490
rect 74373 81432 74423 81456
rect 74709 81490 74759 81514
rect 74709 81456 74717 81490
rect 74751 81456 74759 81490
rect 74709 81432 74759 81456
rect 75045 81490 75095 81514
rect 75045 81456 75053 81490
rect 75087 81456 75095 81490
rect 75045 81432 75095 81456
rect 75381 81490 75431 81514
rect 75381 81456 75389 81490
rect 75423 81456 75431 81490
rect 75381 81432 75431 81456
rect 75717 81490 75767 81514
rect 75717 81456 75725 81490
rect 75759 81456 75767 81490
rect 75717 81432 75767 81456
rect 76053 81490 76103 81514
rect 76053 81456 76061 81490
rect 76095 81456 76103 81490
rect 76053 81432 76103 81456
rect 76389 81490 76439 81514
rect 76389 81456 76397 81490
rect 76431 81456 76439 81490
rect 76389 81432 76439 81456
rect 76725 81490 76775 81514
rect 76725 81456 76733 81490
rect 76767 81456 76775 81490
rect 76725 81432 76775 81456
rect 77061 81490 77111 81514
rect 77061 81456 77069 81490
rect 77103 81456 77111 81490
rect 77061 81432 77111 81456
rect 77397 81490 77447 81514
rect 77397 81456 77405 81490
rect 77439 81456 77447 81490
rect 77397 81432 77447 81456
rect 77733 81490 77783 81514
rect 77733 81456 77741 81490
rect 77775 81456 77783 81490
rect 77733 81432 77783 81456
rect 78069 81490 78119 81514
rect 78069 81456 78077 81490
rect 78111 81456 78119 81490
rect 78069 81432 78119 81456
rect 78405 81490 78455 81514
rect 78405 81456 78413 81490
rect 78447 81456 78455 81490
rect 78405 81432 78455 81456
rect 78741 81490 78791 81514
rect 78741 81456 78749 81490
rect 78783 81456 78791 81490
rect 78741 81432 78791 81456
rect 79077 81490 79127 81514
rect 79077 81456 79085 81490
rect 79119 81456 79127 81490
rect 79077 81432 79127 81456
rect 79413 81490 79463 81514
rect 79413 81456 79421 81490
rect 79455 81456 79463 81490
rect 79413 81432 79463 81456
rect 79749 81490 79799 81514
rect 79749 81456 79757 81490
rect 79791 81456 79799 81490
rect 79749 81432 79799 81456
rect 80085 81490 80135 81514
rect 80085 81456 80093 81490
rect 80127 81456 80135 81490
rect 80085 81432 80135 81456
rect 80421 81490 80471 81514
rect 80421 81456 80429 81490
rect 80463 81456 80471 81490
rect 80421 81432 80471 81456
rect 80757 81490 80807 81514
rect 80757 81456 80765 81490
rect 80799 81456 80807 81490
rect 80757 81432 80807 81456
rect 81093 81490 81143 81514
rect 81093 81456 81101 81490
rect 81135 81456 81143 81490
rect 81093 81432 81143 81456
rect 81429 81490 81479 81514
rect 81429 81456 81437 81490
rect 81471 81456 81479 81490
rect 81429 81432 81479 81456
rect 81765 81490 81815 81514
rect 81765 81456 81773 81490
rect 81807 81456 81815 81490
rect 81765 81432 81815 81456
rect 82101 81490 82151 81514
rect 82101 81456 82109 81490
rect 82143 81456 82151 81490
rect 82101 81432 82151 81456
rect 82437 81490 82487 81514
rect 82437 81456 82445 81490
rect 82479 81456 82487 81490
rect 82437 81432 82487 81456
rect 82773 81490 82823 81514
rect 82773 81456 82781 81490
rect 82815 81456 82823 81490
rect 82773 81432 82823 81456
rect 83109 81490 83159 81514
rect 83109 81456 83117 81490
rect 83151 81456 83159 81490
rect 83109 81432 83159 81456
rect 83445 81490 83495 81514
rect 83445 81456 83453 81490
rect 83487 81456 83495 81490
rect 83445 81432 83495 81456
rect 83781 81490 83831 81514
rect 83781 81456 83789 81490
rect 83823 81456 83831 81490
rect 83781 81432 83831 81456
rect 84117 81490 84167 81514
rect 84117 81456 84125 81490
rect 84159 81456 84167 81490
rect 84117 81432 84167 81456
rect 84453 81490 84503 81514
rect 84453 81456 84461 81490
rect 84495 81456 84503 81490
rect 84453 81432 84503 81456
rect 84789 81490 84839 81514
rect 84789 81456 84797 81490
rect 84831 81456 84839 81490
rect 84789 81432 84839 81456
rect 85125 81490 85175 81514
rect 85125 81456 85133 81490
rect 85167 81456 85175 81490
rect 85125 81432 85175 81456
rect 85461 81490 85511 81514
rect 85461 81456 85469 81490
rect 85503 81456 85511 81490
rect 85461 81432 85511 81456
rect 85797 81490 85847 81514
rect 85797 81456 85805 81490
rect 85839 81456 85847 81490
rect 85797 81432 85847 81456
rect 86133 81490 86183 81514
rect 86133 81456 86141 81490
rect 86175 81456 86183 81490
rect 86133 81432 86183 81456
rect 86469 81490 86519 81514
rect 86469 81456 86477 81490
rect 86511 81456 86519 81490
rect 86469 81432 86519 81456
rect 86805 81490 86855 81514
rect 86805 81456 86813 81490
rect 86847 81456 86855 81490
rect 86805 81432 86855 81456
rect 87141 81490 87191 81514
rect 87141 81456 87149 81490
rect 87183 81456 87191 81490
rect 87141 81432 87191 81456
rect 87477 81490 87527 81514
rect 87477 81456 87485 81490
rect 87519 81456 87527 81490
rect 87477 81432 87527 81456
rect 87813 81490 87863 81514
rect 87813 81456 87821 81490
rect 87855 81456 87863 81490
rect 87813 81432 87863 81456
rect 88149 81490 88199 81514
rect 88149 81456 88157 81490
rect 88191 81456 88199 81490
rect 88149 81432 88199 81456
rect 88485 81490 88535 81514
rect 88485 81456 88493 81490
rect 88527 81456 88535 81490
rect 88485 81432 88535 81456
rect 88821 81490 88871 81514
rect 88821 81456 88829 81490
rect 88863 81456 88871 81490
rect 88821 81432 88871 81456
rect 89157 81490 89207 81514
rect 89157 81456 89165 81490
rect 89199 81456 89207 81490
rect 89157 81432 89207 81456
rect 89493 81490 89543 81514
rect 89493 81456 89501 81490
rect 89535 81456 89543 81490
rect 89493 81432 89543 81456
rect 89829 81490 89879 81514
rect 89829 81456 89837 81490
rect 89871 81456 89879 81490
rect 89829 81432 89879 81456
rect 90165 81490 90215 81514
rect 90165 81456 90173 81490
rect 90207 81456 90215 81490
rect 90165 81432 90215 81456
rect 90501 81490 90551 81514
rect 90501 81456 90509 81490
rect 90543 81456 90551 81490
rect 90501 81432 90551 81456
rect 90837 81490 90887 81514
rect 90837 81456 90845 81490
rect 90879 81456 90887 81490
rect 90837 81432 90887 81456
rect 91173 81490 91223 81514
rect 91173 81456 91181 81490
rect 91215 81456 91223 81490
rect 91173 81432 91223 81456
rect 91509 81490 91559 81514
rect 91509 81456 91517 81490
rect 91551 81456 91559 81490
rect 91509 81432 91559 81456
rect 91845 81490 91895 81514
rect 91845 81456 91853 81490
rect 91887 81456 91895 81490
rect 91845 81432 91895 81456
rect 92181 81490 92231 81514
rect 92181 81456 92189 81490
rect 92223 81456 92231 81490
rect 92181 81432 92231 81456
rect 92517 81490 92567 81514
rect 92517 81456 92525 81490
rect 92559 81456 92567 81490
rect 92517 81432 92567 81456
rect 92853 81490 92903 81514
rect 92853 81456 92861 81490
rect 92895 81456 92903 81490
rect 92853 81432 92903 81456
rect 93189 81490 93239 81514
rect 93189 81456 93197 81490
rect 93231 81456 93239 81490
rect 93189 81432 93239 81456
rect 93525 81490 93575 81514
rect 93525 81456 93533 81490
rect 93567 81456 93575 81490
rect 93525 81432 93575 81456
rect 93861 81490 93911 81514
rect 93861 81456 93869 81490
rect 93903 81456 93911 81490
rect 93861 81432 93911 81456
rect 94197 81490 94247 81514
rect 94197 81456 94205 81490
rect 94239 81456 94247 81490
rect 94197 81432 94247 81456
rect 94533 81490 94583 81514
rect 94533 81456 94541 81490
rect 94575 81456 94583 81490
rect 94533 81432 94583 81456
rect 94869 81490 94919 81514
rect 94869 81456 94877 81490
rect 94911 81456 94919 81490
rect 94869 81432 94919 81456
rect 95205 81490 95255 81514
rect 95205 81456 95213 81490
rect 95247 81456 95255 81490
rect 95205 81432 95255 81456
rect 95541 81490 95591 81514
rect 95541 81456 95549 81490
rect 95583 81456 95591 81490
rect 95541 81432 95591 81456
rect 95877 81490 95927 81514
rect 95877 81456 95885 81490
rect 95919 81456 95927 81490
rect 95877 81432 95927 81456
rect 96213 81490 96263 81514
rect 96213 81456 96221 81490
rect 96255 81456 96263 81490
rect 96213 81432 96263 81456
rect 96549 81490 96599 81514
rect 96549 81456 96557 81490
rect 96591 81456 96599 81490
rect 96549 81432 96599 81456
rect 96885 81490 96935 81514
rect 96885 81456 96893 81490
rect 96927 81456 96935 81490
rect 96885 81432 96935 81456
rect 97221 81490 97271 81514
rect 97221 81456 97229 81490
rect 97263 81456 97271 81490
rect 97221 81432 97271 81456
rect 97557 81490 97607 81514
rect 97557 81456 97565 81490
rect 97599 81456 97607 81490
rect 97557 81432 97607 81456
rect 97893 81490 97943 81514
rect 97893 81456 97901 81490
rect 97935 81456 97943 81490
rect 97893 81432 97943 81456
rect 98229 81490 98279 81514
rect 98229 81456 98237 81490
rect 98271 81456 98279 81490
rect 98229 81432 98279 81456
rect 98565 81490 98615 81514
rect 98565 81456 98573 81490
rect 98607 81456 98615 81490
rect 98565 81432 98615 81456
rect 98901 81490 98951 81514
rect 98901 81456 98909 81490
rect 98943 81456 98951 81490
rect 98901 81432 98951 81456
rect 99237 81490 99287 81514
rect 99237 81456 99245 81490
rect 99279 81456 99287 81490
rect 99237 81432 99287 81456
rect 99573 81490 99623 81514
rect 99573 81456 99581 81490
rect 99615 81456 99623 81490
rect 99573 81432 99623 81456
rect 99909 81490 99959 81514
rect 99909 81456 99917 81490
rect 99951 81456 99959 81490
rect 99909 81432 99959 81456
rect 100245 81490 100295 81514
rect 100245 81456 100253 81490
rect 100287 81456 100295 81490
rect 100245 81432 100295 81456
rect 100581 81490 100631 81514
rect 100581 81456 100589 81490
rect 100623 81456 100631 81490
rect 100581 81432 100631 81456
rect 100917 81490 100967 81514
rect 100917 81456 100925 81490
rect 100959 81456 100967 81490
rect 100917 81432 100967 81456
rect 101253 81490 101303 81514
rect 101253 81456 101261 81490
rect 101295 81456 101303 81490
rect 101253 81432 101303 81456
rect 101589 81490 101639 81514
rect 101589 81456 101597 81490
rect 101631 81456 101639 81490
rect 101589 81432 101639 81456
rect 101925 81490 101975 81514
rect 101925 81456 101933 81490
rect 101967 81456 101975 81490
rect 101925 81432 101975 81456
rect 102261 81490 102311 81514
rect 102261 81456 102269 81490
rect 102303 81456 102311 81490
rect 102261 81432 102311 81456
rect 102597 81490 102647 81514
rect 102597 81456 102605 81490
rect 102639 81456 102647 81490
rect 102597 81432 102647 81456
rect 102933 81490 102983 81514
rect 102933 81456 102941 81490
rect 102975 81456 102983 81490
rect 102933 81432 102983 81456
rect 103269 81490 103319 81514
rect 103269 81456 103277 81490
rect 103311 81456 103319 81490
rect 103269 81432 103319 81456
rect 103605 81490 103655 81514
rect 103605 81456 103613 81490
rect 103647 81456 103655 81490
rect 103605 81432 103655 81456
rect 103941 81490 103991 81514
rect 103941 81456 103949 81490
rect 103983 81456 103991 81490
rect 103941 81432 103991 81456
rect 104277 81490 104327 81514
rect 104277 81456 104285 81490
rect 104319 81456 104327 81490
rect 104277 81432 104327 81456
rect 104613 81490 104663 81514
rect 104613 81456 104621 81490
rect 104655 81456 104663 81490
rect 104613 81432 104663 81456
rect 104949 81490 104999 81514
rect 104949 81456 104957 81490
rect 104991 81456 104999 81490
rect 104949 81432 104999 81456
rect 105285 81490 105335 81514
rect 105285 81456 105293 81490
rect 105327 81456 105335 81490
rect 105285 81432 105335 81456
rect 105621 81490 105671 81514
rect 105621 81456 105629 81490
rect 105663 81456 105671 81490
rect 105621 81432 105671 81456
rect 105957 81490 106007 81514
rect 105957 81456 105965 81490
rect 105999 81456 106007 81490
rect 105957 81432 106007 81456
rect 106293 81490 106343 81514
rect 106293 81456 106301 81490
rect 106335 81456 106343 81490
rect 106293 81432 106343 81456
rect 106629 81490 106679 81514
rect 106629 81456 106637 81490
rect 106671 81456 106679 81490
rect 106629 81432 106679 81456
rect 106965 81490 107015 81514
rect 106965 81456 106973 81490
rect 107007 81456 107015 81490
rect 106965 81432 107015 81456
rect 107301 81490 107351 81514
rect 107301 81456 107309 81490
rect 107343 81456 107351 81490
rect 107301 81432 107351 81456
rect 107637 81490 107687 81514
rect 107637 81456 107645 81490
rect 107679 81456 107687 81490
rect 107637 81432 107687 81456
rect 107973 81490 108023 81514
rect 107973 81456 107981 81490
rect 108015 81456 108023 81490
rect 107973 81432 108023 81456
rect 108309 81490 108359 81514
rect 108309 81456 108317 81490
rect 108351 81456 108359 81490
rect 108309 81432 108359 81456
rect 108645 81490 108695 81514
rect 108645 81456 108653 81490
rect 108687 81456 108695 81490
rect 108645 81432 108695 81456
rect 108981 81490 109031 81514
rect 108981 81456 108989 81490
rect 109023 81456 109031 81490
rect 108981 81432 109031 81456
rect 109317 81490 109367 81514
rect 109317 81456 109325 81490
rect 109359 81456 109367 81490
rect 109317 81432 109367 81456
rect 109653 81490 109703 81514
rect 109653 81456 109661 81490
rect 109695 81456 109703 81490
rect 109653 81432 109703 81456
rect 109989 81490 110039 81514
rect 109989 81456 109997 81490
rect 110031 81456 110039 81490
rect 109989 81432 110039 81456
rect 110325 81490 110375 81514
rect 110325 81456 110333 81490
rect 110367 81456 110375 81490
rect 110325 81432 110375 81456
rect 110661 81490 110711 81514
rect 110661 81456 110669 81490
rect 110703 81456 110711 81490
rect 110661 81432 110711 81456
rect 110997 81490 111047 81514
rect 110997 81456 111005 81490
rect 111039 81456 111047 81490
rect 110997 81432 111047 81456
rect 111333 81490 111383 81514
rect 111333 81456 111341 81490
rect 111375 81456 111383 81490
rect 111333 81432 111383 81456
rect 111669 81490 111719 81514
rect 111669 81456 111677 81490
rect 111711 81456 111719 81490
rect 111669 81432 111719 81456
rect 112005 81490 112055 81514
rect 112005 81456 112013 81490
rect 112047 81456 112055 81490
rect 112005 81432 112055 81456
rect 112341 81490 112391 81514
rect 112341 81456 112349 81490
rect 112383 81456 112391 81490
rect 112341 81432 112391 81456
rect 112677 81490 112727 81514
rect 112677 81456 112685 81490
rect 112719 81456 112727 81490
rect 112677 81432 112727 81456
rect 113013 81490 113063 81514
rect 113013 81456 113021 81490
rect 113055 81456 113063 81490
rect 113013 81432 113063 81456
rect 113349 81490 113399 81514
rect 113349 81456 113357 81490
rect 113391 81456 113399 81490
rect 113349 81432 113399 81456
rect 113685 81490 113735 81514
rect 113685 81456 113693 81490
rect 113727 81456 113735 81490
rect 113685 81432 113735 81456
rect 114021 81490 114071 81514
rect 114021 81456 114029 81490
rect 114063 81456 114071 81490
rect 114021 81432 114071 81456
rect 114357 81490 114407 81514
rect 114357 81456 114365 81490
rect 114399 81456 114407 81490
rect 114357 81432 114407 81456
rect 114693 81490 114743 81514
rect 114693 81456 114701 81490
rect 114735 81456 114743 81490
rect 114693 81432 114743 81456
rect 115029 81490 115079 81514
rect 115029 81456 115037 81490
rect 115071 81456 115079 81490
rect 115029 81432 115079 81456
rect 115365 81490 115415 81514
rect 115365 81456 115373 81490
rect 115407 81456 115415 81490
rect 115365 81432 115415 81456
rect 115701 81490 115751 81514
rect 115701 81456 115709 81490
rect 115743 81456 115751 81490
rect 115701 81432 115751 81456
rect 116037 81490 116087 81514
rect 116037 81456 116045 81490
rect 116079 81456 116087 81490
rect 116037 81432 116087 81456
rect 116373 81490 116423 81514
rect 116373 81456 116381 81490
rect 116415 81456 116423 81490
rect 116373 81432 116423 81456
rect 116709 81490 116759 81514
rect 116709 81456 116717 81490
rect 116751 81456 116759 81490
rect 116709 81432 116759 81456
rect 117045 81490 117095 81514
rect 117045 81456 117053 81490
rect 117087 81456 117095 81490
rect 117045 81432 117095 81456
rect 117381 81490 117431 81514
rect 117381 81456 117389 81490
rect 117423 81456 117431 81490
rect 117381 81432 117431 81456
rect 117717 81490 117767 81514
rect 117717 81456 117725 81490
rect 117759 81456 117767 81490
rect 117717 81432 117767 81456
rect 118053 81490 118103 81514
rect 118053 81456 118061 81490
rect 118095 81456 118103 81490
rect 118053 81432 118103 81456
rect 118389 81490 118439 81514
rect 118389 81456 118397 81490
rect 118431 81456 118439 81490
rect 118389 81432 118439 81456
rect 118725 81490 118775 81514
rect 118725 81456 118733 81490
rect 118767 81456 118775 81490
rect 118725 81432 118775 81456
rect 119061 81490 119111 81514
rect 119061 81456 119069 81490
rect 119103 81456 119111 81490
rect 119061 81432 119111 81456
rect 119397 81490 119447 81514
rect 119397 81456 119405 81490
rect 119439 81456 119447 81490
rect 119397 81432 119447 81456
rect 119733 81490 119783 81514
rect 119733 81456 119741 81490
rect 119775 81456 119783 81490
rect 119733 81432 119783 81456
rect 120069 81490 120119 81514
rect 120069 81456 120077 81490
rect 120111 81456 120119 81490
rect 120069 81432 120119 81456
rect 120405 81490 120455 81514
rect 120405 81456 120413 81490
rect 120447 81456 120455 81490
rect 120405 81432 120455 81456
rect 120741 81490 120791 81514
rect 120741 81456 120749 81490
rect 120783 81456 120791 81490
rect 120741 81432 120791 81456
rect 121077 81490 121127 81514
rect 121077 81456 121085 81490
rect 121119 81456 121127 81490
rect 121077 81432 121127 81456
rect 121413 81490 121463 81514
rect 121413 81456 121421 81490
rect 121455 81456 121463 81490
rect 121413 81432 121463 81456
rect 121749 81490 121799 81514
rect 121749 81456 121757 81490
rect 121791 81456 121799 81490
rect 121749 81432 121799 81456
rect 122085 81490 122135 81514
rect 122085 81456 122093 81490
rect 122127 81456 122135 81490
rect 122085 81432 122135 81456
rect 122421 81490 122471 81514
rect 122421 81456 122429 81490
rect 122463 81456 122471 81490
rect 122421 81432 122471 81456
rect 122757 81490 122807 81514
rect 122757 81456 122765 81490
rect 122799 81456 122807 81490
rect 122757 81432 122807 81456
rect 123093 81490 123143 81514
rect 123093 81456 123101 81490
rect 123135 81456 123143 81490
rect 123093 81432 123143 81456
rect 123429 81490 123479 81514
rect 123429 81456 123437 81490
rect 123471 81456 123479 81490
rect 123429 81432 123479 81456
rect 123765 81490 123815 81514
rect 123765 81456 123773 81490
rect 123807 81456 123815 81490
rect 123765 81432 123815 81456
rect 124101 81490 124151 81514
rect 124101 81456 124109 81490
rect 124143 81456 124151 81490
rect 124101 81432 124151 81456
rect 124437 81490 124487 81514
rect 124437 81456 124445 81490
rect 124479 81456 124487 81490
rect 124437 81432 124487 81456
rect 124773 81490 124823 81514
rect 124773 81456 124781 81490
rect 124815 81456 124823 81490
rect 124773 81432 124823 81456
rect 125109 81490 125159 81514
rect 125109 81456 125117 81490
rect 125151 81456 125159 81490
rect 125109 81432 125159 81456
rect 125445 81490 125495 81514
rect 125445 81456 125453 81490
rect 125487 81456 125495 81490
rect 125445 81432 125495 81456
rect 125781 81490 125831 81514
rect 125781 81456 125789 81490
rect 125823 81456 125831 81490
rect 125781 81432 125831 81456
rect 126117 81490 126167 81514
rect 126117 81456 126125 81490
rect 126159 81456 126167 81490
rect 126117 81432 126167 81456
rect 126453 81490 126503 81514
rect 126453 81456 126461 81490
rect 126495 81456 126503 81490
rect 126453 81432 126503 81456
rect 126789 81490 126839 81514
rect 126789 81456 126797 81490
rect 126831 81456 126839 81490
rect 126789 81432 126839 81456
rect 127125 81490 127175 81514
rect 127125 81456 127133 81490
rect 127167 81456 127175 81490
rect 127125 81432 127175 81456
rect 127461 81490 127511 81514
rect 127461 81456 127469 81490
rect 127503 81456 127511 81490
rect 127461 81432 127511 81456
rect 127797 81490 127847 81514
rect 127797 81456 127805 81490
rect 127839 81456 127847 81490
rect 127797 81432 127847 81456
rect 128133 81490 128183 81514
rect 128133 81456 128141 81490
rect 128175 81456 128183 81490
rect 128133 81432 128183 81456
rect 128469 81490 128519 81514
rect 128469 81456 128477 81490
rect 128511 81456 128519 81490
rect 128469 81432 128519 81456
rect 128805 81490 128855 81514
rect 128805 81456 128813 81490
rect 128847 81456 128855 81490
rect 128805 81432 128855 81456
rect 129141 81490 129191 81514
rect 129141 81456 129149 81490
rect 129183 81456 129191 81490
rect 129141 81432 129191 81456
rect 129477 81490 129527 81514
rect 129477 81456 129485 81490
rect 129519 81456 129527 81490
rect 129477 81432 129527 81456
rect 129813 81490 129863 81514
rect 129813 81456 129821 81490
rect 129855 81456 129863 81490
rect 129813 81432 129863 81456
rect 130149 81490 130199 81514
rect 130149 81456 130157 81490
rect 130191 81456 130199 81490
rect 130149 81432 130199 81456
rect 130485 81490 130535 81514
rect 130485 81456 130493 81490
rect 130527 81456 130535 81490
rect 130485 81432 130535 81456
rect 130821 81490 130871 81514
rect 130821 81456 130829 81490
rect 130863 81456 130871 81490
rect 130821 81432 130871 81456
rect 131157 81490 131207 81514
rect 131157 81456 131165 81490
rect 131199 81456 131207 81490
rect 131157 81432 131207 81456
rect 131493 81490 131543 81514
rect 131493 81456 131501 81490
rect 131535 81456 131543 81490
rect 131493 81432 131543 81456
rect 131829 81490 131879 81514
rect 131829 81456 131837 81490
rect 131871 81456 131879 81490
rect 131829 81432 131879 81456
rect 132165 81490 132215 81514
rect 132165 81456 132173 81490
rect 132207 81456 132215 81490
rect 132165 81432 132215 81456
rect 132501 81490 132551 81514
rect 132501 81456 132509 81490
rect 132543 81456 132551 81490
rect 132501 81432 132551 81456
rect 132837 81490 132887 81514
rect 132837 81456 132845 81490
rect 132879 81456 132887 81490
rect 132837 81432 132887 81456
rect 133173 81490 133223 81514
rect 133173 81456 133181 81490
rect 133215 81456 133223 81490
rect 133173 81432 133223 81456
rect 133509 81490 133559 81514
rect 133509 81456 133517 81490
rect 133551 81456 133559 81490
rect 133509 81432 133559 81456
rect 133845 81490 133895 81514
rect 133845 81456 133853 81490
rect 133887 81456 133895 81490
rect 133845 81432 133895 81456
rect 134181 81490 134231 81514
rect 134181 81456 134189 81490
rect 134223 81456 134231 81490
rect 134181 81432 134231 81456
rect 1797 81037 1847 81061
rect 1797 81003 1805 81037
rect 1839 81003 1847 81037
rect 1797 80979 1847 81003
rect 134847 81037 134897 81061
rect 134847 81003 134855 81037
rect 134889 81003 134897 81037
rect 134847 80979 134897 81003
rect 1797 80701 1847 80725
rect 1797 80667 1805 80701
rect 1839 80667 1847 80701
rect 1797 80643 1847 80667
rect 134847 80701 134897 80725
rect 134847 80667 134855 80701
rect 134889 80667 134897 80701
rect 134847 80643 134897 80667
rect 1797 80365 1847 80389
rect 1797 80331 1805 80365
rect 1839 80331 1847 80365
rect 1797 80307 1847 80331
rect 134847 80365 134897 80389
rect 134847 80331 134855 80365
rect 134889 80331 134897 80365
rect 134847 80307 134897 80331
rect 1797 80029 1847 80053
rect 1797 79995 1805 80029
rect 1839 79995 1847 80029
rect 1797 79971 1847 79995
rect 134847 80029 134897 80053
rect 134847 79995 134855 80029
rect 134889 79995 134897 80029
rect 134847 79971 134897 79995
rect 1797 79693 1847 79717
rect 1797 79659 1805 79693
rect 1839 79659 1847 79693
rect 1797 79635 1847 79659
rect 134847 79693 134897 79717
rect 134847 79659 134855 79693
rect 134889 79659 134897 79693
rect 134847 79635 134897 79659
rect 1797 79357 1847 79381
rect 1797 79323 1805 79357
rect 1839 79323 1847 79357
rect 1797 79299 1847 79323
rect 134847 79357 134897 79381
rect 134847 79323 134855 79357
rect 134889 79323 134897 79357
rect 134847 79299 134897 79323
rect 1797 79021 1847 79045
rect 1797 78987 1805 79021
rect 1839 78987 1847 79021
rect 1797 78963 1847 78987
rect 134847 79021 134897 79045
rect 134847 78987 134855 79021
rect 134889 78987 134897 79021
rect 134847 78963 134897 78987
rect 1797 78685 1847 78709
rect 1797 78651 1805 78685
rect 1839 78651 1847 78685
rect 1797 78627 1847 78651
rect 134847 78685 134897 78709
rect 134847 78651 134855 78685
rect 134889 78651 134897 78685
rect 134847 78627 134897 78651
rect 1797 78349 1847 78373
rect 1797 78315 1805 78349
rect 1839 78315 1847 78349
rect 1797 78291 1847 78315
rect 134847 78349 134897 78373
rect 134847 78315 134855 78349
rect 134889 78315 134897 78349
rect 134847 78291 134897 78315
rect 1797 78013 1847 78037
rect 1797 77979 1805 78013
rect 1839 77979 1847 78013
rect 1797 77955 1847 77979
rect 134847 78013 134897 78037
rect 134847 77979 134855 78013
rect 134889 77979 134897 78013
rect 134847 77955 134897 77979
rect 1797 77677 1847 77701
rect 1797 77643 1805 77677
rect 1839 77643 1847 77677
rect 1797 77619 1847 77643
rect 134847 77677 134897 77701
rect 134847 77643 134855 77677
rect 134889 77643 134897 77677
rect 134847 77619 134897 77643
rect 1797 77341 1847 77365
rect 1797 77307 1805 77341
rect 1839 77307 1847 77341
rect 1797 77283 1847 77307
rect 134847 77341 134897 77365
rect 134847 77307 134855 77341
rect 134889 77307 134897 77341
rect 134847 77283 134897 77307
rect 1797 77005 1847 77029
rect 1797 76971 1805 77005
rect 1839 76971 1847 77005
rect 1797 76947 1847 76971
rect 134847 77005 134897 77029
rect 134847 76971 134855 77005
rect 134889 76971 134897 77005
rect 134847 76947 134897 76971
rect 1797 76669 1847 76693
rect 1797 76635 1805 76669
rect 1839 76635 1847 76669
rect 1797 76611 1847 76635
rect 134847 76669 134897 76693
rect 134847 76635 134855 76669
rect 134889 76635 134897 76669
rect 134847 76611 134897 76635
rect 1797 76333 1847 76357
rect 1797 76299 1805 76333
rect 1839 76299 1847 76333
rect 1797 76275 1847 76299
rect 134847 76333 134897 76357
rect 134847 76299 134855 76333
rect 134889 76299 134897 76333
rect 134847 76275 134897 76299
rect 1797 75997 1847 76021
rect 1797 75963 1805 75997
rect 1839 75963 1847 75997
rect 1797 75939 1847 75963
rect 134847 75997 134897 76021
rect 134847 75963 134855 75997
rect 134889 75963 134897 75997
rect 134847 75939 134897 75963
rect 1797 75661 1847 75685
rect 1797 75627 1805 75661
rect 1839 75627 1847 75661
rect 1797 75603 1847 75627
rect 134847 75661 134897 75685
rect 134847 75627 134855 75661
rect 134889 75627 134897 75661
rect 134847 75603 134897 75627
rect 1797 75325 1847 75349
rect 1797 75291 1805 75325
rect 1839 75291 1847 75325
rect 1797 75267 1847 75291
rect 134847 75325 134897 75349
rect 134847 75291 134855 75325
rect 134889 75291 134897 75325
rect 134847 75267 134897 75291
rect 1797 74989 1847 75013
rect 1797 74955 1805 74989
rect 1839 74955 1847 74989
rect 1797 74931 1847 74955
rect 134847 74989 134897 75013
rect 134847 74955 134855 74989
rect 134889 74955 134897 74989
rect 134847 74931 134897 74955
rect 1797 74653 1847 74677
rect 1797 74619 1805 74653
rect 1839 74619 1847 74653
rect 1797 74595 1847 74619
rect 134847 74653 134897 74677
rect 134847 74619 134855 74653
rect 134889 74619 134897 74653
rect 134847 74595 134897 74619
rect 1797 74317 1847 74341
rect 1797 74283 1805 74317
rect 1839 74283 1847 74317
rect 1797 74259 1847 74283
rect 134847 74317 134897 74341
rect 134847 74283 134855 74317
rect 134889 74283 134897 74317
rect 134847 74259 134897 74283
rect 1797 73981 1847 74005
rect 1797 73947 1805 73981
rect 1839 73947 1847 73981
rect 1797 73923 1847 73947
rect 134847 73981 134897 74005
rect 134847 73947 134855 73981
rect 134889 73947 134897 73981
rect 134847 73923 134897 73947
rect 1797 73645 1847 73669
rect 1797 73611 1805 73645
rect 1839 73611 1847 73645
rect 1797 73587 1847 73611
rect 134847 73645 134897 73669
rect 134847 73611 134855 73645
rect 134889 73611 134897 73645
rect 134847 73587 134897 73611
rect 1797 73309 1847 73333
rect 1797 73275 1805 73309
rect 1839 73275 1847 73309
rect 1797 73251 1847 73275
rect 134847 73309 134897 73333
rect 134847 73275 134855 73309
rect 134889 73275 134897 73309
rect 134847 73251 134897 73275
rect 1797 72973 1847 72997
rect 1797 72939 1805 72973
rect 1839 72939 1847 72973
rect 1797 72915 1847 72939
rect 134847 72973 134897 72997
rect 134847 72939 134855 72973
rect 134889 72939 134897 72973
rect 134847 72915 134897 72939
rect 1797 72637 1847 72661
rect 1797 72603 1805 72637
rect 1839 72603 1847 72637
rect 1797 72579 1847 72603
rect 134847 72637 134897 72661
rect 134847 72603 134855 72637
rect 134889 72603 134897 72637
rect 134847 72579 134897 72603
rect 1797 72301 1847 72325
rect 1797 72267 1805 72301
rect 1839 72267 1847 72301
rect 1797 72243 1847 72267
rect 134847 72301 134897 72325
rect 134847 72267 134855 72301
rect 134889 72267 134897 72301
rect 134847 72243 134897 72267
rect 1797 71965 1847 71989
rect 1797 71931 1805 71965
rect 1839 71931 1847 71965
rect 1797 71907 1847 71931
rect 134847 71965 134897 71989
rect 134847 71931 134855 71965
rect 134889 71931 134897 71965
rect 134847 71907 134897 71931
rect 1797 71629 1847 71653
rect 1797 71595 1805 71629
rect 1839 71595 1847 71629
rect 1797 71571 1847 71595
rect 134847 71629 134897 71653
rect 134847 71595 134855 71629
rect 134889 71595 134897 71629
rect 134847 71571 134897 71595
rect 1797 71293 1847 71317
rect 1797 71259 1805 71293
rect 1839 71259 1847 71293
rect 1797 71235 1847 71259
rect 134847 71293 134897 71317
rect 134847 71259 134855 71293
rect 134889 71259 134897 71293
rect 134847 71235 134897 71259
rect 1797 70957 1847 70981
rect 1797 70923 1805 70957
rect 1839 70923 1847 70957
rect 1797 70899 1847 70923
rect 134847 70957 134897 70981
rect 134847 70923 134855 70957
rect 134889 70923 134897 70957
rect 134847 70899 134897 70923
rect 1797 70621 1847 70645
rect 1797 70587 1805 70621
rect 1839 70587 1847 70621
rect 1797 70563 1847 70587
rect 134847 70621 134897 70645
rect 134847 70587 134855 70621
rect 134889 70587 134897 70621
rect 134847 70563 134897 70587
rect 1797 70285 1847 70309
rect 1797 70251 1805 70285
rect 1839 70251 1847 70285
rect 1797 70227 1847 70251
rect 134847 70285 134897 70309
rect 134847 70251 134855 70285
rect 134889 70251 134897 70285
rect 134847 70227 134897 70251
rect 1797 69949 1847 69973
rect 1797 69915 1805 69949
rect 1839 69915 1847 69949
rect 1797 69891 1847 69915
rect 134847 69949 134897 69973
rect 134847 69915 134855 69949
rect 134889 69915 134897 69949
rect 134847 69891 134897 69915
rect 1797 69613 1847 69637
rect 1797 69579 1805 69613
rect 1839 69579 1847 69613
rect 1797 69555 1847 69579
rect 134847 69613 134897 69637
rect 134847 69579 134855 69613
rect 134889 69579 134897 69613
rect 134847 69555 134897 69579
rect 1797 69277 1847 69301
rect 1797 69243 1805 69277
rect 1839 69243 1847 69277
rect 1797 69219 1847 69243
rect 134847 69277 134897 69301
rect 134847 69243 134855 69277
rect 134889 69243 134897 69277
rect 134847 69219 134897 69243
rect 1797 68941 1847 68965
rect 1797 68907 1805 68941
rect 1839 68907 1847 68941
rect 1797 68883 1847 68907
rect 134847 68941 134897 68965
rect 134847 68907 134855 68941
rect 134889 68907 134897 68941
rect 134847 68883 134897 68907
rect 1797 68605 1847 68629
rect 1797 68571 1805 68605
rect 1839 68571 1847 68605
rect 1797 68547 1847 68571
rect 134847 68605 134897 68629
rect 134847 68571 134855 68605
rect 134889 68571 134897 68605
rect 134847 68547 134897 68571
rect 1797 68269 1847 68293
rect 1797 68235 1805 68269
rect 1839 68235 1847 68269
rect 1797 68211 1847 68235
rect 134847 68269 134897 68293
rect 134847 68235 134855 68269
rect 134889 68235 134897 68269
rect 134847 68211 134897 68235
rect 1797 67933 1847 67957
rect 1797 67899 1805 67933
rect 1839 67899 1847 67933
rect 1797 67875 1847 67899
rect 134847 67933 134897 67957
rect 134847 67899 134855 67933
rect 134889 67899 134897 67933
rect 134847 67875 134897 67899
rect 1797 67597 1847 67621
rect 1797 67563 1805 67597
rect 1839 67563 1847 67597
rect 1797 67539 1847 67563
rect 134847 67597 134897 67621
rect 134847 67563 134855 67597
rect 134889 67563 134897 67597
rect 134847 67539 134897 67563
rect 1797 67261 1847 67285
rect 1797 67227 1805 67261
rect 1839 67227 1847 67261
rect 1797 67203 1847 67227
rect 134847 67261 134897 67285
rect 134847 67227 134855 67261
rect 134889 67227 134897 67261
rect 134847 67203 134897 67227
rect 1797 66925 1847 66949
rect 1797 66891 1805 66925
rect 1839 66891 1847 66925
rect 1797 66867 1847 66891
rect 134847 66925 134897 66949
rect 134847 66891 134855 66925
rect 134889 66891 134897 66925
rect 134847 66867 134897 66891
rect 1797 66589 1847 66613
rect 1797 66555 1805 66589
rect 1839 66555 1847 66589
rect 1797 66531 1847 66555
rect 134847 66589 134897 66613
rect 134847 66555 134855 66589
rect 134889 66555 134897 66589
rect 134847 66531 134897 66555
rect 1797 66253 1847 66277
rect 1797 66219 1805 66253
rect 1839 66219 1847 66253
rect 1797 66195 1847 66219
rect 134847 66253 134897 66277
rect 134847 66219 134855 66253
rect 134889 66219 134897 66253
rect 134847 66195 134897 66219
rect 1797 65917 1847 65941
rect 1797 65883 1805 65917
rect 1839 65883 1847 65917
rect 1797 65859 1847 65883
rect 134847 65917 134897 65941
rect 134847 65883 134855 65917
rect 134889 65883 134897 65917
rect 134847 65859 134897 65883
rect 1797 65581 1847 65605
rect 1797 65547 1805 65581
rect 1839 65547 1847 65581
rect 1797 65523 1847 65547
rect 134847 65581 134897 65605
rect 134847 65547 134855 65581
rect 134889 65547 134897 65581
rect 134847 65523 134897 65547
rect 1797 65245 1847 65269
rect 1797 65211 1805 65245
rect 1839 65211 1847 65245
rect 1797 65187 1847 65211
rect 134847 65245 134897 65269
rect 134847 65211 134855 65245
rect 134889 65211 134897 65245
rect 134847 65187 134897 65211
rect 1797 64909 1847 64933
rect 1797 64875 1805 64909
rect 1839 64875 1847 64909
rect 1797 64851 1847 64875
rect 134847 64909 134897 64933
rect 134847 64875 134855 64909
rect 134889 64875 134897 64909
rect 134847 64851 134897 64875
rect 1797 64573 1847 64597
rect 1797 64539 1805 64573
rect 1839 64539 1847 64573
rect 1797 64515 1847 64539
rect 134847 64573 134897 64597
rect 134847 64539 134855 64573
rect 134889 64539 134897 64573
rect 134847 64515 134897 64539
rect 1797 64237 1847 64261
rect 1797 64203 1805 64237
rect 1839 64203 1847 64237
rect 1797 64179 1847 64203
rect 134847 64237 134897 64261
rect 134847 64203 134855 64237
rect 134889 64203 134897 64237
rect 134847 64179 134897 64203
rect 1797 63901 1847 63925
rect 1797 63867 1805 63901
rect 1839 63867 1847 63901
rect 1797 63843 1847 63867
rect 134847 63901 134897 63925
rect 134847 63867 134855 63901
rect 134889 63867 134897 63901
rect 134847 63843 134897 63867
rect 1797 63565 1847 63589
rect 1797 63531 1805 63565
rect 1839 63531 1847 63565
rect 1797 63507 1847 63531
rect 134847 63565 134897 63589
rect 134847 63531 134855 63565
rect 134889 63531 134897 63565
rect 134847 63507 134897 63531
rect 1797 63229 1847 63253
rect 1797 63195 1805 63229
rect 1839 63195 1847 63229
rect 1797 63171 1847 63195
rect 134847 63229 134897 63253
rect 134847 63195 134855 63229
rect 134889 63195 134897 63229
rect 134847 63171 134897 63195
rect 1797 62893 1847 62917
rect 1797 62859 1805 62893
rect 1839 62859 1847 62893
rect 1797 62835 1847 62859
rect 134847 62893 134897 62917
rect 134847 62859 134855 62893
rect 134889 62859 134897 62893
rect 134847 62835 134897 62859
rect 1797 62557 1847 62581
rect 1797 62523 1805 62557
rect 1839 62523 1847 62557
rect 1797 62499 1847 62523
rect 134847 62557 134897 62581
rect 134847 62523 134855 62557
rect 134889 62523 134897 62557
rect 134847 62499 134897 62523
rect 1797 62221 1847 62245
rect 1797 62187 1805 62221
rect 1839 62187 1847 62221
rect 1797 62163 1847 62187
rect 134847 62221 134897 62245
rect 134847 62187 134855 62221
rect 134889 62187 134897 62221
rect 134847 62163 134897 62187
rect 1797 61885 1847 61909
rect 1797 61851 1805 61885
rect 1839 61851 1847 61885
rect 1797 61827 1847 61851
rect 134847 61885 134897 61909
rect 134847 61851 134855 61885
rect 134889 61851 134897 61885
rect 134847 61827 134897 61851
rect 1797 61549 1847 61573
rect 1797 61515 1805 61549
rect 1839 61515 1847 61549
rect 1797 61491 1847 61515
rect 134847 61549 134897 61573
rect 134847 61515 134855 61549
rect 134889 61515 134897 61549
rect 134847 61491 134897 61515
rect 1797 61213 1847 61237
rect 1797 61179 1805 61213
rect 1839 61179 1847 61213
rect 1797 61155 1847 61179
rect 134847 61213 134897 61237
rect 134847 61179 134855 61213
rect 134889 61179 134897 61213
rect 134847 61155 134897 61179
rect 1797 60877 1847 60901
rect 1797 60843 1805 60877
rect 1839 60843 1847 60877
rect 1797 60819 1847 60843
rect 134847 60877 134897 60901
rect 134847 60843 134855 60877
rect 134889 60843 134897 60877
rect 134847 60819 134897 60843
rect 1797 60541 1847 60565
rect 1797 60507 1805 60541
rect 1839 60507 1847 60541
rect 1797 60483 1847 60507
rect 134847 60541 134897 60565
rect 134847 60507 134855 60541
rect 134889 60507 134897 60541
rect 134847 60483 134897 60507
rect 1797 60205 1847 60229
rect 1797 60171 1805 60205
rect 1839 60171 1847 60205
rect 1797 60147 1847 60171
rect 134847 60205 134897 60229
rect 134847 60171 134855 60205
rect 134889 60171 134897 60205
rect 134847 60147 134897 60171
rect 1797 59869 1847 59893
rect 1797 59835 1805 59869
rect 1839 59835 1847 59869
rect 1797 59811 1847 59835
rect 134847 59869 134897 59893
rect 134847 59835 134855 59869
rect 134889 59835 134897 59869
rect 134847 59811 134897 59835
rect 1797 59533 1847 59557
rect 1797 59499 1805 59533
rect 1839 59499 1847 59533
rect 1797 59475 1847 59499
rect 134847 59533 134897 59557
rect 134847 59499 134855 59533
rect 134889 59499 134897 59533
rect 134847 59475 134897 59499
rect 1797 59197 1847 59221
rect 1797 59163 1805 59197
rect 1839 59163 1847 59197
rect 1797 59139 1847 59163
rect 134847 59197 134897 59221
rect 134847 59163 134855 59197
rect 134889 59163 134897 59197
rect 134847 59139 134897 59163
rect 1797 58861 1847 58885
rect 1797 58827 1805 58861
rect 1839 58827 1847 58861
rect 1797 58803 1847 58827
rect 134847 58861 134897 58885
rect 134847 58827 134855 58861
rect 134889 58827 134897 58861
rect 134847 58803 134897 58827
rect 1797 58525 1847 58549
rect 1797 58491 1805 58525
rect 1839 58491 1847 58525
rect 1797 58467 1847 58491
rect 134847 58525 134897 58549
rect 134847 58491 134855 58525
rect 134889 58491 134897 58525
rect 134847 58467 134897 58491
rect 1797 58189 1847 58213
rect 1797 58155 1805 58189
rect 1839 58155 1847 58189
rect 1797 58131 1847 58155
rect 134847 58189 134897 58213
rect 134847 58155 134855 58189
rect 134889 58155 134897 58189
rect 134847 58131 134897 58155
rect 1797 57853 1847 57877
rect 1797 57819 1805 57853
rect 1839 57819 1847 57853
rect 1797 57795 1847 57819
rect 134847 57853 134897 57877
rect 134847 57819 134855 57853
rect 134889 57819 134897 57853
rect 134847 57795 134897 57819
rect 1797 57517 1847 57541
rect 1797 57483 1805 57517
rect 1839 57483 1847 57517
rect 1797 57459 1847 57483
rect 134847 57517 134897 57541
rect 134847 57483 134855 57517
rect 134889 57483 134897 57517
rect 134847 57459 134897 57483
rect 1797 57181 1847 57205
rect 1797 57147 1805 57181
rect 1839 57147 1847 57181
rect 1797 57123 1847 57147
rect 134847 57181 134897 57205
rect 134847 57147 134855 57181
rect 134889 57147 134897 57181
rect 134847 57123 134897 57147
rect 1797 56845 1847 56869
rect 1797 56811 1805 56845
rect 1839 56811 1847 56845
rect 1797 56787 1847 56811
rect 134847 56845 134897 56869
rect 134847 56811 134855 56845
rect 134889 56811 134897 56845
rect 134847 56787 134897 56811
rect 1797 56509 1847 56533
rect 1797 56475 1805 56509
rect 1839 56475 1847 56509
rect 1797 56451 1847 56475
rect 134847 56509 134897 56533
rect 134847 56475 134855 56509
rect 134889 56475 134897 56509
rect 134847 56451 134897 56475
rect 1797 56173 1847 56197
rect 1797 56139 1805 56173
rect 1839 56139 1847 56173
rect 1797 56115 1847 56139
rect 134847 56173 134897 56197
rect 134847 56139 134855 56173
rect 134889 56139 134897 56173
rect 134847 56115 134897 56139
rect 1797 55837 1847 55861
rect 1797 55803 1805 55837
rect 1839 55803 1847 55837
rect 1797 55779 1847 55803
rect 134847 55837 134897 55861
rect 134847 55803 134855 55837
rect 134889 55803 134897 55837
rect 134847 55779 134897 55803
rect 1797 55501 1847 55525
rect 1797 55467 1805 55501
rect 1839 55467 1847 55501
rect 1797 55443 1847 55467
rect 134847 55501 134897 55525
rect 134847 55467 134855 55501
rect 134889 55467 134897 55501
rect 134847 55443 134897 55467
rect 1797 55165 1847 55189
rect 1797 55131 1805 55165
rect 1839 55131 1847 55165
rect 1797 55107 1847 55131
rect 134847 55165 134897 55189
rect 134847 55131 134855 55165
rect 134889 55131 134897 55165
rect 134847 55107 134897 55131
rect 1797 54829 1847 54853
rect 1797 54795 1805 54829
rect 1839 54795 1847 54829
rect 1797 54771 1847 54795
rect 134847 54829 134897 54853
rect 134847 54795 134855 54829
rect 134889 54795 134897 54829
rect 134847 54771 134897 54795
rect 1797 54493 1847 54517
rect 1797 54459 1805 54493
rect 1839 54459 1847 54493
rect 1797 54435 1847 54459
rect 134847 54493 134897 54517
rect 134847 54459 134855 54493
rect 134889 54459 134897 54493
rect 134847 54435 134897 54459
rect 1797 54157 1847 54181
rect 1797 54123 1805 54157
rect 1839 54123 1847 54157
rect 1797 54099 1847 54123
rect 134847 54157 134897 54181
rect 134847 54123 134855 54157
rect 134889 54123 134897 54157
rect 134847 54099 134897 54123
rect 1797 53821 1847 53845
rect 1797 53787 1805 53821
rect 1839 53787 1847 53821
rect 1797 53763 1847 53787
rect 134847 53821 134897 53845
rect 134847 53787 134855 53821
rect 134889 53787 134897 53821
rect 134847 53763 134897 53787
rect 1797 53485 1847 53509
rect 1797 53451 1805 53485
rect 1839 53451 1847 53485
rect 1797 53427 1847 53451
rect 134847 53485 134897 53509
rect 134847 53451 134855 53485
rect 134889 53451 134897 53485
rect 134847 53427 134897 53451
rect 1797 53149 1847 53173
rect 1797 53115 1805 53149
rect 1839 53115 1847 53149
rect 1797 53091 1847 53115
rect 134847 53149 134897 53173
rect 134847 53115 134855 53149
rect 134889 53115 134897 53149
rect 134847 53091 134897 53115
rect 1797 52813 1847 52837
rect 1797 52779 1805 52813
rect 1839 52779 1847 52813
rect 1797 52755 1847 52779
rect 134847 52813 134897 52837
rect 134847 52779 134855 52813
rect 134889 52779 134897 52813
rect 134847 52755 134897 52779
rect 1797 52477 1847 52501
rect 1797 52443 1805 52477
rect 1839 52443 1847 52477
rect 1797 52419 1847 52443
rect 134847 52477 134897 52501
rect 134847 52443 134855 52477
rect 134889 52443 134897 52477
rect 134847 52419 134897 52443
rect 1797 52141 1847 52165
rect 1797 52107 1805 52141
rect 1839 52107 1847 52141
rect 1797 52083 1847 52107
rect 134847 52141 134897 52165
rect 134847 52107 134855 52141
rect 134889 52107 134897 52141
rect 134847 52083 134897 52107
rect 1797 51805 1847 51829
rect 1797 51771 1805 51805
rect 1839 51771 1847 51805
rect 1797 51747 1847 51771
rect 134847 51805 134897 51829
rect 134847 51771 134855 51805
rect 134889 51771 134897 51805
rect 134847 51747 134897 51771
rect 1797 51469 1847 51493
rect 1797 51435 1805 51469
rect 1839 51435 1847 51469
rect 1797 51411 1847 51435
rect 134847 51469 134897 51493
rect 134847 51435 134855 51469
rect 134889 51435 134897 51469
rect 134847 51411 134897 51435
rect 1797 51133 1847 51157
rect 1797 51099 1805 51133
rect 1839 51099 1847 51133
rect 1797 51075 1847 51099
rect 134847 51133 134897 51157
rect 134847 51099 134855 51133
rect 134889 51099 134897 51133
rect 134847 51075 134897 51099
rect 1797 50797 1847 50821
rect 1797 50763 1805 50797
rect 1839 50763 1847 50797
rect 1797 50739 1847 50763
rect 134847 50797 134897 50821
rect 134847 50763 134855 50797
rect 134889 50763 134897 50797
rect 134847 50739 134897 50763
rect 1797 50461 1847 50485
rect 1797 50427 1805 50461
rect 1839 50427 1847 50461
rect 1797 50403 1847 50427
rect 134847 50461 134897 50485
rect 134847 50427 134855 50461
rect 134889 50427 134897 50461
rect 134847 50403 134897 50427
rect 1797 50125 1847 50149
rect 1797 50091 1805 50125
rect 1839 50091 1847 50125
rect 1797 50067 1847 50091
rect 134847 50125 134897 50149
rect 134847 50091 134855 50125
rect 134889 50091 134897 50125
rect 134847 50067 134897 50091
rect 1797 49789 1847 49813
rect 1797 49755 1805 49789
rect 1839 49755 1847 49789
rect 1797 49731 1847 49755
rect 134847 49789 134897 49813
rect 134847 49755 134855 49789
rect 134889 49755 134897 49789
rect 134847 49731 134897 49755
rect 1797 49453 1847 49477
rect 1797 49419 1805 49453
rect 1839 49419 1847 49453
rect 1797 49395 1847 49419
rect 134847 49453 134897 49477
rect 134847 49419 134855 49453
rect 134889 49419 134897 49453
rect 134847 49395 134897 49419
rect 1797 49117 1847 49141
rect 1797 49083 1805 49117
rect 1839 49083 1847 49117
rect 1797 49059 1847 49083
rect 134847 49117 134897 49141
rect 134847 49083 134855 49117
rect 134889 49083 134897 49117
rect 134847 49059 134897 49083
rect 1797 48781 1847 48805
rect 1797 48747 1805 48781
rect 1839 48747 1847 48781
rect 1797 48723 1847 48747
rect 134847 48781 134897 48805
rect 134847 48747 134855 48781
rect 134889 48747 134897 48781
rect 134847 48723 134897 48747
rect 1797 48445 1847 48469
rect 1797 48411 1805 48445
rect 1839 48411 1847 48445
rect 1797 48387 1847 48411
rect 134847 48445 134897 48469
rect 134847 48411 134855 48445
rect 134889 48411 134897 48445
rect 134847 48387 134897 48411
rect 1797 48109 1847 48133
rect 1797 48075 1805 48109
rect 1839 48075 1847 48109
rect 1797 48051 1847 48075
rect 134847 48109 134897 48133
rect 134847 48075 134855 48109
rect 134889 48075 134897 48109
rect 134847 48051 134897 48075
rect 1797 47773 1847 47797
rect 1797 47739 1805 47773
rect 1839 47739 1847 47773
rect 1797 47715 1847 47739
rect 134847 47773 134897 47797
rect 134847 47739 134855 47773
rect 134889 47739 134897 47773
rect 134847 47715 134897 47739
rect 1797 47437 1847 47461
rect 1797 47403 1805 47437
rect 1839 47403 1847 47437
rect 1797 47379 1847 47403
rect 134847 47437 134897 47461
rect 134847 47403 134855 47437
rect 134889 47403 134897 47437
rect 134847 47379 134897 47403
rect 1797 47101 1847 47125
rect 1797 47067 1805 47101
rect 1839 47067 1847 47101
rect 1797 47043 1847 47067
rect 134847 47101 134897 47125
rect 134847 47067 134855 47101
rect 134889 47067 134897 47101
rect 134847 47043 134897 47067
rect 1797 46765 1847 46789
rect 1797 46731 1805 46765
rect 1839 46731 1847 46765
rect 1797 46707 1847 46731
rect 134847 46765 134897 46789
rect 134847 46731 134855 46765
rect 134889 46731 134897 46765
rect 134847 46707 134897 46731
rect 1797 46429 1847 46453
rect 1797 46395 1805 46429
rect 1839 46395 1847 46429
rect 1797 46371 1847 46395
rect 134847 46429 134897 46453
rect 134847 46395 134855 46429
rect 134889 46395 134897 46429
rect 134847 46371 134897 46395
rect 1797 46093 1847 46117
rect 1797 46059 1805 46093
rect 1839 46059 1847 46093
rect 1797 46035 1847 46059
rect 134847 46093 134897 46117
rect 134847 46059 134855 46093
rect 134889 46059 134897 46093
rect 134847 46035 134897 46059
rect 1797 45757 1847 45781
rect 1797 45723 1805 45757
rect 1839 45723 1847 45757
rect 1797 45699 1847 45723
rect 134847 45757 134897 45781
rect 134847 45723 134855 45757
rect 134889 45723 134897 45757
rect 134847 45699 134897 45723
rect 1797 45421 1847 45445
rect 1797 45387 1805 45421
rect 1839 45387 1847 45421
rect 1797 45363 1847 45387
rect 134847 45421 134897 45445
rect 134847 45387 134855 45421
rect 134889 45387 134897 45421
rect 134847 45363 134897 45387
rect 1797 45085 1847 45109
rect 1797 45051 1805 45085
rect 1839 45051 1847 45085
rect 1797 45027 1847 45051
rect 134847 45085 134897 45109
rect 134847 45051 134855 45085
rect 134889 45051 134897 45085
rect 134847 45027 134897 45051
rect 1797 44749 1847 44773
rect 1797 44715 1805 44749
rect 1839 44715 1847 44749
rect 1797 44691 1847 44715
rect 134847 44749 134897 44773
rect 134847 44715 134855 44749
rect 134889 44715 134897 44749
rect 134847 44691 134897 44715
rect 1797 44413 1847 44437
rect 1797 44379 1805 44413
rect 1839 44379 1847 44413
rect 1797 44355 1847 44379
rect 134847 44413 134897 44437
rect 134847 44379 134855 44413
rect 134889 44379 134897 44413
rect 134847 44355 134897 44379
rect 1797 44077 1847 44101
rect 1797 44043 1805 44077
rect 1839 44043 1847 44077
rect 1797 44019 1847 44043
rect 134847 44077 134897 44101
rect 134847 44043 134855 44077
rect 134889 44043 134897 44077
rect 134847 44019 134897 44043
rect 1797 43741 1847 43765
rect 1797 43707 1805 43741
rect 1839 43707 1847 43741
rect 1797 43683 1847 43707
rect 134847 43741 134897 43765
rect 134847 43707 134855 43741
rect 134889 43707 134897 43741
rect 134847 43683 134897 43707
rect 1797 43405 1847 43429
rect 1797 43371 1805 43405
rect 1839 43371 1847 43405
rect 1797 43347 1847 43371
rect 134847 43405 134897 43429
rect 134847 43371 134855 43405
rect 134889 43371 134897 43405
rect 134847 43347 134897 43371
rect 1797 43069 1847 43093
rect 1797 43035 1805 43069
rect 1839 43035 1847 43069
rect 1797 43011 1847 43035
rect 134847 43069 134897 43093
rect 134847 43035 134855 43069
rect 134889 43035 134897 43069
rect 134847 43011 134897 43035
rect 1797 42733 1847 42757
rect 1797 42699 1805 42733
rect 1839 42699 1847 42733
rect 1797 42675 1847 42699
rect 134847 42733 134897 42757
rect 134847 42699 134855 42733
rect 134889 42699 134897 42733
rect 134847 42675 134897 42699
rect 1797 42397 1847 42421
rect 1797 42363 1805 42397
rect 1839 42363 1847 42397
rect 1797 42339 1847 42363
rect 134847 42397 134897 42421
rect 134847 42363 134855 42397
rect 134889 42363 134897 42397
rect 134847 42339 134897 42363
rect 1797 42061 1847 42085
rect 1797 42027 1805 42061
rect 1839 42027 1847 42061
rect 1797 42003 1847 42027
rect 134847 42061 134897 42085
rect 134847 42027 134855 42061
rect 134889 42027 134897 42061
rect 134847 42003 134897 42027
rect 1797 41725 1847 41749
rect 1797 41691 1805 41725
rect 1839 41691 1847 41725
rect 1797 41667 1847 41691
rect 134847 41725 134897 41749
rect 134847 41691 134855 41725
rect 134889 41691 134897 41725
rect 134847 41667 134897 41691
rect 1797 41389 1847 41413
rect 1797 41355 1805 41389
rect 1839 41355 1847 41389
rect 1797 41331 1847 41355
rect 134847 41389 134897 41413
rect 134847 41355 134855 41389
rect 134889 41355 134897 41389
rect 134847 41331 134897 41355
rect 1797 41053 1847 41077
rect 1797 41019 1805 41053
rect 1839 41019 1847 41053
rect 1797 40995 1847 41019
rect 134847 41053 134897 41077
rect 134847 41019 134855 41053
rect 134889 41019 134897 41053
rect 134847 40995 134897 41019
rect 1797 40717 1847 40741
rect 1797 40683 1805 40717
rect 1839 40683 1847 40717
rect 1797 40659 1847 40683
rect 134847 40717 134897 40741
rect 134847 40683 134855 40717
rect 134889 40683 134897 40717
rect 134847 40659 134897 40683
rect 1797 40381 1847 40405
rect 1797 40347 1805 40381
rect 1839 40347 1847 40381
rect 1797 40323 1847 40347
rect 134847 40381 134897 40405
rect 134847 40347 134855 40381
rect 134889 40347 134897 40381
rect 134847 40323 134897 40347
rect 1797 40045 1847 40069
rect 1797 40011 1805 40045
rect 1839 40011 1847 40045
rect 1797 39987 1847 40011
rect 134847 40045 134897 40069
rect 134847 40011 134855 40045
rect 134889 40011 134897 40045
rect 134847 39987 134897 40011
rect 1797 39709 1847 39733
rect 1797 39675 1805 39709
rect 1839 39675 1847 39709
rect 1797 39651 1847 39675
rect 134847 39709 134897 39733
rect 134847 39675 134855 39709
rect 134889 39675 134897 39709
rect 134847 39651 134897 39675
rect 1797 39373 1847 39397
rect 1797 39339 1805 39373
rect 1839 39339 1847 39373
rect 1797 39315 1847 39339
rect 134847 39373 134897 39397
rect 134847 39339 134855 39373
rect 134889 39339 134897 39373
rect 134847 39315 134897 39339
rect 1797 39037 1847 39061
rect 1797 39003 1805 39037
rect 1839 39003 1847 39037
rect 1797 38979 1847 39003
rect 134847 39037 134897 39061
rect 134847 39003 134855 39037
rect 134889 39003 134897 39037
rect 134847 38979 134897 39003
rect 1797 38701 1847 38725
rect 1797 38667 1805 38701
rect 1839 38667 1847 38701
rect 1797 38643 1847 38667
rect 134847 38701 134897 38725
rect 134847 38667 134855 38701
rect 134889 38667 134897 38701
rect 134847 38643 134897 38667
rect 1797 38365 1847 38389
rect 1797 38331 1805 38365
rect 1839 38331 1847 38365
rect 1797 38307 1847 38331
rect 134847 38365 134897 38389
rect 134847 38331 134855 38365
rect 134889 38331 134897 38365
rect 134847 38307 134897 38331
rect 1797 38029 1847 38053
rect 1797 37995 1805 38029
rect 1839 37995 1847 38029
rect 1797 37971 1847 37995
rect 134847 38029 134897 38053
rect 134847 37995 134855 38029
rect 134889 37995 134897 38029
rect 134847 37971 134897 37995
rect 1797 37693 1847 37717
rect 1797 37659 1805 37693
rect 1839 37659 1847 37693
rect 1797 37635 1847 37659
rect 134847 37693 134897 37717
rect 134847 37659 134855 37693
rect 134889 37659 134897 37693
rect 134847 37635 134897 37659
rect 1797 37357 1847 37381
rect 1797 37323 1805 37357
rect 1839 37323 1847 37357
rect 1797 37299 1847 37323
rect 134847 37357 134897 37381
rect 134847 37323 134855 37357
rect 134889 37323 134897 37357
rect 134847 37299 134897 37323
rect 1797 37021 1847 37045
rect 1797 36987 1805 37021
rect 1839 36987 1847 37021
rect 1797 36963 1847 36987
rect 134847 37021 134897 37045
rect 134847 36987 134855 37021
rect 134889 36987 134897 37021
rect 134847 36963 134897 36987
rect 1797 36685 1847 36709
rect 1797 36651 1805 36685
rect 1839 36651 1847 36685
rect 1797 36627 1847 36651
rect 134847 36685 134897 36709
rect 134847 36651 134855 36685
rect 134889 36651 134897 36685
rect 134847 36627 134897 36651
rect 1797 36349 1847 36373
rect 1797 36315 1805 36349
rect 1839 36315 1847 36349
rect 1797 36291 1847 36315
rect 134847 36349 134897 36373
rect 134847 36315 134855 36349
rect 134889 36315 134897 36349
rect 134847 36291 134897 36315
rect 1797 36013 1847 36037
rect 1797 35979 1805 36013
rect 1839 35979 1847 36013
rect 1797 35955 1847 35979
rect 134847 36013 134897 36037
rect 134847 35979 134855 36013
rect 134889 35979 134897 36013
rect 134847 35955 134897 35979
rect 1797 35677 1847 35701
rect 1797 35643 1805 35677
rect 1839 35643 1847 35677
rect 1797 35619 1847 35643
rect 134847 35677 134897 35701
rect 134847 35643 134855 35677
rect 134889 35643 134897 35677
rect 134847 35619 134897 35643
rect 1797 35341 1847 35365
rect 1797 35307 1805 35341
rect 1839 35307 1847 35341
rect 1797 35283 1847 35307
rect 134847 35341 134897 35365
rect 134847 35307 134855 35341
rect 134889 35307 134897 35341
rect 134847 35283 134897 35307
rect 1797 35005 1847 35029
rect 1797 34971 1805 35005
rect 1839 34971 1847 35005
rect 1797 34947 1847 34971
rect 134847 35005 134897 35029
rect 134847 34971 134855 35005
rect 134889 34971 134897 35005
rect 134847 34947 134897 34971
rect 1797 34669 1847 34693
rect 1797 34635 1805 34669
rect 1839 34635 1847 34669
rect 1797 34611 1847 34635
rect 134847 34669 134897 34693
rect 134847 34635 134855 34669
rect 134889 34635 134897 34669
rect 134847 34611 134897 34635
rect 1797 34333 1847 34357
rect 1797 34299 1805 34333
rect 1839 34299 1847 34333
rect 1797 34275 1847 34299
rect 134847 34333 134897 34357
rect 134847 34299 134855 34333
rect 134889 34299 134897 34333
rect 134847 34275 134897 34299
rect 1797 33997 1847 34021
rect 1797 33963 1805 33997
rect 1839 33963 1847 33997
rect 1797 33939 1847 33963
rect 134847 33997 134897 34021
rect 134847 33963 134855 33997
rect 134889 33963 134897 33997
rect 134847 33939 134897 33963
rect 1797 33661 1847 33685
rect 1797 33627 1805 33661
rect 1839 33627 1847 33661
rect 1797 33603 1847 33627
rect 134847 33661 134897 33685
rect 134847 33627 134855 33661
rect 134889 33627 134897 33661
rect 134847 33603 134897 33627
rect 1797 33325 1847 33349
rect 1797 33291 1805 33325
rect 1839 33291 1847 33325
rect 1797 33267 1847 33291
rect 134847 33325 134897 33349
rect 134847 33291 134855 33325
rect 134889 33291 134897 33325
rect 134847 33267 134897 33291
rect 1797 32989 1847 33013
rect 1797 32955 1805 32989
rect 1839 32955 1847 32989
rect 1797 32931 1847 32955
rect 134847 32989 134897 33013
rect 134847 32955 134855 32989
rect 134889 32955 134897 32989
rect 134847 32931 134897 32955
rect 1797 32653 1847 32677
rect 1797 32619 1805 32653
rect 1839 32619 1847 32653
rect 1797 32595 1847 32619
rect 134847 32653 134897 32677
rect 134847 32619 134855 32653
rect 134889 32619 134897 32653
rect 134847 32595 134897 32619
rect 1797 32317 1847 32341
rect 1797 32283 1805 32317
rect 1839 32283 1847 32317
rect 1797 32259 1847 32283
rect 134847 32317 134897 32341
rect 134847 32283 134855 32317
rect 134889 32283 134897 32317
rect 134847 32259 134897 32283
rect 1797 31981 1847 32005
rect 1797 31947 1805 31981
rect 1839 31947 1847 31981
rect 1797 31923 1847 31947
rect 134847 31981 134897 32005
rect 134847 31947 134855 31981
rect 134889 31947 134897 31981
rect 134847 31923 134897 31947
rect 1797 31645 1847 31669
rect 1797 31611 1805 31645
rect 1839 31611 1847 31645
rect 1797 31587 1847 31611
rect 134847 31645 134897 31669
rect 134847 31611 134855 31645
rect 134889 31611 134897 31645
rect 134847 31587 134897 31611
rect 1797 31309 1847 31333
rect 1797 31275 1805 31309
rect 1839 31275 1847 31309
rect 1797 31251 1847 31275
rect 134847 31309 134897 31333
rect 134847 31275 134855 31309
rect 134889 31275 134897 31309
rect 134847 31251 134897 31275
rect 1797 30973 1847 30997
rect 1797 30939 1805 30973
rect 1839 30939 1847 30973
rect 1797 30915 1847 30939
rect 134847 30973 134897 30997
rect 134847 30939 134855 30973
rect 134889 30939 134897 30973
rect 134847 30915 134897 30939
rect 1797 30637 1847 30661
rect 1797 30603 1805 30637
rect 1839 30603 1847 30637
rect 1797 30579 1847 30603
rect 134847 30637 134897 30661
rect 134847 30603 134855 30637
rect 134889 30603 134897 30637
rect 134847 30579 134897 30603
rect 1797 30301 1847 30325
rect 1797 30267 1805 30301
rect 1839 30267 1847 30301
rect 1797 30243 1847 30267
rect 134847 30301 134897 30325
rect 134847 30267 134855 30301
rect 134889 30267 134897 30301
rect 134847 30243 134897 30267
rect 1797 29965 1847 29989
rect 1797 29931 1805 29965
rect 1839 29931 1847 29965
rect 1797 29907 1847 29931
rect 134847 29965 134897 29989
rect 134847 29931 134855 29965
rect 134889 29931 134897 29965
rect 134847 29907 134897 29931
rect 1797 29629 1847 29653
rect 1797 29595 1805 29629
rect 1839 29595 1847 29629
rect 1797 29571 1847 29595
rect 134847 29629 134897 29653
rect 134847 29595 134855 29629
rect 134889 29595 134897 29629
rect 134847 29571 134897 29595
rect 1797 29293 1847 29317
rect 1797 29259 1805 29293
rect 1839 29259 1847 29293
rect 1797 29235 1847 29259
rect 134847 29293 134897 29317
rect 134847 29259 134855 29293
rect 134889 29259 134897 29293
rect 134847 29235 134897 29259
rect 1797 28957 1847 28981
rect 1797 28923 1805 28957
rect 1839 28923 1847 28957
rect 1797 28899 1847 28923
rect 134847 28957 134897 28981
rect 134847 28923 134855 28957
rect 134889 28923 134897 28957
rect 134847 28899 134897 28923
rect 1797 28621 1847 28645
rect 1797 28587 1805 28621
rect 1839 28587 1847 28621
rect 1797 28563 1847 28587
rect 134847 28621 134897 28645
rect 134847 28587 134855 28621
rect 134889 28587 134897 28621
rect 134847 28563 134897 28587
rect 1797 28285 1847 28309
rect 1797 28251 1805 28285
rect 1839 28251 1847 28285
rect 1797 28227 1847 28251
rect 134847 28285 134897 28309
rect 134847 28251 134855 28285
rect 134889 28251 134897 28285
rect 134847 28227 134897 28251
rect 1797 27949 1847 27973
rect 1797 27915 1805 27949
rect 1839 27915 1847 27949
rect 1797 27891 1847 27915
rect 134847 27949 134897 27973
rect 134847 27915 134855 27949
rect 134889 27915 134897 27949
rect 134847 27891 134897 27915
rect 1797 27613 1847 27637
rect 1797 27579 1805 27613
rect 1839 27579 1847 27613
rect 1797 27555 1847 27579
rect 134847 27613 134897 27637
rect 134847 27579 134855 27613
rect 134889 27579 134897 27613
rect 134847 27555 134897 27579
rect 1797 27277 1847 27301
rect 1797 27243 1805 27277
rect 1839 27243 1847 27277
rect 1797 27219 1847 27243
rect 134847 27277 134897 27301
rect 134847 27243 134855 27277
rect 134889 27243 134897 27277
rect 134847 27219 134897 27243
rect 1797 26941 1847 26965
rect 1797 26907 1805 26941
rect 1839 26907 1847 26941
rect 1797 26883 1847 26907
rect 134847 26941 134897 26965
rect 134847 26907 134855 26941
rect 134889 26907 134897 26941
rect 134847 26883 134897 26907
rect 1797 26605 1847 26629
rect 1797 26571 1805 26605
rect 1839 26571 1847 26605
rect 1797 26547 1847 26571
rect 134847 26605 134897 26629
rect 134847 26571 134855 26605
rect 134889 26571 134897 26605
rect 134847 26547 134897 26571
rect 1797 26269 1847 26293
rect 1797 26235 1805 26269
rect 1839 26235 1847 26269
rect 1797 26211 1847 26235
rect 134847 26269 134897 26293
rect 134847 26235 134855 26269
rect 134889 26235 134897 26269
rect 134847 26211 134897 26235
rect 1797 25933 1847 25957
rect 1797 25899 1805 25933
rect 1839 25899 1847 25933
rect 1797 25875 1847 25899
rect 134847 25933 134897 25957
rect 134847 25899 134855 25933
rect 134889 25899 134897 25933
rect 134847 25875 134897 25899
rect 1797 25597 1847 25621
rect 1797 25563 1805 25597
rect 1839 25563 1847 25597
rect 1797 25539 1847 25563
rect 134847 25597 134897 25621
rect 134847 25563 134855 25597
rect 134889 25563 134897 25597
rect 134847 25539 134897 25563
rect 1797 25261 1847 25285
rect 1797 25227 1805 25261
rect 1839 25227 1847 25261
rect 1797 25203 1847 25227
rect 134847 25261 134897 25285
rect 134847 25227 134855 25261
rect 134889 25227 134897 25261
rect 134847 25203 134897 25227
rect 1797 24925 1847 24949
rect 1797 24891 1805 24925
rect 1839 24891 1847 24925
rect 1797 24867 1847 24891
rect 134847 24925 134897 24949
rect 134847 24891 134855 24925
rect 134889 24891 134897 24925
rect 134847 24867 134897 24891
rect 1797 24589 1847 24613
rect 1797 24555 1805 24589
rect 1839 24555 1847 24589
rect 1797 24531 1847 24555
rect 134847 24589 134897 24613
rect 134847 24555 134855 24589
rect 134889 24555 134897 24589
rect 134847 24531 134897 24555
rect 1797 24253 1847 24277
rect 1797 24219 1805 24253
rect 1839 24219 1847 24253
rect 1797 24195 1847 24219
rect 134847 24253 134897 24277
rect 134847 24219 134855 24253
rect 134889 24219 134897 24253
rect 134847 24195 134897 24219
rect 1797 23917 1847 23941
rect 1797 23883 1805 23917
rect 1839 23883 1847 23917
rect 1797 23859 1847 23883
rect 134847 23917 134897 23941
rect 134847 23883 134855 23917
rect 134889 23883 134897 23917
rect 134847 23859 134897 23883
rect 1797 23581 1847 23605
rect 1797 23547 1805 23581
rect 1839 23547 1847 23581
rect 1797 23523 1847 23547
rect 134847 23581 134897 23605
rect 134847 23547 134855 23581
rect 134889 23547 134897 23581
rect 134847 23523 134897 23547
rect 1797 23245 1847 23269
rect 1797 23211 1805 23245
rect 1839 23211 1847 23245
rect 1797 23187 1847 23211
rect 134847 23245 134897 23269
rect 134847 23211 134855 23245
rect 134889 23211 134897 23245
rect 134847 23187 134897 23211
rect 1797 22909 1847 22933
rect 1797 22875 1805 22909
rect 1839 22875 1847 22909
rect 1797 22851 1847 22875
rect 134847 22909 134897 22933
rect 134847 22875 134855 22909
rect 134889 22875 134897 22909
rect 134847 22851 134897 22875
rect 1797 22573 1847 22597
rect 1797 22539 1805 22573
rect 1839 22539 1847 22573
rect 1797 22515 1847 22539
rect 134847 22573 134897 22597
rect 134847 22539 134855 22573
rect 134889 22539 134897 22573
rect 134847 22515 134897 22539
rect 1797 22237 1847 22261
rect 1797 22203 1805 22237
rect 1839 22203 1847 22237
rect 1797 22179 1847 22203
rect 134847 22237 134897 22261
rect 134847 22203 134855 22237
rect 134889 22203 134897 22237
rect 134847 22179 134897 22203
rect 1797 21901 1847 21925
rect 1797 21867 1805 21901
rect 1839 21867 1847 21901
rect 1797 21843 1847 21867
rect 134847 21901 134897 21925
rect 134847 21867 134855 21901
rect 134889 21867 134897 21901
rect 134847 21843 134897 21867
rect 1797 21565 1847 21589
rect 1797 21531 1805 21565
rect 1839 21531 1847 21565
rect 1797 21507 1847 21531
rect 134847 21565 134897 21589
rect 134847 21531 134855 21565
rect 134889 21531 134897 21565
rect 134847 21507 134897 21531
rect 1797 21229 1847 21253
rect 1797 21195 1805 21229
rect 1839 21195 1847 21229
rect 1797 21171 1847 21195
rect 134847 21229 134897 21253
rect 134847 21195 134855 21229
rect 134889 21195 134897 21229
rect 134847 21171 134897 21195
rect 1797 20893 1847 20917
rect 1797 20859 1805 20893
rect 1839 20859 1847 20893
rect 1797 20835 1847 20859
rect 134847 20893 134897 20917
rect 134847 20859 134855 20893
rect 134889 20859 134897 20893
rect 134847 20835 134897 20859
rect 1797 20557 1847 20581
rect 1797 20523 1805 20557
rect 1839 20523 1847 20557
rect 1797 20499 1847 20523
rect 134847 20557 134897 20581
rect 134847 20523 134855 20557
rect 134889 20523 134897 20557
rect 134847 20499 134897 20523
rect 1797 20221 1847 20245
rect 1797 20187 1805 20221
rect 1839 20187 1847 20221
rect 1797 20163 1847 20187
rect 134847 20221 134897 20245
rect 134847 20187 134855 20221
rect 134889 20187 134897 20221
rect 134847 20163 134897 20187
rect 1797 19885 1847 19909
rect 1797 19851 1805 19885
rect 1839 19851 1847 19885
rect 1797 19827 1847 19851
rect 134847 19885 134897 19909
rect 134847 19851 134855 19885
rect 134889 19851 134897 19885
rect 134847 19827 134897 19851
rect 1797 19549 1847 19573
rect 1797 19515 1805 19549
rect 1839 19515 1847 19549
rect 1797 19491 1847 19515
rect 134847 19549 134897 19573
rect 134847 19515 134855 19549
rect 134889 19515 134897 19549
rect 134847 19491 134897 19515
rect 1797 19213 1847 19237
rect 1797 19179 1805 19213
rect 1839 19179 1847 19213
rect 1797 19155 1847 19179
rect 134847 19213 134897 19237
rect 134847 19179 134855 19213
rect 134889 19179 134897 19213
rect 134847 19155 134897 19179
rect 1797 18877 1847 18901
rect 1797 18843 1805 18877
rect 1839 18843 1847 18877
rect 1797 18819 1847 18843
rect 134847 18877 134897 18901
rect 134847 18843 134855 18877
rect 134889 18843 134897 18877
rect 134847 18819 134897 18843
rect 1797 18541 1847 18565
rect 1797 18507 1805 18541
rect 1839 18507 1847 18541
rect 1797 18483 1847 18507
rect 134847 18541 134897 18565
rect 134847 18507 134855 18541
rect 134889 18507 134897 18541
rect 134847 18483 134897 18507
rect 1797 18205 1847 18229
rect 1797 18171 1805 18205
rect 1839 18171 1847 18205
rect 1797 18147 1847 18171
rect 134847 18205 134897 18229
rect 134847 18171 134855 18205
rect 134889 18171 134897 18205
rect 134847 18147 134897 18171
rect 1797 17869 1847 17893
rect 1797 17835 1805 17869
rect 1839 17835 1847 17869
rect 1797 17811 1847 17835
rect 134847 17869 134897 17893
rect 134847 17835 134855 17869
rect 134889 17835 134897 17869
rect 134847 17811 134897 17835
rect 1797 17533 1847 17557
rect 1797 17499 1805 17533
rect 1839 17499 1847 17533
rect 1797 17475 1847 17499
rect 134847 17533 134897 17557
rect 134847 17499 134855 17533
rect 134889 17499 134897 17533
rect 134847 17475 134897 17499
rect 1797 17197 1847 17221
rect 1797 17163 1805 17197
rect 1839 17163 1847 17197
rect 1797 17139 1847 17163
rect 134847 17197 134897 17221
rect 134847 17163 134855 17197
rect 134889 17163 134897 17197
rect 134847 17139 134897 17163
rect 1797 16861 1847 16885
rect 1797 16827 1805 16861
rect 1839 16827 1847 16861
rect 1797 16803 1847 16827
rect 134847 16861 134897 16885
rect 134847 16827 134855 16861
rect 134889 16827 134897 16861
rect 134847 16803 134897 16827
rect 1797 16525 1847 16549
rect 1797 16491 1805 16525
rect 1839 16491 1847 16525
rect 1797 16467 1847 16491
rect 134847 16525 134897 16549
rect 134847 16491 134855 16525
rect 134889 16491 134897 16525
rect 134847 16467 134897 16491
rect 1797 16189 1847 16213
rect 1797 16155 1805 16189
rect 1839 16155 1847 16189
rect 1797 16131 1847 16155
rect 134847 16189 134897 16213
rect 134847 16155 134855 16189
rect 134889 16155 134897 16189
rect 134847 16131 134897 16155
rect 1797 15853 1847 15877
rect 1797 15819 1805 15853
rect 1839 15819 1847 15853
rect 1797 15795 1847 15819
rect 134847 15853 134897 15877
rect 134847 15819 134855 15853
rect 134889 15819 134897 15853
rect 134847 15795 134897 15819
rect 1797 15517 1847 15541
rect 1797 15483 1805 15517
rect 1839 15483 1847 15517
rect 1797 15459 1847 15483
rect 134847 15517 134897 15541
rect 134847 15483 134855 15517
rect 134889 15483 134897 15517
rect 134847 15459 134897 15483
rect 1797 15181 1847 15205
rect 1797 15147 1805 15181
rect 1839 15147 1847 15181
rect 1797 15123 1847 15147
rect 134847 15181 134897 15205
rect 134847 15147 134855 15181
rect 134889 15147 134897 15181
rect 134847 15123 134897 15147
rect 1797 14845 1847 14869
rect 1797 14811 1805 14845
rect 1839 14811 1847 14845
rect 1797 14787 1847 14811
rect 134847 14845 134897 14869
rect 134847 14811 134855 14845
rect 134889 14811 134897 14845
rect 134847 14787 134897 14811
rect 1797 14509 1847 14533
rect 1797 14475 1805 14509
rect 1839 14475 1847 14509
rect 1797 14451 1847 14475
rect 134847 14509 134897 14533
rect 134847 14475 134855 14509
rect 134889 14475 134897 14509
rect 134847 14451 134897 14475
rect 1797 14173 1847 14197
rect 1797 14139 1805 14173
rect 1839 14139 1847 14173
rect 1797 14115 1847 14139
rect 134847 14173 134897 14197
rect 134847 14139 134855 14173
rect 134889 14139 134897 14173
rect 134847 14115 134897 14139
rect 1797 13837 1847 13861
rect 1797 13803 1805 13837
rect 1839 13803 1847 13837
rect 1797 13779 1847 13803
rect 134847 13837 134897 13861
rect 134847 13803 134855 13837
rect 134889 13803 134897 13837
rect 134847 13779 134897 13803
rect 1797 13501 1847 13525
rect 1797 13467 1805 13501
rect 1839 13467 1847 13501
rect 1797 13443 1847 13467
rect 134847 13501 134897 13525
rect 134847 13467 134855 13501
rect 134889 13467 134897 13501
rect 134847 13443 134897 13467
rect 1797 13165 1847 13189
rect 1797 13131 1805 13165
rect 1839 13131 1847 13165
rect 1797 13107 1847 13131
rect 134847 13165 134897 13189
rect 134847 13131 134855 13165
rect 134889 13131 134897 13165
rect 134847 13107 134897 13131
rect 1797 12829 1847 12853
rect 1797 12795 1805 12829
rect 1839 12795 1847 12829
rect 1797 12771 1847 12795
rect 134847 12829 134897 12853
rect 134847 12795 134855 12829
rect 134889 12795 134897 12829
rect 134847 12771 134897 12795
rect 1797 12493 1847 12517
rect 1797 12459 1805 12493
rect 1839 12459 1847 12493
rect 1797 12435 1847 12459
rect 134847 12493 134897 12517
rect 134847 12459 134855 12493
rect 134889 12459 134897 12493
rect 134847 12435 134897 12459
rect 1797 12157 1847 12181
rect 1797 12123 1805 12157
rect 1839 12123 1847 12157
rect 1797 12099 1847 12123
rect 134847 12157 134897 12181
rect 134847 12123 134855 12157
rect 134889 12123 134897 12157
rect 134847 12099 134897 12123
rect 1797 11821 1847 11845
rect 1797 11787 1805 11821
rect 1839 11787 1847 11821
rect 1797 11763 1847 11787
rect 134847 11821 134897 11845
rect 134847 11787 134855 11821
rect 134889 11787 134897 11821
rect 134847 11763 134897 11787
rect 1797 11485 1847 11509
rect 1797 11451 1805 11485
rect 1839 11451 1847 11485
rect 1797 11427 1847 11451
rect 134847 11485 134897 11509
rect 134847 11451 134855 11485
rect 134889 11451 134897 11485
rect 134847 11427 134897 11451
rect 1797 11149 1847 11173
rect 1797 11115 1805 11149
rect 1839 11115 1847 11149
rect 1797 11091 1847 11115
rect 134847 11149 134897 11173
rect 134847 11115 134855 11149
rect 134889 11115 134897 11149
rect 134847 11091 134897 11115
rect 1797 10813 1847 10837
rect 1797 10779 1805 10813
rect 1839 10779 1847 10813
rect 1797 10755 1847 10779
rect 134847 10813 134897 10837
rect 134847 10779 134855 10813
rect 134889 10779 134897 10813
rect 134847 10755 134897 10779
rect 1797 10477 1847 10501
rect 1797 10443 1805 10477
rect 1839 10443 1847 10477
rect 1797 10419 1847 10443
rect 134847 10477 134897 10501
rect 134847 10443 134855 10477
rect 134889 10443 134897 10477
rect 134847 10419 134897 10443
rect 1797 10141 1847 10165
rect 1797 10107 1805 10141
rect 1839 10107 1847 10141
rect 1797 10083 1847 10107
rect 134847 10141 134897 10165
rect 134847 10107 134855 10141
rect 134889 10107 134897 10141
rect 134847 10083 134897 10107
rect 1797 9805 1847 9829
rect 1797 9771 1805 9805
rect 1839 9771 1847 9805
rect 1797 9747 1847 9771
rect 134847 9805 134897 9829
rect 134847 9771 134855 9805
rect 134889 9771 134897 9805
rect 134847 9747 134897 9771
rect 1797 9469 1847 9493
rect 1797 9435 1805 9469
rect 1839 9435 1847 9469
rect 1797 9411 1847 9435
rect 134847 9469 134897 9493
rect 134847 9435 134855 9469
rect 134889 9435 134897 9469
rect 134847 9411 134897 9435
rect 1797 9133 1847 9157
rect 1797 9099 1805 9133
rect 1839 9099 1847 9133
rect 1797 9075 1847 9099
rect 134847 9133 134897 9157
rect 134847 9099 134855 9133
rect 134889 9099 134897 9133
rect 134847 9075 134897 9099
rect 1797 8797 1847 8821
rect 1797 8763 1805 8797
rect 1839 8763 1847 8797
rect 1797 8739 1847 8763
rect 134847 8797 134897 8821
rect 134847 8763 134855 8797
rect 134889 8763 134897 8797
rect 134847 8739 134897 8763
rect 1797 8461 1847 8485
rect 1797 8427 1805 8461
rect 1839 8427 1847 8461
rect 1797 8403 1847 8427
rect 134847 8461 134897 8485
rect 134847 8427 134855 8461
rect 134889 8427 134897 8461
rect 134847 8403 134897 8427
rect 1797 8125 1847 8149
rect 1797 8091 1805 8125
rect 1839 8091 1847 8125
rect 1797 8067 1847 8091
rect 134847 8125 134897 8149
rect 134847 8091 134855 8125
rect 134889 8091 134897 8125
rect 134847 8067 134897 8091
rect 1797 7789 1847 7813
rect 1797 7755 1805 7789
rect 1839 7755 1847 7789
rect 1797 7731 1847 7755
rect 134847 7789 134897 7813
rect 134847 7755 134855 7789
rect 134889 7755 134897 7789
rect 134847 7731 134897 7755
rect 1797 7453 1847 7477
rect 1797 7419 1805 7453
rect 1839 7419 1847 7453
rect 1797 7395 1847 7419
rect 134847 7453 134897 7477
rect 134847 7419 134855 7453
rect 134889 7419 134897 7453
rect 134847 7395 134897 7419
rect 1797 7117 1847 7141
rect 1797 7083 1805 7117
rect 1839 7083 1847 7117
rect 1797 7059 1847 7083
rect 134847 7117 134897 7141
rect 134847 7083 134855 7117
rect 134889 7083 134897 7117
rect 134847 7059 134897 7083
rect 1797 6781 1847 6805
rect 1797 6747 1805 6781
rect 1839 6747 1847 6781
rect 1797 6723 1847 6747
rect 134847 6781 134897 6805
rect 134847 6747 134855 6781
rect 134889 6747 134897 6781
rect 134847 6723 134897 6747
rect 1797 6445 1847 6469
rect 1797 6411 1805 6445
rect 1839 6411 1847 6445
rect 1797 6387 1847 6411
rect 134847 6445 134897 6469
rect 134847 6411 134855 6445
rect 134889 6411 134897 6445
rect 134847 6387 134897 6411
rect 1797 6109 1847 6133
rect 1797 6075 1805 6109
rect 1839 6075 1847 6109
rect 1797 6051 1847 6075
rect 134847 6109 134897 6133
rect 134847 6075 134855 6109
rect 134889 6075 134897 6109
rect 134847 6051 134897 6075
rect 1797 5773 1847 5797
rect 1797 5739 1805 5773
rect 1839 5739 1847 5773
rect 1797 5715 1847 5739
rect 134847 5773 134897 5797
rect 134847 5739 134855 5773
rect 134889 5739 134897 5773
rect 134847 5715 134897 5739
rect 1797 5437 1847 5461
rect 1797 5403 1805 5437
rect 1839 5403 1847 5437
rect 1797 5379 1847 5403
rect 134847 5437 134897 5461
rect 134847 5403 134855 5437
rect 134889 5403 134897 5437
rect 134847 5379 134897 5403
rect 1797 5101 1847 5125
rect 1797 5067 1805 5101
rect 1839 5067 1847 5101
rect 1797 5043 1847 5067
rect 134847 5101 134897 5125
rect 134847 5067 134855 5101
rect 134889 5067 134897 5101
rect 134847 5043 134897 5067
rect 1797 4765 1847 4789
rect 1797 4731 1805 4765
rect 1839 4731 1847 4765
rect 1797 4707 1847 4731
rect 134847 4765 134897 4789
rect 134847 4731 134855 4765
rect 134889 4731 134897 4765
rect 134847 4707 134897 4731
rect 1797 4429 1847 4453
rect 1797 4395 1805 4429
rect 1839 4395 1847 4429
rect 1797 4371 1847 4395
rect 134847 4429 134897 4453
rect 134847 4395 134855 4429
rect 134889 4395 134897 4429
rect 134847 4371 134897 4395
rect 1797 4093 1847 4117
rect 1797 4059 1805 4093
rect 1839 4059 1847 4093
rect 1797 4035 1847 4059
rect 134847 4093 134897 4117
rect 134847 4059 134855 4093
rect 134889 4059 134897 4093
rect 134847 4035 134897 4059
rect 1797 3757 1847 3781
rect 1797 3723 1805 3757
rect 1839 3723 1847 3757
rect 1797 3699 1847 3723
rect 134847 3757 134897 3781
rect 134847 3723 134855 3757
rect 134889 3723 134897 3757
rect 134847 3699 134897 3723
rect 1797 3421 1847 3445
rect 1797 3387 1805 3421
rect 1839 3387 1847 3421
rect 1797 3363 1847 3387
rect 134847 3421 134897 3445
rect 134847 3387 134855 3421
rect 134889 3387 134897 3421
rect 134847 3363 134897 3387
rect 1797 3085 1847 3109
rect 1797 3051 1805 3085
rect 1839 3051 1847 3085
rect 1797 3027 1847 3051
rect 134847 3085 134897 3109
rect 134847 3051 134855 3085
rect 134889 3051 134897 3085
rect 134847 3027 134897 3051
rect 1797 2749 1847 2773
rect 1797 2715 1805 2749
rect 1839 2715 1847 2749
rect 1797 2691 1847 2715
rect 134847 2749 134897 2773
rect 134847 2715 134855 2749
rect 134889 2715 134897 2749
rect 134847 2691 134897 2715
rect 1797 2413 1847 2437
rect 1797 2379 1805 2413
rect 1839 2379 1847 2413
rect 1797 2355 1847 2379
rect 134847 2413 134897 2437
rect 134847 2379 134855 2413
rect 134889 2379 134897 2413
rect 134847 2355 134897 2379
rect 1797 2077 1847 2101
rect 1797 2043 1805 2077
rect 1839 2043 1847 2077
rect 1797 2019 1847 2043
rect 134847 2077 134897 2101
rect 134847 2043 134855 2077
rect 134889 2043 134897 2077
rect 134847 2019 134897 2043
rect 2133 1741 2183 1765
rect 2133 1707 2141 1741
rect 2175 1707 2183 1741
rect 2133 1683 2183 1707
rect 2469 1741 2519 1765
rect 2469 1707 2477 1741
rect 2511 1707 2519 1741
rect 2469 1683 2519 1707
rect 2805 1741 2855 1765
rect 2805 1707 2813 1741
rect 2847 1707 2855 1741
rect 2805 1683 2855 1707
rect 3141 1741 3191 1765
rect 3141 1707 3149 1741
rect 3183 1707 3191 1741
rect 3141 1683 3191 1707
rect 3477 1741 3527 1765
rect 3477 1707 3485 1741
rect 3519 1707 3527 1741
rect 3477 1683 3527 1707
rect 3813 1741 3863 1765
rect 3813 1707 3821 1741
rect 3855 1707 3863 1741
rect 3813 1683 3863 1707
rect 4149 1741 4199 1765
rect 4149 1707 4157 1741
rect 4191 1707 4199 1741
rect 4149 1683 4199 1707
rect 4485 1741 4535 1765
rect 4485 1707 4493 1741
rect 4527 1707 4535 1741
rect 4485 1683 4535 1707
rect 4821 1741 4871 1765
rect 4821 1707 4829 1741
rect 4863 1707 4871 1741
rect 4821 1683 4871 1707
rect 5157 1741 5207 1765
rect 5157 1707 5165 1741
rect 5199 1707 5207 1741
rect 5157 1683 5207 1707
rect 5493 1741 5543 1765
rect 5493 1707 5501 1741
rect 5535 1707 5543 1741
rect 5493 1683 5543 1707
rect 5829 1741 5879 1765
rect 5829 1707 5837 1741
rect 5871 1707 5879 1741
rect 5829 1683 5879 1707
rect 6165 1741 6215 1765
rect 6165 1707 6173 1741
rect 6207 1707 6215 1741
rect 6165 1683 6215 1707
rect 6501 1741 6551 1765
rect 6501 1707 6509 1741
rect 6543 1707 6551 1741
rect 6501 1683 6551 1707
rect 6837 1741 6887 1765
rect 6837 1707 6845 1741
rect 6879 1707 6887 1741
rect 6837 1683 6887 1707
rect 7173 1741 7223 1765
rect 7173 1707 7181 1741
rect 7215 1707 7223 1741
rect 7173 1683 7223 1707
rect 7509 1741 7559 1765
rect 7509 1707 7517 1741
rect 7551 1707 7559 1741
rect 7509 1683 7559 1707
rect 7845 1741 7895 1765
rect 7845 1707 7853 1741
rect 7887 1707 7895 1741
rect 7845 1683 7895 1707
rect 8181 1741 8231 1765
rect 8181 1707 8189 1741
rect 8223 1707 8231 1741
rect 8181 1683 8231 1707
rect 8517 1741 8567 1765
rect 8517 1707 8525 1741
rect 8559 1707 8567 1741
rect 8517 1683 8567 1707
rect 8853 1741 8903 1765
rect 8853 1707 8861 1741
rect 8895 1707 8903 1741
rect 8853 1683 8903 1707
rect 9189 1741 9239 1765
rect 9189 1707 9197 1741
rect 9231 1707 9239 1741
rect 9189 1683 9239 1707
rect 9525 1741 9575 1765
rect 9525 1707 9533 1741
rect 9567 1707 9575 1741
rect 9525 1683 9575 1707
rect 9861 1741 9911 1765
rect 9861 1707 9869 1741
rect 9903 1707 9911 1741
rect 9861 1683 9911 1707
rect 10197 1741 10247 1765
rect 10197 1707 10205 1741
rect 10239 1707 10247 1741
rect 10197 1683 10247 1707
rect 10533 1741 10583 1765
rect 10533 1707 10541 1741
rect 10575 1707 10583 1741
rect 10533 1683 10583 1707
rect 10869 1741 10919 1765
rect 10869 1707 10877 1741
rect 10911 1707 10919 1741
rect 10869 1683 10919 1707
rect 11205 1741 11255 1765
rect 11205 1707 11213 1741
rect 11247 1707 11255 1741
rect 11205 1683 11255 1707
rect 11541 1741 11591 1765
rect 11541 1707 11549 1741
rect 11583 1707 11591 1741
rect 11541 1683 11591 1707
rect 11877 1741 11927 1765
rect 11877 1707 11885 1741
rect 11919 1707 11927 1741
rect 11877 1683 11927 1707
rect 12213 1741 12263 1765
rect 12213 1707 12221 1741
rect 12255 1707 12263 1741
rect 12213 1683 12263 1707
rect 12549 1741 12599 1765
rect 12549 1707 12557 1741
rect 12591 1707 12599 1741
rect 12549 1683 12599 1707
rect 12885 1741 12935 1765
rect 12885 1707 12893 1741
rect 12927 1707 12935 1741
rect 12885 1683 12935 1707
rect 13221 1741 13271 1765
rect 13221 1707 13229 1741
rect 13263 1707 13271 1741
rect 13221 1683 13271 1707
rect 13557 1741 13607 1765
rect 13557 1707 13565 1741
rect 13599 1707 13607 1741
rect 13557 1683 13607 1707
rect 13893 1741 13943 1765
rect 13893 1707 13901 1741
rect 13935 1707 13943 1741
rect 13893 1683 13943 1707
rect 14229 1741 14279 1765
rect 14229 1707 14237 1741
rect 14271 1707 14279 1741
rect 14229 1683 14279 1707
rect 14565 1741 14615 1765
rect 14565 1707 14573 1741
rect 14607 1707 14615 1741
rect 14565 1683 14615 1707
rect 14901 1741 14951 1765
rect 14901 1707 14909 1741
rect 14943 1707 14951 1741
rect 14901 1683 14951 1707
rect 15237 1741 15287 1765
rect 15237 1707 15245 1741
rect 15279 1707 15287 1741
rect 15237 1683 15287 1707
rect 15573 1741 15623 1765
rect 15573 1707 15581 1741
rect 15615 1707 15623 1741
rect 15573 1683 15623 1707
rect 15909 1741 15959 1765
rect 15909 1707 15917 1741
rect 15951 1707 15959 1741
rect 15909 1683 15959 1707
rect 16245 1741 16295 1765
rect 16245 1707 16253 1741
rect 16287 1707 16295 1741
rect 16245 1683 16295 1707
rect 16581 1741 16631 1765
rect 16581 1707 16589 1741
rect 16623 1707 16631 1741
rect 16581 1683 16631 1707
rect 16917 1741 16967 1765
rect 16917 1707 16925 1741
rect 16959 1707 16967 1741
rect 16917 1683 16967 1707
rect 17253 1741 17303 1765
rect 17253 1707 17261 1741
rect 17295 1707 17303 1741
rect 17253 1683 17303 1707
rect 17589 1741 17639 1765
rect 17589 1707 17597 1741
rect 17631 1707 17639 1741
rect 17589 1683 17639 1707
rect 17925 1741 17975 1765
rect 17925 1707 17933 1741
rect 17967 1707 17975 1741
rect 17925 1683 17975 1707
rect 18261 1741 18311 1765
rect 18261 1707 18269 1741
rect 18303 1707 18311 1741
rect 18261 1683 18311 1707
rect 18597 1741 18647 1765
rect 18597 1707 18605 1741
rect 18639 1707 18647 1741
rect 18597 1683 18647 1707
rect 18933 1741 18983 1765
rect 18933 1707 18941 1741
rect 18975 1707 18983 1741
rect 18933 1683 18983 1707
rect 19269 1741 19319 1765
rect 19269 1707 19277 1741
rect 19311 1707 19319 1741
rect 19269 1683 19319 1707
rect 19605 1741 19655 1765
rect 19605 1707 19613 1741
rect 19647 1707 19655 1741
rect 19605 1683 19655 1707
rect 19941 1741 19991 1765
rect 19941 1707 19949 1741
rect 19983 1707 19991 1741
rect 19941 1683 19991 1707
rect 20277 1741 20327 1765
rect 20277 1707 20285 1741
rect 20319 1707 20327 1741
rect 20277 1683 20327 1707
rect 20613 1741 20663 1765
rect 20613 1707 20621 1741
rect 20655 1707 20663 1741
rect 20613 1683 20663 1707
rect 20949 1741 20999 1765
rect 20949 1707 20957 1741
rect 20991 1707 20999 1741
rect 20949 1683 20999 1707
rect 21285 1741 21335 1765
rect 21285 1707 21293 1741
rect 21327 1707 21335 1741
rect 21285 1683 21335 1707
rect 21621 1741 21671 1765
rect 21621 1707 21629 1741
rect 21663 1707 21671 1741
rect 21621 1683 21671 1707
rect 21957 1741 22007 1765
rect 21957 1707 21965 1741
rect 21999 1707 22007 1741
rect 21957 1683 22007 1707
rect 22293 1741 22343 1765
rect 22293 1707 22301 1741
rect 22335 1707 22343 1741
rect 22293 1683 22343 1707
rect 22629 1741 22679 1765
rect 22629 1707 22637 1741
rect 22671 1707 22679 1741
rect 22629 1683 22679 1707
rect 22965 1741 23015 1765
rect 22965 1707 22973 1741
rect 23007 1707 23015 1741
rect 22965 1683 23015 1707
rect 23301 1741 23351 1765
rect 23301 1707 23309 1741
rect 23343 1707 23351 1741
rect 23301 1683 23351 1707
rect 23637 1741 23687 1765
rect 23637 1707 23645 1741
rect 23679 1707 23687 1741
rect 23637 1683 23687 1707
rect 23973 1741 24023 1765
rect 23973 1707 23981 1741
rect 24015 1707 24023 1741
rect 23973 1683 24023 1707
rect 24309 1741 24359 1765
rect 24309 1707 24317 1741
rect 24351 1707 24359 1741
rect 24309 1683 24359 1707
rect 24645 1741 24695 1765
rect 24645 1707 24653 1741
rect 24687 1707 24695 1741
rect 24645 1683 24695 1707
rect 24981 1741 25031 1765
rect 24981 1707 24989 1741
rect 25023 1707 25031 1741
rect 24981 1683 25031 1707
rect 25317 1741 25367 1765
rect 25317 1707 25325 1741
rect 25359 1707 25367 1741
rect 25317 1683 25367 1707
rect 25653 1741 25703 1765
rect 25653 1707 25661 1741
rect 25695 1707 25703 1741
rect 25653 1683 25703 1707
rect 25989 1741 26039 1765
rect 25989 1707 25997 1741
rect 26031 1707 26039 1741
rect 25989 1683 26039 1707
rect 26325 1741 26375 1765
rect 26325 1707 26333 1741
rect 26367 1707 26375 1741
rect 26325 1683 26375 1707
rect 26661 1741 26711 1765
rect 26661 1707 26669 1741
rect 26703 1707 26711 1741
rect 26661 1683 26711 1707
rect 26997 1741 27047 1765
rect 26997 1707 27005 1741
rect 27039 1707 27047 1741
rect 26997 1683 27047 1707
rect 27333 1741 27383 1765
rect 27333 1707 27341 1741
rect 27375 1707 27383 1741
rect 27333 1683 27383 1707
rect 27669 1741 27719 1765
rect 27669 1707 27677 1741
rect 27711 1707 27719 1741
rect 27669 1683 27719 1707
rect 28005 1741 28055 1765
rect 28005 1707 28013 1741
rect 28047 1707 28055 1741
rect 28005 1683 28055 1707
rect 28341 1741 28391 1765
rect 28341 1707 28349 1741
rect 28383 1707 28391 1741
rect 28341 1683 28391 1707
rect 28677 1741 28727 1765
rect 28677 1707 28685 1741
rect 28719 1707 28727 1741
rect 28677 1683 28727 1707
rect 29013 1741 29063 1765
rect 29013 1707 29021 1741
rect 29055 1707 29063 1741
rect 29013 1683 29063 1707
rect 29349 1741 29399 1765
rect 29349 1707 29357 1741
rect 29391 1707 29399 1741
rect 29349 1683 29399 1707
rect 29685 1741 29735 1765
rect 29685 1707 29693 1741
rect 29727 1707 29735 1741
rect 29685 1683 29735 1707
rect 30021 1741 30071 1765
rect 30021 1707 30029 1741
rect 30063 1707 30071 1741
rect 30021 1683 30071 1707
rect 30357 1741 30407 1765
rect 30357 1707 30365 1741
rect 30399 1707 30407 1741
rect 30357 1683 30407 1707
rect 30693 1741 30743 1765
rect 30693 1707 30701 1741
rect 30735 1707 30743 1741
rect 30693 1683 30743 1707
rect 31029 1741 31079 1765
rect 31029 1707 31037 1741
rect 31071 1707 31079 1741
rect 31029 1683 31079 1707
rect 31365 1741 31415 1765
rect 31365 1707 31373 1741
rect 31407 1707 31415 1741
rect 31365 1683 31415 1707
rect 31701 1741 31751 1765
rect 31701 1707 31709 1741
rect 31743 1707 31751 1741
rect 31701 1683 31751 1707
rect 32037 1741 32087 1765
rect 32037 1707 32045 1741
rect 32079 1707 32087 1741
rect 32037 1683 32087 1707
rect 32373 1741 32423 1765
rect 32373 1707 32381 1741
rect 32415 1707 32423 1741
rect 32373 1683 32423 1707
rect 32709 1741 32759 1765
rect 32709 1707 32717 1741
rect 32751 1707 32759 1741
rect 32709 1683 32759 1707
rect 33045 1741 33095 1765
rect 33045 1707 33053 1741
rect 33087 1707 33095 1741
rect 33045 1683 33095 1707
rect 33381 1741 33431 1765
rect 33381 1707 33389 1741
rect 33423 1707 33431 1741
rect 33381 1683 33431 1707
rect 33717 1741 33767 1765
rect 33717 1707 33725 1741
rect 33759 1707 33767 1741
rect 33717 1683 33767 1707
rect 34053 1741 34103 1765
rect 34053 1707 34061 1741
rect 34095 1707 34103 1741
rect 34053 1683 34103 1707
rect 34389 1741 34439 1765
rect 34389 1707 34397 1741
rect 34431 1707 34439 1741
rect 34389 1683 34439 1707
rect 34725 1741 34775 1765
rect 34725 1707 34733 1741
rect 34767 1707 34775 1741
rect 34725 1683 34775 1707
rect 35061 1741 35111 1765
rect 35061 1707 35069 1741
rect 35103 1707 35111 1741
rect 35061 1683 35111 1707
rect 35397 1741 35447 1765
rect 35397 1707 35405 1741
rect 35439 1707 35447 1741
rect 35397 1683 35447 1707
rect 35733 1741 35783 1765
rect 35733 1707 35741 1741
rect 35775 1707 35783 1741
rect 35733 1683 35783 1707
rect 36069 1741 36119 1765
rect 36069 1707 36077 1741
rect 36111 1707 36119 1741
rect 36069 1683 36119 1707
rect 36405 1741 36455 1765
rect 36405 1707 36413 1741
rect 36447 1707 36455 1741
rect 36405 1683 36455 1707
rect 36741 1741 36791 1765
rect 36741 1707 36749 1741
rect 36783 1707 36791 1741
rect 36741 1683 36791 1707
rect 37077 1741 37127 1765
rect 37077 1707 37085 1741
rect 37119 1707 37127 1741
rect 37077 1683 37127 1707
rect 37413 1741 37463 1765
rect 37413 1707 37421 1741
rect 37455 1707 37463 1741
rect 37413 1683 37463 1707
rect 37749 1741 37799 1765
rect 37749 1707 37757 1741
rect 37791 1707 37799 1741
rect 37749 1683 37799 1707
rect 38085 1741 38135 1765
rect 38085 1707 38093 1741
rect 38127 1707 38135 1741
rect 38085 1683 38135 1707
rect 38421 1741 38471 1765
rect 38421 1707 38429 1741
rect 38463 1707 38471 1741
rect 38421 1683 38471 1707
rect 38757 1741 38807 1765
rect 38757 1707 38765 1741
rect 38799 1707 38807 1741
rect 38757 1683 38807 1707
rect 39093 1741 39143 1765
rect 39093 1707 39101 1741
rect 39135 1707 39143 1741
rect 39093 1683 39143 1707
rect 39429 1741 39479 1765
rect 39429 1707 39437 1741
rect 39471 1707 39479 1741
rect 39429 1683 39479 1707
rect 39765 1741 39815 1765
rect 39765 1707 39773 1741
rect 39807 1707 39815 1741
rect 39765 1683 39815 1707
rect 40101 1741 40151 1765
rect 40101 1707 40109 1741
rect 40143 1707 40151 1741
rect 40101 1683 40151 1707
rect 40437 1741 40487 1765
rect 40437 1707 40445 1741
rect 40479 1707 40487 1741
rect 40437 1683 40487 1707
rect 40773 1741 40823 1765
rect 40773 1707 40781 1741
rect 40815 1707 40823 1741
rect 40773 1683 40823 1707
rect 41109 1741 41159 1765
rect 41109 1707 41117 1741
rect 41151 1707 41159 1741
rect 41109 1683 41159 1707
rect 41445 1741 41495 1765
rect 41445 1707 41453 1741
rect 41487 1707 41495 1741
rect 41445 1683 41495 1707
rect 41781 1741 41831 1765
rect 41781 1707 41789 1741
rect 41823 1707 41831 1741
rect 41781 1683 41831 1707
rect 42117 1741 42167 1765
rect 42117 1707 42125 1741
rect 42159 1707 42167 1741
rect 42117 1683 42167 1707
rect 42453 1741 42503 1765
rect 42453 1707 42461 1741
rect 42495 1707 42503 1741
rect 42453 1683 42503 1707
rect 42789 1741 42839 1765
rect 42789 1707 42797 1741
rect 42831 1707 42839 1741
rect 42789 1683 42839 1707
rect 43125 1741 43175 1765
rect 43125 1707 43133 1741
rect 43167 1707 43175 1741
rect 43125 1683 43175 1707
rect 43461 1741 43511 1765
rect 43461 1707 43469 1741
rect 43503 1707 43511 1741
rect 43461 1683 43511 1707
rect 43797 1741 43847 1765
rect 43797 1707 43805 1741
rect 43839 1707 43847 1741
rect 43797 1683 43847 1707
rect 44133 1741 44183 1765
rect 44133 1707 44141 1741
rect 44175 1707 44183 1741
rect 44133 1683 44183 1707
rect 44469 1741 44519 1765
rect 44469 1707 44477 1741
rect 44511 1707 44519 1741
rect 44469 1683 44519 1707
rect 44805 1741 44855 1765
rect 44805 1707 44813 1741
rect 44847 1707 44855 1741
rect 44805 1683 44855 1707
rect 45141 1741 45191 1765
rect 45141 1707 45149 1741
rect 45183 1707 45191 1741
rect 45141 1683 45191 1707
rect 45477 1741 45527 1765
rect 45477 1707 45485 1741
rect 45519 1707 45527 1741
rect 45477 1683 45527 1707
rect 45813 1741 45863 1765
rect 45813 1707 45821 1741
rect 45855 1707 45863 1741
rect 45813 1683 45863 1707
rect 46149 1741 46199 1765
rect 46149 1707 46157 1741
rect 46191 1707 46199 1741
rect 46149 1683 46199 1707
rect 46485 1741 46535 1765
rect 46485 1707 46493 1741
rect 46527 1707 46535 1741
rect 46485 1683 46535 1707
rect 46821 1741 46871 1765
rect 46821 1707 46829 1741
rect 46863 1707 46871 1741
rect 46821 1683 46871 1707
rect 47157 1741 47207 1765
rect 47157 1707 47165 1741
rect 47199 1707 47207 1741
rect 47157 1683 47207 1707
rect 47493 1741 47543 1765
rect 47493 1707 47501 1741
rect 47535 1707 47543 1741
rect 47493 1683 47543 1707
rect 47829 1741 47879 1765
rect 47829 1707 47837 1741
rect 47871 1707 47879 1741
rect 47829 1683 47879 1707
rect 48165 1741 48215 1765
rect 48165 1707 48173 1741
rect 48207 1707 48215 1741
rect 48165 1683 48215 1707
rect 48501 1741 48551 1765
rect 48501 1707 48509 1741
rect 48543 1707 48551 1741
rect 48501 1683 48551 1707
rect 48837 1741 48887 1765
rect 48837 1707 48845 1741
rect 48879 1707 48887 1741
rect 48837 1683 48887 1707
rect 49173 1741 49223 1765
rect 49173 1707 49181 1741
rect 49215 1707 49223 1741
rect 49173 1683 49223 1707
rect 49509 1741 49559 1765
rect 49509 1707 49517 1741
rect 49551 1707 49559 1741
rect 49509 1683 49559 1707
rect 49845 1741 49895 1765
rect 49845 1707 49853 1741
rect 49887 1707 49895 1741
rect 49845 1683 49895 1707
rect 50181 1741 50231 1765
rect 50181 1707 50189 1741
rect 50223 1707 50231 1741
rect 50181 1683 50231 1707
rect 50517 1741 50567 1765
rect 50517 1707 50525 1741
rect 50559 1707 50567 1741
rect 50517 1683 50567 1707
rect 50853 1741 50903 1765
rect 50853 1707 50861 1741
rect 50895 1707 50903 1741
rect 50853 1683 50903 1707
rect 51189 1741 51239 1765
rect 51189 1707 51197 1741
rect 51231 1707 51239 1741
rect 51189 1683 51239 1707
rect 51525 1741 51575 1765
rect 51525 1707 51533 1741
rect 51567 1707 51575 1741
rect 51525 1683 51575 1707
rect 51861 1741 51911 1765
rect 51861 1707 51869 1741
rect 51903 1707 51911 1741
rect 51861 1683 51911 1707
rect 52197 1741 52247 1765
rect 52197 1707 52205 1741
rect 52239 1707 52247 1741
rect 52197 1683 52247 1707
rect 52533 1741 52583 1765
rect 52533 1707 52541 1741
rect 52575 1707 52583 1741
rect 52533 1683 52583 1707
rect 52869 1741 52919 1765
rect 52869 1707 52877 1741
rect 52911 1707 52919 1741
rect 52869 1683 52919 1707
rect 53205 1741 53255 1765
rect 53205 1707 53213 1741
rect 53247 1707 53255 1741
rect 53205 1683 53255 1707
rect 53541 1741 53591 1765
rect 53541 1707 53549 1741
rect 53583 1707 53591 1741
rect 53541 1683 53591 1707
rect 53877 1741 53927 1765
rect 53877 1707 53885 1741
rect 53919 1707 53927 1741
rect 53877 1683 53927 1707
rect 54213 1741 54263 1765
rect 54213 1707 54221 1741
rect 54255 1707 54263 1741
rect 54213 1683 54263 1707
rect 54549 1741 54599 1765
rect 54549 1707 54557 1741
rect 54591 1707 54599 1741
rect 54549 1683 54599 1707
rect 54885 1741 54935 1765
rect 54885 1707 54893 1741
rect 54927 1707 54935 1741
rect 54885 1683 54935 1707
rect 55221 1741 55271 1765
rect 55221 1707 55229 1741
rect 55263 1707 55271 1741
rect 55221 1683 55271 1707
rect 55557 1741 55607 1765
rect 55557 1707 55565 1741
rect 55599 1707 55607 1741
rect 55557 1683 55607 1707
rect 55893 1741 55943 1765
rect 55893 1707 55901 1741
rect 55935 1707 55943 1741
rect 55893 1683 55943 1707
rect 56229 1741 56279 1765
rect 56229 1707 56237 1741
rect 56271 1707 56279 1741
rect 56229 1683 56279 1707
rect 56565 1741 56615 1765
rect 56565 1707 56573 1741
rect 56607 1707 56615 1741
rect 56565 1683 56615 1707
rect 56901 1741 56951 1765
rect 56901 1707 56909 1741
rect 56943 1707 56951 1741
rect 56901 1683 56951 1707
rect 57237 1741 57287 1765
rect 57237 1707 57245 1741
rect 57279 1707 57287 1741
rect 57237 1683 57287 1707
rect 57573 1741 57623 1765
rect 57573 1707 57581 1741
rect 57615 1707 57623 1741
rect 57573 1683 57623 1707
rect 57909 1741 57959 1765
rect 57909 1707 57917 1741
rect 57951 1707 57959 1741
rect 57909 1683 57959 1707
rect 58245 1741 58295 1765
rect 58245 1707 58253 1741
rect 58287 1707 58295 1741
rect 58245 1683 58295 1707
rect 58581 1741 58631 1765
rect 58581 1707 58589 1741
rect 58623 1707 58631 1741
rect 58581 1683 58631 1707
rect 58917 1741 58967 1765
rect 58917 1707 58925 1741
rect 58959 1707 58967 1741
rect 58917 1683 58967 1707
rect 59253 1741 59303 1765
rect 59253 1707 59261 1741
rect 59295 1707 59303 1741
rect 59253 1683 59303 1707
rect 59589 1741 59639 1765
rect 59589 1707 59597 1741
rect 59631 1707 59639 1741
rect 59589 1683 59639 1707
rect 59925 1741 59975 1765
rect 59925 1707 59933 1741
rect 59967 1707 59975 1741
rect 59925 1683 59975 1707
rect 60261 1741 60311 1765
rect 60261 1707 60269 1741
rect 60303 1707 60311 1741
rect 60261 1683 60311 1707
rect 60597 1741 60647 1765
rect 60597 1707 60605 1741
rect 60639 1707 60647 1741
rect 60597 1683 60647 1707
rect 60933 1741 60983 1765
rect 60933 1707 60941 1741
rect 60975 1707 60983 1741
rect 60933 1683 60983 1707
rect 61269 1741 61319 1765
rect 61269 1707 61277 1741
rect 61311 1707 61319 1741
rect 61269 1683 61319 1707
rect 61605 1741 61655 1765
rect 61605 1707 61613 1741
rect 61647 1707 61655 1741
rect 61605 1683 61655 1707
rect 61941 1741 61991 1765
rect 61941 1707 61949 1741
rect 61983 1707 61991 1741
rect 61941 1683 61991 1707
rect 62277 1741 62327 1765
rect 62277 1707 62285 1741
rect 62319 1707 62327 1741
rect 62277 1683 62327 1707
rect 62613 1741 62663 1765
rect 62613 1707 62621 1741
rect 62655 1707 62663 1741
rect 62613 1683 62663 1707
rect 62949 1741 62999 1765
rect 62949 1707 62957 1741
rect 62991 1707 62999 1741
rect 62949 1683 62999 1707
rect 63285 1741 63335 1765
rect 63285 1707 63293 1741
rect 63327 1707 63335 1741
rect 63285 1683 63335 1707
rect 63621 1741 63671 1765
rect 63621 1707 63629 1741
rect 63663 1707 63671 1741
rect 63621 1683 63671 1707
rect 63957 1741 64007 1765
rect 63957 1707 63965 1741
rect 63999 1707 64007 1741
rect 63957 1683 64007 1707
rect 64293 1741 64343 1765
rect 64293 1707 64301 1741
rect 64335 1707 64343 1741
rect 64293 1683 64343 1707
rect 64629 1741 64679 1765
rect 64629 1707 64637 1741
rect 64671 1707 64679 1741
rect 64629 1683 64679 1707
rect 64965 1741 65015 1765
rect 64965 1707 64973 1741
rect 65007 1707 65015 1741
rect 64965 1683 65015 1707
rect 65301 1741 65351 1765
rect 65301 1707 65309 1741
rect 65343 1707 65351 1741
rect 65301 1683 65351 1707
rect 65637 1741 65687 1765
rect 65637 1707 65645 1741
rect 65679 1707 65687 1741
rect 65637 1683 65687 1707
rect 65973 1741 66023 1765
rect 65973 1707 65981 1741
rect 66015 1707 66023 1741
rect 65973 1683 66023 1707
rect 66309 1741 66359 1765
rect 66309 1707 66317 1741
rect 66351 1707 66359 1741
rect 66309 1683 66359 1707
rect 66645 1741 66695 1765
rect 66645 1707 66653 1741
rect 66687 1707 66695 1741
rect 66645 1683 66695 1707
rect 66981 1741 67031 1765
rect 66981 1707 66989 1741
rect 67023 1707 67031 1741
rect 66981 1683 67031 1707
rect 67317 1741 67367 1765
rect 67317 1707 67325 1741
rect 67359 1707 67367 1741
rect 67317 1683 67367 1707
rect 67653 1741 67703 1765
rect 67653 1707 67661 1741
rect 67695 1707 67703 1741
rect 67653 1683 67703 1707
rect 67989 1741 68039 1765
rect 67989 1707 67997 1741
rect 68031 1707 68039 1741
rect 67989 1683 68039 1707
rect 68325 1741 68375 1765
rect 68325 1707 68333 1741
rect 68367 1707 68375 1741
rect 68325 1683 68375 1707
rect 68661 1741 68711 1765
rect 68661 1707 68669 1741
rect 68703 1707 68711 1741
rect 68661 1683 68711 1707
rect 68997 1741 69047 1765
rect 68997 1707 69005 1741
rect 69039 1707 69047 1741
rect 68997 1683 69047 1707
rect 69333 1741 69383 1765
rect 69333 1707 69341 1741
rect 69375 1707 69383 1741
rect 69333 1683 69383 1707
rect 69669 1741 69719 1765
rect 69669 1707 69677 1741
rect 69711 1707 69719 1741
rect 69669 1683 69719 1707
rect 70005 1741 70055 1765
rect 70005 1707 70013 1741
rect 70047 1707 70055 1741
rect 70005 1683 70055 1707
rect 70341 1741 70391 1765
rect 70341 1707 70349 1741
rect 70383 1707 70391 1741
rect 70341 1683 70391 1707
rect 70677 1741 70727 1765
rect 70677 1707 70685 1741
rect 70719 1707 70727 1741
rect 70677 1683 70727 1707
rect 71013 1741 71063 1765
rect 71013 1707 71021 1741
rect 71055 1707 71063 1741
rect 71013 1683 71063 1707
rect 71349 1741 71399 1765
rect 71349 1707 71357 1741
rect 71391 1707 71399 1741
rect 71349 1683 71399 1707
rect 71685 1741 71735 1765
rect 71685 1707 71693 1741
rect 71727 1707 71735 1741
rect 71685 1683 71735 1707
rect 72021 1741 72071 1765
rect 72021 1707 72029 1741
rect 72063 1707 72071 1741
rect 72021 1683 72071 1707
rect 72357 1741 72407 1765
rect 72357 1707 72365 1741
rect 72399 1707 72407 1741
rect 72357 1683 72407 1707
rect 72693 1741 72743 1765
rect 72693 1707 72701 1741
rect 72735 1707 72743 1741
rect 72693 1683 72743 1707
rect 73029 1741 73079 1765
rect 73029 1707 73037 1741
rect 73071 1707 73079 1741
rect 73029 1683 73079 1707
rect 73365 1741 73415 1765
rect 73365 1707 73373 1741
rect 73407 1707 73415 1741
rect 73365 1683 73415 1707
rect 73701 1741 73751 1765
rect 73701 1707 73709 1741
rect 73743 1707 73751 1741
rect 73701 1683 73751 1707
rect 74037 1741 74087 1765
rect 74037 1707 74045 1741
rect 74079 1707 74087 1741
rect 74037 1683 74087 1707
rect 74373 1741 74423 1765
rect 74373 1707 74381 1741
rect 74415 1707 74423 1741
rect 74373 1683 74423 1707
rect 74709 1741 74759 1765
rect 74709 1707 74717 1741
rect 74751 1707 74759 1741
rect 74709 1683 74759 1707
rect 75045 1741 75095 1765
rect 75045 1707 75053 1741
rect 75087 1707 75095 1741
rect 75045 1683 75095 1707
rect 75381 1741 75431 1765
rect 75381 1707 75389 1741
rect 75423 1707 75431 1741
rect 75381 1683 75431 1707
rect 75717 1741 75767 1765
rect 75717 1707 75725 1741
rect 75759 1707 75767 1741
rect 75717 1683 75767 1707
rect 76053 1741 76103 1765
rect 76053 1707 76061 1741
rect 76095 1707 76103 1741
rect 76053 1683 76103 1707
rect 76389 1741 76439 1765
rect 76389 1707 76397 1741
rect 76431 1707 76439 1741
rect 76389 1683 76439 1707
rect 76725 1741 76775 1765
rect 76725 1707 76733 1741
rect 76767 1707 76775 1741
rect 76725 1683 76775 1707
rect 77061 1741 77111 1765
rect 77061 1707 77069 1741
rect 77103 1707 77111 1741
rect 77061 1683 77111 1707
rect 77397 1741 77447 1765
rect 77397 1707 77405 1741
rect 77439 1707 77447 1741
rect 77397 1683 77447 1707
rect 77733 1741 77783 1765
rect 77733 1707 77741 1741
rect 77775 1707 77783 1741
rect 77733 1683 77783 1707
rect 78069 1741 78119 1765
rect 78069 1707 78077 1741
rect 78111 1707 78119 1741
rect 78069 1683 78119 1707
rect 78405 1741 78455 1765
rect 78405 1707 78413 1741
rect 78447 1707 78455 1741
rect 78405 1683 78455 1707
rect 78741 1741 78791 1765
rect 78741 1707 78749 1741
rect 78783 1707 78791 1741
rect 78741 1683 78791 1707
rect 79077 1741 79127 1765
rect 79077 1707 79085 1741
rect 79119 1707 79127 1741
rect 79077 1683 79127 1707
rect 79413 1741 79463 1765
rect 79413 1707 79421 1741
rect 79455 1707 79463 1741
rect 79413 1683 79463 1707
rect 79749 1741 79799 1765
rect 79749 1707 79757 1741
rect 79791 1707 79799 1741
rect 79749 1683 79799 1707
rect 80085 1741 80135 1765
rect 80085 1707 80093 1741
rect 80127 1707 80135 1741
rect 80085 1683 80135 1707
rect 80421 1741 80471 1765
rect 80421 1707 80429 1741
rect 80463 1707 80471 1741
rect 80421 1683 80471 1707
rect 80757 1741 80807 1765
rect 80757 1707 80765 1741
rect 80799 1707 80807 1741
rect 80757 1683 80807 1707
rect 81093 1741 81143 1765
rect 81093 1707 81101 1741
rect 81135 1707 81143 1741
rect 81093 1683 81143 1707
rect 81429 1741 81479 1765
rect 81429 1707 81437 1741
rect 81471 1707 81479 1741
rect 81429 1683 81479 1707
rect 81765 1741 81815 1765
rect 81765 1707 81773 1741
rect 81807 1707 81815 1741
rect 81765 1683 81815 1707
rect 82101 1741 82151 1765
rect 82101 1707 82109 1741
rect 82143 1707 82151 1741
rect 82101 1683 82151 1707
rect 82437 1741 82487 1765
rect 82437 1707 82445 1741
rect 82479 1707 82487 1741
rect 82437 1683 82487 1707
rect 82773 1741 82823 1765
rect 82773 1707 82781 1741
rect 82815 1707 82823 1741
rect 82773 1683 82823 1707
rect 83109 1741 83159 1765
rect 83109 1707 83117 1741
rect 83151 1707 83159 1741
rect 83109 1683 83159 1707
rect 83445 1741 83495 1765
rect 83445 1707 83453 1741
rect 83487 1707 83495 1741
rect 83445 1683 83495 1707
rect 83781 1741 83831 1765
rect 83781 1707 83789 1741
rect 83823 1707 83831 1741
rect 83781 1683 83831 1707
rect 84117 1741 84167 1765
rect 84117 1707 84125 1741
rect 84159 1707 84167 1741
rect 84117 1683 84167 1707
rect 84453 1741 84503 1765
rect 84453 1707 84461 1741
rect 84495 1707 84503 1741
rect 84453 1683 84503 1707
rect 84789 1741 84839 1765
rect 84789 1707 84797 1741
rect 84831 1707 84839 1741
rect 84789 1683 84839 1707
rect 85125 1741 85175 1765
rect 85125 1707 85133 1741
rect 85167 1707 85175 1741
rect 85125 1683 85175 1707
rect 85461 1741 85511 1765
rect 85461 1707 85469 1741
rect 85503 1707 85511 1741
rect 85461 1683 85511 1707
rect 85797 1741 85847 1765
rect 85797 1707 85805 1741
rect 85839 1707 85847 1741
rect 85797 1683 85847 1707
rect 86133 1741 86183 1765
rect 86133 1707 86141 1741
rect 86175 1707 86183 1741
rect 86133 1683 86183 1707
rect 86469 1741 86519 1765
rect 86469 1707 86477 1741
rect 86511 1707 86519 1741
rect 86469 1683 86519 1707
rect 86805 1741 86855 1765
rect 86805 1707 86813 1741
rect 86847 1707 86855 1741
rect 86805 1683 86855 1707
rect 87141 1741 87191 1765
rect 87141 1707 87149 1741
rect 87183 1707 87191 1741
rect 87141 1683 87191 1707
rect 87477 1741 87527 1765
rect 87477 1707 87485 1741
rect 87519 1707 87527 1741
rect 87477 1683 87527 1707
rect 87813 1741 87863 1765
rect 87813 1707 87821 1741
rect 87855 1707 87863 1741
rect 87813 1683 87863 1707
rect 88149 1741 88199 1765
rect 88149 1707 88157 1741
rect 88191 1707 88199 1741
rect 88149 1683 88199 1707
rect 88485 1741 88535 1765
rect 88485 1707 88493 1741
rect 88527 1707 88535 1741
rect 88485 1683 88535 1707
rect 88821 1741 88871 1765
rect 88821 1707 88829 1741
rect 88863 1707 88871 1741
rect 88821 1683 88871 1707
rect 89157 1741 89207 1765
rect 89157 1707 89165 1741
rect 89199 1707 89207 1741
rect 89157 1683 89207 1707
rect 89493 1741 89543 1765
rect 89493 1707 89501 1741
rect 89535 1707 89543 1741
rect 89493 1683 89543 1707
rect 89829 1741 89879 1765
rect 89829 1707 89837 1741
rect 89871 1707 89879 1741
rect 89829 1683 89879 1707
rect 90165 1741 90215 1765
rect 90165 1707 90173 1741
rect 90207 1707 90215 1741
rect 90165 1683 90215 1707
rect 90501 1741 90551 1765
rect 90501 1707 90509 1741
rect 90543 1707 90551 1741
rect 90501 1683 90551 1707
rect 90837 1741 90887 1765
rect 90837 1707 90845 1741
rect 90879 1707 90887 1741
rect 90837 1683 90887 1707
rect 91173 1741 91223 1765
rect 91173 1707 91181 1741
rect 91215 1707 91223 1741
rect 91173 1683 91223 1707
rect 91509 1741 91559 1765
rect 91509 1707 91517 1741
rect 91551 1707 91559 1741
rect 91509 1683 91559 1707
rect 91845 1741 91895 1765
rect 91845 1707 91853 1741
rect 91887 1707 91895 1741
rect 91845 1683 91895 1707
rect 92181 1741 92231 1765
rect 92181 1707 92189 1741
rect 92223 1707 92231 1741
rect 92181 1683 92231 1707
rect 92517 1741 92567 1765
rect 92517 1707 92525 1741
rect 92559 1707 92567 1741
rect 92517 1683 92567 1707
rect 92853 1741 92903 1765
rect 92853 1707 92861 1741
rect 92895 1707 92903 1741
rect 92853 1683 92903 1707
rect 93189 1741 93239 1765
rect 93189 1707 93197 1741
rect 93231 1707 93239 1741
rect 93189 1683 93239 1707
rect 93525 1741 93575 1765
rect 93525 1707 93533 1741
rect 93567 1707 93575 1741
rect 93525 1683 93575 1707
rect 93861 1741 93911 1765
rect 93861 1707 93869 1741
rect 93903 1707 93911 1741
rect 93861 1683 93911 1707
rect 94197 1741 94247 1765
rect 94197 1707 94205 1741
rect 94239 1707 94247 1741
rect 94197 1683 94247 1707
rect 94533 1741 94583 1765
rect 94533 1707 94541 1741
rect 94575 1707 94583 1741
rect 94533 1683 94583 1707
rect 94869 1741 94919 1765
rect 94869 1707 94877 1741
rect 94911 1707 94919 1741
rect 94869 1683 94919 1707
rect 95205 1741 95255 1765
rect 95205 1707 95213 1741
rect 95247 1707 95255 1741
rect 95205 1683 95255 1707
rect 95541 1741 95591 1765
rect 95541 1707 95549 1741
rect 95583 1707 95591 1741
rect 95541 1683 95591 1707
rect 95877 1741 95927 1765
rect 95877 1707 95885 1741
rect 95919 1707 95927 1741
rect 95877 1683 95927 1707
rect 96213 1741 96263 1765
rect 96213 1707 96221 1741
rect 96255 1707 96263 1741
rect 96213 1683 96263 1707
rect 96549 1741 96599 1765
rect 96549 1707 96557 1741
rect 96591 1707 96599 1741
rect 96549 1683 96599 1707
rect 96885 1741 96935 1765
rect 96885 1707 96893 1741
rect 96927 1707 96935 1741
rect 96885 1683 96935 1707
rect 97221 1741 97271 1765
rect 97221 1707 97229 1741
rect 97263 1707 97271 1741
rect 97221 1683 97271 1707
rect 97557 1741 97607 1765
rect 97557 1707 97565 1741
rect 97599 1707 97607 1741
rect 97557 1683 97607 1707
rect 97893 1741 97943 1765
rect 97893 1707 97901 1741
rect 97935 1707 97943 1741
rect 97893 1683 97943 1707
rect 98229 1741 98279 1765
rect 98229 1707 98237 1741
rect 98271 1707 98279 1741
rect 98229 1683 98279 1707
rect 98565 1741 98615 1765
rect 98565 1707 98573 1741
rect 98607 1707 98615 1741
rect 98565 1683 98615 1707
rect 98901 1741 98951 1765
rect 98901 1707 98909 1741
rect 98943 1707 98951 1741
rect 98901 1683 98951 1707
rect 99237 1741 99287 1765
rect 99237 1707 99245 1741
rect 99279 1707 99287 1741
rect 99237 1683 99287 1707
rect 99573 1741 99623 1765
rect 99573 1707 99581 1741
rect 99615 1707 99623 1741
rect 99573 1683 99623 1707
rect 99909 1741 99959 1765
rect 99909 1707 99917 1741
rect 99951 1707 99959 1741
rect 99909 1683 99959 1707
rect 100245 1741 100295 1765
rect 100245 1707 100253 1741
rect 100287 1707 100295 1741
rect 100245 1683 100295 1707
rect 100581 1741 100631 1765
rect 100581 1707 100589 1741
rect 100623 1707 100631 1741
rect 100581 1683 100631 1707
rect 100917 1741 100967 1765
rect 100917 1707 100925 1741
rect 100959 1707 100967 1741
rect 100917 1683 100967 1707
rect 101253 1741 101303 1765
rect 101253 1707 101261 1741
rect 101295 1707 101303 1741
rect 101253 1683 101303 1707
rect 101589 1741 101639 1765
rect 101589 1707 101597 1741
rect 101631 1707 101639 1741
rect 101589 1683 101639 1707
rect 101925 1741 101975 1765
rect 101925 1707 101933 1741
rect 101967 1707 101975 1741
rect 101925 1683 101975 1707
rect 102261 1741 102311 1765
rect 102261 1707 102269 1741
rect 102303 1707 102311 1741
rect 102261 1683 102311 1707
rect 102597 1741 102647 1765
rect 102597 1707 102605 1741
rect 102639 1707 102647 1741
rect 102597 1683 102647 1707
rect 102933 1741 102983 1765
rect 102933 1707 102941 1741
rect 102975 1707 102983 1741
rect 102933 1683 102983 1707
rect 103269 1741 103319 1765
rect 103269 1707 103277 1741
rect 103311 1707 103319 1741
rect 103269 1683 103319 1707
rect 103605 1741 103655 1765
rect 103605 1707 103613 1741
rect 103647 1707 103655 1741
rect 103605 1683 103655 1707
rect 103941 1741 103991 1765
rect 103941 1707 103949 1741
rect 103983 1707 103991 1741
rect 103941 1683 103991 1707
rect 104277 1741 104327 1765
rect 104277 1707 104285 1741
rect 104319 1707 104327 1741
rect 104277 1683 104327 1707
rect 104613 1741 104663 1765
rect 104613 1707 104621 1741
rect 104655 1707 104663 1741
rect 104613 1683 104663 1707
rect 104949 1741 104999 1765
rect 104949 1707 104957 1741
rect 104991 1707 104999 1741
rect 104949 1683 104999 1707
rect 105285 1741 105335 1765
rect 105285 1707 105293 1741
rect 105327 1707 105335 1741
rect 105285 1683 105335 1707
rect 105621 1741 105671 1765
rect 105621 1707 105629 1741
rect 105663 1707 105671 1741
rect 105621 1683 105671 1707
rect 105957 1741 106007 1765
rect 105957 1707 105965 1741
rect 105999 1707 106007 1741
rect 105957 1683 106007 1707
rect 106293 1741 106343 1765
rect 106293 1707 106301 1741
rect 106335 1707 106343 1741
rect 106293 1683 106343 1707
rect 106629 1741 106679 1765
rect 106629 1707 106637 1741
rect 106671 1707 106679 1741
rect 106629 1683 106679 1707
rect 106965 1741 107015 1765
rect 106965 1707 106973 1741
rect 107007 1707 107015 1741
rect 106965 1683 107015 1707
rect 107301 1741 107351 1765
rect 107301 1707 107309 1741
rect 107343 1707 107351 1741
rect 107301 1683 107351 1707
rect 107637 1741 107687 1765
rect 107637 1707 107645 1741
rect 107679 1707 107687 1741
rect 107637 1683 107687 1707
rect 107973 1741 108023 1765
rect 107973 1707 107981 1741
rect 108015 1707 108023 1741
rect 107973 1683 108023 1707
rect 108309 1741 108359 1765
rect 108309 1707 108317 1741
rect 108351 1707 108359 1741
rect 108309 1683 108359 1707
rect 108645 1741 108695 1765
rect 108645 1707 108653 1741
rect 108687 1707 108695 1741
rect 108645 1683 108695 1707
rect 108981 1741 109031 1765
rect 108981 1707 108989 1741
rect 109023 1707 109031 1741
rect 108981 1683 109031 1707
rect 109317 1741 109367 1765
rect 109317 1707 109325 1741
rect 109359 1707 109367 1741
rect 109317 1683 109367 1707
rect 109653 1741 109703 1765
rect 109653 1707 109661 1741
rect 109695 1707 109703 1741
rect 109653 1683 109703 1707
rect 109989 1741 110039 1765
rect 109989 1707 109997 1741
rect 110031 1707 110039 1741
rect 109989 1683 110039 1707
rect 110325 1741 110375 1765
rect 110325 1707 110333 1741
rect 110367 1707 110375 1741
rect 110325 1683 110375 1707
rect 110661 1741 110711 1765
rect 110661 1707 110669 1741
rect 110703 1707 110711 1741
rect 110661 1683 110711 1707
rect 110997 1741 111047 1765
rect 110997 1707 111005 1741
rect 111039 1707 111047 1741
rect 110997 1683 111047 1707
rect 111333 1741 111383 1765
rect 111333 1707 111341 1741
rect 111375 1707 111383 1741
rect 111333 1683 111383 1707
rect 111669 1741 111719 1765
rect 111669 1707 111677 1741
rect 111711 1707 111719 1741
rect 111669 1683 111719 1707
rect 112005 1741 112055 1765
rect 112005 1707 112013 1741
rect 112047 1707 112055 1741
rect 112005 1683 112055 1707
rect 112341 1741 112391 1765
rect 112341 1707 112349 1741
rect 112383 1707 112391 1741
rect 112341 1683 112391 1707
rect 112677 1741 112727 1765
rect 112677 1707 112685 1741
rect 112719 1707 112727 1741
rect 112677 1683 112727 1707
rect 113013 1741 113063 1765
rect 113013 1707 113021 1741
rect 113055 1707 113063 1741
rect 113013 1683 113063 1707
rect 113349 1741 113399 1765
rect 113349 1707 113357 1741
rect 113391 1707 113399 1741
rect 113349 1683 113399 1707
rect 113685 1741 113735 1765
rect 113685 1707 113693 1741
rect 113727 1707 113735 1741
rect 113685 1683 113735 1707
rect 114021 1741 114071 1765
rect 114021 1707 114029 1741
rect 114063 1707 114071 1741
rect 114021 1683 114071 1707
rect 114357 1741 114407 1765
rect 114357 1707 114365 1741
rect 114399 1707 114407 1741
rect 114357 1683 114407 1707
rect 114693 1741 114743 1765
rect 114693 1707 114701 1741
rect 114735 1707 114743 1741
rect 114693 1683 114743 1707
rect 115029 1741 115079 1765
rect 115029 1707 115037 1741
rect 115071 1707 115079 1741
rect 115029 1683 115079 1707
rect 115365 1741 115415 1765
rect 115365 1707 115373 1741
rect 115407 1707 115415 1741
rect 115365 1683 115415 1707
rect 115701 1741 115751 1765
rect 115701 1707 115709 1741
rect 115743 1707 115751 1741
rect 115701 1683 115751 1707
rect 116037 1741 116087 1765
rect 116037 1707 116045 1741
rect 116079 1707 116087 1741
rect 116037 1683 116087 1707
rect 116373 1741 116423 1765
rect 116373 1707 116381 1741
rect 116415 1707 116423 1741
rect 116373 1683 116423 1707
rect 116709 1741 116759 1765
rect 116709 1707 116717 1741
rect 116751 1707 116759 1741
rect 116709 1683 116759 1707
rect 117045 1741 117095 1765
rect 117045 1707 117053 1741
rect 117087 1707 117095 1741
rect 117045 1683 117095 1707
rect 117381 1741 117431 1765
rect 117381 1707 117389 1741
rect 117423 1707 117431 1741
rect 117381 1683 117431 1707
rect 117717 1741 117767 1765
rect 117717 1707 117725 1741
rect 117759 1707 117767 1741
rect 117717 1683 117767 1707
rect 118053 1741 118103 1765
rect 118053 1707 118061 1741
rect 118095 1707 118103 1741
rect 118053 1683 118103 1707
rect 118389 1741 118439 1765
rect 118389 1707 118397 1741
rect 118431 1707 118439 1741
rect 118389 1683 118439 1707
rect 118725 1741 118775 1765
rect 118725 1707 118733 1741
rect 118767 1707 118775 1741
rect 118725 1683 118775 1707
rect 119061 1741 119111 1765
rect 119061 1707 119069 1741
rect 119103 1707 119111 1741
rect 119061 1683 119111 1707
rect 119397 1741 119447 1765
rect 119397 1707 119405 1741
rect 119439 1707 119447 1741
rect 119397 1683 119447 1707
rect 119733 1741 119783 1765
rect 119733 1707 119741 1741
rect 119775 1707 119783 1741
rect 119733 1683 119783 1707
rect 120069 1741 120119 1765
rect 120069 1707 120077 1741
rect 120111 1707 120119 1741
rect 120069 1683 120119 1707
rect 120405 1741 120455 1765
rect 120405 1707 120413 1741
rect 120447 1707 120455 1741
rect 120405 1683 120455 1707
rect 120741 1741 120791 1765
rect 120741 1707 120749 1741
rect 120783 1707 120791 1741
rect 120741 1683 120791 1707
rect 121077 1741 121127 1765
rect 121077 1707 121085 1741
rect 121119 1707 121127 1741
rect 121077 1683 121127 1707
rect 121413 1741 121463 1765
rect 121413 1707 121421 1741
rect 121455 1707 121463 1741
rect 121413 1683 121463 1707
rect 121749 1741 121799 1765
rect 121749 1707 121757 1741
rect 121791 1707 121799 1741
rect 121749 1683 121799 1707
rect 122085 1741 122135 1765
rect 122085 1707 122093 1741
rect 122127 1707 122135 1741
rect 122085 1683 122135 1707
rect 122421 1741 122471 1765
rect 122421 1707 122429 1741
rect 122463 1707 122471 1741
rect 122421 1683 122471 1707
rect 122757 1741 122807 1765
rect 122757 1707 122765 1741
rect 122799 1707 122807 1741
rect 122757 1683 122807 1707
rect 123093 1741 123143 1765
rect 123093 1707 123101 1741
rect 123135 1707 123143 1741
rect 123093 1683 123143 1707
rect 123429 1741 123479 1765
rect 123429 1707 123437 1741
rect 123471 1707 123479 1741
rect 123429 1683 123479 1707
rect 123765 1741 123815 1765
rect 123765 1707 123773 1741
rect 123807 1707 123815 1741
rect 123765 1683 123815 1707
rect 124101 1741 124151 1765
rect 124101 1707 124109 1741
rect 124143 1707 124151 1741
rect 124101 1683 124151 1707
rect 124437 1741 124487 1765
rect 124437 1707 124445 1741
rect 124479 1707 124487 1741
rect 124437 1683 124487 1707
rect 124773 1741 124823 1765
rect 124773 1707 124781 1741
rect 124815 1707 124823 1741
rect 124773 1683 124823 1707
rect 125109 1741 125159 1765
rect 125109 1707 125117 1741
rect 125151 1707 125159 1741
rect 125109 1683 125159 1707
rect 125445 1741 125495 1765
rect 125445 1707 125453 1741
rect 125487 1707 125495 1741
rect 125445 1683 125495 1707
rect 125781 1741 125831 1765
rect 125781 1707 125789 1741
rect 125823 1707 125831 1741
rect 125781 1683 125831 1707
rect 126117 1741 126167 1765
rect 126117 1707 126125 1741
rect 126159 1707 126167 1741
rect 126117 1683 126167 1707
rect 126453 1741 126503 1765
rect 126453 1707 126461 1741
rect 126495 1707 126503 1741
rect 126453 1683 126503 1707
rect 126789 1741 126839 1765
rect 126789 1707 126797 1741
rect 126831 1707 126839 1741
rect 126789 1683 126839 1707
rect 127125 1741 127175 1765
rect 127125 1707 127133 1741
rect 127167 1707 127175 1741
rect 127125 1683 127175 1707
rect 127461 1741 127511 1765
rect 127461 1707 127469 1741
rect 127503 1707 127511 1741
rect 127461 1683 127511 1707
rect 127797 1741 127847 1765
rect 127797 1707 127805 1741
rect 127839 1707 127847 1741
rect 127797 1683 127847 1707
rect 128133 1741 128183 1765
rect 128133 1707 128141 1741
rect 128175 1707 128183 1741
rect 128133 1683 128183 1707
rect 128469 1741 128519 1765
rect 128469 1707 128477 1741
rect 128511 1707 128519 1741
rect 128469 1683 128519 1707
rect 128805 1741 128855 1765
rect 128805 1707 128813 1741
rect 128847 1707 128855 1741
rect 128805 1683 128855 1707
rect 129141 1741 129191 1765
rect 129141 1707 129149 1741
rect 129183 1707 129191 1741
rect 129141 1683 129191 1707
rect 129477 1741 129527 1765
rect 129477 1707 129485 1741
rect 129519 1707 129527 1741
rect 129477 1683 129527 1707
rect 129813 1741 129863 1765
rect 129813 1707 129821 1741
rect 129855 1707 129863 1741
rect 129813 1683 129863 1707
rect 130149 1741 130199 1765
rect 130149 1707 130157 1741
rect 130191 1707 130199 1741
rect 130149 1683 130199 1707
rect 130485 1741 130535 1765
rect 130485 1707 130493 1741
rect 130527 1707 130535 1741
rect 130485 1683 130535 1707
rect 130821 1741 130871 1765
rect 130821 1707 130829 1741
rect 130863 1707 130871 1741
rect 130821 1683 130871 1707
rect 131157 1741 131207 1765
rect 131157 1707 131165 1741
rect 131199 1707 131207 1741
rect 131157 1683 131207 1707
rect 131493 1741 131543 1765
rect 131493 1707 131501 1741
rect 131535 1707 131543 1741
rect 131493 1683 131543 1707
rect 131829 1741 131879 1765
rect 131829 1707 131837 1741
rect 131871 1707 131879 1741
rect 131829 1683 131879 1707
rect 132165 1741 132215 1765
rect 132165 1707 132173 1741
rect 132207 1707 132215 1741
rect 132165 1683 132215 1707
rect 132501 1741 132551 1765
rect 132501 1707 132509 1741
rect 132543 1707 132551 1741
rect 132501 1683 132551 1707
rect 132837 1741 132887 1765
rect 132837 1707 132845 1741
rect 132879 1707 132887 1741
rect 132837 1683 132887 1707
rect 133173 1741 133223 1765
rect 133173 1707 133181 1741
rect 133215 1707 133223 1741
rect 133173 1683 133223 1707
rect 133509 1741 133559 1765
rect 133509 1707 133517 1741
rect 133551 1707 133559 1741
rect 133509 1683 133559 1707
rect 133845 1741 133895 1765
rect 133845 1707 133853 1741
rect 133887 1707 133895 1741
rect 133845 1683 133895 1707
rect 134181 1741 134231 1765
rect 134181 1707 134189 1741
rect 134223 1707 134231 1741
rect 134181 1683 134231 1707
<< nsubdiffcont >>
rect 2141 81456 2175 81490
rect 2477 81456 2511 81490
rect 2813 81456 2847 81490
rect 3149 81456 3183 81490
rect 3485 81456 3519 81490
rect 3821 81456 3855 81490
rect 4157 81456 4191 81490
rect 4493 81456 4527 81490
rect 4829 81456 4863 81490
rect 5165 81456 5199 81490
rect 5501 81456 5535 81490
rect 5837 81456 5871 81490
rect 6173 81456 6207 81490
rect 6509 81456 6543 81490
rect 6845 81456 6879 81490
rect 7181 81456 7215 81490
rect 7517 81456 7551 81490
rect 7853 81456 7887 81490
rect 8189 81456 8223 81490
rect 8525 81456 8559 81490
rect 8861 81456 8895 81490
rect 9197 81456 9231 81490
rect 9533 81456 9567 81490
rect 9869 81456 9903 81490
rect 10205 81456 10239 81490
rect 10541 81456 10575 81490
rect 10877 81456 10911 81490
rect 11213 81456 11247 81490
rect 11549 81456 11583 81490
rect 11885 81456 11919 81490
rect 12221 81456 12255 81490
rect 12557 81456 12591 81490
rect 12893 81456 12927 81490
rect 13229 81456 13263 81490
rect 13565 81456 13599 81490
rect 13901 81456 13935 81490
rect 14237 81456 14271 81490
rect 14573 81456 14607 81490
rect 14909 81456 14943 81490
rect 15245 81456 15279 81490
rect 15581 81456 15615 81490
rect 15917 81456 15951 81490
rect 16253 81456 16287 81490
rect 16589 81456 16623 81490
rect 16925 81456 16959 81490
rect 17261 81456 17295 81490
rect 17597 81456 17631 81490
rect 17933 81456 17967 81490
rect 18269 81456 18303 81490
rect 18605 81456 18639 81490
rect 18941 81456 18975 81490
rect 19277 81456 19311 81490
rect 19613 81456 19647 81490
rect 19949 81456 19983 81490
rect 20285 81456 20319 81490
rect 20621 81456 20655 81490
rect 20957 81456 20991 81490
rect 21293 81456 21327 81490
rect 21629 81456 21663 81490
rect 21965 81456 21999 81490
rect 22301 81456 22335 81490
rect 22637 81456 22671 81490
rect 22973 81456 23007 81490
rect 23309 81456 23343 81490
rect 23645 81456 23679 81490
rect 23981 81456 24015 81490
rect 24317 81456 24351 81490
rect 24653 81456 24687 81490
rect 24989 81456 25023 81490
rect 25325 81456 25359 81490
rect 25661 81456 25695 81490
rect 25997 81456 26031 81490
rect 26333 81456 26367 81490
rect 26669 81456 26703 81490
rect 27005 81456 27039 81490
rect 27341 81456 27375 81490
rect 27677 81456 27711 81490
rect 28013 81456 28047 81490
rect 28349 81456 28383 81490
rect 28685 81456 28719 81490
rect 29021 81456 29055 81490
rect 29357 81456 29391 81490
rect 29693 81456 29727 81490
rect 30029 81456 30063 81490
rect 30365 81456 30399 81490
rect 30701 81456 30735 81490
rect 31037 81456 31071 81490
rect 31373 81456 31407 81490
rect 31709 81456 31743 81490
rect 32045 81456 32079 81490
rect 32381 81456 32415 81490
rect 32717 81456 32751 81490
rect 33053 81456 33087 81490
rect 33389 81456 33423 81490
rect 33725 81456 33759 81490
rect 34061 81456 34095 81490
rect 34397 81456 34431 81490
rect 34733 81456 34767 81490
rect 35069 81456 35103 81490
rect 35405 81456 35439 81490
rect 35741 81456 35775 81490
rect 36077 81456 36111 81490
rect 36413 81456 36447 81490
rect 36749 81456 36783 81490
rect 37085 81456 37119 81490
rect 37421 81456 37455 81490
rect 37757 81456 37791 81490
rect 38093 81456 38127 81490
rect 38429 81456 38463 81490
rect 38765 81456 38799 81490
rect 39101 81456 39135 81490
rect 39437 81456 39471 81490
rect 39773 81456 39807 81490
rect 40109 81456 40143 81490
rect 40445 81456 40479 81490
rect 40781 81456 40815 81490
rect 41117 81456 41151 81490
rect 41453 81456 41487 81490
rect 41789 81456 41823 81490
rect 42125 81456 42159 81490
rect 42461 81456 42495 81490
rect 42797 81456 42831 81490
rect 43133 81456 43167 81490
rect 43469 81456 43503 81490
rect 43805 81456 43839 81490
rect 44141 81456 44175 81490
rect 44477 81456 44511 81490
rect 44813 81456 44847 81490
rect 45149 81456 45183 81490
rect 45485 81456 45519 81490
rect 45821 81456 45855 81490
rect 46157 81456 46191 81490
rect 46493 81456 46527 81490
rect 46829 81456 46863 81490
rect 47165 81456 47199 81490
rect 47501 81456 47535 81490
rect 47837 81456 47871 81490
rect 48173 81456 48207 81490
rect 48509 81456 48543 81490
rect 48845 81456 48879 81490
rect 49181 81456 49215 81490
rect 49517 81456 49551 81490
rect 49853 81456 49887 81490
rect 50189 81456 50223 81490
rect 50525 81456 50559 81490
rect 50861 81456 50895 81490
rect 51197 81456 51231 81490
rect 51533 81456 51567 81490
rect 51869 81456 51903 81490
rect 52205 81456 52239 81490
rect 52541 81456 52575 81490
rect 52877 81456 52911 81490
rect 53213 81456 53247 81490
rect 53549 81456 53583 81490
rect 53885 81456 53919 81490
rect 54221 81456 54255 81490
rect 54557 81456 54591 81490
rect 54893 81456 54927 81490
rect 55229 81456 55263 81490
rect 55565 81456 55599 81490
rect 55901 81456 55935 81490
rect 56237 81456 56271 81490
rect 56573 81456 56607 81490
rect 56909 81456 56943 81490
rect 57245 81456 57279 81490
rect 57581 81456 57615 81490
rect 57917 81456 57951 81490
rect 58253 81456 58287 81490
rect 58589 81456 58623 81490
rect 58925 81456 58959 81490
rect 59261 81456 59295 81490
rect 59597 81456 59631 81490
rect 59933 81456 59967 81490
rect 60269 81456 60303 81490
rect 60605 81456 60639 81490
rect 60941 81456 60975 81490
rect 61277 81456 61311 81490
rect 61613 81456 61647 81490
rect 61949 81456 61983 81490
rect 62285 81456 62319 81490
rect 62621 81456 62655 81490
rect 62957 81456 62991 81490
rect 63293 81456 63327 81490
rect 63629 81456 63663 81490
rect 63965 81456 63999 81490
rect 64301 81456 64335 81490
rect 64637 81456 64671 81490
rect 64973 81456 65007 81490
rect 65309 81456 65343 81490
rect 65645 81456 65679 81490
rect 65981 81456 66015 81490
rect 66317 81456 66351 81490
rect 66653 81456 66687 81490
rect 66989 81456 67023 81490
rect 67325 81456 67359 81490
rect 67661 81456 67695 81490
rect 67997 81456 68031 81490
rect 68333 81456 68367 81490
rect 68669 81456 68703 81490
rect 69005 81456 69039 81490
rect 69341 81456 69375 81490
rect 69677 81456 69711 81490
rect 70013 81456 70047 81490
rect 70349 81456 70383 81490
rect 70685 81456 70719 81490
rect 71021 81456 71055 81490
rect 71357 81456 71391 81490
rect 71693 81456 71727 81490
rect 72029 81456 72063 81490
rect 72365 81456 72399 81490
rect 72701 81456 72735 81490
rect 73037 81456 73071 81490
rect 73373 81456 73407 81490
rect 73709 81456 73743 81490
rect 74045 81456 74079 81490
rect 74381 81456 74415 81490
rect 74717 81456 74751 81490
rect 75053 81456 75087 81490
rect 75389 81456 75423 81490
rect 75725 81456 75759 81490
rect 76061 81456 76095 81490
rect 76397 81456 76431 81490
rect 76733 81456 76767 81490
rect 77069 81456 77103 81490
rect 77405 81456 77439 81490
rect 77741 81456 77775 81490
rect 78077 81456 78111 81490
rect 78413 81456 78447 81490
rect 78749 81456 78783 81490
rect 79085 81456 79119 81490
rect 79421 81456 79455 81490
rect 79757 81456 79791 81490
rect 80093 81456 80127 81490
rect 80429 81456 80463 81490
rect 80765 81456 80799 81490
rect 81101 81456 81135 81490
rect 81437 81456 81471 81490
rect 81773 81456 81807 81490
rect 82109 81456 82143 81490
rect 82445 81456 82479 81490
rect 82781 81456 82815 81490
rect 83117 81456 83151 81490
rect 83453 81456 83487 81490
rect 83789 81456 83823 81490
rect 84125 81456 84159 81490
rect 84461 81456 84495 81490
rect 84797 81456 84831 81490
rect 85133 81456 85167 81490
rect 85469 81456 85503 81490
rect 85805 81456 85839 81490
rect 86141 81456 86175 81490
rect 86477 81456 86511 81490
rect 86813 81456 86847 81490
rect 87149 81456 87183 81490
rect 87485 81456 87519 81490
rect 87821 81456 87855 81490
rect 88157 81456 88191 81490
rect 88493 81456 88527 81490
rect 88829 81456 88863 81490
rect 89165 81456 89199 81490
rect 89501 81456 89535 81490
rect 89837 81456 89871 81490
rect 90173 81456 90207 81490
rect 90509 81456 90543 81490
rect 90845 81456 90879 81490
rect 91181 81456 91215 81490
rect 91517 81456 91551 81490
rect 91853 81456 91887 81490
rect 92189 81456 92223 81490
rect 92525 81456 92559 81490
rect 92861 81456 92895 81490
rect 93197 81456 93231 81490
rect 93533 81456 93567 81490
rect 93869 81456 93903 81490
rect 94205 81456 94239 81490
rect 94541 81456 94575 81490
rect 94877 81456 94911 81490
rect 95213 81456 95247 81490
rect 95549 81456 95583 81490
rect 95885 81456 95919 81490
rect 96221 81456 96255 81490
rect 96557 81456 96591 81490
rect 96893 81456 96927 81490
rect 97229 81456 97263 81490
rect 97565 81456 97599 81490
rect 97901 81456 97935 81490
rect 98237 81456 98271 81490
rect 98573 81456 98607 81490
rect 98909 81456 98943 81490
rect 99245 81456 99279 81490
rect 99581 81456 99615 81490
rect 99917 81456 99951 81490
rect 100253 81456 100287 81490
rect 100589 81456 100623 81490
rect 100925 81456 100959 81490
rect 101261 81456 101295 81490
rect 101597 81456 101631 81490
rect 101933 81456 101967 81490
rect 102269 81456 102303 81490
rect 102605 81456 102639 81490
rect 102941 81456 102975 81490
rect 103277 81456 103311 81490
rect 103613 81456 103647 81490
rect 103949 81456 103983 81490
rect 104285 81456 104319 81490
rect 104621 81456 104655 81490
rect 104957 81456 104991 81490
rect 105293 81456 105327 81490
rect 105629 81456 105663 81490
rect 105965 81456 105999 81490
rect 106301 81456 106335 81490
rect 106637 81456 106671 81490
rect 106973 81456 107007 81490
rect 107309 81456 107343 81490
rect 107645 81456 107679 81490
rect 107981 81456 108015 81490
rect 108317 81456 108351 81490
rect 108653 81456 108687 81490
rect 108989 81456 109023 81490
rect 109325 81456 109359 81490
rect 109661 81456 109695 81490
rect 109997 81456 110031 81490
rect 110333 81456 110367 81490
rect 110669 81456 110703 81490
rect 111005 81456 111039 81490
rect 111341 81456 111375 81490
rect 111677 81456 111711 81490
rect 112013 81456 112047 81490
rect 112349 81456 112383 81490
rect 112685 81456 112719 81490
rect 113021 81456 113055 81490
rect 113357 81456 113391 81490
rect 113693 81456 113727 81490
rect 114029 81456 114063 81490
rect 114365 81456 114399 81490
rect 114701 81456 114735 81490
rect 115037 81456 115071 81490
rect 115373 81456 115407 81490
rect 115709 81456 115743 81490
rect 116045 81456 116079 81490
rect 116381 81456 116415 81490
rect 116717 81456 116751 81490
rect 117053 81456 117087 81490
rect 117389 81456 117423 81490
rect 117725 81456 117759 81490
rect 118061 81456 118095 81490
rect 118397 81456 118431 81490
rect 118733 81456 118767 81490
rect 119069 81456 119103 81490
rect 119405 81456 119439 81490
rect 119741 81456 119775 81490
rect 120077 81456 120111 81490
rect 120413 81456 120447 81490
rect 120749 81456 120783 81490
rect 121085 81456 121119 81490
rect 121421 81456 121455 81490
rect 121757 81456 121791 81490
rect 122093 81456 122127 81490
rect 122429 81456 122463 81490
rect 122765 81456 122799 81490
rect 123101 81456 123135 81490
rect 123437 81456 123471 81490
rect 123773 81456 123807 81490
rect 124109 81456 124143 81490
rect 124445 81456 124479 81490
rect 124781 81456 124815 81490
rect 125117 81456 125151 81490
rect 125453 81456 125487 81490
rect 125789 81456 125823 81490
rect 126125 81456 126159 81490
rect 126461 81456 126495 81490
rect 126797 81456 126831 81490
rect 127133 81456 127167 81490
rect 127469 81456 127503 81490
rect 127805 81456 127839 81490
rect 128141 81456 128175 81490
rect 128477 81456 128511 81490
rect 128813 81456 128847 81490
rect 129149 81456 129183 81490
rect 129485 81456 129519 81490
rect 129821 81456 129855 81490
rect 130157 81456 130191 81490
rect 130493 81456 130527 81490
rect 130829 81456 130863 81490
rect 131165 81456 131199 81490
rect 131501 81456 131535 81490
rect 131837 81456 131871 81490
rect 132173 81456 132207 81490
rect 132509 81456 132543 81490
rect 132845 81456 132879 81490
rect 133181 81456 133215 81490
rect 133517 81456 133551 81490
rect 133853 81456 133887 81490
rect 134189 81456 134223 81490
rect 1805 81003 1839 81037
rect 134855 81003 134889 81037
rect 1805 80667 1839 80701
rect 134855 80667 134889 80701
rect 1805 80331 1839 80365
rect 134855 80331 134889 80365
rect 1805 79995 1839 80029
rect 134855 79995 134889 80029
rect 1805 79659 1839 79693
rect 134855 79659 134889 79693
rect 1805 79323 1839 79357
rect 134855 79323 134889 79357
rect 1805 78987 1839 79021
rect 134855 78987 134889 79021
rect 1805 78651 1839 78685
rect 134855 78651 134889 78685
rect 1805 78315 1839 78349
rect 134855 78315 134889 78349
rect 1805 77979 1839 78013
rect 134855 77979 134889 78013
rect 1805 77643 1839 77677
rect 134855 77643 134889 77677
rect 1805 77307 1839 77341
rect 134855 77307 134889 77341
rect 1805 76971 1839 77005
rect 134855 76971 134889 77005
rect 1805 76635 1839 76669
rect 134855 76635 134889 76669
rect 1805 76299 1839 76333
rect 134855 76299 134889 76333
rect 1805 75963 1839 75997
rect 134855 75963 134889 75997
rect 1805 75627 1839 75661
rect 134855 75627 134889 75661
rect 1805 75291 1839 75325
rect 134855 75291 134889 75325
rect 1805 74955 1839 74989
rect 134855 74955 134889 74989
rect 1805 74619 1839 74653
rect 134855 74619 134889 74653
rect 1805 74283 1839 74317
rect 134855 74283 134889 74317
rect 1805 73947 1839 73981
rect 134855 73947 134889 73981
rect 1805 73611 1839 73645
rect 134855 73611 134889 73645
rect 1805 73275 1839 73309
rect 134855 73275 134889 73309
rect 1805 72939 1839 72973
rect 134855 72939 134889 72973
rect 1805 72603 1839 72637
rect 134855 72603 134889 72637
rect 1805 72267 1839 72301
rect 134855 72267 134889 72301
rect 1805 71931 1839 71965
rect 134855 71931 134889 71965
rect 1805 71595 1839 71629
rect 134855 71595 134889 71629
rect 1805 71259 1839 71293
rect 134855 71259 134889 71293
rect 1805 70923 1839 70957
rect 134855 70923 134889 70957
rect 1805 70587 1839 70621
rect 134855 70587 134889 70621
rect 1805 70251 1839 70285
rect 134855 70251 134889 70285
rect 1805 69915 1839 69949
rect 134855 69915 134889 69949
rect 1805 69579 1839 69613
rect 134855 69579 134889 69613
rect 1805 69243 1839 69277
rect 134855 69243 134889 69277
rect 1805 68907 1839 68941
rect 134855 68907 134889 68941
rect 1805 68571 1839 68605
rect 134855 68571 134889 68605
rect 1805 68235 1839 68269
rect 134855 68235 134889 68269
rect 1805 67899 1839 67933
rect 134855 67899 134889 67933
rect 1805 67563 1839 67597
rect 134855 67563 134889 67597
rect 1805 67227 1839 67261
rect 134855 67227 134889 67261
rect 1805 66891 1839 66925
rect 134855 66891 134889 66925
rect 1805 66555 1839 66589
rect 134855 66555 134889 66589
rect 1805 66219 1839 66253
rect 134855 66219 134889 66253
rect 1805 65883 1839 65917
rect 134855 65883 134889 65917
rect 1805 65547 1839 65581
rect 134855 65547 134889 65581
rect 1805 65211 1839 65245
rect 134855 65211 134889 65245
rect 1805 64875 1839 64909
rect 134855 64875 134889 64909
rect 1805 64539 1839 64573
rect 134855 64539 134889 64573
rect 1805 64203 1839 64237
rect 134855 64203 134889 64237
rect 1805 63867 1839 63901
rect 134855 63867 134889 63901
rect 1805 63531 1839 63565
rect 134855 63531 134889 63565
rect 1805 63195 1839 63229
rect 134855 63195 134889 63229
rect 1805 62859 1839 62893
rect 134855 62859 134889 62893
rect 1805 62523 1839 62557
rect 134855 62523 134889 62557
rect 1805 62187 1839 62221
rect 134855 62187 134889 62221
rect 1805 61851 1839 61885
rect 134855 61851 134889 61885
rect 1805 61515 1839 61549
rect 134855 61515 134889 61549
rect 1805 61179 1839 61213
rect 134855 61179 134889 61213
rect 1805 60843 1839 60877
rect 134855 60843 134889 60877
rect 1805 60507 1839 60541
rect 134855 60507 134889 60541
rect 1805 60171 1839 60205
rect 134855 60171 134889 60205
rect 1805 59835 1839 59869
rect 134855 59835 134889 59869
rect 1805 59499 1839 59533
rect 134855 59499 134889 59533
rect 1805 59163 1839 59197
rect 134855 59163 134889 59197
rect 1805 58827 1839 58861
rect 134855 58827 134889 58861
rect 1805 58491 1839 58525
rect 134855 58491 134889 58525
rect 1805 58155 1839 58189
rect 134855 58155 134889 58189
rect 1805 57819 1839 57853
rect 134855 57819 134889 57853
rect 1805 57483 1839 57517
rect 134855 57483 134889 57517
rect 1805 57147 1839 57181
rect 134855 57147 134889 57181
rect 1805 56811 1839 56845
rect 134855 56811 134889 56845
rect 1805 56475 1839 56509
rect 134855 56475 134889 56509
rect 1805 56139 1839 56173
rect 134855 56139 134889 56173
rect 1805 55803 1839 55837
rect 134855 55803 134889 55837
rect 1805 55467 1839 55501
rect 134855 55467 134889 55501
rect 1805 55131 1839 55165
rect 134855 55131 134889 55165
rect 1805 54795 1839 54829
rect 134855 54795 134889 54829
rect 1805 54459 1839 54493
rect 134855 54459 134889 54493
rect 1805 54123 1839 54157
rect 134855 54123 134889 54157
rect 1805 53787 1839 53821
rect 134855 53787 134889 53821
rect 1805 53451 1839 53485
rect 134855 53451 134889 53485
rect 1805 53115 1839 53149
rect 134855 53115 134889 53149
rect 1805 52779 1839 52813
rect 134855 52779 134889 52813
rect 1805 52443 1839 52477
rect 134855 52443 134889 52477
rect 1805 52107 1839 52141
rect 134855 52107 134889 52141
rect 1805 51771 1839 51805
rect 134855 51771 134889 51805
rect 1805 51435 1839 51469
rect 134855 51435 134889 51469
rect 1805 51099 1839 51133
rect 134855 51099 134889 51133
rect 1805 50763 1839 50797
rect 134855 50763 134889 50797
rect 1805 50427 1839 50461
rect 134855 50427 134889 50461
rect 1805 50091 1839 50125
rect 134855 50091 134889 50125
rect 1805 49755 1839 49789
rect 134855 49755 134889 49789
rect 1805 49419 1839 49453
rect 134855 49419 134889 49453
rect 1805 49083 1839 49117
rect 134855 49083 134889 49117
rect 1805 48747 1839 48781
rect 134855 48747 134889 48781
rect 1805 48411 1839 48445
rect 134855 48411 134889 48445
rect 1805 48075 1839 48109
rect 134855 48075 134889 48109
rect 1805 47739 1839 47773
rect 134855 47739 134889 47773
rect 1805 47403 1839 47437
rect 134855 47403 134889 47437
rect 1805 47067 1839 47101
rect 134855 47067 134889 47101
rect 1805 46731 1839 46765
rect 134855 46731 134889 46765
rect 1805 46395 1839 46429
rect 134855 46395 134889 46429
rect 1805 46059 1839 46093
rect 134855 46059 134889 46093
rect 1805 45723 1839 45757
rect 134855 45723 134889 45757
rect 1805 45387 1839 45421
rect 134855 45387 134889 45421
rect 1805 45051 1839 45085
rect 134855 45051 134889 45085
rect 1805 44715 1839 44749
rect 134855 44715 134889 44749
rect 1805 44379 1839 44413
rect 134855 44379 134889 44413
rect 1805 44043 1839 44077
rect 134855 44043 134889 44077
rect 1805 43707 1839 43741
rect 134855 43707 134889 43741
rect 1805 43371 1839 43405
rect 134855 43371 134889 43405
rect 1805 43035 1839 43069
rect 134855 43035 134889 43069
rect 1805 42699 1839 42733
rect 134855 42699 134889 42733
rect 1805 42363 1839 42397
rect 134855 42363 134889 42397
rect 1805 42027 1839 42061
rect 134855 42027 134889 42061
rect 1805 41691 1839 41725
rect 134855 41691 134889 41725
rect 1805 41355 1839 41389
rect 134855 41355 134889 41389
rect 1805 41019 1839 41053
rect 134855 41019 134889 41053
rect 1805 40683 1839 40717
rect 134855 40683 134889 40717
rect 1805 40347 1839 40381
rect 134855 40347 134889 40381
rect 1805 40011 1839 40045
rect 134855 40011 134889 40045
rect 1805 39675 1839 39709
rect 134855 39675 134889 39709
rect 1805 39339 1839 39373
rect 134855 39339 134889 39373
rect 1805 39003 1839 39037
rect 134855 39003 134889 39037
rect 1805 38667 1839 38701
rect 134855 38667 134889 38701
rect 1805 38331 1839 38365
rect 134855 38331 134889 38365
rect 1805 37995 1839 38029
rect 134855 37995 134889 38029
rect 1805 37659 1839 37693
rect 134855 37659 134889 37693
rect 1805 37323 1839 37357
rect 134855 37323 134889 37357
rect 1805 36987 1839 37021
rect 134855 36987 134889 37021
rect 1805 36651 1839 36685
rect 134855 36651 134889 36685
rect 1805 36315 1839 36349
rect 134855 36315 134889 36349
rect 1805 35979 1839 36013
rect 134855 35979 134889 36013
rect 1805 35643 1839 35677
rect 134855 35643 134889 35677
rect 1805 35307 1839 35341
rect 134855 35307 134889 35341
rect 1805 34971 1839 35005
rect 134855 34971 134889 35005
rect 1805 34635 1839 34669
rect 134855 34635 134889 34669
rect 1805 34299 1839 34333
rect 134855 34299 134889 34333
rect 1805 33963 1839 33997
rect 134855 33963 134889 33997
rect 1805 33627 1839 33661
rect 134855 33627 134889 33661
rect 1805 33291 1839 33325
rect 134855 33291 134889 33325
rect 1805 32955 1839 32989
rect 134855 32955 134889 32989
rect 1805 32619 1839 32653
rect 134855 32619 134889 32653
rect 1805 32283 1839 32317
rect 134855 32283 134889 32317
rect 1805 31947 1839 31981
rect 134855 31947 134889 31981
rect 1805 31611 1839 31645
rect 134855 31611 134889 31645
rect 1805 31275 1839 31309
rect 134855 31275 134889 31309
rect 1805 30939 1839 30973
rect 134855 30939 134889 30973
rect 1805 30603 1839 30637
rect 134855 30603 134889 30637
rect 1805 30267 1839 30301
rect 134855 30267 134889 30301
rect 1805 29931 1839 29965
rect 134855 29931 134889 29965
rect 1805 29595 1839 29629
rect 134855 29595 134889 29629
rect 1805 29259 1839 29293
rect 134855 29259 134889 29293
rect 1805 28923 1839 28957
rect 134855 28923 134889 28957
rect 1805 28587 1839 28621
rect 134855 28587 134889 28621
rect 1805 28251 1839 28285
rect 134855 28251 134889 28285
rect 1805 27915 1839 27949
rect 134855 27915 134889 27949
rect 1805 27579 1839 27613
rect 134855 27579 134889 27613
rect 1805 27243 1839 27277
rect 134855 27243 134889 27277
rect 1805 26907 1839 26941
rect 134855 26907 134889 26941
rect 1805 26571 1839 26605
rect 134855 26571 134889 26605
rect 1805 26235 1839 26269
rect 134855 26235 134889 26269
rect 1805 25899 1839 25933
rect 134855 25899 134889 25933
rect 1805 25563 1839 25597
rect 134855 25563 134889 25597
rect 1805 25227 1839 25261
rect 134855 25227 134889 25261
rect 1805 24891 1839 24925
rect 134855 24891 134889 24925
rect 1805 24555 1839 24589
rect 134855 24555 134889 24589
rect 1805 24219 1839 24253
rect 134855 24219 134889 24253
rect 1805 23883 1839 23917
rect 134855 23883 134889 23917
rect 1805 23547 1839 23581
rect 134855 23547 134889 23581
rect 1805 23211 1839 23245
rect 134855 23211 134889 23245
rect 1805 22875 1839 22909
rect 134855 22875 134889 22909
rect 1805 22539 1839 22573
rect 134855 22539 134889 22573
rect 1805 22203 1839 22237
rect 134855 22203 134889 22237
rect 1805 21867 1839 21901
rect 134855 21867 134889 21901
rect 1805 21531 1839 21565
rect 134855 21531 134889 21565
rect 1805 21195 1839 21229
rect 134855 21195 134889 21229
rect 1805 20859 1839 20893
rect 134855 20859 134889 20893
rect 1805 20523 1839 20557
rect 134855 20523 134889 20557
rect 1805 20187 1839 20221
rect 134855 20187 134889 20221
rect 1805 19851 1839 19885
rect 134855 19851 134889 19885
rect 1805 19515 1839 19549
rect 134855 19515 134889 19549
rect 1805 19179 1839 19213
rect 134855 19179 134889 19213
rect 1805 18843 1839 18877
rect 134855 18843 134889 18877
rect 1805 18507 1839 18541
rect 134855 18507 134889 18541
rect 1805 18171 1839 18205
rect 134855 18171 134889 18205
rect 1805 17835 1839 17869
rect 134855 17835 134889 17869
rect 1805 17499 1839 17533
rect 134855 17499 134889 17533
rect 1805 17163 1839 17197
rect 134855 17163 134889 17197
rect 1805 16827 1839 16861
rect 134855 16827 134889 16861
rect 1805 16491 1839 16525
rect 134855 16491 134889 16525
rect 1805 16155 1839 16189
rect 134855 16155 134889 16189
rect 1805 15819 1839 15853
rect 134855 15819 134889 15853
rect 1805 15483 1839 15517
rect 134855 15483 134889 15517
rect 1805 15147 1839 15181
rect 134855 15147 134889 15181
rect 1805 14811 1839 14845
rect 134855 14811 134889 14845
rect 1805 14475 1839 14509
rect 134855 14475 134889 14509
rect 1805 14139 1839 14173
rect 134855 14139 134889 14173
rect 1805 13803 1839 13837
rect 134855 13803 134889 13837
rect 1805 13467 1839 13501
rect 134855 13467 134889 13501
rect 1805 13131 1839 13165
rect 134855 13131 134889 13165
rect 1805 12795 1839 12829
rect 134855 12795 134889 12829
rect 1805 12459 1839 12493
rect 134855 12459 134889 12493
rect 1805 12123 1839 12157
rect 134855 12123 134889 12157
rect 1805 11787 1839 11821
rect 134855 11787 134889 11821
rect 1805 11451 1839 11485
rect 134855 11451 134889 11485
rect 1805 11115 1839 11149
rect 134855 11115 134889 11149
rect 1805 10779 1839 10813
rect 134855 10779 134889 10813
rect 1805 10443 1839 10477
rect 134855 10443 134889 10477
rect 1805 10107 1839 10141
rect 134855 10107 134889 10141
rect 1805 9771 1839 9805
rect 134855 9771 134889 9805
rect 1805 9435 1839 9469
rect 134855 9435 134889 9469
rect 1805 9099 1839 9133
rect 134855 9099 134889 9133
rect 1805 8763 1839 8797
rect 134855 8763 134889 8797
rect 1805 8427 1839 8461
rect 134855 8427 134889 8461
rect 1805 8091 1839 8125
rect 134855 8091 134889 8125
rect 1805 7755 1839 7789
rect 134855 7755 134889 7789
rect 1805 7419 1839 7453
rect 134855 7419 134889 7453
rect 1805 7083 1839 7117
rect 134855 7083 134889 7117
rect 1805 6747 1839 6781
rect 134855 6747 134889 6781
rect 1805 6411 1839 6445
rect 134855 6411 134889 6445
rect 1805 6075 1839 6109
rect 134855 6075 134889 6109
rect 1805 5739 1839 5773
rect 134855 5739 134889 5773
rect 1805 5403 1839 5437
rect 134855 5403 134889 5437
rect 1805 5067 1839 5101
rect 134855 5067 134889 5101
rect 1805 4731 1839 4765
rect 134855 4731 134889 4765
rect 1805 4395 1839 4429
rect 134855 4395 134889 4429
rect 1805 4059 1839 4093
rect 134855 4059 134889 4093
rect 1805 3723 1839 3757
rect 134855 3723 134889 3757
rect 1805 3387 1839 3421
rect 134855 3387 134889 3421
rect 1805 3051 1839 3085
rect 134855 3051 134889 3085
rect 1805 2715 1839 2749
rect 134855 2715 134889 2749
rect 1805 2379 1839 2413
rect 134855 2379 134889 2413
rect 1805 2043 1839 2077
rect 134855 2043 134889 2077
rect 2141 1707 2175 1741
rect 2477 1707 2511 1741
rect 2813 1707 2847 1741
rect 3149 1707 3183 1741
rect 3485 1707 3519 1741
rect 3821 1707 3855 1741
rect 4157 1707 4191 1741
rect 4493 1707 4527 1741
rect 4829 1707 4863 1741
rect 5165 1707 5199 1741
rect 5501 1707 5535 1741
rect 5837 1707 5871 1741
rect 6173 1707 6207 1741
rect 6509 1707 6543 1741
rect 6845 1707 6879 1741
rect 7181 1707 7215 1741
rect 7517 1707 7551 1741
rect 7853 1707 7887 1741
rect 8189 1707 8223 1741
rect 8525 1707 8559 1741
rect 8861 1707 8895 1741
rect 9197 1707 9231 1741
rect 9533 1707 9567 1741
rect 9869 1707 9903 1741
rect 10205 1707 10239 1741
rect 10541 1707 10575 1741
rect 10877 1707 10911 1741
rect 11213 1707 11247 1741
rect 11549 1707 11583 1741
rect 11885 1707 11919 1741
rect 12221 1707 12255 1741
rect 12557 1707 12591 1741
rect 12893 1707 12927 1741
rect 13229 1707 13263 1741
rect 13565 1707 13599 1741
rect 13901 1707 13935 1741
rect 14237 1707 14271 1741
rect 14573 1707 14607 1741
rect 14909 1707 14943 1741
rect 15245 1707 15279 1741
rect 15581 1707 15615 1741
rect 15917 1707 15951 1741
rect 16253 1707 16287 1741
rect 16589 1707 16623 1741
rect 16925 1707 16959 1741
rect 17261 1707 17295 1741
rect 17597 1707 17631 1741
rect 17933 1707 17967 1741
rect 18269 1707 18303 1741
rect 18605 1707 18639 1741
rect 18941 1707 18975 1741
rect 19277 1707 19311 1741
rect 19613 1707 19647 1741
rect 19949 1707 19983 1741
rect 20285 1707 20319 1741
rect 20621 1707 20655 1741
rect 20957 1707 20991 1741
rect 21293 1707 21327 1741
rect 21629 1707 21663 1741
rect 21965 1707 21999 1741
rect 22301 1707 22335 1741
rect 22637 1707 22671 1741
rect 22973 1707 23007 1741
rect 23309 1707 23343 1741
rect 23645 1707 23679 1741
rect 23981 1707 24015 1741
rect 24317 1707 24351 1741
rect 24653 1707 24687 1741
rect 24989 1707 25023 1741
rect 25325 1707 25359 1741
rect 25661 1707 25695 1741
rect 25997 1707 26031 1741
rect 26333 1707 26367 1741
rect 26669 1707 26703 1741
rect 27005 1707 27039 1741
rect 27341 1707 27375 1741
rect 27677 1707 27711 1741
rect 28013 1707 28047 1741
rect 28349 1707 28383 1741
rect 28685 1707 28719 1741
rect 29021 1707 29055 1741
rect 29357 1707 29391 1741
rect 29693 1707 29727 1741
rect 30029 1707 30063 1741
rect 30365 1707 30399 1741
rect 30701 1707 30735 1741
rect 31037 1707 31071 1741
rect 31373 1707 31407 1741
rect 31709 1707 31743 1741
rect 32045 1707 32079 1741
rect 32381 1707 32415 1741
rect 32717 1707 32751 1741
rect 33053 1707 33087 1741
rect 33389 1707 33423 1741
rect 33725 1707 33759 1741
rect 34061 1707 34095 1741
rect 34397 1707 34431 1741
rect 34733 1707 34767 1741
rect 35069 1707 35103 1741
rect 35405 1707 35439 1741
rect 35741 1707 35775 1741
rect 36077 1707 36111 1741
rect 36413 1707 36447 1741
rect 36749 1707 36783 1741
rect 37085 1707 37119 1741
rect 37421 1707 37455 1741
rect 37757 1707 37791 1741
rect 38093 1707 38127 1741
rect 38429 1707 38463 1741
rect 38765 1707 38799 1741
rect 39101 1707 39135 1741
rect 39437 1707 39471 1741
rect 39773 1707 39807 1741
rect 40109 1707 40143 1741
rect 40445 1707 40479 1741
rect 40781 1707 40815 1741
rect 41117 1707 41151 1741
rect 41453 1707 41487 1741
rect 41789 1707 41823 1741
rect 42125 1707 42159 1741
rect 42461 1707 42495 1741
rect 42797 1707 42831 1741
rect 43133 1707 43167 1741
rect 43469 1707 43503 1741
rect 43805 1707 43839 1741
rect 44141 1707 44175 1741
rect 44477 1707 44511 1741
rect 44813 1707 44847 1741
rect 45149 1707 45183 1741
rect 45485 1707 45519 1741
rect 45821 1707 45855 1741
rect 46157 1707 46191 1741
rect 46493 1707 46527 1741
rect 46829 1707 46863 1741
rect 47165 1707 47199 1741
rect 47501 1707 47535 1741
rect 47837 1707 47871 1741
rect 48173 1707 48207 1741
rect 48509 1707 48543 1741
rect 48845 1707 48879 1741
rect 49181 1707 49215 1741
rect 49517 1707 49551 1741
rect 49853 1707 49887 1741
rect 50189 1707 50223 1741
rect 50525 1707 50559 1741
rect 50861 1707 50895 1741
rect 51197 1707 51231 1741
rect 51533 1707 51567 1741
rect 51869 1707 51903 1741
rect 52205 1707 52239 1741
rect 52541 1707 52575 1741
rect 52877 1707 52911 1741
rect 53213 1707 53247 1741
rect 53549 1707 53583 1741
rect 53885 1707 53919 1741
rect 54221 1707 54255 1741
rect 54557 1707 54591 1741
rect 54893 1707 54927 1741
rect 55229 1707 55263 1741
rect 55565 1707 55599 1741
rect 55901 1707 55935 1741
rect 56237 1707 56271 1741
rect 56573 1707 56607 1741
rect 56909 1707 56943 1741
rect 57245 1707 57279 1741
rect 57581 1707 57615 1741
rect 57917 1707 57951 1741
rect 58253 1707 58287 1741
rect 58589 1707 58623 1741
rect 58925 1707 58959 1741
rect 59261 1707 59295 1741
rect 59597 1707 59631 1741
rect 59933 1707 59967 1741
rect 60269 1707 60303 1741
rect 60605 1707 60639 1741
rect 60941 1707 60975 1741
rect 61277 1707 61311 1741
rect 61613 1707 61647 1741
rect 61949 1707 61983 1741
rect 62285 1707 62319 1741
rect 62621 1707 62655 1741
rect 62957 1707 62991 1741
rect 63293 1707 63327 1741
rect 63629 1707 63663 1741
rect 63965 1707 63999 1741
rect 64301 1707 64335 1741
rect 64637 1707 64671 1741
rect 64973 1707 65007 1741
rect 65309 1707 65343 1741
rect 65645 1707 65679 1741
rect 65981 1707 66015 1741
rect 66317 1707 66351 1741
rect 66653 1707 66687 1741
rect 66989 1707 67023 1741
rect 67325 1707 67359 1741
rect 67661 1707 67695 1741
rect 67997 1707 68031 1741
rect 68333 1707 68367 1741
rect 68669 1707 68703 1741
rect 69005 1707 69039 1741
rect 69341 1707 69375 1741
rect 69677 1707 69711 1741
rect 70013 1707 70047 1741
rect 70349 1707 70383 1741
rect 70685 1707 70719 1741
rect 71021 1707 71055 1741
rect 71357 1707 71391 1741
rect 71693 1707 71727 1741
rect 72029 1707 72063 1741
rect 72365 1707 72399 1741
rect 72701 1707 72735 1741
rect 73037 1707 73071 1741
rect 73373 1707 73407 1741
rect 73709 1707 73743 1741
rect 74045 1707 74079 1741
rect 74381 1707 74415 1741
rect 74717 1707 74751 1741
rect 75053 1707 75087 1741
rect 75389 1707 75423 1741
rect 75725 1707 75759 1741
rect 76061 1707 76095 1741
rect 76397 1707 76431 1741
rect 76733 1707 76767 1741
rect 77069 1707 77103 1741
rect 77405 1707 77439 1741
rect 77741 1707 77775 1741
rect 78077 1707 78111 1741
rect 78413 1707 78447 1741
rect 78749 1707 78783 1741
rect 79085 1707 79119 1741
rect 79421 1707 79455 1741
rect 79757 1707 79791 1741
rect 80093 1707 80127 1741
rect 80429 1707 80463 1741
rect 80765 1707 80799 1741
rect 81101 1707 81135 1741
rect 81437 1707 81471 1741
rect 81773 1707 81807 1741
rect 82109 1707 82143 1741
rect 82445 1707 82479 1741
rect 82781 1707 82815 1741
rect 83117 1707 83151 1741
rect 83453 1707 83487 1741
rect 83789 1707 83823 1741
rect 84125 1707 84159 1741
rect 84461 1707 84495 1741
rect 84797 1707 84831 1741
rect 85133 1707 85167 1741
rect 85469 1707 85503 1741
rect 85805 1707 85839 1741
rect 86141 1707 86175 1741
rect 86477 1707 86511 1741
rect 86813 1707 86847 1741
rect 87149 1707 87183 1741
rect 87485 1707 87519 1741
rect 87821 1707 87855 1741
rect 88157 1707 88191 1741
rect 88493 1707 88527 1741
rect 88829 1707 88863 1741
rect 89165 1707 89199 1741
rect 89501 1707 89535 1741
rect 89837 1707 89871 1741
rect 90173 1707 90207 1741
rect 90509 1707 90543 1741
rect 90845 1707 90879 1741
rect 91181 1707 91215 1741
rect 91517 1707 91551 1741
rect 91853 1707 91887 1741
rect 92189 1707 92223 1741
rect 92525 1707 92559 1741
rect 92861 1707 92895 1741
rect 93197 1707 93231 1741
rect 93533 1707 93567 1741
rect 93869 1707 93903 1741
rect 94205 1707 94239 1741
rect 94541 1707 94575 1741
rect 94877 1707 94911 1741
rect 95213 1707 95247 1741
rect 95549 1707 95583 1741
rect 95885 1707 95919 1741
rect 96221 1707 96255 1741
rect 96557 1707 96591 1741
rect 96893 1707 96927 1741
rect 97229 1707 97263 1741
rect 97565 1707 97599 1741
rect 97901 1707 97935 1741
rect 98237 1707 98271 1741
rect 98573 1707 98607 1741
rect 98909 1707 98943 1741
rect 99245 1707 99279 1741
rect 99581 1707 99615 1741
rect 99917 1707 99951 1741
rect 100253 1707 100287 1741
rect 100589 1707 100623 1741
rect 100925 1707 100959 1741
rect 101261 1707 101295 1741
rect 101597 1707 101631 1741
rect 101933 1707 101967 1741
rect 102269 1707 102303 1741
rect 102605 1707 102639 1741
rect 102941 1707 102975 1741
rect 103277 1707 103311 1741
rect 103613 1707 103647 1741
rect 103949 1707 103983 1741
rect 104285 1707 104319 1741
rect 104621 1707 104655 1741
rect 104957 1707 104991 1741
rect 105293 1707 105327 1741
rect 105629 1707 105663 1741
rect 105965 1707 105999 1741
rect 106301 1707 106335 1741
rect 106637 1707 106671 1741
rect 106973 1707 107007 1741
rect 107309 1707 107343 1741
rect 107645 1707 107679 1741
rect 107981 1707 108015 1741
rect 108317 1707 108351 1741
rect 108653 1707 108687 1741
rect 108989 1707 109023 1741
rect 109325 1707 109359 1741
rect 109661 1707 109695 1741
rect 109997 1707 110031 1741
rect 110333 1707 110367 1741
rect 110669 1707 110703 1741
rect 111005 1707 111039 1741
rect 111341 1707 111375 1741
rect 111677 1707 111711 1741
rect 112013 1707 112047 1741
rect 112349 1707 112383 1741
rect 112685 1707 112719 1741
rect 113021 1707 113055 1741
rect 113357 1707 113391 1741
rect 113693 1707 113727 1741
rect 114029 1707 114063 1741
rect 114365 1707 114399 1741
rect 114701 1707 114735 1741
rect 115037 1707 115071 1741
rect 115373 1707 115407 1741
rect 115709 1707 115743 1741
rect 116045 1707 116079 1741
rect 116381 1707 116415 1741
rect 116717 1707 116751 1741
rect 117053 1707 117087 1741
rect 117389 1707 117423 1741
rect 117725 1707 117759 1741
rect 118061 1707 118095 1741
rect 118397 1707 118431 1741
rect 118733 1707 118767 1741
rect 119069 1707 119103 1741
rect 119405 1707 119439 1741
rect 119741 1707 119775 1741
rect 120077 1707 120111 1741
rect 120413 1707 120447 1741
rect 120749 1707 120783 1741
rect 121085 1707 121119 1741
rect 121421 1707 121455 1741
rect 121757 1707 121791 1741
rect 122093 1707 122127 1741
rect 122429 1707 122463 1741
rect 122765 1707 122799 1741
rect 123101 1707 123135 1741
rect 123437 1707 123471 1741
rect 123773 1707 123807 1741
rect 124109 1707 124143 1741
rect 124445 1707 124479 1741
rect 124781 1707 124815 1741
rect 125117 1707 125151 1741
rect 125453 1707 125487 1741
rect 125789 1707 125823 1741
rect 126125 1707 126159 1741
rect 126461 1707 126495 1741
rect 126797 1707 126831 1741
rect 127133 1707 127167 1741
rect 127469 1707 127503 1741
rect 127805 1707 127839 1741
rect 128141 1707 128175 1741
rect 128477 1707 128511 1741
rect 128813 1707 128847 1741
rect 129149 1707 129183 1741
rect 129485 1707 129519 1741
rect 129821 1707 129855 1741
rect 130157 1707 130191 1741
rect 130493 1707 130527 1741
rect 130829 1707 130863 1741
rect 131165 1707 131199 1741
rect 131501 1707 131535 1741
rect 131837 1707 131871 1741
rect 132173 1707 132207 1741
rect 132509 1707 132543 1741
rect 132845 1707 132879 1741
rect 133181 1707 133215 1741
rect 133517 1707 133551 1741
rect 133853 1707 133887 1741
rect 134189 1707 134223 1741
<< locali >>
rect 2141 81490 2175 81506
rect 2141 81440 2175 81456
rect 2477 81490 2511 81506
rect 2477 81440 2511 81456
rect 2813 81490 2847 81506
rect 2813 81440 2847 81456
rect 3149 81490 3183 81506
rect 3149 81440 3183 81456
rect 3485 81490 3519 81506
rect 3485 81440 3519 81456
rect 3821 81490 3855 81506
rect 3821 81440 3855 81456
rect 4157 81490 4191 81506
rect 4157 81440 4191 81456
rect 4493 81490 4527 81506
rect 4493 81440 4527 81456
rect 4829 81490 4863 81506
rect 4829 81440 4863 81456
rect 5165 81490 5199 81506
rect 5165 81440 5199 81456
rect 5501 81490 5535 81506
rect 5501 81440 5535 81456
rect 5837 81490 5871 81506
rect 5837 81440 5871 81456
rect 6173 81490 6207 81506
rect 6173 81440 6207 81456
rect 6509 81490 6543 81506
rect 6509 81440 6543 81456
rect 6845 81490 6879 81506
rect 6845 81440 6879 81456
rect 7181 81490 7215 81506
rect 7181 81440 7215 81456
rect 7517 81490 7551 81506
rect 7517 81440 7551 81456
rect 7853 81490 7887 81506
rect 7853 81440 7887 81456
rect 8189 81490 8223 81506
rect 8189 81440 8223 81456
rect 8525 81490 8559 81506
rect 8525 81440 8559 81456
rect 8861 81490 8895 81506
rect 8861 81440 8895 81456
rect 9197 81490 9231 81506
rect 9197 81440 9231 81456
rect 9533 81490 9567 81506
rect 9533 81440 9567 81456
rect 9869 81490 9903 81506
rect 9869 81440 9903 81456
rect 10205 81490 10239 81506
rect 10205 81440 10239 81456
rect 10541 81490 10575 81506
rect 10541 81440 10575 81456
rect 10877 81490 10911 81506
rect 10877 81440 10911 81456
rect 11213 81490 11247 81506
rect 11213 81440 11247 81456
rect 11549 81490 11583 81506
rect 11549 81440 11583 81456
rect 11885 81490 11919 81506
rect 11885 81440 11919 81456
rect 12221 81490 12255 81506
rect 12221 81440 12255 81456
rect 12557 81490 12591 81506
rect 12557 81440 12591 81456
rect 12893 81490 12927 81506
rect 12893 81440 12927 81456
rect 13229 81490 13263 81506
rect 13229 81440 13263 81456
rect 13565 81490 13599 81506
rect 13565 81440 13599 81456
rect 13901 81490 13935 81506
rect 13901 81440 13935 81456
rect 14237 81490 14271 81506
rect 14237 81440 14271 81456
rect 14573 81490 14607 81506
rect 14573 81440 14607 81456
rect 14909 81490 14943 81506
rect 14909 81440 14943 81456
rect 15245 81490 15279 81506
rect 15245 81440 15279 81456
rect 15581 81490 15615 81506
rect 15581 81440 15615 81456
rect 15917 81490 15951 81506
rect 15917 81440 15951 81456
rect 16253 81490 16287 81506
rect 16253 81440 16287 81456
rect 16589 81490 16623 81506
rect 16589 81440 16623 81456
rect 16925 81490 16959 81506
rect 16925 81440 16959 81456
rect 17261 81490 17295 81506
rect 17261 81440 17295 81456
rect 17597 81490 17631 81506
rect 17597 81440 17631 81456
rect 17933 81490 17967 81506
rect 17933 81440 17967 81456
rect 18269 81490 18303 81506
rect 18269 81440 18303 81456
rect 18605 81490 18639 81506
rect 18605 81440 18639 81456
rect 18941 81490 18975 81506
rect 18941 81440 18975 81456
rect 19277 81490 19311 81506
rect 19277 81440 19311 81456
rect 19613 81490 19647 81506
rect 19613 81440 19647 81456
rect 19949 81490 19983 81506
rect 19949 81440 19983 81456
rect 20285 81490 20319 81506
rect 20285 81440 20319 81456
rect 20621 81490 20655 81506
rect 20621 81440 20655 81456
rect 20957 81490 20991 81506
rect 20957 81440 20991 81456
rect 21293 81490 21327 81506
rect 21293 81440 21327 81456
rect 21629 81490 21663 81506
rect 21629 81440 21663 81456
rect 21965 81490 21999 81506
rect 21965 81440 21999 81456
rect 22301 81490 22335 81506
rect 22301 81440 22335 81456
rect 22637 81490 22671 81506
rect 22637 81440 22671 81456
rect 22973 81490 23007 81506
rect 22973 81440 23007 81456
rect 23309 81490 23343 81506
rect 23309 81440 23343 81456
rect 23645 81490 23679 81506
rect 23645 81440 23679 81456
rect 23981 81490 24015 81506
rect 23981 81440 24015 81456
rect 24317 81490 24351 81506
rect 24317 81440 24351 81456
rect 24653 81490 24687 81506
rect 24653 81440 24687 81456
rect 24989 81490 25023 81506
rect 24989 81440 25023 81456
rect 25325 81490 25359 81506
rect 25325 81440 25359 81456
rect 25661 81490 25695 81506
rect 25661 81440 25695 81456
rect 25997 81490 26031 81506
rect 25997 81440 26031 81456
rect 26333 81490 26367 81506
rect 26333 81440 26367 81456
rect 26669 81490 26703 81506
rect 26669 81440 26703 81456
rect 27005 81490 27039 81506
rect 27005 81440 27039 81456
rect 27341 81490 27375 81506
rect 27341 81440 27375 81456
rect 27677 81490 27711 81506
rect 27677 81440 27711 81456
rect 28013 81490 28047 81506
rect 28013 81440 28047 81456
rect 28349 81490 28383 81506
rect 28349 81440 28383 81456
rect 28685 81490 28719 81506
rect 28685 81440 28719 81456
rect 29021 81490 29055 81506
rect 29021 81440 29055 81456
rect 29357 81490 29391 81506
rect 29357 81440 29391 81456
rect 29693 81490 29727 81506
rect 29693 81440 29727 81456
rect 30029 81490 30063 81506
rect 30029 81440 30063 81456
rect 30365 81490 30399 81506
rect 30365 81440 30399 81456
rect 30701 81490 30735 81506
rect 30701 81440 30735 81456
rect 31037 81490 31071 81506
rect 31037 81440 31071 81456
rect 31373 81490 31407 81506
rect 31373 81440 31407 81456
rect 31709 81490 31743 81506
rect 31709 81440 31743 81456
rect 32045 81490 32079 81506
rect 32045 81440 32079 81456
rect 32381 81490 32415 81506
rect 32381 81440 32415 81456
rect 32717 81490 32751 81506
rect 32717 81440 32751 81456
rect 33053 81490 33087 81506
rect 33053 81440 33087 81456
rect 33389 81490 33423 81506
rect 33389 81440 33423 81456
rect 33725 81490 33759 81506
rect 33725 81440 33759 81456
rect 34061 81490 34095 81506
rect 34061 81440 34095 81456
rect 34397 81490 34431 81506
rect 34397 81440 34431 81456
rect 34733 81490 34767 81506
rect 34733 81440 34767 81456
rect 35069 81490 35103 81506
rect 35069 81440 35103 81456
rect 35405 81490 35439 81506
rect 35405 81440 35439 81456
rect 35741 81490 35775 81506
rect 35741 81440 35775 81456
rect 36077 81490 36111 81506
rect 36077 81440 36111 81456
rect 36413 81490 36447 81506
rect 36413 81440 36447 81456
rect 36749 81490 36783 81506
rect 36749 81440 36783 81456
rect 37085 81490 37119 81506
rect 37085 81440 37119 81456
rect 37421 81490 37455 81506
rect 37421 81440 37455 81456
rect 37757 81490 37791 81506
rect 37757 81440 37791 81456
rect 38093 81490 38127 81506
rect 38093 81440 38127 81456
rect 38429 81490 38463 81506
rect 38429 81440 38463 81456
rect 38765 81490 38799 81506
rect 38765 81440 38799 81456
rect 39101 81490 39135 81506
rect 39101 81440 39135 81456
rect 39437 81490 39471 81506
rect 39437 81440 39471 81456
rect 39773 81490 39807 81506
rect 39773 81440 39807 81456
rect 40109 81490 40143 81506
rect 40109 81440 40143 81456
rect 40445 81490 40479 81506
rect 40445 81440 40479 81456
rect 40781 81490 40815 81506
rect 40781 81440 40815 81456
rect 41117 81490 41151 81506
rect 41117 81440 41151 81456
rect 41453 81490 41487 81506
rect 41453 81440 41487 81456
rect 41789 81490 41823 81506
rect 41789 81440 41823 81456
rect 42125 81490 42159 81506
rect 42125 81440 42159 81456
rect 42461 81490 42495 81506
rect 42461 81440 42495 81456
rect 42797 81490 42831 81506
rect 42797 81440 42831 81456
rect 43133 81490 43167 81506
rect 43133 81440 43167 81456
rect 43469 81490 43503 81506
rect 43469 81440 43503 81456
rect 43805 81490 43839 81506
rect 43805 81440 43839 81456
rect 44141 81490 44175 81506
rect 44141 81440 44175 81456
rect 44477 81490 44511 81506
rect 44477 81440 44511 81456
rect 44813 81490 44847 81506
rect 44813 81440 44847 81456
rect 45149 81490 45183 81506
rect 45149 81440 45183 81456
rect 45485 81490 45519 81506
rect 45485 81440 45519 81456
rect 45821 81490 45855 81506
rect 45821 81440 45855 81456
rect 46157 81490 46191 81506
rect 46157 81440 46191 81456
rect 46493 81490 46527 81506
rect 46493 81440 46527 81456
rect 46829 81490 46863 81506
rect 46829 81440 46863 81456
rect 47165 81490 47199 81506
rect 47165 81440 47199 81456
rect 47501 81490 47535 81506
rect 47501 81440 47535 81456
rect 47837 81490 47871 81506
rect 47837 81440 47871 81456
rect 48173 81490 48207 81506
rect 48173 81440 48207 81456
rect 48509 81490 48543 81506
rect 48509 81440 48543 81456
rect 48845 81490 48879 81506
rect 48845 81440 48879 81456
rect 49181 81490 49215 81506
rect 49181 81440 49215 81456
rect 49517 81490 49551 81506
rect 49517 81440 49551 81456
rect 49853 81490 49887 81506
rect 49853 81440 49887 81456
rect 50189 81490 50223 81506
rect 50189 81440 50223 81456
rect 50525 81490 50559 81506
rect 50525 81440 50559 81456
rect 50861 81490 50895 81506
rect 50861 81440 50895 81456
rect 51197 81490 51231 81506
rect 51197 81440 51231 81456
rect 51533 81490 51567 81506
rect 51533 81440 51567 81456
rect 51869 81490 51903 81506
rect 51869 81440 51903 81456
rect 52205 81490 52239 81506
rect 52205 81440 52239 81456
rect 52541 81490 52575 81506
rect 52541 81440 52575 81456
rect 52877 81490 52911 81506
rect 52877 81440 52911 81456
rect 53213 81490 53247 81506
rect 53213 81440 53247 81456
rect 53549 81490 53583 81506
rect 53549 81440 53583 81456
rect 53885 81490 53919 81506
rect 53885 81440 53919 81456
rect 54221 81490 54255 81506
rect 54221 81440 54255 81456
rect 54557 81490 54591 81506
rect 54557 81440 54591 81456
rect 54893 81490 54927 81506
rect 54893 81440 54927 81456
rect 55229 81490 55263 81506
rect 55229 81440 55263 81456
rect 55565 81490 55599 81506
rect 55565 81440 55599 81456
rect 55901 81490 55935 81506
rect 55901 81440 55935 81456
rect 56237 81490 56271 81506
rect 56237 81440 56271 81456
rect 56573 81490 56607 81506
rect 56573 81440 56607 81456
rect 56909 81490 56943 81506
rect 56909 81440 56943 81456
rect 57245 81490 57279 81506
rect 57245 81440 57279 81456
rect 57581 81490 57615 81506
rect 57581 81440 57615 81456
rect 57917 81490 57951 81506
rect 57917 81440 57951 81456
rect 58253 81490 58287 81506
rect 58253 81440 58287 81456
rect 58589 81490 58623 81506
rect 58589 81440 58623 81456
rect 58925 81490 58959 81506
rect 58925 81440 58959 81456
rect 59261 81490 59295 81506
rect 59261 81440 59295 81456
rect 59597 81490 59631 81506
rect 59597 81440 59631 81456
rect 59933 81490 59967 81506
rect 59933 81440 59967 81456
rect 60269 81490 60303 81506
rect 60269 81440 60303 81456
rect 60605 81490 60639 81506
rect 60605 81440 60639 81456
rect 60941 81490 60975 81506
rect 60941 81440 60975 81456
rect 61277 81490 61311 81506
rect 61277 81440 61311 81456
rect 61613 81490 61647 81506
rect 61613 81440 61647 81456
rect 61949 81490 61983 81506
rect 61949 81440 61983 81456
rect 62285 81490 62319 81506
rect 62285 81440 62319 81456
rect 62621 81490 62655 81506
rect 62621 81440 62655 81456
rect 62957 81490 62991 81506
rect 62957 81440 62991 81456
rect 63293 81490 63327 81506
rect 63293 81440 63327 81456
rect 63629 81490 63663 81506
rect 63629 81440 63663 81456
rect 63965 81490 63999 81506
rect 63965 81440 63999 81456
rect 64301 81490 64335 81506
rect 64301 81440 64335 81456
rect 64637 81490 64671 81506
rect 64637 81440 64671 81456
rect 64973 81490 65007 81506
rect 64973 81440 65007 81456
rect 65309 81490 65343 81506
rect 65309 81440 65343 81456
rect 65645 81490 65679 81506
rect 65645 81440 65679 81456
rect 65981 81490 66015 81506
rect 65981 81440 66015 81456
rect 66317 81490 66351 81506
rect 66317 81440 66351 81456
rect 66653 81490 66687 81506
rect 66653 81440 66687 81456
rect 66989 81490 67023 81506
rect 66989 81440 67023 81456
rect 67325 81490 67359 81506
rect 67325 81440 67359 81456
rect 67661 81490 67695 81506
rect 67661 81440 67695 81456
rect 67997 81490 68031 81506
rect 67997 81440 68031 81456
rect 68333 81490 68367 81506
rect 68333 81440 68367 81456
rect 68669 81490 68703 81506
rect 68669 81440 68703 81456
rect 69005 81490 69039 81506
rect 69005 81440 69039 81456
rect 69341 81490 69375 81506
rect 69341 81440 69375 81456
rect 69677 81490 69711 81506
rect 69677 81440 69711 81456
rect 70013 81490 70047 81506
rect 70013 81440 70047 81456
rect 70349 81490 70383 81506
rect 70349 81440 70383 81456
rect 70685 81490 70719 81506
rect 70685 81440 70719 81456
rect 71021 81490 71055 81506
rect 71021 81440 71055 81456
rect 71357 81490 71391 81506
rect 71357 81440 71391 81456
rect 71693 81490 71727 81506
rect 71693 81440 71727 81456
rect 72029 81490 72063 81506
rect 72029 81440 72063 81456
rect 72365 81490 72399 81506
rect 72365 81440 72399 81456
rect 72701 81490 72735 81506
rect 72701 81440 72735 81456
rect 73037 81490 73071 81506
rect 73037 81440 73071 81456
rect 73373 81490 73407 81506
rect 73373 81440 73407 81456
rect 73709 81490 73743 81506
rect 73709 81440 73743 81456
rect 74045 81490 74079 81506
rect 74045 81440 74079 81456
rect 74381 81490 74415 81506
rect 74381 81440 74415 81456
rect 74717 81490 74751 81506
rect 74717 81440 74751 81456
rect 75053 81490 75087 81506
rect 75053 81440 75087 81456
rect 75389 81490 75423 81506
rect 75389 81440 75423 81456
rect 75725 81490 75759 81506
rect 75725 81440 75759 81456
rect 76061 81490 76095 81506
rect 76061 81440 76095 81456
rect 76397 81490 76431 81506
rect 76397 81440 76431 81456
rect 76733 81490 76767 81506
rect 76733 81440 76767 81456
rect 77069 81490 77103 81506
rect 77069 81440 77103 81456
rect 77405 81490 77439 81506
rect 77405 81440 77439 81456
rect 77741 81490 77775 81506
rect 77741 81440 77775 81456
rect 78077 81490 78111 81506
rect 78077 81440 78111 81456
rect 78413 81490 78447 81506
rect 78413 81440 78447 81456
rect 78749 81490 78783 81506
rect 78749 81440 78783 81456
rect 79085 81490 79119 81506
rect 79085 81440 79119 81456
rect 79421 81490 79455 81506
rect 79421 81440 79455 81456
rect 79757 81490 79791 81506
rect 79757 81440 79791 81456
rect 80093 81490 80127 81506
rect 80093 81440 80127 81456
rect 80429 81490 80463 81506
rect 80429 81440 80463 81456
rect 80765 81490 80799 81506
rect 80765 81440 80799 81456
rect 81101 81490 81135 81506
rect 81101 81440 81135 81456
rect 81437 81490 81471 81506
rect 81437 81440 81471 81456
rect 81773 81490 81807 81506
rect 81773 81440 81807 81456
rect 82109 81490 82143 81506
rect 82109 81440 82143 81456
rect 82445 81490 82479 81506
rect 82445 81440 82479 81456
rect 82781 81490 82815 81506
rect 82781 81440 82815 81456
rect 83117 81490 83151 81506
rect 83117 81440 83151 81456
rect 83453 81490 83487 81506
rect 83453 81440 83487 81456
rect 83789 81490 83823 81506
rect 83789 81440 83823 81456
rect 84125 81490 84159 81506
rect 84125 81440 84159 81456
rect 84461 81490 84495 81506
rect 84461 81440 84495 81456
rect 84797 81490 84831 81506
rect 84797 81440 84831 81456
rect 85133 81490 85167 81506
rect 85133 81440 85167 81456
rect 85469 81490 85503 81506
rect 85469 81440 85503 81456
rect 85805 81490 85839 81506
rect 85805 81440 85839 81456
rect 86141 81490 86175 81506
rect 86141 81440 86175 81456
rect 86477 81490 86511 81506
rect 86477 81440 86511 81456
rect 86813 81490 86847 81506
rect 86813 81440 86847 81456
rect 87149 81490 87183 81506
rect 87149 81440 87183 81456
rect 87485 81490 87519 81506
rect 87485 81440 87519 81456
rect 87821 81490 87855 81506
rect 87821 81440 87855 81456
rect 88157 81490 88191 81506
rect 88157 81440 88191 81456
rect 88493 81490 88527 81506
rect 88493 81440 88527 81456
rect 88829 81490 88863 81506
rect 88829 81440 88863 81456
rect 89165 81490 89199 81506
rect 89165 81440 89199 81456
rect 89501 81490 89535 81506
rect 89501 81440 89535 81456
rect 89837 81490 89871 81506
rect 89837 81440 89871 81456
rect 90173 81490 90207 81506
rect 90173 81440 90207 81456
rect 90509 81490 90543 81506
rect 90509 81440 90543 81456
rect 90845 81490 90879 81506
rect 90845 81440 90879 81456
rect 91181 81490 91215 81506
rect 91181 81440 91215 81456
rect 91517 81490 91551 81506
rect 91517 81440 91551 81456
rect 91853 81490 91887 81506
rect 91853 81440 91887 81456
rect 92189 81490 92223 81506
rect 92189 81440 92223 81456
rect 92525 81490 92559 81506
rect 92525 81440 92559 81456
rect 92861 81490 92895 81506
rect 92861 81440 92895 81456
rect 93197 81490 93231 81506
rect 93197 81440 93231 81456
rect 93533 81490 93567 81506
rect 93533 81440 93567 81456
rect 93869 81490 93903 81506
rect 93869 81440 93903 81456
rect 94205 81490 94239 81506
rect 94205 81440 94239 81456
rect 94541 81490 94575 81506
rect 94541 81440 94575 81456
rect 94877 81490 94911 81506
rect 94877 81440 94911 81456
rect 95213 81490 95247 81506
rect 95213 81440 95247 81456
rect 95549 81490 95583 81506
rect 95549 81440 95583 81456
rect 95885 81490 95919 81506
rect 95885 81440 95919 81456
rect 96221 81490 96255 81506
rect 96221 81440 96255 81456
rect 96557 81490 96591 81506
rect 96557 81440 96591 81456
rect 96893 81490 96927 81506
rect 96893 81440 96927 81456
rect 97229 81490 97263 81506
rect 97229 81440 97263 81456
rect 97565 81490 97599 81506
rect 97565 81440 97599 81456
rect 97901 81490 97935 81506
rect 97901 81440 97935 81456
rect 98237 81490 98271 81506
rect 98237 81440 98271 81456
rect 98573 81490 98607 81506
rect 98573 81440 98607 81456
rect 98909 81490 98943 81506
rect 98909 81440 98943 81456
rect 99245 81490 99279 81506
rect 99245 81440 99279 81456
rect 99581 81490 99615 81506
rect 99581 81440 99615 81456
rect 99917 81490 99951 81506
rect 99917 81440 99951 81456
rect 100253 81490 100287 81506
rect 100253 81440 100287 81456
rect 100589 81490 100623 81506
rect 100589 81440 100623 81456
rect 100925 81490 100959 81506
rect 100925 81440 100959 81456
rect 101261 81490 101295 81506
rect 101261 81440 101295 81456
rect 101597 81490 101631 81506
rect 101597 81440 101631 81456
rect 101933 81490 101967 81506
rect 101933 81440 101967 81456
rect 102269 81490 102303 81506
rect 102269 81440 102303 81456
rect 102605 81490 102639 81506
rect 102605 81440 102639 81456
rect 102941 81490 102975 81506
rect 102941 81440 102975 81456
rect 103277 81490 103311 81506
rect 103277 81440 103311 81456
rect 103613 81490 103647 81506
rect 103613 81440 103647 81456
rect 103949 81490 103983 81506
rect 103949 81440 103983 81456
rect 104285 81490 104319 81506
rect 104285 81440 104319 81456
rect 104621 81490 104655 81506
rect 104621 81440 104655 81456
rect 104957 81490 104991 81506
rect 104957 81440 104991 81456
rect 105293 81490 105327 81506
rect 105293 81440 105327 81456
rect 105629 81490 105663 81506
rect 105629 81440 105663 81456
rect 105965 81490 105999 81506
rect 105965 81440 105999 81456
rect 106301 81490 106335 81506
rect 106301 81440 106335 81456
rect 106637 81490 106671 81506
rect 106637 81440 106671 81456
rect 106973 81490 107007 81506
rect 106973 81440 107007 81456
rect 107309 81490 107343 81506
rect 107309 81440 107343 81456
rect 107645 81490 107679 81506
rect 107645 81440 107679 81456
rect 107981 81490 108015 81506
rect 107981 81440 108015 81456
rect 108317 81490 108351 81506
rect 108317 81440 108351 81456
rect 108653 81490 108687 81506
rect 108653 81440 108687 81456
rect 108989 81490 109023 81506
rect 108989 81440 109023 81456
rect 109325 81490 109359 81506
rect 109325 81440 109359 81456
rect 109661 81490 109695 81506
rect 109661 81440 109695 81456
rect 109997 81490 110031 81506
rect 109997 81440 110031 81456
rect 110333 81490 110367 81506
rect 110333 81440 110367 81456
rect 110669 81490 110703 81506
rect 110669 81440 110703 81456
rect 111005 81490 111039 81506
rect 111005 81440 111039 81456
rect 111341 81490 111375 81506
rect 111341 81440 111375 81456
rect 111677 81490 111711 81506
rect 111677 81440 111711 81456
rect 112013 81490 112047 81506
rect 112013 81440 112047 81456
rect 112349 81490 112383 81506
rect 112349 81440 112383 81456
rect 112685 81490 112719 81506
rect 112685 81440 112719 81456
rect 113021 81490 113055 81506
rect 113021 81440 113055 81456
rect 113357 81490 113391 81506
rect 113357 81440 113391 81456
rect 113693 81490 113727 81506
rect 113693 81440 113727 81456
rect 114029 81490 114063 81506
rect 114029 81440 114063 81456
rect 114365 81490 114399 81506
rect 114365 81440 114399 81456
rect 114701 81490 114735 81506
rect 114701 81440 114735 81456
rect 115037 81490 115071 81506
rect 115037 81440 115071 81456
rect 115373 81490 115407 81506
rect 115373 81440 115407 81456
rect 115709 81490 115743 81506
rect 115709 81440 115743 81456
rect 116045 81490 116079 81506
rect 116045 81440 116079 81456
rect 116381 81490 116415 81506
rect 116381 81440 116415 81456
rect 116717 81490 116751 81506
rect 116717 81440 116751 81456
rect 117053 81490 117087 81506
rect 117053 81440 117087 81456
rect 117389 81490 117423 81506
rect 117389 81440 117423 81456
rect 117725 81490 117759 81506
rect 117725 81440 117759 81456
rect 118061 81490 118095 81506
rect 118061 81440 118095 81456
rect 118397 81490 118431 81506
rect 118397 81440 118431 81456
rect 118733 81490 118767 81506
rect 118733 81440 118767 81456
rect 119069 81490 119103 81506
rect 119069 81440 119103 81456
rect 119405 81490 119439 81506
rect 119405 81440 119439 81456
rect 119741 81490 119775 81506
rect 119741 81440 119775 81456
rect 120077 81490 120111 81506
rect 120077 81440 120111 81456
rect 120413 81490 120447 81506
rect 120413 81440 120447 81456
rect 120749 81490 120783 81506
rect 120749 81440 120783 81456
rect 121085 81490 121119 81506
rect 121085 81440 121119 81456
rect 121421 81490 121455 81506
rect 121421 81440 121455 81456
rect 121757 81490 121791 81506
rect 121757 81440 121791 81456
rect 122093 81490 122127 81506
rect 122093 81440 122127 81456
rect 122429 81490 122463 81506
rect 122429 81440 122463 81456
rect 122765 81490 122799 81506
rect 122765 81440 122799 81456
rect 123101 81490 123135 81506
rect 123101 81440 123135 81456
rect 123437 81490 123471 81506
rect 123437 81440 123471 81456
rect 123773 81490 123807 81506
rect 123773 81440 123807 81456
rect 124109 81490 124143 81506
rect 124109 81440 124143 81456
rect 124445 81490 124479 81506
rect 124445 81440 124479 81456
rect 124781 81490 124815 81506
rect 124781 81440 124815 81456
rect 125117 81490 125151 81506
rect 125117 81440 125151 81456
rect 125453 81490 125487 81506
rect 125453 81440 125487 81456
rect 125789 81490 125823 81506
rect 125789 81440 125823 81456
rect 126125 81490 126159 81506
rect 126125 81440 126159 81456
rect 126461 81490 126495 81506
rect 126461 81440 126495 81456
rect 126797 81490 126831 81506
rect 126797 81440 126831 81456
rect 127133 81490 127167 81506
rect 127133 81440 127167 81456
rect 127469 81490 127503 81506
rect 127469 81440 127503 81456
rect 127805 81490 127839 81506
rect 127805 81440 127839 81456
rect 128141 81490 128175 81506
rect 128141 81440 128175 81456
rect 128477 81490 128511 81506
rect 128477 81440 128511 81456
rect 128813 81490 128847 81506
rect 128813 81440 128847 81456
rect 129149 81490 129183 81506
rect 129149 81440 129183 81456
rect 129485 81490 129519 81506
rect 129485 81440 129519 81456
rect 129821 81490 129855 81506
rect 129821 81440 129855 81456
rect 130157 81490 130191 81506
rect 130157 81440 130191 81456
rect 130493 81490 130527 81506
rect 130493 81440 130527 81456
rect 130829 81490 130863 81506
rect 130829 81440 130863 81456
rect 131165 81490 131199 81506
rect 131165 81440 131199 81456
rect 131501 81490 131535 81506
rect 131501 81440 131535 81456
rect 131837 81490 131871 81506
rect 131837 81440 131871 81456
rect 132173 81490 132207 81506
rect 132173 81440 132207 81456
rect 132509 81490 132543 81506
rect 132509 81440 132543 81456
rect 132845 81490 132879 81506
rect 132845 81440 132879 81456
rect 133181 81490 133215 81506
rect 133181 81440 133215 81456
rect 133517 81490 133551 81506
rect 133517 81440 133551 81456
rect 133853 81490 133887 81506
rect 133853 81440 133887 81456
rect 134189 81490 134223 81506
rect 134189 81440 134223 81456
rect 1805 81037 1839 81053
rect 1805 80987 1839 81003
rect 134855 81037 134889 81053
rect 134855 80987 134889 81003
rect 1805 80701 1839 80717
rect 1805 80651 1839 80667
rect 134855 80701 134889 80717
rect 134855 80651 134889 80667
rect 1805 80365 1839 80381
rect 1805 80315 1839 80331
rect 134855 80365 134889 80381
rect 134855 80315 134889 80331
rect 1805 80029 1839 80045
rect 1805 79979 1839 79995
rect 134855 80029 134889 80045
rect 134855 79979 134889 79995
rect 1805 79693 1839 79709
rect 1805 79643 1839 79659
rect 134855 79693 134889 79709
rect 134855 79643 134889 79659
rect 1805 79357 1839 79373
rect 1805 79307 1839 79323
rect 134855 79357 134889 79373
rect 134855 79307 134889 79323
rect 1805 79021 1839 79037
rect 1805 78971 1839 78987
rect 134855 79021 134889 79037
rect 134855 78971 134889 78987
rect 1805 78685 1839 78701
rect 1805 78635 1839 78651
rect 134855 78685 134889 78701
rect 134855 78635 134889 78651
rect 1805 78349 1839 78365
rect 1805 78299 1839 78315
rect 134855 78349 134889 78365
rect 134855 78299 134889 78315
rect 1805 78013 1839 78029
rect 1805 77963 1839 77979
rect 134855 78013 134889 78029
rect 134855 77963 134889 77979
rect 1805 77677 1839 77693
rect 1805 77627 1839 77643
rect 134855 77677 134889 77693
rect 134855 77627 134889 77643
rect 1805 77341 1839 77357
rect 1805 77291 1839 77307
rect 134855 77341 134889 77357
rect 134855 77291 134889 77307
rect 1805 77005 1839 77021
rect 1805 76955 1839 76971
rect 134855 77005 134889 77021
rect 134855 76955 134889 76971
rect 1805 76669 1839 76685
rect 1805 76619 1839 76635
rect 134855 76669 134889 76685
rect 134855 76619 134889 76635
rect 1805 76333 1839 76349
rect 1805 76283 1839 76299
rect 134855 76333 134889 76349
rect 134855 76283 134889 76299
rect 1805 75997 1839 76013
rect 1805 75947 1839 75963
rect 134855 75997 134889 76013
rect 134855 75947 134889 75963
rect 1805 75661 1839 75677
rect 1805 75611 1839 75627
rect 134855 75661 134889 75677
rect 134855 75611 134889 75627
rect 1805 75325 1839 75341
rect 1805 75275 1839 75291
rect 134855 75325 134889 75341
rect 134855 75275 134889 75291
rect 1805 74989 1839 75005
rect 1805 74939 1839 74955
rect 134855 74989 134889 75005
rect 134855 74939 134889 74955
rect 1805 74653 1839 74669
rect 1805 74603 1839 74619
rect 134855 74653 134889 74669
rect 134855 74603 134889 74619
rect 1805 74317 1839 74333
rect 1805 74267 1839 74283
rect 134855 74317 134889 74333
rect 134855 74267 134889 74283
rect 1805 73981 1839 73997
rect 1805 73931 1839 73947
rect 134855 73981 134889 73997
rect 134855 73931 134889 73947
rect 1805 73645 1839 73661
rect 1805 73595 1839 73611
rect 134855 73645 134889 73661
rect 134855 73595 134889 73611
rect 1805 73309 1839 73325
rect 1805 73259 1839 73275
rect 134855 73309 134889 73325
rect 134855 73259 134889 73275
rect 1805 72973 1839 72989
rect 1805 72923 1839 72939
rect 134855 72973 134889 72989
rect 134855 72923 134889 72939
rect 1805 72637 1839 72653
rect 1805 72587 1839 72603
rect 134855 72637 134889 72653
rect 134855 72587 134889 72603
rect 1805 72301 1839 72317
rect 1805 72251 1839 72267
rect 134855 72301 134889 72317
rect 134855 72251 134889 72267
rect 1805 71965 1839 71981
rect 1805 71915 1839 71931
rect 134855 71965 134889 71981
rect 134855 71915 134889 71931
rect 1805 71629 1839 71645
rect 1805 71579 1839 71595
rect 134855 71629 134889 71645
rect 134855 71579 134889 71595
rect 1805 71293 1839 71309
rect 1805 71243 1839 71259
rect 134855 71293 134889 71309
rect 134855 71243 134889 71259
rect 1805 70957 1839 70973
rect 1805 70907 1839 70923
rect 134855 70957 134889 70973
rect 134855 70907 134889 70923
rect 1805 70621 1839 70637
rect 1805 70571 1839 70587
rect 134855 70621 134889 70637
rect 134855 70571 134889 70587
rect 1805 70285 1839 70301
rect 1805 70235 1839 70251
rect 134855 70285 134889 70301
rect 134855 70235 134889 70251
rect 1805 69949 1839 69965
rect 1805 69899 1839 69915
rect 134855 69949 134889 69965
rect 134855 69899 134889 69915
rect 1805 69613 1839 69629
rect 1805 69563 1839 69579
rect 134855 69613 134889 69629
rect 134855 69563 134889 69579
rect 1805 69277 1839 69293
rect 1805 69227 1839 69243
rect 134855 69277 134889 69293
rect 134855 69227 134889 69243
rect 1805 68941 1839 68957
rect 1805 68891 1839 68907
rect 134855 68941 134889 68957
rect 134855 68891 134889 68907
rect 1805 68605 1839 68621
rect 1805 68555 1839 68571
rect 134855 68605 134889 68621
rect 134855 68555 134889 68571
rect 1805 68269 1839 68285
rect 1805 68219 1839 68235
rect 134855 68269 134889 68285
rect 134855 68219 134889 68235
rect 1805 67933 1839 67949
rect 1805 67883 1839 67899
rect 134855 67933 134889 67949
rect 134855 67883 134889 67899
rect 1805 67597 1839 67613
rect 1805 67547 1839 67563
rect 134855 67597 134889 67613
rect 134855 67547 134889 67563
rect 1805 67261 1839 67277
rect 1805 67211 1839 67227
rect 134855 67261 134889 67277
rect 134855 67211 134889 67227
rect 1805 66925 1839 66941
rect 1805 66875 1839 66891
rect 134855 66925 134889 66941
rect 134855 66875 134889 66891
rect 1805 66589 1839 66605
rect 1805 66539 1839 66555
rect 134855 66589 134889 66605
rect 134855 66539 134889 66555
rect 1805 66253 1839 66269
rect 1805 66203 1839 66219
rect 134855 66253 134889 66269
rect 134855 66203 134889 66219
rect 1805 65917 1839 65933
rect 1805 65867 1839 65883
rect 134855 65917 134889 65933
rect 134855 65867 134889 65883
rect 1805 65581 1839 65597
rect 1805 65531 1839 65547
rect 134855 65581 134889 65597
rect 134855 65531 134889 65547
rect 1805 65245 1839 65261
rect 1805 65195 1839 65211
rect 134855 65245 134889 65261
rect 134855 65195 134889 65211
rect 1805 64909 1839 64925
rect 1805 64859 1839 64875
rect 134855 64909 134889 64925
rect 134855 64859 134889 64875
rect 1805 64573 1839 64589
rect 1805 64523 1839 64539
rect 134855 64573 134889 64589
rect 134855 64523 134889 64539
rect 1805 64237 1839 64253
rect 1805 64187 1839 64203
rect 134855 64237 134889 64253
rect 134855 64187 134889 64203
rect 1805 63901 1839 63917
rect 1805 63851 1839 63867
rect 134855 63901 134889 63917
rect 134855 63851 134889 63867
rect 1805 63565 1839 63581
rect 1805 63515 1839 63531
rect 134855 63565 134889 63581
rect 134855 63515 134889 63531
rect 1805 63229 1839 63245
rect 1805 63179 1839 63195
rect 134855 63229 134889 63245
rect 134855 63179 134889 63195
rect 1805 62893 1839 62909
rect 1805 62843 1839 62859
rect 134855 62893 134889 62909
rect 134855 62843 134889 62859
rect 1805 62557 1839 62573
rect 1805 62507 1839 62523
rect 134855 62557 134889 62573
rect 134855 62507 134889 62523
rect 1805 62221 1839 62237
rect 1805 62171 1839 62187
rect 134855 62221 134889 62237
rect 134855 62171 134889 62187
rect 1805 61885 1839 61901
rect 1805 61835 1839 61851
rect 134855 61885 134889 61901
rect 134855 61835 134889 61851
rect 1805 61549 1839 61565
rect 1805 61499 1839 61515
rect 134855 61549 134889 61565
rect 134855 61499 134889 61515
rect 1805 61213 1839 61229
rect 1805 61163 1839 61179
rect 134855 61213 134889 61229
rect 134855 61163 134889 61179
rect 1805 60877 1839 60893
rect 1805 60827 1839 60843
rect 134855 60877 134889 60893
rect 134855 60827 134889 60843
rect 1805 60541 1839 60557
rect 1805 60491 1839 60507
rect 134855 60541 134889 60557
rect 134855 60491 134889 60507
rect 1805 60205 1839 60221
rect 1805 60155 1839 60171
rect 134855 60205 134889 60221
rect 134855 60155 134889 60171
rect 1805 59869 1839 59885
rect 1805 59819 1839 59835
rect 134855 59869 134889 59885
rect 134855 59819 134889 59835
rect 1805 59533 1839 59549
rect 1805 59483 1839 59499
rect 134855 59533 134889 59549
rect 134855 59483 134889 59499
rect 1805 59197 1839 59213
rect 1805 59147 1839 59163
rect 134855 59197 134889 59213
rect 134855 59147 134889 59163
rect 1805 58861 1839 58877
rect 1805 58811 1839 58827
rect 134855 58861 134889 58877
rect 134855 58811 134889 58827
rect 1805 58525 1839 58541
rect 1805 58475 1839 58491
rect 134855 58525 134889 58541
rect 134855 58475 134889 58491
rect 1805 58189 1839 58205
rect 1805 58139 1839 58155
rect 134855 58189 134889 58205
rect 134855 58139 134889 58155
rect 1805 57853 1839 57869
rect 1805 57803 1839 57819
rect 134855 57853 134889 57869
rect 134855 57803 134889 57819
rect 1805 57517 1839 57533
rect 1805 57467 1839 57483
rect 134855 57517 134889 57533
rect 134855 57467 134889 57483
rect 1805 57181 1839 57197
rect 1805 57131 1839 57147
rect 134855 57181 134889 57197
rect 134855 57131 134889 57147
rect 1805 56845 1839 56861
rect 1805 56795 1839 56811
rect 134855 56845 134889 56861
rect 134855 56795 134889 56811
rect 1805 56509 1839 56525
rect 1805 56459 1839 56475
rect 134855 56509 134889 56525
rect 134855 56459 134889 56475
rect 1805 56173 1839 56189
rect 1805 56123 1839 56139
rect 134855 56173 134889 56189
rect 134855 56123 134889 56139
rect 1805 55837 1839 55853
rect 1805 55787 1839 55803
rect 134855 55837 134889 55853
rect 134855 55787 134889 55803
rect 1805 55501 1839 55517
rect 1805 55451 1839 55467
rect 134855 55501 134889 55517
rect 134855 55451 134889 55467
rect 1805 55165 1839 55181
rect 1805 55115 1839 55131
rect 134855 55165 134889 55181
rect 134855 55115 134889 55131
rect 1805 54829 1839 54845
rect 1805 54779 1839 54795
rect 134855 54829 134889 54845
rect 134855 54779 134889 54795
rect 1805 54493 1839 54509
rect 1805 54443 1839 54459
rect 134855 54493 134889 54509
rect 134855 54443 134889 54459
rect 1805 54157 1839 54173
rect 1805 54107 1839 54123
rect 134855 54157 134889 54173
rect 134855 54107 134889 54123
rect 1805 53821 1839 53837
rect 1805 53771 1839 53787
rect 134855 53821 134889 53837
rect 134855 53771 134889 53787
rect 1805 53485 1839 53501
rect 1805 53435 1839 53451
rect 134855 53485 134889 53501
rect 134855 53435 134889 53451
rect 1805 53149 1839 53165
rect 1805 53099 1839 53115
rect 134855 53149 134889 53165
rect 134855 53099 134889 53115
rect 1805 52813 1839 52829
rect 1805 52763 1839 52779
rect 134855 52813 134889 52829
rect 134855 52763 134889 52779
rect 1805 52477 1839 52493
rect 1805 52427 1839 52443
rect 134855 52477 134889 52493
rect 134855 52427 134889 52443
rect 1805 52141 1839 52157
rect 1805 52091 1839 52107
rect 134855 52141 134889 52157
rect 134855 52091 134889 52107
rect 1805 51805 1839 51821
rect 1805 51755 1839 51771
rect 134855 51805 134889 51821
rect 134855 51755 134889 51771
rect 1805 51469 1839 51485
rect 1805 51419 1839 51435
rect 134855 51469 134889 51485
rect 134855 51419 134889 51435
rect 1805 51133 1839 51149
rect 1805 51083 1839 51099
rect 134855 51133 134889 51149
rect 134855 51083 134889 51099
rect 1805 50797 1839 50813
rect 1805 50747 1839 50763
rect 134855 50797 134889 50813
rect 134855 50747 134889 50763
rect 1805 50461 1839 50477
rect 1805 50411 1839 50427
rect 134855 50461 134889 50477
rect 134855 50411 134889 50427
rect 1805 50125 1839 50141
rect 1805 50075 1839 50091
rect 134855 50125 134889 50141
rect 134855 50075 134889 50091
rect 1805 49789 1839 49805
rect 1805 49739 1839 49755
rect 134855 49789 134889 49805
rect 134855 49739 134889 49755
rect 1805 49453 1839 49469
rect 1805 49403 1839 49419
rect 134855 49453 134889 49469
rect 134855 49403 134889 49419
rect 1805 49117 1839 49133
rect 1805 49067 1839 49083
rect 134855 49117 134889 49133
rect 134855 49067 134889 49083
rect 1805 48781 1839 48797
rect 1805 48731 1839 48747
rect 134855 48781 134889 48797
rect 134855 48731 134889 48747
rect 1805 48445 1839 48461
rect 1805 48395 1839 48411
rect 134855 48445 134889 48461
rect 134855 48395 134889 48411
rect 1805 48109 1839 48125
rect 1805 48059 1839 48075
rect 134855 48109 134889 48125
rect 134855 48059 134889 48075
rect 1805 47773 1839 47789
rect 1805 47723 1839 47739
rect 134855 47773 134889 47789
rect 134855 47723 134889 47739
rect 1805 47437 1839 47453
rect 1805 47387 1839 47403
rect 134855 47437 134889 47453
rect 134855 47387 134889 47403
rect 1805 47101 1839 47117
rect 1805 47051 1839 47067
rect 134855 47101 134889 47117
rect 134855 47051 134889 47067
rect 1805 46765 1839 46781
rect 1805 46715 1839 46731
rect 134855 46765 134889 46781
rect 134855 46715 134889 46731
rect 1805 46429 1839 46445
rect 1805 46379 1839 46395
rect 134855 46429 134889 46445
rect 134855 46379 134889 46395
rect 1805 46093 1839 46109
rect 1805 46043 1839 46059
rect 134855 46093 134889 46109
rect 134855 46043 134889 46059
rect 1805 45757 1839 45773
rect 1805 45707 1839 45723
rect 134855 45757 134889 45773
rect 134855 45707 134889 45723
rect 1805 45421 1839 45437
rect 1805 45371 1839 45387
rect 134855 45421 134889 45437
rect 134855 45371 134889 45387
rect 1805 45085 1839 45101
rect 1805 45035 1839 45051
rect 134855 45085 134889 45101
rect 134855 45035 134889 45051
rect 1805 44749 1839 44765
rect 1805 44699 1839 44715
rect 134855 44749 134889 44765
rect 134855 44699 134889 44715
rect 1805 44413 1839 44429
rect 1805 44363 1839 44379
rect 134855 44413 134889 44429
rect 134855 44363 134889 44379
rect 1805 44077 1839 44093
rect 1805 44027 1839 44043
rect 134855 44077 134889 44093
rect 134855 44027 134889 44043
rect 1805 43741 1839 43757
rect 1805 43691 1839 43707
rect 134855 43741 134889 43757
rect 134855 43691 134889 43707
rect 1805 43405 1839 43421
rect 1805 43355 1839 43371
rect 134855 43405 134889 43421
rect 134855 43355 134889 43371
rect 1805 43069 1839 43085
rect 1805 43019 1839 43035
rect 134855 43069 134889 43085
rect 134855 43019 134889 43035
rect 1805 42733 1839 42749
rect 1805 42683 1839 42699
rect 134855 42733 134889 42749
rect 134855 42683 134889 42699
rect 1805 42397 1839 42413
rect 1805 42347 1839 42363
rect 134855 42397 134889 42413
rect 134855 42347 134889 42363
rect 1805 42061 1839 42077
rect 1805 42011 1839 42027
rect 134855 42061 134889 42077
rect 134855 42011 134889 42027
rect 1805 41725 1839 41741
rect 1805 41675 1839 41691
rect 134855 41725 134889 41741
rect 134855 41675 134889 41691
rect 1805 41389 1839 41405
rect 1805 41339 1839 41355
rect 134855 41389 134889 41405
rect 134855 41339 134889 41355
rect 1805 41053 1839 41069
rect 1805 41003 1839 41019
rect 134855 41053 134889 41069
rect 134855 41003 134889 41019
rect 1805 40717 1839 40733
rect 1805 40667 1839 40683
rect 134855 40717 134889 40733
rect 134855 40667 134889 40683
rect 1805 40381 1839 40397
rect 1805 40331 1839 40347
rect 134855 40381 134889 40397
rect 134855 40331 134889 40347
rect 1805 40045 1839 40061
rect 1805 39995 1839 40011
rect 134855 40045 134889 40061
rect 134855 39995 134889 40011
rect 1805 39709 1839 39725
rect 1805 39659 1839 39675
rect 134855 39709 134889 39725
rect 134855 39659 134889 39675
rect 1805 39373 1839 39389
rect 1805 39323 1839 39339
rect 134855 39373 134889 39389
rect 134855 39323 134889 39339
rect 1805 39037 1839 39053
rect 1805 38987 1839 39003
rect 134855 39037 134889 39053
rect 134855 38987 134889 39003
rect 1805 38701 1839 38717
rect 1805 38651 1839 38667
rect 134855 38701 134889 38717
rect 134855 38651 134889 38667
rect 1805 38365 1839 38381
rect 1805 38315 1839 38331
rect 134855 38365 134889 38381
rect 134855 38315 134889 38331
rect 1805 38029 1839 38045
rect 1805 37979 1839 37995
rect 134855 38029 134889 38045
rect 134855 37979 134889 37995
rect 1805 37693 1839 37709
rect 1805 37643 1839 37659
rect 134855 37693 134889 37709
rect 134855 37643 134889 37659
rect 1805 37357 1839 37373
rect 1805 37307 1839 37323
rect 134855 37357 134889 37373
rect 134855 37307 134889 37323
rect 1805 37021 1839 37037
rect 1805 36971 1839 36987
rect 134855 37021 134889 37037
rect 134855 36971 134889 36987
rect 1805 36685 1839 36701
rect 1805 36635 1839 36651
rect 134855 36685 134889 36701
rect 134855 36635 134889 36651
rect 1805 36349 1839 36365
rect 1805 36299 1839 36315
rect 134855 36349 134889 36365
rect 134855 36299 134889 36315
rect 1805 36013 1839 36029
rect 1805 35963 1839 35979
rect 134855 36013 134889 36029
rect 134855 35963 134889 35979
rect 1805 35677 1839 35693
rect 1805 35627 1839 35643
rect 134855 35677 134889 35693
rect 134855 35627 134889 35643
rect 1805 35341 1839 35357
rect 1805 35291 1839 35307
rect 134855 35341 134889 35357
rect 134855 35291 134889 35307
rect 1805 35005 1839 35021
rect 1805 34955 1839 34971
rect 134855 35005 134889 35021
rect 134855 34955 134889 34971
rect 1805 34669 1839 34685
rect 1805 34619 1839 34635
rect 134855 34669 134889 34685
rect 134855 34619 134889 34635
rect 1805 34333 1839 34349
rect 1805 34283 1839 34299
rect 134855 34333 134889 34349
rect 134855 34283 134889 34299
rect 1805 33997 1839 34013
rect 1805 33947 1839 33963
rect 134855 33997 134889 34013
rect 134855 33947 134889 33963
rect 1805 33661 1839 33677
rect 1805 33611 1839 33627
rect 134855 33661 134889 33677
rect 134855 33611 134889 33627
rect 1805 33325 1839 33341
rect 1805 33275 1839 33291
rect 134855 33325 134889 33341
rect 134855 33275 134889 33291
rect 1805 32989 1839 33005
rect 1805 32939 1839 32955
rect 134855 32989 134889 33005
rect 134855 32939 134889 32955
rect 1805 32653 1839 32669
rect 1805 32603 1839 32619
rect 134855 32653 134889 32669
rect 134855 32603 134889 32619
rect 1805 32317 1839 32333
rect 1805 32267 1839 32283
rect 134855 32317 134889 32333
rect 134855 32267 134889 32283
rect 1805 31981 1839 31997
rect 1805 31931 1839 31947
rect 134855 31981 134889 31997
rect 134855 31931 134889 31947
rect 1805 31645 1839 31661
rect 1805 31595 1839 31611
rect 134855 31645 134889 31661
rect 134855 31595 134889 31611
rect 1805 31309 1839 31325
rect 1805 31259 1839 31275
rect 134855 31309 134889 31325
rect 134855 31259 134889 31275
rect 1805 30973 1839 30989
rect 1805 30923 1839 30939
rect 134855 30973 134889 30989
rect 134855 30923 134889 30939
rect 1805 30637 1839 30653
rect 1805 30587 1839 30603
rect 134855 30637 134889 30653
rect 134855 30587 134889 30603
rect 1805 30301 1839 30317
rect 1805 30251 1839 30267
rect 134855 30301 134889 30317
rect 134855 30251 134889 30267
rect 1805 29965 1839 29981
rect 1805 29915 1839 29931
rect 134855 29965 134889 29981
rect 134855 29915 134889 29931
rect 1805 29629 1839 29645
rect 1805 29579 1839 29595
rect 134855 29629 134889 29645
rect 134855 29579 134889 29595
rect 1805 29293 1839 29309
rect 1805 29243 1839 29259
rect 134855 29293 134889 29309
rect 134855 29243 134889 29259
rect 1805 28957 1839 28973
rect 1805 28907 1839 28923
rect 134855 28957 134889 28973
rect 134855 28907 134889 28923
rect 1805 28621 1839 28637
rect 1805 28571 1839 28587
rect 134855 28621 134889 28637
rect 134855 28571 134889 28587
rect 1805 28285 1839 28301
rect 1805 28235 1839 28251
rect 134855 28285 134889 28301
rect 134855 28235 134889 28251
rect 1805 27949 1839 27965
rect 1805 27899 1839 27915
rect 134855 27949 134889 27965
rect 134855 27899 134889 27915
rect 1805 27613 1839 27629
rect 1805 27563 1839 27579
rect 134855 27613 134889 27629
rect 134855 27563 134889 27579
rect 1805 27277 1839 27293
rect 1805 27227 1839 27243
rect 134855 27277 134889 27293
rect 134855 27227 134889 27243
rect 1805 26941 1839 26957
rect 1805 26891 1839 26907
rect 134855 26941 134889 26957
rect 134855 26891 134889 26907
rect 1805 26605 1839 26621
rect 1805 26555 1839 26571
rect 134855 26605 134889 26621
rect 134855 26555 134889 26571
rect 1805 26269 1839 26285
rect 1805 26219 1839 26235
rect 134855 26269 134889 26285
rect 134855 26219 134889 26235
rect 1805 25933 1839 25949
rect 1805 25883 1839 25899
rect 134855 25933 134889 25949
rect 134855 25883 134889 25899
rect 1805 25597 1839 25613
rect 1805 25547 1839 25563
rect 134855 25597 134889 25613
rect 134855 25547 134889 25563
rect 1805 25261 1839 25277
rect 1805 25211 1839 25227
rect 134855 25261 134889 25277
rect 134855 25211 134889 25227
rect 1805 24925 1839 24941
rect 1805 24875 1839 24891
rect 134855 24925 134889 24941
rect 134855 24875 134889 24891
rect 1805 24589 1839 24605
rect 1805 24539 1839 24555
rect 134855 24589 134889 24605
rect 134855 24539 134889 24555
rect 1805 24253 1839 24269
rect 1805 24203 1839 24219
rect 134855 24253 134889 24269
rect 134855 24203 134889 24219
rect 1805 23917 1839 23933
rect 1805 23867 1839 23883
rect 134855 23917 134889 23933
rect 134855 23867 134889 23883
rect 1805 23581 1839 23597
rect 1805 23531 1839 23547
rect 134855 23581 134889 23597
rect 134855 23531 134889 23547
rect 1805 23245 1839 23261
rect 1805 23195 1839 23211
rect 134855 23245 134889 23261
rect 134855 23195 134889 23211
rect 1805 22909 1839 22925
rect 1805 22859 1839 22875
rect 134855 22909 134889 22925
rect 134855 22859 134889 22875
rect 1805 22573 1839 22589
rect 1805 22523 1839 22539
rect 134855 22573 134889 22589
rect 134855 22523 134889 22539
rect 1805 22237 1839 22253
rect 1805 22187 1839 22203
rect 134855 22237 134889 22253
rect 134855 22187 134889 22203
rect 1805 21901 1839 21917
rect 1805 21851 1839 21867
rect 134855 21901 134889 21917
rect 134855 21851 134889 21867
rect 1805 21565 1839 21581
rect 1805 21515 1839 21531
rect 134855 21565 134889 21581
rect 134855 21515 134889 21531
rect 1805 21229 1839 21245
rect 1805 21179 1839 21195
rect 134855 21229 134889 21245
rect 134855 21179 134889 21195
rect 1805 20893 1839 20909
rect 1805 20843 1839 20859
rect 134855 20893 134889 20909
rect 134855 20843 134889 20859
rect 1805 20557 1839 20573
rect 1805 20507 1839 20523
rect 134855 20557 134889 20573
rect 134855 20507 134889 20523
rect 1805 20221 1839 20237
rect 1805 20171 1839 20187
rect 134855 20221 134889 20237
rect 134855 20171 134889 20187
rect 1805 19885 1839 19901
rect 1805 19835 1839 19851
rect 134855 19885 134889 19901
rect 134855 19835 134889 19851
rect 1805 19549 1839 19565
rect 1805 19499 1839 19515
rect 134855 19549 134889 19565
rect 134855 19499 134889 19515
rect 1805 19213 1839 19229
rect 1805 19163 1839 19179
rect 134855 19213 134889 19229
rect 134855 19163 134889 19179
rect 1805 18877 1839 18893
rect 1805 18827 1839 18843
rect 134855 18877 134889 18893
rect 134855 18827 134889 18843
rect 1805 18541 1839 18557
rect 1805 18491 1839 18507
rect 134855 18541 134889 18557
rect 134855 18491 134889 18507
rect 1805 18205 1839 18221
rect 1805 18155 1839 18171
rect 134855 18205 134889 18221
rect 134855 18155 134889 18171
rect 1805 17869 1839 17885
rect 1805 17819 1839 17835
rect 134855 17869 134889 17885
rect 134855 17819 134889 17835
rect 1805 17533 1839 17549
rect 1805 17483 1839 17499
rect 134855 17533 134889 17549
rect 134855 17483 134889 17499
rect 1805 17197 1839 17213
rect 1805 17147 1839 17163
rect 134855 17197 134889 17213
rect 134855 17147 134889 17163
rect 1805 16861 1839 16877
rect 1805 16811 1839 16827
rect 134855 16861 134889 16877
rect 134855 16811 134889 16827
rect 1805 16525 1839 16541
rect 1805 16475 1839 16491
rect 134855 16525 134889 16541
rect 134855 16475 134889 16491
rect 1805 16189 1839 16205
rect 1805 16139 1839 16155
rect 134855 16189 134889 16205
rect 134855 16139 134889 16155
rect 1805 15853 1839 15869
rect 1805 15803 1839 15819
rect 134855 15853 134889 15869
rect 134855 15803 134889 15819
rect 1805 15517 1839 15533
rect 1805 15467 1839 15483
rect 134855 15517 134889 15533
rect 134855 15467 134889 15483
rect 1805 15181 1839 15197
rect 1805 15131 1839 15147
rect 134855 15181 134889 15197
rect 134855 15131 134889 15147
rect 1805 14845 1839 14861
rect 1805 14795 1839 14811
rect 134855 14845 134889 14861
rect 134855 14795 134889 14811
rect 1805 14509 1839 14525
rect 1805 14459 1839 14475
rect 134855 14509 134889 14525
rect 134855 14459 134889 14475
rect 1805 14173 1839 14189
rect 1805 14123 1839 14139
rect 134855 14173 134889 14189
rect 134855 14123 134889 14139
rect 1805 13837 1839 13853
rect 1805 13787 1839 13803
rect 134855 13837 134889 13853
rect 134855 13787 134889 13803
rect 1805 13501 1839 13517
rect 1805 13451 1839 13467
rect 134855 13501 134889 13517
rect 134855 13451 134889 13467
rect 1805 13165 1839 13181
rect 1805 13115 1839 13131
rect 134855 13165 134889 13181
rect 134855 13115 134889 13131
rect 1805 12829 1839 12845
rect 1805 12779 1839 12795
rect 134855 12829 134889 12845
rect 134855 12779 134889 12795
rect 1805 12493 1839 12509
rect 1805 12443 1839 12459
rect 134855 12493 134889 12509
rect 134855 12443 134889 12459
rect 1805 12157 1839 12173
rect 1805 12107 1839 12123
rect 134855 12157 134889 12173
rect 134855 12107 134889 12123
rect 1805 11821 1839 11837
rect 1805 11771 1839 11787
rect 134855 11821 134889 11837
rect 134855 11771 134889 11787
rect 1805 11485 1839 11501
rect 1805 11435 1839 11451
rect 134855 11485 134889 11501
rect 134855 11435 134889 11451
rect 1805 11149 1839 11165
rect 1805 11099 1839 11115
rect 134855 11149 134889 11165
rect 134855 11099 134889 11115
rect 1805 10813 1839 10829
rect 1805 10763 1839 10779
rect 134855 10813 134889 10829
rect 134855 10763 134889 10779
rect 1805 10477 1839 10493
rect 1805 10427 1839 10443
rect 134855 10477 134889 10493
rect 134855 10427 134889 10443
rect 1805 10141 1839 10157
rect 1805 10091 1839 10107
rect 134855 10141 134889 10157
rect 134855 10091 134889 10107
rect 1805 9805 1839 9821
rect 1805 9755 1839 9771
rect 134855 9805 134889 9821
rect 134855 9755 134889 9771
rect 1805 9469 1839 9485
rect 1805 9419 1839 9435
rect 134855 9469 134889 9485
rect 134855 9419 134889 9435
rect 1805 9133 1839 9149
rect 1805 9083 1839 9099
rect 134855 9133 134889 9149
rect 134855 9083 134889 9099
rect 1805 8797 1839 8813
rect 1805 8747 1839 8763
rect 134855 8797 134889 8813
rect 134855 8747 134889 8763
rect 1805 8461 1839 8477
rect 1805 8411 1839 8427
rect 134855 8461 134889 8477
rect 134855 8411 134889 8427
rect 1805 8125 1839 8141
rect 1805 8075 1839 8091
rect 134855 8125 134889 8141
rect 134855 8075 134889 8091
rect 1805 7789 1839 7805
rect 1805 7739 1839 7755
rect 134855 7789 134889 7805
rect 134855 7739 134889 7755
rect 1805 7453 1839 7469
rect 1805 7403 1839 7419
rect 134855 7453 134889 7469
rect 134855 7403 134889 7419
rect 1805 7117 1839 7133
rect 1805 7067 1839 7083
rect 134855 7117 134889 7133
rect 134855 7067 134889 7083
rect 1805 6781 1839 6797
rect 1805 6731 1839 6747
rect 134855 6781 134889 6797
rect 134855 6731 134889 6747
rect 1805 6445 1839 6461
rect 1805 6395 1839 6411
rect 134855 6445 134889 6461
rect 134855 6395 134889 6411
rect 1805 6109 1839 6125
rect 1805 6059 1839 6075
rect 134855 6109 134889 6125
rect 134855 6059 134889 6075
rect 1805 5773 1839 5789
rect 1805 5723 1839 5739
rect 134855 5773 134889 5789
rect 134855 5723 134889 5739
rect 1805 5437 1839 5453
rect 1805 5387 1839 5403
rect 134855 5437 134889 5453
rect 134855 5387 134889 5403
rect 1805 5101 1839 5117
rect 1805 5051 1839 5067
rect 134855 5101 134889 5117
rect 134855 5051 134889 5067
rect 1805 4765 1839 4781
rect 1805 4715 1839 4731
rect 134855 4765 134889 4781
rect 134855 4715 134889 4731
rect 1805 4429 1839 4445
rect 1805 4379 1839 4395
rect 134855 4429 134889 4445
rect 134855 4379 134889 4395
rect 1805 4093 1839 4109
rect 1805 4043 1839 4059
rect 134855 4093 134889 4109
rect 134855 4043 134889 4059
rect 1805 3757 1839 3773
rect 1805 3707 1839 3723
rect 134855 3757 134889 3773
rect 134855 3707 134889 3723
rect 1805 3421 1839 3437
rect 1805 3371 1839 3387
rect 134855 3421 134889 3437
rect 134855 3371 134889 3387
rect 1805 3085 1839 3101
rect 1805 3035 1839 3051
rect 134855 3085 134889 3101
rect 134855 3035 134889 3051
rect 1805 2749 1839 2765
rect 1805 2699 1839 2715
rect 134855 2749 134889 2765
rect 134855 2699 134889 2715
rect 1805 2413 1839 2429
rect 1805 2363 1839 2379
rect 134855 2413 134889 2429
rect 134855 2363 134889 2379
rect 1805 2077 1839 2093
rect 1805 2027 1839 2043
rect 134855 2077 134889 2093
rect 134855 2027 134889 2043
rect 2141 1741 2175 1757
rect 2141 1691 2175 1707
rect 2477 1741 2511 1757
rect 2477 1691 2511 1707
rect 2813 1741 2847 1757
rect 2813 1691 2847 1707
rect 3149 1741 3183 1757
rect 3149 1691 3183 1707
rect 3485 1741 3519 1757
rect 3485 1691 3519 1707
rect 3821 1741 3855 1757
rect 3821 1691 3855 1707
rect 4157 1741 4191 1757
rect 4157 1691 4191 1707
rect 4493 1741 4527 1757
rect 4493 1691 4527 1707
rect 4829 1741 4863 1757
rect 4829 1691 4863 1707
rect 5165 1741 5199 1757
rect 5165 1691 5199 1707
rect 5501 1741 5535 1757
rect 5501 1691 5535 1707
rect 5837 1741 5871 1757
rect 5837 1691 5871 1707
rect 6173 1741 6207 1757
rect 6173 1691 6207 1707
rect 6509 1741 6543 1757
rect 6509 1691 6543 1707
rect 6845 1741 6879 1757
rect 6845 1691 6879 1707
rect 7181 1741 7215 1757
rect 7181 1691 7215 1707
rect 7517 1741 7551 1757
rect 7517 1691 7551 1707
rect 7853 1741 7887 1757
rect 7853 1691 7887 1707
rect 8189 1741 8223 1757
rect 8189 1691 8223 1707
rect 8525 1741 8559 1757
rect 8525 1691 8559 1707
rect 8861 1741 8895 1757
rect 8861 1691 8895 1707
rect 9197 1741 9231 1757
rect 9197 1691 9231 1707
rect 9533 1741 9567 1757
rect 9533 1691 9567 1707
rect 9869 1741 9903 1757
rect 9869 1691 9903 1707
rect 10205 1741 10239 1757
rect 10205 1691 10239 1707
rect 10541 1741 10575 1757
rect 10541 1691 10575 1707
rect 10877 1741 10911 1757
rect 10877 1691 10911 1707
rect 11213 1741 11247 1757
rect 11213 1691 11247 1707
rect 11549 1741 11583 1757
rect 11549 1691 11583 1707
rect 11885 1741 11919 1757
rect 11885 1691 11919 1707
rect 12221 1741 12255 1757
rect 12221 1691 12255 1707
rect 12557 1741 12591 1757
rect 12557 1691 12591 1707
rect 12893 1741 12927 1757
rect 12893 1691 12927 1707
rect 13229 1741 13263 1757
rect 13229 1691 13263 1707
rect 13565 1741 13599 1757
rect 13565 1691 13599 1707
rect 13901 1741 13935 1757
rect 13901 1691 13935 1707
rect 14237 1741 14271 1757
rect 14237 1691 14271 1707
rect 14573 1741 14607 1757
rect 14573 1691 14607 1707
rect 14909 1741 14943 1757
rect 14909 1691 14943 1707
rect 15245 1741 15279 1757
rect 15245 1691 15279 1707
rect 15581 1741 15615 1757
rect 15581 1691 15615 1707
rect 15917 1741 15951 1757
rect 15917 1691 15951 1707
rect 16253 1741 16287 1757
rect 16253 1691 16287 1707
rect 16589 1741 16623 1757
rect 16589 1691 16623 1707
rect 16925 1741 16959 1757
rect 16925 1691 16959 1707
rect 17261 1741 17295 1757
rect 17261 1691 17295 1707
rect 17597 1741 17631 1757
rect 17597 1691 17631 1707
rect 17933 1741 17967 1757
rect 17933 1691 17967 1707
rect 18269 1741 18303 1757
rect 18269 1691 18303 1707
rect 18605 1741 18639 1757
rect 18605 1691 18639 1707
rect 18941 1741 18975 1757
rect 18941 1691 18975 1707
rect 19277 1741 19311 1757
rect 19277 1691 19311 1707
rect 19613 1741 19647 1757
rect 19613 1691 19647 1707
rect 19949 1741 19983 1757
rect 19949 1691 19983 1707
rect 20285 1741 20319 1757
rect 20285 1691 20319 1707
rect 20621 1741 20655 1757
rect 20621 1691 20655 1707
rect 20957 1741 20991 1757
rect 20957 1691 20991 1707
rect 21293 1741 21327 1757
rect 21293 1691 21327 1707
rect 21629 1741 21663 1757
rect 21629 1691 21663 1707
rect 21965 1741 21999 1757
rect 21965 1691 21999 1707
rect 22301 1741 22335 1757
rect 22301 1691 22335 1707
rect 22637 1741 22671 1757
rect 22637 1691 22671 1707
rect 22973 1741 23007 1757
rect 22973 1691 23007 1707
rect 23309 1741 23343 1757
rect 23309 1691 23343 1707
rect 23645 1741 23679 1757
rect 23645 1691 23679 1707
rect 23981 1741 24015 1757
rect 23981 1691 24015 1707
rect 24317 1741 24351 1757
rect 24317 1691 24351 1707
rect 24653 1741 24687 1757
rect 24653 1691 24687 1707
rect 24989 1741 25023 1757
rect 24989 1691 25023 1707
rect 25325 1741 25359 1757
rect 25325 1691 25359 1707
rect 25661 1741 25695 1757
rect 25661 1691 25695 1707
rect 25997 1741 26031 1757
rect 25997 1691 26031 1707
rect 26333 1741 26367 1757
rect 26333 1691 26367 1707
rect 26669 1741 26703 1757
rect 26669 1691 26703 1707
rect 27005 1741 27039 1757
rect 27005 1691 27039 1707
rect 27341 1741 27375 1757
rect 27341 1691 27375 1707
rect 27677 1741 27711 1757
rect 27677 1691 27711 1707
rect 28013 1741 28047 1757
rect 28013 1691 28047 1707
rect 28349 1741 28383 1757
rect 28349 1691 28383 1707
rect 28685 1741 28719 1757
rect 28685 1691 28719 1707
rect 29021 1741 29055 1757
rect 29021 1691 29055 1707
rect 29357 1741 29391 1757
rect 29357 1691 29391 1707
rect 29693 1741 29727 1757
rect 29693 1691 29727 1707
rect 30029 1741 30063 1757
rect 30029 1691 30063 1707
rect 30365 1741 30399 1757
rect 30365 1691 30399 1707
rect 30701 1741 30735 1757
rect 30701 1691 30735 1707
rect 31037 1741 31071 1757
rect 31037 1691 31071 1707
rect 31373 1741 31407 1757
rect 31373 1691 31407 1707
rect 31709 1741 31743 1757
rect 31709 1691 31743 1707
rect 32045 1741 32079 1757
rect 32045 1691 32079 1707
rect 32381 1741 32415 1757
rect 32381 1691 32415 1707
rect 32717 1741 32751 1757
rect 32717 1691 32751 1707
rect 33053 1741 33087 1757
rect 33053 1691 33087 1707
rect 33389 1741 33423 1757
rect 33389 1691 33423 1707
rect 33725 1741 33759 1757
rect 33725 1691 33759 1707
rect 34061 1741 34095 1757
rect 34061 1691 34095 1707
rect 34397 1741 34431 1757
rect 34397 1691 34431 1707
rect 34733 1741 34767 1757
rect 34733 1691 34767 1707
rect 35069 1741 35103 1757
rect 35069 1691 35103 1707
rect 35405 1741 35439 1757
rect 35405 1691 35439 1707
rect 35741 1741 35775 1757
rect 35741 1691 35775 1707
rect 36077 1741 36111 1757
rect 36077 1691 36111 1707
rect 36413 1741 36447 1757
rect 36413 1691 36447 1707
rect 36749 1741 36783 1757
rect 36749 1691 36783 1707
rect 37085 1741 37119 1757
rect 37085 1691 37119 1707
rect 37421 1741 37455 1757
rect 37421 1691 37455 1707
rect 37757 1741 37791 1757
rect 37757 1691 37791 1707
rect 38093 1741 38127 1757
rect 38093 1691 38127 1707
rect 38429 1741 38463 1757
rect 38429 1691 38463 1707
rect 38765 1741 38799 1757
rect 38765 1691 38799 1707
rect 39101 1741 39135 1757
rect 39101 1691 39135 1707
rect 39437 1741 39471 1757
rect 39437 1691 39471 1707
rect 39773 1741 39807 1757
rect 39773 1691 39807 1707
rect 40109 1741 40143 1757
rect 40109 1691 40143 1707
rect 40445 1741 40479 1757
rect 40445 1691 40479 1707
rect 40781 1741 40815 1757
rect 40781 1691 40815 1707
rect 41117 1741 41151 1757
rect 41117 1691 41151 1707
rect 41453 1741 41487 1757
rect 41453 1691 41487 1707
rect 41789 1741 41823 1757
rect 41789 1691 41823 1707
rect 42125 1741 42159 1757
rect 42125 1691 42159 1707
rect 42461 1741 42495 1757
rect 42461 1691 42495 1707
rect 42797 1741 42831 1757
rect 42797 1691 42831 1707
rect 43133 1741 43167 1757
rect 43133 1691 43167 1707
rect 43469 1741 43503 1757
rect 43469 1691 43503 1707
rect 43805 1741 43839 1757
rect 43805 1691 43839 1707
rect 44141 1741 44175 1757
rect 44141 1691 44175 1707
rect 44477 1741 44511 1757
rect 44477 1691 44511 1707
rect 44813 1741 44847 1757
rect 44813 1691 44847 1707
rect 45149 1741 45183 1757
rect 45149 1691 45183 1707
rect 45485 1741 45519 1757
rect 45485 1691 45519 1707
rect 45821 1741 45855 1757
rect 45821 1691 45855 1707
rect 46157 1741 46191 1757
rect 46157 1691 46191 1707
rect 46493 1741 46527 1757
rect 46493 1691 46527 1707
rect 46829 1741 46863 1757
rect 46829 1691 46863 1707
rect 47165 1741 47199 1757
rect 47165 1691 47199 1707
rect 47501 1741 47535 1757
rect 47501 1691 47535 1707
rect 47837 1741 47871 1757
rect 47837 1691 47871 1707
rect 48173 1741 48207 1757
rect 48173 1691 48207 1707
rect 48509 1741 48543 1757
rect 48509 1691 48543 1707
rect 48845 1741 48879 1757
rect 48845 1691 48879 1707
rect 49181 1741 49215 1757
rect 49181 1691 49215 1707
rect 49517 1741 49551 1757
rect 49517 1691 49551 1707
rect 49853 1741 49887 1757
rect 49853 1691 49887 1707
rect 50189 1741 50223 1757
rect 50189 1691 50223 1707
rect 50525 1741 50559 1757
rect 50525 1691 50559 1707
rect 50861 1741 50895 1757
rect 50861 1691 50895 1707
rect 51197 1741 51231 1757
rect 51197 1691 51231 1707
rect 51533 1741 51567 1757
rect 51533 1691 51567 1707
rect 51869 1741 51903 1757
rect 51869 1691 51903 1707
rect 52205 1741 52239 1757
rect 52205 1691 52239 1707
rect 52541 1741 52575 1757
rect 52541 1691 52575 1707
rect 52877 1741 52911 1757
rect 52877 1691 52911 1707
rect 53213 1741 53247 1757
rect 53213 1691 53247 1707
rect 53549 1741 53583 1757
rect 53549 1691 53583 1707
rect 53885 1741 53919 1757
rect 53885 1691 53919 1707
rect 54221 1741 54255 1757
rect 54221 1691 54255 1707
rect 54557 1741 54591 1757
rect 54557 1691 54591 1707
rect 54893 1741 54927 1757
rect 54893 1691 54927 1707
rect 55229 1741 55263 1757
rect 55229 1691 55263 1707
rect 55565 1741 55599 1757
rect 55565 1691 55599 1707
rect 55901 1741 55935 1757
rect 55901 1691 55935 1707
rect 56237 1741 56271 1757
rect 56237 1691 56271 1707
rect 56573 1741 56607 1757
rect 56573 1691 56607 1707
rect 56909 1741 56943 1757
rect 56909 1691 56943 1707
rect 57245 1741 57279 1757
rect 57245 1691 57279 1707
rect 57581 1741 57615 1757
rect 57581 1691 57615 1707
rect 57917 1741 57951 1757
rect 57917 1691 57951 1707
rect 58253 1741 58287 1757
rect 58253 1691 58287 1707
rect 58589 1741 58623 1757
rect 58589 1691 58623 1707
rect 58925 1741 58959 1757
rect 58925 1691 58959 1707
rect 59261 1741 59295 1757
rect 59261 1691 59295 1707
rect 59597 1741 59631 1757
rect 59597 1691 59631 1707
rect 59933 1741 59967 1757
rect 59933 1691 59967 1707
rect 60269 1741 60303 1757
rect 60269 1691 60303 1707
rect 60605 1741 60639 1757
rect 60605 1691 60639 1707
rect 60941 1741 60975 1757
rect 60941 1691 60975 1707
rect 61277 1741 61311 1757
rect 61277 1691 61311 1707
rect 61613 1741 61647 1757
rect 61613 1691 61647 1707
rect 61949 1741 61983 1757
rect 61949 1691 61983 1707
rect 62285 1741 62319 1757
rect 62285 1691 62319 1707
rect 62621 1741 62655 1757
rect 62621 1691 62655 1707
rect 62957 1741 62991 1757
rect 62957 1691 62991 1707
rect 63293 1741 63327 1757
rect 63293 1691 63327 1707
rect 63629 1741 63663 1757
rect 63629 1691 63663 1707
rect 63965 1741 63999 1757
rect 63965 1691 63999 1707
rect 64301 1741 64335 1757
rect 64301 1691 64335 1707
rect 64637 1741 64671 1757
rect 64637 1691 64671 1707
rect 64973 1741 65007 1757
rect 64973 1691 65007 1707
rect 65309 1741 65343 1757
rect 65309 1691 65343 1707
rect 65645 1741 65679 1757
rect 65645 1691 65679 1707
rect 65981 1741 66015 1757
rect 65981 1691 66015 1707
rect 66317 1741 66351 1757
rect 66317 1691 66351 1707
rect 66653 1741 66687 1757
rect 66653 1691 66687 1707
rect 66989 1741 67023 1757
rect 66989 1691 67023 1707
rect 67325 1741 67359 1757
rect 67325 1691 67359 1707
rect 67661 1741 67695 1757
rect 67661 1691 67695 1707
rect 67997 1741 68031 1757
rect 67997 1691 68031 1707
rect 68333 1741 68367 1757
rect 68333 1691 68367 1707
rect 68669 1741 68703 1757
rect 68669 1691 68703 1707
rect 69005 1741 69039 1757
rect 69005 1691 69039 1707
rect 69341 1741 69375 1757
rect 69341 1691 69375 1707
rect 69677 1741 69711 1757
rect 69677 1691 69711 1707
rect 70013 1741 70047 1757
rect 70013 1691 70047 1707
rect 70349 1741 70383 1757
rect 70349 1691 70383 1707
rect 70685 1741 70719 1757
rect 70685 1691 70719 1707
rect 71021 1741 71055 1757
rect 71021 1691 71055 1707
rect 71357 1741 71391 1757
rect 71357 1691 71391 1707
rect 71693 1741 71727 1757
rect 71693 1691 71727 1707
rect 72029 1741 72063 1757
rect 72029 1691 72063 1707
rect 72365 1741 72399 1757
rect 72365 1691 72399 1707
rect 72701 1741 72735 1757
rect 72701 1691 72735 1707
rect 73037 1741 73071 1757
rect 73037 1691 73071 1707
rect 73373 1741 73407 1757
rect 73373 1691 73407 1707
rect 73709 1741 73743 1757
rect 73709 1691 73743 1707
rect 74045 1741 74079 1757
rect 74045 1691 74079 1707
rect 74381 1741 74415 1757
rect 74381 1691 74415 1707
rect 74717 1741 74751 1757
rect 74717 1691 74751 1707
rect 75053 1741 75087 1757
rect 75053 1691 75087 1707
rect 75389 1741 75423 1757
rect 75389 1691 75423 1707
rect 75725 1741 75759 1757
rect 75725 1691 75759 1707
rect 76061 1741 76095 1757
rect 76061 1691 76095 1707
rect 76397 1741 76431 1757
rect 76397 1691 76431 1707
rect 76733 1741 76767 1757
rect 76733 1691 76767 1707
rect 77069 1741 77103 1757
rect 77069 1691 77103 1707
rect 77405 1741 77439 1757
rect 77405 1691 77439 1707
rect 77741 1741 77775 1757
rect 77741 1691 77775 1707
rect 78077 1741 78111 1757
rect 78077 1691 78111 1707
rect 78413 1741 78447 1757
rect 78413 1691 78447 1707
rect 78749 1741 78783 1757
rect 78749 1691 78783 1707
rect 79085 1741 79119 1757
rect 79085 1691 79119 1707
rect 79421 1741 79455 1757
rect 79421 1691 79455 1707
rect 79757 1741 79791 1757
rect 79757 1691 79791 1707
rect 80093 1741 80127 1757
rect 80093 1691 80127 1707
rect 80429 1741 80463 1757
rect 80429 1691 80463 1707
rect 80765 1741 80799 1757
rect 80765 1691 80799 1707
rect 81101 1741 81135 1757
rect 81101 1691 81135 1707
rect 81437 1741 81471 1757
rect 81437 1691 81471 1707
rect 81773 1741 81807 1757
rect 81773 1691 81807 1707
rect 82109 1741 82143 1757
rect 82109 1691 82143 1707
rect 82445 1741 82479 1757
rect 82445 1691 82479 1707
rect 82781 1741 82815 1757
rect 82781 1691 82815 1707
rect 83117 1741 83151 1757
rect 83117 1691 83151 1707
rect 83453 1741 83487 1757
rect 83453 1691 83487 1707
rect 83789 1741 83823 1757
rect 83789 1691 83823 1707
rect 84125 1741 84159 1757
rect 84125 1691 84159 1707
rect 84461 1741 84495 1757
rect 84461 1691 84495 1707
rect 84797 1741 84831 1757
rect 84797 1691 84831 1707
rect 85133 1741 85167 1757
rect 85133 1691 85167 1707
rect 85469 1741 85503 1757
rect 85469 1691 85503 1707
rect 85805 1741 85839 1757
rect 85805 1691 85839 1707
rect 86141 1741 86175 1757
rect 86141 1691 86175 1707
rect 86477 1741 86511 1757
rect 86477 1691 86511 1707
rect 86813 1741 86847 1757
rect 86813 1691 86847 1707
rect 87149 1741 87183 1757
rect 87149 1691 87183 1707
rect 87485 1741 87519 1757
rect 87485 1691 87519 1707
rect 87821 1741 87855 1757
rect 87821 1691 87855 1707
rect 88157 1741 88191 1757
rect 88157 1691 88191 1707
rect 88493 1741 88527 1757
rect 88493 1691 88527 1707
rect 88829 1741 88863 1757
rect 88829 1691 88863 1707
rect 89165 1741 89199 1757
rect 89165 1691 89199 1707
rect 89501 1741 89535 1757
rect 89501 1691 89535 1707
rect 89837 1741 89871 1757
rect 89837 1691 89871 1707
rect 90173 1741 90207 1757
rect 90173 1691 90207 1707
rect 90509 1741 90543 1757
rect 90509 1691 90543 1707
rect 90845 1741 90879 1757
rect 90845 1691 90879 1707
rect 91181 1741 91215 1757
rect 91181 1691 91215 1707
rect 91517 1741 91551 1757
rect 91517 1691 91551 1707
rect 91853 1741 91887 1757
rect 91853 1691 91887 1707
rect 92189 1741 92223 1757
rect 92189 1691 92223 1707
rect 92525 1741 92559 1757
rect 92525 1691 92559 1707
rect 92861 1741 92895 1757
rect 92861 1691 92895 1707
rect 93197 1741 93231 1757
rect 93197 1691 93231 1707
rect 93533 1741 93567 1757
rect 93533 1691 93567 1707
rect 93869 1741 93903 1757
rect 93869 1691 93903 1707
rect 94205 1741 94239 1757
rect 94205 1691 94239 1707
rect 94541 1741 94575 1757
rect 94541 1691 94575 1707
rect 94877 1741 94911 1757
rect 94877 1691 94911 1707
rect 95213 1741 95247 1757
rect 95213 1691 95247 1707
rect 95549 1741 95583 1757
rect 95549 1691 95583 1707
rect 95885 1741 95919 1757
rect 95885 1691 95919 1707
rect 96221 1741 96255 1757
rect 96221 1691 96255 1707
rect 96557 1741 96591 1757
rect 96557 1691 96591 1707
rect 96893 1741 96927 1757
rect 96893 1691 96927 1707
rect 97229 1741 97263 1757
rect 97229 1691 97263 1707
rect 97565 1741 97599 1757
rect 97565 1691 97599 1707
rect 97901 1741 97935 1757
rect 97901 1691 97935 1707
rect 98237 1741 98271 1757
rect 98237 1691 98271 1707
rect 98573 1741 98607 1757
rect 98573 1691 98607 1707
rect 98909 1741 98943 1757
rect 98909 1691 98943 1707
rect 99245 1741 99279 1757
rect 99245 1691 99279 1707
rect 99581 1741 99615 1757
rect 99581 1691 99615 1707
rect 99917 1741 99951 1757
rect 99917 1691 99951 1707
rect 100253 1741 100287 1757
rect 100253 1691 100287 1707
rect 100589 1741 100623 1757
rect 100589 1691 100623 1707
rect 100925 1741 100959 1757
rect 100925 1691 100959 1707
rect 101261 1741 101295 1757
rect 101261 1691 101295 1707
rect 101597 1741 101631 1757
rect 101597 1691 101631 1707
rect 101933 1741 101967 1757
rect 101933 1691 101967 1707
rect 102269 1741 102303 1757
rect 102269 1691 102303 1707
rect 102605 1741 102639 1757
rect 102605 1691 102639 1707
rect 102941 1741 102975 1757
rect 102941 1691 102975 1707
rect 103277 1741 103311 1757
rect 103277 1691 103311 1707
rect 103613 1741 103647 1757
rect 103613 1691 103647 1707
rect 103949 1741 103983 1757
rect 103949 1691 103983 1707
rect 104285 1741 104319 1757
rect 104285 1691 104319 1707
rect 104621 1741 104655 1757
rect 104621 1691 104655 1707
rect 104957 1741 104991 1757
rect 104957 1691 104991 1707
rect 105293 1741 105327 1757
rect 105293 1691 105327 1707
rect 105629 1741 105663 1757
rect 105629 1691 105663 1707
rect 105965 1741 105999 1757
rect 105965 1691 105999 1707
rect 106301 1741 106335 1757
rect 106301 1691 106335 1707
rect 106637 1741 106671 1757
rect 106637 1691 106671 1707
rect 106973 1741 107007 1757
rect 106973 1691 107007 1707
rect 107309 1741 107343 1757
rect 107309 1691 107343 1707
rect 107645 1741 107679 1757
rect 107645 1691 107679 1707
rect 107981 1741 108015 1757
rect 107981 1691 108015 1707
rect 108317 1741 108351 1757
rect 108317 1691 108351 1707
rect 108653 1741 108687 1757
rect 108653 1691 108687 1707
rect 108989 1741 109023 1757
rect 108989 1691 109023 1707
rect 109325 1741 109359 1757
rect 109325 1691 109359 1707
rect 109661 1741 109695 1757
rect 109661 1691 109695 1707
rect 109997 1741 110031 1757
rect 109997 1691 110031 1707
rect 110333 1741 110367 1757
rect 110333 1691 110367 1707
rect 110669 1741 110703 1757
rect 110669 1691 110703 1707
rect 111005 1741 111039 1757
rect 111005 1691 111039 1707
rect 111341 1741 111375 1757
rect 111341 1691 111375 1707
rect 111677 1741 111711 1757
rect 111677 1691 111711 1707
rect 112013 1741 112047 1757
rect 112013 1691 112047 1707
rect 112349 1741 112383 1757
rect 112349 1691 112383 1707
rect 112685 1741 112719 1757
rect 112685 1691 112719 1707
rect 113021 1741 113055 1757
rect 113021 1691 113055 1707
rect 113357 1741 113391 1757
rect 113357 1691 113391 1707
rect 113693 1741 113727 1757
rect 113693 1691 113727 1707
rect 114029 1741 114063 1757
rect 114029 1691 114063 1707
rect 114365 1741 114399 1757
rect 114365 1691 114399 1707
rect 114701 1741 114735 1757
rect 114701 1691 114735 1707
rect 115037 1741 115071 1757
rect 115037 1691 115071 1707
rect 115373 1741 115407 1757
rect 115373 1691 115407 1707
rect 115709 1741 115743 1757
rect 115709 1691 115743 1707
rect 116045 1741 116079 1757
rect 116045 1691 116079 1707
rect 116381 1741 116415 1757
rect 116381 1691 116415 1707
rect 116717 1741 116751 1757
rect 116717 1691 116751 1707
rect 117053 1741 117087 1757
rect 117053 1691 117087 1707
rect 117389 1741 117423 1757
rect 117389 1691 117423 1707
rect 117725 1741 117759 1757
rect 117725 1691 117759 1707
rect 118061 1741 118095 1757
rect 118061 1691 118095 1707
rect 118397 1741 118431 1757
rect 118397 1691 118431 1707
rect 118733 1741 118767 1757
rect 118733 1691 118767 1707
rect 119069 1741 119103 1757
rect 119069 1691 119103 1707
rect 119405 1741 119439 1757
rect 119405 1691 119439 1707
rect 119741 1741 119775 1757
rect 119741 1691 119775 1707
rect 120077 1741 120111 1757
rect 120077 1691 120111 1707
rect 120413 1741 120447 1757
rect 120413 1691 120447 1707
rect 120749 1741 120783 1757
rect 120749 1691 120783 1707
rect 121085 1741 121119 1757
rect 121085 1691 121119 1707
rect 121421 1741 121455 1757
rect 121421 1691 121455 1707
rect 121757 1741 121791 1757
rect 121757 1691 121791 1707
rect 122093 1741 122127 1757
rect 122093 1691 122127 1707
rect 122429 1741 122463 1757
rect 122429 1691 122463 1707
rect 122765 1741 122799 1757
rect 122765 1691 122799 1707
rect 123101 1741 123135 1757
rect 123101 1691 123135 1707
rect 123437 1741 123471 1757
rect 123437 1691 123471 1707
rect 123773 1741 123807 1757
rect 123773 1691 123807 1707
rect 124109 1741 124143 1757
rect 124109 1691 124143 1707
rect 124445 1741 124479 1757
rect 124445 1691 124479 1707
rect 124781 1741 124815 1757
rect 124781 1691 124815 1707
rect 125117 1741 125151 1757
rect 125117 1691 125151 1707
rect 125453 1741 125487 1757
rect 125453 1691 125487 1707
rect 125789 1741 125823 1757
rect 125789 1691 125823 1707
rect 126125 1741 126159 1757
rect 126125 1691 126159 1707
rect 126461 1741 126495 1757
rect 126461 1691 126495 1707
rect 126797 1741 126831 1757
rect 126797 1691 126831 1707
rect 127133 1741 127167 1757
rect 127133 1691 127167 1707
rect 127469 1741 127503 1757
rect 127469 1691 127503 1707
rect 127805 1741 127839 1757
rect 127805 1691 127839 1707
rect 128141 1741 128175 1757
rect 128141 1691 128175 1707
rect 128477 1741 128511 1757
rect 128477 1691 128511 1707
rect 128813 1741 128847 1757
rect 128813 1691 128847 1707
rect 129149 1741 129183 1757
rect 129149 1691 129183 1707
rect 129485 1741 129519 1757
rect 129485 1691 129519 1707
rect 129821 1741 129855 1757
rect 129821 1691 129855 1707
rect 130157 1741 130191 1757
rect 130157 1691 130191 1707
rect 130493 1741 130527 1757
rect 130493 1691 130527 1707
rect 130829 1741 130863 1757
rect 130829 1691 130863 1707
rect 131165 1741 131199 1757
rect 131165 1691 131199 1707
rect 131501 1741 131535 1757
rect 131501 1691 131535 1707
rect 131837 1741 131871 1757
rect 131837 1691 131871 1707
rect 132173 1741 132207 1757
rect 132173 1691 132207 1707
rect 132509 1741 132543 1757
rect 132509 1691 132543 1707
rect 132845 1741 132879 1757
rect 132845 1691 132879 1707
rect 133181 1741 133215 1757
rect 133181 1691 133215 1707
rect 133517 1741 133551 1757
rect 133517 1691 133551 1707
rect 133853 1741 133887 1757
rect 133853 1691 133887 1707
rect 134189 1741 134223 1757
rect 134189 1691 134223 1707
<< viali >>
rect 2141 81456 2175 81490
rect 2477 81456 2511 81490
rect 2813 81456 2847 81490
rect 3149 81456 3183 81490
rect 3485 81456 3519 81490
rect 3821 81456 3855 81490
rect 4157 81456 4191 81490
rect 4493 81456 4527 81490
rect 4829 81456 4863 81490
rect 5165 81456 5199 81490
rect 5501 81456 5535 81490
rect 5837 81456 5871 81490
rect 6173 81456 6207 81490
rect 6509 81456 6543 81490
rect 6845 81456 6879 81490
rect 7181 81456 7215 81490
rect 7517 81456 7551 81490
rect 7853 81456 7887 81490
rect 8189 81456 8223 81490
rect 8525 81456 8559 81490
rect 8861 81456 8895 81490
rect 9197 81456 9231 81490
rect 9533 81456 9567 81490
rect 9869 81456 9903 81490
rect 10205 81456 10239 81490
rect 10541 81456 10575 81490
rect 10877 81456 10911 81490
rect 11213 81456 11247 81490
rect 11549 81456 11583 81490
rect 11885 81456 11919 81490
rect 12221 81456 12255 81490
rect 12557 81456 12591 81490
rect 12893 81456 12927 81490
rect 13229 81456 13263 81490
rect 13565 81456 13599 81490
rect 13901 81456 13935 81490
rect 14237 81456 14271 81490
rect 14573 81456 14607 81490
rect 14909 81456 14943 81490
rect 15245 81456 15279 81490
rect 15581 81456 15615 81490
rect 15917 81456 15951 81490
rect 16253 81456 16287 81490
rect 16589 81456 16623 81490
rect 16925 81456 16959 81490
rect 17261 81456 17295 81490
rect 17597 81456 17631 81490
rect 17933 81456 17967 81490
rect 18269 81456 18303 81490
rect 18605 81456 18639 81490
rect 18941 81456 18975 81490
rect 19277 81456 19311 81490
rect 19613 81456 19647 81490
rect 19949 81456 19983 81490
rect 20285 81456 20319 81490
rect 20621 81456 20655 81490
rect 20957 81456 20991 81490
rect 21293 81456 21327 81490
rect 21629 81456 21663 81490
rect 21965 81456 21999 81490
rect 22301 81456 22335 81490
rect 22637 81456 22671 81490
rect 22973 81456 23007 81490
rect 23309 81456 23343 81490
rect 23645 81456 23679 81490
rect 23981 81456 24015 81490
rect 24317 81456 24351 81490
rect 24653 81456 24687 81490
rect 24989 81456 25023 81490
rect 25325 81456 25359 81490
rect 25661 81456 25695 81490
rect 25997 81456 26031 81490
rect 26333 81456 26367 81490
rect 26669 81456 26703 81490
rect 27005 81456 27039 81490
rect 27341 81456 27375 81490
rect 27677 81456 27711 81490
rect 28013 81456 28047 81490
rect 28349 81456 28383 81490
rect 28685 81456 28719 81490
rect 29021 81456 29055 81490
rect 29357 81456 29391 81490
rect 29693 81456 29727 81490
rect 30029 81456 30063 81490
rect 30365 81456 30399 81490
rect 30701 81456 30735 81490
rect 31037 81456 31071 81490
rect 31373 81456 31407 81490
rect 31709 81456 31743 81490
rect 32045 81456 32079 81490
rect 32381 81456 32415 81490
rect 32717 81456 32751 81490
rect 33053 81456 33087 81490
rect 33389 81456 33423 81490
rect 33725 81456 33759 81490
rect 34061 81456 34095 81490
rect 34397 81456 34431 81490
rect 34733 81456 34767 81490
rect 35069 81456 35103 81490
rect 35405 81456 35439 81490
rect 35741 81456 35775 81490
rect 36077 81456 36111 81490
rect 36413 81456 36447 81490
rect 36749 81456 36783 81490
rect 37085 81456 37119 81490
rect 37421 81456 37455 81490
rect 37757 81456 37791 81490
rect 38093 81456 38127 81490
rect 38429 81456 38463 81490
rect 38765 81456 38799 81490
rect 39101 81456 39135 81490
rect 39437 81456 39471 81490
rect 39773 81456 39807 81490
rect 40109 81456 40143 81490
rect 40445 81456 40479 81490
rect 40781 81456 40815 81490
rect 41117 81456 41151 81490
rect 41453 81456 41487 81490
rect 41789 81456 41823 81490
rect 42125 81456 42159 81490
rect 42461 81456 42495 81490
rect 42797 81456 42831 81490
rect 43133 81456 43167 81490
rect 43469 81456 43503 81490
rect 43805 81456 43839 81490
rect 44141 81456 44175 81490
rect 44477 81456 44511 81490
rect 44813 81456 44847 81490
rect 45149 81456 45183 81490
rect 45485 81456 45519 81490
rect 45821 81456 45855 81490
rect 46157 81456 46191 81490
rect 46493 81456 46527 81490
rect 46829 81456 46863 81490
rect 47165 81456 47199 81490
rect 47501 81456 47535 81490
rect 47837 81456 47871 81490
rect 48173 81456 48207 81490
rect 48509 81456 48543 81490
rect 48845 81456 48879 81490
rect 49181 81456 49215 81490
rect 49517 81456 49551 81490
rect 49853 81456 49887 81490
rect 50189 81456 50223 81490
rect 50525 81456 50559 81490
rect 50861 81456 50895 81490
rect 51197 81456 51231 81490
rect 51533 81456 51567 81490
rect 51869 81456 51903 81490
rect 52205 81456 52239 81490
rect 52541 81456 52575 81490
rect 52877 81456 52911 81490
rect 53213 81456 53247 81490
rect 53549 81456 53583 81490
rect 53885 81456 53919 81490
rect 54221 81456 54255 81490
rect 54557 81456 54591 81490
rect 54893 81456 54927 81490
rect 55229 81456 55263 81490
rect 55565 81456 55599 81490
rect 55901 81456 55935 81490
rect 56237 81456 56271 81490
rect 56573 81456 56607 81490
rect 56909 81456 56943 81490
rect 57245 81456 57279 81490
rect 57581 81456 57615 81490
rect 57917 81456 57951 81490
rect 58253 81456 58287 81490
rect 58589 81456 58623 81490
rect 58925 81456 58959 81490
rect 59261 81456 59295 81490
rect 59597 81456 59631 81490
rect 59933 81456 59967 81490
rect 60269 81456 60303 81490
rect 60605 81456 60639 81490
rect 60941 81456 60975 81490
rect 61277 81456 61311 81490
rect 61613 81456 61647 81490
rect 61949 81456 61983 81490
rect 62285 81456 62319 81490
rect 62621 81456 62655 81490
rect 62957 81456 62991 81490
rect 63293 81456 63327 81490
rect 63629 81456 63663 81490
rect 63965 81456 63999 81490
rect 64301 81456 64335 81490
rect 64637 81456 64671 81490
rect 64973 81456 65007 81490
rect 65309 81456 65343 81490
rect 65645 81456 65679 81490
rect 65981 81456 66015 81490
rect 66317 81456 66351 81490
rect 66653 81456 66687 81490
rect 66989 81456 67023 81490
rect 67325 81456 67359 81490
rect 67661 81456 67695 81490
rect 67997 81456 68031 81490
rect 68333 81456 68367 81490
rect 68669 81456 68703 81490
rect 69005 81456 69039 81490
rect 69341 81456 69375 81490
rect 69677 81456 69711 81490
rect 70013 81456 70047 81490
rect 70349 81456 70383 81490
rect 70685 81456 70719 81490
rect 71021 81456 71055 81490
rect 71357 81456 71391 81490
rect 71693 81456 71727 81490
rect 72029 81456 72063 81490
rect 72365 81456 72399 81490
rect 72701 81456 72735 81490
rect 73037 81456 73071 81490
rect 73373 81456 73407 81490
rect 73709 81456 73743 81490
rect 74045 81456 74079 81490
rect 74381 81456 74415 81490
rect 74717 81456 74751 81490
rect 75053 81456 75087 81490
rect 75389 81456 75423 81490
rect 75725 81456 75759 81490
rect 76061 81456 76095 81490
rect 76397 81456 76431 81490
rect 76733 81456 76767 81490
rect 77069 81456 77103 81490
rect 77405 81456 77439 81490
rect 77741 81456 77775 81490
rect 78077 81456 78111 81490
rect 78413 81456 78447 81490
rect 78749 81456 78783 81490
rect 79085 81456 79119 81490
rect 79421 81456 79455 81490
rect 79757 81456 79791 81490
rect 80093 81456 80127 81490
rect 80429 81456 80463 81490
rect 80765 81456 80799 81490
rect 81101 81456 81135 81490
rect 81437 81456 81471 81490
rect 81773 81456 81807 81490
rect 82109 81456 82143 81490
rect 82445 81456 82479 81490
rect 82781 81456 82815 81490
rect 83117 81456 83151 81490
rect 83453 81456 83487 81490
rect 83789 81456 83823 81490
rect 84125 81456 84159 81490
rect 84461 81456 84495 81490
rect 84797 81456 84831 81490
rect 85133 81456 85167 81490
rect 85469 81456 85503 81490
rect 85805 81456 85839 81490
rect 86141 81456 86175 81490
rect 86477 81456 86511 81490
rect 86813 81456 86847 81490
rect 87149 81456 87183 81490
rect 87485 81456 87519 81490
rect 87821 81456 87855 81490
rect 88157 81456 88191 81490
rect 88493 81456 88527 81490
rect 88829 81456 88863 81490
rect 89165 81456 89199 81490
rect 89501 81456 89535 81490
rect 89837 81456 89871 81490
rect 90173 81456 90207 81490
rect 90509 81456 90543 81490
rect 90845 81456 90879 81490
rect 91181 81456 91215 81490
rect 91517 81456 91551 81490
rect 91853 81456 91887 81490
rect 92189 81456 92223 81490
rect 92525 81456 92559 81490
rect 92861 81456 92895 81490
rect 93197 81456 93231 81490
rect 93533 81456 93567 81490
rect 93869 81456 93903 81490
rect 94205 81456 94239 81490
rect 94541 81456 94575 81490
rect 94877 81456 94911 81490
rect 95213 81456 95247 81490
rect 95549 81456 95583 81490
rect 95885 81456 95919 81490
rect 96221 81456 96255 81490
rect 96557 81456 96591 81490
rect 96893 81456 96927 81490
rect 97229 81456 97263 81490
rect 97565 81456 97599 81490
rect 97901 81456 97935 81490
rect 98237 81456 98271 81490
rect 98573 81456 98607 81490
rect 98909 81456 98943 81490
rect 99245 81456 99279 81490
rect 99581 81456 99615 81490
rect 99917 81456 99951 81490
rect 100253 81456 100287 81490
rect 100589 81456 100623 81490
rect 100925 81456 100959 81490
rect 101261 81456 101295 81490
rect 101597 81456 101631 81490
rect 101933 81456 101967 81490
rect 102269 81456 102303 81490
rect 102605 81456 102639 81490
rect 102941 81456 102975 81490
rect 103277 81456 103311 81490
rect 103613 81456 103647 81490
rect 103949 81456 103983 81490
rect 104285 81456 104319 81490
rect 104621 81456 104655 81490
rect 104957 81456 104991 81490
rect 105293 81456 105327 81490
rect 105629 81456 105663 81490
rect 105965 81456 105999 81490
rect 106301 81456 106335 81490
rect 106637 81456 106671 81490
rect 106973 81456 107007 81490
rect 107309 81456 107343 81490
rect 107645 81456 107679 81490
rect 107981 81456 108015 81490
rect 108317 81456 108351 81490
rect 108653 81456 108687 81490
rect 108989 81456 109023 81490
rect 109325 81456 109359 81490
rect 109661 81456 109695 81490
rect 109997 81456 110031 81490
rect 110333 81456 110367 81490
rect 110669 81456 110703 81490
rect 111005 81456 111039 81490
rect 111341 81456 111375 81490
rect 111677 81456 111711 81490
rect 112013 81456 112047 81490
rect 112349 81456 112383 81490
rect 112685 81456 112719 81490
rect 113021 81456 113055 81490
rect 113357 81456 113391 81490
rect 113693 81456 113727 81490
rect 114029 81456 114063 81490
rect 114365 81456 114399 81490
rect 114701 81456 114735 81490
rect 115037 81456 115071 81490
rect 115373 81456 115407 81490
rect 115709 81456 115743 81490
rect 116045 81456 116079 81490
rect 116381 81456 116415 81490
rect 116717 81456 116751 81490
rect 117053 81456 117087 81490
rect 117389 81456 117423 81490
rect 117725 81456 117759 81490
rect 118061 81456 118095 81490
rect 118397 81456 118431 81490
rect 118733 81456 118767 81490
rect 119069 81456 119103 81490
rect 119405 81456 119439 81490
rect 119741 81456 119775 81490
rect 120077 81456 120111 81490
rect 120413 81456 120447 81490
rect 120749 81456 120783 81490
rect 121085 81456 121119 81490
rect 121421 81456 121455 81490
rect 121757 81456 121791 81490
rect 122093 81456 122127 81490
rect 122429 81456 122463 81490
rect 122765 81456 122799 81490
rect 123101 81456 123135 81490
rect 123437 81456 123471 81490
rect 123773 81456 123807 81490
rect 124109 81456 124143 81490
rect 124445 81456 124479 81490
rect 124781 81456 124815 81490
rect 125117 81456 125151 81490
rect 125453 81456 125487 81490
rect 125789 81456 125823 81490
rect 126125 81456 126159 81490
rect 126461 81456 126495 81490
rect 126797 81456 126831 81490
rect 127133 81456 127167 81490
rect 127469 81456 127503 81490
rect 127805 81456 127839 81490
rect 128141 81456 128175 81490
rect 128477 81456 128511 81490
rect 128813 81456 128847 81490
rect 129149 81456 129183 81490
rect 129485 81456 129519 81490
rect 129821 81456 129855 81490
rect 130157 81456 130191 81490
rect 130493 81456 130527 81490
rect 130829 81456 130863 81490
rect 131165 81456 131199 81490
rect 131501 81456 131535 81490
rect 131837 81456 131871 81490
rect 132173 81456 132207 81490
rect 132509 81456 132543 81490
rect 132845 81456 132879 81490
rect 133181 81456 133215 81490
rect 133517 81456 133551 81490
rect 133853 81456 133887 81490
rect 134189 81456 134223 81490
rect 1805 81003 1839 81037
rect 134855 81003 134889 81037
rect 1805 80667 1839 80701
rect 134855 80667 134889 80701
rect 1805 80331 1839 80365
rect 134855 80331 134889 80365
rect 1805 79995 1839 80029
rect 134855 79995 134889 80029
rect 1805 79659 1839 79693
rect 134855 79659 134889 79693
rect 1805 79323 1839 79357
rect 134855 79323 134889 79357
rect 1805 78987 1839 79021
rect 134855 78987 134889 79021
rect 1805 78651 1839 78685
rect 134855 78651 134889 78685
rect 1805 78315 1839 78349
rect 134855 78315 134889 78349
rect 1805 77979 1839 78013
rect 134855 77979 134889 78013
rect 1805 77643 1839 77677
rect 134855 77643 134889 77677
rect 1805 77307 1839 77341
rect 134855 77307 134889 77341
rect 1805 76971 1839 77005
rect 134855 76971 134889 77005
rect 1805 76635 1839 76669
rect 134855 76635 134889 76669
rect 1805 76299 1839 76333
rect 134855 76299 134889 76333
rect 1805 75963 1839 75997
rect 134855 75963 134889 75997
rect 1805 75627 1839 75661
rect 134855 75627 134889 75661
rect 1805 75291 1839 75325
rect 134855 75291 134889 75325
rect 1805 74955 1839 74989
rect 134855 74955 134889 74989
rect 1805 74619 1839 74653
rect 134855 74619 134889 74653
rect 1805 74283 1839 74317
rect 134855 74283 134889 74317
rect 1805 73947 1839 73981
rect 134855 73947 134889 73981
rect 1805 73611 1839 73645
rect 134855 73611 134889 73645
rect 1805 73275 1839 73309
rect 134855 73275 134889 73309
rect 1805 72939 1839 72973
rect 134855 72939 134889 72973
rect 1805 72603 1839 72637
rect 134855 72603 134889 72637
rect 1805 72267 1839 72301
rect 134855 72267 134889 72301
rect 1805 71931 1839 71965
rect 134855 71931 134889 71965
rect 1805 71595 1839 71629
rect 134855 71595 134889 71629
rect 1805 71259 1839 71293
rect 134855 71259 134889 71293
rect 1805 70923 1839 70957
rect 134855 70923 134889 70957
rect 1805 70587 1839 70621
rect 134855 70587 134889 70621
rect 1805 70251 1839 70285
rect 134855 70251 134889 70285
rect 1805 69915 1839 69949
rect 134855 69915 134889 69949
rect 1805 69579 1839 69613
rect 134855 69579 134889 69613
rect 1805 69243 1839 69277
rect 134855 69243 134889 69277
rect 1805 68907 1839 68941
rect 134855 68907 134889 68941
rect 1805 68571 1839 68605
rect 134855 68571 134889 68605
rect 1805 68235 1839 68269
rect 134855 68235 134889 68269
rect 1805 67899 1839 67933
rect 134855 67899 134889 67933
rect 1805 67563 1839 67597
rect 134855 67563 134889 67597
rect 1805 67227 1839 67261
rect 134855 67227 134889 67261
rect 1805 66891 1839 66925
rect 134855 66891 134889 66925
rect 1805 66555 1839 66589
rect 134855 66555 134889 66589
rect 1805 66219 1839 66253
rect 134855 66219 134889 66253
rect 1805 65883 1839 65917
rect 134855 65883 134889 65917
rect 1805 65547 1839 65581
rect 134855 65547 134889 65581
rect 1805 65211 1839 65245
rect 134855 65211 134889 65245
rect 1805 64875 1839 64909
rect 134855 64875 134889 64909
rect 1805 64539 1839 64573
rect 134855 64539 134889 64573
rect 1805 64203 1839 64237
rect 134855 64203 134889 64237
rect 1805 63867 1839 63901
rect 134855 63867 134889 63901
rect 1805 63531 1839 63565
rect 134855 63531 134889 63565
rect 1805 63195 1839 63229
rect 134855 63195 134889 63229
rect 1805 62859 1839 62893
rect 134855 62859 134889 62893
rect 1805 62523 1839 62557
rect 134855 62523 134889 62557
rect 1805 62187 1839 62221
rect 134855 62187 134889 62221
rect 1805 61851 1839 61885
rect 134855 61851 134889 61885
rect 1805 61515 1839 61549
rect 134855 61515 134889 61549
rect 1805 61179 1839 61213
rect 134855 61179 134889 61213
rect 1805 60843 1839 60877
rect 134855 60843 134889 60877
rect 1805 60507 1839 60541
rect 134855 60507 134889 60541
rect 1805 60171 1839 60205
rect 134855 60171 134889 60205
rect 1805 59835 1839 59869
rect 134855 59835 134889 59869
rect 1805 59499 1839 59533
rect 134855 59499 134889 59533
rect 1805 59163 1839 59197
rect 134855 59163 134889 59197
rect 1805 58827 1839 58861
rect 134855 58827 134889 58861
rect 1805 58491 1839 58525
rect 134855 58491 134889 58525
rect 1805 58155 1839 58189
rect 134855 58155 134889 58189
rect 1805 57819 1839 57853
rect 134855 57819 134889 57853
rect 1805 57483 1839 57517
rect 134855 57483 134889 57517
rect 1805 57147 1839 57181
rect 134855 57147 134889 57181
rect 1805 56811 1839 56845
rect 134855 56811 134889 56845
rect 1805 56475 1839 56509
rect 134855 56475 134889 56509
rect 1805 56139 1839 56173
rect 134855 56139 134889 56173
rect 1805 55803 1839 55837
rect 134855 55803 134889 55837
rect 1805 55467 1839 55501
rect 134855 55467 134889 55501
rect 1805 55131 1839 55165
rect 134855 55131 134889 55165
rect 1805 54795 1839 54829
rect 134855 54795 134889 54829
rect 1805 54459 1839 54493
rect 134855 54459 134889 54493
rect 1805 54123 1839 54157
rect 134855 54123 134889 54157
rect 1805 53787 1839 53821
rect 134855 53787 134889 53821
rect 1805 53451 1839 53485
rect 134855 53451 134889 53485
rect 1805 53115 1839 53149
rect 134855 53115 134889 53149
rect 1805 52779 1839 52813
rect 134855 52779 134889 52813
rect 1805 52443 1839 52477
rect 134855 52443 134889 52477
rect 1805 52107 1839 52141
rect 134855 52107 134889 52141
rect 1805 51771 1839 51805
rect 134855 51771 134889 51805
rect 1805 51435 1839 51469
rect 134855 51435 134889 51469
rect 1805 51099 1839 51133
rect 134855 51099 134889 51133
rect 1805 50763 1839 50797
rect 134855 50763 134889 50797
rect 1805 50427 1839 50461
rect 134855 50427 134889 50461
rect 1805 50091 1839 50125
rect 134855 50091 134889 50125
rect 1805 49755 1839 49789
rect 134855 49755 134889 49789
rect 1805 49419 1839 49453
rect 134855 49419 134889 49453
rect 1805 49083 1839 49117
rect 134855 49083 134889 49117
rect 1805 48747 1839 48781
rect 134855 48747 134889 48781
rect 1805 48411 1839 48445
rect 134855 48411 134889 48445
rect 1805 48075 1839 48109
rect 134855 48075 134889 48109
rect 1805 47739 1839 47773
rect 134855 47739 134889 47773
rect 1805 47403 1839 47437
rect 134855 47403 134889 47437
rect 1805 47067 1839 47101
rect 134855 47067 134889 47101
rect 1805 46731 1839 46765
rect 134855 46731 134889 46765
rect 1805 46395 1839 46429
rect 134855 46395 134889 46429
rect 1805 46059 1839 46093
rect 134855 46059 134889 46093
rect 1805 45723 1839 45757
rect 134855 45723 134889 45757
rect 1805 45387 1839 45421
rect 134855 45387 134889 45421
rect 1805 45051 1839 45085
rect 134855 45051 134889 45085
rect 1805 44715 1839 44749
rect 134855 44715 134889 44749
rect 1805 44379 1839 44413
rect 134855 44379 134889 44413
rect 1805 44043 1839 44077
rect 134855 44043 134889 44077
rect 1805 43707 1839 43741
rect 134855 43707 134889 43741
rect 1805 43371 1839 43405
rect 134855 43371 134889 43405
rect 1805 43035 1839 43069
rect 134855 43035 134889 43069
rect 1805 42699 1839 42733
rect 134855 42699 134889 42733
rect 1805 42363 1839 42397
rect 134855 42363 134889 42397
rect 1805 42027 1839 42061
rect 134855 42027 134889 42061
rect 1805 41691 1839 41725
rect 134855 41691 134889 41725
rect 1805 41355 1839 41389
rect 134855 41355 134889 41389
rect 1805 41019 1839 41053
rect 134855 41019 134889 41053
rect 1805 40683 1839 40717
rect 134855 40683 134889 40717
rect 1805 40347 1839 40381
rect 134855 40347 134889 40381
rect 1805 40011 1839 40045
rect 134855 40011 134889 40045
rect 1805 39675 1839 39709
rect 134855 39675 134889 39709
rect 1805 39339 1839 39373
rect 134855 39339 134889 39373
rect 1805 39003 1839 39037
rect 134855 39003 134889 39037
rect 1805 38667 1839 38701
rect 134855 38667 134889 38701
rect 1805 38331 1839 38365
rect 134855 38331 134889 38365
rect 1805 37995 1839 38029
rect 134855 37995 134889 38029
rect 1805 37659 1839 37693
rect 134855 37659 134889 37693
rect 1805 37323 1839 37357
rect 134855 37323 134889 37357
rect 1805 36987 1839 37021
rect 134855 36987 134889 37021
rect 1805 36651 1839 36685
rect 134855 36651 134889 36685
rect 1805 36315 1839 36349
rect 134855 36315 134889 36349
rect 1805 35979 1839 36013
rect 134855 35979 134889 36013
rect 1805 35643 1839 35677
rect 134855 35643 134889 35677
rect 1805 35307 1839 35341
rect 134855 35307 134889 35341
rect 1805 34971 1839 35005
rect 134855 34971 134889 35005
rect 1805 34635 1839 34669
rect 134855 34635 134889 34669
rect 1805 34299 1839 34333
rect 134855 34299 134889 34333
rect 1805 33963 1839 33997
rect 134855 33963 134889 33997
rect 1805 33627 1839 33661
rect 134855 33627 134889 33661
rect 1805 33291 1839 33325
rect 134855 33291 134889 33325
rect 1805 32955 1839 32989
rect 134855 32955 134889 32989
rect 1805 32619 1839 32653
rect 134855 32619 134889 32653
rect 1805 32283 1839 32317
rect 134855 32283 134889 32317
rect 1805 31947 1839 31981
rect 134855 31947 134889 31981
rect 1805 31611 1839 31645
rect 134855 31611 134889 31645
rect 1805 31275 1839 31309
rect 134855 31275 134889 31309
rect 1805 30939 1839 30973
rect 134855 30939 134889 30973
rect 1805 30603 1839 30637
rect 134855 30603 134889 30637
rect 1805 30267 1839 30301
rect 134855 30267 134889 30301
rect 1805 29931 1839 29965
rect 134855 29931 134889 29965
rect 1805 29595 1839 29629
rect 134855 29595 134889 29629
rect 1805 29259 1839 29293
rect 134855 29259 134889 29293
rect 1805 28923 1839 28957
rect 134855 28923 134889 28957
rect 1805 28587 1839 28621
rect 134855 28587 134889 28621
rect 1805 28251 1839 28285
rect 134855 28251 134889 28285
rect 1805 27915 1839 27949
rect 134855 27915 134889 27949
rect 1805 27579 1839 27613
rect 134855 27579 134889 27613
rect 1805 27243 1839 27277
rect 134855 27243 134889 27277
rect 1805 26907 1839 26941
rect 134855 26907 134889 26941
rect 1805 26571 1839 26605
rect 134855 26571 134889 26605
rect 1805 26235 1839 26269
rect 134855 26235 134889 26269
rect 1805 25899 1839 25933
rect 134855 25899 134889 25933
rect 1805 25563 1839 25597
rect 134855 25563 134889 25597
rect 1805 25227 1839 25261
rect 134855 25227 134889 25261
rect 1805 24891 1839 24925
rect 134855 24891 134889 24925
rect 1805 24555 1839 24589
rect 134855 24555 134889 24589
rect 1805 24219 1839 24253
rect 134855 24219 134889 24253
rect 1805 23883 1839 23917
rect 134855 23883 134889 23917
rect 1805 23547 1839 23581
rect 134855 23547 134889 23581
rect 1805 23211 1839 23245
rect 134855 23211 134889 23245
rect 1805 22875 1839 22909
rect 134855 22875 134889 22909
rect 1805 22539 1839 22573
rect 134855 22539 134889 22573
rect 1805 22203 1839 22237
rect 134855 22203 134889 22237
rect 1805 21867 1839 21901
rect 134855 21867 134889 21901
rect 1805 21531 1839 21565
rect 134855 21531 134889 21565
rect 1805 21195 1839 21229
rect 134855 21195 134889 21229
rect 1805 20859 1839 20893
rect 134855 20859 134889 20893
rect 1805 20523 1839 20557
rect 134855 20523 134889 20557
rect 1805 20187 1839 20221
rect 134855 20187 134889 20221
rect 1805 19851 1839 19885
rect 134855 19851 134889 19885
rect 1805 19515 1839 19549
rect 134855 19515 134889 19549
rect 1805 19179 1839 19213
rect 134855 19179 134889 19213
rect 1805 18843 1839 18877
rect 134855 18843 134889 18877
rect 1805 18507 1839 18541
rect 134855 18507 134889 18541
rect 1805 18171 1839 18205
rect 134855 18171 134889 18205
rect 1805 17835 1839 17869
rect 134855 17835 134889 17869
rect 1805 17499 1839 17533
rect 134855 17499 134889 17533
rect 1805 17163 1839 17197
rect 134855 17163 134889 17197
rect 1805 16827 1839 16861
rect 134855 16827 134889 16861
rect 1805 16491 1839 16525
rect 134855 16491 134889 16525
rect 1805 16155 1839 16189
rect 134855 16155 134889 16189
rect 1805 15819 1839 15853
rect 134855 15819 134889 15853
rect 1805 15483 1839 15517
rect 134855 15483 134889 15517
rect 1805 15147 1839 15181
rect 134855 15147 134889 15181
rect 1805 14811 1839 14845
rect 134855 14811 134889 14845
rect 1805 14475 1839 14509
rect 134855 14475 134889 14509
rect 1805 14139 1839 14173
rect 134855 14139 134889 14173
rect 1805 13803 1839 13837
rect 134855 13803 134889 13837
rect 1805 13467 1839 13501
rect 134855 13467 134889 13501
rect 1805 13131 1839 13165
rect 134855 13131 134889 13165
rect 1805 12795 1839 12829
rect 134855 12795 134889 12829
rect 1805 12459 1839 12493
rect 134855 12459 134889 12493
rect 1805 12123 1839 12157
rect 134855 12123 134889 12157
rect 1805 11787 1839 11821
rect 134855 11787 134889 11821
rect 1805 11451 1839 11485
rect 134855 11451 134889 11485
rect 1805 11115 1839 11149
rect 134855 11115 134889 11149
rect 1805 10779 1839 10813
rect 134855 10779 134889 10813
rect 1805 10443 1839 10477
rect 134855 10443 134889 10477
rect 1805 10107 1839 10141
rect 134855 10107 134889 10141
rect 1805 9771 1839 9805
rect 134855 9771 134889 9805
rect 1805 9435 1839 9469
rect 134855 9435 134889 9469
rect 1805 9099 1839 9133
rect 134855 9099 134889 9133
rect 1805 8763 1839 8797
rect 134855 8763 134889 8797
rect 1805 8427 1839 8461
rect 134855 8427 134889 8461
rect 1805 8091 1839 8125
rect 134855 8091 134889 8125
rect 1805 7755 1839 7789
rect 134855 7755 134889 7789
rect 1805 7419 1839 7453
rect 134855 7419 134889 7453
rect 1805 7083 1839 7117
rect 134855 7083 134889 7117
rect 1805 6747 1839 6781
rect 134855 6747 134889 6781
rect 1805 6411 1839 6445
rect 134855 6411 134889 6445
rect 1805 6075 1839 6109
rect 134855 6075 134889 6109
rect 1805 5739 1839 5773
rect 134855 5739 134889 5773
rect 1805 5403 1839 5437
rect 134855 5403 134889 5437
rect 1805 5067 1839 5101
rect 134855 5067 134889 5101
rect 1805 4731 1839 4765
rect 134855 4731 134889 4765
rect 1805 4395 1839 4429
rect 134855 4395 134889 4429
rect 1805 4059 1839 4093
rect 134855 4059 134889 4093
rect 1805 3723 1839 3757
rect 134855 3723 134889 3757
rect 1805 3387 1839 3421
rect 134855 3387 134889 3421
rect 1805 3051 1839 3085
rect 134855 3051 134889 3085
rect 1805 2715 1839 2749
rect 134855 2715 134889 2749
rect 1805 2379 1839 2413
rect 134855 2379 134889 2413
rect 1805 2043 1839 2077
rect 134855 2043 134889 2077
rect 2141 1707 2175 1741
rect 2477 1707 2511 1741
rect 2813 1707 2847 1741
rect 3149 1707 3183 1741
rect 3485 1707 3519 1741
rect 3821 1707 3855 1741
rect 4157 1707 4191 1741
rect 4493 1707 4527 1741
rect 4829 1707 4863 1741
rect 5165 1707 5199 1741
rect 5501 1707 5535 1741
rect 5837 1707 5871 1741
rect 6173 1707 6207 1741
rect 6509 1707 6543 1741
rect 6845 1707 6879 1741
rect 7181 1707 7215 1741
rect 7517 1707 7551 1741
rect 7853 1707 7887 1741
rect 8189 1707 8223 1741
rect 8525 1707 8559 1741
rect 8861 1707 8895 1741
rect 9197 1707 9231 1741
rect 9533 1707 9567 1741
rect 9869 1707 9903 1741
rect 10205 1707 10239 1741
rect 10541 1707 10575 1741
rect 10877 1707 10911 1741
rect 11213 1707 11247 1741
rect 11549 1707 11583 1741
rect 11885 1707 11919 1741
rect 12221 1707 12255 1741
rect 12557 1707 12591 1741
rect 12893 1707 12927 1741
rect 13229 1707 13263 1741
rect 13565 1707 13599 1741
rect 13901 1707 13935 1741
rect 14237 1707 14271 1741
rect 14573 1707 14607 1741
rect 14909 1707 14943 1741
rect 15245 1707 15279 1741
rect 15581 1707 15615 1741
rect 15917 1707 15951 1741
rect 16253 1707 16287 1741
rect 16589 1707 16623 1741
rect 16925 1707 16959 1741
rect 17261 1707 17295 1741
rect 17597 1707 17631 1741
rect 17933 1707 17967 1741
rect 18269 1707 18303 1741
rect 18605 1707 18639 1741
rect 18941 1707 18975 1741
rect 19277 1707 19311 1741
rect 19613 1707 19647 1741
rect 19949 1707 19983 1741
rect 20285 1707 20319 1741
rect 20621 1707 20655 1741
rect 20957 1707 20991 1741
rect 21293 1707 21327 1741
rect 21629 1707 21663 1741
rect 21965 1707 21999 1741
rect 22301 1707 22335 1741
rect 22637 1707 22671 1741
rect 22973 1707 23007 1741
rect 23309 1707 23343 1741
rect 23645 1707 23679 1741
rect 23981 1707 24015 1741
rect 24317 1707 24351 1741
rect 24653 1707 24687 1741
rect 24989 1707 25023 1741
rect 25325 1707 25359 1741
rect 25661 1707 25695 1741
rect 25997 1707 26031 1741
rect 26333 1707 26367 1741
rect 26669 1707 26703 1741
rect 27005 1707 27039 1741
rect 27341 1707 27375 1741
rect 27677 1707 27711 1741
rect 28013 1707 28047 1741
rect 28349 1707 28383 1741
rect 28685 1707 28719 1741
rect 29021 1707 29055 1741
rect 29357 1707 29391 1741
rect 29693 1707 29727 1741
rect 30029 1707 30063 1741
rect 30365 1707 30399 1741
rect 30701 1707 30735 1741
rect 31037 1707 31071 1741
rect 31373 1707 31407 1741
rect 31709 1707 31743 1741
rect 32045 1707 32079 1741
rect 32381 1707 32415 1741
rect 32717 1707 32751 1741
rect 33053 1707 33087 1741
rect 33389 1707 33423 1741
rect 33725 1707 33759 1741
rect 34061 1707 34095 1741
rect 34397 1707 34431 1741
rect 34733 1707 34767 1741
rect 35069 1707 35103 1741
rect 35405 1707 35439 1741
rect 35741 1707 35775 1741
rect 36077 1707 36111 1741
rect 36413 1707 36447 1741
rect 36749 1707 36783 1741
rect 37085 1707 37119 1741
rect 37421 1707 37455 1741
rect 37757 1707 37791 1741
rect 38093 1707 38127 1741
rect 38429 1707 38463 1741
rect 38765 1707 38799 1741
rect 39101 1707 39135 1741
rect 39437 1707 39471 1741
rect 39773 1707 39807 1741
rect 40109 1707 40143 1741
rect 40445 1707 40479 1741
rect 40781 1707 40815 1741
rect 41117 1707 41151 1741
rect 41453 1707 41487 1741
rect 41789 1707 41823 1741
rect 42125 1707 42159 1741
rect 42461 1707 42495 1741
rect 42797 1707 42831 1741
rect 43133 1707 43167 1741
rect 43469 1707 43503 1741
rect 43805 1707 43839 1741
rect 44141 1707 44175 1741
rect 44477 1707 44511 1741
rect 44813 1707 44847 1741
rect 45149 1707 45183 1741
rect 45485 1707 45519 1741
rect 45821 1707 45855 1741
rect 46157 1707 46191 1741
rect 46493 1707 46527 1741
rect 46829 1707 46863 1741
rect 47165 1707 47199 1741
rect 47501 1707 47535 1741
rect 47837 1707 47871 1741
rect 48173 1707 48207 1741
rect 48509 1707 48543 1741
rect 48845 1707 48879 1741
rect 49181 1707 49215 1741
rect 49517 1707 49551 1741
rect 49853 1707 49887 1741
rect 50189 1707 50223 1741
rect 50525 1707 50559 1741
rect 50861 1707 50895 1741
rect 51197 1707 51231 1741
rect 51533 1707 51567 1741
rect 51869 1707 51903 1741
rect 52205 1707 52239 1741
rect 52541 1707 52575 1741
rect 52877 1707 52911 1741
rect 53213 1707 53247 1741
rect 53549 1707 53583 1741
rect 53885 1707 53919 1741
rect 54221 1707 54255 1741
rect 54557 1707 54591 1741
rect 54893 1707 54927 1741
rect 55229 1707 55263 1741
rect 55565 1707 55599 1741
rect 55901 1707 55935 1741
rect 56237 1707 56271 1741
rect 56573 1707 56607 1741
rect 56909 1707 56943 1741
rect 57245 1707 57279 1741
rect 57581 1707 57615 1741
rect 57917 1707 57951 1741
rect 58253 1707 58287 1741
rect 58589 1707 58623 1741
rect 58925 1707 58959 1741
rect 59261 1707 59295 1741
rect 59597 1707 59631 1741
rect 59933 1707 59967 1741
rect 60269 1707 60303 1741
rect 60605 1707 60639 1741
rect 60941 1707 60975 1741
rect 61277 1707 61311 1741
rect 61613 1707 61647 1741
rect 61949 1707 61983 1741
rect 62285 1707 62319 1741
rect 62621 1707 62655 1741
rect 62957 1707 62991 1741
rect 63293 1707 63327 1741
rect 63629 1707 63663 1741
rect 63965 1707 63999 1741
rect 64301 1707 64335 1741
rect 64637 1707 64671 1741
rect 64973 1707 65007 1741
rect 65309 1707 65343 1741
rect 65645 1707 65679 1741
rect 65981 1707 66015 1741
rect 66317 1707 66351 1741
rect 66653 1707 66687 1741
rect 66989 1707 67023 1741
rect 67325 1707 67359 1741
rect 67661 1707 67695 1741
rect 67997 1707 68031 1741
rect 68333 1707 68367 1741
rect 68669 1707 68703 1741
rect 69005 1707 69039 1741
rect 69341 1707 69375 1741
rect 69677 1707 69711 1741
rect 70013 1707 70047 1741
rect 70349 1707 70383 1741
rect 70685 1707 70719 1741
rect 71021 1707 71055 1741
rect 71357 1707 71391 1741
rect 71693 1707 71727 1741
rect 72029 1707 72063 1741
rect 72365 1707 72399 1741
rect 72701 1707 72735 1741
rect 73037 1707 73071 1741
rect 73373 1707 73407 1741
rect 73709 1707 73743 1741
rect 74045 1707 74079 1741
rect 74381 1707 74415 1741
rect 74717 1707 74751 1741
rect 75053 1707 75087 1741
rect 75389 1707 75423 1741
rect 75725 1707 75759 1741
rect 76061 1707 76095 1741
rect 76397 1707 76431 1741
rect 76733 1707 76767 1741
rect 77069 1707 77103 1741
rect 77405 1707 77439 1741
rect 77741 1707 77775 1741
rect 78077 1707 78111 1741
rect 78413 1707 78447 1741
rect 78749 1707 78783 1741
rect 79085 1707 79119 1741
rect 79421 1707 79455 1741
rect 79757 1707 79791 1741
rect 80093 1707 80127 1741
rect 80429 1707 80463 1741
rect 80765 1707 80799 1741
rect 81101 1707 81135 1741
rect 81437 1707 81471 1741
rect 81773 1707 81807 1741
rect 82109 1707 82143 1741
rect 82445 1707 82479 1741
rect 82781 1707 82815 1741
rect 83117 1707 83151 1741
rect 83453 1707 83487 1741
rect 83789 1707 83823 1741
rect 84125 1707 84159 1741
rect 84461 1707 84495 1741
rect 84797 1707 84831 1741
rect 85133 1707 85167 1741
rect 85469 1707 85503 1741
rect 85805 1707 85839 1741
rect 86141 1707 86175 1741
rect 86477 1707 86511 1741
rect 86813 1707 86847 1741
rect 87149 1707 87183 1741
rect 87485 1707 87519 1741
rect 87821 1707 87855 1741
rect 88157 1707 88191 1741
rect 88493 1707 88527 1741
rect 88829 1707 88863 1741
rect 89165 1707 89199 1741
rect 89501 1707 89535 1741
rect 89837 1707 89871 1741
rect 90173 1707 90207 1741
rect 90509 1707 90543 1741
rect 90845 1707 90879 1741
rect 91181 1707 91215 1741
rect 91517 1707 91551 1741
rect 91853 1707 91887 1741
rect 92189 1707 92223 1741
rect 92525 1707 92559 1741
rect 92861 1707 92895 1741
rect 93197 1707 93231 1741
rect 93533 1707 93567 1741
rect 93869 1707 93903 1741
rect 94205 1707 94239 1741
rect 94541 1707 94575 1741
rect 94877 1707 94911 1741
rect 95213 1707 95247 1741
rect 95549 1707 95583 1741
rect 95885 1707 95919 1741
rect 96221 1707 96255 1741
rect 96557 1707 96591 1741
rect 96893 1707 96927 1741
rect 97229 1707 97263 1741
rect 97565 1707 97599 1741
rect 97901 1707 97935 1741
rect 98237 1707 98271 1741
rect 98573 1707 98607 1741
rect 98909 1707 98943 1741
rect 99245 1707 99279 1741
rect 99581 1707 99615 1741
rect 99917 1707 99951 1741
rect 100253 1707 100287 1741
rect 100589 1707 100623 1741
rect 100925 1707 100959 1741
rect 101261 1707 101295 1741
rect 101597 1707 101631 1741
rect 101933 1707 101967 1741
rect 102269 1707 102303 1741
rect 102605 1707 102639 1741
rect 102941 1707 102975 1741
rect 103277 1707 103311 1741
rect 103613 1707 103647 1741
rect 103949 1707 103983 1741
rect 104285 1707 104319 1741
rect 104621 1707 104655 1741
rect 104957 1707 104991 1741
rect 105293 1707 105327 1741
rect 105629 1707 105663 1741
rect 105965 1707 105999 1741
rect 106301 1707 106335 1741
rect 106637 1707 106671 1741
rect 106973 1707 107007 1741
rect 107309 1707 107343 1741
rect 107645 1707 107679 1741
rect 107981 1707 108015 1741
rect 108317 1707 108351 1741
rect 108653 1707 108687 1741
rect 108989 1707 109023 1741
rect 109325 1707 109359 1741
rect 109661 1707 109695 1741
rect 109997 1707 110031 1741
rect 110333 1707 110367 1741
rect 110669 1707 110703 1741
rect 111005 1707 111039 1741
rect 111341 1707 111375 1741
rect 111677 1707 111711 1741
rect 112013 1707 112047 1741
rect 112349 1707 112383 1741
rect 112685 1707 112719 1741
rect 113021 1707 113055 1741
rect 113357 1707 113391 1741
rect 113693 1707 113727 1741
rect 114029 1707 114063 1741
rect 114365 1707 114399 1741
rect 114701 1707 114735 1741
rect 115037 1707 115071 1741
rect 115373 1707 115407 1741
rect 115709 1707 115743 1741
rect 116045 1707 116079 1741
rect 116381 1707 116415 1741
rect 116717 1707 116751 1741
rect 117053 1707 117087 1741
rect 117389 1707 117423 1741
rect 117725 1707 117759 1741
rect 118061 1707 118095 1741
rect 118397 1707 118431 1741
rect 118733 1707 118767 1741
rect 119069 1707 119103 1741
rect 119405 1707 119439 1741
rect 119741 1707 119775 1741
rect 120077 1707 120111 1741
rect 120413 1707 120447 1741
rect 120749 1707 120783 1741
rect 121085 1707 121119 1741
rect 121421 1707 121455 1741
rect 121757 1707 121791 1741
rect 122093 1707 122127 1741
rect 122429 1707 122463 1741
rect 122765 1707 122799 1741
rect 123101 1707 123135 1741
rect 123437 1707 123471 1741
rect 123773 1707 123807 1741
rect 124109 1707 124143 1741
rect 124445 1707 124479 1741
rect 124781 1707 124815 1741
rect 125117 1707 125151 1741
rect 125453 1707 125487 1741
rect 125789 1707 125823 1741
rect 126125 1707 126159 1741
rect 126461 1707 126495 1741
rect 126797 1707 126831 1741
rect 127133 1707 127167 1741
rect 127469 1707 127503 1741
rect 127805 1707 127839 1741
rect 128141 1707 128175 1741
rect 128477 1707 128511 1741
rect 128813 1707 128847 1741
rect 129149 1707 129183 1741
rect 129485 1707 129519 1741
rect 129821 1707 129855 1741
rect 130157 1707 130191 1741
rect 130493 1707 130527 1741
rect 130829 1707 130863 1741
rect 131165 1707 131199 1741
rect 131501 1707 131535 1741
rect 131837 1707 131871 1741
rect 132173 1707 132207 1741
rect 132509 1707 132543 1741
rect 132845 1707 132879 1741
rect 133181 1707 133215 1741
rect 133517 1707 133551 1741
rect 133853 1707 133887 1741
rect 134189 1707 134223 1741
<< metal1 >>
rect 1710 81499 134984 81585
rect 1710 81447 2132 81499
rect 2184 81490 3812 81499
rect 3864 81490 5492 81499
rect 5544 81490 7172 81499
rect 7224 81490 8852 81499
rect 8904 81490 10532 81499
rect 10584 81490 12212 81499
rect 12264 81490 13892 81499
rect 13944 81490 15572 81499
rect 15624 81490 17252 81499
rect 17304 81490 18932 81499
rect 18984 81490 20612 81499
rect 20664 81490 22292 81499
rect 22344 81490 23972 81499
rect 24024 81490 25652 81499
rect 25704 81490 27332 81499
rect 27384 81490 29012 81499
rect 29064 81490 30692 81499
rect 30744 81490 32372 81499
rect 32424 81490 34052 81499
rect 34104 81490 35732 81499
rect 35784 81490 37412 81499
rect 37464 81490 39092 81499
rect 39144 81490 40772 81499
rect 40824 81490 42452 81499
rect 42504 81490 44132 81499
rect 44184 81490 45812 81499
rect 45864 81490 47492 81499
rect 47544 81490 49172 81499
rect 49224 81490 50852 81499
rect 50904 81490 52532 81499
rect 52584 81490 54212 81499
rect 54264 81490 55892 81499
rect 55944 81490 57572 81499
rect 57624 81490 59252 81499
rect 59304 81490 60932 81499
rect 60984 81490 62612 81499
rect 62664 81490 64292 81499
rect 64344 81490 65972 81499
rect 66024 81490 67652 81499
rect 67704 81490 69332 81499
rect 69384 81490 71012 81499
rect 71064 81490 72692 81499
rect 72744 81490 74372 81499
rect 74424 81490 76052 81499
rect 76104 81490 77732 81499
rect 77784 81490 79412 81499
rect 79464 81490 81092 81499
rect 81144 81490 82772 81499
rect 82824 81490 84452 81499
rect 84504 81490 86132 81499
rect 86184 81490 87812 81499
rect 87864 81490 89492 81499
rect 89544 81490 91172 81499
rect 91224 81490 92852 81499
rect 92904 81490 94532 81499
rect 94584 81490 96212 81499
rect 96264 81490 97892 81499
rect 97944 81490 99572 81499
rect 99624 81490 101252 81499
rect 101304 81490 102932 81499
rect 102984 81490 104612 81499
rect 104664 81490 106292 81499
rect 106344 81490 107972 81499
rect 108024 81490 109652 81499
rect 109704 81490 111332 81499
rect 111384 81490 113012 81499
rect 113064 81490 114692 81499
rect 114744 81490 116372 81499
rect 116424 81490 118052 81499
rect 118104 81490 119732 81499
rect 119784 81490 121412 81499
rect 121464 81490 123092 81499
rect 123144 81490 124772 81499
rect 124824 81490 126452 81499
rect 126504 81490 128132 81499
rect 128184 81490 129812 81499
rect 129864 81490 131492 81499
rect 131544 81490 133172 81499
rect 133224 81490 134984 81499
rect 2184 81456 2477 81490
rect 2511 81456 2813 81490
rect 2847 81456 3149 81490
rect 3183 81456 3485 81490
rect 3519 81456 3812 81490
rect 3864 81456 4157 81490
rect 4191 81456 4493 81490
rect 4527 81456 4829 81490
rect 4863 81456 5165 81490
rect 5199 81456 5492 81490
rect 5544 81456 5837 81490
rect 5871 81456 6173 81490
rect 6207 81456 6509 81490
rect 6543 81456 6845 81490
rect 6879 81456 7172 81490
rect 7224 81456 7517 81490
rect 7551 81456 7853 81490
rect 7887 81456 8189 81490
rect 8223 81456 8525 81490
rect 8559 81456 8852 81490
rect 8904 81456 9197 81490
rect 9231 81456 9533 81490
rect 9567 81456 9869 81490
rect 9903 81456 10205 81490
rect 10239 81456 10532 81490
rect 10584 81456 10877 81490
rect 10911 81456 11213 81490
rect 11247 81456 11549 81490
rect 11583 81456 11885 81490
rect 11919 81456 12212 81490
rect 12264 81456 12557 81490
rect 12591 81456 12893 81490
rect 12927 81456 13229 81490
rect 13263 81456 13565 81490
rect 13599 81456 13892 81490
rect 13944 81456 14237 81490
rect 14271 81456 14573 81490
rect 14607 81456 14909 81490
rect 14943 81456 15245 81490
rect 15279 81456 15572 81490
rect 15624 81456 15917 81490
rect 15951 81456 16253 81490
rect 16287 81456 16589 81490
rect 16623 81456 16925 81490
rect 16959 81456 17252 81490
rect 17304 81456 17597 81490
rect 17631 81456 17933 81490
rect 17967 81456 18269 81490
rect 18303 81456 18605 81490
rect 18639 81456 18932 81490
rect 18984 81456 19277 81490
rect 19311 81456 19613 81490
rect 19647 81456 19949 81490
rect 19983 81456 20285 81490
rect 20319 81456 20612 81490
rect 20664 81456 20957 81490
rect 20991 81456 21293 81490
rect 21327 81456 21629 81490
rect 21663 81456 21965 81490
rect 21999 81456 22292 81490
rect 22344 81456 22637 81490
rect 22671 81456 22973 81490
rect 23007 81456 23309 81490
rect 23343 81456 23645 81490
rect 23679 81456 23972 81490
rect 24024 81456 24317 81490
rect 24351 81456 24653 81490
rect 24687 81456 24989 81490
rect 25023 81456 25325 81490
rect 25359 81456 25652 81490
rect 25704 81456 25997 81490
rect 26031 81456 26333 81490
rect 26367 81456 26669 81490
rect 26703 81456 27005 81490
rect 27039 81456 27332 81490
rect 27384 81456 27677 81490
rect 27711 81456 28013 81490
rect 28047 81456 28349 81490
rect 28383 81456 28685 81490
rect 28719 81456 29012 81490
rect 29064 81456 29357 81490
rect 29391 81456 29693 81490
rect 29727 81456 30029 81490
rect 30063 81456 30365 81490
rect 30399 81456 30692 81490
rect 30744 81456 31037 81490
rect 31071 81456 31373 81490
rect 31407 81456 31709 81490
rect 31743 81456 32045 81490
rect 32079 81456 32372 81490
rect 32424 81456 32717 81490
rect 32751 81456 33053 81490
rect 33087 81456 33389 81490
rect 33423 81456 33725 81490
rect 33759 81456 34052 81490
rect 34104 81456 34397 81490
rect 34431 81456 34733 81490
rect 34767 81456 35069 81490
rect 35103 81456 35405 81490
rect 35439 81456 35732 81490
rect 35784 81456 36077 81490
rect 36111 81456 36413 81490
rect 36447 81456 36749 81490
rect 36783 81456 37085 81490
rect 37119 81456 37412 81490
rect 37464 81456 37757 81490
rect 37791 81456 38093 81490
rect 38127 81456 38429 81490
rect 38463 81456 38765 81490
rect 38799 81456 39092 81490
rect 39144 81456 39437 81490
rect 39471 81456 39773 81490
rect 39807 81456 40109 81490
rect 40143 81456 40445 81490
rect 40479 81456 40772 81490
rect 40824 81456 41117 81490
rect 41151 81456 41453 81490
rect 41487 81456 41789 81490
rect 41823 81456 42125 81490
rect 42159 81456 42452 81490
rect 42504 81456 42797 81490
rect 42831 81456 43133 81490
rect 43167 81456 43469 81490
rect 43503 81456 43805 81490
rect 43839 81456 44132 81490
rect 44184 81456 44477 81490
rect 44511 81456 44813 81490
rect 44847 81456 45149 81490
rect 45183 81456 45485 81490
rect 45519 81456 45812 81490
rect 45864 81456 46157 81490
rect 46191 81456 46493 81490
rect 46527 81456 46829 81490
rect 46863 81456 47165 81490
rect 47199 81456 47492 81490
rect 47544 81456 47837 81490
rect 47871 81456 48173 81490
rect 48207 81456 48509 81490
rect 48543 81456 48845 81490
rect 48879 81456 49172 81490
rect 49224 81456 49517 81490
rect 49551 81456 49853 81490
rect 49887 81456 50189 81490
rect 50223 81456 50525 81490
rect 50559 81456 50852 81490
rect 50904 81456 51197 81490
rect 51231 81456 51533 81490
rect 51567 81456 51869 81490
rect 51903 81456 52205 81490
rect 52239 81456 52532 81490
rect 52584 81456 52877 81490
rect 52911 81456 53213 81490
rect 53247 81456 53549 81490
rect 53583 81456 53885 81490
rect 53919 81456 54212 81490
rect 54264 81456 54557 81490
rect 54591 81456 54893 81490
rect 54927 81456 55229 81490
rect 55263 81456 55565 81490
rect 55599 81456 55892 81490
rect 55944 81456 56237 81490
rect 56271 81456 56573 81490
rect 56607 81456 56909 81490
rect 56943 81456 57245 81490
rect 57279 81456 57572 81490
rect 57624 81456 57917 81490
rect 57951 81456 58253 81490
rect 58287 81456 58589 81490
rect 58623 81456 58925 81490
rect 58959 81456 59252 81490
rect 59304 81456 59597 81490
rect 59631 81456 59933 81490
rect 59967 81456 60269 81490
rect 60303 81456 60605 81490
rect 60639 81456 60932 81490
rect 60984 81456 61277 81490
rect 61311 81456 61613 81490
rect 61647 81456 61949 81490
rect 61983 81456 62285 81490
rect 62319 81456 62612 81490
rect 62664 81456 62957 81490
rect 62991 81456 63293 81490
rect 63327 81456 63629 81490
rect 63663 81456 63965 81490
rect 63999 81456 64292 81490
rect 64344 81456 64637 81490
rect 64671 81456 64973 81490
rect 65007 81456 65309 81490
rect 65343 81456 65645 81490
rect 65679 81456 65972 81490
rect 66024 81456 66317 81490
rect 66351 81456 66653 81490
rect 66687 81456 66989 81490
rect 67023 81456 67325 81490
rect 67359 81456 67652 81490
rect 67704 81456 67997 81490
rect 68031 81456 68333 81490
rect 68367 81456 68669 81490
rect 68703 81456 69005 81490
rect 69039 81456 69332 81490
rect 69384 81456 69677 81490
rect 69711 81456 70013 81490
rect 70047 81456 70349 81490
rect 70383 81456 70685 81490
rect 70719 81456 71012 81490
rect 71064 81456 71357 81490
rect 71391 81456 71693 81490
rect 71727 81456 72029 81490
rect 72063 81456 72365 81490
rect 72399 81456 72692 81490
rect 72744 81456 73037 81490
rect 73071 81456 73373 81490
rect 73407 81456 73709 81490
rect 73743 81456 74045 81490
rect 74079 81456 74372 81490
rect 74424 81456 74717 81490
rect 74751 81456 75053 81490
rect 75087 81456 75389 81490
rect 75423 81456 75725 81490
rect 75759 81456 76052 81490
rect 76104 81456 76397 81490
rect 76431 81456 76733 81490
rect 76767 81456 77069 81490
rect 77103 81456 77405 81490
rect 77439 81456 77732 81490
rect 77784 81456 78077 81490
rect 78111 81456 78413 81490
rect 78447 81456 78749 81490
rect 78783 81456 79085 81490
rect 79119 81456 79412 81490
rect 79464 81456 79757 81490
rect 79791 81456 80093 81490
rect 80127 81456 80429 81490
rect 80463 81456 80765 81490
rect 80799 81456 81092 81490
rect 81144 81456 81437 81490
rect 81471 81456 81773 81490
rect 81807 81456 82109 81490
rect 82143 81456 82445 81490
rect 82479 81456 82772 81490
rect 82824 81456 83117 81490
rect 83151 81456 83453 81490
rect 83487 81456 83789 81490
rect 83823 81456 84125 81490
rect 84159 81456 84452 81490
rect 84504 81456 84797 81490
rect 84831 81456 85133 81490
rect 85167 81456 85469 81490
rect 85503 81456 85805 81490
rect 85839 81456 86132 81490
rect 86184 81456 86477 81490
rect 86511 81456 86813 81490
rect 86847 81456 87149 81490
rect 87183 81456 87485 81490
rect 87519 81456 87812 81490
rect 87864 81456 88157 81490
rect 88191 81456 88493 81490
rect 88527 81456 88829 81490
rect 88863 81456 89165 81490
rect 89199 81456 89492 81490
rect 89544 81456 89837 81490
rect 89871 81456 90173 81490
rect 90207 81456 90509 81490
rect 90543 81456 90845 81490
rect 90879 81456 91172 81490
rect 91224 81456 91517 81490
rect 91551 81456 91853 81490
rect 91887 81456 92189 81490
rect 92223 81456 92525 81490
rect 92559 81456 92852 81490
rect 92904 81456 93197 81490
rect 93231 81456 93533 81490
rect 93567 81456 93869 81490
rect 93903 81456 94205 81490
rect 94239 81456 94532 81490
rect 94584 81456 94877 81490
rect 94911 81456 95213 81490
rect 95247 81456 95549 81490
rect 95583 81456 95885 81490
rect 95919 81456 96212 81490
rect 96264 81456 96557 81490
rect 96591 81456 96893 81490
rect 96927 81456 97229 81490
rect 97263 81456 97565 81490
rect 97599 81456 97892 81490
rect 97944 81456 98237 81490
rect 98271 81456 98573 81490
rect 98607 81456 98909 81490
rect 98943 81456 99245 81490
rect 99279 81456 99572 81490
rect 99624 81456 99917 81490
rect 99951 81456 100253 81490
rect 100287 81456 100589 81490
rect 100623 81456 100925 81490
rect 100959 81456 101252 81490
rect 101304 81456 101597 81490
rect 101631 81456 101933 81490
rect 101967 81456 102269 81490
rect 102303 81456 102605 81490
rect 102639 81456 102932 81490
rect 102984 81456 103277 81490
rect 103311 81456 103613 81490
rect 103647 81456 103949 81490
rect 103983 81456 104285 81490
rect 104319 81456 104612 81490
rect 104664 81456 104957 81490
rect 104991 81456 105293 81490
rect 105327 81456 105629 81490
rect 105663 81456 105965 81490
rect 105999 81456 106292 81490
rect 106344 81456 106637 81490
rect 106671 81456 106973 81490
rect 107007 81456 107309 81490
rect 107343 81456 107645 81490
rect 107679 81456 107972 81490
rect 108024 81456 108317 81490
rect 108351 81456 108653 81490
rect 108687 81456 108989 81490
rect 109023 81456 109325 81490
rect 109359 81456 109652 81490
rect 109704 81456 109997 81490
rect 110031 81456 110333 81490
rect 110367 81456 110669 81490
rect 110703 81456 111005 81490
rect 111039 81456 111332 81490
rect 111384 81456 111677 81490
rect 111711 81456 112013 81490
rect 112047 81456 112349 81490
rect 112383 81456 112685 81490
rect 112719 81456 113012 81490
rect 113064 81456 113357 81490
rect 113391 81456 113693 81490
rect 113727 81456 114029 81490
rect 114063 81456 114365 81490
rect 114399 81456 114692 81490
rect 114744 81456 115037 81490
rect 115071 81456 115373 81490
rect 115407 81456 115709 81490
rect 115743 81456 116045 81490
rect 116079 81456 116372 81490
rect 116424 81456 116717 81490
rect 116751 81456 117053 81490
rect 117087 81456 117389 81490
rect 117423 81456 117725 81490
rect 117759 81456 118052 81490
rect 118104 81456 118397 81490
rect 118431 81456 118733 81490
rect 118767 81456 119069 81490
rect 119103 81456 119405 81490
rect 119439 81456 119732 81490
rect 119784 81456 120077 81490
rect 120111 81456 120413 81490
rect 120447 81456 120749 81490
rect 120783 81456 121085 81490
rect 121119 81456 121412 81490
rect 121464 81456 121757 81490
rect 121791 81456 122093 81490
rect 122127 81456 122429 81490
rect 122463 81456 122765 81490
rect 122799 81456 123092 81490
rect 123144 81456 123437 81490
rect 123471 81456 123773 81490
rect 123807 81456 124109 81490
rect 124143 81456 124445 81490
rect 124479 81456 124772 81490
rect 124824 81456 125117 81490
rect 125151 81456 125453 81490
rect 125487 81456 125789 81490
rect 125823 81456 126125 81490
rect 126159 81456 126452 81490
rect 126504 81456 126797 81490
rect 126831 81456 127133 81490
rect 127167 81456 127469 81490
rect 127503 81456 127805 81490
rect 127839 81456 128132 81490
rect 128184 81456 128477 81490
rect 128511 81456 128813 81490
rect 128847 81456 129149 81490
rect 129183 81456 129485 81490
rect 129519 81456 129812 81490
rect 129864 81456 130157 81490
rect 130191 81456 130493 81490
rect 130527 81456 130829 81490
rect 130863 81456 131165 81490
rect 131199 81456 131492 81490
rect 131544 81456 131837 81490
rect 131871 81456 132173 81490
rect 132207 81456 132509 81490
rect 132543 81456 132845 81490
rect 132879 81456 133172 81490
rect 133224 81456 133517 81490
rect 133551 81456 133853 81490
rect 133887 81456 134189 81490
rect 134223 81456 134984 81490
rect 2184 81447 3812 81456
rect 3864 81447 5492 81456
rect 5544 81447 7172 81456
rect 7224 81447 8852 81456
rect 8904 81447 10532 81456
rect 10584 81447 12212 81456
rect 12264 81447 13892 81456
rect 13944 81447 15572 81456
rect 15624 81447 17252 81456
rect 17304 81447 18932 81456
rect 18984 81447 20612 81456
rect 20664 81447 22292 81456
rect 22344 81447 23972 81456
rect 24024 81447 25652 81456
rect 25704 81447 27332 81456
rect 27384 81447 29012 81456
rect 29064 81447 30692 81456
rect 30744 81447 32372 81456
rect 32424 81447 34052 81456
rect 34104 81447 35732 81456
rect 35784 81447 37412 81456
rect 37464 81447 39092 81456
rect 39144 81447 40772 81456
rect 40824 81447 42452 81456
rect 42504 81447 44132 81456
rect 44184 81447 45812 81456
rect 45864 81447 47492 81456
rect 47544 81447 49172 81456
rect 49224 81447 50852 81456
rect 50904 81447 52532 81456
rect 52584 81447 54212 81456
rect 54264 81447 55892 81456
rect 55944 81447 57572 81456
rect 57624 81447 59252 81456
rect 59304 81447 60932 81456
rect 60984 81447 62612 81456
rect 62664 81447 64292 81456
rect 64344 81447 65972 81456
rect 66024 81447 67652 81456
rect 67704 81447 69332 81456
rect 69384 81447 71012 81456
rect 71064 81447 72692 81456
rect 72744 81447 74372 81456
rect 74424 81447 76052 81456
rect 76104 81447 77732 81456
rect 77784 81447 79412 81456
rect 79464 81447 81092 81456
rect 81144 81447 82772 81456
rect 82824 81447 84452 81456
rect 84504 81447 86132 81456
rect 86184 81447 87812 81456
rect 87864 81447 89492 81456
rect 89544 81447 91172 81456
rect 91224 81447 92852 81456
rect 92904 81447 94532 81456
rect 94584 81447 96212 81456
rect 96264 81447 97892 81456
rect 97944 81447 99572 81456
rect 99624 81447 101252 81456
rect 101304 81447 102932 81456
rect 102984 81447 104612 81456
rect 104664 81447 106292 81456
rect 106344 81447 107972 81456
rect 108024 81447 109652 81456
rect 109704 81447 111332 81456
rect 111384 81447 113012 81456
rect 113064 81447 114692 81456
rect 114744 81447 116372 81456
rect 116424 81447 118052 81456
rect 118104 81447 119732 81456
rect 119784 81447 121412 81456
rect 121464 81447 123092 81456
rect 123144 81447 124772 81456
rect 124824 81447 126452 81456
rect 126504 81447 128132 81456
rect 128184 81447 129812 81456
rect 129864 81447 131492 81456
rect 131544 81447 133172 81456
rect 133224 81447 134984 81456
rect 1710 81361 134984 81447
rect 1790 80994 1796 81046
rect 1848 80994 1854 81046
rect 134840 80994 134846 81046
rect 134898 80994 134904 81046
rect 1790 80658 1796 80710
rect 1848 80658 1854 80710
rect 134840 80658 134846 80710
rect 134898 80658 134904 80710
rect 1790 80322 1796 80374
rect 1848 80322 1854 80374
rect 134840 80322 134846 80374
rect 134898 80322 134904 80374
rect 1790 79986 1796 80038
rect 1848 79986 1854 80038
rect 134840 79986 134846 80038
rect 134898 79986 134904 80038
rect 1790 79650 1796 79702
rect 1848 79650 1854 79702
rect 134840 79650 134846 79702
rect 134898 79650 134904 79702
rect 1790 79314 1796 79366
rect 1848 79314 1854 79366
rect 134840 79314 134846 79366
rect 134898 79314 134904 79366
rect 1790 78978 1796 79030
rect 1848 78978 1854 79030
rect 134840 78978 134846 79030
rect 134898 78978 134904 79030
rect 1790 78642 1796 78694
rect 1848 78642 1854 78694
rect 134840 78642 134846 78694
rect 134898 78642 134904 78694
rect 1790 78306 1796 78358
rect 1848 78306 1854 78358
rect 134840 78306 134846 78358
rect 134898 78306 134904 78358
rect 1790 77970 1796 78022
rect 1848 77970 1854 78022
rect 134840 77970 134846 78022
rect 134898 77970 134904 78022
rect 1790 77634 1796 77686
rect 1848 77634 1854 77686
rect 134840 77634 134846 77686
rect 134898 77634 134904 77686
rect 1790 77298 1796 77350
rect 1848 77298 1854 77350
rect 134840 77298 134846 77350
rect 134898 77298 134904 77350
rect 1790 76962 1796 77014
rect 1848 76962 1854 77014
rect 28614 76993 28620 77045
rect 28672 76993 28678 77045
rect 31110 76993 31116 77045
rect 31168 76993 31174 77045
rect 33606 76993 33612 77045
rect 33664 76993 33670 77045
rect 36102 76993 36108 77045
rect 36160 76993 36166 77045
rect 38598 76993 38604 77045
rect 38656 76993 38662 77045
rect 41094 76993 41100 77045
rect 41152 76993 41158 77045
rect 43590 76993 43596 77045
rect 43648 76993 43654 77045
rect 46086 76993 46092 77045
rect 46144 76993 46150 77045
rect 48582 76993 48588 77045
rect 48640 76993 48646 77045
rect 51078 76993 51084 77045
rect 51136 76993 51142 77045
rect 53574 76993 53580 77045
rect 53632 76993 53638 77045
rect 56070 76993 56076 77045
rect 56128 76993 56134 77045
rect 58566 76993 58572 77045
rect 58624 76993 58630 77045
rect 61062 76993 61068 77045
rect 61120 76993 61126 77045
rect 63558 76993 63564 77045
rect 63616 76993 63622 77045
rect 66054 76993 66060 77045
rect 66112 76993 66118 77045
rect 68550 76993 68556 77045
rect 68608 76993 68614 77045
rect 71046 76993 71052 77045
rect 71104 76993 71110 77045
rect 73542 76993 73548 77045
rect 73600 76993 73606 77045
rect 76038 76993 76044 77045
rect 76096 76993 76102 77045
rect 78534 76993 78540 77045
rect 78592 76993 78598 77045
rect 81030 76993 81036 77045
rect 81088 76993 81094 77045
rect 83526 76993 83532 77045
rect 83584 76993 83590 77045
rect 86022 76993 86028 77045
rect 86080 76993 86086 77045
rect 88518 76993 88524 77045
rect 88576 76993 88582 77045
rect 91014 76993 91020 77045
rect 91072 76993 91078 77045
rect 93510 76993 93516 77045
rect 93568 76993 93574 77045
rect 96006 76993 96012 77045
rect 96064 76993 96070 77045
rect 98502 76993 98508 77045
rect 98560 76993 98566 77045
rect 100998 76993 101004 77045
rect 101056 76993 101062 77045
rect 103494 76993 103500 77045
rect 103552 76993 103558 77045
rect 105990 76993 105996 77045
rect 106048 76993 106054 77045
rect 134840 76962 134846 77014
rect 134898 76962 134904 77014
rect 1790 76626 1796 76678
rect 1848 76626 1854 76678
rect 134840 76626 134846 76678
rect 134898 76626 134904 76678
rect 1790 76290 1796 76342
rect 1848 76290 1854 76342
rect 134840 76290 134846 76342
rect 134898 76290 134904 76342
rect 1790 75954 1796 76006
rect 1848 75954 1854 76006
rect 134840 75954 134846 76006
rect 134898 75954 134904 76006
rect 1790 75618 1796 75670
rect 1848 75618 1854 75670
rect 134840 75618 134846 75670
rect 134898 75618 134904 75670
rect 1790 75282 1796 75334
rect 1848 75282 1854 75334
rect 134840 75282 134846 75334
rect 134898 75282 134904 75334
rect 1790 74946 1796 74998
rect 1848 74946 1854 74998
rect 134840 74946 134846 74998
rect 134898 74946 134904 74998
rect 1790 74610 1796 74662
rect 1848 74610 1854 74662
rect 134840 74610 134846 74662
rect 134898 74610 134904 74662
rect 1790 74274 1796 74326
rect 1848 74274 1854 74326
rect 134840 74274 134846 74326
rect 134898 74274 134904 74326
rect 1790 73938 1796 73990
rect 1848 73938 1854 73990
rect 134840 73938 134846 73990
rect 134898 73938 134904 73990
rect 1790 73602 1796 73654
rect 1848 73602 1854 73654
rect 134840 73602 134846 73654
rect 134898 73602 134904 73654
rect 1790 73266 1796 73318
rect 1848 73266 1854 73318
rect 134840 73266 134846 73318
rect 134898 73266 134904 73318
rect 1790 72930 1796 72982
rect 1848 72930 1854 72982
rect 134840 72930 134846 72982
rect 134898 72930 134904 72982
rect 1790 72594 1796 72646
rect 1848 72594 1854 72646
rect 134840 72594 134846 72646
rect 134898 72594 134904 72646
rect 1790 72258 1796 72310
rect 1848 72258 1854 72310
rect 134840 72258 134846 72310
rect 134898 72258 134904 72310
rect 1790 71922 1796 71974
rect 1848 71922 1854 71974
rect 134840 71922 134846 71974
rect 134898 71922 134904 71974
rect 1790 71586 1796 71638
rect 1848 71586 1854 71638
rect 134840 71586 134846 71638
rect 134898 71586 134904 71638
rect 1790 71250 1796 71302
rect 1848 71250 1854 71302
rect 134840 71250 134846 71302
rect 134898 71250 134904 71302
rect 1790 70914 1796 70966
rect 1848 70914 1854 70966
rect 134840 70914 134846 70966
rect 134898 70914 134904 70966
rect 1790 70578 1796 70630
rect 1848 70578 1854 70630
rect 134840 70578 134846 70630
rect 134898 70578 134904 70630
rect 1790 70242 1796 70294
rect 1848 70242 1854 70294
rect 134840 70242 134846 70294
rect 134898 70242 134904 70294
rect 1790 69906 1796 69958
rect 1848 69906 1854 69958
rect 134840 69906 134846 69958
rect 134898 69906 134904 69958
rect 1790 69570 1796 69622
rect 1848 69570 1854 69622
rect 134840 69570 134846 69622
rect 134898 69570 134904 69622
rect 1790 69234 1796 69286
rect 1848 69234 1854 69286
rect 134840 69234 134846 69286
rect 134898 69234 134904 69286
rect 1790 68898 1796 68950
rect 1848 68898 1854 68950
rect 134840 68898 134846 68950
rect 134898 68898 134904 68950
rect 1790 68562 1796 68614
rect 1848 68562 1854 68614
rect 134840 68562 134846 68614
rect 134898 68562 134904 68614
rect 1790 68226 1796 68278
rect 1848 68226 1854 68278
rect 134840 68226 134846 68278
rect 134898 68226 134904 68278
rect 1790 67890 1796 67942
rect 1848 67890 1854 67942
rect 134840 67890 134846 67942
rect 134898 67890 134904 67942
rect 1790 67554 1796 67606
rect 1848 67554 1854 67606
rect 134840 67554 134846 67606
rect 134898 67554 134904 67606
rect 1790 67218 1796 67270
rect 1848 67218 1854 67270
rect 134840 67218 134846 67270
rect 134898 67218 134904 67270
rect 1790 66882 1796 66934
rect 1848 66882 1854 66934
rect 134840 66882 134846 66934
rect 134898 66882 134904 66934
rect 1790 66546 1796 66598
rect 1848 66546 1854 66598
rect 134840 66546 134846 66598
rect 134898 66546 134904 66598
rect 1790 66210 1796 66262
rect 1848 66210 1854 66262
rect 134840 66210 134846 66262
rect 134898 66210 134904 66262
rect 1790 65874 1796 65926
rect 1848 65874 1854 65926
rect 134840 65874 134846 65926
rect 134898 65874 134904 65926
rect 1790 65538 1796 65590
rect 1848 65538 1854 65590
rect 134840 65538 134846 65590
rect 134898 65538 134904 65590
rect 1790 65202 1796 65254
rect 1848 65202 1854 65254
rect 134840 65202 134846 65254
rect 134898 65202 134904 65254
rect 1790 64866 1796 64918
rect 1848 64866 1854 64918
rect 134840 64866 134846 64918
rect 134898 64866 134904 64918
rect 1790 64530 1796 64582
rect 1848 64530 1854 64582
rect 134840 64530 134846 64582
rect 134898 64530 134904 64582
rect 1790 64194 1796 64246
rect 1848 64194 1854 64246
rect 134840 64194 134846 64246
rect 134898 64194 134904 64246
rect 1790 63858 1796 63910
rect 1848 63858 1854 63910
rect 134840 63858 134846 63910
rect 134898 63858 134904 63910
rect 1790 63522 1796 63574
rect 1848 63522 1854 63574
rect 134840 63522 134846 63574
rect 134898 63522 134904 63574
rect 1790 63186 1796 63238
rect 1848 63186 1854 63238
rect 134840 63186 134846 63238
rect 134898 63186 134904 63238
rect 1790 62850 1796 62902
rect 1848 62850 1854 62902
rect 134840 62850 134846 62902
rect 134898 62850 134904 62902
rect 1790 62514 1796 62566
rect 1848 62514 1854 62566
rect 134840 62514 134846 62566
rect 134898 62514 134904 62566
rect 1790 62178 1796 62230
rect 1848 62178 1854 62230
rect 134840 62178 134846 62230
rect 134898 62178 134904 62230
rect 1790 61842 1796 61894
rect 1848 61842 1854 61894
rect 134840 61842 134846 61894
rect 134898 61842 134904 61894
rect 1790 61506 1796 61558
rect 1848 61506 1854 61558
rect 134840 61506 134846 61558
rect 134898 61506 134904 61558
rect 1790 61170 1796 61222
rect 1848 61170 1854 61222
rect 134840 61170 134846 61222
rect 134898 61170 134904 61222
rect 1790 60834 1796 60886
rect 1848 60834 1854 60886
rect 134840 60834 134846 60886
rect 134898 60834 134904 60886
rect 1790 60498 1796 60550
rect 1848 60498 1854 60550
rect 134840 60498 134846 60550
rect 134898 60498 134904 60550
rect 1790 60162 1796 60214
rect 1848 60162 1854 60214
rect 134840 60162 134846 60214
rect 134898 60162 134904 60214
rect 1790 59826 1796 59878
rect 1848 59826 1854 59878
rect 134840 59826 134846 59878
rect 134898 59826 134904 59878
rect 1790 59490 1796 59542
rect 1848 59490 1854 59542
rect 134840 59490 134846 59542
rect 134898 59490 134904 59542
rect 1790 59154 1796 59206
rect 1848 59154 1854 59206
rect 134840 59154 134846 59206
rect 134898 59154 134904 59206
rect 1790 58818 1796 58870
rect 1848 58818 1854 58870
rect 134840 58818 134846 58870
rect 134898 58818 134904 58870
rect 1790 58482 1796 58534
rect 1848 58482 1854 58534
rect 134840 58482 134846 58534
rect 134898 58482 134904 58534
rect 1790 58146 1796 58198
rect 1848 58146 1854 58198
rect 134840 58146 134846 58198
rect 134898 58146 134904 58198
rect 1790 57810 1796 57862
rect 1848 57810 1854 57862
rect 134840 57810 134846 57862
rect 134898 57810 134904 57862
rect 1790 57474 1796 57526
rect 1848 57474 1854 57526
rect 134840 57474 134846 57526
rect 134898 57474 134904 57526
rect 1790 57138 1796 57190
rect 1848 57138 1854 57190
rect 134840 57138 134846 57190
rect 134898 57138 134904 57190
rect 1790 56802 1796 56854
rect 1848 56802 1854 56854
rect 134840 56802 134846 56854
rect 134898 56802 134904 56854
rect 1790 56466 1796 56518
rect 1848 56466 1854 56518
rect 134840 56466 134846 56518
rect 134898 56466 134904 56518
rect 1790 56130 1796 56182
rect 1848 56130 1854 56182
rect 134840 56130 134846 56182
rect 134898 56130 134904 56182
rect 1790 55794 1796 55846
rect 1848 55794 1854 55846
rect 134840 55794 134846 55846
rect 134898 55794 134904 55846
rect 1790 55458 1796 55510
rect 1848 55458 1854 55510
rect 134840 55458 134846 55510
rect 134898 55458 134904 55510
rect 1790 55122 1796 55174
rect 1848 55122 1854 55174
rect 134840 55122 134846 55174
rect 134898 55122 134904 55174
rect 1790 54786 1796 54838
rect 1848 54786 1854 54838
rect 134840 54786 134846 54838
rect 134898 54786 134904 54838
rect 1790 54450 1796 54502
rect 1848 54450 1854 54502
rect 134840 54450 134846 54502
rect 134898 54450 134904 54502
rect 1790 54114 1796 54166
rect 1848 54114 1854 54166
rect 134840 54114 134846 54166
rect 134898 54114 134904 54166
rect 1790 53778 1796 53830
rect 1848 53778 1854 53830
rect 134840 53778 134846 53830
rect 134898 53778 134904 53830
rect 1790 53442 1796 53494
rect 1848 53442 1854 53494
rect 134840 53442 134846 53494
rect 134898 53442 134904 53494
rect 1790 53106 1796 53158
rect 1848 53106 1854 53158
rect 134840 53106 134846 53158
rect 134898 53106 134904 53158
rect 1790 52770 1796 52822
rect 1848 52770 1854 52822
rect 134840 52770 134846 52822
rect 134898 52770 134904 52822
rect 1790 52434 1796 52486
rect 1848 52434 1854 52486
rect 134840 52434 134846 52486
rect 134898 52434 134904 52486
rect 1790 52098 1796 52150
rect 1848 52098 1854 52150
rect 134840 52098 134846 52150
rect 134898 52098 134904 52150
rect 1790 51762 1796 51814
rect 1848 51762 1854 51814
rect 134840 51762 134846 51814
rect 134898 51762 134904 51814
rect 1790 51426 1796 51478
rect 1848 51426 1854 51478
rect 134840 51426 134846 51478
rect 134898 51426 134904 51478
rect 1790 51090 1796 51142
rect 1848 51090 1854 51142
rect 134840 51090 134846 51142
rect 134898 51090 134904 51142
rect 1790 50754 1796 50806
rect 1848 50754 1854 50806
rect 134840 50754 134846 50806
rect 134898 50754 134904 50806
rect 1790 50418 1796 50470
rect 1848 50418 1854 50470
rect 134840 50418 134846 50470
rect 134898 50418 134904 50470
rect 1790 50082 1796 50134
rect 1848 50082 1854 50134
rect 134840 50082 134846 50134
rect 134898 50082 134904 50134
rect 1790 49746 1796 49798
rect 1848 49746 1854 49798
rect 134840 49746 134846 49798
rect 134898 49746 134904 49798
rect 1790 49410 1796 49462
rect 1848 49410 1854 49462
rect 134840 49410 134846 49462
rect 134898 49410 134904 49462
rect 1790 49074 1796 49126
rect 1848 49074 1854 49126
rect 134840 49074 134846 49126
rect 134898 49074 134904 49126
rect 1790 48738 1796 48790
rect 1848 48738 1854 48790
rect 134840 48738 134846 48790
rect 134898 48738 134904 48790
rect 1790 48402 1796 48454
rect 1848 48402 1854 48454
rect 134840 48402 134846 48454
rect 134898 48402 134904 48454
rect 1790 48066 1796 48118
rect 1848 48066 1854 48118
rect 134840 48066 134846 48118
rect 134898 48066 134904 48118
rect 1790 47730 1796 47782
rect 1848 47730 1854 47782
rect 134840 47730 134846 47782
rect 134898 47730 134904 47782
rect 1790 47394 1796 47446
rect 1848 47394 1854 47446
rect 134840 47394 134846 47446
rect 134898 47394 134904 47446
rect 1790 47058 1796 47110
rect 1848 47058 1854 47110
rect 134840 47058 134846 47110
rect 134898 47058 134904 47110
rect 1790 46722 1796 46774
rect 1848 46722 1854 46774
rect 134840 46722 134846 46774
rect 134898 46722 134904 46774
rect 1790 46386 1796 46438
rect 1848 46386 1854 46438
rect 134840 46386 134846 46438
rect 134898 46386 134904 46438
rect 1790 46050 1796 46102
rect 1848 46050 1854 46102
rect 134840 46050 134846 46102
rect 134898 46050 134904 46102
rect 1790 45714 1796 45766
rect 1848 45714 1854 45766
rect 134840 45714 134846 45766
rect 134898 45714 134904 45766
rect 1790 45378 1796 45430
rect 1848 45378 1854 45430
rect 134840 45378 134846 45430
rect 134898 45378 134904 45430
rect 1790 45042 1796 45094
rect 1848 45042 1854 45094
rect 134840 45042 134846 45094
rect 134898 45042 134904 45094
rect 1790 44706 1796 44758
rect 1848 44706 1854 44758
rect 134840 44706 134846 44758
rect 134898 44706 134904 44758
rect 1790 44370 1796 44422
rect 1848 44370 1854 44422
rect 134840 44370 134846 44422
rect 134898 44370 134904 44422
rect 1790 44034 1796 44086
rect 1848 44034 1854 44086
rect 134840 44034 134846 44086
rect 134898 44034 134904 44086
rect 1790 43698 1796 43750
rect 1848 43698 1854 43750
rect 134840 43698 134846 43750
rect 134898 43698 134904 43750
rect 1790 43362 1796 43414
rect 1848 43362 1854 43414
rect 134840 43362 134846 43414
rect 134898 43362 134904 43414
rect 1790 43026 1796 43078
rect 1848 43026 1854 43078
rect 134840 43026 134846 43078
rect 134898 43026 134904 43078
rect 1790 42690 1796 42742
rect 1848 42690 1854 42742
rect 134840 42690 134846 42742
rect 134898 42690 134904 42742
rect 1790 42354 1796 42406
rect 1848 42354 1854 42406
rect 134840 42354 134846 42406
rect 134898 42354 134904 42406
rect 1790 42018 1796 42070
rect 1848 42018 1854 42070
rect 134840 42018 134846 42070
rect 134898 42018 134904 42070
rect 1790 41682 1796 41734
rect 1848 41682 1854 41734
rect 134840 41682 134846 41734
rect 134898 41682 134904 41734
rect 1790 41346 1796 41398
rect 1848 41346 1854 41398
rect 134840 41346 134846 41398
rect 134898 41346 134904 41398
rect 1790 41010 1796 41062
rect 1848 41010 1854 41062
rect 134840 41010 134846 41062
rect 134898 41010 134904 41062
rect 1790 40674 1796 40726
rect 1848 40674 1854 40726
rect 134840 40674 134846 40726
rect 134898 40674 134904 40726
rect 1790 40338 1796 40390
rect 1848 40338 1854 40390
rect 134840 40338 134846 40390
rect 134898 40338 134904 40390
rect 1790 40002 1796 40054
rect 1848 40002 1854 40054
rect 134840 40002 134846 40054
rect 134898 40002 134904 40054
rect 1790 39666 1796 39718
rect 1848 39666 1854 39718
rect 134840 39666 134846 39718
rect 134898 39666 134904 39718
rect 1790 39330 1796 39382
rect 1848 39330 1854 39382
rect 134840 39330 134846 39382
rect 134898 39330 134904 39382
rect 1790 38994 1796 39046
rect 1848 38994 1854 39046
rect 134840 38994 134846 39046
rect 134898 38994 134904 39046
rect 1790 38658 1796 38710
rect 1848 38658 1854 38710
rect 134840 38658 134846 38710
rect 134898 38658 134904 38710
rect 1790 38322 1796 38374
rect 1848 38322 1854 38374
rect 134840 38322 134846 38374
rect 134898 38322 134904 38374
rect 1790 37986 1796 38038
rect 1848 37986 1854 38038
rect 134840 37986 134846 38038
rect 134898 37986 134904 38038
rect 1790 37650 1796 37702
rect 1848 37650 1854 37702
rect 134840 37650 134846 37702
rect 134898 37650 134904 37702
rect 1790 37314 1796 37366
rect 1848 37314 1854 37366
rect 134840 37314 134846 37366
rect 134898 37314 134904 37366
rect 1790 36978 1796 37030
rect 1848 36978 1854 37030
rect 134840 36978 134846 37030
rect 134898 36978 134904 37030
rect 15343 36839 15349 36891
rect 15401 36839 15407 36891
rect 1790 36642 1796 36694
rect 1848 36642 1854 36694
rect 1790 36306 1796 36358
rect 1848 36306 1854 36358
rect 1790 35970 1796 36022
rect 1848 35970 1854 36022
rect 1790 35634 1796 35686
rect 1848 35634 1854 35686
rect 15263 35569 15269 35621
rect 15321 35569 15327 35621
rect 1790 35298 1796 35350
rect 1848 35298 1854 35350
rect 1790 34962 1796 35014
rect 1848 34962 1854 35014
rect 1790 34626 1796 34678
rect 1848 34626 1854 34678
rect 1790 34290 1796 34342
rect 1848 34290 1854 34342
rect 15183 34011 15189 34063
rect 15241 34011 15247 34063
rect 1790 33954 1796 34006
rect 1848 33954 1854 34006
rect 1790 33618 1796 33670
rect 1848 33618 1854 33670
rect 1790 33282 1796 33334
rect 1848 33282 1854 33334
rect 1790 32946 1796 32998
rect 1848 32946 1854 32998
rect 15103 32741 15109 32793
rect 15161 32741 15167 32793
rect 1790 32610 1796 32662
rect 1848 32610 1854 32662
rect 1790 32274 1796 32326
rect 1848 32274 1854 32326
rect 1790 31938 1796 31990
rect 1848 31938 1854 31990
rect 1790 31602 1796 31654
rect 1848 31602 1854 31654
rect 1790 31266 1796 31318
rect 1848 31266 1854 31318
rect 15023 31183 15029 31235
rect 15081 31183 15087 31235
rect 1790 30930 1796 30982
rect 1848 30930 1854 30982
rect 1790 30594 1796 30646
rect 1848 30594 1854 30646
rect 1790 30258 1796 30310
rect 1848 30258 1854 30310
rect 1790 29922 1796 29974
rect 1848 29922 1854 29974
rect 14943 29913 14949 29965
rect 15001 29913 15007 29965
rect 1790 29586 1796 29638
rect 1848 29586 1854 29638
rect 1790 29250 1796 29302
rect 1848 29250 1854 29302
rect 1790 28914 1796 28966
rect 1848 28914 1854 28966
rect 1790 28578 1796 28630
rect 1848 28578 1854 28630
rect 14863 28355 14869 28407
rect 14921 28355 14927 28407
rect 1790 28242 1796 28294
rect 1848 28242 1854 28294
rect 1790 27906 1796 27958
rect 1848 27906 1854 27958
rect 1790 27570 1796 27622
rect 1848 27570 1854 27622
rect 1790 27234 1796 27286
rect 1848 27234 1854 27286
rect 1790 26898 1796 26950
rect 1848 26898 1854 26950
rect 1790 26562 1796 26614
rect 1848 26562 1854 26614
rect 1790 26226 1796 26278
rect 1848 26226 1854 26278
rect 1790 25890 1796 25942
rect 1848 25890 1854 25942
rect 1790 25554 1796 25606
rect 1848 25554 1854 25606
rect 1790 25218 1796 25270
rect 1848 25218 1854 25270
rect 1790 24882 1796 24934
rect 1848 24882 1854 24934
rect 1790 24546 1796 24598
rect 1848 24546 1854 24598
rect 1790 24210 1796 24262
rect 1848 24210 1854 24262
rect 1790 23874 1796 23926
rect 1848 23874 1854 23926
rect 14881 23796 14909 28355
rect 14961 23796 14989 29913
rect 15041 23796 15069 31183
rect 15121 23796 15149 32741
rect 15201 23796 15229 34011
rect 15281 23796 15309 35569
rect 15361 23796 15389 36839
rect 134840 36642 134846 36694
rect 134898 36642 134904 36694
rect 134840 36306 134846 36358
rect 134898 36306 134904 36358
rect 134840 35970 134846 36022
rect 134898 35970 134904 36022
rect 134840 35634 134846 35686
rect 134898 35634 134904 35686
rect 134840 35298 134846 35350
rect 134898 35298 134904 35350
rect 134840 34962 134846 35014
rect 134898 34962 134904 35014
rect 134840 34626 134846 34678
rect 134898 34626 134904 34678
rect 134840 34290 134846 34342
rect 134898 34290 134904 34342
rect 134840 33954 134846 34006
rect 134898 33954 134904 34006
rect 134840 33618 134846 33670
rect 134898 33618 134904 33670
rect 134840 33282 134846 33334
rect 134898 33282 134904 33334
rect 134840 32946 134846 32998
rect 134898 32946 134904 32998
rect 134840 32610 134846 32662
rect 134898 32610 134904 32662
rect 134840 32274 134846 32326
rect 134898 32274 134904 32326
rect 134840 31938 134846 31990
rect 134898 31938 134904 31990
rect 134840 31602 134846 31654
rect 134898 31602 134904 31654
rect 134840 31266 134846 31318
rect 134898 31266 134904 31318
rect 134840 30930 134846 30982
rect 134898 30930 134904 30982
rect 134840 30594 134846 30646
rect 134898 30594 134904 30646
rect 134840 30258 134846 30310
rect 134898 30258 134904 30310
rect 134840 29922 134846 29974
rect 134898 29922 134904 29974
rect 134840 29586 134846 29638
rect 134898 29586 134904 29638
rect 134840 29250 134846 29302
rect 134898 29250 134904 29302
rect 134840 28914 134846 28966
rect 134898 28914 134904 28966
rect 134840 28578 134846 28630
rect 134898 28578 134904 28630
rect 134840 28242 134846 28294
rect 134898 28242 134904 28294
rect 134840 27906 134846 27958
rect 134898 27906 134904 27958
rect 134840 27570 134846 27622
rect 134898 27570 134904 27622
rect 134840 27234 134846 27286
rect 134898 27234 134904 27286
rect 134840 26898 134846 26950
rect 134898 26898 134904 26950
rect 134840 26562 134846 26614
rect 134898 26562 134904 26614
rect 134840 26226 134846 26278
rect 134898 26226 134904 26278
rect 134840 25890 134846 25942
rect 134898 25890 134904 25942
rect 134840 25554 134846 25606
rect 134898 25554 134904 25606
rect 134840 25218 134846 25270
rect 134898 25218 134904 25270
rect 134840 24882 134846 24934
rect 134898 24882 134904 24934
rect 134840 24546 134846 24598
rect 134898 24546 134904 24598
rect 134840 24210 134846 24262
rect 134898 24210 134904 24262
rect 134840 23874 134846 23926
rect 134898 23874 134904 23926
rect 1790 23538 1796 23590
rect 1848 23538 1854 23590
rect 1790 23202 1796 23254
rect 1848 23202 1854 23254
rect 1790 22866 1796 22918
rect 1848 22866 1854 22918
rect 1790 22530 1796 22582
rect 1848 22530 1854 22582
rect 1790 22194 1796 22246
rect 1848 22194 1854 22246
rect 1790 21858 1796 21910
rect 1848 21858 1854 21910
rect 1790 21522 1796 21574
rect 1848 21522 1854 21574
rect 1790 21186 1796 21238
rect 1848 21186 1854 21238
rect 1790 20850 1796 20902
rect 1848 20850 1854 20902
rect 1790 20514 1796 20566
rect 1848 20514 1854 20566
rect 1790 20178 1796 20230
rect 1848 20178 1854 20230
rect 1790 19842 1796 19894
rect 1848 19842 1854 19894
rect 1790 19506 1796 19558
rect 1848 19506 1854 19558
rect 1790 19170 1796 19222
rect 1848 19170 1854 19222
rect 1790 18834 1796 18886
rect 1848 18834 1854 18886
rect 1790 18498 1796 18550
rect 1848 18498 1854 18550
rect 1790 18162 1796 18214
rect 1848 18162 1854 18214
rect 1790 17826 1796 17878
rect 1848 17826 1854 17878
rect 1790 17490 1796 17542
rect 1848 17490 1854 17542
rect 1790 17154 1796 17206
rect 1848 17154 1854 17206
rect 1790 16818 1796 16870
rect 1848 16818 1854 16870
rect 1790 16482 1796 16534
rect 1848 16482 1854 16534
rect 1790 16146 1796 16198
rect 1848 16146 1854 16198
rect 1790 15810 1796 15862
rect 1848 15810 1854 15862
rect 1790 15474 1796 15526
rect 1848 15474 1854 15526
rect 1790 15138 1796 15190
rect 1848 15138 1854 15190
rect 1790 14802 1796 14854
rect 1848 14802 1854 14854
rect 1790 14466 1796 14518
rect 1848 14466 1854 14518
rect 1790 14130 1796 14182
rect 1848 14130 1854 14182
rect 1790 13794 1796 13846
rect 1848 13794 1854 13846
rect 1790 13458 1796 13510
rect 1848 13458 1854 13510
rect 28614 13207 28620 13259
rect 28672 13207 28678 13259
rect 31110 13207 31116 13259
rect 31168 13207 31174 13259
rect 33606 13207 33612 13259
rect 33664 13207 33670 13259
rect 36102 13207 36108 13259
rect 36160 13207 36166 13259
rect 38598 13207 38604 13259
rect 38656 13207 38662 13259
rect 41094 13207 41100 13259
rect 41152 13207 41158 13259
rect 43590 13207 43596 13259
rect 43648 13207 43654 13259
rect 46086 13207 46092 13259
rect 46144 13207 46150 13259
rect 48582 13207 48588 13259
rect 48640 13207 48646 13259
rect 51078 13207 51084 13259
rect 51136 13207 51142 13259
rect 53574 13207 53580 13259
rect 53632 13207 53638 13259
rect 56070 13207 56076 13259
rect 56128 13207 56134 13259
rect 58566 13207 58572 13259
rect 58624 13207 58630 13259
rect 61062 13207 61068 13259
rect 61120 13207 61126 13259
rect 63558 13207 63564 13259
rect 63616 13207 63622 13259
rect 66054 13207 66060 13259
rect 66112 13207 66118 13259
rect 68550 13207 68556 13259
rect 68608 13207 68614 13259
rect 71046 13207 71052 13259
rect 71104 13207 71110 13259
rect 73542 13207 73548 13259
rect 73600 13207 73606 13259
rect 76038 13207 76044 13259
rect 76096 13207 76102 13259
rect 78534 13207 78540 13259
rect 78592 13207 78598 13259
rect 81030 13207 81036 13259
rect 81088 13207 81094 13259
rect 83526 13207 83532 13259
rect 83584 13207 83590 13259
rect 86022 13207 86028 13259
rect 86080 13207 86086 13259
rect 88518 13207 88524 13259
rect 88576 13207 88582 13259
rect 91014 13207 91020 13259
rect 91072 13207 91078 13259
rect 93510 13207 93516 13259
rect 93568 13207 93574 13259
rect 96006 13207 96012 13259
rect 96064 13207 96070 13259
rect 98502 13207 98508 13259
rect 98560 13207 98566 13259
rect 100998 13207 101004 13259
rect 101056 13207 101062 13259
rect 103494 13207 103500 13259
rect 103552 13207 103558 13259
rect 105990 13207 105996 13259
rect 106048 13207 106054 13259
rect 1790 13122 1796 13174
rect 1848 13122 1854 13174
rect 1790 12786 1796 12838
rect 1848 12786 1854 12838
rect 1790 12450 1796 12502
rect 1848 12450 1854 12502
rect 1790 12114 1796 12166
rect 1848 12114 1854 12166
rect 1790 11778 1796 11830
rect 1848 11778 1854 11830
rect 1790 11442 1796 11494
rect 1848 11442 1854 11494
rect 1790 11106 1796 11158
rect 1848 11106 1854 11158
rect 1790 10770 1796 10822
rect 1848 10770 1854 10822
rect 121521 10753 121549 23796
rect 121601 12023 121629 23796
rect 121681 13581 121709 23796
rect 121761 14851 121789 23796
rect 121841 16409 121869 23796
rect 121921 17679 121949 23796
rect 122001 19237 122029 23796
rect 134840 23538 134846 23590
rect 134898 23538 134904 23590
rect 134840 23202 134846 23254
rect 134898 23202 134904 23254
rect 134840 22866 134846 22918
rect 134898 22866 134904 22918
rect 134840 22530 134846 22582
rect 134898 22530 134904 22582
rect 134840 22194 134846 22246
rect 134898 22194 134904 22246
rect 134840 21858 134846 21910
rect 134898 21858 134904 21910
rect 134840 21522 134846 21574
rect 134898 21522 134904 21574
rect 134840 21186 134846 21238
rect 134898 21186 134904 21238
rect 134840 20850 134846 20902
rect 134898 20850 134904 20902
rect 134840 20514 134846 20566
rect 134898 20514 134904 20566
rect 134840 20178 134846 20230
rect 134898 20178 134904 20230
rect 134840 19842 134846 19894
rect 134898 19842 134904 19894
rect 134840 19506 134846 19558
rect 134898 19506 134904 19558
rect 121983 19185 121989 19237
rect 122041 19185 122047 19237
rect 134840 19170 134846 19222
rect 134898 19170 134904 19222
rect 134840 18834 134846 18886
rect 134898 18834 134904 18886
rect 134840 18498 134846 18550
rect 134898 18498 134904 18550
rect 134840 18162 134846 18214
rect 134898 18162 134904 18214
rect 134840 17826 134846 17878
rect 134898 17826 134904 17878
rect 121903 17627 121909 17679
rect 121961 17627 121967 17679
rect 134840 17490 134846 17542
rect 134898 17490 134904 17542
rect 134840 17154 134846 17206
rect 134898 17154 134904 17206
rect 134840 16818 134846 16870
rect 134898 16818 134904 16870
rect 134840 16482 134846 16534
rect 134898 16482 134904 16534
rect 121823 16357 121829 16409
rect 121881 16357 121887 16409
rect 134840 16146 134846 16198
rect 134898 16146 134904 16198
rect 134840 15810 134846 15862
rect 134898 15810 134904 15862
rect 134840 15474 134846 15526
rect 134898 15474 134904 15526
rect 134840 15138 134846 15190
rect 134898 15138 134904 15190
rect 121743 14799 121749 14851
rect 121801 14799 121807 14851
rect 134840 14802 134846 14854
rect 134898 14802 134904 14854
rect 134840 14466 134846 14518
rect 134898 14466 134904 14518
rect 134840 14130 134846 14182
rect 134898 14130 134904 14182
rect 134840 13794 134846 13846
rect 134898 13794 134904 13846
rect 121663 13529 121669 13581
rect 121721 13529 121727 13581
rect 134840 13458 134846 13510
rect 134898 13458 134904 13510
rect 134840 13122 134846 13174
rect 134898 13122 134904 13174
rect 134840 12786 134846 12838
rect 134898 12786 134904 12838
rect 134840 12450 134846 12502
rect 134898 12450 134904 12502
rect 134840 12114 134846 12166
rect 134898 12114 134904 12166
rect 121583 11971 121589 12023
rect 121641 11971 121647 12023
rect 134840 11778 134846 11830
rect 134898 11778 134904 11830
rect 134840 11442 134846 11494
rect 134898 11442 134904 11494
rect 134840 11106 134846 11158
rect 134898 11106 134904 11158
rect 134840 10770 134846 10822
rect 134898 10770 134904 10822
rect 121503 10701 121509 10753
rect 121561 10701 121567 10753
rect 1790 10434 1796 10486
rect 1848 10434 1854 10486
rect 134840 10434 134846 10486
rect 134898 10434 134904 10486
rect 1790 10098 1796 10150
rect 1848 10098 1854 10150
rect 134840 10098 134846 10150
rect 134898 10098 134904 10150
rect 1790 9762 1796 9814
rect 1848 9762 1854 9814
rect 134840 9762 134846 9814
rect 134898 9762 134904 9814
rect 1790 9426 1796 9478
rect 1848 9426 1854 9478
rect 134840 9426 134846 9478
rect 134898 9426 134904 9478
rect 1790 9090 1796 9142
rect 1848 9090 1854 9142
rect 134840 9090 134846 9142
rect 134898 9090 134904 9142
rect 1790 8754 1796 8806
rect 1848 8754 1854 8806
rect 134840 8754 134846 8806
rect 134898 8754 134904 8806
rect 1790 8418 1796 8470
rect 1848 8418 1854 8470
rect 134840 8418 134846 8470
rect 134898 8418 134904 8470
rect 1790 8082 1796 8134
rect 1848 8082 1854 8134
rect 134840 8082 134846 8134
rect 134898 8082 134904 8134
rect 1790 7746 1796 7798
rect 1848 7746 1854 7798
rect 134840 7746 134846 7798
rect 134898 7746 134904 7798
rect 1790 7410 1796 7462
rect 1848 7410 1854 7462
rect 134840 7410 134846 7462
rect 134898 7410 134904 7462
rect 1790 7074 1796 7126
rect 1848 7074 1854 7126
rect 134840 7074 134846 7126
rect 134898 7074 134904 7126
rect 1790 6738 1796 6790
rect 1848 6738 1854 6790
rect 134840 6738 134846 6790
rect 134898 6738 134904 6790
rect 1790 6402 1796 6454
rect 1848 6402 1854 6454
rect 134840 6402 134846 6454
rect 134898 6402 134904 6454
rect 1790 6066 1796 6118
rect 1848 6066 1854 6118
rect 134840 6066 134846 6118
rect 134898 6066 134904 6118
rect 1790 5730 1796 5782
rect 1848 5730 1854 5782
rect 134840 5730 134846 5782
rect 134898 5730 134904 5782
rect 1790 5394 1796 5446
rect 1848 5394 1854 5446
rect 134840 5394 134846 5446
rect 134898 5394 134904 5446
rect 1790 5058 1796 5110
rect 1848 5058 1854 5110
rect 134840 5058 134846 5110
rect 134898 5058 134904 5110
rect 1790 4722 1796 4774
rect 1848 4722 1854 4774
rect 134840 4722 134846 4774
rect 134898 4722 134904 4774
rect 1790 4386 1796 4438
rect 1848 4386 1854 4438
rect 134840 4386 134846 4438
rect 134898 4386 134904 4438
rect 1790 4050 1796 4102
rect 1848 4050 1854 4102
rect 134840 4050 134846 4102
rect 134898 4050 134904 4102
rect 1790 3714 1796 3766
rect 1848 3714 1854 3766
rect 134840 3714 134846 3766
rect 134898 3714 134904 3766
rect 1790 3378 1796 3430
rect 1848 3378 1854 3430
rect 134840 3378 134846 3430
rect 134898 3378 134904 3430
rect 1790 3042 1796 3094
rect 1848 3042 1854 3094
rect 134840 3042 134846 3094
rect 134898 3042 134904 3094
rect 1790 2706 1796 2758
rect 1848 2706 1854 2758
rect 134840 2706 134846 2758
rect 134898 2706 134904 2758
rect 1790 2370 1796 2422
rect 1848 2370 1854 2422
rect 134840 2370 134846 2422
rect 134898 2370 134904 2422
rect 1790 2034 1796 2086
rect 1848 2034 1854 2086
rect 134840 2034 134846 2086
rect 134898 2034 134904 2086
rect 1710 1750 134984 1836
rect 1710 1698 2132 1750
rect 2184 1741 3812 1750
rect 3864 1741 5492 1750
rect 5544 1741 7172 1750
rect 7224 1741 8852 1750
rect 8904 1741 10532 1750
rect 10584 1741 12212 1750
rect 12264 1741 13892 1750
rect 13944 1741 15572 1750
rect 15624 1741 17252 1750
rect 17304 1741 18932 1750
rect 18984 1741 20612 1750
rect 20664 1741 22292 1750
rect 22344 1741 23972 1750
rect 24024 1741 25652 1750
rect 25704 1741 27332 1750
rect 27384 1741 29012 1750
rect 29064 1741 30692 1750
rect 30744 1741 32372 1750
rect 32424 1741 34052 1750
rect 34104 1741 35732 1750
rect 35784 1741 37412 1750
rect 37464 1741 39092 1750
rect 39144 1741 40772 1750
rect 40824 1741 42452 1750
rect 42504 1741 44132 1750
rect 44184 1741 45812 1750
rect 45864 1741 47492 1750
rect 47544 1741 49172 1750
rect 49224 1741 50852 1750
rect 50904 1741 52532 1750
rect 52584 1741 54212 1750
rect 54264 1741 55892 1750
rect 55944 1741 57572 1750
rect 57624 1741 59252 1750
rect 59304 1741 60932 1750
rect 60984 1741 62612 1750
rect 62664 1741 64292 1750
rect 64344 1741 65972 1750
rect 66024 1741 67652 1750
rect 67704 1741 69332 1750
rect 69384 1741 71012 1750
rect 71064 1741 72692 1750
rect 72744 1741 74372 1750
rect 74424 1741 76052 1750
rect 76104 1741 77732 1750
rect 77784 1741 79412 1750
rect 79464 1741 81092 1750
rect 81144 1741 82772 1750
rect 82824 1741 84452 1750
rect 84504 1741 86132 1750
rect 86184 1741 87812 1750
rect 87864 1741 89492 1750
rect 89544 1741 91172 1750
rect 91224 1741 92852 1750
rect 92904 1741 94532 1750
rect 94584 1741 96212 1750
rect 96264 1741 97892 1750
rect 97944 1741 99572 1750
rect 99624 1741 101252 1750
rect 101304 1741 102932 1750
rect 102984 1741 104612 1750
rect 104664 1741 106292 1750
rect 106344 1741 107972 1750
rect 108024 1741 109652 1750
rect 109704 1741 111332 1750
rect 111384 1741 113012 1750
rect 113064 1741 114692 1750
rect 114744 1741 116372 1750
rect 116424 1741 118052 1750
rect 118104 1741 119732 1750
rect 119784 1741 121412 1750
rect 121464 1741 123092 1750
rect 123144 1741 124772 1750
rect 124824 1741 126452 1750
rect 126504 1741 128132 1750
rect 128184 1741 129812 1750
rect 129864 1741 131492 1750
rect 131544 1741 133172 1750
rect 133224 1741 134984 1750
rect 2184 1707 2477 1741
rect 2511 1707 2813 1741
rect 2847 1707 3149 1741
rect 3183 1707 3485 1741
rect 3519 1707 3812 1741
rect 3864 1707 4157 1741
rect 4191 1707 4493 1741
rect 4527 1707 4829 1741
rect 4863 1707 5165 1741
rect 5199 1707 5492 1741
rect 5544 1707 5837 1741
rect 5871 1707 6173 1741
rect 6207 1707 6509 1741
rect 6543 1707 6845 1741
rect 6879 1707 7172 1741
rect 7224 1707 7517 1741
rect 7551 1707 7853 1741
rect 7887 1707 8189 1741
rect 8223 1707 8525 1741
rect 8559 1707 8852 1741
rect 8904 1707 9197 1741
rect 9231 1707 9533 1741
rect 9567 1707 9869 1741
rect 9903 1707 10205 1741
rect 10239 1707 10532 1741
rect 10584 1707 10877 1741
rect 10911 1707 11213 1741
rect 11247 1707 11549 1741
rect 11583 1707 11885 1741
rect 11919 1707 12212 1741
rect 12264 1707 12557 1741
rect 12591 1707 12893 1741
rect 12927 1707 13229 1741
rect 13263 1707 13565 1741
rect 13599 1707 13892 1741
rect 13944 1707 14237 1741
rect 14271 1707 14573 1741
rect 14607 1707 14909 1741
rect 14943 1707 15245 1741
rect 15279 1707 15572 1741
rect 15624 1707 15917 1741
rect 15951 1707 16253 1741
rect 16287 1707 16589 1741
rect 16623 1707 16925 1741
rect 16959 1707 17252 1741
rect 17304 1707 17597 1741
rect 17631 1707 17933 1741
rect 17967 1707 18269 1741
rect 18303 1707 18605 1741
rect 18639 1707 18932 1741
rect 18984 1707 19277 1741
rect 19311 1707 19613 1741
rect 19647 1707 19949 1741
rect 19983 1707 20285 1741
rect 20319 1707 20612 1741
rect 20664 1707 20957 1741
rect 20991 1707 21293 1741
rect 21327 1707 21629 1741
rect 21663 1707 21965 1741
rect 21999 1707 22292 1741
rect 22344 1707 22637 1741
rect 22671 1707 22973 1741
rect 23007 1707 23309 1741
rect 23343 1707 23645 1741
rect 23679 1707 23972 1741
rect 24024 1707 24317 1741
rect 24351 1707 24653 1741
rect 24687 1707 24989 1741
rect 25023 1707 25325 1741
rect 25359 1707 25652 1741
rect 25704 1707 25997 1741
rect 26031 1707 26333 1741
rect 26367 1707 26669 1741
rect 26703 1707 27005 1741
rect 27039 1707 27332 1741
rect 27384 1707 27677 1741
rect 27711 1707 28013 1741
rect 28047 1707 28349 1741
rect 28383 1707 28685 1741
rect 28719 1707 29012 1741
rect 29064 1707 29357 1741
rect 29391 1707 29693 1741
rect 29727 1707 30029 1741
rect 30063 1707 30365 1741
rect 30399 1707 30692 1741
rect 30744 1707 31037 1741
rect 31071 1707 31373 1741
rect 31407 1707 31709 1741
rect 31743 1707 32045 1741
rect 32079 1707 32372 1741
rect 32424 1707 32717 1741
rect 32751 1707 33053 1741
rect 33087 1707 33389 1741
rect 33423 1707 33725 1741
rect 33759 1707 34052 1741
rect 34104 1707 34397 1741
rect 34431 1707 34733 1741
rect 34767 1707 35069 1741
rect 35103 1707 35405 1741
rect 35439 1707 35732 1741
rect 35784 1707 36077 1741
rect 36111 1707 36413 1741
rect 36447 1707 36749 1741
rect 36783 1707 37085 1741
rect 37119 1707 37412 1741
rect 37464 1707 37757 1741
rect 37791 1707 38093 1741
rect 38127 1707 38429 1741
rect 38463 1707 38765 1741
rect 38799 1707 39092 1741
rect 39144 1707 39437 1741
rect 39471 1707 39773 1741
rect 39807 1707 40109 1741
rect 40143 1707 40445 1741
rect 40479 1707 40772 1741
rect 40824 1707 41117 1741
rect 41151 1707 41453 1741
rect 41487 1707 41789 1741
rect 41823 1707 42125 1741
rect 42159 1707 42452 1741
rect 42504 1707 42797 1741
rect 42831 1707 43133 1741
rect 43167 1707 43469 1741
rect 43503 1707 43805 1741
rect 43839 1707 44132 1741
rect 44184 1707 44477 1741
rect 44511 1707 44813 1741
rect 44847 1707 45149 1741
rect 45183 1707 45485 1741
rect 45519 1707 45812 1741
rect 45864 1707 46157 1741
rect 46191 1707 46493 1741
rect 46527 1707 46829 1741
rect 46863 1707 47165 1741
rect 47199 1707 47492 1741
rect 47544 1707 47837 1741
rect 47871 1707 48173 1741
rect 48207 1707 48509 1741
rect 48543 1707 48845 1741
rect 48879 1707 49172 1741
rect 49224 1707 49517 1741
rect 49551 1707 49853 1741
rect 49887 1707 50189 1741
rect 50223 1707 50525 1741
rect 50559 1707 50852 1741
rect 50904 1707 51197 1741
rect 51231 1707 51533 1741
rect 51567 1707 51869 1741
rect 51903 1707 52205 1741
rect 52239 1707 52532 1741
rect 52584 1707 52877 1741
rect 52911 1707 53213 1741
rect 53247 1707 53549 1741
rect 53583 1707 53885 1741
rect 53919 1707 54212 1741
rect 54264 1707 54557 1741
rect 54591 1707 54893 1741
rect 54927 1707 55229 1741
rect 55263 1707 55565 1741
rect 55599 1707 55892 1741
rect 55944 1707 56237 1741
rect 56271 1707 56573 1741
rect 56607 1707 56909 1741
rect 56943 1707 57245 1741
rect 57279 1707 57572 1741
rect 57624 1707 57917 1741
rect 57951 1707 58253 1741
rect 58287 1707 58589 1741
rect 58623 1707 58925 1741
rect 58959 1707 59252 1741
rect 59304 1707 59597 1741
rect 59631 1707 59933 1741
rect 59967 1707 60269 1741
rect 60303 1707 60605 1741
rect 60639 1707 60932 1741
rect 60984 1707 61277 1741
rect 61311 1707 61613 1741
rect 61647 1707 61949 1741
rect 61983 1707 62285 1741
rect 62319 1707 62612 1741
rect 62664 1707 62957 1741
rect 62991 1707 63293 1741
rect 63327 1707 63629 1741
rect 63663 1707 63965 1741
rect 63999 1707 64292 1741
rect 64344 1707 64637 1741
rect 64671 1707 64973 1741
rect 65007 1707 65309 1741
rect 65343 1707 65645 1741
rect 65679 1707 65972 1741
rect 66024 1707 66317 1741
rect 66351 1707 66653 1741
rect 66687 1707 66989 1741
rect 67023 1707 67325 1741
rect 67359 1707 67652 1741
rect 67704 1707 67997 1741
rect 68031 1707 68333 1741
rect 68367 1707 68669 1741
rect 68703 1707 69005 1741
rect 69039 1707 69332 1741
rect 69384 1707 69677 1741
rect 69711 1707 70013 1741
rect 70047 1707 70349 1741
rect 70383 1707 70685 1741
rect 70719 1707 71012 1741
rect 71064 1707 71357 1741
rect 71391 1707 71693 1741
rect 71727 1707 72029 1741
rect 72063 1707 72365 1741
rect 72399 1707 72692 1741
rect 72744 1707 73037 1741
rect 73071 1707 73373 1741
rect 73407 1707 73709 1741
rect 73743 1707 74045 1741
rect 74079 1707 74372 1741
rect 74424 1707 74717 1741
rect 74751 1707 75053 1741
rect 75087 1707 75389 1741
rect 75423 1707 75725 1741
rect 75759 1707 76052 1741
rect 76104 1707 76397 1741
rect 76431 1707 76733 1741
rect 76767 1707 77069 1741
rect 77103 1707 77405 1741
rect 77439 1707 77732 1741
rect 77784 1707 78077 1741
rect 78111 1707 78413 1741
rect 78447 1707 78749 1741
rect 78783 1707 79085 1741
rect 79119 1707 79412 1741
rect 79464 1707 79757 1741
rect 79791 1707 80093 1741
rect 80127 1707 80429 1741
rect 80463 1707 80765 1741
rect 80799 1707 81092 1741
rect 81144 1707 81437 1741
rect 81471 1707 81773 1741
rect 81807 1707 82109 1741
rect 82143 1707 82445 1741
rect 82479 1707 82772 1741
rect 82824 1707 83117 1741
rect 83151 1707 83453 1741
rect 83487 1707 83789 1741
rect 83823 1707 84125 1741
rect 84159 1707 84452 1741
rect 84504 1707 84797 1741
rect 84831 1707 85133 1741
rect 85167 1707 85469 1741
rect 85503 1707 85805 1741
rect 85839 1707 86132 1741
rect 86184 1707 86477 1741
rect 86511 1707 86813 1741
rect 86847 1707 87149 1741
rect 87183 1707 87485 1741
rect 87519 1707 87812 1741
rect 87864 1707 88157 1741
rect 88191 1707 88493 1741
rect 88527 1707 88829 1741
rect 88863 1707 89165 1741
rect 89199 1707 89492 1741
rect 89544 1707 89837 1741
rect 89871 1707 90173 1741
rect 90207 1707 90509 1741
rect 90543 1707 90845 1741
rect 90879 1707 91172 1741
rect 91224 1707 91517 1741
rect 91551 1707 91853 1741
rect 91887 1707 92189 1741
rect 92223 1707 92525 1741
rect 92559 1707 92852 1741
rect 92904 1707 93197 1741
rect 93231 1707 93533 1741
rect 93567 1707 93869 1741
rect 93903 1707 94205 1741
rect 94239 1707 94532 1741
rect 94584 1707 94877 1741
rect 94911 1707 95213 1741
rect 95247 1707 95549 1741
rect 95583 1707 95885 1741
rect 95919 1707 96212 1741
rect 96264 1707 96557 1741
rect 96591 1707 96893 1741
rect 96927 1707 97229 1741
rect 97263 1707 97565 1741
rect 97599 1707 97892 1741
rect 97944 1707 98237 1741
rect 98271 1707 98573 1741
rect 98607 1707 98909 1741
rect 98943 1707 99245 1741
rect 99279 1707 99572 1741
rect 99624 1707 99917 1741
rect 99951 1707 100253 1741
rect 100287 1707 100589 1741
rect 100623 1707 100925 1741
rect 100959 1707 101252 1741
rect 101304 1707 101597 1741
rect 101631 1707 101933 1741
rect 101967 1707 102269 1741
rect 102303 1707 102605 1741
rect 102639 1707 102932 1741
rect 102984 1707 103277 1741
rect 103311 1707 103613 1741
rect 103647 1707 103949 1741
rect 103983 1707 104285 1741
rect 104319 1707 104612 1741
rect 104664 1707 104957 1741
rect 104991 1707 105293 1741
rect 105327 1707 105629 1741
rect 105663 1707 105965 1741
rect 105999 1707 106292 1741
rect 106344 1707 106637 1741
rect 106671 1707 106973 1741
rect 107007 1707 107309 1741
rect 107343 1707 107645 1741
rect 107679 1707 107972 1741
rect 108024 1707 108317 1741
rect 108351 1707 108653 1741
rect 108687 1707 108989 1741
rect 109023 1707 109325 1741
rect 109359 1707 109652 1741
rect 109704 1707 109997 1741
rect 110031 1707 110333 1741
rect 110367 1707 110669 1741
rect 110703 1707 111005 1741
rect 111039 1707 111332 1741
rect 111384 1707 111677 1741
rect 111711 1707 112013 1741
rect 112047 1707 112349 1741
rect 112383 1707 112685 1741
rect 112719 1707 113012 1741
rect 113064 1707 113357 1741
rect 113391 1707 113693 1741
rect 113727 1707 114029 1741
rect 114063 1707 114365 1741
rect 114399 1707 114692 1741
rect 114744 1707 115037 1741
rect 115071 1707 115373 1741
rect 115407 1707 115709 1741
rect 115743 1707 116045 1741
rect 116079 1707 116372 1741
rect 116424 1707 116717 1741
rect 116751 1707 117053 1741
rect 117087 1707 117389 1741
rect 117423 1707 117725 1741
rect 117759 1707 118052 1741
rect 118104 1707 118397 1741
rect 118431 1707 118733 1741
rect 118767 1707 119069 1741
rect 119103 1707 119405 1741
rect 119439 1707 119732 1741
rect 119784 1707 120077 1741
rect 120111 1707 120413 1741
rect 120447 1707 120749 1741
rect 120783 1707 121085 1741
rect 121119 1707 121412 1741
rect 121464 1707 121757 1741
rect 121791 1707 122093 1741
rect 122127 1707 122429 1741
rect 122463 1707 122765 1741
rect 122799 1707 123092 1741
rect 123144 1707 123437 1741
rect 123471 1707 123773 1741
rect 123807 1707 124109 1741
rect 124143 1707 124445 1741
rect 124479 1707 124772 1741
rect 124824 1707 125117 1741
rect 125151 1707 125453 1741
rect 125487 1707 125789 1741
rect 125823 1707 126125 1741
rect 126159 1707 126452 1741
rect 126504 1707 126797 1741
rect 126831 1707 127133 1741
rect 127167 1707 127469 1741
rect 127503 1707 127805 1741
rect 127839 1707 128132 1741
rect 128184 1707 128477 1741
rect 128511 1707 128813 1741
rect 128847 1707 129149 1741
rect 129183 1707 129485 1741
rect 129519 1707 129812 1741
rect 129864 1707 130157 1741
rect 130191 1707 130493 1741
rect 130527 1707 130829 1741
rect 130863 1707 131165 1741
rect 131199 1707 131492 1741
rect 131544 1707 131837 1741
rect 131871 1707 132173 1741
rect 132207 1707 132509 1741
rect 132543 1707 132845 1741
rect 132879 1707 133172 1741
rect 133224 1707 133517 1741
rect 133551 1707 133853 1741
rect 133887 1707 134189 1741
rect 134223 1707 134984 1741
rect 2184 1698 3812 1707
rect 3864 1698 5492 1707
rect 5544 1698 7172 1707
rect 7224 1698 8852 1707
rect 8904 1698 10532 1707
rect 10584 1698 12212 1707
rect 12264 1698 13892 1707
rect 13944 1698 15572 1707
rect 15624 1698 17252 1707
rect 17304 1698 18932 1707
rect 18984 1698 20612 1707
rect 20664 1698 22292 1707
rect 22344 1698 23972 1707
rect 24024 1698 25652 1707
rect 25704 1698 27332 1707
rect 27384 1698 29012 1707
rect 29064 1698 30692 1707
rect 30744 1698 32372 1707
rect 32424 1698 34052 1707
rect 34104 1698 35732 1707
rect 35784 1698 37412 1707
rect 37464 1698 39092 1707
rect 39144 1698 40772 1707
rect 40824 1698 42452 1707
rect 42504 1698 44132 1707
rect 44184 1698 45812 1707
rect 45864 1698 47492 1707
rect 47544 1698 49172 1707
rect 49224 1698 50852 1707
rect 50904 1698 52532 1707
rect 52584 1698 54212 1707
rect 54264 1698 55892 1707
rect 55944 1698 57572 1707
rect 57624 1698 59252 1707
rect 59304 1698 60932 1707
rect 60984 1698 62612 1707
rect 62664 1698 64292 1707
rect 64344 1698 65972 1707
rect 66024 1698 67652 1707
rect 67704 1698 69332 1707
rect 69384 1698 71012 1707
rect 71064 1698 72692 1707
rect 72744 1698 74372 1707
rect 74424 1698 76052 1707
rect 76104 1698 77732 1707
rect 77784 1698 79412 1707
rect 79464 1698 81092 1707
rect 81144 1698 82772 1707
rect 82824 1698 84452 1707
rect 84504 1698 86132 1707
rect 86184 1698 87812 1707
rect 87864 1698 89492 1707
rect 89544 1698 91172 1707
rect 91224 1698 92852 1707
rect 92904 1698 94532 1707
rect 94584 1698 96212 1707
rect 96264 1698 97892 1707
rect 97944 1698 99572 1707
rect 99624 1698 101252 1707
rect 101304 1698 102932 1707
rect 102984 1698 104612 1707
rect 104664 1698 106292 1707
rect 106344 1698 107972 1707
rect 108024 1698 109652 1707
rect 109704 1698 111332 1707
rect 111384 1698 113012 1707
rect 113064 1698 114692 1707
rect 114744 1698 116372 1707
rect 116424 1698 118052 1707
rect 118104 1698 119732 1707
rect 119784 1698 121412 1707
rect 121464 1698 123092 1707
rect 123144 1698 124772 1707
rect 124824 1698 126452 1707
rect 126504 1698 128132 1707
rect 128184 1698 129812 1707
rect 129864 1698 131492 1707
rect 131544 1698 133172 1707
rect 133224 1698 134984 1707
rect 1710 1612 134984 1698
<< via1 >>
rect 2132 81490 2184 81499
rect 3812 81490 3864 81499
rect 5492 81490 5544 81499
rect 7172 81490 7224 81499
rect 8852 81490 8904 81499
rect 10532 81490 10584 81499
rect 12212 81490 12264 81499
rect 13892 81490 13944 81499
rect 15572 81490 15624 81499
rect 17252 81490 17304 81499
rect 18932 81490 18984 81499
rect 20612 81490 20664 81499
rect 22292 81490 22344 81499
rect 23972 81490 24024 81499
rect 25652 81490 25704 81499
rect 27332 81490 27384 81499
rect 29012 81490 29064 81499
rect 30692 81490 30744 81499
rect 32372 81490 32424 81499
rect 34052 81490 34104 81499
rect 35732 81490 35784 81499
rect 37412 81490 37464 81499
rect 39092 81490 39144 81499
rect 40772 81490 40824 81499
rect 42452 81490 42504 81499
rect 44132 81490 44184 81499
rect 45812 81490 45864 81499
rect 47492 81490 47544 81499
rect 49172 81490 49224 81499
rect 50852 81490 50904 81499
rect 52532 81490 52584 81499
rect 54212 81490 54264 81499
rect 55892 81490 55944 81499
rect 57572 81490 57624 81499
rect 59252 81490 59304 81499
rect 60932 81490 60984 81499
rect 62612 81490 62664 81499
rect 64292 81490 64344 81499
rect 65972 81490 66024 81499
rect 67652 81490 67704 81499
rect 69332 81490 69384 81499
rect 71012 81490 71064 81499
rect 72692 81490 72744 81499
rect 74372 81490 74424 81499
rect 76052 81490 76104 81499
rect 77732 81490 77784 81499
rect 79412 81490 79464 81499
rect 81092 81490 81144 81499
rect 82772 81490 82824 81499
rect 84452 81490 84504 81499
rect 86132 81490 86184 81499
rect 87812 81490 87864 81499
rect 89492 81490 89544 81499
rect 91172 81490 91224 81499
rect 92852 81490 92904 81499
rect 94532 81490 94584 81499
rect 96212 81490 96264 81499
rect 97892 81490 97944 81499
rect 99572 81490 99624 81499
rect 101252 81490 101304 81499
rect 102932 81490 102984 81499
rect 104612 81490 104664 81499
rect 106292 81490 106344 81499
rect 107972 81490 108024 81499
rect 109652 81490 109704 81499
rect 111332 81490 111384 81499
rect 113012 81490 113064 81499
rect 114692 81490 114744 81499
rect 116372 81490 116424 81499
rect 118052 81490 118104 81499
rect 119732 81490 119784 81499
rect 121412 81490 121464 81499
rect 123092 81490 123144 81499
rect 124772 81490 124824 81499
rect 126452 81490 126504 81499
rect 128132 81490 128184 81499
rect 129812 81490 129864 81499
rect 131492 81490 131544 81499
rect 133172 81490 133224 81499
rect 2132 81456 2141 81490
rect 2141 81456 2175 81490
rect 2175 81456 2184 81490
rect 3812 81456 3821 81490
rect 3821 81456 3855 81490
rect 3855 81456 3864 81490
rect 5492 81456 5501 81490
rect 5501 81456 5535 81490
rect 5535 81456 5544 81490
rect 7172 81456 7181 81490
rect 7181 81456 7215 81490
rect 7215 81456 7224 81490
rect 8852 81456 8861 81490
rect 8861 81456 8895 81490
rect 8895 81456 8904 81490
rect 10532 81456 10541 81490
rect 10541 81456 10575 81490
rect 10575 81456 10584 81490
rect 12212 81456 12221 81490
rect 12221 81456 12255 81490
rect 12255 81456 12264 81490
rect 13892 81456 13901 81490
rect 13901 81456 13935 81490
rect 13935 81456 13944 81490
rect 15572 81456 15581 81490
rect 15581 81456 15615 81490
rect 15615 81456 15624 81490
rect 17252 81456 17261 81490
rect 17261 81456 17295 81490
rect 17295 81456 17304 81490
rect 18932 81456 18941 81490
rect 18941 81456 18975 81490
rect 18975 81456 18984 81490
rect 20612 81456 20621 81490
rect 20621 81456 20655 81490
rect 20655 81456 20664 81490
rect 22292 81456 22301 81490
rect 22301 81456 22335 81490
rect 22335 81456 22344 81490
rect 23972 81456 23981 81490
rect 23981 81456 24015 81490
rect 24015 81456 24024 81490
rect 25652 81456 25661 81490
rect 25661 81456 25695 81490
rect 25695 81456 25704 81490
rect 27332 81456 27341 81490
rect 27341 81456 27375 81490
rect 27375 81456 27384 81490
rect 29012 81456 29021 81490
rect 29021 81456 29055 81490
rect 29055 81456 29064 81490
rect 30692 81456 30701 81490
rect 30701 81456 30735 81490
rect 30735 81456 30744 81490
rect 32372 81456 32381 81490
rect 32381 81456 32415 81490
rect 32415 81456 32424 81490
rect 34052 81456 34061 81490
rect 34061 81456 34095 81490
rect 34095 81456 34104 81490
rect 35732 81456 35741 81490
rect 35741 81456 35775 81490
rect 35775 81456 35784 81490
rect 37412 81456 37421 81490
rect 37421 81456 37455 81490
rect 37455 81456 37464 81490
rect 39092 81456 39101 81490
rect 39101 81456 39135 81490
rect 39135 81456 39144 81490
rect 40772 81456 40781 81490
rect 40781 81456 40815 81490
rect 40815 81456 40824 81490
rect 42452 81456 42461 81490
rect 42461 81456 42495 81490
rect 42495 81456 42504 81490
rect 44132 81456 44141 81490
rect 44141 81456 44175 81490
rect 44175 81456 44184 81490
rect 45812 81456 45821 81490
rect 45821 81456 45855 81490
rect 45855 81456 45864 81490
rect 47492 81456 47501 81490
rect 47501 81456 47535 81490
rect 47535 81456 47544 81490
rect 49172 81456 49181 81490
rect 49181 81456 49215 81490
rect 49215 81456 49224 81490
rect 50852 81456 50861 81490
rect 50861 81456 50895 81490
rect 50895 81456 50904 81490
rect 52532 81456 52541 81490
rect 52541 81456 52575 81490
rect 52575 81456 52584 81490
rect 54212 81456 54221 81490
rect 54221 81456 54255 81490
rect 54255 81456 54264 81490
rect 55892 81456 55901 81490
rect 55901 81456 55935 81490
rect 55935 81456 55944 81490
rect 57572 81456 57581 81490
rect 57581 81456 57615 81490
rect 57615 81456 57624 81490
rect 59252 81456 59261 81490
rect 59261 81456 59295 81490
rect 59295 81456 59304 81490
rect 60932 81456 60941 81490
rect 60941 81456 60975 81490
rect 60975 81456 60984 81490
rect 62612 81456 62621 81490
rect 62621 81456 62655 81490
rect 62655 81456 62664 81490
rect 64292 81456 64301 81490
rect 64301 81456 64335 81490
rect 64335 81456 64344 81490
rect 65972 81456 65981 81490
rect 65981 81456 66015 81490
rect 66015 81456 66024 81490
rect 67652 81456 67661 81490
rect 67661 81456 67695 81490
rect 67695 81456 67704 81490
rect 69332 81456 69341 81490
rect 69341 81456 69375 81490
rect 69375 81456 69384 81490
rect 71012 81456 71021 81490
rect 71021 81456 71055 81490
rect 71055 81456 71064 81490
rect 72692 81456 72701 81490
rect 72701 81456 72735 81490
rect 72735 81456 72744 81490
rect 74372 81456 74381 81490
rect 74381 81456 74415 81490
rect 74415 81456 74424 81490
rect 76052 81456 76061 81490
rect 76061 81456 76095 81490
rect 76095 81456 76104 81490
rect 77732 81456 77741 81490
rect 77741 81456 77775 81490
rect 77775 81456 77784 81490
rect 79412 81456 79421 81490
rect 79421 81456 79455 81490
rect 79455 81456 79464 81490
rect 81092 81456 81101 81490
rect 81101 81456 81135 81490
rect 81135 81456 81144 81490
rect 82772 81456 82781 81490
rect 82781 81456 82815 81490
rect 82815 81456 82824 81490
rect 84452 81456 84461 81490
rect 84461 81456 84495 81490
rect 84495 81456 84504 81490
rect 86132 81456 86141 81490
rect 86141 81456 86175 81490
rect 86175 81456 86184 81490
rect 87812 81456 87821 81490
rect 87821 81456 87855 81490
rect 87855 81456 87864 81490
rect 89492 81456 89501 81490
rect 89501 81456 89535 81490
rect 89535 81456 89544 81490
rect 91172 81456 91181 81490
rect 91181 81456 91215 81490
rect 91215 81456 91224 81490
rect 92852 81456 92861 81490
rect 92861 81456 92895 81490
rect 92895 81456 92904 81490
rect 94532 81456 94541 81490
rect 94541 81456 94575 81490
rect 94575 81456 94584 81490
rect 96212 81456 96221 81490
rect 96221 81456 96255 81490
rect 96255 81456 96264 81490
rect 97892 81456 97901 81490
rect 97901 81456 97935 81490
rect 97935 81456 97944 81490
rect 99572 81456 99581 81490
rect 99581 81456 99615 81490
rect 99615 81456 99624 81490
rect 101252 81456 101261 81490
rect 101261 81456 101295 81490
rect 101295 81456 101304 81490
rect 102932 81456 102941 81490
rect 102941 81456 102975 81490
rect 102975 81456 102984 81490
rect 104612 81456 104621 81490
rect 104621 81456 104655 81490
rect 104655 81456 104664 81490
rect 106292 81456 106301 81490
rect 106301 81456 106335 81490
rect 106335 81456 106344 81490
rect 107972 81456 107981 81490
rect 107981 81456 108015 81490
rect 108015 81456 108024 81490
rect 109652 81456 109661 81490
rect 109661 81456 109695 81490
rect 109695 81456 109704 81490
rect 111332 81456 111341 81490
rect 111341 81456 111375 81490
rect 111375 81456 111384 81490
rect 113012 81456 113021 81490
rect 113021 81456 113055 81490
rect 113055 81456 113064 81490
rect 114692 81456 114701 81490
rect 114701 81456 114735 81490
rect 114735 81456 114744 81490
rect 116372 81456 116381 81490
rect 116381 81456 116415 81490
rect 116415 81456 116424 81490
rect 118052 81456 118061 81490
rect 118061 81456 118095 81490
rect 118095 81456 118104 81490
rect 119732 81456 119741 81490
rect 119741 81456 119775 81490
rect 119775 81456 119784 81490
rect 121412 81456 121421 81490
rect 121421 81456 121455 81490
rect 121455 81456 121464 81490
rect 123092 81456 123101 81490
rect 123101 81456 123135 81490
rect 123135 81456 123144 81490
rect 124772 81456 124781 81490
rect 124781 81456 124815 81490
rect 124815 81456 124824 81490
rect 126452 81456 126461 81490
rect 126461 81456 126495 81490
rect 126495 81456 126504 81490
rect 128132 81456 128141 81490
rect 128141 81456 128175 81490
rect 128175 81456 128184 81490
rect 129812 81456 129821 81490
rect 129821 81456 129855 81490
rect 129855 81456 129864 81490
rect 131492 81456 131501 81490
rect 131501 81456 131535 81490
rect 131535 81456 131544 81490
rect 133172 81456 133181 81490
rect 133181 81456 133215 81490
rect 133215 81456 133224 81490
rect 2132 81447 2184 81456
rect 3812 81447 3864 81456
rect 5492 81447 5544 81456
rect 7172 81447 7224 81456
rect 8852 81447 8904 81456
rect 10532 81447 10584 81456
rect 12212 81447 12264 81456
rect 13892 81447 13944 81456
rect 15572 81447 15624 81456
rect 17252 81447 17304 81456
rect 18932 81447 18984 81456
rect 20612 81447 20664 81456
rect 22292 81447 22344 81456
rect 23972 81447 24024 81456
rect 25652 81447 25704 81456
rect 27332 81447 27384 81456
rect 29012 81447 29064 81456
rect 30692 81447 30744 81456
rect 32372 81447 32424 81456
rect 34052 81447 34104 81456
rect 35732 81447 35784 81456
rect 37412 81447 37464 81456
rect 39092 81447 39144 81456
rect 40772 81447 40824 81456
rect 42452 81447 42504 81456
rect 44132 81447 44184 81456
rect 45812 81447 45864 81456
rect 47492 81447 47544 81456
rect 49172 81447 49224 81456
rect 50852 81447 50904 81456
rect 52532 81447 52584 81456
rect 54212 81447 54264 81456
rect 55892 81447 55944 81456
rect 57572 81447 57624 81456
rect 59252 81447 59304 81456
rect 60932 81447 60984 81456
rect 62612 81447 62664 81456
rect 64292 81447 64344 81456
rect 65972 81447 66024 81456
rect 67652 81447 67704 81456
rect 69332 81447 69384 81456
rect 71012 81447 71064 81456
rect 72692 81447 72744 81456
rect 74372 81447 74424 81456
rect 76052 81447 76104 81456
rect 77732 81447 77784 81456
rect 79412 81447 79464 81456
rect 81092 81447 81144 81456
rect 82772 81447 82824 81456
rect 84452 81447 84504 81456
rect 86132 81447 86184 81456
rect 87812 81447 87864 81456
rect 89492 81447 89544 81456
rect 91172 81447 91224 81456
rect 92852 81447 92904 81456
rect 94532 81447 94584 81456
rect 96212 81447 96264 81456
rect 97892 81447 97944 81456
rect 99572 81447 99624 81456
rect 101252 81447 101304 81456
rect 102932 81447 102984 81456
rect 104612 81447 104664 81456
rect 106292 81447 106344 81456
rect 107972 81447 108024 81456
rect 109652 81447 109704 81456
rect 111332 81447 111384 81456
rect 113012 81447 113064 81456
rect 114692 81447 114744 81456
rect 116372 81447 116424 81456
rect 118052 81447 118104 81456
rect 119732 81447 119784 81456
rect 121412 81447 121464 81456
rect 123092 81447 123144 81456
rect 124772 81447 124824 81456
rect 126452 81447 126504 81456
rect 128132 81447 128184 81456
rect 129812 81447 129864 81456
rect 131492 81447 131544 81456
rect 133172 81447 133224 81456
rect 1796 81037 1848 81046
rect 1796 81003 1805 81037
rect 1805 81003 1839 81037
rect 1839 81003 1848 81037
rect 1796 80994 1848 81003
rect 134846 81037 134898 81046
rect 134846 81003 134855 81037
rect 134855 81003 134889 81037
rect 134889 81003 134898 81037
rect 134846 80994 134898 81003
rect 1796 80701 1848 80710
rect 1796 80667 1805 80701
rect 1805 80667 1839 80701
rect 1839 80667 1848 80701
rect 1796 80658 1848 80667
rect 134846 80701 134898 80710
rect 134846 80667 134855 80701
rect 134855 80667 134889 80701
rect 134889 80667 134898 80701
rect 134846 80658 134898 80667
rect 1796 80365 1848 80374
rect 1796 80331 1805 80365
rect 1805 80331 1839 80365
rect 1839 80331 1848 80365
rect 1796 80322 1848 80331
rect 134846 80365 134898 80374
rect 134846 80331 134855 80365
rect 134855 80331 134889 80365
rect 134889 80331 134898 80365
rect 134846 80322 134898 80331
rect 1796 80029 1848 80038
rect 1796 79995 1805 80029
rect 1805 79995 1839 80029
rect 1839 79995 1848 80029
rect 1796 79986 1848 79995
rect 134846 80029 134898 80038
rect 134846 79995 134855 80029
rect 134855 79995 134889 80029
rect 134889 79995 134898 80029
rect 134846 79986 134898 79995
rect 1796 79693 1848 79702
rect 1796 79659 1805 79693
rect 1805 79659 1839 79693
rect 1839 79659 1848 79693
rect 1796 79650 1848 79659
rect 134846 79693 134898 79702
rect 134846 79659 134855 79693
rect 134855 79659 134889 79693
rect 134889 79659 134898 79693
rect 134846 79650 134898 79659
rect 1796 79357 1848 79366
rect 1796 79323 1805 79357
rect 1805 79323 1839 79357
rect 1839 79323 1848 79357
rect 1796 79314 1848 79323
rect 134846 79357 134898 79366
rect 134846 79323 134855 79357
rect 134855 79323 134889 79357
rect 134889 79323 134898 79357
rect 134846 79314 134898 79323
rect 1796 79021 1848 79030
rect 1796 78987 1805 79021
rect 1805 78987 1839 79021
rect 1839 78987 1848 79021
rect 1796 78978 1848 78987
rect 134846 79021 134898 79030
rect 134846 78987 134855 79021
rect 134855 78987 134889 79021
rect 134889 78987 134898 79021
rect 134846 78978 134898 78987
rect 1796 78685 1848 78694
rect 1796 78651 1805 78685
rect 1805 78651 1839 78685
rect 1839 78651 1848 78685
rect 1796 78642 1848 78651
rect 134846 78685 134898 78694
rect 134846 78651 134855 78685
rect 134855 78651 134889 78685
rect 134889 78651 134898 78685
rect 134846 78642 134898 78651
rect 1796 78349 1848 78358
rect 1796 78315 1805 78349
rect 1805 78315 1839 78349
rect 1839 78315 1848 78349
rect 1796 78306 1848 78315
rect 134846 78349 134898 78358
rect 134846 78315 134855 78349
rect 134855 78315 134889 78349
rect 134889 78315 134898 78349
rect 134846 78306 134898 78315
rect 1796 78013 1848 78022
rect 1796 77979 1805 78013
rect 1805 77979 1839 78013
rect 1839 77979 1848 78013
rect 1796 77970 1848 77979
rect 134846 78013 134898 78022
rect 134846 77979 134855 78013
rect 134855 77979 134889 78013
rect 134889 77979 134898 78013
rect 134846 77970 134898 77979
rect 1796 77677 1848 77686
rect 1796 77643 1805 77677
rect 1805 77643 1839 77677
rect 1839 77643 1848 77677
rect 1796 77634 1848 77643
rect 134846 77677 134898 77686
rect 134846 77643 134855 77677
rect 134855 77643 134889 77677
rect 134889 77643 134898 77677
rect 134846 77634 134898 77643
rect 1796 77341 1848 77350
rect 1796 77307 1805 77341
rect 1805 77307 1839 77341
rect 1839 77307 1848 77341
rect 1796 77298 1848 77307
rect 134846 77341 134898 77350
rect 134846 77307 134855 77341
rect 134855 77307 134889 77341
rect 134889 77307 134898 77341
rect 134846 77298 134898 77307
rect 1796 77005 1848 77014
rect 1796 76971 1805 77005
rect 1805 76971 1839 77005
rect 1839 76971 1848 77005
rect 1796 76962 1848 76971
rect 28620 76993 28672 77045
rect 31116 76993 31168 77045
rect 33612 76993 33664 77045
rect 36108 76993 36160 77045
rect 38604 76993 38656 77045
rect 41100 76993 41152 77045
rect 43596 76993 43648 77045
rect 46092 76993 46144 77045
rect 48588 76993 48640 77045
rect 51084 76993 51136 77045
rect 53580 76993 53632 77045
rect 56076 76993 56128 77045
rect 58572 76993 58624 77045
rect 61068 76993 61120 77045
rect 63564 76993 63616 77045
rect 66060 76993 66112 77045
rect 68556 76993 68608 77045
rect 71052 76993 71104 77045
rect 73548 76993 73600 77045
rect 76044 76993 76096 77045
rect 78540 76993 78592 77045
rect 81036 76993 81088 77045
rect 83532 76993 83584 77045
rect 86028 76993 86080 77045
rect 88524 76993 88576 77045
rect 91020 76993 91072 77045
rect 93516 76993 93568 77045
rect 96012 76993 96064 77045
rect 98508 76993 98560 77045
rect 101004 76993 101056 77045
rect 103500 76993 103552 77045
rect 105996 76993 106048 77045
rect 134846 77005 134898 77014
rect 134846 76971 134855 77005
rect 134855 76971 134889 77005
rect 134889 76971 134898 77005
rect 134846 76962 134898 76971
rect 1796 76669 1848 76678
rect 1796 76635 1805 76669
rect 1805 76635 1839 76669
rect 1839 76635 1848 76669
rect 1796 76626 1848 76635
rect 134846 76669 134898 76678
rect 134846 76635 134855 76669
rect 134855 76635 134889 76669
rect 134889 76635 134898 76669
rect 134846 76626 134898 76635
rect 1796 76333 1848 76342
rect 1796 76299 1805 76333
rect 1805 76299 1839 76333
rect 1839 76299 1848 76333
rect 1796 76290 1848 76299
rect 134846 76333 134898 76342
rect 134846 76299 134855 76333
rect 134855 76299 134889 76333
rect 134889 76299 134898 76333
rect 134846 76290 134898 76299
rect 1796 75997 1848 76006
rect 1796 75963 1805 75997
rect 1805 75963 1839 75997
rect 1839 75963 1848 75997
rect 1796 75954 1848 75963
rect 134846 75997 134898 76006
rect 134846 75963 134855 75997
rect 134855 75963 134889 75997
rect 134889 75963 134898 75997
rect 134846 75954 134898 75963
rect 1796 75661 1848 75670
rect 1796 75627 1805 75661
rect 1805 75627 1839 75661
rect 1839 75627 1848 75661
rect 1796 75618 1848 75627
rect 134846 75661 134898 75670
rect 134846 75627 134855 75661
rect 134855 75627 134889 75661
rect 134889 75627 134898 75661
rect 134846 75618 134898 75627
rect 1796 75325 1848 75334
rect 1796 75291 1805 75325
rect 1805 75291 1839 75325
rect 1839 75291 1848 75325
rect 1796 75282 1848 75291
rect 134846 75325 134898 75334
rect 134846 75291 134855 75325
rect 134855 75291 134889 75325
rect 134889 75291 134898 75325
rect 134846 75282 134898 75291
rect 1796 74989 1848 74998
rect 1796 74955 1805 74989
rect 1805 74955 1839 74989
rect 1839 74955 1848 74989
rect 1796 74946 1848 74955
rect 134846 74989 134898 74998
rect 134846 74955 134855 74989
rect 134855 74955 134889 74989
rect 134889 74955 134898 74989
rect 134846 74946 134898 74955
rect 1796 74653 1848 74662
rect 1796 74619 1805 74653
rect 1805 74619 1839 74653
rect 1839 74619 1848 74653
rect 1796 74610 1848 74619
rect 134846 74653 134898 74662
rect 134846 74619 134855 74653
rect 134855 74619 134889 74653
rect 134889 74619 134898 74653
rect 134846 74610 134898 74619
rect 1796 74317 1848 74326
rect 1796 74283 1805 74317
rect 1805 74283 1839 74317
rect 1839 74283 1848 74317
rect 1796 74274 1848 74283
rect 134846 74317 134898 74326
rect 134846 74283 134855 74317
rect 134855 74283 134889 74317
rect 134889 74283 134898 74317
rect 134846 74274 134898 74283
rect 1796 73981 1848 73990
rect 1796 73947 1805 73981
rect 1805 73947 1839 73981
rect 1839 73947 1848 73981
rect 1796 73938 1848 73947
rect 134846 73981 134898 73990
rect 134846 73947 134855 73981
rect 134855 73947 134889 73981
rect 134889 73947 134898 73981
rect 134846 73938 134898 73947
rect 1796 73645 1848 73654
rect 1796 73611 1805 73645
rect 1805 73611 1839 73645
rect 1839 73611 1848 73645
rect 1796 73602 1848 73611
rect 134846 73645 134898 73654
rect 134846 73611 134855 73645
rect 134855 73611 134889 73645
rect 134889 73611 134898 73645
rect 134846 73602 134898 73611
rect 1796 73309 1848 73318
rect 1796 73275 1805 73309
rect 1805 73275 1839 73309
rect 1839 73275 1848 73309
rect 1796 73266 1848 73275
rect 134846 73309 134898 73318
rect 134846 73275 134855 73309
rect 134855 73275 134889 73309
rect 134889 73275 134898 73309
rect 134846 73266 134898 73275
rect 1796 72973 1848 72982
rect 1796 72939 1805 72973
rect 1805 72939 1839 72973
rect 1839 72939 1848 72973
rect 1796 72930 1848 72939
rect 134846 72973 134898 72982
rect 134846 72939 134855 72973
rect 134855 72939 134889 72973
rect 134889 72939 134898 72973
rect 134846 72930 134898 72939
rect 1796 72637 1848 72646
rect 1796 72603 1805 72637
rect 1805 72603 1839 72637
rect 1839 72603 1848 72637
rect 1796 72594 1848 72603
rect 134846 72637 134898 72646
rect 134846 72603 134855 72637
rect 134855 72603 134889 72637
rect 134889 72603 134898 72637
rect 134846 72594 134898 72603
rect 1796 72301 1848 72310
rect 1796 72267 1805 72301
rect 1805 72267 1839 72301
rect 1839 72267 1848 72301
rect 1796 72258 1848 72267
rect 134846 72301 134898 72310
rect 134846 72267 134855 72301
rect 134855 72267 134889 72301
rect 134889 72267 134898 72301
rect 134846 72258 134898 72267
rect 1796 71965 1848 71974
rect 1796 71931 1805 71965
rect 1805 71931 1839 71965
rect 1839 71931 1848 71965
rect 1796 71922 1848 71931
rect 134846 71965 134898 71974
rect 134846 71931 134855 71965
rect 134855 71931 134889 71965
rect 134889 71931 134898 71965
rect 134846 71922 134898 71931
rect 1796 71629 1848 71638
rect 1796 71595 1805 71629
rect 1805 71595 1839 71629
rect 1839 71595 1848 71629
rect 1796 71586 1848 71595
rect 134846 71629 134898 71638
rect 134846 71595 134855 71629
rect 134855 71595 134889 71629
rect 134889 71595 134898 71629
rect 134846 71586 134898 71595
rect 1796 71293 1848 71302
rect 1796 71259 1805 71293
rect 1805 71259 1839 71293
rect 1839 71259 1848 71293
rect 1796 71250 1848 71259
rect 134846 71293 134898 71302
rect 134846 71259 134855 71293
rect 134855 71259 134889 71293
rect 134889 71259 134898 71293
rect 134846 71250 134898 71259
rect 1796 70957 1848 70966
rect 1796 70923 1805 70957
rect 1805 70923 1839 70957
rect 1839 70923 1848 70957
rect 1796 70914 1848 70923
rect 134846 70957 134898 70966
rect 134846 70923 134855 70957
rect 134855 70923 134889 70957
rect 134889 70923 134898 70957
rect 134846 70914 134898 70923
rect 1796 70621 1848 70630
rect 1796 70587 1805 70621
rect 1805 70587 1839 70621
rect 1839 70587 1848 70621
rect 1796 70578 1848 70587
rect 134846 70621 134898 70630
rect 134846 70587 134855 70621
rect 134855 70587 134889 70621
rect 134889 70587 134898 70621
rect 134846 70578 134898 70587
rect 1796 70285 1848 70294
rect 1796 70251 1805 70285
rect 1805 70251 1839 70285
rect 1839 70251 1848 70285
rect 1796 70242 1848 70251
rect 134846 70285 134898 70294
rect 134846 70251 134855 70285
rect 134855 70251 134889 70285
rect 134889 70251 134898 70285
rect 134846 70242 134898 70251
rect 1796 69949 1848 69958
rect 1796 69915 1805 69949
rect 1805 69915 1839 69949
rect 1839 69915 1848 69949
rect 1796 69906 1848 69915
rect 134846 69949 134898 69958
rect 134846 69915 134855 69949
rect 134855 69915 134889 69949
rect 134889 69915 134898 69949
rect 134846 69906 134898 69915
rect 1796 69613 1848 69622
rect 1796 69579 1805 69613
rect 1805 69579 1839 69613
rect 1839 69579 1848 69613
rect 1796 69570 1848 69579
rect 134846 69613 134898 69622
rect 134846 69579 134855 69613
rect 134855 69579 134889 69613
rect 134889 69579 134898 69613
rect 134846 69570 134898 69579
rect 1796 69277 1848 69286
rect 1796 69243 1805 69277
rect 1805 69243 1839 69277
rect 1839 69243 1848 69277
rect 1796 69234 1848 69243
rect 134846 69277 134898 69286
rect 134846 69243 134855 69277
rect 134855 69243 134889 69277
rect 134889 69243 134898 69277
rect 134846 69234 134898 69243
rect 1796 68941 1848 68950
rect 1796 68907 1805 68941
rect 1805 68907 1839 68941
rect 1839 68907 1848 68941
rect 1796 68898 1848 68907
rect 134846 68941 134898 68950
rect 134846 68907 134855 68941
rect 134855 68907 134889 68941
rect 134889 68907 134898 68941
rect 134846 68898 134898 68907
rect 1796 68605 1848 68614
rect 1796 68571 1805 68605
rect 1805 68571 1839 68605
rect 1839 68571 1848 68605
rect 1796 68562 1848 68571
rect 134846 68605 134898 68614
rect 134846 68571 134855 68605
rect 134855 68571 134889 68605
rect 134889 68571 134898 68605
rect 134846 68562 134898 68571
rect 1796 68269 1848 68278
rect 1796 68235 1805 68269
rect 1805 68235 1839 68269
rect 1839 68235 1848 68269
rect 1796 68226 1848 68235
rect 134846 68269 134898 68278
rect 134846 68235 134855 68269
rect 134855 68235 134889 68269
rect 134889 68235 134898 68269
rect 134846 68226 134898 68235
rect 1796 67933 1848 67942
rect 1796 67899 1805 67933
rect 1805 67899 1839 67933
rect 1839 67899 1848 67933
rect 1796 67890 1848 67899
rect 134846 67933 134898 67942
rect 134846 67899 134855 67933
rect 134855 67899 134889 67933
rect 134889 67899 134898 67933
rect 134846 67890 134898 67899
rect 1796 67597 1848 67606
rect 1796 67563 1805 67597
rect 1805 67563 1839 67597
rect 1839 67563 1848 67597
rect 1796 67554 1848 67563
rect 134846 67597 134898 67606
rect 134846 67563 134855 67597
rect 134855 67563 134889 67597
rect 134889 67563 134898 67597
rect 134846 67554 134898 67563
rect 1796 67261 1848 67270
rect 1796 67227 1805 67261
rect 1805 67227 1839 67261
rect 1839 67227 1848 67261
rect 1796 67218 1848 67227
rect 134846 67261 134898 67270
rect 134846 67227 134855 67261
rect 134855 67227 134889 67261
rect 134889 67227 134898 67261
rect 134846 67218 134898 67227
rect 1796 66925 1848 66934
rect 1796 66891 1805 66925
rect 1805 66891 1839 66925
rect 1839 66891 1848 66925
rect 1796 66882 1848 66891
rect 134846 66925 134898 66934
rect 134846 66891 134855 66925
rect 134855 66891 134889 66925
rect 134889 66891 134898 66925
rect 134846 66882 134898 66891
rect 1796 66589 1848 66598
rect 1796 66555 1805 66589
rect 1805 66555 1839 66589
rect 1839 66555 1848 66589
rect 1796 66546 1848 66555
rect 134846 66589 134898 66598
rect 134846 66555 134855 66589
rect 134855 66555 134889 66589
rect 134889 66555 134898 66589
rect 134846 66546 134898 66555
rect 1796 66253 1848 66262
rect 1796 66219 1805 66253
rect 1805 66219 1839 66253
rect 1839 66219 1848 66253
rect 1796 66210 1848 66219
rect 134846 66253 134898 66262
rect 134846 66219 134855 66253
rect 134855 66219 134889 66253
rect 134889 66219 134898 66253
rect 134846 66210 134898 66219
rect 1796 65917 1848 65926
rect 1796 65883 1805 65917
rect 1805 65883 1839 65917
rect 1839 65883 1848 65917
rect 1796 65874 1848 65883
rect 134846 65917 134898 65926
rect 134846 65883 134855 65917
rect 134855 65883 134889 65917
rect 134889 65883 134898 65917
rect 134846 65874 134898 65883
rect 1796 65581 1848 65590
rect 1796 65547 1805 65581
rect 1805 65547 1839 65581
rect 1839 65547 1848 65581
rect 1796 65538 1848 65547
rect 134846 65581 134898 65590
rect 134846 65547 134855 65581
rect 134855 65547 134889 65581
rect 134889 65547 134898 65581
rect 134846 65538 134898 65547
rect 1796 65245 1848 65254
rect 1796 65211 1805 65245
rect 1805 65211 1839 65245
rect 1839 65211 1848 65245
rect 1796 65202 1848 65211
rect 134846 65245 134898 65254
rect 134846 65211 134855 65245
rect 134855 65211 134889 65245
rect 134889 65211 134898 65245
rect 134846 65202 134898 65211
rect 1796 64909 1848 64918
rect 1796 64875 1805 64909
rect 1805 64875 1839 64909
rect 1839 64875 1848 64909
rect 1796 64866 1848 64875
rect 134846 64909 134898 64918
rect 134846 64875 134855 64909
rect 134855 64875 134889 64909
rect 134889 64875 134898 64909
rect 134846 64866 134898 64875
rect 1796 64573 1848 64582
rect 1796 64539 1805 64573
rect 1805 64539 1839 64573
rect 1839 64539 1848 64573
rect 1796 64530 1848 64539
rect 134846 64573 134898 64582
rect 134846 64539 134855 64573
rect 134855 64539 134889 64573
rect 134889 64539 134898 64573
rect 134846 64530 134898 64539
rect 1796 64237 1848 64246
rect 1796 64203 1805 64237
rect 1805 64203 1839 64237
rect 1839 64203 1848 64237
rect 1796 64194 1848 64203
rect 134846 64237 134898 64246
rect 134846 64203 134855 64237
rect 134855 64203 134889 64237
rect 134889 64203 134898 64237
rect 134846 64194 134898 64203
rect 1796 63901 1848 63910
rect 1796 63867 1805 63901
rect 1805 63867 1839 63901
rect 1839 63867 1848 63901
rect 1796 63858 1848 63867
rect 134846 63901 134898 63910
rect 134846 63867 134855 63901
rect 134855 63867 134889 63901
rect 134889 63867 134898 63901
rect 134846 63858 134898 63867
rect 1796 63565 1848 63574
rect 1796 63531 1805 63565
rect 1805 63531 1839 63565
rect 1839 63531 1848 63565
rect 1796 63522 1848 63531
rect 134846 63565 134898 63574
rect 134846 63531 134855 63565
rect 134855 63531 134889 63565
rect 134889 63531 134898 63565
rect 134846 63522 134898 63531
rect 1796 63229 1848 63238
rect 1796 63195 1805 63229
rect 1805 63195 1839 63229
rect 1839 63195 1848 63229
rect 1796 63186 1848 63195
rect 134846 63229 134898 63238
rect 134846 63195 134855 63229
rect 134855 63195 134889 63229
rect 134889 63195 134898 63229
rect 134846 63186 134898 63195
rect 1796 62893 1848 62902
rect 1796 62859 1805 62893
rect 1805 62859 1839 62893
rect 1839 62859 1848 62893
rect 1796 62850 1848 62859
rect 134846 62893 134898 62902
rect 134846 62859 134855 62893
rect 134855 62859 134889 62893
rect 134889 62859 134898 62893
rect 134846 62850 134898 62859
rect 1796 62557 1848 62566
rect 1796 62523 1805 62557
rect 1805 62523 1839 62557
rect 1839 62523 1848 62557
rect 1796 62514 1848 62523
rect 134846 62557 134898 62566
rect 134846 62523 134855 62557
rect 134855 62523 134889 62557
rect 134889 62523 134898 62557
rect 134846 62514 134898 62523
rect 1796 62221 1848 62230
rect 1796 62187 1805 62221
rect 1805 62187 1839 62221
rect 1839 62187 1848 62221
rect 1796 62178 1848 62187
rect 134846 62221 134898 62230
rect 134846 62187 134855 62221
rect 134855 62187 134889 62221
rect 134889 62187 134898 62221
rect 134846 62178 134898 62187
rect 1796 61885 1848 61894
rect 1796 61851 1805 61885
rect 1805 61851 1839 61885
rect 1839 61851 1848 61885
rect 1796 61842 1848 61851
rect 134846 61885 134898 61894
rect 134846 61851 134855 61885
rect 134855 61851 134889 61885
rect 134889 61851 134898 61885
rect 134846 61842 134898 61851
rect 1796 61549 1848 61558
rect 1796 61515 1805 61549
rect 1805 61515 1839 61549
rect 1839 61515 1848 61549
rect 1796 61506 1848 61515
rect 134846 61549 134898 61558
rect 134846 61515 134855 61549
rect 134855 61515 134889 61549
rect 134889 61515 134898 61549
rect 134846 61506 134898 61515
rect 1796 61213 1848 61222
rect 1796 61179 1805 61213
rect 1805 61179 1839 61213
rect 1839 61179 1848 61213
rect 1796 61170 1848 61179
rect 134846 61213 134898 61222
rect 134846 61179 134855 61213
rect 134855 61179 134889 61213
rect 134889 61179 134898 61213
rect 134846 61170 134898 61179
rect 1796 60877 1848 60886
rect 1796 60843 1805 60877
rect 1805 60843 1839 60877
rect 1839 60843 1848 60877
rect 1796 60834 1848 60843
rect 134846 60877 134898 60886
rect 134846 60843 134855 60877
rect 134855 60843 134889 60877
rect 134889 60843 134898 60877
rect 134846 60834 134898 60843
rect 1796 60541 1848 60550
rect 1796 60507 1805 60541
rect 1805 60507 1839 60541
rect 1839 60507 1848 60541
rect 1796 60498 1848 60507
rect 134846 60541 134898 60550
rect 134846 60507 134855 60541
rect 134855 60507 134889 60541
rect 134889 60507 134898 60541
rect 134846 60498 134898 60507
rect 1796 60205 1848 60214
rect 1796 60171 1805 60205
rect 1805 60171 1839 60205
rect 1839 60171 1848 60205
rect 1796 60162 1848 60171
rect 134846 60205 134898 60214
rect 134846 60171 134855 60205
rect 134855 60171 134889 60205
rect 134889 60171 134898 60205
rect 134846 60162 134898 60171
rect 1796 59869 1848 59878
rect 1796 59835 1805 59869
rect 1805 59835 1839 59869
rect 1839 59835 1848 59869
rect 1796 59826 1848 59835
rect 134846 59869 134898 59878
rect 134846 59835 134855 59869
rect 134855 59835 134889 59869
rect 134889 59835 134898 59869
rect 134846 59826 134898 59835
rect 1796 59533 1848 59542
rect 1796 59499 1805 59533
rect 1805 59499 1839 59533
rect 1839 59499 1848 59533
rect 1796 59490 1848 59499
rect 134846 59533 134898 59542
rect 134846 59499 134855 59533
rect 134855 59499 134889 59533
rect 134889 59499 134898 59533
rect 134846 59490 134898 59499
rect 1796 59197 1848 59206
rect 1796 59163 1805 59197
rect 1805 59163 1839 59197
rect 1839 59163 1848 59197
rect 1796 59154 1848 59163
rect 134846 59197 134898 59206
rect 134846 59163 134855 59197
rect 134855 59163 134889 59197
rect 134889 59163 134898 59197
rect 134846 59154 134898 59163
rect 1796 58861 1848 58870
rect 1796 58827 1805 58861
rect 1805 58827 1839 58861
rect 1839 58827 1848 58861
rect 1796 58818 1848 58827
rect 134846 58861 134898 58870
rect 134846 58827 134855 58861
rect 134855 58827 134889 58861
rect 134889 58827 134898 58861
rect 134846 58818 134898 58827
rect 1796 58525 1848 58534
rect 1796 58491 1805 58525
rect 1805 58491 1839 58525
rect 1839 58491 1848 58525
rect 1796 58482 1848 58491
rect 134846 58525 134898 58534
rect 134846 58491 134855 58525
rect 134855 58491 134889 58525
rect 134889 58491 134898 58525
rect 134846 58482 134898 58491
rect 1796 58189 1848 58198
rect 1796 58155 1805 58189
rect 1805 58155 1839 58189
rect 1839 58155 1848 58189
rect 1796 58146 1848 58155
rect 134846 58189 134898 58198
rect 134846 58155 134855 58189
rect 134855 58155 134889 58189
rect 134889 58155 134898 58189
rect 134846 58146 134898 58155
rect 1796 57853 1848 57862
rect 1796 57819 1805 57853
rect 1805 57819 1839 57853
rect 1839 57819 1848 57853
rect 1796 57810 1848 57819
rect 134846 57853 134898 57862
rect 134846 57819 134855 57853
rect 134855 57819 134889 57853
rect 134889 57819 134898 57853
rect 134846 57810 134898 57819
rect 1796 57517 1848 57526
rect 1796 57483 1805 57517
rect 1805 57483 1839 57517
rect 1839 57483 1848 57517
rect 1796 57474 1848 57483
rect 134846 57517 134898 57526
rect 134846 57483 134855 57517
rect 134855 57483 134889 57517
rect 134889 57483 134898 57517
rect 134846 57474 134898 57483
rect 1796 57181 1848 57190
rect 1796 57147 1805 57181
rect 1805 57147 1839 57181
rect 1839 57147 1848 57181
rect 1796 57138 1848 57147
rect 134846 57181 134898 57190
rect 134846 57147 134855 57181
rect 134855 57147 134889 57181
rect 134889 57147 134898 57181
rect 134846 57138 134898 57147
rect 1796 56845 1848 56854
rect 1796 56811 1805 56845
rect 1805 56811 1839 56845
rect 1839 56811 1848 56845
rect 1796 56802 1848 56811
rect 134846 56845 134898 56854
rect 134846 56811 134855 56845
rect 134855 56811 134889 56845
rect 134889 56811 134898 56845
rect 134846 56802 134898 56811
rect 1796 56509 1848 56518
rect 1796 56475 1805 56509
rect 1805 56475 1839 56509
rect 1839 56475 1848 56509
rect 1796 56466 1848 56475
rect 134846 56509 134898 56518
rect 134846 56475 134855 56509
rect 134855 56475 134889 56509
rect 134889 56475 134898 56509
rect 134846 56466 134898 56475
rect 1796 56173 1848 56182
rect 1796 56139 1805 56173
rect 1805 56139 1839 56173
rect 1839 56139 1848 56173
rect 1796 56130 1848 56139
rect 134846 56173 134898 56182
rect 134846 56139 134855 56173
rect 134855 56139 134889 56173
rect 134889 56139 134898 56173
rect 134846 56130 134898 56139
rect 1796 55837 1848 55846
rect 1796 55803 1805 55837
rect 1805 55803 1839 55837
rect 1839 55803 1848 55837
rect 1796 55794 1848 55803
rect 134846 55837 134898 55846
rect 134846 55803 134855 55837
rect 134855 55803 134889 55837
rect 134889 55803 134898 55837
rect 134846 55794 134898 55803
rect 1796 55501 1848 55510
rect 1796 55467 1805 55501
rect 1805 55467 1839 55501
rect 1839 55467 1848 55501
rect 1796 55458 1848 55467
rect 134846 55501 134898 55510
rect 134846 55467 134855 55501
rect 134855 55467 134889 55501
rect 134889 55467 134898 55501
rect 134846 55458 134898 55467
rect 1796 55165 1848 55174
rect 1796 55131 1805 55165
rect 1805 55131 1839 55165
rect 1839 55131 1848 55165
rect 1796 55122 1848 55131
rect 134846 55165 134898 55174
rect 134846 55131 134855 55165
rect 134855 55131 134889 55165
rect 134889 55131 134898 55165
rect 134846 55122 134898 55131
rect 1796 54829 1848 54838
rect 1796 54795 1805 54829
rect 1805 54795 1839 54829
rect 1839 54795 1848 54829
rect 1796 54786 1848 54795
rect 134846 54829 134898 54838
rect 134846 54795 134855 54829
rect 134855 54795 134889 54829
rect 134889 54795 134898 54829
rect 134846 54786 134898 54795
rect 1796 54493 1848 54502
rect 1796 54459 1805 54493
rect 1805 54459 1839 54493
rect 1839 54459 1848 54493
rect 1796 54450 1848 54459
rect 134846 54493 134898 54502
rect 134846 54459 134855 54493
rect 134855 54459 134889 54493
rect 134889 54459 134898 54493
rect 134846 54450 134898 54459
rect 1796 54157 1848 54166
rect 1796 54123 1805 54157
rect 1805 54123 1839 54157
rect 1839 54123 1848 54157
rect 1796 54114 1848 54123
rect 134846 54157 134898 54166
rect 134846 54123 134855 54157
rect 134855 54123 134889 54157
rect 134889 54123 134898 54157
rect 134846 54114 134898 54123
rect 1796 53821 1848 53830
rect 1796 53787 1805 53821
rect 1805 53787 1839 53821
rect 1839 53787 1848 53821
rect 1796 53778 1848 53787
rect 134846 53821 134898 53830
rect 134846 53787 134855 53821
rect 134855 53787 134889 53821
rect 134889 53787 134898 53821
rect 134846 53778 134898 53787
rect 1796 53485 1848 53494
rect 1796 53451 1805 53485
rect 1805 53451 1839 53485
rect 1839 53451 1848 53485
rect 1796 53442 1848 53451
rect 134846 53485 134898 53494
rect 134846 53451 134855 53485
rect 134855 53451 134889 53485
rect 134889 53451 134898 53485
rect 134846 53442 134898 53451
rect 1796 53149 1848 53158
rect 1796 53115 1805 53149
rect 1805 53115 1839 53149
rect 1839 53115 1848 53149
rect 1796 53106 1848 53115
rect 134846 53149 134898 53158
rect 134846 53115 134855 53149
rect 134855 53115 134889 53149
rect 134889 53115 134898 53149
rect 134846 53106 134898 53115
rect 1796 52813 1848 52822
rect 1796 52779 1805 52813
rect 1805 52779 1839 52813
rect 1839 52779 1848 52813
rect 1796 52770 1848 52779
rect 134846 52813 134898 52822
rect 134846 52779 134855 52813
rect 134855 52779 134889 52813
rect 134889 52779 134898 52813
rect 134846 52770 134898 52779
rect 1796 52477 1848 52486
rect 1796 52443 1805 52477
rect 1805 52443 1839 52477
rect 1839 52443 1848 52477
rect 1796 52434 1848 52443
rect 134846 52477 134898 52486
rect 134846 52443 134855 52477
rect 134855 52443 134889 52477
rect 134889 52443 134898 52477
rect 134846 52434 134898 52443
rect 1796 52141 1848 52150
rect 1796 52107 1805 52141
rect 1805 52107 1839 52141
rect 1839 52107 1848 52141
rect 1796 52098 1848 52107
rect 134846 52141 134898 52150
rect 134846 52107 134855 52141
rect 134855 52107 134889 52141
rect 134889 52107 134898 52141
rect 134846 52098 134898 52107
rect 1796 51805 1848 51814
rect 1796 51771 1805 51805
rect 1805 51771 1839 51805
rect 1839 51771 1848 51805
rect 1796 51762 1848 51771
rect 134846 51805 134898 51814
rect 134846 51771 134855 51805
rect 134855 51771 134889 51805
rect 134889 51771 134898 51805
rect 134846 51762 134898 51771
rect 1796 51469 1848 51478
rect 1796 51435 1805 51469
rect 1805 51435 1839 51469
rect 1839 51435 1848 51469
rect 1796 51426 1848 51435
rect 134846 51469 134898 51478
rect 134846 51435 134855 51469
rect 134855 51435 134889 51469
rect 134889 51435 134898 51469
rect 134846 51426 134898 51435
rect 1796 51133 1848 51142
rect 1796 51099 1805 51133
rect 1805 51099 1839 51133
rect 1839 51099 1848 51133
rect 1796 51090 1848 51099
rect 134846 51133 134898 51142
rect 134846 51099 134855 51133
rect 134855 51099 134889 51133
rect 134889 51099 134898 51133
rect 134846 51090 134898 51099
rect 1796 50797 1848 50806
rect 1796 50763 1805 50797
rect 1805 50763 1839 50797
rect 1839 50763 1848 50797
rect 1796 50754 1848 50763
rect 134846 50797 134898 50806
rect 134846 50763 134855 50797
rect 134855 50763 134889 50797
rect 134889 50763 134898 50797
rect 134846 50754 134898 50763
rect 1796 50461 1848 50470
rect 1796 50427 1805 50461
rect 1805 50427 1839 50461
rect 1839 50427 1848 50461
rect 1796 50418 1848 50427
rect 134846 50461 134898 50470
rect 134846 50427 134855 50461
rect 134855 50427 134889 50461
rect 134889 50427 134898 50461
rect 134846 50418 134898 50427
rect 1796 50125 1848 50134
rect 1796 50091 1805 50125
rect 1805 50091 1839 50125
rect 1839 50091 1848 50125
rect 1796 50082 1848 50091
rect 134846 50125 134898 50134
rect 134846 50091 134855 50125
rect 134855 50091 134889 50125
rect 134889 50091 134898 50125
rect 134846 50082 134898 50091
rect 1796 49789 1848 49798
rect 1796 49755 1805 49789
rect 1805 49755 1839 49789
rect 1839 49755 1848 49789
rect 1796 49746 1848 49755
rect 134846 49789 134898 49798
rect 134846 49755 134855 49789
rect 134855 49755 134889 49789
rect 134889 49755 134898 49789
rect 134846 49746 134898 49755
rect 1796 49453 1848 49462
rect 1796 49419 1805 49453
rect 1805 49419 1839 49453
rect 1839 49419 1848 49453
rect 1796 49410 1848 49419
rect 134846 49453 134898 49462
rect 134846 49419 134855 49453
rect 134855 49419 134889 49453
rect 134889 49419 134898 49453
rect 134846 49410 134898 49419
rect 1796 49117 1848 49126
rect 1796 49083 1805 49117
rect 1805 49083 1839 49117
rect 1839 49083 1848 49117
rect 1796 49074 1848 49083
rect 134846 49117 134898 49126
rect 134846 49083 134855 49117
rect 134855 49083 134889 49117
rect 134889 49083 134898 49117
rect 134846 49074 134898 49083
rect 1796 48781 1848 48790
rect 1796 48747 1805 48781
rect 1805 48747 1839 48781
rect 1839 48747 1848 48781
rect 1796 48738 1848 48747
rect 134846 48781 134898 48790
rect 134846 48747 134855 48781
rect 134855 48747 134889 48781
rect 134889 48747 134898 48781
rect 134846 48738 134898 48747
rect 1796 48445 1848 48454
rect 1796 48411 1805 48445
rect 1805 48411 1839 48445
rect 1839 48411 1848 48445
rect 1796 48402 1848 48411
rect 134846 48445 134898 48454
rect 134846 48411 134855 48445
rect 134855 48411 134889 48445
rect 134889 48411 134898 48445
rect 134846 48402 134898 48411
rect 1796 48109 1848 48118
rect 1796 48075 1805 48109
rect 1805 48075 1839 48109
rect 1839 48075 1848 48109
rect 1796 48066 1848 48075
rect 134846 48109 134898 48118
rect 134846 48075 134855 48109
rect 134855 48075 134889 48109
rect 134889 48075 134898 48109
rect 134846 48066 134898 48075
rect 1796 47773 1848 47782
rect 1796 47739 1805 47773
rect 1805 47739 1839 47773
rect 1839 47739 1848 47773
rect 1796 47730 1848 47739
rect 134846 47773 134898 47782
rect 134846 47739 134855 47773
rect 134855 47739 134889 47773
rect 134889 47739 134898 47773
rect 134846 47730 134898 47739
rect 1796 47437 1848 47446
rect 1796 47403 1805 47437
rect 1805 47403 1839 47437
rect 1839 47403 1848 47437
rect 1796 47394 1848 47403
rect 134846 47437 134898 47446
rect 134846 47403 134855 47437
rect 134855 47403 134889 47437
rect 134889 47403 134898 47437
rect 134846 47394 134898 47403
rect 1796 47101 1848 47110
rect 1796 47067 1805 47101
rect 1805 47067 1839 47101
rect 1839 47067 1848 47101
rect 1796 47058 1848 47067
rect 134846 47101 134898 47110
rect 134846 47067 134855 47101
rect 134855 47067 134889 47101
rect 134889 47067 134898 47101
rect 134846 47058 134898 47067
rect 1796 46765 1848 46774
rect 1796 46731 1805 46765
rect 1805 46731 1839 46765
rect 1839 46731 1848 46765
rect 1796 46722 1848 46731
rect 134846 46765 134898 46774
rect 134846 46731 134855 46765
rect 134855 46731 134889 46765
rect 134889 46731 134898 46765
rect 134846 46722 134898 46731
rect 1796 46429 1848 46438
rect 1796 46395 1805 46429
rect 1805 46395 1839 46429
rect 1839 46395 1848 46429
rect 1796 46386 1848 46395
rect 134846 46429 134898 46438
rect 134846 46395 134855 46429
rect 134855 46395 134889 46429
rect 134889 46395 134898 46429
rect 134846 46386 134898 46395
rect 1796 46093 1848 46102
rect 1796 46059 1805 46093
rect 1805 46059 1839 46093
rect 1839 46059 1848 46093
rect 1796 46050 1848 46059
rect 134846 46093 134898 46102
rect 134846 46059 134855 46093
rect 134855 46059 134889 46093
rect 134889 46059 134898 46093
rect 134846 46050 134898 46059
rect 1796 45757 1848 45766
rect 1796 45723 1805 45757
rect 1805 45723 1839 45757
rect 1839 45723 1848 45757
rect 1796 45714 1848 45723
rect 134846 45757 134898 45766
rect 134846 45723 134855 45757
rect 134855 45723 134889 45757
rect 134889 45723 134898 45757
rect 134846 45714 134898 45723
rect 1796 45421 1848 45430
rect 1796 45387 1805 45421
rect 1805 45387 1839 45421
rect 1839 45387 1848 45421
rect 1796 45378 1848 45387
rect 134846 45421 134898 45430
rect 134846 45387 134855 45421
rect 134855 45387 134889 45421
rect 134889 45387 134898 45421
rect 134846 45378 134898 45387
rect 1796 45085 1848 45094
rect 1796 45051 1805 45085
rect 1805 45051 1839 45085
rect 1839 45051 1848 45085
rect 1796 45042 1848 45051
rect 134846 45085 134898 45094
rect 134846 45051 134855 45085
rect 134855 45051 134889 45085
rect 134889 45051 134898 45085
rect 134846 45042 134898 45051
rect 1796 44749 1848 44758
rect 1796 44715 1805 44749
rect 1805 44715 1839 44749
rect 1839 44715 1848 44749
rect 1796 44706 1848 44715
rect 134846 44749 134898 44758
rect 134846 44715 134855 44749
rect 134855 44715 134889 44749
rect 134889 44715 134898 44749
rect 134846 44706 134898 44715
rect 1796 44413 1848 44422
rect 1796 44379 1805 44413
rect 1805 44379 1839 44413
rect 1839 44379 1848 44413
rect 1796 44370 1848 44379
rect 134846 44413 134898 44422
rect 134846 44379 134855 44413
rect 134855 44379 134889 44413
rect 134889 44379 134898 44413
rect 134846 44370 134898 44379
rect 1796 44077 1848 44086
rect 1796 44043 1805 44077
rect 1805 44043 1839 44077
rect 1839 44043 1848 44077
rect 1796 44034 1848 44043
rect 134846 44077 134898 44086
rect 134846 44043 134855 44077
rect 134855 44043 134889 44077
rect 134889 44043 134898 44077
rect 134846 44034 134898 44043
rect 1796 43741 1848 43750
rect 1796 43707 1805 43741
rect 1805 43707 1839 43741
rect 1839 43707 1848 43741
rect 1796 43698 1848 43707
rect 134846 43741 134898 43750
rect 134846 43707 134855 43741
rect 134855 43707 134889 43741
rect 134889 43707 134898 43741
rect 134846 43698 134898 43707
rect 1796 43405 1848 43414
rect 1796 43371 1805 43405
rect 1805 43371 1839 43405
rect 1839 43371 1848 43405
rect 1796 43362 1848 43371
rect 134846 43405 134898 43414
rect 134846 43371 134855 43405
rect 134855 43371 134889 43405
rect 134889 43371 134898 43405
rect 134846 43362 134898 43371
rect 1796 43069 1848 43078
rect 1796 43035 1805 43069
rect 1805 43035 1839 43069
rect 1839 43035 1848 43069
rect 1796 43026 1848 43035
rect 134846 43069 134898 43078
rect 134846 43035 134855 43069
rect 134855 43035 134889 43069
rect 134889 43035 134898 43069
rect 134846 43026 134898 43035
rect 1796 42733 1848 42742
rect 1796 42699 1805 42733
rect 1805 42699 1839 42733
rect 1839 42699 1848 42733
rect 1796 42690 1848 42699
rect 134846 42733 134898 42742
rect 134846 42699 134855 42733
rect 134855 42699 134889 42733
rect 134889 42699 134898 42733
rect 134846 42690 134898 42699
rect 1796 42397 1848 42406
rect 1796 42363 1805 42397
rect 1805 42363 1839 42397
rect 1839 42363 1848 42397
rect 1796 42354 1848 42363
rect 134846 42397 134898 42406
rect 134846 42363 134855 42397
rect 134855 42363 134889 42397
rect 134889 42363 134898 42397
rect 134846 42354 134898 42363
rect 1796 42061 1848 42070
rect 1796 42027 1805 42061
rect 1805 42027 1839 42061
rect 1839 42027 1848 42061
rect 1796 42018 1848 42027
rect 134846 42061 134898 42070
rect 134846 42027 134855 42061
rect 134855 42027 134889 42061
rect 134889 42027 134898 42061
rect 134846 42018 134898 42027
rect 1796 41725 1848 41734
rect 1796 41691 1805 41725
rect 1805 41691 1839 41725
rect 1839 41691 1848 41725
rect 1796 41682 1848 41691
rect 134846 41725 134898 41734
rect 134846 41691 134855 41725
rect 134855 41691 134889 41725
rect 134889 41691 134898 41725
rect 134846 41682 134898 41691
rect 1796 41389 1848 41398
rect 1796 41355 1805 41389
rect 1805 41355 1839 41389
rect 1839 41355 1848 41389
rect 1796 41346 1848 41355
rect 134846 41389 134898 41398
rect 134846 41355 134855 41389
rect 134855 41355 134889 41389
rect 134889 41355 134898 41389
rect 134846 41346 134898 41355
rect 1796 41053 1848 41062
rect 1796 41019 1805 41053
rect 1805 41019 1839 41053
rect 1839 41019 1848 41053
rect 1796 41010 1848 41019
rect 134846 41053 134898 41062
rect 134846 41019 134855 41053
rect 134855 41019 134889 41053
rect 134889 41019 134898 41053
rect 134846 41010 134898 41019
rect 1796 40717 1848 40726
rect 1796 40683 1805 40717
rect 1805 40683 1839 40717
rect 1839 40683 1848 40717
rect 1796 40674 1848 40683
rect 134846 40717 134898 40726
rect 134846 40683 134855 40717
rect 134855 40683 134889 40717
rect 134889 40683 134898 40717
rect 134846 40674 134898 40683
rect 1796 40381 1848 40390
rect 1796 40347 1805 40381
rect 1805 40347 1839 40381
rect 1839 40347 1848 40381
rect 1796 40338 1848 40347
rect 134846 40381 134898 40390
rect 134846 40347 134855 40381
rect 134855 40347 134889 40381
rect 134889 40347 134898 40381
rect 134846 40338 134898 40347
rect 1796 40045 1848 40054
rect 1796 40011 1805 40045
rect 1805 40011 1839 40045
rect 1839 40011 1848 40045
rect 1796 40002 1848 40011
rect 134846 40045 134898 40054
rect 134846 40011 134855 40045
rect 134855 40011 134889 40045
rect 134889 40011 134898 40045
rect 134846 40002 134898 40011
rect 1796 39709 1848 39718
rect 1796 39675 1805 39709
rect 1805 39675 1839 39709
rect 1839 39675 1848 39709
rect 1796 39666 1848 39675
rect 134846 39709 134898 39718
rect 134846 39675 134855 39709
rect 134855 39675 134889 39709
rect 134889 39675 134898 39709
rect 134846 39666 134898 39675
rect 1796 39373 1848 39382
rect 1796 39339 1805 39373
rect 1805 39339 1839 39373
rect 1839 39339 1848 39373
rect 1796 39330 1848 39339
rect 134846 39373 134898 39382
rect 134846 39339 134855 39373
rect 134855 39339 134889 39373
rect 134889 39339 134898 39373
rect 134846 39330 134898 39339
rect 1796 39037 1848 39046
rect 1796 39003 1805 39037
rect 1805 39003 1839 39037
rect 1839 39003 1848 39037
rect 1796 38994 1848 39003
rect 134846 39037 134898 39046
rect 134846 39003 134855 39037
rect 134855 39003 134889 39037
rect 134889 39003 134898 39037
rect 134846 38994 134898 39003
rect 1796 38701 1848 38710
rect 1796 38667 1805 38701
rect 1805 38667 1839 38701
rect 1839 38667 1848 38701
rect 1796 38658 1848 38667
rect 134846 38701 134898 38710
rect 134846 38667 134855 38701
rect 134855 38667 134889 38701
rect 134889 38667 134898 38701
rect 134846 38658 134898 38667
rect 1796 38365 1848 38374
rect 1796 38331 1805 38365
rect 1805 38331 1839 38365
rect 1839 38331 1848 38365
rect 1796 38322 1848 38331
rect 134846 38365 134898 38374
rect 134846 38331 134855 38365
rect 134855 38331 134889 38365
rect 134889 38331 134898 38365
rect 134846 38322 134898 38331
rect 1796 38029 1848 38038
rect 1796 37995 1805 38029
rect 1805 37995 1839 38029
rect 1839 37995 1848 38029
rect 1796 37986 1848 37995
rect 134846 38029 134898 38038
rect 134846 37995 134855 38029
rect 134855 37995 134889 38029
rect 134889 37995 134898 38029
rect 134846 37986 134898 37995
rect 1796 37693 1848 37702
rect 1796 37659 1805 37693
rect 1805 37659 1839 37693
rect 1839 37659 1848 37693
rect 1796 37650 1848 37659
rect 134846 37693 134898 37702
rect 134846 37659 134855 37693
rect 134855 37659 134889 37693
rect 134889 37659 134898 37693
rect 134846 37650 134898 37659
rect 1796 37357 1848 37366
rect 1796 37323 1805 37357
rect 1805 37323 1839 37357
rect 1839 37323 1848 37357
rect 1796 37314 1848 37323
rect 134846 37357 134898 37366
rect 134846 37323 134855 37357
rect 134855 37323 134889 37357
rect 134889 37323 134898 37357
rect 134846 37314 134898 37323
rect 1796 37021 1848 37030
rect 1796 36987 1805 37021
rect 1805 36987 1839 37021
rect 1839 36987 1848 37021
rect 1796 36978 1848 36987
rect 134846 37021 134898 37030
rect 134846 36987 134855 37021
rect 134855 36987 134889 37021
rect 134889 36987 134898 37021
rect 134846 36978 134898 36987
rect 15349 36839 15401 36891
rect 1796 36685 1848 36694
rect 1796 36651 1805 36685
rect 1805 36651 1839 36685
rect 1839 36651 1848 36685
rect 1796 36642 1848 36651
rect 1796 36349 1848 36358
rect 1796 36315 1805 36349
rect 1805 36315 1839 36349
rect 1839 36315 1848 36349
rect 1796 36306 1848 36315
rect 1796 36013 1848 36022
rect 1796 35979 1805 36013
rect 1805 35979 1839 36013
rect 1839 35979 1848 36013
rect 1796 35970 1848 35979
rect 1796 35677 1848 35686
rect 1796 35643 1805 35677
rect 1805 35643 1839 35677
rect 1839 35643 1848 35677
rect 1796 35634 1848 35643
rect 15269 35569 15321 35621
rect 1796 35341 1848 35350
rect 1796 35307 1805 35341
rect 1805 35307 1839 35341
rect 1839 35307 1848 35341
rect 1796 35298 1848 35307
rect 1796 35005 1848 35014
rect 1796 34971 1805 35005
rect 1805 34971 1839 35005
rect 1839 34971 1848 35005
rect 1796 34962 1848 34971
rect 1796 34669 1848 34678
rect 1796 34635 1805 34669
rect 1805 34635 1839 34669
rect 1839 34635 1848 34669
rect 1796 34626 1848 34635
rect 1796 34333 1848 34342
rect 1796 34299 1805 34333
rect 1805 34299 1839 34333
rect 1839 34299 1848 34333
rect 1796 34290 1848 34299
rect 15189 34011 15241 34063
rect 1796 33997 1848 34006
rect 1796 33963 1805 33997
rect 1805 33963 1839 33997
rect 1839 33963 1848 33997
rect 1796 33954 1848 33963
rect 1796 33661 1848 33670
rect 1796 33627 1805 33661
rect 1805 33627 1839 33661
rect 1839 33627 1848 33661
rect 1796 33618 1848 33627
rect 1796 33325 1848 33334
rect 1796 33291 1805 33325
rect 1805 33291 1839 33325
rect 1839 33291 1848 33325
rect 1796 33282 1848 33291
rect 1796 32989 1848 32998
rect 1796 32955 1805 32989
rect 1805 32955 1839 32989
rect 1839 32955 1848 32989
rect 1796 32946 1848 32955
rect 15109 32741 15161 32793
rect 1796 32653 1848 32662
rect 1796 32619 1805 32653
rect 1805 32619 1839 32653
rect 1839 32619 1848 32653
rect 1796 32610 1848 32619
rect 1796 32317 1848 32326
rect 1796 32283 1805 32317
rect 1805 32283 1839 32317
rect 1839 32283 1848 32317
rect 1796 32274 1848 32283
rect 1796 31981 1848 31990
rect 1796 31947 1805 31981
rect 1805 31947 1839 31981
rect 1839 31947 1848 31981
rect 1796 31938 1848 31947
rect 1796 31645 1848 31654
rect 1796 31611 1805 31645
rect 1805 31611 1839 31645
rect 1839 31611 1848 31645
rect 1796 31602 1848 31611
rect 1796 31309 1848 31318
rect 1796 31275 1805 31309
rect 1805 31275 1839 31309
rect 1839 31275 1848 31309
rect 1796 31266 1848 31275
rect 15029 31183 15081 31235
rect 1796 30973 1848 30982
rect 1796 30939 1805 30973
rect 1805 30939 1839 30973
rect 1839 30939 1848 30973
rect 1796 30930 1848 30939
rect 1796 30637 1848 30646
rect 1796 30603 1805 30637
rect 1805 30603 1839 30637
rect 1839 30603 1848 30637
rect 1796 30594 1848 30603
rect 1796 30301 1848 30310
rect 1796 30267 1805 30301
rect 1805 30267 1839 30301
rect 1839 30267 1848 30301
rect 1796 30258 1848 30267
rect 1796 29965 1848 29974
rect 1796 29931 1805 29965
rect 1805 29931 1839 29965
rect 1839 29931 1848 29965
rect 1796 29922 1848 29931
rect 14949 29913 15001 29965
rect 1796 29629 1848 29638
rect 1796 29595 1805 29629
rect 1805 29595 1839 29629
rect 1839 29595 1848 29629
rect 1796 29586 1848 29595
rect 1796 29293 1848 29302
rect 1796 29259 1805 29293
rect 1805 29259 1839 29293
rect 1839 29259 1848 29293
rect 1796 29250 1848 29259
rect 1796 28957 1848 28966
rect 1796 28923 1805 28957
rect 1805 28923 1839 28957
rect 1839 28923 1848 28957
rect 1796 28914 1848 28923
rect 1796 28621 1848 28630
rect 1796 28587 1805 28621
rect 1805 28587 1839 28621
rect 1839 28587 1848 28621
rect 1796 28578 1848 28587
rect 14869 28355 14921 28407
rect 1796 28285 1848 28294
rect 1796 28251 1805 28285
rect 1805 28251 1839 28285
rect 1839 28251 1848 28285
rect 1796 28242 1848 28251
rect 1796 27949 1848 27958
rect 1796 27915 1805 27949
rect 1805 27915 1839 27949
rect 1839 27915 1848 27949
rect 1796 27906 1848 27915
rect 1796 27613 1848 27622
rect 1796 27579 1805 27613
rect 1805 27579 1839 27613
rect 1839 27579 1848 27613
rect 1796 27570 1848 27579
rect 1796 27277 1848 27286
rect 1796 27243 1805 27277
rect 1805 27243 1839 27277
rect 1839 27243 1848 27277
rect 1796 27234 1848 27243
rect 1796 26941 1848 26950
rect 1796 26907 1805 26941
rect 1805 26907 1839 26941
rect 1839 26907 1848 26941
rect 1796 26898 1848 26907
rect 1796 26605 1848 26614
rect 1796 26571 1805 26605
rect 1805 26571 1839 26605
rect 1839 26571 1848 26605
rect 1796 26562 1848 26571
rect 1796 26269 1848 26278
rect 1796 26235 1805 26269
rect 1805 26235 1839 26269
rect 1839 26235 1848 26269
rect 1796 26226 1848 26235
rect 1796 25933 1848 25942
rect 1796 25899 1805 25933
rect 1805 25899 1839 25933
rect 1839 25899 1848 25933
rect 1796 25890 1848 25899
rect 1796 25597 1848 25606
rect 1796 25563 1805 25597
rect 1805 25563 1839 25597
rect 1839 25563 1848 25597
rect 1796 25554 1848 25563
rect 1796 25261 1848 25270
rect 1796 25227 1805 25261
rect 1805 25227 1839 25261
rect 1839 25227 1848 25261
rect 1796 25218 1848 25227
rect 1796 24925 1848 24934
rect 1796 24891 1805 24925
rect 1805 24891 1839 24925
rect 1839 24891 1848 24925
rect 1796 24882 1848 24891
rect 1796 24589 1848 24598
rect 1796 24555 1805 24589
rect 1805 24555 1839 24589
rect 1839 24555 1848 24589
rect 1796 24546 1848 24555
rect 1796 24253 1848 24262
rect 1796 24219 1805 24253
rect 1805 24219 1839 24253
rect 1839 24219 1848 24253
rect 1796 24210 1848 24219
rect 1796 23917 1848 23926
rect 1796 23883 1805 23917
rect 1805 23883 1839 23917
rect 1839 23883 1848 23917
rect 1796 23874 1848 23883
rect 134846 36685 134898 36694
rect 134846 36651 134855 36685
rect 134855 36651 134889 36685
rect 134889 36651 134898 36685
rect 134846 36642 134898 36651
rect 134846 36349 134898 36358
rect 134846 36315 134855 36349
rect 134855 36315 134889 36349
rect 134889 36315 134898 36349
rect 134846 36306 134898 36315
rect 134846 36013 134898 36022
rect 134846 35979 134855 36013
rect 134855 35979 134889 36013
rect 134889 35979 134898 36013
rect 134846 35970 134898 35979
rect 134846 35677 134898 35686
rect 134846 35643 134855 35677
rect 134855 35643 134889 35677
rect 134889 35643 134898 35677
rect 134846 35634 134898 35643
rect 134846 35341 134898 35350
rect 134846 35307 134855 35341
rect 134855 35307 134889 35341
rect 134889 35307 134898 35341
rect 134846 35298 134898 35307
rect 134846 35005 134898 35014
rect 134846 34971 134855 35005
rect 134855 34971 134889 35005
rect 134889 34971 134898 35005
rect 134846 34962 134898 34971
rect 134846 34669 134898 34678
rect 134846 34635 134855 34669
rect 134855 34635 134889 34669
rect 134889 34635 134898 34669
rect 134846 34626 134898 34635
rect 134846 34333 134898 34342
rect 134846 34299 134855 34333
rect 134855 34299 134889 34333
rect 134889 34299 134898 34333
rect 134846 34290 134898 34299
rect 134846 33997 134898 34006
rect 134846 33963 134855 33997
rect 134855 33963 134889 33997
rect 134889 33963 134898 33997
rect 134846 33954 134898 33963
rect 134846 33661 134898 33670
rect 134846 33627 134855 33661
rect 134855 33627 134889 33661
rect 134889 33627 134898 33661
rect 134846 33618 134898 33627
rect 134846 33325 134898 33334
rect 134846 33291 134855 33325
rect 134855 33291 134889 33325
rect 134889 33291 134898 33325
rect 134846 33282 134898 33291
rect 134846 32989 134898 32998
rect 134846 32955 134855 32989
rect 134855 32955 134889 32989
rect 134889 32955 134898 32989
rect 134846 32946 134898 32955
rect 134846 32653 134898 32662
rect 134846 32619 134855 32653
rect 134855 32619 134889 32653
rect 134889 32619 134898 32653
rect 134846 32610 134898 32619
rect 134846 32317 134898 32326
rect 134846 32283 134855 32317
rect 134855 32283 134889 32317
rect 134889 32283 134898 32317
rect 134846 32274 134898 32283
rect 134846 31981 134898 31990
rect 134846 31947 134855 31981
rect 134855 31947 134889 31981
rect 134889 31947 134898 31981
rect 134846 31938 134898 31947
rect 134846 31645 134898 31654
rect 134846 31611 134855 31645
rect 134855 31611 134889 31645
rect 134889 31611 134898 31645
rect 134846 31602 134898 31611
rect 134846 31309 134898 31318
rect 134846 31275 134855 31309
rect 134855 31275 134889 31309
rect 134889 31275 134898 31309
rect 134846 31266 134898 31275
rect 134846 30973 134898 30982
rect 134846 30939 134855 30973
rect 134855 30939 134889 30973
rect 134889 30939 134898 30973
rect 134846 30930 134898 30939
rect 134846 30637 134898 30646
rect 134846 30603 134855 30637
rect 134855 30603 134889 30637
rect 134889 30603 134898 30637
rect 134846 30594 134898 30603
rect 134846 30301 134898 30310
rect 134846 30267 134855 30301
rect 134855 30267 134889 30301
rect 134889 30267 134898 30301
rect 134846 30258 134898 30267
rect 134846 29965 134898 29974
rect 134846 29931 134855 29965
rect 134855 29931 134889 29965
rect 134889 29931 134898 29965
rect 134846 29922 134898 29931
rect 134846 29629 134898 29638
rect 134846 29595 134855 29629
rect 134855 29595 134889 29629
rect 134889 29595 134898 29629
rect 134846 29586 134898 29595
rect 134846 29293 134898 29302
rect 134846 29259 134855 29293
rect 134855 29259 134889 29293
rect 134889 29259 134898 29293
rect 134846 29250 134898 29259
rect 134846 28957 134898 28966
rect 134846 28923 134855 28957
rect 134855 28923 134889 28957
rect 134889 28923 134898 28957
rect 134846 28914 134898 28923
rect 134846 28621 134898 28630
rect 134846 28587 134855 28621
rect 134855 28587 134889 28621
rect 134889 28587 134898 28621
rect 134846 28578 134898 28587
rect 134846 28285 134898 28294
rect 134846 28251 134855 28285
rect 134855 28251 134889 28285
rect 134889 28251 134898 28285
rect 134846 28242 134898 28251
rect 134846 27949 134898 27958
rect 134846 27915 134855 27949
rect 134855 27915 134889 27949
rect 134889 27915 134898 27949
rect 134846 27906 134898 27915
rect 134846 27613 134898 27622
rect 134846 27579 134855 27613
rect 134855 27579 134889 27613
rect 134889 27579 134898 27613
rect 134846 27570 134898 27579
rect 134846 27277 134898 27286
rect 134846 27243 134855 27277
rect 134855 27243 134889 27277
rect 134889 27243 134898 27277
rect 134846 27234 134898 27243
rect 134846 26941 134898 26950
rect 134846 26907 134855 26941
rect 134855 26907 134889 26941
rect 134889 26907 134898 26941
rect 134846 26898 134898 26907
rect 134846 26605 134898 26614
rect 134846 26571 134855 26605
rect 134855 26571 134889 26605
rect 134889 26571 134898 26605
rect 134846 26562 134898 26571
rect 134846 26269 134898 26278
rect 134846 26235 134855 26269
rect 134855 26235 134889 26269
rect 134889 26235 134898 26269
rect 134846 26226 134898 26235
rect 134846 25933 134898 25942
rect 134846 25899 134855 25933
rect 134855 25899 134889 25933
rect 134889 25899 134898 25933
rect 134846 25890 134898 25899
rect 134846 25597 134898 25606
rect 134846 25563 134855 25597
rect 134855 25563 134889 25597
rect 134889 25563 134898 25597
rect 134846 25554 134898 25563
rect 134846 25261 134898 25270
rect 134846 25227 134855 25261
rect 134855 25227 134889 25261
rect 134889 25227 134898 25261
rect 134846 25218 134898 25227
rect 134846 24925 134898 24934
rect 134846 24891 134855 24925
rect 134855 24891 134889 24925
rect 134889 24891 134898 24925
rect 134846 24882 134898 24891
rect 134846 24589 134898 24598
rect 134846 24555 134855 24589
rect 134855 24555 134889 24589
rect 134889 24555 134898 24589
rect 134846 24546 134898 24555
rect 134846 24253 134898 24262
rect 134846 24219 134855 24253
rect 134855 24219 134889 24253
rect 134889 24219 134898 24253
rect 134846 24210 134898 24219
rect 134846 23917 134898 23926
rect 134846 23883 134855 23917
rect 134855 23883 134889 23917
rect 134889 23883 134898 23917
rect 134846 23874 134898 23883
rect 1796 23581 1848 23590
rect 1796 23547 1805 23581
rect 1805 23547 1839 23581
rect 1839 23547 1848 23581
rect 1796 23538 1848 23547
rect 1796 23245 1848 23254
rect 1796 23211 1805 23245
rect 1805 23211 1839 23245
rect 1839 23211 1848 23245
rect 1796 23202 1848 23211
rect 1796 22909 1848 22918
rect 1796 22875 1805 22909
rect 1805 22875 1839 22909
rect 1839 22875 1848 22909
rect 1796 22866 1848 22875
rect 1796 22573 1848 22582
rect 1796 22539 1805 22573
rect 1805 22539 1839 22573
rect 1839 22539 1848 22573
rect 1796 22530 1848 22539
rect 1796 22237 1848 22246
rect 1796 22203 1805 22237
rect 1805 22203 1839 22237
rect 1839 22203 1848 22237
rect 1796 22194 1848 22203
rect 1796 21901 1848 21910
rect 1796 21867 1805 21901
rect 1805 21867 1839 21901
rect 1839 21867 1848 21901
rect 1796 21858 1848 21867
rect 1796 21565 1848 21574
rect 1796 21531 1805 21565
rect 1805 21531 1839 21565
rect 1839 21531 1848 21565
rect 1796 21522 1848 21531
rect 1796 21229 1848 21238
rect 1796 21195 1805 21229
rect 1805 21195 1839 21229
rect 1839 21195 1848 21229
rect 1796 21186 1848 21195
rect 1796 20893 1848 20902
rect 1796 20859 1805 20893
rect 1805 20859 1839 20893
rect 1839 20859 1848 20893
rect 1796 20850 1848 20859
rect 1796 20557 1848 20566
rect 1796 20523 1805 20557
rect 1805 20523 1839 20557
rect 1839 20523 1848 20557
rect 1796 20514 1848 20523
rect 1796 20221 1848 20230
rect 1796 20187 1805 20221
rect 1805 20187 1839 20221
rect 1839 20187 1848 20221
rect 1796 20178 1848 20187
rect 1796 19885 1848 19894
rect 1796 19851 1805 19885
rect 1805 19851 1839 19885
rect 1839 19851 1848 19885
rect 1796 19842 1848 19851
rect 1796 19549 1848 19558
rect 1796 19515 1805 19549
rect 1805 19515 1839 19549
rect 1839 19515 1848 19549
rect 1796 19506 1848 19515
rect 1796 19213 1848 19222
rect 1796 19179 1805 19213
rect 1805 19179 1839 19213
rect 1839 19179 1848 19213
rect 1796 19170 1848 19179
rect 1796 18877 1848 18886
rect 1796 18843 1805 18877
rect 1805 18843 1839 18877
rect 1839 18843 1848 18877
rect 1796 18834 1848 18843
rect 1796 18541 1848 18550
rect 1796 18507 1805 18541
rect 1805 18507 1839 18541
rect 1839 18507 1848 18541
rect 1796 18498 1848 18507
rect 1796 18205 1848 18214
rect 1796 18171 1805 18205
rect 1805 18171 1839 18205
rect 1839 18171 1848 18205
rect 1796 18162 1848 18171
rect 1796 17869 1848 17878
rect 1796 17835 1805 17869
rect 1805 17835 1839 17869
rect 1839 17835 1848 17869
rect 1796 17826 1848 17835
rect 1796 17533 1848 17542
rect 1796 17499 1805 17533
rect 1805 17499 1839 17533
rect 1839 17499 1848 17533
rect 1796 17490 1848 17499
rect 1796 17197 1848 17206
rect 1796 17163 1805 17197
rect 1805 17163 1839 17197
rect 1839 17163 1848 17197
rect 1796 17154 1848 17163
rect 1796 16861 1848 16870
rect 1796 16827 1805 16861
rect 1805 16827 1839 16861
rect 1839 16827 1848 16861
rect 1796 16818 1848 16827
rect 1796 16525 1848 16534
rect 1796 16491 1805 16525
rect 1805 16491 1839 16525
rect 1839 16491 1848 16525
rect 1796 16482 1848 16491
rect 1796 16189 1848 16198
rect 1796 16155 1805 16189
rect 1805 16155 1839 16189
rect 1839 16155 1848 16189
rect 1796 16146 1848 16155
rect 1796 15853 1848 15862
rect 1796 15819 1805 15853
rect 1805 15819 1839 15853
rect 1839 15819 1848 15853
rect 1796 15810 1848 15819
rect 1796 15517 1848 15526
rect 1796 15483 1805 15517
rect 1805 15483 1839 15517
rect 1839 15483 1848 15517
rect 1796 15474 1848 15483
rect 1796 15181 1848 15190
rect 1796 15147 1805 15181
rect 1805 15147 1839 15181
rect 1839 15147 1848 15181
rect 1796 15138 1848 15147
rect 1796 14845 1848 14854
rect 1796 14811 1805 14845
rect 1805 14811 1839 14845
rect 1839 14811 1848 14845
rect 1796 14802 1848 14811
rect 1796 14509 1848 14518
rect 1796 14475 1805 14509
rect 1805 14475 1839 14509
rect 1839 14475 1848 14509
rect 1796 14466 1848 14475
rect 1796 14173 1848 14182
rect 1796 14139 1805 14173
rect 1805 14139 1839 14173
rect 1839 14139 1848 14173
rect 1796 14130 1848 14139
rect 1796 13837 1848 13846
rect 1796 13803 1805 13837
rect 1805 13803 1839 13837
rect 1839 13803 1848 13837
rect 1796 13794 1848 13803
rect 1796 13501 1848 13510
rect 1796 13467 1805 13501
rect 1805 13467 1839 13501
rect 1839 13467 1848 13501
rect 1796 13458 1848 13467
rect 28620 13207 28672 13259
rect 31116 13207 31168 13259
rect 33612 13207 33664 13259
rect 36108 13207 36160 13259
rect 38604 13207 38656 13259
rect 41100 13207 41152 13259
rect 43596 13207 43648 13259
rect 46092 13207 46144 13259
rect 48588 13207 48640 13259
rect 51084 13207 51136 13259
rect 53580 13207 53632 13259
rect 56076 13207 56128 13259
rect 58572 13207 58624 13259
rect 61068 13207 61120 13259
rect 63564 13207 63616 13259
rect 66060 13207 66112 13259
rect 68556 13207 68608 13259
rect 71052 13207 71104 13259
rect 73548 13207 73600 13259
rect 76044 13207 76096 13259
rect 78540 13207 78592 13259
rect 81036 13207 81088 13259
rect 83532 13207 83584 13259
rect 86028 13207 86080 13259
rect 88524 13207 88576 13259
rect 91020 13207 91072 13259
rect 93516 13207 93568 13259
rect 96012 13207 96064 13259
rect 98508 13207 98560 13259
rect 101004 13207 101056 13259
rect 103500 13207 103552 13259
rect 105996 13207 106048 13259
rect 1796 13165 1848 13174
rect 1796 13131 1805 13165
rect 1805 13131 1839 13165
rect 1839 13131 1848 13165
rect 1796 13122 1848 13131
rect 1796 12829 1848 12838
rect 1796 12795 1805 12829
rect 1805 12795 1839 12829
rect 1839 12795 1848 12829
rect 1796 12786 1848 12795
rect 1796 12493 1848 12502
rect 1796 12459 1805 12493
rect 1805 12459 1839 12493
rect 1839 12459 1848 12493
rect 1796 12450 1848 12459
rect 1796 12157 1848 12166
rect 1796 12123 1805 12157
rect 1805 12123 1839 12157
rect 1839 12123 1848 12157
rect 1796 12114 1848 12123
rect 1796 11821 1848 11830
rect 1796 11787 1805 11821
rect 1805 11787 1839 11821
rect 1839 11787 1848 11821
rect 1796 11778 1848 11787
rect 1796 11485 1848 11494
rect 1796 11451 1805 11485
rect 1805 11451 1839 11485
rect 1839 11451 1848 11485
rect 1796 11442 1848 11451
rect 1796 11149 1848 11158
rect 1796 11115 1805 11149
rect 1805 11115 1839 11149
rect 1839 11115 1848 11149
rect 1796 11106 1848 11115
rect 1796 10813 1848 10822
rect 1796 10779 1805 10813
rect 1805 10779 1839 10813
rect 1839 10779 1848 10813
rect 1796 10770 1848 10779
rect 134846 23581 134898 23590
rect 134846 23547 134855 23581
rect 134855 23547 134889 23581
rect 134889 23547 134898 23581
rect 134846 23538 134898 23547
rect 134846 23245 134898 23254
rect 134846 23211 134855 23245
rect 134855 23211 134889 23245
rect 134889 23211 134898 23245
rect 134846 23202 134898 23211
rect 134846 22909 134898 22918
rect 134846 22875 134855 22909
rect 134855 22875 134889 22909
rect 134889 22875 134898 22909
rect 134846 22866 134898 22875
rect 134846 22573 134898 22582
rect 134846 22539 134855 22573
rect 134855 22539 134889 22573
rect 134889 22539 134898 22573
rect 134846 22530 134898 22539
rect 134846 22237 134898 22246
rect 134846 22203 134855 22237
rect 134855 22203 134889 22237
rect 134889 22203 134898 22237
rect 134846 22194 134898 22203
rect 134846 21901 134898 21910
rect 134846 21867 134855 21901
rect 134855 21867 134889 21901
rect 134889 21867 134898 21901
rect 134846 21858 134898 21867
rect 134846 21565 134898 21574
rect 134846 21531 134855 21565
rect 134855 21531 134889 21565
rect 134889 21531 134898 21565
rect 134846 21522 134898 21531
rect 134846 21229 134898 21238
rect 134846 21195 134855 21229
rect 134855 21195 134889 21229
rect 134889 21195 134898 21229
rect 134846 21186 134898 21195
rect 134846 20893 134898 20902
rect 134846 20859 134855 20893
rect 134855 20859 134889 20893
rect 134889 20859 134898 20893
rect 134846 20850 134898 20859
rect 134846 20557 134898 20566
rect 134846 20523 134855 20557
rect 134855 20523 134889 20557
rect 134889 20523 134898 20557
rect 134846 20514 134898 20523
rect 134846 20221 134898 20230
rect 134846 20187 134855 20221
rect 134855 20187 134889 20221
rect 134889 20187 134898 20221
rect 134846 20178 134898 20187
rect 134846 19885 134898 19894
rect 134846 19851 134855 19885
rect 134855 19851 134889 19885
rect 134889 19851 134898 19885
rect 134846 19842 134898 19851
rect 134846 19549 134898 19558
rect 134846 19515 134855 19549
rect 134855 19515 134889 19549
rect 134889 19515 134898 19549
rect 134846 19506 134898 19515
rect 121989 19185 122041 19237
rect 134846 19213 134898 19222
rect 134846 19179 134855 19213
rect 134855 19179 134889 19213
rect 134889 19179 134898 19213
rect 134846 19170 134898 19179
rect 134846 18877 134898 18886
rect 134846 18843 134855 18877
rect 134855 18843 134889 18877
rect 134889 18843 134898 18877
rect 134846 18834 134898 18843
rect 134846 18541 134898 18550
rect 134846 18507 134855 18541
rect 134855 18507 134889 18541
rect 134889 18507 134898 18541
rect 134846 18498 134898 18507
rect 134846 18205 134898 18214
rect 134846 18171 134855 18205
rect 134855 18171 134889 18205
rect 134889 18171 134898 18205
rect 134846 18162 134898 18171
rect 134846 17869 134898 17878
rect 134846 17835 134855 17869
rect 134855 17835 134889 17869
rect 134889 17835 134898 17869
rect 134846 17826 134898 17835
rect 121909 17627 121961 17679
rect 134846 17533 134898 17542
rect 134846 17499 134855 17533
rect 134855 17499 134889 17533
rect 134889 17499 134898 17533
rect 134846 17490 134898 17499
rect 134846 17197 134898 17206
rect 134846 17163 134855 17197
rect 134855 17163 134889 17197
rect 134889 17163 134898 17197
rect 134846 17154 134898 17163
rect 134846 16861 134898 16870
rect 134846 16827 134855 16861
rect 134855 16827 134889 16861
rect 134889 16827 134898 16861
rect 134846 16818 134898 16827
rect 134846 16525 134898 16534
rect 134846 16491 134855 16525
rect 134855 16491 134889 16525
rect 134889 16491 134898 16525
rect 134846 16482 134898 16491
rect 121829 16357 121881 16409
rect 134846 16189 134898 16198
rect 134846 16155 134855 16189
rect 134855 16155 134889 16189
rect 134889 16155 134898 16189
rect 134846 16146 134898 16155
rect 134846 15853 134898 15862
rect 134846 15819 134855 15853
rect 134855 15819 134889 15853
rect 134889 15819 134898 15853
rect 134846 15810 134898 15819
rect 134846 15517 134898 15526
rect 134846 15483 134855 15517
rect 134855 15483 134889 15517
rect 134889 15483 134898 15517
rect 134846 15474 134898 15483
rect 134846 15181 134898 15190
rect 134846 15147 134855 15181
rect 134855 15147 134889 15181
rect 134889 15147 134898 15181
rect 134846 15138 134898 15147
rect 121749 14799 121801 14851
rect 134846 14845 134898 14854
rect 134846 14811 134855 14845
rect 134855 14811 134889 14845
rect 134889 14811 134898 14845
rect 134846 14802 134898 14811
rect 134846 14509 134898 14518
rect 134846 14475 134855 14509
rect 134855 14475 134889 14509
rect 134889 14475 134898 14509
rect 134846 14466 134898 14475
rect 134846 14173 134898 14182
rect 134846 14139 134855 14173
rect 134855 14139 134889 14173
rect 134889 14139 134898 14173
rect 134846 14130 134898 14139
rect 134846 13837 134898 13846
rect 134846 13803 134855 13837
rect 134855 13803 134889 13837
rect 134889 13803 134898 13837
rect 134846 13794 134898 13803
rect 121669 13529 121721 13581
rect 134846 13501 134898 13510
rect 134846 13467 134855 13501
rect 134855 13467 134889 13501
rect 134889 13467 134898 13501
rect 134846 13458 134898 13467
rect 134846 13165 134898 13174
rect 134846 13131 134855 13165
rect 134855 13131 134889 13165
rect 134889 13131 134898 13165
rect 134846 13122 134898 13131
rect 134846 12829 134898 12838
rect 134846 12795 134855 12829
rect 134855 12795 134889 12829
rect 134889 12795 134898 12829
rect 134846 12786 134898 12795
rect 134846 12493 134898 12502
rect 134846 12459 134855 12493
rect 134855 12459 134889 12493
rect 134889 12459 134898 12493
rect 134846 12450 134898 12459
rect 134846 12157 134898 12166
rect 134846 12123 134855 12157
rect 134855 12123 134889 12157
rect 134889 12123 134898 12157
rect 134846 12114 134898 12123
rect 121589 11971 121641 12023
rect 134846 11821 134898 11830
rect 134846 11787 134855 11821
rect 134855 11787 134889 11821
rect 134889 11787 134898 11821
rect 134846 11778 134898 11787
rect 134846 11485 134898 11494
rect 134846 11451 134855 11485
rect 134855 11451 134889 11485
rect 134889 11451 134898 11485
rect 134846 11442 134898 11451
rect 134846 11149 134898 11158
rect 134846 11115 134855 11149
rect 134855 11115 134889 11149
rect 134889 11115 134898 11149
rect 134846 11106 134898 11115
rect 134846 10813 134898 10822
rect 134846 10779 134855 10813
rect 134855 10779 134889 10813
rect 134889 10779 134898 10813
rect 134846 10770 134898 10779
rect 121509 10701 121561 10753
rect 1796 10477 1848 10486
rect 1796 10443 1805 10477
rect 1805 10443 1839 10477
rect 1839 10443 1848 10477
rect 1796 10434 1848 10443
rect 134846 10477 134898 10486
rect 134846 10443 134855 10477
rect 134855 10443 134889 10477
rect 134889 10443 134898 10477
rect 134846 10434 134898 10443
rect 1796 10141 1848 10150
rect 1796 10107 1805 10141
rect 1805 10107 1839 10141
rect 1839 10107 1848 10141
rect 1796 10098 1848 10107
rect 134846 10141 134898 10150
rect 134846 10107 134855 10141
rect 134855 10107 134889 10141
rect 134889 10107 134898 10141
rect 134846 10098 134898 10107
rect 1796 9805 1848 9814
rect 1796 9771 1805 9805
rect 1805 9771 1839 9805
rect 1839 9771 1848 9805
rect 1796 9762 1848 9771
rect 134846 9805 134898 9814
rect 134846 9771 134855 9805
rect 134855 9771 134889 9805
rect 134889 9771 134898 9805
rect 134846 9762 134898 9771
rect 1796 9469 1848 9478
rect 1796 9435 1805 9469
rect 1805 9435 1839 9469
rect 1839 9435 1848 9469
rect 1796 9426 1848 9435
rect 134846 9469 134898 9478
rect 134846 9435 134855 9469
rect 134855 9435 134889 9469
rect 134889 9435 134898 9469
rect 134846 9426 134898 9435
rect 1796 9133 1848 9142
rect 1796 9099 1805 9133
rect 1805 9099 1839 9133
rect 1839 9099 1848 9133
rect 1796 9090 1848 9099
rect 134846 9133 134898 9142
rect 134846 9099 134855 9133
rect 134855 9099 134889 9133
rect 134889 9099 134898 9133
rect 134846 9090 134898 9099
rect 1796 8797 1848 8806
rect 1796 8763 1805 8797
rect 1805 8763 1839 8797
rect 1839 8763 1848 8797
rect 1796 8754 1848 8763
rect 134846 8797 134898 8806
rect 134846 8763 134855 8797
rect 134855 8763 134889 8797
rect 134889 8763 134898 8797
rect 134846 8754 134898 8763
rect 1796 8461 1848 8470
rect 1796 8427 1805 8461
rect 1805 8427 1839 8461
rect 1839 8427 1848 8461
rect 1796 8418 1848 8427
rect 134846 8461 134898 8470
rect 134846 8427 134855 8461
rect 134855 8427 134889 8461
rect 134889 8427 134898 8461
rect 134846 8418 134898 8427
rect 1796 8125 1848 8134
rect 1796 8091 1805 8125
rect 1805 8091 1839 8125
rect 1839 8091 1848 8125
rect 1796 8082 1848 8091
rect 134846 8125 134898 8134
rect 134846 8091 134855 8125
rect 134855 8091 134889 8125
rect 134889 8091 134898 8125
rect 134846 8082 134898 8091
rect 1796 7789 1848 7798
rect 1796 7755 1805 7789
rect 1805 7755 1839 7789
rect 1839 7755 1848 7789
rect 1796 7746 1848 7755
rect 134846 7789 134898 7798
rect 134846 7755 134855 7789
rect 134855 7755 134889 7789
rect 134889 7755 134898 7789
rect 134846 7746 134898 7755
rect 1796 7453 1848 7462
rect 1796 7419 1805 7453
rect 1805 7419 1839 7453
rect 1839 7419 1848 7453
rect 1796 7410 1848 7419
rect 134846 7453 134898 7462
rect 134846 7419 134855 7453
rect 134855 7419 134889 7453
rect 134889 7419 134898 7453
rect 134846 7410 134898 7419
rect 1796 7117 1848 7126
rect 1796 7083 1805 7117
rect 1805 7083 1839 7117
rect 1839 7083 1848 7117
rect 1796 7074 1848 7083
rect 134846 7117 134898 7126
rect 134846 7083 134855 7117
rect 134855 7083 134889 7117
rect 134889 7083 134898 7117
rect 134846 7074 134898 7083
rect 1796 6781 1848 6790
rect 1796 6747 1805 6781
rect 1805 6747 1839 6781
rect 1839 6747 1848 6781
rect 1796 6738 1848 6747
rect 134846 6781 134898 6790
rect 134846 6747 134855 6781
rect 134855 6747 134889 6781
rect 134889 6747 134898 6781
rect 134846 6738 134898 6747
rect 1796 6445 1848 6454
rect 1796 6411 1805 6445
rect 1805 6411 1839 6445
rect 1839 6411 1848 6445
rect 1796 6402 1848 6411
rect 134846 6445 134898 6454
rect 134846 6411 134855 6445
rect 134855 6411 134889 6445
rect 134889 6411 134898 6445
rect 134846 6402 134898 6411
rect 1796 6109 1848 6118
rect 1796 6075 1805 6109
rect 1805 6075 1839 6109
rect 1839 6075 1848 6109
rect 1796 6066 1848 6075
rect 134846 6109 134898 6118
rect 134846 6075 134855 6109
rect 134855 6075 134889 6109
rect 134889 6075 134898 6109
rect 134846 6066 134898 6075
rect 1796 5773 1848 5782
rect 1796 5739 1805 5773
rect 1805 5739 1839 5773
rect 1839 5739 1848 5773
rect 1796 5730 1848 5739
rect 134846 5773 134898 5782
rect 134846 5739 134855 5773
rect 134855 5739 134889 5773
rect 134889 5739 134898 5773
rect 134846 5730 134898 5739
rect 1796 5437 1848 5446
rect 1796 5403 1805 5437
rect 1805 5403 1839 5437
rect 1839 5403 1848 5437
rect 1796 5394 1848 5403
rect 134846 5437 134898 5446
rect 134846 5403 134855 5437
rect 134855 5403 134889 5437
rect 134889 5403 134898 5437
rect 134846 5394 134898 5403
rect 1796 5101 1848 5110
rect 1796 5067 1805 5101
rect 1805 5067 1839 5101
rect 1839 5067 1848 5101
rect 1796 5058 1848 5067
rect 134846 5101 134898 5110
rect 134846 5067 134855 5101
rect 134855 5067 134889 5101
rect 134889 5067 134898 5101
rect 134846 5058 134898 5067
rect 1796 4765 1848 4774
rect 1796 4731 1805 4765
rect 1805 4731 1839 4765
rect 1839 4731 1848 4765
rect 1796 4722 1848 4731
rect 134846 4765 134898 4774
rect 134846 4731 134855 4765
rect 134855 4731 134889 4765
rect 134889 4731 134898 4765
rect 134846 4722 134898 4731
rect 1796 4429 1848 4438
rect 1796 4395 1805 4429
rect 1805 4395 1839 4429
rect 1839 4395 1848 4429
rect 1796 4386 1848 4395
rect 134846 4429 134898 4438
rect 134846 4395 134855 4429
rect 134855 4395 134889 4429
rect 134889 4395 134898 4429
rect 134846 4386 134898 4395
rect 1796 4093 1848 4102
rect 1796 4059 1805 4093
rect 1805 4059 1839 4093
rect 1839 4059 1848 4093
rect 1796 4050 1848 4059
rect 134846 4093 134898 4102
rect 134846 4059 134855 4093
rect 134855 4059 134889 4093
rect 134889 4059 134898 4093
rect 134846 4050 134898 4059
rect 1796 3757 1848 3766
rect 1796 3723 1805 3757
rect 1805 3723 1839 3757
rect 1839 3723 1848 3757
rect 1796 3714 1848 3723
rect 134846 3757 134898 3766
rect 134846 3723 134855 3757
rect 134855 3723 134889 3757
rect 134889 3723 134898 3757
rect 134846 3714 134898 3723
rect 1796 3421 1848 3430
rect 1796 3387 1805 3421
rect 1805 3387 1839 3421
rect 1839 3387 1848 3421
rect 1796 3378 1848 3387
rect 134846 3421 134898 3430
rect 134846 3387 134855 3421
rect 134855 3387 134889 3421
rect 134889 3387 134898 3421
rect 134846 3378 134898 3387
rect 1796 3085 1848 3094
rect 1796 3051 1805 3085
rect 1805 3051 1839 3085
rect 1839 3051 1848 3085
rect 1796 3042 1848 3051
rect 134846 3085 134898 3094
rect 134846 3051 134855 3085
rect 134855 3051 134889 3085
rect 134889 3051 134898 3085
rect 134846 3042 134898 3051
rect 1796 2749 1848 2758
rect 1796 2715 1805 2749
rect 1805 2715 1839 2749
rect 1839 2715 1848 2749
rect 1796 2706 1848 2715
rect 134846 2749 134898 2758
rect 134846 2715 134855 2749
rect 134855 2715 134889 2749
rect 134889 2715 134898 2749
rect 134846 2706 134898 2715
rect 1796 2413 1848 2422
rect 1796 2379 1805 2413
rect 1805 2379 1839 2413
rect 1839 2379 1848 2413
rect 1796 2370 1848 2379
rect 134846 2413 134898 2422
rect 134846 2379 134855 2413
rect 134855 2379 134889 2413
rect 134889 2379 134898 2413
rect 134846 2370 134898 2379
rect 1796 2077 1848 2086
rect 1796 2043 1805 2077
rect 1805 2043 1839 2077
rect 1839 2043 1848 2077
rect 1796 2034 1848 2043
rect 134846 2077 134898 2086
rect 134846 2043 134855 2077
rect 134855 2043 134889 2077
rect 134889 2043 134898 2077
rect 134846 2034 134898 2043
rect 2132 1741 2184 1750
rect 3812 1741 3864 1750
rect 5492 1741 5544 1750
rect 7172 1741 7224 1750
rect 8852 1741 8904 1750
rect 10532 1741 10584 1750
rect 12212 1741 12264 1750
rect 13892 1741 13944 1750
rect 15572 1741 15624 1750
rect 17252 1741 17304 1750
rect 18932 1741 18984 1750
rect 20612 1741 20664 1750
rect 22292 1741 22344 1750
rect 23972 1741 24024 1750
rect 25652 1741 25704 1750
rect 27332 1741 27384 1750
rect 29012 1741 29064 1750
rect 30692 1741 30744 1750
rect 32372 1741 32424 1750
rect 34052 1741 34104 1750
rect 35732 1741 35784 1750
rect 37412 1741 37464 1750
rect 39092 1741 39144 1750
rect 40772 1741 40824 1750
rect 42452 1741 42504 1750
rect 44132 1741 44184 1750
rect 45812 1741 45864 1750
rect 47492 1741 47544 1750
rect 49172 1741 49224 1750
rect 50852 1741 50904 1750
rect 52532 1741 52584 1750
rect 54212 1741 54264 1750
rect 55892 1741 55944 1750
rect 57572 1741 57624 1750
rect 59252 1741 59304 1750
rect 60932 1741 60984 1750
rect 62612 1741 62664 1750
rect 64292 1741 64344 1750
rect 65972 1741 66024 1750
rect 67652 1741 67704 1750
rect 69332 1741 69384 1750
rect 71012 1741 71064 1750
rect 72692 1741 72744 1750
rect 74372 1741 74424 1750
rect 76052 1741 76104 1750
rect 77732 1741 77784 1750
rect 79412 1741 79464 1750
rect 81092 1741 81144 1750
rect 82772 1741 82824 1750
rect 84452 1741 84504 1750
rect 86132 1741 86184 1750
rect 87812 1741 87864 1750
rect 89492 1741 89544 1750
rect 91172 1741 91224 1750
rect 92852 1741 92904 1750
rect 94532 1741 94584 1750
rect 96212 1741 96264 1750
rect 97892 1741 97944 1750
rect 99572 1741 99624 1750
rect 101252 1741 101304 1750
rect 102932 1741 102984 1750
rect 104612 1741 104664 1750
rect 106292 1741 106344 1750
rect 107972 1741 108024 1750
rect 109652 1741 109704 1750
rect 111332 1741 111384 1750
rect 113012 1741 113064 1750
rect 114692 1741 114744 1750
rect 116372 1741 116424 1750
rect 118052 1741 118104 1750
rect 119732 1741 119784 1750
rect 121412 1741 121464 1750
rect 123092 1741 123144 1750
rect 124772 1741 124824 1750
rect 126452 1741 126504 1750
rect 128132 1741 128184 1750
rect 129812 1741 129864 1750
rect 131492 1741 131544 1750
rect 133172 1741 133224 1750
rect 2132 1707 2141 1741
rect 2141 1707 2175 1741
rect 2175 1707 2184 1741
rect 3812 1707 3821 1741
rect 3821 1707 3855 1741
rect 3855 1707 3864 1741
rect 5492 1707 5501 1741
rect 5501 1707 5535 1741
rect 5535 1707 5544 1741
rect 7172 1707 7181 1741
rect 7181 1707 7215 1741
rect 7215 1707 7224 1741
rect 8852 1707 8861 1741
rect 8861 1707 8895 1741
rect 8895 1707 8904 1741
rect 10532 1707 10541 1741
rect 10541 1707 10575 1741
rect 10575 1707 10584 1741
rect 12212 1707 12221 1741
rect 12221 1707 12255 1741
rect 12255 1707 12264 1741
rect 13892 1707 13901 1741
rect 13901 1707 13935 1741
rect 13935 1707 13944 1741
rect 15572 1707 15581 1741
rect 15581 1707 15615 1741
rect 15615 1707 15624 1741
rect 17252 1707 17261 1741
rect 17261 1707 17295 1741
rect 17295 1707 17304 1741
rect 18932 1707 18941 1741
rect 18941 1707 18975 1741
rect 18975 1707 18984 1741
rect 20612 1707 20621 1741
rect 20621 1707 20655 1741
rect 20655 1707 20664 1741
rect 22292 1707 22301 1741
rect 22301 1707 22335 1741
rect 22335 1707 22344 1741
rect 23972 1707 23981 1741
rect 23981 1707 24015 1741
rect 24015 1707 24024 1741
rect 25652 1707 25661 1741
rect 25661 1707 25695 1741
rect 25695 1707 25704 1741
rect 27332 1707 27341 1741
rect 27341 1707 27375 1741
rect 27375 1707 27384 1741
rect 29012 1707 29021 1741
rect 29021 1707 29055 1741
rect 29055 1707 29064 1741
rect 30692 1707 30701 1741
rect 30701 1707 30735 1741
rect 30735 1707 30744 1741
rect 32372 1707 32381 1741
rect 32381 1707 32415 1741
rect 32415 1707 32424 1741
rect 34052 1707 34061 1741
rect 34061 1707 34095 1741
rect 34095 1707 34104 1741
rect 35732 1707 35741 1741
rect 35741 1707 35775 1741
rect 35775 1707 35784 1741
rect 37412 1707 37421 1741
rect 37421 1707 37455 1741
rect 37455 1707 37464 1741
rect 39092 1707 39101 1741
rect 39101 1707 39135 1741
rect 39135 1707 39144 1741
rect 40772 1707 40781 1741
rect 40781 1707 40815 1741
rect 40815 1707 40824 1741
rect 42452 1707 42461 1741
rect 42461 1707 42495 1741
rect 42495 1707 42504 1741
rect 44132 1707 44141 1741
rect 44141 1707 44175 1741
rect 44175 1707 44184 1741
rect 45812 1707 45821 1741
rect 45821 1707 45855 1741
rect 45855 1707 45864 1741
rect 47492 1707 47501 1741
rect 47501 1707 47535 1741
rect 47535 1707 47544 1741
rect 49172 1707 49181 1741
rect 49181 1707 49215 1741
rect 49215 1707 49224 1741
rect 50852 1707 50861 1741
rect 50861 1707 50895 1741
rect 50895 1707 50904 1741
rect 52532 1707 52541 1741
rect 52541 1707 52575 1741
rect 52575 1707 52584 1741
rect 54212 1707 54221 1741
rect 54221 1707 54255 1741
rect 54255 1707 54264 1741
rect 55892 1707 55901 1741
rect 55901 1707 55935 1741
rect 55935 1707 55944 1741
rect 57572 1707 57581 1741
rect 57581 1707 57615 1741
rect 57615 1707 57624 1741
rect 59252 1707 59261 1741
rect 59261 1707 59295 1741
rect 59295 1707 59304 1741
rect 60932 1707 60941 1741
rect 60941 1707 60975 1741
rect 60975 1707 60984 1741
rect 62612 1707 62621 1741
rect 62621 1707 62655 1741
rect 62655 1707 62664 1741
rect 64292 1707 64301 1741
rect 64301 1707 64335 1741
rect 64335 1707 64344 1741
rect 65972 1707 65981 1741
rect 65981 1707 66015 1741
rect 66015 1707 66024 1741
rect 67652 1707 67661 1741
rect 67661 1707 67695 1741
rect 67695 1707 67704 1741
rect 69332 1707 69341 1741
rect 69341 1707 69375 1741
rect 69375 1707 69384 1741
rect 71012 1707 71021 1741
rect 71021 1707 71055 1741
rect 71055 1707 71064 1741
rect 72692 1707 72701 1741
rect 72701 1707 72735 1741
rect 72735 1707 72744 1741
rect 74372 1707 74381 1741
rect 74381 1707 74415 1741
rect 74415 1707 74424 1741
rect 76052 1707 76061 1741
rect 76061 1707 76095 1741
rect 76095 1707 76104 1741
rect 77732 1707 77741 1741
rect 77741 1707 77775 1741
rect 77775 1707 77784 1741
rect 79412 1707 79421 1741
rect 79421 1707 79455 1741
rect 79455 1707 79464 1741
rect 81092 1707 81101 1741
rect 81101 1707 81135 1741
rect 81135 1707 81144 1741
rect 82772 1707 82781 1741
rect 82781 1707 82815 1741
rect 82815 1707 82824 1741
rect 84452 1707 84461 1741
rect 84461 1707 84495 1741
rect 84495 1707 84504 1741
rect 86132 1707 86141 1741
rect 86141 1707 86175 1741
rect 86175 1707 86184 1741
rect 87812 1707 87821 1741
rect 87821 1707 87855 1741
rect 87855 1707 87864 1741
rect 89492 1707 89501 1741
rect 89501 1707 89535 1741
rect 89535 1707 89544 1741
rect 91172 1707 91181 1741
rect 91181 1707 91215 1741
rect 91215 1707 91224 1741
rect 92852 1707 92861 1741
rect 92861 1707 92895 1741
rect 92895 1707 92904 1741
rect 94532 1707 94541 1741
rect 94541 1707 94575 1741
rect 94575 1707 94584 1741
rect 96212 1707 96221 1741
rect 96221 1707 96255 1741
rect 96255 1707 96264 1741
rect 97892 1707 97901 1741
rect 97901 1707 97935 1741
rect 97935 1707 97944 1741
rect 99572 1707 99581 1741
rect 99581 1707 99615 1741
rect 99615 1707 99624 1741
rect 101252 1707 101261 1741
rect 101261 1707 101295 1741
rect 101295 1707 101304 1741
rect 102932 1707 102941 1741
rect 102941 1707 102975 1741
rect 102975 1707 102984 1741
rect 104612 1707 104621 1741
rect 104621 1707 104655 1741
rect 104655 1707 104664 1741
rect 106292 1707 106301 1741
rect 106301 1707 106335 1741
rect 106335 1707 106344 1741
rect 107972 1707 107981 1741
rect 107981 1707 108015 1741
rect 108015 1707 108024 1741
rect 109652 1707 109661 1741
rect 109661 1707 109695 1741
rect 109695 1707 109704 1741
rect 111332 1707 111341 1741
rect 111341 1707 111375 1741
rect 111375 1707 111384 1741
rect 113012 1707 113021 1741
rect 113021 1707 113055 1741
rect 113055 1707 113064 1741
rect 114692 1707 114701 1741
rect 114701 1707 114735 1741
rect 114735 1707 114744 1741
rect 116372 1707 116381 1741
rect 116381 1707 116415 1741
rect 116415 1707 116424 1741
rect 118052 1707 118061 1741
rect 118061 1707 118095 1741
rect 118095 1707 118104 1741
rect 119732 1707 119741 1741
rect 119741 1707 119775 1741
rect 119775 1707 119784 1741
rect 121412 1707 121421 1741
rect 121421 1707 121455 1741
rect 121455 1707 121464 1741
rect 123092 1707 123101 1741
rect 123101 1707 123135 1741
rect 123135 1707 123144 1741
rect 124772 1707 124781 1741
rect 124781 1707 124815 1741
rect 124815 1707 124824 1741
rect 126452 1707 126461 1741
rect 126461 1707 126495 1741
rect 126495 1707 126504 1741
rect 128132 1707 128141 1741
rect 128141 1707 128175 1741
rect 128175 1707 128184 1741
rect 129812 1707 129821 1741
rect 129821 1707 129855 1741
rect 129855 1707 129864 1741
rect 131492 1707 131501 1741
rect 131501 1707 131535 1741
rect 131535 1707 131544 1741
rect 133172 1707 133181 1741
rect 133181 1707 133215 1741
rect 133215 1707 133224 1741
rect 2132 1698 2184 1707
rect 3812 1698 3864 1707
rect 5492 1698 5544 1707
rect 7172 1698 7224 1707
rect 8852 1698 8904 1707
rect 10532 1698 10584 1707
rect 12212 1698 12264 1707
rect 13892 1698 13944 1707
rect 15572 1698 15624 1707
rect 17252 1698 17304 1707
rect 18932 1698 18984 1707
rect 20612 1698 20664 1707
rect 22292 1698 22344 1707
rect 23972 1698 24024 1707
rect 25652 1698 25704 1707
rect 27332 1698 27384 1707
rect 29012 1698 29064 1707
rect 30692 1698 30744 1707
rect 32372 1698 32424 1707
rect 34052 1698 34104 1707
rect 35732 1698 35784 1707
rect 37412 1698 37464 1707
rect 39092 1698 39144 1707
rect 40772 1698 40824 1707
rect 42452 1698 42504 1707
rect 44132 1698 44184 1707
rect 45812 1698 45864 1707
rect 47492 1698 47544 1707
rect 49172 1698 49224 1707
rect 50852 1698 50904 1707
rect 52532 1698 52584 1707
rect 54212 1698 54264 1707
rect 55892 1698 55944 1707
rect 57572 1698 57624 1707
rect 59252 1698 59304 1707
rect 60932 1698 60984 1707
rect 62612 1698 62664 1707
rect 64292 1698 64344 1707
rect 65972 1698 66024 1707
rect 67652 1698 67704 1707
rect 69332 1698 69384 1707
rect 71012 1698 71064 1707
rect 72692 1698 72744 1707
rect 74372 1698 74424 1707
rect 76052 1698 76104 1707
rect 77732 1698 77784 1707
rect 79412 1698 79464 1707
rect 81092 1698 81144 1707
rect 82772 1698 82824 1707
rect 84452 1698 84504 1707
rect 86132 1698 86184 1707
rect 87812 1698 87864 1707
rect 89492 1698 89544 1707
rect 91172 1698 91224 1707
rect 92852 1698 92904 1707
rect 94532 1698 94584 1707
rect 96212 1698 96264 1707
rect 97892 1698 97944 1707
rect 99572 1698 99624 1707
rect 101252 1698 101304 1707
rect 102932 1698 102984 1707
rect 104612 1698 104664 1707
rect 106292 1698 106344 1707
rect 107972 1698 108024 1707
rect 109652 1698 109704 1707
rect 111332 1698 111384 1707
rect 113012 1698 113064 1707
rect 114692 1698 114744 1707
rect 116372 1698 116424 1707
rect 118052 1698 118104 1707
rect 119732 1698 119784 1707
rect 121412 1698 121464 1707
rect 123092 1698 123144 1707
rect 124772 1698 124824 1707
rect 126452 1698 126504 1707
rect 128132 1698 128184 1707
rect 129812 1698 129864 1707
rect 131492 1698 131544 1707
rect 133172 1698 133224 1707
<< metal2 >>
rect 1710 81048 1934 81585
rect 2130 81501 2186 81510
rect 2130 81436 2186 81445
rect 3810 81501 3866 81510
rect 3810 81436 3866 81445
rect 5490 81501 5546 81510
rect 5490 81436 5546 81445
rect 7170 81501 7226 81510
rect 7170 81436 7226 81445
rect 8850 81501 8906 81510
rect 8850 81436 8906 81445
rect 10530 81501 10586 81510
rect 10530 81436 10586 81445
rect 12210 81501 12266 81510
rect 12210 81436 12266 81445
rect 13890 81501 13946 81510
rect 13890 81436 13946 81445
rect 15570 81501 15626 81510
rect 15570 81436 15626 81445
rect 17250 81501 17306 81510
rect 17250 81436 17306 81445
rect 18930 81501 18986 81510
rect 18930 81436 18986 81445
rect 20610 81501 20666 81510
rect 20610 81436 20666 81445
rect 22290 81501 22346 81510
rect 22290 81436 22346 81445
rect 23970 81501 24026 81510
rect 23970 81436 24026 81445
rect 25650 81501 25706 81510
rect 25650 81436 25706 81445
rect 27330 81501 27386 81510
rect 27330 81436 27386 81445
rect 29010 81501 29066 81510
rect 29010 81436 29066 81445
rect 30690 81501 30746 81510
rect 30690 81436 30746 81445
rect 32370 81501 32426 81510
rect 32370 81436 32426 81445
rect 34050 81501 34106 81510
rect 34050 81436 34106 81445
rect 35730 81501 35786 81510
rect 35730 81436 35786 81445
rect 37410 81501 37466 81510
rect 37410 81436 37466 81445
rect 39090 81501 39146 81510
rect 39090 81436 39146 81445
rect 40770 81501 40826 81510
rect 40770 81436 40826 81445
rect 42450 81501 42506 81510
rect 42450 81436 42506 81445
rect 44130 81501 44186 81510
rect 44130 81436 44186 81445
rect 45810 81501 45866 81510
rect 45810 81436 45866 81445
rect 47490 81501 47546 81510
rect 47490 81436 47546 81445
rect 49170 81501 49226 81510
rect 49170 81436 49226 81445
rect 50850 81501 50906 81510
rect 50850 81436 50906 81445
rect 52530 81501 52586 81510
rect 52530 81436 52586 81445
rect 54210 81501 54266 81510
rect 54210 81436 54266 81445
rect 55890 81501 55946 81510
rect 55890 81436 55946 81445
rect 57570 81501 57626 81510
rect 57570 81436 57626 81445
rect 59250 81501 59306 81510
rect 59250 81436 59306 81445
rect 60930 81501 60986 81510
rect 60930 81436 60986 81445
rect 62610 81501 62666 81510
rect 62610 81436 62666 81445
rect 64290 81501 64346 81510
rect 64290 81436 64346 81445
rect 65970 81501 66026 81510
rect 65970 81436 66026 81445
rect 67650 81501 67706 81510
rect 67650 81436 67706 81445
rect 69330 81501 69386 81510
rect 69330 81436 69386 81445
rect 71010 81501 71066 81510
rect 71010 81436 71066 81445
rect 72690 81501 72746 81510
rect 72690 81436 72746 81445
rect 74370 81501 74426 81510
rect 74370 81436 74426 81445
rect 76050 81501 76106 81510
rect 76050 81436 76106 81445
rect 77730 81501 77786 81510
rect 77730 81436 77786 81445
rect 79410 81501 79466 81510
rect 79410 81436 79466 81445
rect 81090 81501 81146 81510
rect 81090 81436 81146 81445
rect 82770 81501 82826 81510
rect 82770 81436 82826 81445
rect 84450 81501 84506 81510
rect 84450 81436 84506 81445
rect 86130 81501 86186 81510
rect 86130 81436 86186 81445
rect 87810 81501 87866 81510
rect 87810 81436 87866 81445
rect 89490 81501 89546 81510
rect 89490 81436 89546 81445
rect 91170 81501 91226 81510
rect 91170 81436 91226 81445
rect 92850 81501 92906 81510
rect 92850 81436 92906 81445
rect 94530 81501 94586 81510
rect 94530 81436 94586 81445
rect 96210 81501 96266 81510
rect 96210 81436 96266 81445
rect 97890 81501 97946 81510
rect 97890 81436 97946 81445
rect 99570 81501 99626 81510
rect 99570 81436 99626 81445
rect 101250 81501 101306 81510
rect 101250 81436 101306 81445
rect 102930 81501 102986 81510
rect 102930 81436 102986 81445
rect 104610 81501 104666 81510
rect 104610 81436 104666 81445
rect 106290 81501 106346 81510
rect 106290 81436 106346 81445
rect 107970 81501 108026 81510
rect 107970 81436 108026 81445
rect 109650 81501 109706 81510
rect 109650 81436 109706 81445
rect 111330 81501 111386 81510
rect 111330 81436 111386 81445
rect 113010 81501 113066 81510
rect 113010 81436 113066 81445
rect 114690 81501 114746 81510
rect 114690 81436 114746 81445
rect 116370 81501 116426 81510
rect 116370 81436 116426 81445
rect 118050 81501 118106 81510
rect 118050 81436 118106 81445
rect 119730 81501 119786 81510
rect 119730 81436 119786 81445
rect 121410 81501 121466 81510
rect 121410 81436 121466 81445
rect 123090 81501 123146 81510
rect 123090 81436 123146 81445
rect 124770 81501 124826 81510
rect 124770 81436 124826 81445
rect 126450 81501 126506 81510
rect 126450 81436 126506 81445
rect 128130 81501 128186 81510
rect 128130 81436 128186 81445
rect 129810 81501 129866 81510
rect 129810 81436 129866 81445
rect 131490 81501 131546 81510
rect 131490 81436 131546 81445
rect 133170 81501 133226 81510
rect 133170 81436 133226 81445
rect 1710 80992 1794 81048
rect 1850 80992 1934 81048
rect 1710 80710 1934 80992
rect 1710 80658 1796 80710
rect 1848 80658 1934 80710
rect 1710 80374 1934 80658
rect 134760 81048 134984 81585
rect 134760 80992 134844 81048
rect 134900 80992 134984 81048
rect 134760 80710 134984 80992
rect 134760 80658 134846 80710
rect 134898 80658 134984 80710
rect 122188 80521 122244 80530
rect 122188 80456 122244 80465
rect 1710 80322 1796 80374
rect 1848 80322 1934 80374
rect 1710 80038 1934 80322
rect 118598 80265 118654 80274
rect 118598 80200 118654 80209
rect 119766 80265 119822 80274
rect 119766 80200 119822 80209
rect 1710 79986 1796 80038
rect 1848 79986 1934 80038
rect 1710 79702 1934 79986
rect 1710 79650 1796 79702
rect 1848 79650 1934 79702
rect 1710 79368 1934 79650
rect 1710 79312 1794 79368
rect 1850 79312 1934 79368
rect 1710 79030 1934 79312
rect 1710 78978 1796 79030
rect 1848 78978 1934 79030
rect 1710 78694 1934 78978
rect 1710 78642 1796 78694
rect 1848 78642 1934 78694
rect 1710 78358 1934 78642
rect 1710 78306 1796 78358
rect 1848 78306 1934 78358
rect 1710 78022 1934 78306
rect 1710 77970 1796 78022
rect 1848 77970 1934 78022
rect 1710 77688 1934 77970
rect 1710 77632 1794 77688
rect 1850 77632 1934 77688
rect 1710 77350 1934 77632
rect 1710 77298 1796 77350
rect 1848 77298 1934 77350
rect 1710 77014 1934 77298
rect 122202 79111 122230 80456
rect 134760 80374 134984 80658
rect 134760 80322 134846 80374
rect 134898 80322 134984 80374
rect 134760 80038 134984 80322
rect 134760 79986 134846 80038
rect 134898 79986 134984 80038
rect 134760 79702 134984 79986
rect 134760 79650 134846 79702
rect 134898 79650 134984 79702
rect 134760 79368 134984 79650
rect 134760 79312 134844 79368
rect 134900 79312 134984 79368
rect 133884 79268 133940 79277
rect 133884 79203 133940 79212
rect 130747 79163 130803 79172
rect 122202 79083 122300 79111
rect 130747 79098 130803 79107
rect 1710 76962 1796 77014
rect 1848 76962 1934 77014
rect 28618 77047 28674 77056
rect 28618 76982 28674 76991
rect 31114 77047 31170 77056
rect 31114 76982 31170 76991
rect 33610 77047 33666 77056
rect 33610 76982 33666 76991
rect 36106 77047 36162 77056
rect 36106 76982 36162 76991
rect 38602 77047 38658 77056
rect 38602 76982 38658 76991
rect 41098 77047 41154 77056
rect 41098 76982 41154 76991
rect 43594 77047 43650 77056
rect 43594 76982 43650 76991
rect 46090 77047 46146 77056
rect 46090 76982 46146 76991
rect 48586 77047 48642 77056
rect 48586 76982 48642 76991
rect 51082 77047 51138 77056
rect 51082 76982 51138 76991
rect 53578 77047 53634 77056
rect 53578 76982 53634 76991
rect 56074 77047 56130 77056
rect 56074 76982 56130 76991
rect 58570 77047 58626 77056
rect 58570 76982 58626 76991
rect 61066 77047 61122 77056
rect 61066 76982 61122 76991
rect 63562 77047 63618 77056
rect 63562 76982 63618 76991
rect 66058 77047 66114 77056
rect 66058 76982 66114 76991
rect 68554 77047 68610 77056
rect 68554 76982 68610 76991
rect 71050 77047 71106 77056
rect 71050 76982 71106 76991
rect 73546 77047 73602 77056
rect 73546 76982 73602 76991
rect 76042 77047 76098 77056
rect 76042 76982 76098 76991
rect 78538 77047 78594 77056
rect 78538 76982 78594 76991
rect 81034 77047 81090 77056
rect 81034 76982 81090 76991
rect 83530 77047 83586 77056
rect 83530 76982 83586 76991
rect 86026 77047 86082 77056
rect 86026 76982 86082 76991
rect 88522 77047 88578 77056
rect 88522 76982 88578 76991
rect 91018 77047 91074 77056
rect 91018 76982 91074 76991
rect 93514 77047 93570 77056
rect 93514 76982 93570 76991
rect 96010 77047 96066 77056
rect 96010 76982 96066 76991
rect 98506 77047 98562 77056
rect 98506 76982 98562 76991
rect 101002 77047 101058 77056
rect 101002 76982 101058 76991
rect 103498 77047 103554 77056
rect 103498 76982 103554 76991
rect 105994 77047 106050 77056
rect 105994 76982 106050 76991
rect 1710 76678 1934 76962
rect 1710 76626 1796 76678
rect 1848 76626 1934 76678
rect 1710 76342 1934 76626
rect 1710 76290 1796 76342
rect 1848 76290 1934 76342
rect 1710 76008 1934 76290
rect 1710 75952 1794 76008
rect 1850 75952 1934 76008
rect 1710 75670 1934 75952
rect 1710 75618 1796 75670
rect 1848 75618 1934 75670
rect 1710 75334 1934 75618
rect 1710 75282 1796 75334
rect 1848 75282 1934 75334
rect 1710 74998 1934 75282
rect 1710 74946 1796 74998
rect 1848 74946 1934 74998
rect 1710 74662 1934 74946
rect 110061 74883 110117 74915
rect 110061 74818 110117 74827
rect 1710 74610 1796 74662
rect 1848 74610 1934 74662
rect 1710 74328 1934 74610
rect 1710 74272 1794 74328
rect 1850 74272 1934 74328
rect 1710 73990 1934 74272
rect 1710 73938 1796 73990
rect 1848 73938 1934 73990
rect 1710 73654 1934 73938
rect 1710 73602 1796 73654
rect 1848 73602 1934 73654
rect 1710 73318 1934 73602
rect 1710 73266 1796 73318
rect 1848 73266 1934 73318
rect 1710 72982 1934 73266
rect 1710 72930 1796 72982
rect 1848 72930 1934 72982
rect 1710 72648 1934 72930
rect 1710 72592 1794 72648
rect 1850 72592 1934 72648
rect 1710 72310 1934 72592
rect 1710 72258 1796 72310
rect 1848 72258 1934 72310
rect 1710 71974 1934 72258
rect 1710 71922 1796 71974
rect 1848 71922 1934 71974
rect 1710 71638 1934 71922
rect 1710 71586 1796 71638
rect 1848 71586 1934 71638
rect 1710 71302 1934 71586
rect 1710 71250 1796 71302
rect 1848 71250 1934 71302
rect 1710 70968 1934 71250
rect 110075 71182 110103 74818
rect 110185 73469 110241 73478
rect 110185 73404 110241 73413
rect 110199 71182 110227 73404
rect 114046 72055 114102 72064
rect 114046 71990 114102 71999
rect 1710 70912 1794 70968
rect 1850 70912 1934 70968
rect 1710 70630 1934 70912
rect 114060 70705 114088 71990
rect 1710 70578 1796 70630
rect 1848 70578 1934 70630
rect 1710 70294 1934 70578
rect 1710 70242 1796 70294
rect 1848 70242 1934 70294
rect 1710 69958 1934 70242
rect 1710 69906 1796 69958
rect 1848 69906 1934 69958
rect 1710 69622 1934 69906
rect 1710 69570 1796 69622
rect 1848 69570 1934 69622
rect 1710 69288 1934 69570
rect 1710 69232 1794 69288
rect 1850 69232 1934 69288
rect 1710 68950 1934 69232
rect 1710 68898 1796 68950
rect 1848 68898 1934 68950
rect 1710 68614 1934 68898
rect 1710 68562 1796 68614
rect 1848 68562 1934 68614
rect 1710 68278 1934 68562
rect 1710 68226 1796 68278
rect 1848 68226 1934 68278
rect 1710 67942 1934 68226
rect 1710 67890 1796 67942
rect 1848 67890 1934 67942
rect 1710 67608 1934 67890
rect 1710 67552 1794 67608
rect 1850 67552 1934 67608
rect 1710 67270 1934 67552
rect 1710 67218 1796 67270
rect 1848 67218 1934 67270
rect 1710 66934 1934 67218
rect 1710 66882 1796 66934
rect 1848 66882 1934 66934
rect 1710 66598 1934 66882
rect 1710 66546 1796 66598
rect 1848 66546 1934 66598
rect 1710 66262 1934 66546
rect 1710 66210 1796 66262
rect 1848 66210 1934 66262
rect 1710 65928 1934 66210
rect 1710 65872 1794 65928
rect 1850 65872 1934 65928
rect 1710 65590 1934 65872
rect 1710 65538 1796 65590
rect 1848 65538 1934 65590
rect 1710 65254 1934 65538
rect 1710 65202 1796 65254
rect 1848 65202 1934 65254
rect 1710 64918 1934 65202
rect 1710 64866 1796 64918
rect 1848 64866 1934 64918
rect 1710 64582 1934 64866
rect 1710 64530 1796 64582
rect 1848 64530 1934 64582
rect 1710 64248 1934 64530
rect 1710 64192 1794 64248
rect 1850 64192 1934 64248
rect 1710 63910 1934 64192
rect 1710 63858 1796 63910
rect 1848 63858 1934 63910
rect 1710 63574 1934 63858
rect 1710 63522 1796 63574
rect 1848 63522 1934 63574
rect 1710 63238 1934 63522
rect 1710 63186 1796 63238
rect 1848 63186 1934 63238
rect 1710 62902 1934 63186
rect 1710 62850 1796 62902
rect 1848 62850 1934 62902
rect 1710 62568 1934 62850
rect 1710 62512 1794 62568
rect 1850 62512 1934 62568
rect 1710 62230 1934 62512
rect 1710 62178 1796 62230
rect 1848 62178 1934 62230
rect 1710 61894 1934 62178
rect 1710 61842 1796 61894
rect 1848 61842 1934 61894
rect 1710 61558 1934 61842
rect 1710 61506 1796 61558
rect 1848 61506 1934 61558
rect 1710 61222 1934 61506
rect 1710 61170 1796 61222
rect 1848 61170 1934 61222
rect 1710 60888 1934 61170
rect 1710 60832 1794 60888
rect 1850 60832 1934 60888
rect 1710 60550 1934 60832
rect 1710 60498 1796 60550
rect 1848 60498 1934 60550
rect 1710 60214 1934 60498
rect 1710 60162 1796 60214
rect 1848 60162 1934 60214
rect 1710 59878 1934 60162
rect 1710 59826 1796 59878
rect 1848 59826 1934 59878
rect 1710 59542 1934 59826
rect 1710 59490 1796 59542
rect 1848 59490 1934 59542
rect 1710 59208 1934 59490
rect 1710 59152 1794 59208
rect 1850 59152 1934 59208
rect 1710 58870 1934 59152
rect 1710 58818 1796 58870
rect 1848 58818 1934 58870
rect 1710 58534 1934 58818
rect 1710 58482 1796 58534
rect 1848 58482 1934 58534
rect 1710 58198 1934 58482
rect 1710 58146 1796 58198
rect 1848 58146 1934 58198
rect 1710 57862 1934 58146
rect 1710 57810 1796 57862
rect 1848 57810 1934 57862
rect 1710 57528 1934 57810
rect 1710 57472 1794 57528
rect 1850 57472 1934 57528
rect 1710 57190 1934 57472
rect 1710 57138 1796 57190
rect 1848 57138 1934 57190
rect 1710 56854 1934 57138
rect 1710 56802 1796 56854
rect 1848 56802 1934 56854
rect 1710 56518 1934 56802
rect 1710 56466 1796 56518
rect 1848 56466 1934 56518
rect 1710 56182 1934 56466
rect 1710 56130 1796 56182
rect 1848 56130 1934 56182
rect 1710 55848 1934 56130
rect 1710 55792 1794 55848
rect 1850 55792 1934 55848
rect 1710 55510 1934 55792
rect 1710 55458 1796 55510
rect 1848 55458 1934 55510
rect 1710 55174 1934 55458
rect 1710 55122 1796 55174
rect 1848 55122 1934 55174
rect 1710 54838 1934 55122
rect 1710 54786 1796 54838
rect 1848 54786 1934 54838
rect 1710 54502 1934 54786
rect 1710 54450 1796 54502
rect 1848 54450 1934 54502
rect 1710 54168 1934 54450
rect 1710 54112 1794 54168
rect 1850 54112 1934 54168
rect 1710 53830 1934 54112
rect 1710 53778 1796 53830
rect 1848 53778 1934 53830
rect 1710 53494 1934 53778
rect 1710 53442 1796 53494
rect 1848 53442 1934 53494
rect 1710 53158 1934 53442
rect 1710 53106 1796 53158
rect 1848 53106 1934 53158
rect 1710 52822 1934 53106
rect 1710 52770 1796 52822
rect 1848 52770 1934 52822
rect 1710 52488 1934 52770
rect 1710 52432 1794 52488
rect 1850 52432 1934 52488
rect 1710 52150 1934 52432
rect 1710 52098 1796 52150
rect 1848 52098 1934 52150
rect 1710 51814 1934 52098
rect 1710 51762 1796 51814
rect 1848 51762 1934 51814
rect 1710 51478 1934 51762
rect 1710 51426 1796 51478
rect 1848 51426 1934 51478
rect 1710 51142 1934 51426
rect 1710 51090 1796 51142
rect 1848 51090 1934 51142
rect 1710 50808 1934 51090
rect 1710 50752 1794 50808
rect 1850 50752 1934 50808
rect 1710 50470 1934 50752
rect 1710 50418 1796 50470
rect 1848 50418 1934 50470
rect 1710 50134 1934 50418
rect 1710 50082 1796 50134
rect 1848 50082 1934 50134
rect 1710 49798 1934 50082
rect 1710 49746 1796 49798
rect 1848 49746 1934 49798
rect 1710 49462 1934 49746
rect 1710 49410 1796 49462
rect 1848 49410 1934 49462
rect 1710 49128 1934 49410
rect 1710 49072 1794 49128
rect 1850 49072 1934 49128
rect 1710 48790 1934 49072
rect 1710 48738 1796 48790
rect 1848 48738 1934 48790
rect 1710 48454 1934 48738
rect 1710 48402 1796 48454
rect 1848 48402 1934 48454
rect 1710 48118 1934 48402
rect 1710 48066 1796 48118
rect 1848 48066 1934 48118
rect 1710 47782 1934 48066
rect 1710 47730 1796 47782
rect 1848 47730 1934 47782
rect 1710 47448 1934 47730
rect 1710 47392 1794 47448
rect 1850 47392 1934 47448
rect 1710 47110 1934 47392
rect 1710 47058 1796 47110
rect 1848 47058 1934 47110
rect 1710 46774 1934 47058
rect 1710 46722 1796 46774
rect 1848 46722 1934 46774
rect 1710 46438 1934 46722
rect 1710 46386 1796 46438
rect 1848 46386 1934 46438
rect 1710 46102 1934 46386
rect 1710 46050 1796 46102
rect 1848 46050 1934 46102
rect 1710 45768 1934 46050
rect 1710 45712 1794 45768
rect 1850 45712 1934 45768
rect 1710 45430 1934 45712
rect 1710 45378 1796 45430
rect 1848 45378 1934 45430
rect 1710 45094 1934 45378
rect 1710 45042 1796 45094
rect 1848 45042 1934 45094
rect 1710 44758 1934 45042
rect 1710 44706 1796 44758
rect 1848 44706 1934 44758
rect 1710 44422 1934 44706
rect 1710 44370 1796 44422
rect 1848 44370 1934 44422
rect 1710 44088 1934 44370
rect 1710 44032 1794 44088
rect 1850 44032 1934 44088
rect 1710 43750 1934 44032
rect 1710 43698 1796 43750
rect 1848 43698 1934 43750
rect 1710 43414 1934 43698
rect 1710 43362 1796 43414
rect 1848 43362 1934 43414
rect 1710 43078 1934 43362
rect 1710 43026 1796 43078
rect 1848 43026 1934 43078
rect 1710 42742 1934 43026
rect 1710 42690 1796 42742
rect 1848 42690 1934 42742
rect 1710 42408 1934 42690
rect 1710 42352 1794 42408
rect 1850 42352 1934 42408
rect 1710 42070 1934 42352
rect 1710 42018 1796 42070
rect 1848 42018 1934 42070
rect 1710 41734 1934 42018
rect 1710 41682 1796 41734
rect 1848 41682 1934 41734
rect 1710 41398 1934 41682
rect 1710 41346 1796 41398
rect 1848 41346 1934 41398
rect 1710 41062 1934 41346
rect 1710 41010 1796 41062
rect 1848 41010 1934 41062
rect 1710 40728 1934 41010
rect 1710 40672 1794 40728
rect 1850 40672 1934 40728
rect 1710 40390 1934 40672
rect 1710 40338 1796 40390
rect 1848 40338 1934 40390
rect 1710 40054 1934 40338
rect 1710 40002 1796 40054
rect 1848 40002 1934 40054
rect 1710 39718 1934 40002
rect 1710 39666 1796 39718
rect 1848 39666 1934 39718
rect 1710 39382 1934 39666
rect 1710 39330 1796 39382
rect 1848 39330 1934 39382
rect 1710 39048 1934 39330
rect 1710 38992 1794 39048
rect 1850 38992 1934 39048
rect 1710 38710 1934 38992
rect 1710 38658 1796 38710
rect 1848 38658 1934 38710
rect 1710 38374 1934 38658
rect 1710 38322 1796 38374
rect 1848 38322 1934 38374
rect 1710 38038 1934 38322
rect 1710 37986 1796 38038
rect 1848 37986 1934 38038
rect 1710 37702 1934 37986
rect 1710 37650 1796 37702
rect 1848 37650 1934 37702
rect 1710 37368 1934 37650
rect 1710 37312 1794 37368
rect 1850 37312 1934 37368
rect 1710 37030 1934 37312
rect 1710 36978 1796 37030
rect 1848 36978 1934 37030
rect 1710 36694 1934 36978
rect 14613 36893 14669 36902
rect 13668 36822 13724 36831
rect 14613 36828 14669 36837
rect 15347 36893 15403 36902
rect 15347 36828 15403 36837
rect 13668 36757 13724 36766
rect 1710 36642 1796 36694
rect 1848 36642 1934 36694
rect 1710 36358 1934 36642
rect 1710 36306 1796 36358
rect 1848 36306 1934 36358
rect 1710 36022 1934 36306
rect 1710 35970 1796 36022
rect 1848 35970 1934 36022
rect 1710 35688 1934 35970
rect 1710 35632 1794 35688
rect 1850 35632 1934 35688
rect 1710 35350 1934 35632
rect 13668 35694 13724 35703
rect 13668 35629 13724 35638
rect 14613 35623 14669 35632
rect 14613 35558 14669 35567
rect 15267 35623 15323 35632
rect 15267 35558 15323 35567
rect 1710 35298 1796 35350
rect 1848 35298 1934 35350
rect 1710 35014 1934 35298
rect 1710 34962 1796 35014
rect 1848 34962 1934 35014
rect 1710 34678 1934 34962
rect 1710 34626 1796 34678
rect 1848 34626 1934 34678
rect 1710 34342 1934 34626
rect 1710 34290 1796 34342
rect 1848 34290 1934 34342
rect 1710 34008 1934 34290
rect 1710 33952 1794 34008
rect 1850 33952 1934 34008
rect 14613 34065 14669 34074
rect 1710 33670 1934 33952
rect 13668 33994 13724 34003
rect 14613 34000 14669 34009
rect 15187 34065 15243 34074
rect 15187 34000 15243 34009
rect 13668 33929 13724 33938
rect 1710 33618 1796 33670
rect 1848 33618 1934 33670
rect 1710 33334 1934 33618
rect 1710 33282 1796 33334
rect 1848 33282 1934 33334
rect 1710 32998 1934 33282
rect 1710 32946 1796 32998
rect 1848 32946 1934 32998
rect 1710 32662 1934 32946
rect 13668 32866 13724 32875
rect 13668 32801 13724 32810
rect 14613 32795 14669 32804
rect 14613 32730 14669 32739
rect 15107 32795 15163 32804
rect 15107 32730 15163 32739
rect 1710 32610 1796 32662
rect 1848 32610 1934 32662
rect 1710 32328 1934 32610
rect 1710 32272 1794 32328
rect 1850 32272 1934 32328
rect 1710 31990 1934 32272
rect 1710 31938 1796 31990
rect 1848 31938 1934 31990
rect 1710 31654 1934 31938
rect 1710 31602 1796 31654
rect 1848 31602 1934 31654
rect 1710 31318 1934 31602
rect 1710 31266 1796 31318
rect 1848 31266 1934 31318
rect 1710 30982 1934 31266
rect 14613 31237 14669 31246
rect 13668 31166 13724 31175
rect 14613 31172 14669 31181
rect 15027 31237 15083 31246
rect 15027 31172 15083 31181
rect 13668 31101 13724 31110
rect 1710 30930 1796 30982
rect 1848 30930 1934 30982
rect 1710 30648 1934 30930
rect 1710 30592 1794 30648
rect 1850 30592 1934 30648
rect 1710 30310 1934 30592
rect 1710 30258 1796 30310
rect 1848 30258 1934 30310
rect 1710 29974 1934 30258
rect 1710 29922 1796 29974
rect 1848 29922 1934 29974
rect 13668 30038 13724 30047
rect 13668 29973 13724 29982
rect 1710 29638 1934 29922
rect 14613 29967 14669 29976
rect 14613 29902 14669 29911
rect 14947 29967 15003 29976
rect 14947 29902 15003 29911
rect 1710 29586 1796 29638
rect 1848 29586 1934 29638
rect 1710 29302 1934 29586
rect 1710 29250 1796 29302
rect 1848 29250 1934 29302
rect 1710 28968 1934 29250
rect 1710 28912 1794 28968
rect 1850 28912 1934 28968
rect 1710 28630 1934 28912
rect 1710 28578 1796 28630
rect 1848 28578 1934 28630
rect 1710 28294 1934 28578
rect 14613 28409 14669 28418
rect 1710 28242 1796 28294
rect 1848 28242 1934 28294
rect 13668 28338 13724 28347
rect 14613 28344 14669 28353
rect 14867 28409 14923 28418
rect 14867 28344 14923 28353
rect 13668 28273 13724 28282
rect 1710 27958 1934 28242
rect 14750 28082 14806 28091
rect 14750 28017 14806 28026
rect 1710 27906 1796 27958
rect 1848 27906 1934 27958
rect 1710 27622 1934 27906
rect 1710 27570 1796 27622
rect 1848 27570 1934 27622
rect 1710 27288 1934 27570
rect 1710 27232 1794 27288
rect 1850 27232 1934 27288
rect 1710 26950 1934 27232
rect 1710 26898 1796 26950
rect 1848 26898 1934 26950
rect 1710 26614 1934 26898
rect 1710 26562 1796 26614
rect 1848 26562 1934 26614
rect 1710 26278 1934 26562
rect 1710 26226 1796 26278
rect 1848 26226 1934 26278
rect 1710 25942 1934 26226
rect 1710 25890 1796 25942
rect 1848 25890 1934 25942
rect 1710 25608 1934 25890
rect 1710 25552 1794 25608
rect 1850 25552 1934 25608
rect 1710 25270 1934 25552
rect 2541 25361 2597 25370
rect 2541 25296 2597 25305
rect 1710 25218 1796 25270
rect 1848 25218 1934 25270
rect 1710 24934 1934 25218
rect 1710 24882 1796 24934
rect 1848 24882 1934 24934
rect 1710 24598 1934 24882
rect 1710 24546 1796 24598
rect 1848 24546 1934 24598
rect 1710 24262 1934 24546
rect 1710 24210 1796 24262
rect 1848 24210 1934 24262
rect 1710 23928 1934 24210
rect 1710 23872 1794 23928
rect 1850 23872 1934 23928
rect 1710 23590 1934 23872
rect 1710 23538 1796 23590
rect 1848 23538 1934 23590
rect 1710 23254 1934 23538
rect 1710 23202 1796 23254
rect 1848 23202 1934 23254
rect 1710 22918 1934 23202
rect 1710 22866 1796 22918
rect 1848 22866 1934 22918
rect 1710 22582 1934 22866
rect 1710 22530 1796 22582
rect 1848 22530 1934 22582
rect 1710 22248 1934 22530
rect 1710 22192 1794 22248
rect 1850 22192 1934 22248
rect 1710 21910 1934 22192
rect 1710 21858 1796 21910
rect 1848 21858 1934 21910
rect 1710 21574 1934 21858
rect 1710 21522 1796 21574
rect 1848 21522 1934 21574
rect 1710 21238 1934 21522
rect 1710 21186 1796 21238
rect 1848 21186 1934 21238
rect 1710 20902 1934 21186
rect 1710 20850 1796 20902
rect 1848 20850 1934 20902
rect 1710 20568 1934 20850
rect 1710 20512 1794 20568
rect 1850 20512 1934 20568
rect 1710 20230 1934 20512
rect 1710 20178 1796 20230
rect 1848 20178 1934 20230
rect 1710 19894 1934 20178
rect 1710 19842 1796 19894
rect 1848 19842 1934 19894
rect 1710 19558 1934 19842
rect 1710 19506 1796 19558
rect 1848 19506 1934 19558
rect 1710 19222 1934 19506
rect 1710 19170 1796 19222
rect 1848 19170 1934 19222
rect 1710 18888 1934 19170
rect 1710 18832 1794 18888
rect 1850 18832 1934 18888
rect 1710 18550 1934 18832
rect 1710 18498 1796 18550
rect 1848 18498 1934 18550
rect 1710 18214 1934 18498
rect 1710 18162 1796 18214
rect 1848 18162 1934 18214
rect 14666 18253 14722 18262
rect 14666 18188 14722 18197
rect 1710 17878 1934 18162
rect 1710 17826 1796 17878
rect 1848 17826 1934 17878
rect 1710 17542 1934 17826
rect 1710 17490 1796 17542
rect 1848 17490 1934 17542
rect 1710 17208 1934 17490
rect 1710 17152 1794 17208
rect 1850 17152 1934 17208
rect 1710 16870 1934 17152
rect 1710 16818 1796 16870
rect 1848 16818 1934 16870
rect 1710 16534 1934 16818
rect 1710 16482 1796 16534
rect 1848 16482 1934 16534
rect 1710 16198 1934 16482
rect 1710 16146 1796 16198
rect 1848 16146 1934 16198
rect 1710 15862 1934 16146
rect 1710 15810 1796 15862
rect 1848 15810 1934 15862
rect 1710 15528 1934 15810
rect 1710 15472 1794 15528
rect 1850 15472 1934 15528
rect 1710 15190 1934 15472
rect 14666 15425 14722 15434
rect 14666 15360 14722 15369
rect 1710 15138 1796 15190
rect 1848 15138 1934 15190
rect 1710 14854 1934 15138
rect 1710 14802 1796 14854
rect 1848 14802 1934 14854
rect 1710 14518 1934 14802
rect 1710 14466 1796 14518
rect 1848 14466 1934 14518
rect 1710 14182 1934 14466
rect 1710 14130 1796 14182
rect 1848 14130 1934 14182
rect 1710 13848 1934 14130
rect 14666 14011 14722 14020
rect 14666 13946 14722 13955
rect 1710 13792 1794 13848
rect 1850 13792 1934 13848
rect 1710 13510 1934 13792
rect 1710 13458 1796 13510
rect 1848 13458 1934 13510
rect 1710 13174 1934 13458
rect 1710 13122 1796 13174
rect 1848 13122 1934 13174
rect 1710 12838 1934 13122
rect 1710 12786 1796 12838
rect 1848 12786 1934 12838
rect 1710 12502 1934 12786
rect 14666 12597 14722 12606
rect 14666 12532 14722 12541
rect 1710 12450 1796 12502
rect 1848 12450 1934 12502
rect 1710 12168 1934 12450
rect 1710 12112 1794 12168
rect 1850 12112 1934 12168
rect 1710 11830 1934 12112
rect 1710 11778 1796 11830
rect 1848 11778 1934 11830
rect 1710 11494 1934 11778
rect 1710 11442 1796 11494
rect 1848 11442 1934 11494
rect 1710 11158 1934 11442
rect 1710 11106 1796 11158
rect 1848 11106 1934 11158
rect 1710 10822 1934 11106
rect 1710 10770 1796 10822
rect 1848 10770 1934 10822
rect 1710 10488 1934 10770
rect 1710 10432 1794 10488
rect 1850 10432 1934 10488
rect 1710 10150 1934 10432
rect 1710 10098 1796 10150
rect 1848 10098 1934 10150
rect 1710 9814 1934 10098
rect 2754 9912 2810 9921
rect 2754 9847 2810 9856
rect 1710 9762 1796 9814
rect 1848 9762 1934 9814
rect 1710 9478 1934 9762
rect 1710 9426 1796 9478
rect 1848 9426 1934 9478
rect 1710 9142 1934 9426
rect 1710 9090 1796 9142
rect 1848 9090 1934 9142
rect 1710 8808 1934 9090
rect 1710 8752 1794 8808
rect 1850 8752 1934 8808
rect 1710 8470 1934 8752
rect 1710 8418 1796 8470
rect 1848 8418 1934 8470
rect 1710 8134 1934 8418
rect 14764 8341 14792 28017
rect 122202 19575 122230 79083
rect 134760 79030 134984 79312
rect 134760 78978 134846 79030
rect 134898 78978 134984 79030
rect 134760 78694 134984 78978
rect 134760 78642 134846 78694
rect 134898 78642 134984 78694
rect 134760 78358 134984 78642
rect 134760 78306 134846 78358
rect 134898 78306 134984 78358
rect 134760 78022 134984 78306
rect 134760 77970 134846 78022
rect 134898 77970 134984 78022
rect 134760 77688 134984 77970
rect 134760 77632 134844 77688
rect 134900 77632 134984 77688
rect 134760 77350 134984 77632
rect 134760 77298 134846 77350
rect 134898 77298 134984 77350
rect 134760 77014 134984 77298
rect 134760 76962 134846 77014
rect 134898 76962 134984 77014
rect 134760 76678 134984 76962
rect 134760 76626 134846 76678
rect 134898 76626 134984 76678
rect 134760 76342 134984 76626
rect 134760 76290 134846 76342
rect 134898 76290 134984 76342
rect 134760 76008 134984 76290
rect 134760 75952 134844 76008
rect 134900 75952 134984 76008
rect 134760 75670 134984 75952
rect 134760 75618 134846 75670
rect 134898 75618 134984 75670
rect 134760 75334 134984 75618
rect 134760 75282 134846 75334
rect 134898 75282 134984 75334
rect 134760 74998 134984 75282
rect 134760 74946 134846 74998
rect 134898 74946 134984 74998
rect 122272 74883 122328 74892
rect 122272 74818 122328 74827
rect 134760 74662 134984 74946
rect 134760 74610 134846 74662
rect 134898 74610 134984 74662
rect 134760 74328 134984 74610
rect 134760 74272 134844 74328
rect 134900 74272 134984 74328
rect 134760 73990 134984 74272
rect 134760 73938 134846 73990
rect 134898 73938 134984 73990
rect 134760 73654 134984 73938
rect 134760 73602 134846 73654
rect 134898 73602 134984 73654
rect 122272 73469 122328 73478
rect 122272 73404 122328 73413
rect 134760 73318 134984 73602
rect 134760 73266 134846 73318
rect 134898 73266 134984 73318
rect 134760 72982 134984 73266
rect 134760 72930 134846 72982
rect 134898 72930 134984 72982
rect 134760 72648 134984 72930
rect 134760 72592 134844 72648
rect 134900 72592 134984 72648
rect 134760 72310 134984 72592
rect 134760 72258 134846 72310
rect 134898 72258 134984 72310
rect 122272 72055 122328 72064
rect 122272 71990 122328 71999
rect 134760 71974 134984 72258
rect 134760 71922 134846 71974
rect 134898 71922 134984 71974
rect 134760 71638 134984 71922
rect 134760 71586 134846 71638
rect 134898 71586 134984 71638
rect 134760 71302 134984 71586
rect 134760 71250 134846 71302
rect 134898 71250 134984 71302
rect 134760 70968 134984 71250
rect 134760 70912 134844 70968
rect 134900 70912 134984 70968
rect 134760 70630 134984 70912
rect 134760 70578 134846 70630
rect 134898 70578 134984 70630
rect 134760 70294 134984 70578
rect 134760 70242 134846 70294
rect 134898 70242 134984 70294
rect 134760 69958 134984 70242
rect 134760 69906 134846 69958
rect 134898 69906 134984 69958
rect 134760 69622 134984 69906
rect 134760 69570 134846 69622
rect 134898 69570 134984 69622
rect 134760 69288 134984 69570
rect 134760 69232 134844 69288
rect 134900 69232 134984 69288
rect 134760 68950 134984 69232
rect 134760 68898 134846 68950
rect 134898 68898 134984 68950
rect 134760 68614 134984 68898
rect 134760 68562 134846 68614
rect 134898 68562 134984 68614
rect 134760 68278 134984 68562
rect 134760 68226 134846 68278
rect 134898 68226 134984 68278
rect 134760 67942 134984 68226
rect 134760 67890 134846 67942
rect 134898 67890 134984 67942
rect 134760 67608 134984 67890
rect 134760 67552 134844 67608
rect 134900 67552 134984 67608
rect 134760 67270 134984 67552
rect 134760 67218 134846 67270
rect 134898 67218 134984 67270
rect 134760 66934 134984 67218
rect 134760 66882 134846 66934
rect 134898 66882 134984 66934
rect 134760 66598 134984 66882
rect 134760 66546 134846 66598
rect 134898 66546 134984 66598
rect 134760 66262 134984 66546
rect 134760 66210 134846 66262
rect 134898 66210 134984 66262
rect 134760 65928 134984 66210
rect 134760 65872 134844 65928
rect 134900 65872 134984 65928
rect 134760 65590 134984 65872
rect 134760 65538 134846 65590
rect 134898 65538 134984 65590
rect 134760 65254 134984 65538
rect 134760 65202 134846 65254
rect 134898 65202 134984 65254
rect 134760 64918 134984 65202
rect 134760 64866 134846 64918
rect 134898 64866 134984 64918
rect 134760 64582 134984 64866
rect 134760 64530 134846 64582
rect 134898 64530 134984 64582
rect 134760 64248 134984 64530
rect 134760 64192 134844 64248
rect 134900 64192 134984 64248
rect 134760 63910 134984 64192
rect 134760 63858 134846 63910
rect 134898 63858 134984 63910
rect 134760 63574 134984 63858
rect 134760 63522 134846 63574
rect 134898 63522 134984 63574
rect 134760 63238 134984 63522
rect 134760 63186 134846 63238
rect 134898 63186 134984 63238
rect 134760 62902 134984 63186
rect 134760 62850 134846 62902
rect 134898 62850 134984 62902
rect 134760 62568 134984 62850
rect 134760 62512 134844 62568
rect 134900 62512 134984 62568
rect 134760 62230 134984 62512
rect 134760 62178 134846 62230
rect 134898 62178 134984 62230
rect 134097 62119 134153 62128
rect 134097 62054 134153 62063
rect 134760 61894 134984 62178
rect 134760 61842 134846 61894
rect 134898 61842 134984 61894
rect 134760 61558 134984 61842
rect 134760 61506 134846 61558
rect 134898 61506 134984 61558
rect 134760 61222 134984 61506
rect 134760 61170 134846 61222
rect 134898 61170 134984 61222
rect 134760 60888 134984 61170
rect 134760 60832 134844 60888
rect 134900 60832 134984 60888
rect 134760 60550 134984 60832
rect 134760 60498 134846 60550
rect 134898 60498 134984 60550
rect 134760 60214 134984 60498
rect 134760 60162 134846 60214
rect 134898 60162 134984 60214
rect 134760 59878 134984 60162
rect 134760 59826 134846 59878
rect 134898 59826 134984 59878
rect 134760 59542 134984 59826
rect 134760 59490 134846 59542
rect 134898 59490 134984 59542
rect 134760 59208 134984 59490
rect 134760 59152 134844 59208
rect 134900 59152 134984 59208
rect 134760 58870 134984 59152
rect 134760 58818 134846 58870
rect 134898 58818 134984 58870
rect 134760 58534 134984 58818
rect 134760 58482 134846 58534
rect 134898 58482 134984 58534
rect 134760 58198 134984 58482
rect 134760 58146 134846 58198
rect 134898 58146 134984 58198
rect 134760 57862 134984 58146
rect 134760 57810 134846 57862
rect 134898 57810 134984 57862
rect 134760 57528 134984 57810
rect 134760 57472 134844 57528
rect 134900 57472 134984 57528
rect 134760 57190 134984 57472
rect 134760 57138 134846 57190
rect 134898 57138 134984 57190
rect 134760 56854 134984 57138
rect 134760 56802 134846 56854
rect 134898 56802 134984 56854
rect 134760 56518 134984 56802
rect 134760 56466 134846 56518
rect 134898 56466 134984 56518
rect 134760 56182 134984 56466
rect 134760 56130 134846 56182
rect 134898 56130 134984 56182
rect 134760 55848 134984 56130
rect 134760 55792 134844 55848
rect 134900 55792 134984 55848
rect 134760 55510 134984 55792
rect 134760 55458 134846 55510
rect 134898 55458 134984 55510
rect 134760 55174 134984 55458
rect 134760 55122 134846 55174
rect 134898 55122 134984 55174
rect 134760 54838 134984 55122
rect 134760 54786 134846 54838
rect 134898 54786 134984 54838
rect 134760 54502 134984 54786
rect 134760 54450 134846 54502
rect 134898 54450 134984 54502
rect 134760 54168 134984 54450
rect 134760 54112 134844 54168
rect 134900 54112 134984 54168
rect 134760 53830 134984 54112
rect 134760 53778 134846 53830
rect 134898 53778 134984 53830
rect 134760 53494 134984 53778
rect 134760 53442 134846 53494
rect 134898 53442 134984 53494
rect 134760 53158 134984 53442
rect 134760 53106 134846 53158
rect 134898 53106 134984 53158
rect 134760 52822 134984 53106
rect 134760 52770 134846 52822
rect 134898 52770 134984 52822
rect 134760 52488 134984 52770
rect 134760 52432 134844 52488
rect 134900 52432 134984 52488
rect 134760 52150 134984 52432
rect 134760 52098 134846 52150
rect 134898 52098 134984 52150
rect 134760 51814 134984 52098
rect 134760 51762 134846 51814
rect 134898 51762 134984 51814
rect 134760 51478 134984 51762
rect 134760 51426 134846 51478
rect 134898 51426 134984 51478
rect 134760 51142 134984 51426
rect 134760 51090 134846 51142
rect 134898 51090 134984 51142
rect 134760 50808 134984 51090
rect 134760 50752 134844 50808
rect 134900 50752 134984 50808
rect 134760 50470 134984 50752
rect 134760 50418 134846 50470
rect 134898 50418 134984 50470
rect 134760 50134 134984 50418
rect 134760 50082 134846 50134
rect 134898 50082 134984 50134
rect 134760 49798 134984 50082
rect 134760 49746 134846 49798
rect 134898 49746 134984 49798
rect 134760 49462 134984 49746
rect 134760 49410 134846 49462
rect 134898 49410 134984 49462
rect 134760 49128 134984 49410
rect 134760 49072 134844 49128
rect 134900 49072 134984 49128
rect 134760 48790 134984 49072
rect 134760 48738 134846 48790
rect 134898 48738 134984 48790
rect 134760 48454 134984 48738
rect 134760 48402 134846 48454
rect 134898 48402 134984 48454
rect 134760 48118 134984 48402
rect 134760 48066 134846 48118
rect 134898 48066 134984 48118
rect 134760 47782 134984 48066
rect 134760 47730 134846 47782
rect 134898 47730 134984 47782
rect 134760 47448 134984 47730
rect 134760 47392 134844 47448
rect 134900 47392 134984 47448
rect 134760 47110 134984 47392
rect 134760 47058 134846 47110
rect 134898 47058 134984 47110
rect 134760 46774 134984 47058
rect 134760 46722 134846 46774
rect 134898 46722 134984 46774
rect 134760 46438 134984 46722
rect 134760 46386 134846 46438
rect 134898 46386 134984 46438
rect 134760 46102 134984 46386
rect 134760 46050 134846 46102
rect 134898 46050 134984 46102
rect 134760 45768 134984 46050
rect 134760 45712 134844 45768
rect 134900 45712 134984 45768
rect 134760 45430 134984 45712
rect 134760 45378 134846 45430
rect 134898 45378 134984 45430
rect 134760 45094 134984 45378
rect 134760 45042 134846 45094
rect 134898 45042 134984 45094
rect 134760 44758 134984 45042
rect 134760 44706 134846 44758
rect 134898 44706 134984 44758
rect 134760 44422 134984 44706
rect 134760 44370 134846 44422
rect 134898 44370 134984 44422
rect 134760 44088 134984 44370
rect 134760 44032 134844 44088
rect 134900 44032 134984 44088
rect 134760 43750 134984 44032
rect 134760 43698 134846 43750
rect 134898 43698 134984 43750
rect 134760 43414 134984 43698
rect 134760 43362 134846 43414
rect 134898 43362 134984 43414
rect 134760 43078 134984 43362
rect 134760 43026 134846 43078
rect 134898 43026 134984 43078
rect 134760 42742 134984 43026
rect 134760 42690 134846 42742
rect 134898 42690 134984 42742
rect 134760 42408 134984 42690
rect 134760 42352 134844 42408
rect 134900 42352 134984 42408
rect 134760 42070 134984 42352
rect 134760 42018 134846 42070
rect 134898 42018 134984 42070
rect 134760 41734 134984 42018
rect 134760 41682 134846 41734
rect 134898 41682 134984 41734
rect 134760 41398 134984 41682
rect 134760 41346 134846 41398
rect 134898 41346 134984 41398
rect 134760 41062 134984 41346
rect 134760 41010 134846 41062
rect 134898 41010 134984 41062
rect 134760 40728 134984 41010
rect 134760 40672 134844 40728
rect 134900 40672 134984 40728
rect 134760 40390 134984 40672
rect 134760 40338 134846 40390
rect 134898 40338 134984 40390
rect 134760 40054 134984 40338
rect 134760 40002 134846 40054
rect 134898 40002 134984 40054
rect 134760 39718 134984 40002
rect 134760 39666 134846 39718
rect 134898 39666 134984 39718
rect 134760 39382 134984 39666
rect 134760 39330 134846 39382
rect 134898 39330 134984 39382
rect 134760 39048 134984 39330
rect 134760 38992 134844 39048
rect 134900 38992 134984 39048
rect 134760 38710 134984 38992
rect 134760 38658 134846 38710
rect 134898 38658 134984 38710
rect 134760 38374 134984 38658
rect 134760 38322 134846 38374
rect 134898 38322 134984 38374
rect 134760 38038 134984 38322
rect 134760 37986 134846 38038
rect 134898 37986 134984 38038
rect 134760 37702 134984 37986
rect 134760 37650 134846 37702
rect 134898 37650 134984 37702
rect 134760 37368 134984 37650
rect 134760 37312 134844 37368
rect 134900 37312 134984 37368
rect 134760 37030 134984 37312
rect 134760 36978 134846 37030
rect 134898 36978 134984 37030
rect 134760 36694 134984 36978
rect 134760 36642 134846 36694
rect 134898 36642 134984 36694
rect 134760 36358 134984 36642
rect 134760 36306 134846 36358
rect 134898 36306 134984 36358
rect 134760 36022 134984 36306
rect 134760 35970 134846 36022
rect 134898 35970 134984 36022
rect 134760 35688 134984 35970
rect 134760 35632 134844 35688
rect 134900 35632 134984 35688
rect 134760 35350 134984 35632
rect 134760 35298 134846 35350
rect 134898 35298 134984 35350
rect 134760 35014 134984 35298
rect 134760 34962 134846 35014
rect 134898 34962 134984 35014
rect 134760 34678 134984 34962
rect 134760 34626 134846 34678
rect 134898 34626 134984 34678
rect 134760 34342 134984 34626
rect 134760 34290 134846 34342
rect 134898 34290 134984 34342
rect 134760 34008 134984 34290
rect 134760 33952 134844 34008
rect 134900 33952 134984 34008
rect 134760 33670 134984 33952
rect 134760 33618 134846 33670
rect 134898 33618 134984 33670
rect 134760 33334 134984 33618
rect 134760 33282 134846 33334
rect 134898 33282 134984 33334
rect 134760 32998 134984 33282
rect 134760 32946 134846 32998
rect 134898 32946 134984 32998
rect 134760 32662 134984 32946
rect 134760 32610 134846 32662
rect 134898 32610 134984 32662
rect 134760 32328 134984 32610
rect 134760 32272 134844 32328
rect 134900 32272 134984 32328
rect 134760 31990 134984 32272
rect 134760 31938 134846 31990
rect 134898 31938 134984 31990
rect 134760 31654 134984 31938
rect 134760 31602 134846 31654
rect 134898 31602 134984 31654
rect 134760 31318 134984 31602
rect 134760 31266 134846 31318
rect 134898 31266 134984 31318
rect 134760 30982 134984 31266
rect 134760 30930 134846 30982
rect 134898 30930 134984 30982
rect 134760 30648 134984 30930
rect 134760 30592 134844 30648
rect 134900 30592 134984 30648
rect 134760 30310 134984 30592
rect 134760 30258 134846 30310
rect 134898 30258 134984 30310
rect 134760 29974 134984 30258
rect 134760 29922 134846 29974
rect 134898 29922 134984 29974
rect 134760 29638 134984 29922
rect 134760 29586 134846 29638
rect 134898 29586 134984 29638
rect 134760 29302 134984 29586
rect 134760 29250 134846 29302
rect 134898 29250 134984 29302
rect 134760 28968 134984 29250
rect 134760 28912 134844 28968
rect 134900 28912 134984 28968
rect 134760 28630 134984 28912
rect 134760 28578 134846 28630
rect 134898 28578 134984 28630
rect 134760 28294 134984 28578
rect 134760 28242 134846 28294
rect 134898 28242 134984 28294
rect 134760 27958 134984 28242
rect 134760 27906 134846 27958
rect 134898 27906 134984 27958
rect 134760 27622 134984 27906
rect 134760 27570 134846 27622
rect 134898 27570 134984 27622
rect 134760 27288 134984 27570
rect 134760 27232 134844 27288
rect 134900 27232 134984 27288
rect 134760 26950 134984 27232
rect 134760 26898 134846 26950
rect 134898 26898 134984 26950
rect 134760 26614 134984 26898
rect 134760 26562 134846 26614
rect 134898 26562 134984 26614
rect 134760 26278 134984 26562
rect 134760 26226 134846 26278
rect 134898 26226 134984 26278
rect 134760 25942 134984 26226
rect 134760 25890 134846 25942
rect 134898 25890 134984 25942
rect 134760 25608 134984 25890
rect 134760 25552 134844 25608
rect 134900 25552 134984 25608
rect 134760 25270 134984 25552
rect 134760 25218 134846 25270
rect 134898 25218 134984 25270
rect 134760 24934 134984 25218
rect 134760 24882 134846 24934
rect 134898 24882 134984 24934
rect 134760 24598 134984 24882
rect 134760 24546 134846 24598
rect 134898 24546 134984 24598
rect 134760 24262 134984 24546
rect 134760 24210 134846 24262
rect 134898 24210 134984 24262
rect 134760 23928 134984 24210
rect 134760 23872 134844 23928
rect 134900 23872 134984 23928
rect 134760 23590 134984 23872
rect 134760 23538 134846 23590
rect 134898 23538 134984 23590
rect 134760 23254 134984 23538
rect 134760 23202 134846 23254
rect 134898 23202 134984 23254
rect 134760 22918 134984 23202
rect 134760 22866 134846 22918
rect 134898 22866 134984 22918
rect 134760 22582 134984 22866
rect 134760 22530 134846 22582
rect 134898 22530 134984 22582
rect 134760 22248 134984 22530
rect 134760 22192 134844 22248
rect 134900 22192 134984 22248
rect 134760 21910 134984 22192
rect 134760 21858 134846 21910
rect 134898 21858 134984 21910
rect 134760 21574 134984 21858
rect 134760 21522 134846 21574
rect 134898 21522 134984 21574
rect 134760 21238 134984 21522
rect 134760 21186 134846 21238
rect 134898 21186 134984 21238
rect 134760 20902 134984 21186
rect 134760 20850 134846 20902
rect 134898 20850 134984 20902
rect 134760 20568 134984 20850
rect 134760 20512 134844 20568
rect 134900 20512 134984 20568
rect 134760 20230 134984 20512
rect 134760 20178 134846 20230
rect 134898 20178 134984 20230
rect 134760 19894 134984 20178
rect 134760 19842 134846 19894
rect 134898 19842 134984 19894
rect 122188 19566 122244 19575
rect 22822 18262 22850 19547
rect 122188 19501 122244 19510
rect 134760 19558 134984 19842
rect 134760 19506 134846 19558
rect 134898 19506 134984 19558
rect 123270 19310 123326 19319
rect 121987 19239 122043 19248
rect 121987 19174 122043 19183
rect 122325 19239 122381 19248
rect 123270 19245 123326 19254
rect 122325 19174 122381 19183
rect 134760 19222 134984 19506
rect 134760 19170 134846 19222
rect 134898 19170 134984 19222
rect 22808 18253 22864 18262
rect 22808 18188 22864 18197
rect 26525 15434 26553 19070
rect 134760 18888 134984 19170
rect 134760 18832 134844 18888
rect 134900 18832 134984 18888
rect 134760 18550 134984 18832
rect 134760 18498 134846 18550
rect 134898 18498 134984 18550
rect 134760 18214 134984 18498
rect 134760 18162 134846 18214
rect 134898 18162 134984 18214
rect 134760 17878 134984 18162
rect 134760 17826 134846 17878
rect 134898 17826 134984 17878
rect 121907 17681 121963 17690
rect 121907 17616 121963 17625
rect 122325 17681 122381 17690
rect 122325 17616 122381 17625
rect 123270 17610 123326 17619
rect 123270 17545 123326 17554
rect 134760 17542 134984 17826
rect 134760 17490 134846 17542
rect 134898 17490 134984 17542
rect 134760 17208 134984 17490
rect 134760 17152 134844 17208
rect 134900 17152 134984 17208
rect 134760 16870 134984 17152
rect 134760 16818 134846 16870
rect 134898 16818 134984 16870
rect 134760 16534 134984 16818
rect 123270 16482 123326 16491
rect 121827 16411 121883 16420
rect 121827 16346 121883 16355
rect 122325 16411 122381 16420
rect 123270 16417 123326 16426
rect 134760 16482 134846 16534
rect 134898 16482 134984 16534
rect 122325 16346 122381 16355
rect 134760 16198 134984 16482
rect 134760 16146 134846 16198
rect 134898 16146 134984 16198
rect 134760 15862 134984 16146
rect 134760 15810 134846 15862
rect 134898 15810 134984 15862
rect 134760 15528 134984 15810
rect 134760 15472 134844 15528
rect 134900 15472 134984 15528
rect 26511 15425 26567 15434
rect 26511 15360 26567 15369
rect 134760 15190 134984 15472
rect 134760 15138 134846 15190
rect 134898 15138 134984 15190
rect 121747 14853 121803 14862
rect 121747 14788 121803 14797
rect 122325 14853 122381 14862
rect 122325 14788 122381 14797
rect 134760 14854 134984 15138
rect 134760 14802 134846 14854
rect 134898 14802 134984 14854
rect 123270 14782 123326 14791
rect 123270 14717 123326 14726
rect 134760 14518 134984 14802
rect 134760 14466 134846 14518
rect 134898 14466 134984 14518
rect 134760 14182 134984 14466
rect 134760 14130 134846 14182
rect 134898 14130 134984 14182
rect 26759 14011 26815 14020
rect 26759 13946 26815 13955
rect 26635 12597 26691 12606
rect 26635 12532 26691 12541
rect 26649 9457 26677 12532
rect 26773 9457 26801 13946
rect 134760 13848 134984 14130
rect 134760 13792 134844 13848
rect 134900 13792 134984 13848
rect 123270 13654 123326 13663
rect 121667 13583 121723 13592
rect 121667 13518 121723 13527
rect 122325 13583 122381 13592
rect 123270 13589 123326 13598
rect 122325 13518 122381 13527
rect 134760 13510 134984 13792
rect 134760 13458 134846 13510
rect 134898 13458 134984 13510
rect 28618 13261 28674 13270
rect 28618 13196 28674 13205
rect 31114 13261 31170 13270
rect 31114 13196 31170 13205
rect 33610 13261 33666 13270
rect 33610 13196 33666 13205
rect 36106 13261 36162 13270
rect 36106 13196 36162 13205
rect 38602 13261 38658 13270
rect 38602 13196 38658 13205
rect 41098 13261 41154 13270
rect 41098 13196 41154 13205
rect 43594 13261 43650 13270
rect 43594 13196 43650 13205
rect 46090 13261 46146 13270
rect 46090 13196 46146 13205
rect 48586 13261 48642 13270
rect 48586 13196 48642 13205
rect 51082 13261 51138 13270
rect 51082 13196 51138 13205
rect 53578 13261 53634 13270
rect 53578 13196 53634 13205
rect 56074 13261 56130 13270
rect 56074 13196 56130 13205
rect 58570 13261 58626 13270
rect 58570 13196 58626 13205
rect 61066 13261 61122 13270
rect 61066 13196 61122 13205
rect 63562 13261 63618 13270
rect 63562 13196 63618 13205
rect 66058 13261 66114 13270
rect 66058 13196 66114 13205
rect 68554 13261 68610 13270
rect 68554 13196 68610 13205
rect 71050 13261 71106 13270
rect 71050 13196 71106 13205
rect 73546 13261 73602 13270
rect 73546 13196 73602 13205
rect 76042 13261 76098 13270
rect 76042 13196 76098 13205
rect 78538 13261 78594 13270
rect 78538 13196 78594 13205
rect 81034 13261 81090 13270
rect 81034 13196 81090 13205
rect 83530 13261 83586 13270
rect 83530 13196 83586 13205
rect 86026 13261 86082 13270
rect 86026 13196 86082 13205
rect 88522 13261 88578 13270
rect 88522 13196 88578 13205
rect 91018 13261 91074 13270
rect 91018 13196 91074 13205
rect 93514 13261 93570 13270
rect 93514 13196 93570 13205
rect 96010 13261 96066 13270
rect 96010 13196 96066 13205
rect 98506 13261 98562 13270
rect 98506 13196 98562 13205
rect 101002 13261 101058 13270
rect 101002 13196 101058 13205
rect 103498 13261 103554 13270
rect 103498 13196 103554 13205
rect 105994 13261 106050 13270
rect 105994 13196 106050 13205
rect 134760 13174 134984 13458
rect 134760 13122 134846 13174
rect 134898 13122 134984 13174
rect 134760 12838 134984 13122
rect 134760 12786 134846 12838
rect 134898 12786 134984 12838
rect 134760 12502 134984 12786
rect 134760 12450 134846 12502
rect 134898 12450 134984 12502
rect 134760 12168 134984 12450
rect 134760 12112 134844 12168
rect 134900 12112 134984 12168
rect 121587 12025 121643 12034
rect 121587 11960 121643 11969
rect 122325 12025 122381 12034
rect 122325 11960 122381 11969
rect 123270 11954 123326 11963
rect 123270 11889 123326 11898
rect 134760 11830 134984 12112
rect 134760 11778 134846 11830
rect 134898 11778 134984 11830
rect 134760 11494 134984 11778
rect 134760 11442 134846 11494
rect 134898 11442 134984 11494
rect 134760 11158 134984 11442
rect 134760 11106 134846 11158
rect 134898 11106 134984 11158
rect 123270 10826 123326 10835
rect 121507 10755 121563 10764
rect 121507 10690 121563 10699
rect 122325 10755 122381 10764
rect 123270 10761 123326 10770
rect 134760 10822 134984 11106
rect 134760 10770 134846 10822
rect 134898 10770 134984 10822
rect 122325 10690 122381 10699
rect 134760 10488 134984 10770
rect 134760 10432 134844 10488
rect 134900 10432 134984 10488
rect 134760 10150 134984 10432
rect 134760 10098 134846 10150
rect 134898 10098 134984 10150
rect 134760 9814 134984 10098
rect 134760 9762 134846 9814
rect 134898 9762 134984 9814
rect 134760 9478 134984 9762
rect 5975 8317 6031 8326
rect 14694 8313 14792 8341
rect 5975 8252 6031 8261
rect 2754 8212 2810 8221
rect 2754 8147 2810 8156
rect 1710 8082 1796 8134
rect 1848 8082 1934 8134
rect 1710 7798 1934 8082
rect 1710 7746 1796 7798
rect 1848 7746 1934 7798
rect 1710 7462 1934 7746
rect 1710 7410 1796 7462
rect 1848 7410 1934 7462
rect 1710 7128 1934 7410
rect 1710 7072 1794 7128
rect 1850 7072 1934 7128
rect 1710 6790 1934 7072
rect 1710 6738 1796 6790
rect 1848 6738 1934 6790
rect 1710 6454 1934 6738
rect 1710 6402 1796 6454
rect 1848 6402 1934 6454
rect 1710 6118 1934 6402
rect 1710 6066 1796 6118
rect 1848 6066 1934 6118
rect 1710 5782 1934 6066
rect 1710 5730 1796 5782
rect 1848 5730 1934 5782
rect 1710 5448 1934 5730
rect 1710 5392 1794 5448
rect 1850 5392 1934 5448
rect 1710 5110 1934 5392
rect 1710 5058 1796 5110
rect 1848 5058 1934 5110
rect 1710 4774 1934 5058
rect 1710 4722 1796 4774
rect 1848 4722 1934 4774
rect 1710 4438 1934 4722
rect 1710 4386 1796 4438
rect 1848 4386 1934 4438
rect 1710 4102 1934 4386
rect 1710 4050 1796 4102
rect 1848 4050 1934 4102
rect 1710 3768 1934 4050
rect 1710 3712 1794 3768
rect 1850 3712 1934 3768
rect 1710 3430 1934 3712
rect 1710 3378 1796 3430
rect 1848 3378 1934 3430
rect 1710 3094 1934 3378
rect 1710 3042 1796 3094
rect 1848 3042 1934 3094
rect 1710 2758 1934 3042
rect 1710 2706 1796 2758
rect 1848 2706 1934 2758
rect 14764 2741 14792 8313
rect 134760 9426 134846 9478
rect 134898 9426 134984 9478
rect 134760 9142 134984 9426
rect 134760 9090 134846 9142
rect 134898 9090 134984 9142
rect 134760 8808 134984 9090
rect 134760 8752 134844 8808
rect 134900 8752 134984 8808
rect 134760 8470 134984 8752
rect 134760 8418 134846 8470
rect 134898 8418 134984 8470
rect 134760 8134 134984 8418
rect 134760 8082 134846 8134
rect 134898 8082 134984 8134
rect 134760 7798 134984 8082
rect 134760 7746 134846 7798
rect 134898 7746 134984 7798
rect 134760 7462 134984 7746
rect 134760 7410 134846 7462
rect 134898 7410 134984 7462
rect 134760 7128 134984 7410
rect 134760 7072 134844 7128
rect 134900 7072 134984 7128
rect 134760 6790 134984 7072
rect 134760 6738 134846 6790
rect 134898 6738 134984 6790
rect 134760 6454 134984 6738
rect 134760 6402 134846 6454
rect 134898 6402 134984 6454
rect 134760 6118 134984 6402
rect 134760 6066 134846 6118
rect 134898 6066 134984 6118
rect 134760 5782 134984 6066
rect 134760 5730 134846 5782
rect 134898 5730 134984 5782
rect 134760 5448 134984 5730
rect 134760 5392 134844 5448
rect 134900 5392 134984 5448
rect 134760 5110 134984 5392
rect 134760 5058 134846 5110
rect 134898 5058 134984 5110
rect 134760 4774 134984 5058
rect 134760 4722 134846 4774
rect 134898 4722 134984 4774
rect 134760 4438 134984 4722
rect 134760 4386 134846 4438
rect 134898 4386 134984 4438
rect 134760 4102 134984 4386
rect 134760 4050 134846 4102
rect 134898 4050 134984 4102
rect 134760 3768 134984 4050
rect 134760 3712 134844 3768
rect 134900 3712 134984 3768
rect 134760 3430 134984 3712
rect 134760 3378 134846 3430
rect 134898 3378 134984 3430
rect 134760 3094 134984 3378
rect 134760 3042 134846 3094
rect 134898 3042 134984 3094
rect 16004 2988 16060 2997
rect 16004 2923 16060 2932
rect 17172 2988 17228 2997
rect 17172 2923 17228 2932
rect 18340 2988 18396 2997
rect 18340 2923 18396 2932
rect 19508 2988 19564 2997
rect 19508 2923 19564 2932
rect 20676 2988 20732 2997
rect 20676 2923 20732 2932
rect 21844 2988 21900 2997
rect 21844 2923 21900 2932
rect 23012 2988 23068 2997
rect 23012 2923 23068 2932
rect 24180 2988 24236 2997
rect 24180 2923 24236 2932
rect 25348 2988 25404 2997
rect 25348 2923 25404 2932
rect 26516 2988 26572 2997
rect 26516 2923 26572 2932
rect 27684 2988 27740 2997
rect 27684 2923 27740 2932
rect 28852 2988 28908 2997
rect 28852 2923 28908 2932
rect 30020 2988 30076 2997
rect 30020 2923 30076 2932
rect 31188 2988 31244 2997
rect 31188 2923 31244 2932
rect 32356 2988 32412 2997
rect 32356 2923 32412 2932
rect 33524 2988 33580 2997
rect 33524 2923 33580 2932
rect 34692 2988 34748 2997
rect 34692 2923 34748 2932
rect 35860 2988 35916 2997
rect 35860 2923 35916 2932
rect 37028 2988 37084 2997
rect 37028 2923 37084 2932
rect 38196 2988 38252 2997
rect 38196 2923 38252 2932
rect 39364 2988 39420 2997
rect 39364 2923 39420 2932
rect 40532 2988 40588 2997
rect 40532 2923 40588 2932
rect 41700 2988 41756 2997
rect 41700 2923 41756 2932
rect 42868 2988 42924 2997
rect 42868 2923 42924 2932
rect 44036 2988 44092 2997
rect 44036 2923 44092 2932
rect 45204 2988 45260 2997
rect 45204 2923 45260 2932
rect 46372 2988 46428 2997
rect 46372 2923 46428 2932
rect 47540 2988 47596 2997
rect 47540 2923 47596 2932
rect 48708 2988 48764 2997
rect 48708 2923 48764 2932
rect 49876 2988 49932 2997
rect 49876 2923 49932 2932
rect 51044 2988 51100 2997
rect 51044 2923 51100 2932
rect 52212 2988 52268 2997
rect 52212 2923 52268 2932
rect 53380 2988 53436 2997
rect 53380 2923 53436 2932
rect 54548 2988 54604 2997
rect 54548 2923 54604 2932
rect 55716 2988 55772 2997
rect 55716 2923 55772 2932
rect 56884 2988 56940 2997
rect 56884 2923 56940 2932
rect 58052 2988 58108 2997
rect 58052 2923 58108 2932
rect 59220 2988 59276 2997
rect 59220 2923 59276 2932
rect 134760 2758 134984 3042
rect 1710 2422 1934 2706
rect 14750 2732 14806 2741
rect 14750 2667 14806 2676
rect 134760 2706 134846 2758
rect 134898 2706 134984 2758
rect 1710 2370 1796 2422
rect 1848 2370 1934 2422
rect 1710 2088 1934 2370
rect 1710 2032 1794 2088
rect 1850 2032 1934 2088
rect 1710 1612 1934 2032
rect 134760 2422 134984 2706
rect 134760 2370 134846 2422
rect 134898 2370 134984 2422
rect 134760 2088 134984 2370
rect 134760 2032 134844 2088
rect 134900 2032 134984 2088
rect 2130 1752 2186 1761
rect 2130 1687 2186 1696
rect 3810 1752 3866 1761
rect 3810 1687 3866 1696
rect 5490 1752 5546 1761
rect 5490 1687 5546 1696
rect 7170 1752 7226 1761
rect 7170 1687 7226 1696
rect 8850 1752 8906 1761
rect 8850 1687 8906 1696
rect 10530 1752 10586 1761
rect 10530 1687 10586 1696
rect 12210 1752 12266 1761
rect 12210 1687 12266 1696
rect 13890 1752 13946 1761
rect 13890 1687 13946 1696
rect 15570 1752 15626 1761
rect 15570 1687 15626 1696
rect 17250 1752 17306 1761
rect 17250 1687 17306 1696
rect 18930 1752 18986 1761
rect 18930 1687 18986 1696
rect 20610 1752 20666 1761
rect 20610 1687 20666 1696
rect 22290 1752 22346 1761
rect 22290 1687 22346 1696
rect 23970 1752 24026 1761
rect 23970 1687 24026 1696
rect 25650 1752 25706 1761
rect 25650 1687 25706 1696
rect 27330 1752 27386 1761
rect 27330 1687 27386 1696
rect 29010 1752 29066 1761
rect 29010 1687 29066 1696
rect 30690 1752 30746 1761
rect 30690 1687 30746 1696
rect 32370 1752 32426 1761
rect 32370 1687 32426 1696
rect 34050 1752 34106 1761
rect 34050 1687 34106 1696
rect 35730 1752 35786 1761
rect 35730 1687 35786 1696
rect 37410 1752 37466 1761
rect 37410 1687 37466 1696
rect 39090 1752 39146 1761
rect 39090 1687 39146 1696
rect 40770 1752 40826 1761
rect 40770 1687 40826 1696
rect 42450 1752 42506 1761
rect 42450 1687 42506 1696
rect 44130 1752 44186 1761
rect 44130 1687 44186 1696
rect 45810 1752 45866 1761
rect 45810 1687 45866 1696
rect 47490 1752 47546 1761
rect 47490 1687 47546 1696
rect 49170 1752 49226 1761
rect 49170 1687 49226 1696
rect 50850 1752 50906 1761
rect 50850 1687 50906 1696
rect 52530 1752 52586 1761
rect 52530 1687 52586 1696
rect 54210 1752 54266 1761
rect 54210 1687 54266 1696
rect 55890 1752 55946 1761
rect 55890 1687 55946 1696
rect 57570 1752 57626 1761
rect 57570 1687 57626 1696
rect 59250 1752 59306 1761
rect 59250 1687 59306 1696
rect 60930 1752 60986 1761
rect 60930 1687 60986 1696
rect 62610 1752 62666 1761
rect 62610 1687 62666 1696
rect 64290 1752 64346 1761
rect 64290 1687 64346 1696
rect 65970 1752 66026 1761
rect 65970 1687 66026 1696
rect 67650 1752 67706 1761
rect 67650 1687 67706 1696
rect 69330 1752 69386 1761
rect 69330 1687 69386 1696
rect 71010 1752 71066 1761
rect 71010 1687 71066 1696
rect 72690 1752 72746 1761
rect 72690 1687 72746 1696
rect 74370 1752 74426 1761
rect 74370 1687 74426 1696
rect 76050 1752 76106 1761
rect 76050 1687 76106 1696
rect 77730 1752 77786 1761
rect 77730 1687 77786 1696
rect 79410 1752 79466 1761
rect 79410 1687 79466 1696
rect 81090 1752 81146 1761
rect 81090 1687 81146 1696
rect 82770 1752 82826 1761
rect 82770 1687 82826 1696
rect 84450 1752 84506 1761
rect 84450 1687 84506 1696
rect 86130 1752 86186 1761
rect 86130 1687 86186 1696
rect 87810 1752 87866 1761
rect 87810 1687 87866 1696
rect 89490 1752 89546 1761
rect 89490 1687 89546 1696
rect 91170 1752 91226 1761
rect 91170 1687 91226 1696
rect 92850 1752 92906 1761
rect 92850 1687 92906 1696
rect 94530 1752 94586 1761
rect 94530 1687 94586 1696
rect 96210 1752 96266 1761
rect 96210 1687 96266 1696
rect 97890 1752 97946 1761
rect 97890 1687 97946 1696
rect 99570 1752 99626 1761
rect 99570 1687 99626 1696
rect 101250 1752 101306 1761
rect 101250 1687 101306 1696
rect 102930 1752 102986 1761
rect 102930 1687 102986 1696
rect 104610 1752 104666 1761
rect 104610 1687 104666 1696
rect 106290 1752 106346 1761
rect 106290 1687 106346 1696
rect 107970 1752 108026 1761
rect 107970 1687 108026 1696
rect 109650 1752 109706 1761
rect 109650 1687 109706 1696
rect 111330 1752 111386 1761
rect 111330 1687 111386 1696
rect 113010 1752 113066 1761
rect 113010 1687 113066 1696
rect 114690 1752 114746 1761
rect 114690 1687 114746 1696
rect 116370 1752 116426 1761
rect 116370 1687 116426 1696
rect 118050 1752 118106 1761
rect 118050 1687 118106 1696
rect 119730 1752 119786 1761
rect 119730 1687 119786 1696
rect 121410 1752 121466 1761
rect 121410 1687 121466 1696
rect 123090 1752 123146 1761
rect 123090 1687 123146 1696
rect 124770 1752 124826 1761
rect 124770 1687 124826 1696
rect 126450 1752 126506 1761
rect 126450 1687 126506 1696
rect 128130 1752 128186 1761
rect 128130 1687 128186 1696
rect 129810 1752 129866 1761
rect 129810 1687 129866 1696
rect 131490 1752 131546 1761
rect 131490 1687 131546 1696
rect 133170 1752 133226 1761
rect 133170 1687 133226 1696
rect 134760 1612 134984 2032
<< via2 >>
rect 2130 81499 2186 81501
rect 2130 81447 2132 81499
rect 2132 81447 2184 81499
rect 2184 81447 2186 81499
rect 2130 81445 2186 81447
rect 3810 81499 3866 81501
rect 3810 81447 3812 81499
rect 3812 81447 3864 81499
rect 3864 81447 3866 81499
rect 3810 81445 3866 81447
rect 5490 81499 5546 81501
rect 5490 81447 5492 81499
rect 5492 81447 5544 81499
rect 5544 81447 5546 81499
rect 5490 81445 5546 81447
rect 7170 81499 7226 81501
rect 7170 81447 7172 81499
rect 7172 81447 7224 81499
rect 7224 81447 7226 81499
rect 7170 81445 7226 81447
rect 8850 81499 8906 81501
rect 8850 81447 8852 81499
rect 8852 81447 8904 81499
rect 8904 81447 8906 81499
rect 8850 81445 8906 81447
rect 10530 81499 10586 81501
rect 10530 81447 10532 81499
rect 10532 81447 10584 81499
rect 10584 81447 10586 81499
rect 10530 81445 10586 81447
rect 12210 81499 12266 81501
rect 12210 81447 12212 81499
rect 12212 81447 12264 81499
rect 12264 81447 12266 81499
rect 12210 81445 12266 81447
rect 13890 81499 13946 81501
rect 13890 81447 13892 81499
rect 13892 81447 13944 81499
rect 13944 81447 13946 81499
rect 13890 81445 13946 81447
rect 15570 81499 15626 81501
rect 15570 81447 15572 81499
rect 15572 81447 15624 81499
rect 15624 81447 15626 81499
rect 15570 81445 15626 81447
rect 17250 81499 17306 81501
rect 17250 81447 17252 81499
rect 17252 81447 17304 81499
rect 17304 81447 17306 81499
rect 17250 81445 17306 81447
rect 18930 81499 18986 81501
rect 18930 81447 18932 81499
rect 18932 81447 18984 81499
rect 18984 81447 18986 81499
rect 18930 81445 18986 81447
rect 20610 81499 20666 81501
rect 20610 81447 20612 81499
rect 20612 81447 20664 81499
rect 20664 81447 20666 81499
rect 20610 81445 20666 81447
rect 22290 81499 22346 81501
rect 22290 81447 22292 81499
rect 22292 81447 22344 81499
rect 22344 81447 22346 81499
rect 22290 81445 22346 81447
rect 23970 81499 24026 81501
rect 23970 81447 23972 81499
rect 23972 81447 24024 81499
rect 24024 81447 24026 81499
rect 23970 81445 24026 81447
rect 25650 81499 25706 81501
rect 25650 81447 25652 81499
rect 25652 81447 25704 81499
rect 25704 81447 25706 81499
rect 25650 81445 25706 81447
rect 27330 81499 27386 81501
rect 27330 81447 27332 81499
rect 27332 81447 27384 81499
rect 27384 81447 27386 81499
rect 27330 81445 27386 81447
rect 29010 81499 29066 81501
rect 29010 81447 29012 81499
rect 29012 81447 29064 81499
rect 29064 81447 29066 81499
rect 29010 81445 29066 81447
rect 30690 81499 30746 81501
rect 30690 81447 30692 81499
rect 30692 81447 30744 81499
rect 30744 81447 30746 81499
rect 30690 81445 30746 81447
rect 32370 81499 32426 81501
rect 32370 81447 32372 81499
rect 32372 81447 32424 81499
rect 32424 81447 32426 81499
rect 32370 81445 32426 81447
rect 34050 81499 34106 81501
rect 34050 81447 34052 81499
rect 34052 81447 34104 81499
rect 34104 81447 34106 81499
rect 34050 81445 34106 81447
rect 35730 81499 35786 81501
rect 35730 81447 35732 81499
rect 35732 81447 35784 81499
rect 35784 81447 35786 81499
rect 35730 81445 35786 81447
rect 37410 81499 37466 81501
rect 37410 81447 37412 81499
rect 37412 81447 37464 81499
rect 37464 81447 37466 81499
rect 37410 81445 37466 81447
rect 39090 81499 39146 81501
rect 39090 81447 39092 81499
rect 39092 81447 39144 81499
rect 39144 81447 39146 81499
rect 39090 81445 39146 81447
rect 40770 81499 40826 81501
rect 40770 81447 40772 81499
rect 40772 81447 40824 81499
rect 40824 81447 40826 81499
rect 40770 81445 40826 81447
rect 42450 81499 42506 81501
rect 42450 81447 42452 81499
rect 42452 81447 42504 81499
rect 42504 81447 42506 81499
rect 42450 81445 42506 81447
rect 44130 81499 44186 81501
rect 44130 81447 44132 81499
rect 44132 81447 44184 81499
rect 44184 81447 44186 81499
rect 44130 81445 44186 81447
rect 45810 81499 45866 81501
rect 45810 81447 45812 81499
rect 45812 81447 45864 81499
rect 45864 81447 45866 81499
rect 45810 81445 45866 81447
rect 47490 81499 47546 81501
rect 47490 81447 47492 81499
rect 47492 81447 47544 81499
rect 47544 81447 47546 81499
rect 47490 81445 47546 81447
rect 49170 81499 49226 81501
rect 49170 81447 49172 81499
rect 49172 81447 49224 81499
rect 49224 81447 49226 81499
rect 49170 81445 49226 81447
rect 50850 81499 50906 81501
rect 50850 81447 50852 81499
rect 50852 81447 50904 81499
rect 50904 81447 50906 81499
rect 50850 81445 50906 81447
rect 52530 81499 52586 81501
rect 52530 81447 52532 81499
rect 52532 81447 52584 81499
rect 52584 81447 52586 81499
rect 52530 81445 52586 81447
rect 54210 81499 54266 81501
rect 54210 81447 54212 81499
rect 54212 81447 54264 81499
rect 54264 81447 54266 81499
rect 54210 81445 54266 81447
rect 55890 81499 55946 81501
rect 55890 81447 55892 81499
rect 55892 81447 55944 81499
rect 55944 81447 55946 81499
rect 55890 81445 55946 81447
rect 57570 81499 57626 81501
rect 57570 81447 57572 81499
rect 57572 81447 57624 81499
rect 57624 81447 57626 81499
rect 57570 81445 57626 81447
rect 59250 81499 59306 81501
rect 59250 81447 59252 81499
rect 59252 81447 59304 81499
rect 59304 81447 59306 81499
rect 59250 81445 59306 81447
rect 60930 81499 60986 81501
rect 60930 81447 60932 81499
rect 60932 81447 60984 81499
rect 60984 81447 60986 81499
rect 60930 81445 60986 81447
rect 62610 81499 62666 81501
rect 62610 81447 62612 81499
rect 62612 81447 62664 81499
rect 62664 81447 62666 81499
rect 62610 81445 62666 81447
rect 64290 81499 64346 81501
rect 64290 81447 64292 81499
rect 64292 81447 64344 81499
rect 64344 81447 64346 81499
rect 64290 81445 64346 81447
rect 65970 81499 66026 81501
rect 65970 81447 65972 81499
rect 65972 81447 66024 81499
rect 66024 81447 66026 81499
rect 65970 81445 66026 81447
rect 67650 81499 67706 81501
rect 67650 81447 67652 81499
rect 67652 81447 67704 81499
rect 67704 81447 67706 81499
rect 67650 81445 67706 81447
rect 69330 81499 69386 81501
rect 69330 81447 69332 81499
rect 69332 81447 69384 81499
rect 69384 81447 69386 81499
rect 69330 81445 69386 81447
rect 71010 81499 71066 81501
rect 71010 81447 71012 81499
rect 71012 81447 71064 81499
rect 71064 81447 71066 81499
rect 71010 81445 71066 81447
rect 72690 81499 72746 81501
rect 72690 81447 72692 81499
rect 72692 81447 72744 81499
rect 72744 81447 72746 81499
rect 72690 81445 72746 81447
rect 74370 81499 74426 81501
rect 74370 81447 74372 81499
rect 74372 81447 74424 81499
rect 74424 81447 74426 81499
rect 74370 81445 74426 81447
rect 76050 81499 76106 81501
rect 76050 81447 76052 81499
rect 76052 81447 76104 81499
rect 76104 81447 76106 81499
rect 76050 81445 76106 81447
rect 77730 81499 77786 81501
rect 77730 81447 77732 81499
rect 77732 81447 77784 81499
rect 77784 81447 77786 81499
rect 77730 81445 77786 81447
rect 79410 81499 79466 81501
rect 79410 81447 79412 81499
rect 79412 81447 79464 81499
rect 79464 81447 79466 81499
rect 79410 81445 79466 81447
rect 81090 81499 81146 81501
rect 81090 81447 81092 81499
rect 81092 81447 81144 81499
rect 81144 81447 81146 81499
rect 81090 81445 81146 81447
rect 82770 81499 82826 81501
rect 82770 81447 82772 81499
rect 82772 81447 82824 81499
rect 82824 81447 82826 81499
rect 82770 81445 82826 81447
rect 84450 81499 84506 81501
rect 84450 81447 84452 81499
rect 84452 81447 84504 81499
rect 84504 81447 84506 81499
rect 84450 81445 84506 81447
rect 86130 81499 86186 81501
rect 86130 81447 86132 81499
rect 86132 81447 86184 81499
rect 86184 81447 86186 81499
rect 86130 81445 86186 81447
rect 87810 81499 87866 81501
rect 87810 81447 87812 81499
rect 87812 81447 87864 81499
rect 87864 81447 87866 81499
rect 87810 81445 87866 81447
rect 89490 81499 89546 81501
rect 89490 81447 89492 81499
rect 89492 81447 89544 81499
rect 89544 81447 89546 81499
rect 89490 81445 89546 81447
rect 91170 81499 91226 81501
rect 91170 81447 91172 81499
rect 91172 81447 91224 81499
rect 91224 81447 91226 81499
rect 91170 81445 91226 81447
rect 92850 81499 92906 81501
rect 92850 81447 92852 81499
rect 92852 81447 92904 81499
rect 92904 81447 92906 81499
rect 92850 81445 92906 81447
rect 94530 81499 94586 81501
rect 94530 81447 94532 81499
rect 94532 81447 94584 81499
rect 94584 81447 94586 81499
rect 94530 81445 94586 81447
rect 96210 81499 96266 81501
rect 96210 81447 96212 81499
rect 96212 81447 96264 81499
rect 96264 81447 96266 81499
rect 96210 81445 96266 81447
rect 97890 81499 97946 81501
rect 97890 81447 97892 81499
rect 97892 81447 97944 81499
rect 97944 81447 97946 81499
rect 97890 81445 97946 81447
rect 99570 81499 99626 81501
rect 99570 81447 99572 81499
rect 99572 81447 99624 81499
rect 99624 81447 99626 81499
rect 99570 81445 99626 81447
rect 101250 81499 101306 81501
rect 101250 81447 101252 81499
rect 101252 81447 101304 81499
rect 101304 81447 101306 81499
rect 101250 81445 101306 81447
rect 102930 81499 102986 81501
rect 102930 81447 102932 81499
rect 102932 81447 102984 81499
rect 102984 81447 102986 81499
rect 102930 81445 102986 81447
rect 104610 81499 104666 81501
rect 104610 81447 104612 81499
rect 104612 81447 104664 81499
rect 104664 81447 104666 81499
rect 104610 81445 104666 81447
rect 106290 81499 106346 81501
rect 106290 81447 106292 81499
rect 106292 81447 106344 81499
rect 106344 81447 106346 81499
rect 106290 81445 106346 81447
rect 107970 81499 108026 81501
rect 107970 81447 107972 81499
rect 107972 81447 108024 81499
rect 108024 81447 108026 81499
rect 107970 81445 108026 81447
rect 109650 81499 109706 81501
rect 109650 81447 109652 81499
rect 109652 81447 109704 81499
rect 109704 81447 109706 81499
rect 109650 81445 109706 81447
rect 111330 81499 111386 81501
rect 111330 81447 111332 81499
rect 111332 81447 111384 81499
rect 111384 81447 111386 81499
rect 111330 81445 111386 81447
rect 113010 81499 113066 81501
rect 113010 81447 113012 81499
rect 113012 81447 113064 81499
rect 113064 81447 113066 81499
rect 113010 81445 113066 81447
rect 114690 81499 114746 81501
rect 114690 81447 114692 81499
rect 114692 81447 114744 81499
rect 114744 81447 114746 81499
rect 114690 81445 114746 81447
rect 116370 81499 116426 81501
rect 116370 81447 116372 81499
rect 116372 81447 116424 81499
rect 116424 81447 116426 81499
rect 116370 81445 116426 81447
rect 118050 81499 118106 81501
rect 118050 81447 118052 81499
rect 118052 81447 118104 81499
rect 118104 81447 118106 81499
rect 118050 81445 118106 81447
rect 119730 81499 119786 81501
rect 119730 81447 119732 81499
rect 119732 81447 119784 81499
rect 119784 81447 119786 81499
rect 119730 81445 119786 81447
rect 121410 81499 121466 81501
rect 121410 81447 121412 81499
rect 121412 81447 121464 81499
rect 121464 81447 121466 81499
rect 121410 81445 121466 81447
rect 123090 81499 123146 81501
rect 123090 81447 123092 81499
rect 123092 81447 123144 81499
rect 123144 81447 123146 81499
rect 123090 81445 123146 81447
rect 124770 81499 124826 81501
rect 124770 81447 124772 81499
rect 124772 81447 124824 81499
rect 124824 81447 124826 81499
rect 124770 81445 124826 81447
rect 126450 81499 126506 81501
rect 126450 81447 126452 81499
rect 126452 81447 126504 81499
rect 126504 81447 126506 81499
rect 126450 81445 126506 81447
rect 128130 81499 128186 81501
rect 128130 81447 128132 81499
rect 128132 81447 128184 81499
rect 128184 81447 128186 81499
rect 128130 81445 128186 81447
rect 129810 81499 129866 81501
rect 129810 81447 129812 81499
rect 129812 81447 129864 81499
rect 129864 81447 129866 81499
rect 129810 81445 129866 81447
rect 131490 81499 131546 81501
rect 131490 81447 131492 81499
rect 131492 81447 131544 81499
rect 131544 81447 131546 81499
rect 131490 81445 131546 81447
rect 133170 81499 133226 81501
rect 133170 81447 133172 81499
rect 133172 81447 133224 81499
rect 133224 81447 133226 81499
rect 133170 81445 133226 81447
rect 1794 81046 1850 81048
rect 1794 80994 1796 81046
rect 1796 80994 1848 81046
rect 1848 80994 1850 81046
rect 1794 80992 1850 80994
rect 134844 81046 134900 81048
rect 134844 80994 134846 81046
rect 134846 80994 134898 81046
rect 134898 80994 134900 81046
rect 134844 80992 134900 80994
rect 122188 80465 122244 80521
rect 118598 80209 118654 80265
rect 119766 80209 119822 80265
rect 1794 79366 1850 79368
rect 1794 79314 1796 79366
rect 1796 79314 1848 79366
rect 1848 79314 1850 79366
rect 1794 79312 1850 79314
rect 1794 77686 1850 77688
rect 1794 77634 1796 77686
rect 1796 77634 1848 77686
rect 1848 77634 1850 77686
rect 1794 77632 1850 77634
rect 134844 79366 134900 79368
rect 134844 79314 134846 79366
rect 134846 79314 134898 79366
rect 134898 79314 134900 79366
rect 134844 79312 134900 79314
rect 133884 79212 133940 79268
rect 130747 79107 130803 79163
rect 28618 77045 28674 77047
rect 28618 76993 28620 77045
rect 28620 76993 28672 77045
rect 28672 76993 28674 77045
rect 28618 76991 28674 76993
rect 31114 77045 31170 77047
rect 31114 76993 31116 77045
rect 31116 76993 31168 77045
rect 31168 76993 31170 77045
rect 31114 76991 31170 76993
rect 33610 77045 33666 77047
rect 33610 76993 33612 77045
rect 33612 76993 33664 77045
rect 33664 76993 33666 77045
rect 33610 76991 33666 76993
rect 36106 77045 36162 77047
rect 36106 76993 36108 77045
rect 36108 76993 36160 77045
rect 36160 76993 36162 77045
rect 36106 76991 36162 76993
rect 38602 77045 38658 77047
rect 38602 76993 38604 77045
rect 38604 76993 38656 77045
rect 38656 76993 38658 77045
rect 38602 76991 38658 76993
rect 41098 77045 41154 77047
rect 41098 76993 41100 77045
rect 41100 76993 41152 77045
rect 41152 76993 41154 77045
rect 41098 76991 41154 76993
rect 43594 77045 43650 77047
rect 43594 76993 43596 77045
rect 43596 76993 43648 77045
rect 43648 76993 43650 77045
rect 43594 76991 43650 76993
rect 46090 77045 46146 77047
rect 46090 76993 46092 77045
rect 46092 76993 46144 77045
rect 46144 76993 46146 77045
rect 46090 76991 46146 76993
rect 48586 77045 48642 77047
rect 48586 76993 48588 77045
rect 48588 76993 48640 77045
rect 48640 76993 48642 77045
rect 48586 76991 48642 76993
rect 51082 77045 51138 77047
rect 51082 76993 51084 77045
rect 51084 76993 51136 77045
rect 51136 76993 51138 77045
rect 51082 76991 51138 76993
rect 53578 77045 53634 77047
rect 53578 76993 53580 77045
rect 53580 76993 53632 77045
rect 53632 76993 53634 77045
rect 53578 76991 53634 76993
rect 56074 77045 56130 77047
rect 56074 76993 56076 77045
rect 56076 76993 56128 77045
rect 56128 76993 56130 77045
rect 56074 76991 56130 76993
rect 58570 77045 58626 77047
rect 58570 76993 58572 77045
rect 58572 76993 58624 77045
rect 58624 76993 58626 77045
rect 58570 76991 58626 76993
rect 61066 77045 61122 77047
rect 61066 76993 61068 77045
rect 61068 76993 61120 77045
rect 61120 76993 61122 77045
rect 61066 76991 61122 76993
rect 63562 77045 63618 77047
rect 63562 76993 63564 77045
rect 63564 76993 63616 77045
rect 63616 76993 63618 77045
rect 63562 76991 63618 76993
rect 66058 77045 66114 77047
rect 66058 76993 66060 77045
rect 66060 76993 66112 77045
rect 66112 76993 66114 77045
rect 66058 76991 66114 76993
rect 68554 77045 68610 77047
rect 68554 76993 68556 77045
rect 68556 76993 68608 77045
rect 68608 76993 68610 77045
rect 68554 76991 68610 76993
rect 71050 77045 71106 77047
rect 71050 76993 71052 77045
rect 71052 76993 71104 77045
rect 71104 76993 71106 77045
rect 71050 76991 71106 76993
rect 73546 77045 73602 77047
rect 73546 76993 73548 77045
rect 73548 76993 73600 77045
rect 73600 76993 73602 77045
rect 73546 76991 73602 76993
rect 76042 77045 76098 77047
rect 76042 76993 76044 77045
rect 76044 76993 76096 77045
rect 76096 76993 76098 77045
rect 76042 76991 76098 76993
rect 78538 77045 78594 77047
rect 78538 76993 78540 77045
rect 78540 76993 78592 77045
rect 78592 76993 78594 77045
rect 78538 76991 78594 76993
rect 81034 77045 81090 77047
rect 81034 76993 81036 77045
rect 81036 76993 81088 77045
rect 81088 76993 81090 77045
rect 81034 76991 81090 76993
rect 83530 77045 83586 77047
rect 83530 76993 83532 77045
rect 83532 76993 83584 77045
rect 83584 76993 83586 77045
rect 83530 76991 83586 76993
rect 86026 77045 86082 77047
rect 86026 76993 86028 77045
rect 86028 76993 86080 77045
rect 86080 76993 86082 77045
rect 86026 76991 86082 76993
rect 88522 77045 88578 77047
rect 88522 76993 88524 77045
rect 88524 76993 88576 77045
rect 88576 76993 88578 77045
rect 88522 76991 88578 76993
rect 91018 77045 91074 77047
rect 91018 76993 91020 77045
rect 91020 76993 91072 77045
rect 91072 76993 91074 77045
rect 91018 76991 91074 76993
rect 93514 77045 93570 77047
rect 93514 76993 93516 77045
rect 93516 76993 93568 77045
rect 93568 76993 93570 77045
rect 93514 76991 93570 76993
rect 96010 77045 96066 77047
rect 96010 76993 96012 77045
rect 96012 76993 96064 77045
rect 96064 76993 96066 77045
rect 96010 76991 96066 76993
rect 98506 77045 98562 77047
rect 98506 76993 98508 77045
rect 98508 76993 98560 77045
rect 98560 76993 98562 77045
rect 98506 76991 98562 76993
rect 101002 77045 101058 77047
rect 101002 76993 101004 77045
rect 101004 76993 101056 77045
rect 101056 76993 101058 77045
rect 101002 76991 101058 76993
rect 103498 77045 103554 77047
rect 103498 76993 103500 77045
rect 103500 76993 103552 77045
rect 103552 76993 103554 77045
rect 103498 76991 103554 76993
rect 105994 77045 106050 77047
rect 105994 76993 105996 77045
rect 105996 76993 106048 77045
rect 106048 76993 106050 77045
rect 105994 76991 106050 76993
rect 1794 76006 1850 76008
rect 1794 75954 1796 76006
rect 1796 75954 1848 76006
rect 1848 75954 1850 76006
rect 1794 75952 1850 75954
rect 110061 74827 110117 74883
rect 1794 74326 1850 74328
rect 1794 74274 1796 74326
rect 1796 74274 1848 74326
rect 1848 74274 1850 74326
rect 1794 74272 1850 74274
rect 1794 72646 1850 72648
rect 1794 72594 1796 72646
rect 1796 72594 1848 72646
rect 1848 72594 1850 72646
rect 1794 72592 1850 72594
rect 110185 73413 110241 73469
rect 114046 71999 114102 72055
rect 1794 70966 1850 70968
rect 1794 70914 1796 70966
rect 1796 70914 1848 70966
rect 1848 70914 1850 70966
rect 1794 70912 1850 70914
rect 1794 69286 1850 69288
rect 1794 69234 1796 69286
rect 1796 69234 1848 69286
rect 1848 69234 1850 69286
rect 1794 69232 1850 69234
rect 1794 67606 1850 67608
rect 1794 67554 1796 67606
rect 1796 67554 1848 67606
rect 1848 67554 1850 67606
rect 1794 67552 1850 67554
rect 1794 65926 1850 65928
rect 1794 65874 1796 65926
rect 1796 65874 1848 65926
rect 1848 65874 1850 65926
rect 1794 65872 1850 65874
rect 1794 64246 1850 64248
rect 1794 64194 1796 64246
rect 1796 64194 1848 64246
rect 1848 64194 1850 64246
rect 1794 64192 1850 64194
rect 1794 62566 1850 62568
rect 1794 62514 1796 62566
rect 1796 62514 1848 62566
rect 1848 62514 1850 62566
rect 1794 62512 1850 62514
rect 1794 60886 1850 60888
rect 1794 60834 1796 60886
rect 1796 60834 1848 60886
rect 1848 60834 1850 60886
rect 1794 60832 1850 60834
rect 1794 59206 1850 59208
rect 1794 59154 1796 59206
rect 1796 59154 1848 59206
rect 1848 59154 1850 59206
rect 1794 59152 1850 59154
rect 1794 57526 1850 57528
rect 1794 57474 1796 57526
rect 1796 57474 1848 57526
rect 1848 57474 1850 57526
rect 1794 57472 1850 57474
rect 1794 55846 1850 55848
rect 1794 55794 1796 55846
rect 1796 55794 1848 55846
rect 1848 55794 1850 55846
rect 1794 55792 1850 55794
rect 1794 54166 1850 54168
rect 1794 54114 1796 54166
rect 1796 54114 1848 54166
rect 1848 54114 1850 54166
rect 1794 54112 1850 54114
rect 1794 52486 1850 52488
rect 1794 52434 1796 52486
rect 1796 52434 1848 52486
rect 1848 52434 1850 52486
rect 1794 52432 1850 52434
rect 1794 50806 1850 50808
rect 1794 50754 1796 50806
rect 1796 50754 1848 50806
rect 1848 50754 1850 50806
rect 1794 50752 1850 50754
rect 1794 49126 1850 49128
rect 1794 49074 1796 49126
rect 1796 49074 1848 49126
rect 1848 49074 1850 49126
rect 1794 49072 1850 49074
rect 1794 47446 1850 47448
rect 1794 47394 1796 47446
rect 1796 47394 1848 47446
rect 1848 47394 1850 47446
rect 1794 47392 1850 47394
rect 1794 45766 1850 45768
rect 1794 45714 1796 45766
rect 1796 45714 1848 45766
rect 1848 45714 1850 45766
rect 1794 45712 1850 45714
rect 1794 44086 1850 44088
rect 1794 44034 1796 44086
rect 1796 44034 1848 44086
rect 1848 44034 1850 44086
rect 1794 44032 1850 44034
rect 1794 42406 1850 42408
rect 1794 42354 1796 42406
rect 1796 42354 1848 42406
rect 1848 42354 1850 42406
rect 1794 42352 1850 42354
rect 1794 40726 1850 40728
rect 1794 40674 1796 40726
rect 1796 40674 1848 40726
rect 1848 40674 1850 40726
rect 1794 40672 1850 40674
rect 1794 39046 1850 39048
rect 1794 38994 1796 39046
rect 1796 38994 1848 39046
rect 1848 38994 1850 39046
rect 1794 38992 1850 38994
rect 1794 37366 1850 37368
rect 1794 37314 1796 37366
rect 1796 37314 1848 37366
rect 1848 37314 1850 37366
rect 1794 37312 1850 37314
rect 14613 36837 14669 36893
rect 15347 36891 15403 36893
rect 15347 36839 15349 36891
rect 15349 36839 15401 36891
rect 15401 36839 15403 36891
rect 15347 36837 15403 36839
rect 13668 36766 13724 36822
rect 1794 35686 1850 35688
rect 1794 35634 1796 35686
rect 1796 35634 1848 35686
rect 1848 35634 1850 35686
rect 1794 35632 1850 35634
rect 13668 35638 13724 35694
rect 14613 35567 14669 35623
rect 15267 35621 15323 35623
rect 15267 35569 15269 35621
rect 15269 35569 15321 35621
rect 15321 35569 15323 35621
rect 15267 35567 15323 35569
rect 1794 34006 1850 34008
rect 1794 33954 1796 34006
rect 1796 33954 1848 34006
rect 1848 33954 1850 34006
rect 1794 33952 1850 33954
rect 14613 34009 14669 34065
rect 15187 34063 15243 34065
rect 15187 34011 15189 34063
rect 15189 34011 15241 34063
rect 15241 34011 15243 34063
rect 15187 34009 15243 34011
rect 13668 33938 13724 33994
rect 13668 32810 13724 32866
rect 14613 32739 14669 32795
rect 15107 32793 15163 32795
rect 15107 32741 15109 32793
rect 15109 32741 15161 32793
rect 15161 32741 15163 32793
rect 15107 32739 15163 32741
rect 1794 32326 1850 32328
rect 1794 32274 1796 32326
rect 1796 32274 1848 32326
rect 1848 32274 1850 32326
rect 1794 32272 1850 32274
rect 14613 31181 14669 31237
rect 15027 31235 15083 31237
rect 15027 31183 15029 31235
rect 15029 31183 15081 31235
rect 15081 31183 15083 31235
rect 15027 31181 15083 31183
rect 13668 31110 13724 31166
rect 1794 30646 1850 30648
rect 1794 30594 1796 30646
rect 1796 30594 1848 30646
rect 1848 30594 1850 30646
rect 1794 30592 1850 30594
rect 13668 29982 13724 30038
rect 14613 29911 14669 29967
rect 14947 29965 15003 29967
rect 14947 29913 14949 29965
rect 14949 29913 15001 29965
rect 15001 29913 15003 29965
rect 14947 29911 15003 29913
rect 1794 28966 1850 28968
rect 1794 28914 1796 28966
rect 1796 28914 1848 28966
rect 1848 28914 1850 28966
rect 1794 28912 1850 28914
rect 14613 28353 14669 28409
rect 14867 28407 14923 28409
rect 14867 28355 14869 28407
rect 14869 28355 14921 28407
rect 14921 28355 14923 28407
rect 14867 28353 14923 28355
rect 13668 28282 13724 28338
rect 14750 28026 14806 28082
rect 1794 27286 1850 27288
rect 1794 27234 1796 27286
rect 1796 27234 1848 27286
rect 1848 27234 1850 27286
rect 1794 27232 1850 27234
rect 1794 25606 1850 25608
rect 1794 25554 1796 25606
rect 1796 25554 1848 25606
rect 1848 25554 1850 25606
rect 1794 25552 1850 25554
rect 2541 25305 2597 25361
rect 1794 23926 1850 23928
rect 1794 23874 1796 23926
rect 1796 23874 1848 23926
rect 1848 23874 1850 23926
rect 1794 23872 1850 23874
rect 1794 22246 1850 22248
rect 1794 22194 1796 22246
rect 1796 22194 1848 22246
rect 1848 22194 1850 22246
rect 1794 22192 1850 22194
rect 1794 20566 1850 20568
rect 1794 20514 1796 20566
rect 1796 20514 1848 20566
rect 1848 20514 1850 20566
rect 1794 20512 1850 20514
rect 1794 18886 1850 18888
rect 1794 18834 1796 18886
rect 1796 18834 1848 18886
rect 1848 18834 1850 18886
rect 1794 18832 1850 18834
rect 14666 18197 14722 18253
rect 1794 17206 1850 17208
rect 1794 17154 1796 17206
rect 1796 17154 1848 17206
rect 1848 17154 1850 17206
rect 1794 17152 1850 17154
rect 1794 15526 1850 15528
rect 1794 15474 1796 15526
rect 1796 15474 1848 15526
rect 1848 15474 1850 15526
rect 1794 15472 1850 15474
rect 14666 15369 14722 15425
rect 14666 13955 14722 14011
rect 1794 13846 1850 13848
rect 1794 13794 1796 13846
rect 1796 13794 1848 13846
rect 1848 13794 1850 13846
rect 1794 13792 1850 13794
rect 14666 12541 14722 12597
rect 1794 12166 1850 12168
rect 1794 12114 1796 12166
rect 1796 12114 1848 12166
rect 1848 12114 1850 12166
rect 1794 12112 1850 12114
rect 1794 10486 1850 10488
rect 1794 10434 1796 10486
rect 1796 10434 1848 10486
rect 1848 10434 1850 10486
rect 1794 10432 1850 10434
rect 2754 9856 2810 9912
rect 1794 8806 1850 8808
rect 1794 8754 1796 8806
rect 1796 8754 1848 8806
rect 1848 8754 1850 8806
rect 1794 8752 1850 8754
rect 134844 77686 134900 77688
rect 134844 77634 134846 77686
rect 134846 77634 134898 77686
rect 134898 77634 134900 77686
rect 134844 77632 134900 77634
rect 134844 76006 134900 76008
rect 134844 75954 134846 76006
rect 134846 75954 134898 76006
rect 134898 75954 134900 76006
rect 134844 75952 134900 75954
rect 122272 74827 122328 74883
rect 134844 74326 134900 74328
rect 134844 74274 134846 74326
rect 134846 74274 134898 74326
rect 134898 74274 134900 74326
rect 134844 74272 134900 74274
rect 122272 73413 122328 73469
rect 134844 72646 134900 72648
rect 134844 72594 134846 72646
rect 134846 72594 134898 72646
rect 134898 72594 134900 72646
rect 134844 72592 134900 72594
rect 122272 71999 122328 72055
rect 134844 70966 134900 70968
rect 134844 70914 134846 70966
rect 134846 70914 134898 70966
rect 134898 70914 134900 70966
rect 134844 70912 134900 70914
rect 134844 69286 134900 69288
rect 134844 69234 134846 69286
rect 134846 69234 134898 69286
rect 134898 69234 134900 69286
rect 134844 69232 134900 69234
rect 134844 67606 134900 67608
rect 134844 67554 134846 67606
rect 134846 67554 134898 67606
rect 134898 67554 134900 67606
rect 134844 67552 134900 67554
rect 134844 65926 134900 65928
rect 134844 65874 134846 65926
rect 134846 65874 134898 65926
rect 134898 65874 134900 65926
rect 134844 65872 134900 65874
rect 134844 64246 134900 64248
rect 134844 64194 134846 64246
rect 134846 64194 134898 64246
rect 134898 64194 134900 64246
rect 134844 64192 134900 64194
rect 134844 62566 134900 62568
rect 134844 62514 134846 62566
rect 134846 62514 134898 62566
rect 134898 62514 134900 62566
rect 134844 62512 134900 62514
rect 134097 62063 134153 62119
rect 134844 60886 134900 60888
rect 134844 60834 134846 60886
rect 134846 60834 134898 60886
rect 134898 60834 134900 60886
rect 134844 60832 134900 60834
rect 134844 59206 134900 59208
rect 134844 59154 134846 59206
rect 134846 59154 134898 59206
rect 134898 59154 134900 59206
rect 134844 59152 134900 59154
rect 134844 57526 134900 57528
rect 134844 57474 134846 57526
rect 134846 57474 134898 57526
rect 134898 57474 134900 57526
rect 134844 57472 134900 57474
rect 134844 55846 134900 55848
rect 134844 55794 134846 55846
rect 134846 55794 134898 55846
rect 134898 55794 134900 55846
rect 134844 55792 134900 55794
rect 134844 54166 134900 54168
rect 134844 54114 134846 54166
rect 134846 54114 134898 54166
rect 134898 54114 134900 54166
rect 134844 54112 134900 54114
rect 134844 52486 134900 52488
rect 134844 52434 134846 52486
rect 134846 52434 134898 52486
rect 134898 52434 134900 52486
rect 134844 52432 134900 52434
rect 134844 50806 134900 50808
rect 134844 50754 134846 50806
rect 134846 50754 134898 50806
rect 134898 50754 134900 50806
rect 134844 50752 134900 50754
rect 134844 49126 134900 49128
rect 134844 49074 134846 49126
rect 134846 49074 134898 49126
rect 134898 49074 134900 49126
rect 134844 49072 134900 49074
rect 134844 47446 134900 47448
rect 134844 47394 134846 47446
rect 134846 47394 134898 47446
rect 134898 47394 134900 47446
rect 134844 47392 134900 47394
rect 134844 45766 134900 45768
rect 134844 45714 134846 45766
rect 134846 45714 134898 45766
rect 134898 45714 134900 45766
rect 134844 45712 134900 45714
rect 134844 44086 134900 44088
rect 134844 44034 134846 44086
rect 134846 44034 134898 44086
rect 134898 44034 134900 44086
rect 134844 44032 134900 44034
rect 134844 42406 134900 42408
rect 134844 42354 134846 42406
rect 134846 42354 134898 42406
rect 134898 42354 134900 42406
rect 134844 42352 134900 42354
rect 134844 40726 134900 40728
rect 134844 40674 134846 40726
rect 134846 40674 134898 40726
rect 134898 40674 134900 40726
rect 134844 40672 134900 40674
rect 134844 39046 134900 39048
rect 134844 38994 134846 39046
rect 134846 38994 134898 39046
rect 134898 38994 134900 39046
rect 134844 38992 134900 38994
rect 134844 37366 134900 37368
rect 134844 37314 134846 37366
rect 134846 37314 134898 37366
rect 134898 37314 134900 37366
rect 134844 37312 134900 37314
rect 134844 35686 134900 35688
rect 134844 35634 134846 35686
rect 134846 35634 134898 35686
rect 134898 35634 134900 35686
rect 134844 35632 134900 35634
rect 134844 34006 134900 34008
rect 134844 33954 134846 34006
rect 134846 33954 134898 34006
rect 134898 33954 134900 34006
rect 134844 33952 134900 33954
rect 134844 32326 134900 32328
rect 134844 32274 134846 32326
rect 134846 32274 134898 32326
rect 134898 32274 134900 32326
rect 134844 32272 134900 32274
rect 134844 30646 134900 30648
rect 134844 30594 134846 30646
rect 134846 30594 134898 30646
rect 134898 30594 134900 30646
rect 134844 30592 134900 30594
rect 134844 28966 134900 28968
rect 134844 28914 134846 28966
rect 134846 28914 134898 28966
rect 134898 28914 134900 28966
rect 134844 28912 134900 28914
rect 134844 27286 134900 27288
rect 134844 27234 134846 27286
rect 134846 27234 134898 27286
rect 134898 27234 134900 27286
rect 134844 27232 134900 27234
rect 134844 25606 134900 25608
rect 134844 25554 134846 25606
rect 134846 25554 134898 25606
rect 134898 25554 134900 25606
rect 134844 25552 134900 25554
rect 134844 23926 134900 23928
rect 134844 23874 134846 23926
rect 134846 23874 134898 23926
rect 134898 23874 134900 23926
rect 134844 23872 134900 23874
rect 134844 22246 134900 22248
rect 134844 22194 134846 22246
rect 134846 22194 134898 22246
rect 134898 22194 134900 22246
rect 134844 22192 134900 22194
rect 134844 20566 134900 20568
rect 134844 20514 134846 20566
rect 134846 20514 134898 20566
rect 134898 20514 134900 20566
rect 134844 20512 134900 20514
rect 122188 19510 122244 19566
rect 123270 19254 123326 19310
rect 121987 19237 122043 19239
rect 121987 19185 121989 19237
rect 121989 19185 122041 19237
rect 122041 19185 122043 19237
rect 121987 19183 122043 19185
rect 122325 19183 122381 19239
rect 22808 18197 22864 18253
rect 134844 18886 134900 18888
rect 134844 18834 134846 18886
rect 134846 18834 134898 18886
rect 134898 18834 134900 18886
rect 134844 18832 134900 18834
rect 121907 17679 121963 17681
rect 121907 17627 121909 17679
rect 121909 17627 121961 17679
rect 121961 17627 121963 17679
rect 121907 17625 121963 17627
rect 122325 17625 122381 17681
rect 123270 17554 123326 17610
rect 134844 17206 134900 17208
rect 134844 17154 134846 17206
rect 134846 17154 134898 17206
rect 134898 17154 134900 17206
rect 134844 17152 134900 17154
rect 123270 16426 123326 16482
rect 121827 16409 121883 16411
rect 121827 16357 121829 16409
rect 121829 16357 121881 16409
rect 121881 16357 121883 16409
rect 121827 16355 121883 16357
rect 122325 16355 122381 16411
rect 134844 15526 134900 15528
rect 134844 15474 134846 15526
rect 134846 15474 134898 15526
rect 134898 15474 134900 15526
rect 134844 15472 134900 15474
rect 26511 15369 26567 15425
rect 121747 14851 121803 14853
rect 121747 14799 121749 14851
rect 121749 14799 121801 14851
rect 121801 14799 121803 14851
rect 121747 14797 121803 14799
rect 122325 14797 122381 14853
rect 123270 14726 123326 14782
rect 26759 13955 26815 14011
rect 26635 12541 26691 12597
rect 134844 13846 134900 13848
rect 134844 13794 134846 13846
rect 134846 13794 134898 13846
rect 134898 13794 134900 13846
rect 134844 13792 134900 13794
rect 123270 13598 123326 13654
rect 121667 13581 121723 13583
rect 121667 13529 121669 13581
rect 121669 13529 121721 13581
rect 121721 13529 121723 13581
rect 121667 13527 121723 13529
rect 122325 13527 122381 13583
rect 28618 13259 28674 13261
rect 28618 13207 28620 13259
rect 28620 13207 28672 13259
rect 28672 13207 28674 13259
rect 28618 13205 28674 13207
rect 31114 13259 31170 13261
rect 31114 13207 31116 13259
rect 31116 13207 31168 13259
rect 31168 13207 31170 13259
rect 31114 13205 31170 13207
rect 33610 13259 33666 13261
rect 33610 13207 33612 13259
rect 33612 13207 33664 13259
rect 33664 13207 33666 13259
rect 33610 13205 33666 13207
rect 36106 13259 36162 13261
rect 36106 13207 36108 13259
rect 36108 13207 36160 13259
rect 36160 13207 36162 13259
rect 36106 13205 36162 13207
rect 38602 13259 38658 13261
rect 38602 13207 38604 13259
rect 38604 13207 38656 13259
rect 38656 13207 38658 13259
rect 38602 13205 38658 13207
rect 41098 13259 41154 13261
rect 41098 13207 41100 13259
rect 41100 13207 41152 13259
rect 41152 13207 41154 13259
rect 41098 13205 41154 13207
rect 43594 13259 43650 13261
rect 43594 13207 43596 13259
rect 43596 13207 43648 13259
rect 43648 13207 43650 13259
rect 43594 13205 43650 13207
rect 46090 13259 46146 13261
rect 46090 13207 46092 13259
rect 46092 13207 46144 13259
rect 46144 13207 46146 13259
rect 46090 13205 46146 13207
rect 48586 13259 48642 13261
rect 48586 13207 48588 13259
rect 48588 13207 48640 13259
rect 48640 13207 48642 13259
rect 48586 13205 48642 13207
rect 51082 13259 51138 13261
rect 51082 13207 51084 13259
rect 51084 13207 51136 13259
rect 51136 13207 51138 13259
rect 51082 13205 51138 13207
rect 53578 13259 53634 13261
rect 53578 13207 53580 13259
rect 53580 13207 53632 13259
rect 53632 13207 53634 13259
rect 53578 13205 53634 13207
rect 56074 13259 56130 13261
rect 56074 13207 56076 13259
rect 56076 13207 56128 13259
rect 56128 13207 56130 13259
rect 56074 13205 56130 13207
rect 58570 13259 58626 13261
rect 58570 13207 58572 13259
rect 58572 13207 58624 13259
rect 58624 13207 58626 13259
rect 58570 13205 58626 13207
rect 61066 13259 61122 13261
rect 61066 13207 61068 13259
rect 61068 13207 61120 13259
rect 61120 13207 61122 13259
rect 61066 13205 61122 13207
rect 63562 13259 63618 13261
rect 63562 13207 63564 13259
rect 63564 13207 63616 13259
rect 63616 13207 63618 13259
rect 63562 13205 63618 13207
rect 66058 13259 66114 13261
rect 66058 13207 66060 13259
rect 66060 13207 66112 13259
rect 66112 13207 66114 13259
rect 66058 13205 66114 13207
rect 68554 13259 68610 13261
rect 68554 13207 68556 13259
rect 68556 13207 68608 13259
rect 68608 13207 68610 13259
rect 68554 13205 68610 13207
rect 71050 13259 71106 13261
rect 71050 13207 71052 13259
rect 71052 13207 71104 13259
rect 71104 13207 71106 13259
rect 71050 13205 71106 13207
rect 73546 13259 73602 13261
rect 73546 13207 73548 13259
rect 73548 13207 73600 13259
rect 73600 13207 73602 13259
rect 73546 13205 73602 13207
rect 76042 13259 76098 13261
rect 76042 13207 76044 13259
rect 76044 13207 76096 13259
rect 76096 13207 76098 13259
rect 76042 13205 76098 13207
rect 78538 13259 78594 13261
rect 78538 13207 78540 13259
rect 78540 13207 78592 13259
rect 78592 13207 78594 13259
rect 78538 13205 78594 13207
rect 81034 13259 81090 13261
rect 81034 13207 81036 13259
rect 81036 13207 81088 13259
rect 81088 13207 81090 13259
rect 81034 13205 81090 13207
rect 83530 13259 83586 13261
rect 83530 13207 83532 13259
rect 83532 13207 83584 13259
rect 83584 13207 83586 13259
rect 83530 13205 83586 13207
rect 86026 13259 86082 13261
rect 86026 13207 86028 13259
rect 86028 13207 86080 13259
rect 86080 13207 86082 13259
rect 86026 13205 86082 13207
rect 88522 13259 88578 13261
rect 88522 13207 88524 13259
rect 88524 13207 88576 13259
rect 88576 13207 88578 13259
rect 88522 13205 88578 13207
rect 91018 13259 91074 13261
rect 91018 13207 91020 13259
rect 91020 13207 91072 13259
rect 91072 13207 91074 13259
rect 91018 13205 91074 13207
rect 93514 13259 93570 13261
rect 93514 13207 93516 13259
rect 93516 13207 93568 13259
rect 93568 13207 93570 13259
rect 93514 13205 93570 13207
rect 96010 13259 96066 13261
rect 96010 13207 96012 13259
rect 96012 13207 96064 13259
rect 96064 13207 96066 13259
rect 96010 13205 96066 13207
rect 98506 13259 98562 13261
rect 98506 13207 98508 13259
rect 98508 13207 98560 13259
rect 98560 13207 98562 13259
rect 98506 13205 98562 13207
rect 101002 13259 101058 13261
rect 101002 13207 101004 13259
rect 101004 13207 101056 13259
rect 101056 13207 101058 13259
rect 101002 13205 101058 13207
rect 103498 13259 103554 13261
rect 103498 13207 103500 13259
rect 103500 13207 103552 13259
rect 103552 13207 103554 13259
rect 103498 13205 103554 13207
rect 105994 13259 106050 13261
rect 105994 13207 105996 13259
rect 105996 13207 106048 13259
rect 106048 13207 106050 13259
rect 105994 13205 106050 13207
rect 134844 12166 134900 12168
rect 134844 12114 134846 12166
rect 134846 12114 134898 12166
rect 134898 12114 134900 12166
rect 134844 12112 134900 12114
rect 121587 12023 121643 12025
rect 121587 11971 121589 12023
rect 121589 11971 121641 12023
rect 121641 11971 121643 12023
rect 121587 11969 121643 11971
rect 122325 11969 122381 12025
rect 123270 11898 123326 11954
rect 123270 10770 123326 10826
rect 121507 10753 121563 10755
rect 121507 10701 121509 10753
rect 121509 10701 121561 10753
rect 121561 10701 121563 10753
rect 121507 10699 121563 10701
rect 122325 10699 122381 10755
rect 134844 10486 134900 10488
rect 134844 10434 134846 10486
rect 134846 10434 134898 10486
rect 134898 10434 134900 10486
rect 134844 10432 134900 10434
rect 5975 8261 6031 8317
rect 2754 8156 2810 8212
rect 1794 7126 1850 7128
rect 1794 7074 1796 7126
rect 1796 7074 1848 7126
rect 1848 7074 1850 7126
rect 1794 7072 1850 7074
rect 1794 5446 1850 5448
rect 1794 5394 1796 5446
rect 1796 5394 1848 5446
rect 1848 5394 1850 5446
rect 1794 5392 1850 5394
rect 1794 3766 1850 3768
rect 1794 3714 1796 3766
rect 1796 3714 1848 3766
rect 1848 3714 1850 3766
rect 1794 3712 1850 3714
rect 134844 8806 134900 8808
rect 134844 8754 134846 8806
rect 134846 8754 134898 8806
rect 134898 8754 134900 8806
rect 134844 8752 134900 8754
rect 134844 7126 134900 7128
rect 134844 7074 134846 7126
rect 134846 7074 134898 7126
rect 134898 7074 134900 7126
rect 134844 7072 134900 7074
rect 134844 5446 134900 5448
rect 134844 5394 134846 5446
rect 134846 5394 134898 5446
rect 134898 5394 134900 5446
rect 134844 5392 134900 5394
rect 134844 3766 134900 3768
rect 134844 3714 134846 3766
rect 134846 3714 134898 3766
rect 134898 3714 134900 3766
rect 134844 3712 134900 3714
rect 16004 2932 16060 2988
rect 17172 2932 17228 2988
rect 18340 2932 18396 2988
rect 19508 2932 19564 2988
rect 20676 2932 20732 2988
rect 21844 2932 21900 2988
rect 23012 2932 23068 2988
rect 24180 2932 24236 2988
rect 25348 2932 25404 2988
rect 26516 2932 26572 2988
rect 27684 2932 27740 2988
rect 28852 2932 28908 2988
rect 30020 2932 30076 2988
rect 31188 2932 31244 2988
rect 32356 2932 32412 2988
rect 33524 2932 33580 2988
rect 34692 2932 34748 2988
rect 35860 2932 35916 2988
rect 37028 2932 37084 2988
rect 38196 2932 38252 2988
rect 39364 2932 39420 2988
rect 40532 2932 40588 2988
rect 41700 2932 41756 2988
rect 42868 2932 42924 2988
rect 44036 2932 44092 2988
rect 45204 2932 45260 2988
rect 46372 2932 46428 2988
rect 47540 2932 47596 2988
rect 48708 2932 48764 2988
rect 49876 2932 49932 2988
rect 51044 2932 51100 2988
rect 52212 2932 52268 2988
rect 53380 2932 53436 2988
rect 54548 2932 54604 2988
rect 55716 2932 55772 2988
rect 56884 2932 56940 2988
rect 58052 2932 58108 2988
rect 59220 2932 59276 2988
rect 14750 2676 14806 2732
rect 1794 2086 1850 2088
rect 1794 2034 1796 2086
rect 1796 2034 1848 2086
rect 1848 2034 1850 2086
rect 1794 2032 1850 2034
rect 134844 2086 134900 2088
rect 134844 2034 134846 2086
rect 134846 2034 134898 2086
rect 134898 2034 134900 2086
rect 134844 2032 134900 2034
rect 2130 1750 2186 1752
rect 2130 1698 2132 1750
rect 2132 1698 2184 1750
rect 2184 1698 2186 1750
rect 2130 1696 2186 1698
rect 3810 1750 3866 1752
rect 3810 1698 3812 1750
rect 3812 1698 3864 1750
rect 3864 1698 3866 1750
rect 3810 1696 3866 1698
rect 5490 1750 5546 1752
rect 5490 1698 5492 1750
rect 5492 1698 5544 1750
rect 5544 1698 5546 1750
rect 5490 1696 5546 1698
rect 7170 1750 7226 1752
rect 7170 1698 7172 1750
rect 7172 1698 7224 1750
rect 7224 1698 7226 1750
rect 7170 1696 7226 1698
rect 8850 1750 8906 1752
rect 8850 1698 8852 1750
rect 8852 1698 8904 1750
rect 8904 1698 8906 1750
rect 8850 1696 8906 1698
rect 10530 1750 10586 1752
rect 10530 1698 10532 1750
rect 10532 1698 10584 1750
rect 10584 1698 10586 1750
rect 10530 1696 10586 1698
rect 12210 1750 12266 1752
rect 12210 1698 12212 1750
rect 12212 1698 12264 1750
rect 12264 1698 12266 1750
rect 12210 1696 12266 1698
rect 13890 1750 13946 1752
rect 13890 1698 13892 1750
rect 13892 1698 13944 1750
rect 13944 1698 13946 1750
rect 13890 1696 13946 1698
rect 15570 1750 15626 1752
rect 15570 1698 15572 1750
rect 15572 1698 15624 1750
rect 15624 1698 15626 1750
rect 15570 1696 15626 1698
rect 17250 1750 17306 1752
rect 17250 1698 17252 1750
rect 17252 1698 17304 1750
rect 17304 1698 17306 1750
rect 17250 1696 17306 1698
rect 18930 1750 18986 1752
rect 18930 1698 18932 1750
rect 18932 1698 18984 1750
rect 18984 1698 18986 1750
rect 18930 1696 18986 1698
rect 20610 1750 20666 1752
rect 20610 1698 20612 1750
rect 20612 1698 20664 1750
rect 20664 1698 20666 1750
rect 20610 1696 20666 1698
rect 22290 1750 22346 1752
rect 22290 1698 22292 1750
rect 22292 1698 22344 1750
rect 22344 1698 22346 1750
rect 22290 1696 22346 1698
rect 23970 1750 24026 1752
rect 23970 1698 23972 1750
rect 23972 1698 24024 1750
rect 24024 1698 24026 1750
rect 23970 1696 24026 1698
rect 25650 1750 25706 1752
rect 25650 1698 25652 1750
rect 25652 1698 25704 1750
rect 25704 1698 25706 1750
rect 25650 1696 25706 1698
rect 27330 1750 27386 1752
rect 27330 1698 27332 1750
rect 27332 1698 27384 1750
rect 27384 1698 27386 1750
rect 27330 1696 27386 1698
rect 29010 1750 29066 1752
rect 29010 1698 29012 1750
rect 29012 1698 29064 1750
rect 29064 1698 29066 1750
rect 29010 1696 29066 1698
rect 30690 1750 30746 1752
rect 30690 1698 30692 1750
rect 30692 1698 30744 1750
rect 30744 1698 30746 1750
rect 30690 1696 30746 1698
rect 32370 1750 32426 1752
rect 32370 1698 32372 1750
rect 32372 1698 32424 1750
rect 32424 1698 32426 1750
rect 32370 1696 32426 1698
rect 34050 1750 34106 1752
rect 34050 1698 34052 1750
rect 34052 1698 34104 1750
rect 34104 1698 34106 1750
rect 34050 1696 34106 1698
rect 35730 1750 35786 1752
rect 35730 1698 35732 1750
rect 35732 1698 35784 1750
rect 35784 1698 35786 1750
rect 35730 1696 35786 1698
rect 37410 1750 37466 1752
rect 37410 1698 37412 1750
rect 37412 1698 37464 1750
rect 37464 1698 37466 1750
rect 37410 1696 37466 1698
rect 39090 1750 39146 1752
rect 39090 1698 39092 1750
rect 39092 1698 39144 1750
rect 39144 1698 39146 1750
rect 39090 1696 39146 1698
rect 40770 1750 40826 1752
rect 40770 1698 40772 1750
rect 40772 1698 40824 1750
rect 40824 1698 40826 1750
rect 40770 1696 40826 1698
rect 42450 1750 42506 1752
rect 42450 1698 42452 1750
rect 42452 1698 42504 1750
rect 42504 1698 42506 1750
rect 42450 1696 42506 1698
rect 44130 1750 44186 1752
rect 44130 1698 44132 1750
rect 44132 1698 44184 1750
rect 44184 1698 44186 1750
rect 44130 1696 44186 1698
rect 45810 1750 45866 1752
rect 45810 1698 45812 1750
rect 45812 1698 45864 1750
rect 45864 1698 45866 1750
rect 45810 1696 45866 1698
rect 47490 1750 47546 1752
rect 47490 1698 47492 1750
rect 47492 1698 47544 1750
rect 47544 1698 47546 1750
rect 47490 1696 47546 1698
rect 49170 1750 49226 1752
rect 49170 1698 49172 1750
rect 49172 1698 49224 1750
rect 49224 1698 49226 1750
rect 49170 1696 49226 1698
rect 50850 1750 50906 1752
rect 50850 1698 50852 1750
rect 50852 1698 50904 1750
rect 50904 1698 50906 1750
rect 50850 1696 50906 1698
rect 52530 1750 52586 1752
rect 52530 1698 52532 1750
rect 52532 1698 52584 1750
rect 52584 1698 52586 1750
rect 52530 1696 52586 1698
rect 54210 1750 54266 1752
rect 54210 1698 54212 1750
rect 54212 1698 54264 1750
rect 54264 1698 54266 1750
rect 54210 1696 54266 1698
rect 55890 1750 55946 1752
rect 55890 1698 55892 1750
rect 55892 1698 55944 1750
rect 55944 1698 55946 1750
rect 55890 1696 55946 1698
rect 57570 1750 57626 1752
rect 57570 1698 57572 1750
rect 57572 1698 57624 1750
rect 57624 1698 57626 1750
rect 57570 1696 57626 1698
rect 59250 1750 59306 1752
rect 59250 1698 59252 1750
rect 59252 1698 59304 1750
rect 59304 1698 59306 1750
rect 59250 1696 59306 1698
rect 60930 1750 60986 1752
rect 60930 1698 60932 1750
rect 60932 1698 60984 1750
rect 60984 1698 60986 1750
rect 60930 1696 60986 1698
rect 62610 1750 62666 1752
rect 62610 1698 62612 1750
rect 62612 1698 62664 1750
rect 62664 1698 62666 1750
rect 62610 1696 62666 1698
rect 64290 1750 64346 1752
rect 64290 1698 64292 1750
rect 64292 1698 64344 1750
rect 64344 1698 64346 1750
rect 64290 1696 64346 1698
rect 65970 1750 66026 1752
rect 65970 1698 65972 1750
rect 65972 1698 66024 1750
rect 66024 1698 66026 1750
rect 65970 1696 66026 1698
rect 67650 1750 67706 1752
rect 67650 1698 67652 1750
rect 67652 1698 67704 1750
rect 67704 1698 67706 1750
rect 67650 1696 67706 1698
rect 69330 1750 69386 1752
rect 69330 1698 69332 1750
rect 69332 1698 69384 1750
rect 69384 1698 69386 1750
rect 69330 1696 69386 1698
rect 71010 1750 71066 1752
rect 71010 1698 71012 1750
rect 71012 1698 71064 1750
rect 71064 1698 71066 1750
rect 71010 1696 71066 1698
rect 72690 1750 72746 1752
rect 72690 1698 72692 1750
rect 72692 1698 72744 1750
rect 72744 1698 72746 1750
rect 72690 1696 72746 1698
rect 74370 1750 74426 1752
rect 74370 1698 74372 1750
rect 74372 1698 74424 1750
rect 74424 1698 74426 1750
rect 74370 1696 74426 1698
rect 76050 1750 76106 1752
rect 76050 1698 76052 1750
rect 76052 1698 76104 1750
rect 76104 1698 76106 1750
rect 76050 1696 76106 1698
rect 77730 1750 77786 1752
rect 77730 1698 77732 1750
rect 77732 1698 77784 1750
rect 77784 1698 77786 1750
rect 77730 1696 77786 1698
rect 79410 1750 79466 1752
rect 79410 1698 79412 1750
rect 79412 1698 79464 1750
rect 79464 1698 79466 1750
rect 79410 1696 79466 1698
rect 81090 1750 81146 1752
rect 81090 1698 81092 1750
rect 81092 1698 81144 1750
rect 81144 1698 81146 1750
rect 81090 1696 81146 1698
rect 82770 1750 82826 1752
rect 82770 1698 82772 1750
rect 82772 1698 82824 1750
rect 82824 1698 82826 1750
rect 82770 1696 82826 1698
rect 84450 1750 84506 1752
rect 84450 1698 84452 1750
rect 84452 1698 84504 1750
rect 84504 1698 84506 1750
rect 84450 1696 84506 1698
rect 86130 1750 86186 1752
rect 86130 1698 86132 1750
rect 86132 1698 86184 1750
rect 86184 1698 86186 1750
rect 86130 1696 86186 1698
rect 87810 1750 87866 1752
rect 87810 1698 87812 1750
rect 87812 1698 87864 1750
rect 87864 1698 87866 1750
rect 87810 1696 87866 1698
rect 89490 1750 89546 1752
rect 89490 1698 89492 1750
rect 89492 1698 89544 1750
rect 89544 1698 89546 1750
rect 89490 1696 89546 1698
rect 91170 1750 91226 1752
rect 91170 1698 91172 1750
rect 91172 1698 91224 1750
rect 91224 1698 91226 1750
rect 91170 1696 91226 1698
rect 92850 1750 92906 1752
rect 92850 1698 92852 1750
rect 92852 1698 92904 1750
rect 92904 1698 92906 1750
rect 92850 1696 92906 1698
rect 94530 1750 94586 1752
rect 94530 1698 94532 1750
rect 94532 1698 94584 1750
rect 94584 1698 94586 1750
rect 94530 1696 94586 1698
rect 96210 1750 96266 1752
rect 96210 1698 96212 1750
rect 96212 1698 96264 1750
rect 96264 1698 96266 1750
rect 96210 1696 96266 1698
rect 97890 1750 97946 1752
rect 97890 1698 97892 1750
rect 97892 1698 97944 1750
rect 97944 1698 97946 1750
rect 97890 1696 97946 1698
rect 99570 1750 99626 1752
rect 99570 1698 99572 1750
rect 99572 1698 99624 1750
rect 99624 1698 99626 1750
rect 99570 1696 99626 1698
rect 101250 1750 101306 1752
rect 101250 1698 101252 1750
rect 101252 1698 101304 1750
rect 101304 1698 101306 1750
rect 101250 1696 101306 1698
rect 102930 1750 102986 1752
rect 102930 1698 102932 1750
rect 102932 1698 102984 1750
rect 102984 1698 102986 1750
rect 102930 1696 102986 1698
rect 104610 1750 104666 1752
rect 104610 1698 104612 1750
rect 104612 1698 104664 1750
rect 104664 1698 104666 1750
rect 104610 1696 104666 1698
rect 106290 1750 106346 1752
rect 106290 1698 106292 1750
rect 106292 1698 106344 1750
rect 106344 1698 106346 1750
rect 106290 1696 106346 1698
rect 107970 1750 108026 1752
rect 107970 1698 107972 1750
rect 107972 1698 108024 1750
rect 108024 1698 108026 1750
rect 107970 1696 108026 1698
rect 109650 1750 109706 1752
rect 109650 1698 109652 1750
rect 109652 1698 109704 1750
rect 109704 1698 109706 1750
rect 109650 1696 109706 1698
rect 111330 1750 111386 1752
rect 111330 1698 111332 1750
rect 111332 1698 111384 1750
rect 111384 1698 111386 1750
rect 111330 1696 111386 1698
rect 113010 1750 113066 1752
rect 113010 1698 113012 1750
rect 113012 1698 113064 1750
rect 113064 1698 113066 1750
rect 113010 1696 113066 1698
rect 114690 1750 114746 1752
rect 114690 1698 114692 1750
rect 114692 1698 114744 1750
rect 114744 1698 114746 1750
rect 114690 1696 114746 1698
rect 116370 1750 116426 1752
rect 116370 1698 116372 1750
rect 116372 1698 116424 1750
rect 116424 1698 116426 1750
rect 116370 1696 116426 1698
rect 118050 1750 118106 1752
rect 118050 1698 118052 1750
rect 118052 1698 118104 1750
rect 118104 1698 118106 1750
rect 118050 1696 118106 1698
rect 119730 1750 119786 1752
rect 119730 1698 119732 1750
rect 119732 1698 119784 1750
rect 119784 1698 119786 1750
rect 119730 1696 119786 1698
rect 121410 1750 121466 1752
rect 121410 1698 121412 1750
rect 121412 1698 121464 1750
rect 121464 1698 121466 1750
rect 121410 1696 121466 1698
rect 123090 1750 123146 1752
rect 123090 1698 123092 1750
rect 123092 1698 123144 1750
rect 123144 1698 123146 1750
rect 123090 1696 123146 1698
rect 124770 1750 124826 1752
rect 124770 1698 124772 1750
rect 124772 1698 124824 1750
rect 124824 1698 124826 1750
rect 124770 1696 124826 1698
rect 126450 1750 126506 1752
rect 126450 1698 126452 1750
rect 126452 1698 126504 1750
rect 126504 1698 126506 1750
rect 126450 1696 126506 1698
rect 128130 1750 128186 1752
rect 128130 1698 128132 1750
rect 128132 1698 128184 1750
rect 128184 1698 128186 1750
rect 128130 1696 128186 1698
rect 129810 1750 129866 1752
rect 129810 1698 129812 1750
rect 129812 1698 129864 1750
rect 129864 1698 129866 1750
rect 129810 1696 129866 1698
rect 131490 1750 131546 1752
rect 131490 1698 131492 1750
rect 131492 1698 131544 1750
rect 131544 1698 131546 1750
rect 131490 1696 131546 1698
rect 133170 1750 133226 1752
rect 133170 1698 133172 1750
rect 133172 1698 133224 1750
rect 133224 1698 133226 1750
rect 133170 1696 133226 1698
<< metal3 >>
rect 272 83030 136348 83036
rect 272 82966 278 83030
rect 342 82966 414 83030
rect 478 82966 550 83030
rect 614 82966 136006 83030
rect 136070 82966 136142 83030
rect 136206 82966 136278 83030
rect 136342 82966 136348 83030
rect 272 82894 136348 82966
rect 272 82830 278 82894
rect 342 82830 414 82894
rect 478 82830 550 82894
rect 614 82830 136006 82894
rect 136070 82830 136142 82894
rect 136206 82830 136278 82894
rect 136342 82830 136348 82894
rect 272 82758 136348 82830
rect 272 82694 278 82758
rect 342 82694 414 82758
rect 478 82694 550 82758
rect 614 82694 118054 82758
rect 118118 82694 136006 82758
rect 136070 82694 136142 82758
rect 136206 82694 136278 82758
rect 136342 82694 136348 82758
rect 272 82688 136348 82694
rect 952 82350 135668 82356
rect 952 82286 958 82350
rect 1022 82286 1094 82350
rect 1158 82286 1230 82350
rect 1294 82286 135326 82350
rect 135390 82286 135462 82350
rect 135526 82286 135598 82350
rect 135662 82286 135668 82350
rect 952 82214 135668 82286
rect 952 82150 958 82214
rect 1022 82150 1094 82214
rect 1158 82150 1230 82214
rect 1294 82150 135326 82214
rect 135390 82150 135462 82214
rect 135526 82150 135598 82214
rect 135662 82150 135668 82214
rect 952 82078 135668 82150
rect 952 82014 958 82078
rect 1022 82014 1094 82078
rect 1158 82014 1230 82078
rect 1294 82014 2182 82078
rect 2246 82014 3950 82078
rect 4014 82014 5446 82078
rect 5510 82014 7214 82078
rect 7278 82014 8710 82078
rect 8774 82014 10478 82078
rect 10542 82014 12110 82078
rect 12174 82014 14014 82078
rect 14078 82014 15646 82078
rect 15710 82014 17142 82078
rect 17206 82014 18910 82078
rect 18974 82014 20678 82078
rect 20742 82014 22174 82078
rect 22238 82014 23942 82078
rect 24006 82014 25710 82078
rect 25774 82014 27206 82078
rect 27270 82014 28974 82078
rect 29038 82014 30606 82078
rect 30670 82014 32374 82078
rect 32438 82014 34142 82078
rect 34206 82014 35638 82078
rect 35702 82014 37542 82078
rect 37606 82014 39174 82078
rect 39238 82014 40670 82078
rect 40734 82014 42438 82078
rect 42502 82014 44206 82078
rect 44270 82014 45702 82078
rect 45766 82014 47470 82078
rect 47534 82014 49238 82078
rect 49302 82014 50734 82078
rect 50798 82014 52638 82078
rect 52702 82014 54134 82078
rect 54198 82014 55902 82078
rect 55966 82014 57670 82078
rect 57734 82014 59166 82078
rect 59230 82014 60798 82078
rect 60862 82014 62702 82078
rect 62766 82014 64198 82078
rect 64262 82014 65830 82078
rect 65894 82014 67598 82078
rect 67662 82014 69230 82078
rect 69294 82014 70862 82078
rect 70926 82014 72630 82078
rect 72694 82014 74398 82078
rect 74462 82014 76166 82078
rect 76230 82014 77662 82078
rect 77726 82014 79430 82078
rect 79494 82014 81334 82078
rect 81398 82014 82694 82078
rect 82758 82014 84462 82078
rect 84526 82014 86230 82078
rect 86294 82014 87726 82078
rect 87790 82014 89358 82078
rect 89422 82014 91126 82078
rect 91190 82014 92894 82078
rect 92958 82014 94390 82078
rect 94454 82014 96294 82078
rect 96358 82014 97926 82078
rect 97990 82014 99694 82078
rect 99758 82014 101326 82078
rect 101390 82014 102958 82078
rect 103022 82014 104590 82078
rect 104654 82014 106358 82078
rect 106422 82014 107854 82078
rect 107918 82014 109622 82078
rect 109686 82014 111390 82078
rect 111454 82014 112886 82078
rect 112950 82014 114654 82078
rect 114718 82014 116422 82078
rect 116486 82014 117918 82078
rect 117982 82014 119550 82078
rect 119614 82014 121454 82078
rect 121518 82014 123222 82078
rect 123286 82014 124718 82078
rect 124782 82014 126350 82078
rect 126414 82014 128118 82078
rect 128182 82014 129886 82078
rect 129950 82014 131382 82078
rect 131446 82014 133150 82078
rect 133214 82014 135326 82078
rect 135390 82014 135462 82078
rect 135526 82014 135598 82078
rect 135662 82014 135668 82078
rect 952 82008 135668 82014
rect 2040 81534 2252 81540
rect 2040 81501 2182 81534
rect 2040 81445 2130 81501
rect 2246 81470 2252 81534
rect 2186 81445 2252 81470
rect 2040 81398 2252 81445
rect 2040 81334 2046 81398
rect 2110 81334 2252 81398
rect 2040 81328 2252 81334
rect 3672 81534 4020 81540
rect 3672 81501 3950 81534
rect 3672 81445 3810 81501
rect 3866 81470 3950 81501
rect 4014 81470 4020 81534
rect 3866 81445 4020 81470
rect 3672 81328 4020 81445
rect 5440 81534 5652 81540
rect 5440 81470 5446 81534
rect 5510 81501 5652 81534
rect 5440 81445 5490 81470
rect 5546 81445 5652 81501
rect 5440 81328 5652 81445
rect 7072 81534 7284 81540
rect 7072 81501 7214 81534
rect 7072 81445 7170 81501
rect 7278 81470 7284 81534
rect 7226 81445 7284 81470
rect 7072 81328 7284 81445
rect 8704 81534 9052 81540
rect 8704 81470 8710 81534
rect 8774 81501 9052 81534
rect 8774 81470 8850 81501
rect 8704 81445 8850 81470
rect 8906 81445 9052 81501
rect 8704 81328 9052 81445
rect 10472 81534 10684 81540
rect 10472 81470 10478 81534
rect 10542 81501 10684 81534
rect 10472 81445 10530 81470
rect 10586 81445 10684 81501
rect 10472 81328 10684 81445
rect 12104 81534 12316 81540
rect 12104 81470 12110 81534
rect 12174 81501 12316 81534
rect 12174 81470 12210 81501
rect 12104 81445 12210 81470
rect 12266 81445 12316 81501
rect 12104 81328 12316 81445
rect 13736 81534 14084 81540
rect 13736 81501 14014 81534
rect 13736 81445 13890 81501
rect 13946 81470 14014 81501
rect 14078 81470 14084 81534
rect 13946 81445 14084 81470
rect 13736 81328 14084 81445
rect 15504 81534 15716 81540
rect 15504 81501 15646 81534
rect 15504 81445 15570 81501
rect 15626 81470 15646 81501
rect 15710 81470 15716 81534
rect 15626 81445 15716 81470
rect 15504 81328 15716 81445
rect 17136 81534 17348 81540
rect 17136 81470 17142 81534
rect 17206 81501 17348 81534
rect 17206 81470 17250 81501
rect 17136 81445 17250 81470
rect 17306 81445 17348 81501
rect 17136 81328 17348 81445
rect 18904 81534 19116 81540
rect 18904 81470 18910 81534
rect 18974 81501 19116 81534
rect 18904 81445 18930 81470
rect 18986 81445 19116 81501
rect 18904 81328 19116 81445
rect 20536 81534 20748 81540
rect 20536 81501 20678 81534
rect 20536 81445 20610 81501
rect 20666 81470 20678 81501
rect 20742 81470 20748 81534
rect 20666 81445 20748 81470
rect 20536 81328 20748 81445
rect 22168 81534 22380 81540
rect 22168 81470 22174 81534
rect 22238 81501 22380 81534
rect 22238 81470 22290 81501
rect 22168 81445 22290 81470
rect 22346 81445 22380 81501
rect 22168 81328 22380 81445
rect 23936 81534 24148 81540
rect 23936 81470 23942 81534
rect 24006 81501 24148 81534
rect 23936 81445 23970 81470
rect 24026 81445 24148 81501
rect 23936 81328 24148 81445
rect 25568 81534 25780 81540
rect 25568 81501 25710 81534
rect 25568 81445 25650 81501
rect 25706 81470 25710 81501
rect 25774 81470 25780 81534
rect 25706 81445 25780 81470
rect 25568 81328 25780 81445
rect 27200 81534 27412 81540
rect 27200 81470 27206 81534
rect 27270 81501 27412 81534
rect 27270 81470 27330 81501
rect 27200 81445 27330 81470
rect 27386 81445 27412 81501
rect 27200 81328 27412 81445
rect 28968 81534 29180 81540
rect 28968 81470 28974 81534
rect 29038 81501 29180 81534
rect 28968 81445 29010 81470
rect 29066 81445 29180 81501
rect 28968 81328 29180 81445
rect 30600 81534 30812 81540
rect 30600 81470 30606 81534
rect 30670 81501 30812 81534
rect 30670 81470 30690 81501
rect 30600 81445 30690 81470
rect 30746 81445 30812 81501
rect 30600 81328 30812 81445
rect 32232 81534 32580 81540
rect 32232 81501 32374 81534
rect 32232 81445 32370 81501
rect 32438 81470 32580 81534
rect 32426 81445 32580 81470
rect 32232 81328 32580 81445
rect 34000 81534 34212 81540
rect 34000 81501 34142 81534
rect 34000 81445 34050 81501
rect 34106 81470 34142 81501
rect 34206 81470 34212 81534
rect 34106 81445 34212 81470
rect 34000 81328 34212 81445
rect 35632 81534 35844 81540
rect 35632 81470 35638 81534
rect 35702 81501 35844 81534
rect 35702 81470 35730 81501
rect 35632 81445 35730 81470
rect 35786 81445 35844 81501
rect 35632 81328 35844 81445
rect 37264 81534 37612 81540
rect 37264 81501 37542 81534
rect 37264 81445 37410 81501
rect 37466 81470 37542 81501
rect 37606 81470 37612 81534
rect 37466 81445 37612 81470
rect 37264 81328 37612 81445
rect 39032 81534 39244 81540
rect 39032 81501 39174 81534
rect 39032 81445 39090 81501
rect 39146 81470 39174 81501
rect 39238 81470 39244 81534
rect 39146 81445 39244 81470
rect 39032 81328 39244 81445
rect 40664 81534 40876 81540
rect 40664 81470 40670 81534
rect 40734 81501 40876 81534
rect 40734 81470 40770 81501
rect 40664 81445 40770 81470
rect 40826 81445 40876 81501
rect 40664 81328 40876 81445
rect 42296 81534 42644 81540
rect 42296 81470 42438 81534
rect 42502 81501 42644 81534
rect 42296 81445 42450 81470
rect 42506 81445 42644 81501
rect 42296 81328 42644 81445
rect 44064 81534 44276 81540
rect 44064 81501 44206 81534
rect 44064 81445 44130 81501
rect 44186 81470 44206 81501
rect 44270 81470 44276 81534
rect 44186 81445 44276 81470
rect 44064 81328 44276 81445
rect 45696 81534 45908 81540
rect 45696 81470 45702 81534
rect 45766 81501 45908 81534
rect 45766 81470 45810 81501
rect 45696 81445 45810 81470
rect 45866 81445 45908 81501
rect 45696 81328 45908 81445
rect 47464 81534 47676 81540
rect 47464 81470 47470 81534
rect 47534 81501 47676 81534
rect 47464 81445 47490 81470
rect 47546 81445 47676 81501
rect 47464 81328 47676 81445
rect 49096 81534 49308 81540
rect 49096 81501 49238 81534
rect 49096 81445 49170 81501
rect 49226 81470 49238 81501
rect 49302 81470 49308 81534
rect 49226 81445 49308 81470
rect 49096 81328 49308 81445
rect 50728 81534 50940 81540
rect 50728 81470 50734 81534
rect 50798 81501 50940 81534
rect 50798 81470 50850 81501
rect 50728 81445 50850 81470
rect 50906 81445 50940 81501
rect 50728 81328 50940 81445
rect 52496 81534 52708 81540
rect 52496 81501 52638 81534
rect 52496 81445 52530 81501
rect 52586 81470 52638 81501
rect 52702 81470 52708 81534
rect 52586 81445 52708 81470
rect 52496 81328 52708 81445
rect 54128 81534 54340 81540
rect 54128 81470 54134 81534
rect 54198 81501 54340 81534
rect 54198 81470 54210 81501
rect 54128 81445 54210 81470
rect 54266 81445 54340 81501
rect 54128 81328 54340 81445
rect 55760 81534 55972 81540
rect 55760 81501 55902 81534
rect 55760 81445 55890 81501
rect 55966 81470 55972 81534
rect 55946 81445 55972 81470
rect 55760 81328 55972 81445
rect 57528 81534 57740 81540
rect 57528 81501 57670 81534
rect 57528 81445 57570 81501
rect 57626 81470 57670 81501
rect 57734 81470 57740 81534
rect 57626 81445 57740 81470
rect 57528 81328 57740 81445
rect 59160 81534 59372 81540
rect 59160 81470 59166 81534
rect 59230 81501 59372 81534
rect 59230 81470 59250 81501
rect 59160 81445 59250 81470
rect 59306 81445 59372 81501
rect 59160 81328 59372 81445
rect 60792 81534 61140 81540
rect 60792 81470 60798 81534
rect 60862 81501 61140 81534
rect 60862 81470 60930 81501
rect 60792 81445 60930 81470
rect 60986 81445 61140 81501
rect 60792 81328 61140 81445
rect 62560 81534 62772 81540
rect 62560 81501 62702 81534
rect 62560 81445 62610 81501
rect 62666 81470 62702 81501
rect 62766 81470 62772 81534
rect 62666 81445 62772 81470
rect 62560 81328 62772 81445
rect 64192 81534 64404 81540
rect 64192 81470 64198 81534
rect 64262 81501 64404 81534
rect 64262 81470 64290 81501
rect 64192 81445 64290 81470
rect 64346 81445 64404 81501
rect 64192 81328 64404 81445
rect 65824 81534 66172 81540
rect 65824 81470 65830 81534
rect 65894 81501 66172 81534
rect 65894 81470 65970 81501
rect 65824 81445 65970 81470
rect 66026 81445 66172 81501
rect 65824 81328 66172 81445
rect 67592 81534 67804 81540
rect 67592 81470 67598 81534
rect 67662 81501 67804 81534
rect 67592 81445 67650 81470
rect 67706 81445 67804 81501
rect 67592 81328 67804 81445
rect 69224 81534 69436 81540
rect 69224 81470 69230 81534
rect 69294 81501 69436 81534
rect 69294 81470 69330 81501
rect 69224 81445 69330 81470
rect 69386 81445 69436 81501
rect 69224 81328 69436 81445
rect 70856 81534 71204 81540
rect 70856 81470 70862 81534
rect 70926 81501 71204 81534
rect 70926 81470 71010 81501
rect 70856 81445 71010 81470
rect 71066 81445 71204 81501
rect 70856 81328 71204 81445
rect 72624 81534 72836 81540
rect 72624 81470 72630 81534
rect 72694 81501 72836 81534
rect 72624 81445 72690 81470
rect 72746 81445 72836 81501
rect 72624 81328 72836 81445
rect 74256 81534 74468 81540
rect 74256 81501 74398 81534
rect 74256 81445 74370 81501
rect 74462 81470 74468 81534
rect 74426 81445 74468 81470
rect 74256 81328 74468 81445
rect 76024 81534 76236 81540
rect 76024 81501 76166 81534
rect 76024 81445 76050 81501
rect 76106 81470 76166 81501
rect 76230 81470 76236 81534
rect 76106 81445 76236 81470
rect 76024 81328 76236 81445
rect 77656 81534 77868 81540
rect 77656 81470 77662 81534
rect 77726 81501 77868 81534
rect 77726 81470 77730 81501
rect 77656 81445 77730 81470
rect 77786 81445 77868 81501
rect 77656 81328 77868 81445
rect 79288 81534 79500 81540
rect 79288 81501 79430 81534
rect 79288 81445 79410 81501
rect 79494 81470 79500 81534
rect 79466 81445 79500 81470
rect 79288 81328 79500 81445
rect 81056 81534 81404 81540
rect 81056 81501 81334 81534
rect 81056 81445 81090 81501
rect 81146 81470 81334 81501
rect 81398 81470 81404 81534
rect 81146 81464 81404 81470
rect 82688 81534 82900 81540
rect 82688 81470 82694 81534
rect 82758 81501 82900 81534
rect 82758 81470 82770 81501
rect 81146 81445 81268 81464
rect 81056 81328 81268 81445
rect 82688 81445 82770 81470
rect 82826 81445 82900 81501
rect 82688 81328 82900 81445
rect 84320 81534 84532 81540
rect 84320 81501 84462 81534
rect 84320 81445 84450 81501
rect 84526 81470 84532 81534
rect 84506 81445 84532 81470
rect 84320 81328 84532 81445
rect 86088 81534 86300 81540
rect 86088 81501 86230 81534
rect 86088 81445 86130 81501
rect 86186 81470 86230 81501
rect 86294 81470 86300 81534
rect 86186 81445 86300 81470
rect 86088 81328 86300 81445
rect 87720 81534 87932 81540
rect 87720 81470 87726 81534
rect 87790 81501 87932 81534
rect 87790 81470 87810 81501
rect 87720 81445 87810 81470
rect 87866 81445 87932 81501
rect 87720 81328 87932 81445
rect 89352 81534 89700 81540
rect 89352 81470 89358 81534
rect 89422 81501 89700 81534
rect 89422 81470 89490 81501
rect 89352 81445 89490 81470
rect 89546 81445 89700 81501
rect 89352 81328 89700 81445
rect 91120 81534 91332 81540
rect 91120 81470 91126 81534
rect 91190 81501 91332 81534
rect 91120 81445 91170 81470
rect 91226 81445 91332 81501
rect 91120 81328 91332 81445
rect 92752 81534 92964 81540
rect 92752 81501 92894 81534
rect 92752 81445 92850 81501
rect 92958 81470 92964 81534
rect 92906 81445 92964 81470
rect 92752 81328 92964 81445
rect 94384 81534 94732 81540
rect 94384 81470 94390 81534
rect 94454 81501 94732 81534
rect 94454 81470 94530 81501
rect 94384 81445 94530 81470
rect 94586 81445 94732 81501
rect 94384 81328 94732 81445
rect 96152 81534 96364 81540
rect 96152 81501 96294 81534
rect 96152 81445 96210 81501
rect 96266 81470 96294 81501
rect 96358 81470 96364 81534
rect 96266 81445 96364 81470
rect 96152 81328 96364 81445
rect 97784 81534 97996 81540
rect 97784 81501 97926 81534
rect 97784 81445 97890 81501
rect 97990 81470 97996 81534
rect 97946 81445 97996 81470
rect 97784 81328 97996 81445
rect 99416 81534 99764 81540
rect 99416 81501 99694 81534
rect 99416 81445 99570 81501
rect 99626 81470 99694 81501
rect 99758 81470 99764 81534
rect 99626 81445 99764 81470
rect 99416 81328 99764 81445
rect 101184 81534 101396 81540
rect 101184 81501 101326 81534
rect 101184 81445 101250 81501
rect 101306 81470 101326 81501
rect 101390 81470 101396 81534
rect 101306 81445 101396 81470
rect 101184 81328 101396 81445
rect 102816 81534 103028 81540
rect 102816 81501 102958 81534
rect 102816 81445 102930 81501
rect 103022 81470 103028 81534
rect 102986 81445 103028 81470
rect 102816 81328 103028 81445
rect 104584 81534 104796 81540
rect 104584 81470 104590 81534
rect 104654 81501 104796 81534
rect 104584 81445 104610 81470
rect 104666 81445 104796 81501
rect 104584 81328 104796 81445
rect 106216 81534 106428 81540
rect 106216 81501 106358 81534
rect 106216 81445 106290 81501
rect 106346 81470 106358 81501
rect 106422 81470 106428 81534
rect 106346 81445 106428 81470
rect 106216 81328 106428 81445
rect 107848 81534 108060 81540
rect 107848 81470 107854 81534
rect 107918 81501 108060 81534
rect 107918 81470 107970 81501
rect 107848 81445 107970 81470
rect 108026 81445 108060 81501
rect 107848 81328 108060 81445
rect 109616 81534 109828 81540
rect 109616 81470 109622 81534
rect 109686 81501 109828 81534
rect 109616 81445 109650 81470
rect 109706 81445 109828 81501
rect 109616 81328 109828 81445
rect 111248 81534 111460 81540
rect 111248 81501 111390 81534
rect 111248 81445 111330 81501
rect 111386 81470 111390 81501
rect 111454 81470 111460 81534
rect 111386 81445 111460 81470
rect 111248 81328 111460 81445
rect 112880 81534 113092 81540
rect 112880 81470 112886 81534
rect 112950 81501 113092 81534
rect 112950 81470 113010 81501
rect 112880 81445 113010 81470
rect 113066 81445 113092 81501
rect 112880 81328 113092 81445
rect 114648 81534 114860 81540
rect 114648 81470 114654 81534
rect 114718 81501 114860 81534
rect 114648 81445 114690 81470
rect 114746 81445 114860 81501
rect 114648 81328 114860 81445
rect 116280 81534 116492 81540
rect 116280 81501 116422 81534
rect 116280 81445 116370 81501
rect 116486 81470 116492 81534
rect 116426 81445 116492 81470
rect 116280 81328 116492 81445
rect 117912 81534 118260 81540
rect 117912 81470 117918 81534
rect 117982 81501 118260 81534
rect 117982 81470 118050 81501
rect 117912 81445 118050 81470
rect 118106 81445 118260 81501
rect 119544 81534 119892 81540
rect 119544 81470 119550 81534
rect 119614 81501 119892 81534
rect 119614 81470 119730 81501
rect 119544 81464 119730 81470
rect 117912 81398 118260 81445
rect 117912 81334 118190 81398
rect 118254 81334 118260 81398
rect 117912 81328 118260 81334
rect 119680 81445 119730 81464
rect 119786 81445 119892 81501
rect 119680 81328 119892 81445
rect 121312 81534 121524 81540
rect 121312 81501 121454 81534
rect 121312 81445 121410 81501
rect 121518 81470 121524 81534
rect 121466 81445 121524 81470
rect 121312 81328 121524 81445
rect 122944 81534 123292 81540
rect 122944 81501 123222 81534
rect 122944 81445 123090 81501
rect 123146 81470 123222 81501
rect 123286 81470 123292 81534
rect 123146 81445 123292 81470
rect 122944 81398 123292 81445
rect 122944 81334 122950 81398
rect 123014 81334 123292 81398
rect 122944 81328 123292 81334
rect 124712 81534 124924 81540
rect 124712 81470 124718 81534
rect 124782 81501 124924 81534
rect 124712 81445 124770 81470
rect 124826 81445 124924 81501
rect 124712 81328 124924 81445
rect 126344 81534 126556 81540
rect 126344 81470 126350 81534
rect 126414 81501 126556 81534
rect 126414 81470 126450 81501
rect 126344 81445 126450 81470
rect 126506 81445 126556 81501
rect 126344 81328 126556 81445
rect 127976 81534 128324 81540
rect 127976 81470 128118 81534
rect 128182 81501 128324 81534
rect 127976 81445 128130 81470
rect 128186 81445 128324 81501
rect 127976 81328 128324 81445
rect 129744 81534 129956 81540
rect 129744 81501 129886 81534
rect 129744 81445 129810 81501
rect 129866 81470 129886 81501
rect 129950 81470 129956 81534
rect 129866 81445 129956 81470
rect 129744 81328 129956 81445
rect 131376 81534 131588 81540
rect 131376 81470 131382 81534
rect 131446 81501 131588 81534
rect 131446 81470 131490 81501
rect 131376 81445 131490 81470
rect 131546 81445 131588 81501
rect 131376 81328 131588 81445
rect 133144 81534 133356 81540
rect 133144 81470 133150 81534
rect 133214 81501 133356 81534
rect 133144 81445 133170 81470
rect 133226 81445 133356 81501
rect 133144 81328 133356 81445
rect 1768 81126 2116 81132
rect 1768 81062 2046 81126
rect 2110 81062 2116 81126
rect 1768 81056 2116 81062
rect 1768 81048 1980 81056
rect 1768 80992 1794 81048
rect 1850 80992 1980 81048
rect 1768 80920 1980 80992
rect 134776 81048 134988 81132
rect 134776 80992 134844 81048
rect 134900 80996 134988 81048
rect 134900 80992 135396 80996
rect 134776 80990 135396 80992
rect 134776 80926 135326 80990
rect 135390 80926 135396 80990
rect 134776 80920 135396 80926
rect 118048 80854 118396 80860
rect 118048 80790 118054 80854
rect 118118 80790 118396 80854
rect 118048 80724 118396 80790
rect 119272 80724 119484 80860
rect 117950 80718 122340 80724
rect 117912 80654 117918 80718
rect 117982 80654 122270 80718
rect 122334 80654 122340 80718
rect 117950 80648 122340 80654
rect 122183 80523 122249 80526
rect 118796 80521 122249 80523
rect 118796 80465 122188 80521
rect 122244 80465 122249 80521
rect 118796 80463 122249 80465
rect 122183 80460 122249 80463
rect 118456 80310 118804 80316
rect 118456 80246 118462 80310
rect 118526 80265 118804 80310
rect 118526 80246 118598 80265
rect 118456 80209 118598 80246
rect 118654 80209 118804 80265
rect 118456 80104 118804 80209
rect 119680 80310 119892 80316
rect 119680 80246 119686 80310
rect 119750 80265 119892 80310
rect 119750 80246 119766 80265
rect 119680 80209 119766 80246
rect 119822 80209 119892 80265
rect 119680 80104 119892 80209
rect 122264 79902 122476 79908
rect 122264 79838 122270 79902
rect 122334 79838 122476 79902
rect 122264 79766 122476 79838
rect 122264 79702 122406 79766
rect 122470 79702 122476 79766
rect 122264 79696 122476 79702
rect 133960 79902 136076 79908
rect 133960 79838 136006 79902
rect 136070 79838 136076 79902
rect 133960 79832 136076 79838
rect 133960 79696 134172 79832
rect 1224 79494 1980 79500
rect 1224 79430 1230 79494
rect 1294 79430 1980 79494
rect 1224 79424 1980 79430
rect 1768 79368 1980 79424
rect 1768 79312 1794 79368
rect 1850 79312 1980 79368
rect 1768 79288 1980 79312
rect 118048 79494 118396 79500
rect 118048 79430 118190 79494
rect 118254 79430 118396 79494
rect 118048 79364 118396 79430
rect 119272 79364 119484 79500
rect 134776 79494 135396 79500
rect 134776 79430 135326 79494
rect 135390 79430 135396 79494
rect 134776 79424 135396 79430
rect 134823 79368 134921 79424
rect 118048 79358 119484 79364
rect 118048 79294 118054 79358
rect 118118 79294 119484 79358
rect 118048 79288 119484 79294
rect 133824 79268 134036 79364
rect 134823 79312 134844 79368
rect 134900 79312 134921 79368
rect 134823 79291 134921 79312
rect 130696 79222 130908 79228
rect 130696 79163 130838 79222
rect 130696 79107 130747 79163
rect 130803 79158 130838 79163
rect 130902 79158 130908 79222
rect 130803 79107 130908 79158
rect 133824 79212 133884 79268
rect 133940 79228 134036 79268
rect 133940 79212 136620 79228
rect 133824 79152 136620 79212
rect 130696 79016 130908 79107
rect 115328 78678 117988 78684
rect 115328 78614 117918 78678
rect 117982 78614 117988 78678
rect 115328 78608 117988 78614
rect 115328 78472 115540 78608
rect 116416 78542 116628 78608
rect 116416 78478 116558 78542
rect 116622 78478 116628 78542
rect 116416 78472 116628 78478
rect 122264 78542 123020 78548
rect 122264 78478 122950 78542
rect 123014 78478 123020 78542
rect 122264 78472 123020 78478
rect 122264 78406 122476 78472
rect 122264 78342 122270 78406
rect 122334 78342 122476 78406
rect 122264 78336 122476 78342
rect 133960 78412 134172 78548
rect 133960 78406 134852 78412
rect 133960 78342 134782 78406
rect 134846 78342 134852 78406
rect 133960 78336 134852 78342
rect 1768 77688 1980 77732
rect 1768 77632 1794 77688
rect 1850 77632 1980 77688
rect 1768 77596 1980 77632
rect 1224 77590 1980 77596
rect 1224 77526 1230 77590
rect 1294 77526 1980 77590
rect 1224 77520 1980 77526
rect 134776 77726 135396 77732
rect 134776 77662 134782 77726
rect 134846 77688 135326 77726
rect 134900 77662 135326 77688
rect 135390 77662 135396 77726
rect 134776 77632 134844 77662
rect 134900 77656 135396 77662
rect 134900 77632 134988 77656
rect 134776 77520 134988 77632
rect 115328 77318 118124 77324
rect 115328 77254 118054 77318
rect 118118 77254 118124 77318
rect 115328 77248 118124 77254
rect 28560 77182 28772 77188
rect 28560 77118 28702 77182
rect 28766 77118 28772 77182
rect 28560 77047 28772 77118
rect 28968 77087 29044 77188
rect 28560 76991 28618 77047
rect 28674 76991 28772 77047
rect 28560 76840 28772 76991
rect 28851 77046 29044 77087
rect 28851 76989 28974 77046
rect 28968 76982 28974 76989
rect 29038 76982 29044 77046
rect 28968 76976 29044 76982
rect 31008 77182 31220 77188
rect 31008 77118 31014 77182
rect 31078 77118 31220 77182
rect 31008 77047 31220 77118
rect 31008 76991 31114 77047
rect 31170 76991 31220 77047
rect 31008 76840 31220 76991
rect 31280 77046 31492 77188
rect 31280 76982 31422 77046
rect 31486 76982 31492 77046
rect 31280 76976 31492 76982
rect 33456 77182 33668 77188
rect 33456 77118 33462 77182
rect 33526 77118 33668 77182
rect 33456 77068 33668 77118
rect 33864 77087 34076 77188
rect 33456 77047 33687 77068
rect 33456 76991 33610 77047
rect 33666 76991 33687 77047
rect 33456 76916 33687 76991
rect 33843 77046 34076 77087
rect 33843 76989 34006 77046
rect 34000 76982 34006 76989
rect 34070 76982 34076 77046
rect 34000 76976 34076 76982
rect 36040 77182 36252 77188
rect 36040 77118 36182 77182
rect 36246 77118 36252 77182
rect 36040 77047 36252 77118
rect 36448 77087 36524 77188
rect 36040 76991 36106 77047
rect 36162 76991 36252 77047
rect 33456 76840 33804 76916
rect 36040 76840 36252 76991
rect 36339 77046 36524 77087
rect 36339 76989 36454 77046
rect 36448 76982 36454 76989
rect 36518 76982 36524 77046
rect 36448 76976 36524 76982
rect 38488 77182 38700 77188
rect 38488 77118 38494 77182
rect 38558 77118 38700 77182
rect 38488 77047 38700 77118
rect 38896 77087 38972 77188
rect 38488 76991 38602 77047
rect 38658 76991 38700 77047
rect 38488 76840 38700 76991
rect 38835 77052 38972 77087
rect 41072 77182 41148 77188
rect 41072 77118 41078 77182
rect 41142 77118 41148 77182
rect 41072 77068 41148 77118
rect 41344 77087 41556 77188
rect 38835 77046 39108 77052
rect 38835 76989 39038 77046
rect 38896 76982 39038 76989
rect 39102 76982 39108 77046
rect 38896 76976 39108 76982
rect 41072 77047 41175 77068
rect 41072 76991 41098 77047
rect 41154 76991 41175 77047
rect 41072 76916 41175 76991
rect 41331 77046 41556 77087
rect 41331 76989 41486 77046
rect 41344 76982 41486 76989
rect 41550 76982 41556 77046
rect 41344 76976 41556 76982
rect 43520 77182 43732 77188
rect 43520 77118 43526 77182
rect 43590 77118 43732 77182
rect 43520 77047 43732 77118
rect 43928 77087 44004 77188
rect 43520 76991 43594 77047
rect 43650 76991 43732 77047
rect 41072 76840 41284 76916
rect 43520 76840 43732 76991
rect 43827 77046 44004 77087
rect 43827 76989 43934 77046
rect 43928 76982 43934 76989
rect 43998 76982 44004 77046
rect 43928 76976 44004 76982
rect 45968 77182 46180 77188
rect 45968 77118 46110 77182
rect 46174 77118 46180 77182
rect 45968 77047 46180 77118
rect 46376 77087 46452 77188
rect 45968 76991 46090 77047
rect 46146 76991 46180 77047
rect 45968 76840 46180 76991
rect 46323 77052 46452 77087
rect 48552 77182 48628 77188
rect 48552 77118 48558 77182
rect 48622 77118 48628 77182
rect 48552 77068 48628 77118
rect 48824 77087 49036 77188
rect 46323 77046 46588 77052
rect 46323 76989 46518 77046
rect 46376 76982 46518 76989
rect 46582 76982 46588 77046
rect 46376 76976 46588 76982
rect 48552 77047 48663 77068
rect 48552 76991 48586 77047
rect 48642 76991 48663 77047
rect 48552 76916 48663 76991
rect 48819 77046 49036 77087
rect 48819 76989 48966 77046
rect 48960 76982 48966 76989
rect 49030 76982 49036 77046
rect 48960 76976 49036 76982
rect 51000 77182 51212 77188
rect 51000 77118 51142 77182
rect 51206 77118 51212 77182
rect 51000 77047 51212 77118
rect 51408 77087 51484 77188
rect 51000 76991 51082 77047
rect 51138 76991 51212 77047
rect 48552 76840 48764 76916
rect 51000 76840 51212 76991
rect 51315 77046 51484 77087
rect 51315 76989 51414 77046
rect 51408 76982 51414 76989
rect 51478 76982 51484 77046
rect 51408 76976 51484 76982
rect 53448 77182 53660 77188
rect 53448 77118 53590 77182
rect 53654 77118 53660 77182
rect 53448 77047 53660 77118
rect 53856 77087 53932 77188
rect 53448 76991 53578 77047
rect 53634 76991 53660 77047
rect 53448 76840 53660 76991
rect 53811 77046 53932 77087
rect 53811 76989 53862 77046
rect 53856 76982 53862 76989
rect 53926 76982 53932 77046
rect 53856 76976 53932 76982
rect 56032 77182 56244 77188
rect 56032 77118 56174 77182
rect 56238 77118 56244 77182
rect 56032 77047 56244 77118
rect 56032 76991 56074 77047
rect 56130 76991 56244 77047
rect 56032 76840 56244 76991
rect 56304 77046 56516 77188
rect 56304 76982 56446 77046
rect 56510 76982 56516 77046
rect 56304 76976 56516 76982
rect 58480 77182 58692 77188
rect 58480 77118 58486 77182
rect 58550 77118 58692 77182
rect 58480 77047 58692 77118
rect 58888 77087 58964 77188
rect 58480 76991 58570 77047
rect 58626 76991 58692 77047
rect 58480 76840 58692 76991
rect 58803 77046 58964 77087
rect 58803 76989 58894 77046
rect 58888 76982 58894 76989
rect 58958 76982 58964 77046
rect 58888 76976 58964 76982
rect 60928 77182 61140 77188
rect 60928 77118 60934 77182
rect 60998 77118 61140 77182
rect 61336 77182 61548 77188
rect 61336 77150 61478 77182
rect 60928 77068 61140 77118
rect 61299 77118 61478 77150
rect 61542 77118 61548 77182
rect 61299 77112 61548 77118
rect 63512 77182 63724 77188
rect 63512 77118 63654 77182
rect 63718 77118 63724 77182
rect 60928 77047 61143 77068
rect 60928 76991 61066 77047
rect 61122 76991 61143 77047
rect 60928 76916 61143 76991
rect 61299 76989 61397 77112
rect 63512 77047 63724 77118
rect 63920 77087 63996 77188
rect 63512 76991 63562 77047
rect 63618 76991 63724 77047
rect 60928 76840 61276 76916
rect 63512 76840 63724 76991
rect 63795 77046 63996 77087
rect 63795 76989 63926 77046
rect 63920 76982 63926 76989
rect 63990 76982 63996 77046
rect 63920 76976 63996 76982
rect 65960 77182 66172 77188
rect 65960 77118 66102 77182
rect 66166 77118 66172 77182
rect 65960 77047 66172 77118
rect 66368 77087 66444 77188
rect 65960 76991 66058 77047
rect 66114 76991 66172 77047
rect 65960 76840 66172 76991
rect 66291 77052 66444 77087
rect 68408 77182 68620 77188
rect 68408 77118 68550 77182
rect 68614 77118 68620 77182
rect 68816 77182 69028 77188
rect 68816 77150 68958 77182
rect 68408 77068 68620 77118
rect 68787 77118 68958 77150
rect 69022 77118 69028 77182
rect 68787 77112 69028 77118
rect 70992 77182 71204 77188
rect 70992 77118 70998 77182
rect 71062 77118 71204 77182
rect 66291 77046 66580 77052
rect 66291 76989 66510 77046
rect 66368 76982 66510 76989
rect 66574 76982 66580 77046
rect 66368 76976 66580 76982
rect 68408 77047 68631 77068
rect 68408 76991 68554 77047
rect 68610 76991 68631 77047
rect 68408 76916 68631 76991
rect 68787 76989 68885 77112
rect 70992 77047 71204 77118
rect 71400 77087 71476 77188
rect 70992 76991 71050 77047
rect 71106 76991 71204 77047
rect 68408 76840 68756 76916
rect 70992 76840 71204 76991
rect 71283 77046 71476 77087
rect 71283 76989 71406 77046
rect 71400 76982 71406 76989
rect 71470 76982 71476 77046
rect 71400 76976 71476 76982
rect 73440 77182 73652 77188
rect 73440 77118 73582 77182
rect 73646 77118 73652 77182
rect 73440 77047 73652 77118
rect 73848 77087 73924 77188
rect 73440 76991 73546 77047
rect 73602 76991 73652 77047
rect 73440 76840 73652 76991
rect 73779 77046 73924 77087
rect 73779 76989 73854 77046
rect 73848 76982 73854 76989
rect 73918 76982 73924 77046
rect 73848 76976 73924 76982
rect 75888 77182 76100 77188
rect 75888 77118 75894 77182
rect 75958 77118 76100 77182
rect 75888 77068 76100 77118
rect 76296 77087 76508 77188
rect 75888 77047 76119 77068
rect 75888 76991 76042 77047
rect 76098 76991 76119 77047
rect 75888 76916 76119 76991
rect 76275 77046 76508 77087
rect 76275 76989 76438 77046
rect 76432 76982 76438 76989
rect 76502 76982 76508 77046
rect 76432 76976 76508 76982
rect 78472 77182 78684 77188
rect 78472 77118 78614 77182
rect 78678 77118 78684 77182
rect 78472 77047 78684 77118
rect 78880 77087 78956 77188
rect 78472 76991 78538 77047
rect 78594 76991 78684 77047
rect 75888 76840 76236 76916
rect 78472 76840 78684 76991
rect 78771 77046 78956 77087
rect 78771 76989 78886 77046
rect 78880 76982 78886 76989
rect 78950 76982 78956 77046
rect 78880 76976 78956 76982
rect 80920 77182 81132 77188
rect 80920 77118 81062 77182
rect 81126 77118 81132 77182
rect 80920 77047 81132 77118
rect 81328 77087 81404 77188
rect 80920 76991 81034 77047
rect 81090 76991 81132 77047
rect 80920 76840 81132 76991
rect 81267 77052 81404 77087
rect 83504 77182 83580 77188
rect 83504 77118 83510 77182
rect 83574 77118 83580 77182
rect 83504 77068 83580 77118
rect 83776 77087 83988 77188
rect 81267 77046 81540 77052
rect 81267 76989 81470 77046
rect 81328 76982 81470 76989
rect 81534 76982 81540 77046
rect 81328 76976 81540 76982
rect 83504 77047 83607 77068
rect 83504 76991 83530 77047
rect 83586 76991 83607 77047
rect 83504 76916 83607 76991
rect 83763 77046 83988 77087
rect 83763 76989 83918 77046
rect 83912 76982 83918 76989
rect 83982 76982 83988 77046
rect 83912 76976 83988 76982
rect 85952 77182 86164 77188
rect 85952 77118 85958 77182
rect 86022 77118 86164 77182
rect 85952 77047 86164 77118
rect 86360 77087 86436 77188
rect 85952 76991 86026 77047
rect 86082 76991 86164 77047
rect 83504 76840 83716 76916
rect 85952 76840 86164 76991
rect 86259 77046 86436 77087
rect 86259 76989 86366 77046
rect 86360 76982 86366 76989
rect 86430 76982 86436 77046
rect 86360 76976 86436 76982
rect 88400 77182 88612 77188
rect 88400 77118 88406 77182
rect 88470 77118 88612 77182
rect 88400 77047 88612 77118
rect 88808 77087 88884 77188
rect 88400 76991 88522 77047
rect 88578 76991 88612 77047
rect 88400 76840 88612 76991
rect 88755 77052 88884 77087
rect 90984 77182 91060 77188
rect 90984 77118 90990 77182
rect 91054 77118 91060 77182
rect 90984 77068 91060 77118
rect 91256 77182 91468 77188
rect 91256 77118 91262 77182
rect 91326 77118 91468 77182
rect 91256 77087 91468 77118
rect 88755 77046 89020 77052
rect 88755 76989 88950 77046
rect 88808 76982 88950 76989
rect 89014 76982 89020 77046
rect 88808 76976 89020 76982
rect 90984 77047 91095 77068
rect 90984 76991 91018 77047
rect 91074 76991 91095 77047
rect 90984 76916 91095 76991
rect 91251 76989 91468 77087
rect 91392 76976 91468 76989
rect 93432 77182 93644 77188
rect 93432 77118 93574 77182
rect 93638 77118 93644 77182
rect 93432 77047 93644 77118
rect 93840 77087 93916 77188
rect 93432 76991 93514 77047
rect 93570 76991 93644 77047
rect 90984 76840 91196 76916
rect 93432 76840 93644 76991
rect 93747 77046 93916 77087
rect 93747 76989 93846 77046
rect 93840 76982 93846 76989
rect 93910 76982 93916 77046
rect 93840 76976 93916 76982
rect 95880 77182 96092 77188
rect 95880 77118 96022 77182
rect 96086 77118 96092 77182
rect 95880 77047 96092 77118
rect 96288 77087 96364 77188
rect 95880 76991 96010 77047
rect 96066 76991 96092 77047
rect 95880 76840 96092 76991
rect 96243 77046 96364 77087
rect 96243 76989 96294 77046
rect 96288 76982 96294 76989
rect 96358 76982 96364 77046
rect 96288 76976 96364 76982
rect 98464 77182 98676 77188
rect 98464 77118 98470 77182
rect 98534 77118 98676 77182
rect 98464 77047 98676 77118
rect 98872 77087 98948 77188
rect 98464 76991 98506 77047
rect 98562 76991 98676 77047
rect 98464 76840 98676 76991
rect 98739 77046 98948 77087
rect 98739 76989 98878 77046
rect 98872 76982 98878 76989
rect 98942 76982 98948 77046
rect 98872 76976 98948 76982
rect 100912 77182 101124 77188
rect 100912 77118 101054 77182
rect 101118 77118 101124 77182
rect 100912 77047 101124 77118
rect 101320 77087 101396 77188
rect 100912 76991 101002 77047
rect 101058 76991 101124 77047
rect 100912 76840 101124 76991
rect 101235 77046 101396 77087
rect 101235 76989 101326 77046
rect 101320 76982 101326 76989
rect 101390 76982 101396 77046
rect 101320 76976 101396 76982
rect 103360 77182 103572 77188
rect 103360 77118 103366 77182
rect 103430 77118 103572 77182
rect 103768 77182 103980 77188
rect 103768 77150 103910 77182
rect 103360 77068 103572 77118
rect 103731 77118 103910 77150
rect 103974 77118 103980 77182
rect 103731 77112 103980 77118
rect 105944 77182 106156 77188
rect 105944 77118 106086 77182
rect 106150 77118 106156 77182
rect 103360 77047 103575 77068
rect 103360 76991 103498 77047
rect 103554 76991 103575 77047
rect 103360 76916 103575 76991
rect 103731 76989 103829 77112
rect 105944 77047 106156 77118
rect 106352 77087 106428 77188
rect 115328 77182 115540 77248
rect 115328 77118 115334 77182
rect 115398 77118 115540 77182
rect 115328 77112 115540 77118
rect 116416 77112 116628 77248
rect 105944 76991 105994 77047
rect 106050 76991 106156 77047
rect 103360 76840 103708 76916
rect 105944 76840 106156 76991
rect 106227 77046 106428 77087
rect 106227 76989 106358 77046
rect 106352 76982 106358 76989
rect 106422 76982 106428 77046
rect 106352 76976 106428 76982
rect 122264 77046 122476 77052
rect 122264 76982 122406 77046
rect 122470 76982 122476 77046
rect 122264 76910 122476 76982
rect 122264 76846 122406 76910
rect 122470 76846 122476 76910
rect 122264 76840 122476 76846
rect 28832 76638 29044 76780
rect 28832 76574 28974 76638
rect 29038 76574 29044 76638
rect 28832 76568 29044 76574
rect 31280 76704 36524 76780
rect 31280 76638 31492 76704
rect 31280 76574 31286 76638
rect 31350 76574 31492 76638
rect 31280 76568 31492 76574
rect 33728 76638 34076 76704
rect 33728 76574 33734 76638
rect 33798 76574 34076 76638
rect 33728 76568 34076 76574
rect 36312 76644 36524 76704
rect 36312 76638 38700 76644
rect 36312 76574 36318 76638
rect 36382 76574 38630 76638
rect 38694 76574 38700 76638
rect 36312 76568 38700 76574
rect 38760 76638 38972 76780
rect 38760 76574 38902 76638
rect 38966 76574 38972 76638
rect 38760 76568 38972 76574
rect 41208 76644 41556 76780
rect 41208 76638 43732 76644
rect 41208 76574 41350 76638
rect 41414 76574 43662 76638
rect 43726 76574 43732 76638
rect 41208 76568 43732 76574
rect 43792 76638 44004 76780
rect 43792 76574 43934 76638
rect 43998 76574 44004 76638
rect 43792 76568 44004 76574
rect 46240 76638 46452 76780
rect 46240 76574 46382 76638
rect 46446 76574 46452 76638
rect 46240 76568 46452 76574
rect 48688 76704 51484 76780
rect 48688 76638 49036 76704
rect 48688 76574 48694 76638
rect 48758 76574 49036 76638
rect 48688 76568 49036 76574
rect 51272 76638 51484 76704
rect 51272 76574 51414 76638
rect 51478 76574 51484 76638
rect 51272 76568 51484 76574
rect 53720 76644 53932 76780
rect 56304 76704 61412 76780
rect 53720 76638 56244 76644
rect 53720 76574 53726 76638
rect 53790 76574 56174 76638
rect 56238 76574 56244 76638
rect 53720 76568 56244 76574
rect 56304 76638 56516 76704
rect 56304 76574 56310 76638
rect 56374 76574 56516 76638
rect 56304 76568 56516 76574
rect 58752 76638 58964 76704
rect 58752 76574 58758 76638
rect 58822 76574 58964 76638
rect 58752 76568 58964 76574
rect 61200 76638 61412 76704
rect 61200 76574 61342 76638
rect 61406 76574 61412 76638
rect 61200 76568 61412 76574
rect 63784 76638 63996 76780
rect 63784 76574 63790 76638
rect 63854 76574 63996 76638
rect 63784 76568 63996 76574
rect 66232 76638 66444 76780
rect 66232 76574 66374 76638
rect 66438 76574 66444 76638
rect 66232 76568 66444 76574
rect 68680 76638 68892 76780
rect 71264 76644 71476 76780
rect 71166 76638 71476 76644
rect 68680 76574 68822 76638
rect 68886 76574 68892 76638
rect 71128 76574 71134 76638
rect 71198 76574 71406 76638
rect 71470 76574 71476 76638
rect 68680 76568 68892 76574
rect 71166 76568 71476 76574
rect 73712 76704 76508 76780
rect 73712 76638 73924 76704
rect 73712 76574 73718 76638
rect 73782 76574 73924 76638
rect 73712 76568 73924 76574
rect 76160 76644 76508 76704
rect 78744 76644 78956 76780
rect 81192 76644 81404 76780
rect 76160 76638 78684 76644
rect 76160 76574 76166 76638
rect 76230 76574 78614 76638
rect 78678 76574 78684 76638
rect 76160 76568 78684 76574
rect 78744 76638 81404 76644
rect 78744 76574 78750 76638
rect 78814 76574 81334 76638
rect 81398 76574 81404 76638
rect 78744 76568 81404 76574
rect 83640 76644 83988 76780
rect 86224 76644 86436 76780
rect 88672 76644 88884 76780
rect 83640 76638 86436 76644
rect 88574 76638 88884 76644
rect 83640 76574 83782 76638
rect 83846 76574 86366 76638
rect 86430 76574 86436 76638
rect 88536 76574 88542 76638
rect 88606 76574 88814 76638
rect 88878 76574 88884 76638
rect 83640 76568 86436 76574
rect 88574 76568 88884 76574
rect 91120 76644 91468 76780
rect 91120 76638 93644 76644
rect 91120 76574 91398 76638
rect 91462 76574 93574 76638
rect 93638 76574 93644 76638
rect 91120 76568 93644 76574
rect 93704 76638 93916 76780
rect 93704 76574 93846 76638
rect 93910 76574 93916 76638
rect 93704 76568 93916 76574
rect 96152 76644 96364 76780
rect 98736 76704 103844 76780
rect 96152 76638 98676 76644
rect 96152 76574 96158 76638
rect 96222 76574 98606 76638
rect 98670 76574 98676 76638
rect 96152 76568 98676 76574
rect 98736 76638 98948 76704
rect 98736 76574 98742 76638
rect 98806 76574 98948 76638
rect 98736 76568 98948 76574
rect 101184 76638 101396 76704
rect 101184 76574 101190 76638
rect 101254 76574 101396 76638
rect 101184 76568 101396 76574
rect 103632 76638 103844 76704
rect 103632 76574 103774 76638
rect 103838 76574 103844 76638
rect 103632 76568 103844 76574
rect 106216 76638 106428 76780
rect 106216 76574 106222 76638
rect 106286 76574 106428 76638
rect 106216 76568 106428 76574
rect 1224 76094 1980 76100
rect 1224 76030 1230 76094
rect 1294 76030 1980 76094
rect 1224 76024 1980 76030
rect 1768 76008 1980 76024
rect 1768 75952 1794 76008
rect 1850 75952 1980 76008
rect 134776 76094 135396 76100
rect 134776 76030 135326 76094
rect 135390 76030 135396 76094
rect 134776 76024 135396 76030
rect 134776 76008 134988 76024
rect 1768 75888 1980 75952
rect 28832 75958 31492 75964
rect 28832 75894 28974 75958
rect 29038 75894 31286 75958
rect 31350 75894 31492 75958
rect 28832 75888 31492 75894
rect 28832 75752 29044 75888
rect 31280 75752 31492 75888
rect 33728 75958 33940 75964
rect 33728 75894 33734 75958
rect 33798 75894 33940 75958
rect 33728 75752 33940 75894
rect 36312 75958 36524 75964
rect 38662 75958 38972 75964
rect 36312 75894 36318 75958
rect 36382 75894 36524 75958
rect 38624 75894 38630 75958
rect 38694 75894 38902 75958
rect 38966 75894 38972 75958
rect 36312 75752 36524 75894
rect 38662 75888 38972 75894
rect 38760 75828 38972 75888
rect 41208 75958 41420 75964
rect 43694 75958 49036 75964
rect 41208 75894 41350 75958
rect 41414 75894 41420 75958
rect 43656 75894 43662 75958
rect 43726 75894 43934 75958
rect 43998 75894 46382 75958
rect 46446 75894 48694 75958
rect 48758 75894 49036 75958
rect 41208 75828 41420 75894
rect 43694 75888 49036 75894
rect 38760 75752 41420 75828
rect 43792 75752 44004 75888
rect 46240 75752 46452 75888
rect 48688 75752 49036 75888
rect 51272 75958 51484 75964
rect 51272 75894 51414 75958
rect 51478 75894 51484 75958
rect 51272 75828 51484 75894
rect 53720 75958 53932 75964
rect 53720 75894 53726 75958
rect 53790 75894 53932 75958
rect 53720 75828 53932 75894
rect 51272 75752 53932 75828
rect 56168 75958 56516 75964
rect 56168 75894 56174 75958
rect 56238 75894 56310 75958
rect 56374 75894 56516 75958
rect 56168 75752 56516 75894
rect 58752 75958 58964 75964
rect 58752 75894 58758 75958
rect 58822 75894 58964 75958
rect 58752 75828 58964 75894
rect 61200 75958 66444 75964
rect 61200 75894 61342 75958
rect 61406 75894 63790 75958
rect 63854 75894 66374 75958
rect 66438 75894 66444 75958
rect 61200 75888 66444 75894
rect 58752 75822 59508 75828
rect 58752 75758 59438 75822
rect 59502 75758 59508 75822
rect 58752 75752 59508 75758
rect 61200 75752 61412 75888
rect 63648 75752 63996 75888
rect 66232 75828 66444 75888
rect 68680 75958 71204 75964
rect 68680 75894 68822 75958
rect 68886 75894 71134 75958
rect 71198 75894 71204 75958
rect 68680 75888 71204 75894
rect 71264 75958 73924 75964
rect 71264 75894 71406 75958
rect 71470 75894 73718 75958
rect 73782 75894 73924 75958
rect 71264 75888 73924 75894
rect 68680 75828 68892 75888
rect 66232 75752 68892 75828
rect 71264 75752 71476 75888
rect 73712 75752 73924 75888
rect 76160 75958 76372 75964
rect 78646 75958 78956 75964
rect 76160 75894 76166 75958
rect 76230 75894 76372 75958
rect 78608 75894 78614 75958
rect 78678 75894 78750 75958
rect 78814 75894 78956 75958
rect 76160 75752 76372 75894
rect 78646 75888 78956 75894
rect 78744 75752 78956 75888
rect 81192 75958 81404 75964
rect 81192 75894 81334 75958
rect 81398 75894 81404 75958
rect 81192 75828 81404 75894
rect 83640 75958 83852 75964
rect 83640 75894 83782 75958
rect 83846 75894 83852 75958
rect 83640 75828 83852 75894
rect 81192 75752 83852 75828
rect 86224 75958 88612 75964
rect 86224 75894 86366 75958
rect 86430 75894 88542 75958
rect 88606 75894 88612 75958
rect 86224 75888 88612 75894
rect 88672 75958 91468 75964
rect 93606 75958 93916 75964
rect 88672 75894 88814 75958
rect 88878 75894 91398 75958
rect 91462 75894 91468 75958
rect 93568 75894 93574 75958
rect 93638 75894 93846 75958
rect 93910 75894 93916 75958
rect 88672 75888 91468 75894
rect 93606 75888 93916 75894
rect 86224 75752 86436 75888
rect 88672 75752 88884 75888
rect 91120 75752 91468 75888
rect 93704 75828 93916 75888
rect 96152 75958 96364 75964
rect 96152 75894 96158 75958
rect 96222 75894 96364 75958
rect 96152 75828 96364 75894
rect 93704 75752 96364 75828
rect 98600 75958 98948 75964
rect 98600 75894 98606 75958
rect 98670 75894 98742 75958
rect 98806 75894 98948 75958
rect 98600 75752 98948 75894
rect 101184 75958 101396 75964
rect 101184 75894 101190 75958
rect 101254 75894 101396 75958
rect 101184 75752 101396 75894
rect 103632 75958 106428 75964
rect 103632 75894 103774 75958
rect 103838 75894 106222 75958
rect 106286 75894 106428 75958
rect 103632 75888 106428 75894
rect 103632 75752 103844 75888
rect 106080 75752 106428 75888
rect 115328 75692 115540 75964
rect 116416 75958 116628 75964
rect 116416 75894 116558 75958
rect 116622 75894 116628 75958
rect 116416 75692 116628 75894
rect 134776 75952 134844 76008
rect 134900 75952 134988 76008
rect 134776 75888 134988 75952
rect 115328 75686 116628 75692
rect 115328 75622 115470 75686
rect 115534 75622 116628 75686
rect 115328 75616 116628 75622
rect 122264 75686 122476 75692
rect 122264 75622 122270 75686
rect 122334 75622 122476 75686
rect 122264 75550 122476 75622
rect 122264 75486 122270 75550
rect 122334 75486 122476 75550
rect 122264 75480 122476 75486
rect 28832 75278 29044 75284
rect 28832 75214 28838 75278
rect 28902 75214 29044 75278
rect 28832 75142 29044 75214
rect 28832 75078 28974 75142
rect 29038 75078 29044 75142
rect 28832 75072 29044 75078
rect 31416 75278 31628 75284
rect 31416 75214 31422 75278
rect 31486 75214 31628 75278
rect 31416 75142 31628 75214
rect 31416 75078 31558 75142
rect 31622 75078 31628 75142
rect 31416 75072 31628 75078
rect 33864 75278 34076 75284
rect 33864 75214 34006 75278
rect 34070 75214 34076 75278
rect 33864 75142 34076 75214
rect 33864 75078 34006 75142
rect 34070 75078 34076 75142
rect 33864 75072 34076 75078
rect 36312 75278 36524 75284
rect 36312 75214 36454 75278
rect 36518 75214 36524 75278
rect 36312 75142 36524 75214
rect 36312 75078 36454 75142
rect 36518 75078 36524 75142
rect 36312 75072 36524 75078
rect 38896 75278 39108 75284
rect 38896 75214 39038 75278
rect 39102 75214 39108 75278
rect 38896 75142 39108 75214
rect 38896 75078 39038 75142
rect 39102 75078 39108 75142
rect 38896 75072 39108 75078
rect 41344 75278 41556 75284
rect 41344 75214 41486 75278
rect 41550 75214 41556 75278
rect 41344 75142 41556 75214
rect 41344 75078 41486 75142
rect 41550 75078 41556 75142
rect 41344 75072 41556 75078
rect 43792 75278 44004 75284
rect 43792 75214 43798 75278
rect 43862 75214 44004 75278
rect 43792 75148 44004 75214
rect 46376 75278 46588 75284
rect 46376 75214 46518 75278
rect 46582 75214 46588 75278
rect 43792 75142 44140 75148
rect 43792 75078 44070 75142
rect 44134 75078 44140 75142
rect 43792 75072 44140 75078
rect 46376 75142 46588 75214
rect 46376 75078 46518 75142
rect 46582 75078 46588 75142
rect 46376 75072 46588 75078
rect 48824 75278 49036 75284
rect 48824 75214 48966 75278
rect 49030 75214 49036 75278
rect 48824 75142 49036 75214
rect 48824 75078 48966 75142
rect 49030 75078 49036 75142
rect 48824 75072 49036 75078
rect 51272 75278 51484 75284
rect 51272 75214 51278 75278
rect 51342 75214 51484 75278
rect 51272 75148 51484 75214
rect 53856 75278 54068 75284
rect 53856 75214 53862 75278
rect 53926 75214 54068 75278
rect 51272 75142 51620 75148
rect 51272 75078 51550 75142
rect 51614 75078 51620 75142
rect 51272 75072 51620 75078
rect 53856 75142 54068 75214
rect 53856 75078 53998 75142
rect 54062 75078 54068 75142
rect 53856 75072 54068 75078
rect 56304 75278 56516 75284
rect 56304 75214 56446 75278
rect 56510 75214 56516 75278
rect 56304 75142 56516 75214
rect 56304 75078 56310 75142
rect 56374 75078 56516 75142
rect 56304 75072 56516 75078
rect 58752 75278 59100 75284
rect 58752 75214 58894 75278
rect 58958 75214 59100 75278
rect 58752 75142 59100 75214
rect 58752 75078 59030 75142
rect 59094 75078 59100 75142
rect 58752 75072 59100 75078
rect 61336 75278 61548 75284
rect 61336 75214 61478 75278
rect 61542 75214 61548 75278
rect 61336 75142 61548 75214
rect 61336 75078 61478 75142
rect 61542 75078 61548 75142
rect 61336 75072 61548 75078
rect 63784 75278 63996 75284
rect 63784 75214 63926 75278
rect 63990 75214 63996 75278
rect 63784 75142 63996 75214
rect 63784 75078 63926 75142
rect 63990 75078 63996 75142
rect 63784 75072 63996 75078
rect 66232 75278 66580 75284
rect 66232 75214 66510 75278
rect 66574 75214 66580 75278
rect 66232 75142 66580 75214
rect 66232 75078 66510 75142
rect 66574 75078 66580 75142
rect 66232 75072 66580 75078
rect 68816 75278 69028 75284
rect 68816 75214 68958 75278
rect 69022 75214 69028 75278
rect 68816 75142 69028 75214
rect 68816 75078 68958 75142
rect 69022 75078 69028 75142
rect 68816 75072 69028 75078
rect 71264 75278 71476 75284
rect 71264 75214 71270 75278
rect 71334 75214 71476 75278
rect 71264 75142 71476 75214
rect 71264 75078 71406 75142
rect 71470 75078 71476 75142
rect 71264 75072 71476 75078
rect 73848 75278 74060 75284
rect 73848 75214 73854 75278
rect 73918 75214 74060 75278
rect 73848 75142 74060 75214
rect 73848 75078 73990 75142
rect 74054 75078 74060 75142
rect 73848 75072 74060 75078
rect 76296 75278 76508 75284
rect 76296 75214 76438 75278
rect 76502 75214 76508 75278
rect 76296 75142 76508 75214
rect 76296 75078 76438 75142
rect 76502 75078 76508 75142
rect 76296 75072 76508 75078
rect 78744 75278 78956 75284
rect 78744 75214 78886 75278
rect 78950 75214 78956 75278
rect 78744 75142 78956 75214
rect 78744 75078 78886 75142
rect 78950 75078 78956 75142
rect 78744 75072 78956 75078
rect 81328 75278 81540 75284
rect 81328 75214 81470 75278
rect 81534 75214 81540 75278
rect 81328 75142 81540 75214
rect 81328 75078 81470 75142
rect 81534 75078 81540 75142
rect 81328 75072 81540 75078
rect 83776 75278 83988 75284
rect 83776 75214 83918 75278
rect 83982 75214 83988 75278
rect 83776 75142 83988 75214
rect 83776 75078 83918 75142
rect 83982 75078 83988 75142
rect 83776 75072 83988 75078
rect 86224 75278 86436 75284
rect 86224 75214 86230 75278
rect 86294 75214 86436 75278
rect 86224 75148 86436 75214
rect 88808 75278 89020 75284
rect 88808 75214 88950 75278
rect 89014 75214 89020 75278
rect 86224 75142 86572 75148
rect 86224 75078 86502 75142
rect 86566 75078 86572 75142
rect 86224 75072 86572 75078
rect 88808 75142 89020 75214
rect 88808 75078 88950 75142
rect 89014 75078 89020 75142
rect 88808 75072 89020 75078
rect 91256 75278 91468 75284
rect 91256 75214 91262 75278
rect 91326 75214 91468 75278
rect 91256 75142 91468 75214
rect 91256 75078 91398 75142
rect 91462 75078 91468 75142
rect 91256 75072 91468 75078
rect 93704 75278 93916 75284
rect 93704 75214 93710 75278
rect 93774 75214 93916 75278
rect 93704 75142 93916 75214
rect 93704 75078 93710 75142
rect 93774 75078 93916 75142
rect 93704 75072 93916 75078
rect 96288 75278 96500 75284
rect 96288 75214 96294 75278
rect 96358 75214 96500 75278
rect 96288 75142 96500 75214
rect 96288 75078 96430 75142
rect 96494 75078 96500 75142
rect 96288 75072 96500 75078
rect 98736 75278 98948 75284
rect 98736 75214 98878 75278
rect 98942 75214 98948 75278
rect 98736 75142 98948 75214
rect 98736 75078 98878 75142
rect 98942 75078 98948 75142
rect 98736 75072 98948 75078
rect 101184 75278 101532 75284
rect 101184 75214 101326 75278
rect 101390 75214 101532 75278
rect 101184 75142 101532 75214
rect 101184 75078 101462 75142
rect 101526 75078 101532 75142
rect 101184 75072 101532 75078
rect 103768 75278 103980 75284
rect 103768 75214 103910 75278
rect 103974 75214 103980 75278
rect 103768 75142 103980 75214
rect 103768 75078 103910 75142
rect 103974 75078 103980 75142
rect 103768 75072 103980 75078
rect 106216 75278 106428 75284
rect 106216 75214 106358 75278
rect 106422 75214 106428 75278
rect 106216 75142 106428 75214
rect 106216 75078 106358 75142
rect 106422 75078 106428 75142
rect 106216 75072 106428 75078
rect 28921 75055 29019 75072
rect 31417 75055 31515 75072
rect 33913 75055 34011 75072
rect 36409 75055 36507 75072
rect 38905 75055 39003 75072
rect 41401 75055 41499 75072
rect 43897 75055 43995 75072
rect 46393 75055 46491 75072
rect 48889 75055 48987 75072
rect 51385 75055 51483 75072
rect 53881 75055 53979 75072
rect 56377 75055 56475 75072
rect 58873 75055 58971 75072
rect 61369 75055 61467 75072
rect 63865 75055 63963 75072
rect 66361 75055 66459 75072
rect 68857 75055 68955 75072
rect 71353 75055 71451 75072
rect 73849 75055 73947 75072
rect 76345 75055 76443 75072
rect 78841 75055 78939 75072
rect 81337 75055 81435 75072
rect 83833 75055 83931 75072
rect 86329 75055 86427 75072
rect 88825 75055 88923 75072
rect 91321 75055 91419 75072
rect 93817 75055 93915 75072
rect 96313 75055 96411 75072
rect 98809 75055 98907 75072
rect 101305 75055 101403 75072
rect 103801 75055 103899 75072
rect 106297 75055 106395 75072
rect 110056 74885 110122 74919
rect 122267 74885 122333 74888
rect 110056 74883 122333 74885
rect 110056 74827 110061 74883
rect 110117 74827 122272 74883
rect 122328 74827 122333 74883
rect 110056 74825 122333 74827
rect 110056 74822 110122 74825
rect 122267 74822 122333 74825
rect 1768 74328 1980 74468
rect 1768 74272 1794 74328
rect 1850 74272 1980 74328
rect 1768 74196 1980 74272
rect 115328 74462 116628 74468
rect 115328 74398 115334 74462
rect 115398 74398 116628 74462
rect 115328 74392 116628 74398
rect 115328 74326 115540 74392
rect 115328 74262 115334 74326
rect 115398 74262 115540 74326
rect 115328 74256 115540 74262
rect 116416 74256 116628 74392
rect 122264 74326 122476 74332
rect 122264 74262 122406 74326
rect 122470 74262 122476 74326
rect 1224 74190 1980 74196
rect 1224 74126 1230 74190
rect 1294 74126 1980 74190
rect 1224 74120 1980 74126
rect 122264 74054 122476 74262
rect 122264 73990 122406 74054
rect 122470 73990 122476 74054
rect 122264 73984 122476 73990
rect 132600 74060 132812 74332
rect 133280 74196 133492 74332
rect 134776 74328 134988 74468
rect 134776 74272 134844 74328
rect 134900 74272 134988 74328
rect 134776 74196 134988 74272
rect 133280 74190 135396 74196
rect 133280 74126 135326 74190
rect 135390 74126 135396 74190
rect 133280 74120 135396 74126
rect 133280 74060 133492 74120
rect 132600 73984 133492 74060
rect 110180 73471 110246 73474
rect 122267 73471 122333 73474
rect 110180 73469 122333 73471
rect 110180 73413 110185 73469
rect 110241 73413 122272 73469
rect 122328 73413 122333 73469
rect 110180 73411 122333 73413
rect 110180 73408 110246 73411
rect 122267 73408 122333 73411
rect 28968 73238 29316 73244
rect 28968 73174 28974 73238
rect 29038 73174 29316 73238
rect 28968 73108 29316 73174
rect 30328 73108 30540 73244
rect 31552 73238 32988 73244
rect 31552 73174 31558 73238
rect 31622 73174 32988 73238
rect 31552 73168 32988 73174
rect 31552 73108 31764 73168
rect 28968 73102 31764 73108
rect 28968 73038 28974 73102
rect 29038 73038 31764 73102
rect 28968 73032 31764 73038
rect 32776 73108 32988 73168
rect 34000 73238 35436 73244
rect 34000 73174 34006 73238
rect 34070 73174 35436 73238
rect 34000 73168 35436 73174
rect 34000 73108 34212 73168
rect 32776 73032 34212 73108
rect 35224 73108 35436 73168
rect 36448 73238 39244 73244
rect 36448 73174 36454 73238
rect 36518 73174 39038 73238
rect 39102 73174 39244 73238
rect 36448 73168 39244 73174
rect 36448 73108 36796 73168
rect 35224 73032 36796 73108
rect 37808 73032 38020 73168
rect 39032 73108 39244 73168
rect 40256 73238 41692 73244
rect 40256 73174 41486 73238
rect 41550 73174 41692 73238
rect 40256 73168 41692 73174
rect 40256 73108 40468 73168
rect 39032 73032 40468 73108
rect 41480 73108 41692 73168
rect 42704 73238 45500 73244
rect 42704 73174 44070 73238
rect 44134 73174 45500 73238
rect 42704 73168 45500 73174
rect 42704 73108 43052 73168
rect 41480 73032 43052 73108
rect 44064 73032 44276 73168
rect 45288 73108 45500 73168
rect 46512 73238 47948 73244
rect 46512 73174 46518 73238
rect 46582 73174 47948 73238
rect 46512 73168 47948 73174
rect 46512 73108 46724 73168
rect 45288 73032 46724 73108
rect 47736 73108 47948 73168
rect 48960 73238 51756 73244
rect 48960 73174 48966 73238
rect 49030 73174 51550 73238
rect 51614 73174 51756 73238
rect 48960 73168 51756 73174
rect 48960 73108 49172 73168
rect 47736 73032 49172 73108
rect 50184 73032 50532 73168
rect 51544 73108 51756 73168
rect 52768 73238 54204 73244
rect 52768 73174 53998 73238
rect 54062 73174 54204 73238
rect 52768 73168 54204 73174
rect 52768 73108 52980 73168
rect 51544 73032 52980 73108
rect 53992 73108 54204 73168
rect 55216 73238 56380 73244
rect 55216 73174 56310 73238
rect 56374 73174 56380 73238
rect 55216 73168 56380 73174
rect 55216 73108 55428 73168
rect 56440 73108 56652 73244
rect 57664 73238 60460 73244
rect 57664 73174 59030 73238
rect 59094 73174 60460 73238
rect 57664 73168 60460 73174
rect 57664 73108 58012 73168
rect 53992 73032 58012 73108
rect 59024 73032 59236 73168
rect 60248 73108 60460 73168
rect 61472 73238 62908 73244
rect 61472 73174 61478 73238
rect 61542 73174 62908 73238
rect 61472 73168 62908 73174
rect 61472 73108 61684 73168
rect 60248 73032 61684 73108
rect 62696 73108 62908 73168
rect 63920 73238 66716 73244
rect 63920 73174 63926 73238
rect 63990 73174 66510 73238
rect 66574 73174 66716 73238
rect 63920 73168 66716 73174
rect 63920 73108 64268 73168
rect 62696 73032 64268 73108
rect 65280 73032 65492 73168
rect 66504 73108 66716 73168
rect 67728 73238 69164 73244
rect 67728 73174 68958 73238
rect 69022 73174 69164 73238
rect 67728 73168 69164 73174
rect 67728 73108 67940 73168
rect 66504 73032 67940 73108
rect 68952 73108 69164 73168
rect 70176 73238 71748 73244
rect 70176 73174 71406 73238
rect 71470 73174 71748 73238
rect 70176 73168 71748 73174
rect 70176 73108 70388 73168
rect 68952 73032 70388 73108
rect 71400 73108 71748 73168
rect 72760 73108 72972 73244
rect 73984 73238 75420 73244
rect 73984 73174 73990 73238
rect 74054 73174 75420 73238
rect 73984 73168 75420 73174
rect 73984 73108 74196 73168
rect 71400 73032 74196 73108
rect 75208 73108 75420 73168
rect 76432 73238 77868 73244
rect 76432 73174 76438 73238
rect 76502 73174 77868 73238
rect 76432 73168 77868 73174
rect 76432 73108 76644 73168
rect 75208 73032 76644 73108
rect 77656 73108 77868 73168
rect 78880 73238 81676 73244
rect 78880 73174 78886 73238
rect 78950 73174 81470 73238
rect 81534 73174 81676 73238
rect 78880 73168 81676 73174
rect 78880 73108 79228 73168
rect 77656 73032 79228 73108
rect 80240 73032 80452 73168
rect 81464 73108 81676 73168
rect 82688 73238 84124 73244
rect 82688 73174 83918 73238
rect 83982 73174 84124 73238
rect 82688 73168 84124 73174
rect 82688 73108 82900 73168
rect 81464 73032 82900 73108
rect 83912 73108 84124 73168
rect 85136 73238 87932 73244
rect 85136 73174 86502 73238
rect 86566 73174 87932 73238
rect 85136 73168 87932 73174
rect 85136 73108 85484 73168
rect 83912 73032 85484 73108
rect 86496 73032 86708 73168
rect 87720 73108 87932 73168
rect 88944 73238 90380 73244
rect 88944 73174 88950 73238
rect 89014 73174 90380 73238
rect 88944 73168 90380 73174
rect 88944 73108 89156 73168
rect 87720 73032 89156 73108
rect 90168 73108 90380 73168
rect 91392 73238 93780 73244
rect 91392 73174 91398 73238
rect 91462 73174 93710 73238
rect 93774 73174 93780 73238
rect 91392 73168 93780 73174
rect 91392 73108 91604 73168
rect 90168 73032 91604 73108
rect 92616 73108 92964 73168
rect 93976 73108 94188 73244
rect 95200 73238 96636 73244
rect 95200 73174 96430 73238
rect 96494 73174 96636 73238
rect 95200 73168 96636 73174
rect 95200 73108 95412 73168
rect 92616 73032 95412 73108
rect 96424 73108 96636 73168
rect 97648 73238 99084 73244
rect 97648 73174 98878 73238
rect 98942 73174 99084 73238
rect 97648 73168 99084 73174
rect 97648 73108 97860 73168
rect 96424 73032 97860 73108
rect 98872 73108 99084 73168
rect 100096 73108 100444 73244
rect 101456 73238 102892 73244
rect 101456 73174 101462 73238
rect 101526 73174 102892 73238
rect 101456 73168 102892 73174
rect 101456 73108 101668 73168
rect 98872 73032 101668 73108
rect 102680 73108 102892 73168
rect 103904 73238 105340 73244
rect 103904 73174 103910 73238
rect 103974 73174 105340 73238
rect 103904 73168 105340 73174
rect 103904 73108 104116 73168
rect 102680 73032 104116 73108
rect 105128 73108 105340 73168
rect 106352 73238 107924 73244
rect 106352 73174 106358 73238
rect 106422 73174 107924 73238
rect 106352 73168 107924 73174
rect 106352 73108 106700 73168
rect 105128 73032 106700 73108
rect 107712 73108 107924 73168
rect 107712 73102 109692 73108
rect 107712 73038 109622 73102
rect 109686 73038 109692 73102
rect 107712 73032 109692 73038
rect 115328 73102 116628 73108
rect 115328 73038 115470 73102
rect 115534 73038 116628 73102
rect 115328 73032 116628 73038
rect 115328 72972 115540 73032
rect 115328 72966 115948 72972
rect 115328 72902 115878 72966
rect 115942 72902 115948 72966
rect 115328 72896 115948 72902
rect 116416 72896 116628 73032
rect 122264 72830 122476 72836
rect 122264 72766 122270 72830
rect 122334 72766 122476 72830
rect 1224 72694 1980 72700
rect 1224 72630 1230 72694
rect 1294 72648 1980 72694
rect 1294 72630 1794 72648
rect 1224 72624 1794 72630
rect 1768 72592 1794 72624
rect 1850 72592 1980 72648
rect 122264 72624 122476 72766
rect 132600 72830 136076 72836
rect 132600 72766 136006 72830
rect 136070 72766 136076 72830
rect 132600 72760 136076 72766
rect 132600 72624 132812 72760
rect 133280 72624 133492 72760
rect 134776 72648 134988 72700
rect 1768 72488 1980 72592
rect 134776 72592 134844 72648
rect 134900 72592 134988 72648
rect 134776 72564 134988 72592
rect 134776 72558 135396 72564
rect 134776 72494 135326 72558
rect 135390 72494 135396 72558
rect 134776 72488 135396 72494
rect 134087 72356 134093 72358
rect 115272 72296 115332 72356
rect 122132 72296 134093 72356
rect 134087 72294 134093 72296
rect 134157 72294 134163 72358
rect 114041 72057 114107 72060
rect 122267 72057 122333 72060
rect 114041 72055 122333 72057
rect 114041 71999 114046 72055
rect 114102 71999 122272 72055
rect 122328 71999 122333 72055
rect 114041 71997 122333 71999
rect 114041 71994 114107 71997
rect 122267 71994 122333 71997
rect 28560 71470 28772 71612
rect 28560 71406 28566 71470
rect 28630 71406 28702 71470
rect 28766 71406 28772 71470
rect 28560 71400 28772 71406
rect 29512 71476 29724 71612
rect 29784 71476 30132 71612
rect 29512 71470 30132 71476
rect 29512 71406 29790 71470
rect 29854 71406 30132 71470
rect 29512 71400 30132 71406
rect 30736 71536 31356 71612
rect 30736 71400 30948 71536
rect 31144 71470 31356 71536
rect 31144 71406 31286 71470
rect 31350 71406 31356 71470
rect 31144 71400 31356 71406
rect 31960 71476 32172 71612
rect 32368 71476 32580 71612
rect 31960 71470 32580 71476
rect 31960 71406 31966 71470
rect 32030 71406 32510 71470
rect 32574 71406 32580 71470
rect 31960 71400 32580 71406
rect 33184 71536 33804 71612
rect 33184 71400 33396 71536
rect 33592 71470 33804 71536
rect 33592 71406 33734 71470
rect 33798 71406 33804 71470
rect 33592 71400 33804 71406
rect 34408 71476 34620 71612
rect 34816 71476 35028 71612
rect 34408 71470 35028 71476
rect 34408 71406 34414 71470
rect 34478 71406 34958 71470
rect 35022 71406 35028 71470
rect 34408 71400 35028 71406
rect 35632 71476 35980 71612
rect 36040 71476 36252 71612
rect 35632 71470 36252 71476
rect 35632 71406 35774 71470
rect 35838 71406 36182 71470
rect 36246 71406 36252 71470
rect 35632 71400 36252 71406
rect 36992 71536 37612 71612
rect 36992 71470 37204 71536
rect 36992 71406 36998 71470
rect 37062 71406 37204 71470
rect 36992 71400 37204 71406
rect 37264 71470 37612 71536
rect 37264 71406 37542 71470
rect 37606 71406 37612 71470
rect 37264 71400 37612 71406
rect 38216 71476 38428 71612
rect 38624 71476 38836 71612
rect 38216 71470 38836 71476
rect 38216 71406 38222 71470
rect 38286 71406 38836 71470
rect 38216 71400 38836 71406
rect 39440 71536 40060 71612
rect 39440 71400 39652 71536
rect 39848 71470 40060 71536
rect 39848 71406 39990 71470
rect 40054 71406 40060 71470
rect 39848 71400 40060 71406
rect 40664 71476 40876 71612
rect 41072 71476 41284 71612
rect 40664 71470 41284 71476
rect 40664 71406 40670 71470
rect 40734 71406 41214 71470
rect 41278 71406 41284 71470
rect 40664 71400 41284 71406
rect 41888 71536 42508 71612
rect 41888 71470 42236 71536
rect 41888 71406 41894 71470
rect 41958 71406 42236 71470
rect 41888 71400 42236 71406
rect 42296 71470 42508 71536
rect 42296 71406 42438 71470
rect 42502 71406 42508 71470
rect 42296 71400 42508 71406
rect 43248 71536 43868 71612
rect 43248 71470 43460 71536
rect 43248 71406 43254 71470
rect 43318 71406 43460 71470
rect 43248 71400 43460 71406
rect 43520 71400 43868 71536
rect 44472 71476 44684 71612
rect 44880 71536 46316 71612
rect 44880 71476 45092 71536
rect 44472 71470 45092 71476
rect 44472 71406 44614 71470
rect 44678 71406 45092 71470
rect 44472 71400 45092 71406
rect 45696 71470 45908 71536
rect 45696 71406 45702 71470
rect 45766 71406 45908 71470
rect 45696 71400 45908 71406
rect 46104 71470 46316 71536
rect 46104 71406 46246 71470
rect 46310 71406 46316 71470
rect 46104 71400 46316 71406
rect 46920 71476 47132 71612
rect 47328 71476 47540 71612
rect 46920 71470 47540 71476
rect 46920 71406 46926 71470
rect 46990 71406 47540 71470
rect 46920 71400 47540 71406
rect 48144 71536 48764 71612
rect 48144 71400 48356 71536
rect 48552 71470 48764 71536
rect 48552 71406 48694 71470
rect 48758 71406 48764 71470
rect 48552 71400 48764 71406
rect 49368 71536 49988 71612
rect 49368 71400 49716 71536
rect 49776 71470 49988 71536
rect 49776 71406 49918 71470
rect 49982 71406 49988 71470
rect 49776 71400 49988 71406
rect 50728 71476 50940 71612
rect 51000 71476 51348 71612
rect 50728 71470 51348 71476
rect 50728 71406 50734 71470
rect 50798 71406 51278 71470
rect 51342 71406 51348 71470
rect 50728 71400 51348 71406
rect 51952 71536 52572 71612
rect 51952 71400 52164 71536
rect 52360 71470 52572 71536
rect 52360 71406 52502 71470
rect 52566 71406 52572 71470
rect 52360 71400 52572 71406
rect 53176 71476 53388 71612
rect 53584 71476 53796 71612
rect 53176 71470 53796 71476
rect 53176 71406 53182 71470
rect 53246 71406 53318 71470
rect 53382 71406 53796 71470
rect 53176 71400 53796 71406
rect 54400 71536 55020 71612
rect 54400 71470 54612 71536
rect 54400 71406 54406 71470
rect 54470 71406 54612 71470
rect 54400 71400 54612 71406
rect 54808 71470 55020 71536
rect 54808 71406 54950 71470
rect 55014 71406 55020 71470
rect 54808 71400 55020 71406
rect 55624 71476 55836 71612
rect 56032 71476 56244 71612
rect 55624 71470 56244 71476
rect 55624 71406 56038 71470
rect 56102 71406 56244 71470
rect 55624 71400 56244 71406
rect 56848 71536 57468 71612
rect 56848 71400 57196 71536
rect 57256 71470 57468 71536
rect 57256 71406 57398 71470
rect 57462 71406 57468 71470
rect 57256 71400 57468 71406
rect 58208 71536 58828 71612
rect 58208 71400 58420 71536
rect 58480 71470 58828 71536
rect 58480 71406 58622 71470
rect 58686 71406 58828 71470
rect 58480 71400 58828 71406
rect 59432 71606 59644 71612
rect 59432 71542 59438 71606
rect 59502 71542 59644 71606
rect 59432 71476 59644 71542
rect 59840 71476 60052 71612
rect 59432 71470 60052 71476
rect 59432 71406 59438 71470
rect 59502 71406 59982 71470
rect 60046 71406 60052 71470
rect 59432 71400 60052 71406
rect 60656 71536 61276 71612
rect 60656 71400 60868 71536
rect 61064 71470 61276 71536
rect 61064 71406 61206 71470
rect 61270 71406 61276 71470
rect 61064 71400 61276 71406
rect 61880 71476 62092 71612
rect 62288 71476 62500 71612
rect 61880 71470 62500 71476
rect 61880 71406 61886 71470
rect 61950 71406 62430 71470
rect 62494 71406 62500 71470
rect 61880 71400 62500 71406
rect 63104 71536 63724 71612
rect 63104 71470 63452 71536
rect 63104 71406 63110 71470
rect 63174 71406 63452 71470
rect 63104 71400 63452 71406
rect 63512 71470 63724 71536
rect 63512 71406 63654 71470
rect 63718 71406 63724 71470
rect 63512 71400 63724 71406
rect 64464 71536 65084 71612
rect 64464 71400 64676 71536
rect 64736 71470 65084 71536
rect 64736 71406 65014 71470
rect 65078 71406 65084 71470
rect 64736 71400 65084 71406
rect 65688 71476 65900 71612
rect 66096 71476 66308 71612
rect 65688 71470 66308 71476
rect 65688 71406 66102 71470
rect 66166 71406 66308 71470
rect 65688 71400 66308 71406
rect 66912 71536 67532 71612
rect 66912 71470 67124 71536
rect 66912 71406 66918 71470
rect 66982 71406 67124 71470
rect 66912 71400 67124 71406
rect 67320 71470 67532 71536
rect 67320 71406 67462 71470
rect 67526 71406 67532 71470
rect 67320 71400 67532 71406
rect 68136 71476 68348 71612
rect 68544 71476 68756 71612
rect 68136 71470 68756 71476
rect 68136 71406 68142 71470
rect 68206 71406 68686 71470
rect 68750 71406 68756 71470
rect 68136 71400 68756 71406
rect 69360 71536 69980 71612
rect 69360 71400 69572 71536
rect 69768 71470 69980 71536
rect 69768 71406 69910 71470
rect 69974 71406 69980 71470
rect 69768 71400 69980 71406
rect 70584 71476 70932 71612
rect 70992 71476 71204 71612
rect 70584 71470 71204 71476
rect 70584 71406 70590 71470
rect 70654 71406 71204 71470
rect 70584 71400 71204 71406
rect 71944 71476 72156 71612
rect 72216 71476 72564 71612
rect 71944 71470 72564 71476
rect 71944 71406 72086 71470
rect 72150 71406 72222 71470
rect 72286 71406 72564 71470
rect 71944 71400 72564 71406
rect 73168 71536 73788 71612
rect 73168 71400 73380 71536
rect 73576 71470 73788 71536
rect 73576 71406 73718 71470
rect 73782 71406 73788 71470
rect 73576 71400 73788 71406
rect 74392 71476 74604 71612
rect 74800 71476 75012 71612
rect 74392 71470 75012 71476
rect 74392 71406 74398 71470
rect 74462 71406 74942 71470
rect 75006 71406 75012 71470
rect 74392 71400 75012 71406
rect 75616 71536 76236 71612
rect 75616 71470 75828 71536
rect 75616 71406 75622 71470
rect 75686 71406 75828 71470
rect 75616 71400 75828 71406
rect 76024 71470 76236 71536
rect 76024 71406 76166 71470
rect 76230 71406 76236 71470
rect 76024 71400 76236 71406
rect 76840 71476 77052 71612
rect 77248 71476 77460 71612
rect 76840 71470 77460 71476
rect 76840 71406 76846 71470
rect 76910 71406 77390 71470
rect 77454 71406 77460 71470
rect 76840 71400 77460 71406
rect 78064 71470 78412 71612
rect 78064 71406 78206 71470
rect 78270 71406 78412 71470
rect 78064 71400 78412 71406
rect 78472 71470 78684 71612
rect 78472 71406 78478 71470
rect 78542 71406 78684 71470
rect 78472 71400 78684 71406
rect 79424 71536 80044 71612
rect 79424 71470 79636 71536
rect 79424 71406 79430 71470
rect 79494 71406 79636 71470
rect 79424 71400 79636 71406
rect 79696 71470 80044 71536
rect 79696 71406 79974 71470
rect 80038 71406 80044 71470
rect 79696 71400 80044 71406
rect 80648 71476 80860 71612
rect 81056 71476 81268 71612
rect 80648 71470 81268 71476
rect 80648 71406 80654 71470
rect 80718 71406 81268 71470
rect 80648 71400 81268 71406
rect 81872 71536 82492 71612
rect 81872 71470 82084 71536
rect 81872 71406 81878 71470
rect 81942 71406 82084 71470
rect 81872 71400 82084 71406
rect 82280 71470 82492 71536
rect 82280 71406 82422 71470
rect 82486 71406 82492 71470
rect 82280 71400 82492 71406
rect 83096 71476 83308 71612
rect 83504 71476 83716 71612
rect 83096 71470 83716 71476
rect 83096 71406 83102 71470
rect 83166 71406 83646 71470
rect 83710 71406 83716 71470
rect 83096 71400 83716 71406
rect 84320 71536 84940 71612
rect 84320 71470 84668 71536
rect 84320 71406 84598 71470
rect 84662 71406 84668 71470
rect 84320 71400 84668 71406
rect 84728 71400 84940 71536
rect 85680 71536 86300 71612
rect 85680 71400 85892 71536
rect 85952 71470 86300 71536
rect 85952 71406 86094 71470
rect 86158 71406 86300 71470
rect 85952 71400 86300 71406
rect 86904 71476 87116 71612
rect 87312 71476 87524 71612
rect 86904 71470 87524 71476
rect 86904 71406 86910 71470
rect 86974 71406 87524 71470
rect 86904 71400 87524 71406
rect 88128 71536 88748 71612
rect 88128 71470 88340 71536
rect 88128 71406 88134 71470
rect 88198 71406 88340 71470
rect 88128 71400 88340 71406
rect 88536 71470 88748 71536
rect 88536 71406 88678 71470
rect 88742 71406 88748 71470
rect 88536 71400 88748 71406
rect 89352 71476 89564 71612
rect 89760 71476 89972 71612
rect 89352 71470 89972 71476
rect 89352 71406 89358 71470
rect 89422 71406 89902 71470
rect 89966 71406 89972 71470
rect 89352 71400 89972 71406
rect 90576 71536 91196 71612
rect 90576 71470 90788 71536
rect 90576 71406 90718 71470
rect 90782 71406 90788 71470
rect 90576 71400 90788 71406
rect 90984 71470 91196 71536
rect 90984 71406 91126 71470
rect 91190 71406 91196 71470
rect 90984 71400 91196 71406
rect 91800 71476 92148 71612
rect 92208 71476 92420 71612
rect 91800 71470 92420 71476
rect 91800 71406 92350 71470
rect 92414 71406 92420 71470
rect 91800 71400 92420 71406
rect 93160 71476 93372 71612
rect 93432 71476 93780 71612
rect 93160 71470 93780 71476
rect 93160 71406 93302 71470
rect 93366 71406 93780 71470
rect 93160 71400 93780 71406
rect 94384 71536 95004 71612
rect 94384 71400 94596 71536
rect 94792 71470 95004 71536
rect 94792 71406 94934 71470
rect 94998 71406 95004 71470
rect 94792 71400 95004 71406
rect 95608 71476 95820 71612
rect 96016 71476 96228 71612
rect 95608 71470 96228 71476
rect 95608 71406 95614 71470
rect 95678 71406 96228 71470
rect 95608 71400 96228 71406
rect 96832 71536 97452 71612
rect 96832 71470 97044 71536
rect 96832 71406 96838 71470
rect 96902 71406 97044 71470
rect 96832 71400 97044 71406
rect 97240 71470 97452 71536
rect 97240 71406 97382 71470
rect 97446 71406 97452 71470
rect 97240 71400 97452 71406
rect 98056 71476 98268 71612
rect 98464 71476 98676 71612
rect 98056 71400 98676 71476
rect 99280 71536 99900 71612
rect 99280 71400 99628 71536
rect 99688 71470 99900 71536
rect 99688 71406 99830 71470
rect 99894 71406 99900 71470
rect 99688 71400 99900 71406
rect 100640 71536 101260 71612
rect 100640 71400 100852 71536
rect 100912 71470 101260 71536
rect 100912 71406 100918 71470
rect 100982 71406 101260 71470
rect 100912 71400 101260 71406
rect 101864 71476 102076 71612
rect 102272 71476 102484 71612
rect 101864 71470 102484 71476
rect 101864 71406 101870 71470
rect 101934 71406 102414 71470
rect 102478 71406 102484 71470
rect 101864 71400 102484 71406
rect 103088 71536 103708 71612
rect 103088 71470 103300 71536
rect 103088 71406 103094 71470
rect 103158 71406 103300 71470
rect 103088 71400 103300 71406
rect 103496 71470 103708 71536
rect 103496 71406 103638 71470
rect 103702 71406 103708 71470
rect 103496 71400 103708 71406
rect 104312 71476 104524 71612
rect 104720 71476 104932 71612
rect 104312 71470 104932 71476
rect 104312 71406 104318 71470
rect 104382 71406 104862 71470
rect 104926 71406 104932 71470
rect 104312 71400 104932 71406
rect 105536 71536 106156 71612
rect 105536 71470 105884 71536
rect 105536 71406 105542 71470
rect 105606 71406 105884 71470
rect 105536 71400 105884 71406
rect 105944 71470 106156 71536
rect 105944 71406 106086 71470
rect 106150 71406 106156 71470
rect 105944 71400 106156 71406
rect 106896 71536 107516 71612
rect 106896 71400 107108 71536
rect 107168 71470 107516 71536
rect 107168 71406 107310 71470
rect 107374 71406 107516 71470
rect 107168 71400 107516 71406
rect 108120 71476 108332 71612
rect 108528 71476 108740 71612
rect 108120 71470 108740 71476
rect 108120 71406 108534 71470
rect 108598 71406 108740 71470
rect 108120 71400 108740 71406
rect 122264 71470 122476 71476
rect 122264 71406 122406 71470
rect 122470 71406 122476 71470
rect 98192 71340 98268 71400
rect 98192 71334 98676 71340
rect 98192 71270 98606 71334
rect 98670 71270 98676 71334
rect 98192 71264 98676 71270
rect 122264 71264 122476 71406
rect 132600 71340 132812 71476
rect 133280 71340 133492 71476
rect 132600 71334 134852 71340
rect 132600 71270 134782 71334
rect 134846 71270 134852 71334
rect 132600 71264 134852 71270
rect 1224 71062 1980 71068
rect 1224 70998 1230 71062
rect 1294 70998 1980 71062
rect 1224 70992 1980 70998
rect 1768 70968 1980 70992
rect 1768 70912 1794 70968
rect 1850 70912 1980 70968
rect 28152 71062 28636 71068
rect 28152 70998 28566 71062
rect 28630 70998 28636 71062
rect 28152 70992 28636 70998
rect 28696 71062 28908 71068
rect 28696 70998 28702 71062
rect 28766 70998 28908 71062
rect 1768 70856 1980 70912
rect 27064 70796 27276 70932
rect 28152 70856 28364 70992
rect 28696 70932 28908 70998
rect 29376 71062 29860 71068
rect 29376 70998 29790 71062
rect 29854 70998 29860 71062
rect 29376 70992 29860 70998
rect 29920 70992 30812 71068
rect 29376 70932 29588 70992
rect 29920 70932 30132 70992
rect 28696 70856 30132 70932
rect 30600 70932 30812 70992
rect 31144 71062 31492 71068
rect 31144 70998 31286 71062
rect 31350 70998 31492 71062
rect 31144 70932 31492 70998
rect 31824 71062 32036 71068
rect 31824 70998 31966 71062
rect 32030 70998 32036 71062
rect 31824 70932 32036 70998
rect 30600 70856 32036 70932
rect 32504 71062 32716 71068
rect 32504 70998 32510 71062
rect 32574 70998 32716 71062
rect 32504 70932 32716 70998
rect 33048 70932 33260 71068
rect 33728 71062 34620 71068
rect 33728 70998 33734 71062
rect 33798 70998 34414 71062
rect 34478 70998 34620 71062
rect 33728 70992 34620 70998
rect 33728 70932 33940 70992
rect 32504 70856 33940 70932
rect 34272 70856 34620 70992
rect 34952 71062 35164 71068
rect 34952 70998 34958 71062
rect 35022 70998 35164 71062
rect 34952 70932 35164 70998
rect 35632 71062 35844 71068
rect 35632 70998 35774 71062
rect 35838 70998 35844 71062
rect 35632 70932 35844 70998
rect 34952 70856 35844 70932
rect 36176 71062 37068 71068
rect 36176 70998 36182 71062
rect 36246 70998 36998 71062
rect 37062 70998 37068 71062
rect 36176 70992 37068 70998
rect 36176 70856 36388 70992
rect 36856 70856 37068 70992
rect 37400 71062 37748 71068
rect 37400 70998 37542 71062
rect 37606 70998 37748 71062
rect 37400 70932 37748 70998
rect 38080 71062 38972 71068
rect 38080 70998 38222 71062
rect 38286 70998 38972 71062
rect 38080 70992 38972 70998
rect 38080 70932 38292 70992
rect 37400 70856 38292 70932
rect 38760 70932 38972 70992
rect 39304 70932 39516 71068
rect 39984 71062 40740 71068
rect 39984 70998 39990 71062
rect 40054 70998 40670 71062
rect 40734 70998 40740 71062
rect 39984 70992 40740 70998
rect 39984 70932 40196 70992
rect 38760 70856 40196 70932
rect 40528 70856 40740 70992
rect 41208 71062 41420 71068
rect 41208 70998 41214 71062
rect 41278 70998 41420 71062
rect 41208 70932 41420 70998
rect 41752 71062 42100 71068
rect 41752 70998 41894 71062
rect 41958 70998 42100 71062
rect 41752 70932 42100 70998
rect 41208 70856 42100 70932
rect 42432 71062 43324 71068
rect 42432 70998 42438 71062
rect 42502 70998 43254 71062
rect 43318 70998 43324 71062
rect 42432 70992 43324 70998
rect 42432 70856 42644 70992
rect 43112 70932 43324 70992
rect 43656 70932 43868 71068
rect 44336 70992 45228 71068
rect 44336 70932 44548 70992
rect 44880 70932 45228 70992
rect 43112 70856 44548 70932
rect 44646 70926 45228 70932
rect 44608 70862 44614 70926
rect 44678 70862 45228 70926
rect 44646 70856 45228 70862
rect 45560 71062 45772 71068
rect 45560 70998 45702 71062
rect 45766 70998 45772 71062
rect 45560 70856 45772 70998
rect 46240 71062 47676 71068
rect 46240 70998 46246 71062
rect 46310 70998 46926 71062
rect 46990 70998 47676 71062
rect 46240 70992 47676 70998
rect 46240 70856 46452 70992
rect 46784 70856 46996 70992
rect 47464 70932 47676 70992
rect 48008 71062 49580 71068
rect 48008 70998 48694 71062
rect 48758 70998 49580 71062
rect 48008 70992 49580 70998
rect 48008 70932 48356 70992
rect 47464 70856 48356 70932
rect 48688 70856 48900 70992
rect 49368 70932 49580 70992
rect 49912 71062 50124 71068
rect 49912 70998 49918 71062
rect 49982 70998 50124 71062
rect 49912 70932 50124 70998
rect 50592 71062 50804 71068
rect 50592 70998 50734 71062
rect 50798 70998 50804 71062
rect 50592 70932 50804 70998
rect 49368 70856 50804 70932
rect 51136 71062 52028 71068
rect 51136 70998 51278 71062
rect 51342 70998 52028 71062
rect 51136 70992 52028 70998
rect 51136 70856 51348 70992
rect 51816 70932 52028 70992
rect 52360 71062 53252 71068
rect 53350 71062 53932 71068
rect 52360 70998 52502 71062
rect 52566 70998 53182 71062
rect 53246 70998 53252 71062
rect 53312 70998 53318 71062
rect 53382 70998 53932 71062
rect 52360 70992 53252 70998
rect 53350 70992 53932 70998
rect 52360 70932 52708 70992
rect 51816 70856 52708 70932
rect 53040 70856 53252 70992
rect 53720 70932 53932 70992
rect 54264 71062 54476 71068
rect 54264 70998 54406 71062
rect 54470 70998 54476 71062
rect 54264 70932 54476 70998
rect 53720 70856 54476 70932
rect 54944 71062 56108 71068
rect 54944 70998 54950 71062
rect 55014 70998 56038 71062
rect 56102 70998 56108 71062
rect 54944 70992 56108 70998
rect 54944 70856 55156 70992
rect 55488 70932 55836 70992
rect 56168 70932 56380 71068
rect 56848 71062 58284 71068
rect 56848 70998 57398 71062
rect 57462 70998 58284 71062
rect 56848 70992 58284 70998
rect 56848 70932 57060 70992
rect 55488 70856 57060 70932
rect 57392 70856 57604 70992
rect 58072 70932 58284 70992
rect 58616 71062 58964 71068
rect 58616 70998 58622 71062
rect 58686 70998 58964 71062
rect 58616 70932 58964 70998
rect 59296 71062 59508 71068
rect 59296 70998 59438 71062
rect 59502 70998 59508 71062
rect 59296 70932 59508 70998
rect 58072 70856 59508 70932
rect 59976 71062 60188 71068
rect 59976 70998 59982 71062
rect 60046 70998 60188 71062
rect 59976 70932 60188 70998
rect 60520 70932 60732 71068
rect 61200 71062 61956 71068
rect 61200 70998 61206 71062
rect 61270 70998 61886 71062
rect 61950 70998 61956 71062
rect 61200 70992 61956 70998
rect 61200 70932 61412 70992
rect 59976 70856 61412 70932
rect 61744 70856 61956 70992
rect 62424 71062 62636 71068
rect 62424 70998 62430 71062
rect 62494 70998 62636 71062
rect 62424 70932 62636 70998
rect 62968 71062 63316 71068
rect 62968 70998 63110 71062
rect 63174 70998 63316 71062
rect 62968 70932 63316 70998
rect 62424 70856 63316 70932
rect 63648 71062 64540 71068
rect 63648 70998 63654 71062
rect 63718 70998 64540 71062
rect 63648 70992 64540 70998
rect 63648 70856 63860 70992
rect 64328 70932 64540 70992
rect 64872 71062 65084 71068
rect 64872 70998 65014 71062
rect 65078 70998 65084 71062
rect 64872 70932 65084 70998
rect 65552 71062 66988 71068
rect 65552 70998 66102 71062
rect 66166 70998 66918 71062
rect 66982 70998 66988 71062
rect 65552 70992 66988 70998
rect 65552 70932 65764 70992
rect 64328 70856 65764 70932
rect 66096 70856 66444 70992
rect 66776 70856 66988 70992
rect 67456 71062 68212 71068
rect 67456 70998 67462 71062
rect 67526 70998 68142 71062
rect 68206 70998 68212 71062
rect 67456 70992 68212 70998
rect 67456 70856 67668 70992
rect 68000 70856 68212 70992
rect 68680 71062 68892 71068
rect 68680 70998 68686 71062
rect 68750 70998 68892 71062
rect 68680 70932 68892 70998
rect 69224 70932 69572 71068
rect 69904 71062 70796 71068
rect 69904 70998 69910 71062
rect 69974 70998 70590 71062
rect 70654 70998 70796 71062
rect 69904 70992 70796 70998
rect 69904 70932 70116 70992
rect 68680 70856 70116 70932
rect 70584 70932 70796 70992
rect 71128 70932 71340 71068
rect 71808 71062 72292 71068
rect 71808 70998 72222 71062
rect 72286 70998 72292 71062
rect 71808 70992 72292 70998
rect 72352 70992 73244 71068
rect 71808 70932 72020 70992
rect 72352 70932 72564 70992
rect 70584 70856 72020 70932
rect 72118 70926 72564 70932
rect 72080 70862 72086 70926
rect 72150 70862 72564 70926
rect 72118 70856 72564 70862
rect 73032 70932 73244 70992
rect 73576 71062 73924 71068
rect 73576 70998 73718 71062
rect 73782 70998 73924 71062
rect 73576 70932 73924 70998
rect 74256 71062 74468 71068
rect 74256 70998 74398 71062
rect 74462 70998 74468 71062
rect 74256 70932 74468 70998
rect 73032 70856 74468 70932
rect 74936 71062 75148 71068
rect 74936 70998 74942 71062
rect 75006 70998 75148 71062
rect 74936 70932 75148 70998
rect 75480 71062 75692 71068
rect 75480 70998 75622 71062
rect 75686 70998 75692 71062
rect 75480 70932 75692 70998
rect 74936 70856 75692 70932
rect 76160 71062 77052 71068
rect 76160 70998 76166 71062
rect 76230 70998 76846 71062
rect 76910 70998 77052 71062
rect 76160 70992 77052 70998
rect 76160 70856 76372 70992
rect 76704 70856 77052 70992
rect 77384 71062 77596 71068
rect 77384 70998 77390 71062
rect 77454 70998 77596 71062
rect 77384 70932 77596 70998
rect 78064 71062 78548 71068
rect 78064 70998 78206 71062
rect 78270 70998 78478 71062
rect 78542 70998 78548 71062
rect 78064 70992 78548 70998
rect 78608 71062 79500 71068
rect 78608 70998 79430 71062
rect 79494 70998 79500 71062
rect 78608 70992 79500 70998
rect 78064 70932 78276 70992
rect 78608 70932 78820 70992
rect 77384 70856 78820 70932
rect 79288 70856 79500 70992
rect 79832 71062 80180 71068
rect 79832 70998 79974 71062
rect 80038 70998 80180 71062
rect 79832 70932 80180 70998
rect 80512 71062 81404 71068
rect 80512 70998 80654 71062
rect 80718 70998 81404 71062
rect 80512 70992 81404 70998
rect 80512 70932 80724 70992
rect 79832 70856 80724 70932
rect 81192 70932 81404 70992
rect 81736 71062 81948 71068
rect 81736 70998 81878 71062
rect 81942 70998 81948 71062
rect 81736 70932 81948 70998
rect 81192 70856 81948 70932
rect 82416 71062 83172 71068
rect 82416 70998 82422 71062
rect 82486 70998 83102 71062
rect 83166 70998 83172 71062
rect 82416 70992 83172 70998
rect 82416 70856 82628 70992
rect 82960 70856 83172 70992
rect 83640 71062 83852 71068
rect 83640 70998 83646 71062
rect 83710 70998 83852 71062
rect 83640 70932 83852 70998
rect 84184 70932 84532 71068
rect 84630 71062 85756 71068
rect 84592 70998 84598 71062
rect 84662 70998 85756 71062
rect 84630 70992 85756 70998
rect 84864 70932 85076 70992
rect 83640 70856 85076 70932
rect 85544 70932 85756 70992
rect 86088 71062 86300 71068
rect 86088 70998 86094 71062
rect 86158 70998 86300 71062
rect 86088 70932 86300 70998
rect 86768 71062 88204 71068
rect 86768 70998 86910 71062
rect 86974 70998 88134 71062
rect 88198 70998 88204 71062
rect 86768 70992 88204 70998
rect 86768 70932 86980 70992
rect 85544 70856 86980 70932
rect 87312 70856 87660 70992
rect 87992 70856 88204 70992
rect 88672 71062 89428 71068
rect 88672 70998 88678 71062
rect 88742 70998 89358 71062
rect 89422 70998 89428 71062
rect 88672 70992 89428 70998
rect 88672 70856 88884 70992
rect 89216 70856 89428 70992
rect 89896 71062 90108 71068
rect 89896 70998 89902 71062
rect 89966 70998 90108 71062
rect 89896 70932 90108 70998
rect 90440 71062 90788 71068
rect 90440 70998 90718 71062
rect 90782 70998 90788 71062
rect 90440 70932 90788 70998
rect 89896 70856 90788 70932
rect 91120 71062 92012 71068
rect 91120 70998 91126 71062
rect 91190 70998 92012 71062
rect 91120 70992 92012 70998
rect 91120 70856 91332 70992
rect 91800 70932 92012 70992
rect 92344 71062 92556 71068
rect 92344 70998 92350 71062
rect 92414 70998 92556 71062
rect 92344 70932 92556 70998
rect 93024 70992 94460 71068
rect 93024 70932 93236 70992
rect 93568 70932 93780 70992
rect 91800 70856 93236 70932
rect 93334 70926 93780 70932
rect 93296 70862 93302 70926
rect 93366 70862 93780 70926
rect 93334 70856 93780 70862
rect 94248 70932 94460 70992
rect 94792 71062 95140 71068
rect 94792 70998 94934 71062
rect 94998 70998 95140 71062
rect 94792 70932 95140 70998
rect 95472 71062 96364 71068
rect 95472 70998 95614 71062
rect 95678 70998 96364 71062
rect 95472 70992 96364 70998
rect 95472 70932 95684 70992
rect 94248 70856 95684 70932
rect 96152 70932 96364 70992
rect 96696 71062 96908 71068
rect 96696 70998 96838 71062
rect 96902 70998 96908 71062
rect 96696 70932 96908 70998
rect 96152 70856 96908 70932
rect 97376 71062 98268 71068
rect 97376 70998 97382 71062
rect 97446 70998 98268 71062
rect 97376 70992 98268 70998
rect 97376 70856 97588 70992
rect 97920 70932 98268 70992
rect 98600 71062 98812 71068
rect 98600 70998 98606 71062
rect 98670 70998 98812 71062
rect 98600 70932 98812 70998
rect 99280 71062 100988 71068
rect 99280 70998 99830 71062
rect 99894 70998 100918 71062
rect 100982 70998 100988 71062
rect 99280 70992 100988 70998
rect 99280 70932 99492 70992
rect 97920 70856 99492 70932
rect 99824 70856 100036 70992
rect 100504 70932 100716 70992
rect 101048 70932 101396 71068
rect 101728 71062 101940 71068
rect 101728 70998 101870 71062
rect 101934 70998 101940 71062
rect 101728 70932 101940 70998
rect 100504 70856 101940 70932
rect 102408 71062 102620 71068
rect 102408 70998 102414 71062
rect 102478 70998 102620 71062
rect 102408 70932 102620 70998
rect 102952 71062 103164 71068
rect 102952 70998 103094 71062
rect 103158 70998 103164 71062
rect 102952 70932 103164 70998
rect 102408 70856 103164 70932
rect 103632 71062 104388 71068
rect 103632 70998 103638 71062
rect 103702 70998 104318 71062
rect 104382 70998 104388 71062
rect 103632 70992 104388 70998
rect 103632 70856 103844 70992
rect 104176 70856 104388 70992
rect 104856 71062 105068 71068
rect 104856 70998 104862 71062
rect 104926 70998 105068 71062
rect 104856 70932 105068 70998
rect 105400 71062 105748 71068
rect 105400 70998 105542 71062
rect 105606 70998 105748 71062
rect 105400 70932 105748 70998
rect 104856 70856 105748 70932
rect 106080 71062 106972 71068
rect 106080 70998 106086 71062
rect 106150 70998 106972 71062
rect 106080 70992 106972 70998
rect 106080 70856 106292 70992
rect 106760 70932 106972 70992
rect 107304 71062 107516 71068
rect 107304 70998 107310 71062
rect 107374 70998 107516 71062
rect 107304 70932 107516 70998
rect 107984 71062 110780 71068
rect 107984 70998 108534 71062
rect 108598 70998 110710 71062
rect 110774 70998 110780 71062
rect 107984 70992 110780 70998
rect 134776 71062 134988 71068
rect 134776 70998 134782 71062
rect 134846 70998 134988 71062
rect 107984 70932 108196 70992
rect 106760 70856 108196 70932
rect 108528 70856 108876 70992
rect 134776 70968 134988 70998
rect 109616 70926 109828 70932
rect 109616 70862 109622 70926
rect 109686 70862 109828 70926
rect 27064 70790 29044 70796
rect 27064 70726 28974 70790
rect 29038 70726 29044 70790
rect 27064 70720 29044 70726
rect 27064 70660 27276 70720
rect 27064 70584 27412 70660
rect 27336 70524 27412 70584
rect 109616 70584 109828 70862
rect 134776 70912 134844 70968
rect 134900 70932 134988 70968
rect 134900 70926 135396 70932
rect 134900 70912 135326 70926
rect 134776 70862 135326 70912
rect 135390 70862 135396 70926
rect 134776 70856 135396 70862
rect 110704 70654 110916 70660
rect 110704 70590 110710 70654
rect 110774 70590 110916 70654
rect 109616 70524 109692 70584
rect 27336 70312 27684 70524
rect 109344 70448 109692 70524
rect 110704 70524 110916 70590
rect 113424 70524 113636 70660
rect 114240 70654 115404 70660
rect 114240 70590 115334 70654
rect 115398 70590 115404 70654
rect 114240 70584 115404 70590
rect 114240 70524 114452 70584
rect 110704 70518 114452 70524
rect 110704 70454 114246 70518
rect 114310 70454 114452 70518
rect 110704 70448 114452 70454
rect 109344 70312 109556 70448
rect 27336 70252 27412 70312
rect 109480 70252 109556 70312
rect 20808 69904 21020 70116
rect 21216 70040 21972 70116
rect 21216 69904 21428 70040
rect 21624 69904 21972 70040
rect 22032 69974 22244 70116
rect 22032 69910 22174 69974
rect 22238 69910 22244 69974
rect 22032 69904 22244 69910
rect 22440 69974 22652 70116
rect 27336 70040 27684 70252
rect 27608 69980 27684 70040
rect 22440 69910 22446 69974
rect 22510 69910 22652 69974
rect 22440 69904 22652 69910
rect 20944 69844 21020 69904
rect 21624 69844 21700 69904
rect 20808 69566 21020 69844
rect 21352 69768 21700 69844
rect 27336 69768 27684 69980
rect 109344 70040 109556 70252
rect 114240 70110 114452 70116
rect 114240 70046 114246 70110
rect 114310 70046 114452 70110
rect 109344 69980 109420 70040
rect 109344 69768 109556 69980
rect 114240 69974 114452 70046
rect 114240 69910 114382 69974
rect 114446 69910 114452 69974
rect 114240 69904 114452 69910
rect 114648 69974 114860 70116
rect 114648 69910 114654 69974
rect 114718 69910 114860 69974
rect 114648 69904 114860 69910
rect 115056 69980 115268 70116
rect 115056 69974 115404 69980
rect 115056 69910 115334 69974
rect 115398 69910 115404 69974
rect 115056 69904 115404 69910
rect 115464 69974 115676 70116
rect 115464 69910 115470 69974
rect 115534 69910 115676 69974
rect 115464 69904 115676 69910
rect 115872 70110 116084 70116
rect 115872 70046 115878 70110
rect 115942 70046 116084 70110
rect 115872 69904 116084 70046
rect 132600 69904 133492 69980
rect 115872 69844 115948 69904
rect 21352 69708 21428 69768
rect 27472 69708 27548 69768
rect 109344 69708 109420 69768
rect 20808 69502 20814 69566
rect 20878 69502 21020 69566
rect 20808 69496 21020 69502
rect 21216 69632 21972 69708
rect 21216 69566 21428 69632
rect 21216 69502 21358 69566
rect 21422 69502 21428 69566
rect 21216 69496 21428 69502
rect 21624 69566 21972 69632
rect 21624 69502 21630 69566
rect 21694 69502 21972 69566
rect 21624 69496 21972 69502
rect 22032 69702 22244 69708
rect 22032 69638 22174 69702
rect 22238 69638 22244 69702
rect 22032 69566 22244 69638
rect 22032 69502 22174 69566
rect 22238 69502 22244 69566
rect 22032 69496 22244 69502
rect 22440 69702 22652 69708
rect 22440 69638 22446 69702
rect 22510 69638 22652 69702
rect 22440 69566 22652 69638
rect 22440 69502 22446 69566
rect 22510 69502 22652 69566
rect 22440 69496 22652 69502
rect 27336 69496 27684 69708
rect 109344 69496 109556 69708
rect 114240 69702 114452 69708
rect 114240 69638 114382 69702
rect 114446 69638 114452 69702
rect 114240 69566 114452 69638
rect 114240 69502 114246 69566
rect 114310 69502 114452 69566
rect 114240 69496 114452 69502
rect 114648 69702 114860 69708
rect 114648 69638 114654 69702
rect 114718 69638 114860 69702
rect 114648 69566 114860 69638
rect 114648 69502 114654 69566
rect 114718 69502 114860 69566
rect 114648 69496 114860 69502
rect 115056 69566 115268 69708
rect 115366 69702 115676 69708
rect 115328 69638 115334 69702
rect 115398 69638 115470 69702
rect 115534 69638 115676 69702
rect 115366 69632 115676 69638
rect 115056 69502 115062 69566
rect 115126 69502 115268 69566
rect 115056 69496 115268 69502
rect 115464 69566 115676 69632
rect 115464 69502 115606 69566
rect 115670 69502 115676 69566
rect 115464 69496 115676 69502
rect 115872 69566 116084 69844
rect 132600 69768 132812 69904
rect 133280 69844 133492 69904
rect 133182 69838 133492 69844
rect 133144 69774 133150 69838
rect 133214 69774 133492 69838
rect 133182 69768 133492 69774
rect 115872 69502 116014 69566
rect 116078 69502 116084 69566
rect 115872 69496 116084 69502
rect 27472 69436 27548 69496
rect 109480 69436 109556 69496
rect 1768 69300 1980 69436
rect 1224 69294 1980 69300
rect 1224 69230 1230 69294
rect 1294 69288 1980 69294
rect 1294 69232 1794 69288
rect 1850 69232 1980 69288
rect 1294 69230 1980 69232
rect 1224 69224 1980 69230
rect 1768 69088 1980 69224
rect 20808 69294 21020 69300
rect 20808 69230 20814 69294
rect 20878 69230 21020 69294
rect 20808 69088 21020 69230
rect 21216 69294 21428 69300
rect 21216 69230 21358 69294
rect 21422 69230 21428 69294
rect 21216 69088 21428 69230
rect 21624 69294 21972 69300
rect 21624 69230 21630 69294
rect 21694 69230 21972 69294
rect 21624 69158 21972 69230
rect 21624 69094 21766 69158
rect 21830 69094 21972 69158
rect 21624 69088 21972 69094
rect 22032 69294 22244 69300
rect 22032 69230 22174 69294
rect 22238 69230 22244 69294
rect 22032 69158 22244 69230
rect 22032 69094 22038 69158
rect 22102 69094 22244 69158
rect 22032 69088 22244 69094
rect 22440 69294 22652 69300
rect 22440 69230 22446 69294
rect 22510 69230 22652 69294
rect 22440 69158 22652 69230
rect 27336 69224 27684 69436
rect 109344 69224 109556 69436
rect 134776 69430 135396 69436
rect 134776 69366 135326 69430
rect 135390 69366 135396 69430
rect 134776 69360 135396 69366
rect 27472 69164 27548 69224
rect 109480 69164 109556 69224
rect 22440 69094 22446 69158
rect 22510 69094 22652 69158
rect 22440 69088 22652 69094
rect 20808 69028 20884 69088
rect 20808 68886 21020 69028
rect 27336 68952 27684 69164
rect 109344 68952 109556 69164
rect 114240 69294 114452 69300
rect 114240 69230 114246 69294
rect 114310 69230 114452 69294
rect 114240 69158 114452 69230
rect 114240 69094 114382 69158
rect 114446 69094 114452 69158
rect 114240 69088 114452 69094
rect 114648 69294 114860 69300
rect 114648 69230 114654 69294
rect 114718 69230 114860 69294
rect 114648 69158 114860 69230
rect 114648 69094 114790 69158
rect 114854 69094 114860 69158
rect 114648 69088 114860 69094
rect 115056 69294 115268 69300
rect 115056 69230 115062 69294
rect 115126 69230 115268 69294
rect 115056 69158 115268 69230
rect 115056 69094 115198 69158
rect 115262 69094 115268 69158
rect 115056 69088 115268 69094
rect 115464 69294 115676 69300
rect 115464 69230 115606 69294
rect 115670 69230 115676 69294
rect 115464 69088 115676 69230
rect 115872 69294 116084 69300
rect 115872 69230 116014 69294
rect 116078 69230 116084 69294
rect 115872 69088 116084 69230
rect 134776 69288 134988 69360
rect 134776 69232 134844 69288
rect 134900 69232 134988 69288
rect 134776 69158 134988 69232
rect 134776 69094 134782 69158
rect 134846 69094 134988 69158
rect 134776 69088 134988 69094
rect 115464 69028 115540 69088
rect 115192 68952 115540 69028
rect 115872 69028 115948 69088
rect 27472 68892 27548 68952
rect 109344 68892 109420 68952
rect 115192 68892 115268 68952
rect 20808 68822 20814 68886
rect 20878 68822 21020 68886
rect 20808 68816 21020 68822
rect 21216 68680 21428 68892
rect 21624 68886 21972 68892
rect 21624 68822 21766 68886
rect 21830 68822 21972 68886
rect 21624 68756 21972 68822
rect 21488 68680 21972 68756
rect 22032 68886 22244 68892
rect 22032 68822 22038 68886
rect 22102 68822 22244 68886
rect 22032 68750 22244 68822
rect 22032 68686 22038 68750
rect 22102 68686 22244 68750
rect 22032 68680 22244 68686
rect 22440 68886 22652 68892
rect 22440 68822 22446 68886
rect 22510 68822 22652 68886
rect 22440 68750 22652 68822
rect 22440 68686 22446 68750
rect 22510 68686 22652 68750
rect 22440 68680 22652 68686
rect 21216 68620 21292 68680
rect 21488 68620 21564 68680
rect 20808 68614 21020 68620
rect 20808 68550 20814 68614
rect 20878 68550 21020 68614
rect 20808 68272 21020 68550
rect 21216 68544 21564 68620
rect 21624 68620 21700 68680
rect 21216 68272 21428 68544
rect 21624 68342 21972 68620
rect 21624 68278 21902 68342
rect 21966 68278 21972 68342
rect 21624 68272 21972 68278
rect 22032 68478 22244 68484
rect 22032 68414 22038 68478
rect 22102 68414 22244 68478
rect 22032 68272 22244 68414
rect 22440 68478 22652 68484
rect 22440 68414 22446 68478
rect 22510 68414 22652 68478
rect 22440 68272 22652 68414
rect 27336 68408 27684 68892
rect 109344 68408 109556 68892
rect 114240 68886 114452 68892
rect 114240 68822 114382 68886
rect 114446 68822 114452 68886
rect 114240 68756 114452 68822
rect 114648 68886 114860 68892
rect 114648 68822 114790 68886
rect 114854 68822 114860 68886
rect 114240 68750 114588 68756
rect 114240 68686 114382 68750
rect 114446 68686 114588 68750
rect 114240 68680 114588 68686
rect 114648 68750 114860 68822
rect 114648 68686 114654 68750
rect 114718 68686 114860 68750
rect 114648 68680 114860 68686
rect 115056 68886 115676 68892
rect 115056 68822 115198 68886
rect 115262 68822 115676 68886
rect 115056 68816 115676 68822
rect 115872 68886 116084 69028
rect 115872 68822 116014 68886
rect 116078 68822 116084 68886
rect 115872 68816 116084 68822
rect 115056 68680 115268 68816
rect 114512 68620 114588 68680
rect 115192 68620 115268 68680
rect 114512 68544 115268 68620
rect 27472 68348 27548 68408
rect 109480 68348 109556 68408
rect 20944 68212 21020 68272
rect 22168 68212 22244 68272
rect 22576 68212 22652 68272
rect 20808 68070 21020 68212
rect 20808 68006 20814 68070
rect 20878 68006 21020 68070
rect 20808 68000 21020 68006
rect 21216 67864 21428 68076
rect 21624 68070 21972 68076
rect 21624 68006 21902 68070
rect 21966 68006 21972 68070
rect 21624 67864 21972 68006
rect 21216 67804 21292 67864
rect 21896 67804 21972 67864
rect 20808 67798 21020 67804
rect 20808 67734 20814 67798
rect 20878 67734 21020 67798
rect 1768 67608 1980 67668
rect 1768 67552 1794 67608
rect 1850 67552 1980 67608
rect 20808 67662 21020 67734
rect 20808 67598 20814 67662
rect 20878 67598 21020 67662
rect 20808 67592 21020 67598
rect 21216 67662 21428 67804
rect 21216 67598 21222 67662
rect 21286 67598 21428 67662
rect 21216 67592 21428 67598
rect 21624 67662 21972 67804
rect 21624 67598 21630 67662
rect 21694 67598 21972 67662
rect 21624 67592 21972 67598
rect 22032 67864 22244 68212
rect 22440 67864 22652 68212
rect 27336 68206 27684 68348
rect 27336 68142 27478 68206
rect 27542 68142 27684 68206
rect 27336 67934 27684 68142
rect 27336 67870 27342 67934
rect 27406 67870 27478 67934
rect 27542 67870 27684 67934
rect 22032 67804 22108 67864
rect 22440 67804 22516 67864
rect 1768 67532 1980 67552
rect 1224 67526 1980 67532
rect 1224 67462 1230 67526
rect 1294 67462 1980 67526
rect 1224 67456 1980 67462
rect 22032 67456 22244 67804
rect 22168 67396 22244 67456
rect 20808 67390 21020 67396
rect 20808 67326 20814 67390
rect 20878 67326 21020 67390
rect 20808 67254 21020 67326
rect 20808 67190 20814 67254
rect 20878 67190 21020 67254
rect 20808 67184 21020 67190
rect 21216 67390 21428 67396
rect 21216 67326 21222 67390
rect 21286 67326 21428 67390
rect 21216 67260 21428 67326
rect 21624 67390 21972 67396
rect 21624 67326 21630 67390
rect 21694 67326 21972 67390
rect 21216 67254 21564 67260
rect 21216 67190 21494 67254
rect 21558 67190 21564 67254
rect 21216 67184 21564 67190
rect 21216 67124 21428 67184
rect 21624 67124 21972 67326
rect 22032 67254 22244 67396
rect 22032 67190 22038 67254
rect 22102 67190 22244 67254
rect 22032 67184 22244 67190
rect 22440 67456 22652 67804
rect 27336 67728 27684 67870
rect 109344 68206 109556 68348
rect 109344 68142 109486 68206
rect 109550 68142 109556 68206
rect 109344 67934 109556 68142
rect 109344 67870 109486 67934
rect 109550 67870 109556 67934
rect 109344 67798 109556 67870
rect 114240 68478 114452 68484
rect 114240 68414 114382 68478
rect 114446 68414 114452 68478
rect 114240 68272 114452 68414
rect 114648 68478 114860 68484
rect 114648 68414 114654 68478
rect 114718 68414 114860 68478
rect 114648 68272 114860 68414
rect 115056 68272 115268 68544
rect 115464 68680 115676 68816
rect 115464 68620 115540 68680
rect 115464 68348 115676 68620
rect 115366 68342 115676 68348
rect 115328 68278 115334 68342
rect 115398 68278 115676 68342
rect 115366 68272 115676 68278
rect 115872 68614 116084 68620
rect 115872 68550 116014 68614
rect 116078 68550 116084 68614
rect 115872 68272 116084 68550
rect 132600 68484 132812 68620
rect 133280 68614 134852 68620
rect 133280 68550 134782 68614
rect 134846 68550 134852 68614
rect 133280 68544 134852 68550
rect 133280 68484 133492 68544
rect 132600 68408 133492 68484
rect 114240 68212 114316 68272
rect 114648 68212 114724 68272
rect 116008 68212 116084 68272
rect 114240 67864 114452 68212
rect 114648 67864 114860 68212
rect 115056 68070 115404 68076
rect 115056 68006 115334 68070
rect 115398 68006 115404 68070
rect 115056 68000 115404 68006
rect 115056 67864 115268 68000
rect 115464 67940 115676 68076
rect 115872 68070 116084 68212
rect 115872 68006 115878 68070
rect 115942 68006 116084 68070
rect 115872 68000 116084 68006
rect 114376 67804 114452 67864
rect 114784 67804 114860 67864
rect 115192 67804 115268 67864
rect 115328 67864 115676 67940
rect 115328 67804 115404 67864
rect 109344 67734 109350 67798
rect 109414 67734 109556 67798
rect 109344 67728 109556 67734
rect 27336 67668 27412 67728
rect 27336 67662 27684 67668
rect 27336 67598 27342 67662
rect 27406 67598 27684 67662
rect 27336 67592 27684 67598
rect 109344 67592 109556 67668
rect 22440 67396 22516 67456
rect 27462 67396 27560 67592
rect 109344 67396 109448 67592
rect 114240 67456 114452 67804
rect 114648 67456 114860 67804
rect 115056 67728 115404 67804
rect 115056 67668 115268 67728
rect 115464 67668 115676 67804
rect 115056 67662 115676 67668
rect 115056 67598 115606 67662
rect 115670 67598 115676 67662
rect 115056 67592 115676 67598
rect 115872 67798 116084 67804
rect 115872 67734 115878 67798
rect 115942 67734 116084 67798
rect 115872 67662 116084 67734
rect 115872 67598 116014 67662
rect 116078 67598 116084 67662
rect 115872 67592 116084 67598
rect 134776 67662 135396 67668
rect 134776 67608 135326 67662
rect 134776 67552 134844 67608
rect 134900 67598 135326 67608
rect 135390 67598 135396 67662
rect 134900 67592 135396 67598
rect 134900 67552 134988 67592
rect 134776 67456 134988 67552
rect 114240 67396 114316 67456
rect 114648 67396 114724 67456
rect 22440 67254 22652 67396
rect 22440 67190 22446 67254
rect 22510 67190 22652 67254
rect 22440 67184 22652 67190
rect 27336 67184 27684 67396
rect 109344 67390 109556 67396
rect 109344 67326 109350 67390
rect 109414 67326 109486 67390
rect 109550 67326 109556 67390
rect 109344 67184 109556 67326
rect 114240 67254 114452 67396
rect 114240 67190 114382 67254
rect 114446 67190 114452 67254
rect 114240 67184 114452 67190
rect 114648 67254 114860 67396
rect 114648 67190 114654 67254
rect 114718 67190 114860 67254
rect 114648 67184 114860 67190
rect 27472 67124 27548 67184
rect 109480 67124 109556 67184
rect 21216 67048 21972 67124
rect 21352 66988 21428 67048
rect 20808 66982 21020 66988
rect 20808 66918 20814 66982
rect 20878 66918 21020 66982
rect 20808 66846 21020 66918
rect 20808 66782 20814 66846
rect 20878 66782 21020 66846
rect 20808 66776 21020 66782
rect 21216 66776 21428 66988
rect 21526 66982 21972 66988
rect 21488 66918 21494 66982
rect 21558 66918 21972 66982
rect 21526 66912 21972 66918
rect 21624 66846 21972 66912
rect 21624 66782 21630 66846
rect 21694 66782 21972 66846
rect 21624 66776 21972 66782
rect 22032 66982 22244 66988
rect 22032 66918 22038 66982
rect 22102 66918 22244 66982
rect 22032 66846 22244 66918
rect 22032 66782 22038 66846
rect 22102 66782 22244 66846
rect 22032 66776 22244 66782
rect 22440 66982 22652 66988
rect 22440 66918 22446 66982
rect 22510 66918 22652 66982
rect 22440 66846 22652 66918
rect 22440 66782 22446 66846
rect 22510 66782 22652 66846
rect 22440 66776 22652 66782
rect 27336 66912 27684 67124
rect 109344 67118 109556 67124
rect 109344 67054 109486 67118
rect 109550 67054 109556 67118
rect 109344 66912 109556 67054
rect 115056 67048 115268 67396
rect 115464 67390 115676 67396
rect 115464 67326 115606 67390
rect 115670 67326 115676 67390
rect 115464 67124 115676 67326
rect 115872 67390 116084 67396
rect 115872 67326 116014 67390
rect 116078 67326 116084 67390
rect 115872 67254 116084 67326
rect 115872 67190 115878 67254
rect 115942 67190 116084 67254
rect 115872 67184 116084 67190
rect 132600 67184 133492 67260
rect 115192 66988 115268 67048
rect 115328 67048 115676 67124
rect 132600 67124 132812 67184
rect 132600 67118 133220 67124
rect 132600 67054 133150 67118
rect 133214 67054 133220 67118
rect 132600 67048 133220 67054
rect 115328 66988 115404 67048
rect 114240 66982 114452 66988
rect 114240 66918 114382 66982
rect 114446 66918 114452 66982
rect 27336 66852 27412 66912
rect 109344 66852 109420 66912
rect 27336 66640 27684 66852
rect 109344 66640 109556 66852
rect 114240 66846 114452 66918
rect 114240 66782 114382 66846
rect 114446 66782 114452 66846
rect 114240 66776 114452 66782
rect 114648 66982 114860 66988
rect 114648 66918 114654 66982
rect 114718 66918 114860 66982
rect 114648 66846 114860 66918
rect 114648 66782 114790 66846
rect 114854 66782 114860 66846
rect 114648 66776 114860 66782
rect 115056 66912 115404 66988
rect 115056 66852 115268 66912
rect 115464 66852 115676 66988
rect 115056 66846 115676 66852
rect 115056 66782 115606 66846
rect 115670 66782 115676 66846
rect 115056 66776 115676 66782
rect 115872 66982 116084 66988
rect 115872 66918 115878 66982
rect 115942 66918 116084 66982
rect 115872 66846 116084 66918
rect 132600 66982 132812 67048
rect 132600 66918 132606 66982
rect 132670 66918 132812 66982
rect 132600 66912 132812 66918
rect 133280 66912 133492 67184
rect 115872 66782 115878 66846
rect 115942 66782 116084 66846
rect 115872 66776 116084 66782
rect 27472 66580 27548 66640
rect 109344 66580 109420 66640
rect 20808 66574 21020 66580
rect 20808 66510 20814 66574
rect 20878 66510 21020 66574
rect 20808 66438 21020 66510
rect 20808 66374 20950 66438
rect 21014 66374 21020 66438
rect 20808 66368 21020 66374
rect 21216 66574 21972 66580
rect 21216 66510 21630 66574
rect 21694 66510 21972 66574
rect 21216 66504 21972 66510
rect 21216 66444 21428 66504
rect 21216 66438 21564 66444
rect 21216 66374 21358 66438
rect 21422 66374 21494 66438
rect 21558 66374 21564 66438
rect 21216 66368 21564 66374
rect 21624 66368 21972 66504
rect 22032 66574 22244 66580
rect 22032 66510 22038 66574
rect 22102 66510 22244 66574
rect 22032 66438 22244 66510
rect 22032 66374 22174 66438
rect 22238 66374 22244 66438
rect 22032 66368 22244 66374
rect 22440 66574 22652 66580
rect 22440 66510 22446 66574
rect 22510 66510 22652 66574
rect 22440 66438 22652 66510
rect 22440 66374 22582 66438
rect 22646 66374 22652 66438
rect 22440 66368 22652 66374
rect 27336 66368 27684 66580
rect 109344 66368 109556 66580
rect 114240 66574 114452 66580
rect 114240 66510 114382 66574
rect 114446 66510 114452 66574
rect 114240 66438 114452 66510
rect 114240 66374 114246 66438
rect 114310 66374 114452 66438
rect 114240 66368 114452 66374
rect 114648 66574 114860 66580
rect 114648 66510 114790 66574
rect 114854 66510 114860 66574
rect 114648 66438 114860 66510
rect 114648 66374 114654 66438
rect 114718 66374 114860 66438
rect 114648 66368 114860 66374
rect 115056 66574 115676 66580
rect 115056 66510 115606 66574
rect 115670 66510 115676 66574
rect 115056 66504 115676 66510
rect 115056 66444 115268 66504
rect 115056 66438 115404 66444
rect 115056 66374 115062 66438
rect 115126 66374 115334 66438
rect 115398 66374 115404 66438
rect 115056 66368 115404 66374
rect 115464 66368 115676 66504
rect 115872 66574 116084 66580
rect 115872 66510 115878 66574
rect 115942 66510 116084 66574
rect 115872 66438 116084 66510
rect 115872 66374 116014 66438
rect 116078 66374 116084 66438
rect 115872 66368 116084 66374
rect 27608 66308 27684 66368
rect 109480 66308 109556 66368
rect 20808 66166 21020 66172
rect 20808 66102 20950 66166
rect 21014 66102 21020 66166
rect 1224 66030 1980 66036
rect 1224 65966 1230 66030
rect 1294 65966 1980 66030
rect 1224 65960 1980 65966
rect 20808 66030 21020 66102
rect 20808 65966 20814 66030
rect 20878 65966 21020 66030
rect 20808 65960 21020 65966
rect 21216 66166 21428 66172
rect 21526 66166 21972 66172
rect 21216 66102 21358 66166
rect 21422 66102 21428 66166
rect 21488 66102 21494 66166
rect 21558 66102 21972 66166
rect 21216 65960 21428 66102
rect 21526 66096 21972 66102
rect 21624 66030 21972 66096
rect 21624 65966 21766 66030
rect 21830 65966 21972 66030
rect 21624 65960 21972 65966
rect 22032 66166 22244 66172
rect 22032 66102 22174 66166
rect 22238 66102 22244 66166
rect 22032 66030 22244 66102
rect 22032 65966 22038 66030
rect 22102 65966 22244 66030
rect 22032 65960 22244 65966
rect 22440 66166 22652 66172
rect 22440 66102 22582 66166
rect 22646 66102 22652 66166
rect 22440 66030 22652 66102
rect 27336 66096 27684 66308
rect 109344 66096 109556 66308
rect 27608 66036 27684 66096
rect 109480 66036 109556 66096
rect 22440 65966 22582 66030
rect 22646 65966 22652 66030
rect 22440 65960 22652 65966
rect 1768 65928 1980 65960
rect 1768 65872 1794 65928
rect 1850 65872 1980 65928
rect 1768 65824 1980 65872
rect 27336 65824 27684 66036
rect 27608 65764 27684 65824
rect 20808 65758 21020 65764
rect 20808 65694 20814 65758
rect 20878 65694 21020 65758
rect 20808 65622 21020 65694
rect 20808 65558 20950 65622
rect 21014 65558 21020 65622
rect 20808 65552 21020 65558
rect 21216 65622 21428 65764
rect 21624 65758 21972 65764
rect 21624 65694 21766 65758
rect 21830 65694 21972 65758
rect 21624 65628 21972 65694
rect 21526 65622 21972 65628
rect 21216 65558 21358 65622
rect 21422 65558 21428 65622
rect 21488 65558 21494 65622
rect 21558 65558 21972 65622
rect 21216 65552 21428 65558
rect 21526 65552 21972 65558
rect 22032 65758 22244 65764
rect 22032 65694 22038 65758
rect 22102 65694 22244 65758
rect 22032 65622 22244 65694
rect 22032 65558 22038 65622
rect 22102 65558 22244 65622
rect 22032 65552 22244 65558
rect 22440 65758 22652 65764
rect 22440 65694 22582 65758
rect 22646 65694 22652 65758
rect 22440 65622 22652 65694
rect 22440 65558 22446 65622
rect 22510 65558 22652 65622
rect 22440 65552 22652 65558
rect 27336 65552 27684 65764
rect 27608 65492 27684 65552
rect 20808 65350 21020 65356
rect 20808 65286 20950 65350
rect 21014 65286 21020 65350
rect 20808 65144 21020 65286
rect 21216 65350 21564 65356
rect 21216 65286 21358 65350
rect 21422 65286 21494 65350
rect 21558 65286 21564 65350
rect 21216 65280 21564 65286
rect 21216 65220 21428 65280
rect 21624 65220 21972 65356
rect 21216 65214 21972 65220
rect 21216 65150 21902 65214
rect 21966 65150 21972 65214
rect 21216 65144 21972 65150
rect 22032 65350 22244 65356
rect 22032 65286 22038 65350
rect 22102 65286 22244 65350
rect 22032 65214 22244 65286
rect 22032 65150 22174 65214
rect 22238 65150 22244 65214
rect 22032 65144 22244 65150
rect 22440 65350 22652 65356
rect 22440 65286 22446 65350
rect 22510 65286 22652 65350
rect 22440 65214 22652 65286
rect 27336 65280 27684 65492
rect 109344 65824 109556 66036
rect 114240 66166 114452 66172
rect 114240 66102 114246 66166
rect 114310 66102 114452 66166
rect 114240 66030 114452 66102
rect 114240 65966 114382 66030
rect 114446 65966 114452 66030
rect 114240 65960 114452 65966
rect 114648 66166 114860 66172
rect 114648 66102 114654 66166
rect 114718 66102 114860 66166
rect 114648 66030 114860 66102
rect 114648 65966 114654 66030
rect 114718 65966 114860 66030
rect 114648 65960 114860 65966
rect 115056 66166 115268 66172
rect 115366 66166 115676 66172
rect 115056 66102 115062 66166
rect 115126 66102 115268 66166
rect 115328 66102 115334 66166
rect 115398 66102 115676 66166
rect 115056 65960 115268 66102
rect 115366 66096 115676 66102
rect 115464 66030 115676 66096
rect 115464 65966 115606 66030
rect 115670 65966 115676 66030
rect 115464 65960 115676 65966
rect 115872 66166 116084 66172
rect 115872 66102 116014 66166
rect 116078 66102 116084 66166
rect 115872 66030 116084 66102
rect 115872 65966 116014 66030
rect 116078 65966 116084 66030
rect 115872 65960 116084 65966
rect 134776 65928 134988 66036
rect 134776 65872 134844 65928
rect 134900 65900 134988 65928
rect 134900 65894 135396 65900
rect 134900 65872 135326 65894
rect 134776 65830 135326 65872
rect 135390 65830 135396 65894
rect 134776 65824 135396 65830
rect 109344 65764 109420 65824
rect 134776 65764 134852 65824
rect 109344 65552 109556 65764
rect 114240 65758 114452 65764
rect 114240 65694 114382 65758
rect 114446 65694 114452 65758
rect 114240 65622 114452 65694
rect 114240 65558 114382 65622
rect 114446 65558 114452 65622
rect 114240 65552 114452 65558
rect 114648 65758 114860 65764
rect 114648 65694 114654 65758
rect 114718 65694 114860 65758
rect 114648 65622 114860 65694
rect 114648 65558 114654 65622
rect 114718 65558 114860 65622
rect 114648 65552 114860 65558
rect 115056 65758 115676 65764
rect 115056 65694 115606 65758
rect 115670 65694 115676 65758
rect 115056 65688 115676 65694
rect 115056 65628 115268 65688
rect 115056 65622 115404 65628
rect 115056 65558 115198 65622
rect 115262 65558 115334 65622
rect 115398 65558 115404 65622
rect 115056 65552 115404 65558
rect 115464 65552 115676 65688
rect 115872 65758 116084 65764
rect 115872 65694 116014 65758
rect 116078 65694 116084 65758
rect 115872 65622 116084 65694
rect 115872 65558 115878 65622
rect 115942 65558 116084 65622
rect 115872 65552 116084 65558
rect 132600 65688 134852 65764
rect 132600 65552 132812 65688
rect 133280 65552 133492 65688
rect 109344 65492 109420 65552
rect 109344 65280 109556 65492
rect 27472 65220 27548 65280
rect 109480 65220 109556 65280
rect 22440 65150 22446 65214
rect 22510 65150 22652 65214
rect 22440 65144 22652 65150
rect 20944 65084 21020 65144
rect 20808 65078 22108 65084
rect 20808 65014 22038 65078
rect 22102 65014 22108 65078
rect 20808 65008 22108 65014
rect 27336 65078 27684 65220
rect 27336 65014 27614 65078
rect 27678 65014 27684 65078
rect 27336 65008 27684 65014
rect 109344 65008 109556 65220
rect 114240 65350 114452 65356
rect 114240 65286 114382 65350
rect 114446 65286 114452 65350
rect 114240 65214 114452 65286
rect 114240 65150 114246 65214
rect 114310 65150 114452 65214
rect 114240 65144 114452 65150
rect 114648 65350 114860 65356
rect 114648 65286 114654 65350
rect 114718 65286 114860 65350
rect 114648 65214 114860 65286
rect 114648 65150 114654 65214
rect 114718 65150 114860 65214
rect 114648 65144 114860 65150
rect 115056 65350 115268 65356
rect 115366 65350 115676 65356
rect 115056 65286 115198 65350
rect 115262 65286 115268 65350
rect 115328 65286 115334 65350
rect 115398 65286 115676 65350
rect 115056 65214 115268 65286
rect 115366 65280 115676 65286
rect 115056 65150 115062 65214
rect 115126 65150 115268 65214
rect 115056 65144 115268 65150
rect 115464 65214 115676 65280
rect 115464 65150 115470 65214
rect 115534 65150 115676 65214
rect 115464 65144 115676 65150
rect 115872 65350 116084 65356
rect 115872 65286 115878 65350
rect 115942 65286 116084 65350
rect 115872 65144 116084 65286
rect 20808 64736 21020 65008
rect 27608 64948 27684 65008
rect 109480 64948 109556 65008
rect 115872 65084 115948 65144
rect 21216 64736 21428 64948
rect 21624 64942 21972 64948
rect 21624 64878 21902 64942
rect 21966 64878 21972 64942
rect 21624 64812 21972 64878
rect 21488 64736 21972 64812
rect 22032 64942 22244 64948
rect 22032 64878 22174 64942
rect 22238 64878 22244 64942
rect 22032 64806 22244 64878
rect 22032 64742 22174 64806
rect 22238 64742 22244 64806
rect 22032 64736 22244 64742
rect 22440 64942 22652 64948
rect 22440 64878 22446 64942
rect 22510 64878 22652 64942
rect 22440 64806 22652 64878
rect 22440 64742 22582 64806
rect 22646 64742 22652 64806
rect 22440 64736 22652 64742
rect 27336 64806 27684 64948
rect 27336 64742 27614 64806
rect 27678 64742 27684 64806
rect 20808 64676 20884 64736
rect 21216 64676 21292 64736
rect 21488 64676 21564 64736
rect 1768 64248 1980 64404
rect 1768 64192 1794 64248
rect 1850 64192 1980 64248
rect 1768 64132 1980 64192
rect 1224 64126 1980 64132
rect 1224 64062 1230 64126
rect 1294 64062 1980 64126
rect 1224 64056 1980 64062
rect 20808 64328 21020 64676
rect 21216 64600 21564 64676
rect 21216 64404 21428 64600
rect 21624 64404 21972 64676
rect 21216 64398 21972 64404
rect 21216 64334 21766 64398
rect 21830 64334 21972 64398
rect 21216 64328 21972 64334
rect 22032 64534 22244 64540
rect 22032 64470 22038 64534
rect 22102 64470 22174 64534
rect 22238 64470 22244 64534
rect 22032 64328 22244 64470
rect 22440 64534 22652 64540
rect 22440 64470 22582 64534
rect 22646 64470 22652 64534
rect 22440 64328 22652 64470
rect 27336 64534 27684 64742
rect 27336 64470 27342 64534
rect 27406 64470 27684 64534
rect 27336 64464 27684 64470
rect 109344 64806 109556 64948
rect 109344 64742 109350 64806
rect 109414 64742 109556 64806
rect 109344 64464 109556 64742
rect 114240 64942 114452 64948
rect 114240 64878 114246 64942
rect 114310 64878 114452 64942
rect 114240 64806 114452 64878
rect 114240 64742 114382 64806
rect 114446 64742 114452 64806
rect 114240 64736 114452 64742
rect 114648 64942 114860 64948
rect 114648 64878 114654 64942
rect 114718 64878 114860 64942
rect 114648 64806 114860 64878
rect 114648 64742 114654 64806
rect 114718 64742 114860 64806
rect 114648 64736 114860 64742
rect 115056 64942 115268 64948
rect 115056 64878 115062 64942
rect 115126 64878 115268 64942
rect 115056 64736 115268 64878
rect 115464 64942 115676 64948
rect 115464 64878 115470 64942
rect 115534 64878 115676 64942
rect 115464 64736 115676 64878
rect 115600 64676 115676 64736
rect 115056 64600 115676 64676
rect 114240 64534 114452 64540
rect 114240 64470 114382 64534
rect 114446 64470 114452 64534
rect 109344 64404 109420 64464
rect 20808 64268 20884 64328
rect 22032 64268 22108 64328
rect 22440 64268 22516 64328
rect 20808 64126 21020 64268
rect 20808 64062 20814 64126
rect 20878 64062 21020 64126
rect 20808 64056 21020 64062
rect 21216 63996 21428 64132
rect 21624 64126 21972 64132
rect 21624 64062 21766 64126
rect 21830 64062 21972 64126
rect 21216 63920 21564 63996
rect 21624 63920 21972 64062
rect 22032 63920 22244 64268
rect 21352 63860 21428 63920
rect 20808 63854 21020 63860
rect 20808 63790 20814 63854
rect 20878 63790 21020 63854
rect 20808 63718 21020 63790
rect 20808 63654 20814 63718
rect 20878 63654 21020 63718
rect 20808 63648 21020 63654
rect 21216 63648 21428 63860
rect 21488 63860 21564 63920
rect 21896 63860 21972 63920
rect 22168 63860 22244 63920
rect 21488 63784 21972 63860
rect 21624 63718 21972 63784
rect 21624 63654 21902 63718
rect 21966 63654 21972 63718
rect 21624 63648 21972 63654
rect 22032 63512 22244 63860
rect 22440 63920 22652 64268
rect 27336 64262 27684 64404
rect 27336 64198 27342 64262
rect 27406 64198 27614 64262
rect 27678 64198 27684 64262
rect 27336 63990 27684 64198
rect 109344 64398 109556 64404
rect 109344 64334 109350 64398
rect 109414 64334 109556 64398
rect 109344 64262 109556 64334
rect 114240 64328 114452 64470
rect 114376 64268 114452 64328
rect 109344 64198 109486 64262
rect 109550 64198 109556 64262
rect 109344 63996 109556 64198
rect 109246 63990 109556 63996
rect 27336 63926 27614 63990
rect 27678 63926 27684 63990
rect 109208 63926 109214 63990
rect 109278 63926 109486 63990
rect 109550 63926 109556 63990
rect 22440 63860 22516 63920
rect 22440 63512 22652 63860
rect 27336 63854 27684 63926
rect 109246 63920 109556 63926
rect 27336 63790 27478 63854
rect 27542 63790 27684 63854
rect 27336 63784 27684 63790
rect 109344 63854 109556 63920
rect 109344 63790 109350 63854
rect 109414 63790 109556 63854
rect 109344 63784 109556 63790
rect 114240 63920 114452 64268
rect 114648 64534 114860 64540
rect 114648 64470 114654 64534
rect 114718 64470 114860 64534
rect 114648 64328 114860 64470
rect 115056 64404 115268 64600
rect 115056 64398 115404 64404
rect 115056 64334 115334 64398
rect 115398 64334 115404 64398
rect 115056 64328 115404 64334
rect 115464 64328 115676 64600
rect 115872 64736 116084 65084
rect 115872 64676 115948 64736
rect 115872 64328 116084 64676
rect 134640 64534 136076 64540
rect 134640 64470 136006 64534
rect 136070 64470 136076 64534
rect 134640 64464 136076 64470
rect 134640 64404 134716 64464
rect 114648 64268 114724 64328
rect 116008 64268 116084 64328
rect 114648 63920 114860 64268
rect 115056 63996 115268 64132
rect 115366 64126 115676 64132
rect 115328 64062 115334 64126
rect 115398 64062 115676 64126
rect 115366 64056 115676 64062
rect 115872 64126 116084 64268
rect 132600 64398 132812 64404
rect 132600 64334 132606 64398
rect 132670 64334 132812 64398
rect 132600 64268 132812 64334
rect 133280 64328 134716 64404
rect 133280 64268 133492 64328
rect 132600 64262 133492 64268
rect 132600 64198 133422 64262
rect 133486 64198 133492 64262
rect 132600 64192 133492 64198
rect 134776 64248 134988 64404
rect 134776 64192 134844 64248
rect 134900 64192 134988 64248
rect 115872 64062 116014 64126
rect 116078 64062 116084 64126
rect 115872 64056 116084 64062
rect 134776 64132 134988 64192
rect 134776 64126 135396 64132
rect 134776 64062 135326 64126
rect 135390 64062 135396 64126
rect 134776 64056 135396 64062
rect 115056 63920 115404 63996
rect 114240 63860 114316 63920
rect 114648 63860 114724 63920
rect 115056 63860 115132 63920
rect 115328 63860 115404 63920
rect 115464 63920 115676 64056
rect 115464 63860 115540 63920
rect 22032 63452 22108 63512
rect 22576 63452 22652 63512
rect 20808 63446 21020 63452
rect 20808 63382 20814 63446
rect 20878 63382 21020 63446
rect 20808 63310 21020 63382
rect 20808 63246 20814 63310
rect 20878 63246 21020 63310
rect 20808 63240 21020 63246
rect 21216 63316 21428 63452
rect 21624 63446 21972 63452
rect 21624 63382 21902 63446
rect 21966 63382 21972 63446
rect 21624 63316 21972 63382
rect 21216 63240 21972 63316
rect 22032 63310 22244 63452
rect 22032 63246 22038 63310
rect 22102 63246 22244 63310
rect 22032 63240 22244 63246
rect 22440 63310 22652 63452
rect 22440 63246 22582 63310
rect 22646 63246 22652 63310
rect 22440 63240 22652 63246
rect 27336 63582 27684 63588
rect 27336 63518 27478 63582
rect 27542 63518 27684 63582
rect 27336 63240 27684 63518
rect 109208 63582 109556 63588
rect 109208 63518 109214 63582
rect 109278 63518 109350 63582
rect 109414 63518 109556 63582
rect 109208 63512 109556 63518
rect 114240 63512 114452 63860
rect 114648 63512 114860 63860
rect 115056 63648 115268 63860
rect 115328 63784 115676 63860
rect 115464 63718 115676 63784
rect 115464 63654 115470 63718
rect 115534 63654 115676 63718
rect 115464 63648 115676 63654
rect 115872 63854 116084 63860
rect 115872 63790 116014 63854
rect 116078 63790 116084 63854
rect 115872 63718 116084 63790
rect 115872 63654 115878 63718
rect 115942 63654 116084 63718
rect 115872 63648 116084 63654
rect 109344 63240 109556 63512
rect 114376 63452 114452 63512
rect 114784 63452 114860 63512
rect 114240 63310 114452 63452
rect 114240 63246 114246 63310
rect 114310 63246 114452 63310
rect 114240 63240 114452 63246
rect 114648 63310 114860 63452
rect 114648 63246 114790 63310
rect 114854 63246 114860 63310
rect 114648 63240 114860 63246
rect 21216 63180 21428 63240
rect 21216 63104 21564 63180
rect 21624 63104 21972 63240
rect 27608 63180 27684 63240
rect 109480 63180 109556 63240
rect 21352 63044 21428 63104
rect 20808 63038 21020 63044
rect 20808 62974 20814 63038
rect 20878 62974 21020 63038
rect 20808 62902 21020 62974
rect 20808 62838 20814 62902
rect 20878 62838 21020 62902
rect 20808 62832 21020 62838
rect 21216 62832 21428 63044
rect 21488 63044 21564 63104
rect 21488 62968 21972 63044
rect 21624 62902 21972 62968
rect 21624 62838 21766 62902
rect 21830 62838 21972 62902
rect 21624 62832 21972 62838
rect 22032 63038 22244 63044
rect 22032 62974 22038 63038
rect 22102 62974 22244 63038
rect 22032 62902 22244 62974
rect 22032 62838 22038 62902
rect 22102 62838 22244 62902
rect 22032 62832 22244 62838
rect 22440 63038 22652 63044
rect 22440 62974 22582 63038
rect 22646 62974 22652 63038
rect 22440 62902 22652 62974
rect 27336 62968 27684 63180
rect 109344 62968 109556 63180
rect 115056 63104 115268 63452
rect 115464 63446 115676 63452
rect 115464 63382 115470 63446
rect 115534 63382 115676 63446
rect 115464 63104 115676 63382
rect 115872 63446 116084 63452
rect 115872 63382 115878 63446
rect 115942 63382 116084 63446
rect 115872 63310 116084 63382
rect 115872 63246 116014 63310
rect 116078 63246 116084 63310
rect 115872 63240 116084 63246
rect 115056 63044 115132 63104
rect 115464 63044 115540 63104
rect 27608 62908 27684 62968
rect 109480 62908 109556 62968
rect 22440 62838 22446 62902
rect 22510 62838 22652 62902
rect 22440 62832 22652 62838
rect 1224 62630 1980 62636
rect 1224 62566 1230 62630
rect 1294 62568 1980 62630
rect 1294 62566 1794 62568
rect 1224 62560 1794 62566
rect 1768 62512 1794 62560
rect 1850 62512 1980 62568
rect 1768 62424 1980 62512
rect 20808 62630 21020 62636
rect 20808 62566 20814 62630
rect 20878 62566 21020 62630
rect 20808 62494 21020 62566
rect 20808 62430 20814 62494
rect 20878 62430 21020 62494
rect 20808 62424 21020 62430
rect 21216 62494 21428 62636
rect 21216 62430 21222 62494
rect 21286 62430 21428 62494
rect 21216 62424 21428 62430
rect 21624 62630 21972 62636
rect 21624 62566 21766 62630
rect 21830 62566 21972 62630
rect 21624 62494 21972 62566
rect 21624 62430 21630 62494
rect 21694 62430 21972 62494
rect 21624 62424 21972 62430
rect 22032 62630 22244 62636
rect 22032 62566 22038 62630
rect 22102 62566 22244 62630
rect 22032 62494 22244 62566
rect 22032 62430 22038 62494
rect 22102 62430 22244 62494
rect 22032 62424 22244 62430
rect 22440 62630 22652 62636
rect 22440 62566 22446 62630
rect 22510 62566 22652 62630
rect 22440 62494 22652 62566
rect 22440 62430 22582 62494
rect 22646 62430 22652 62494
rect 22440 62424 22652 62430
rect 27336 62424 27684 62908
rect 109344 62630 109556 62908
rect 114240 63038 114452 63044
rect 114240 62974 114246 63038
rect 114310 62974 114452 63038
rect 114240 62902 114452 62974
rect 114240 62838 114246 62902
rect 114310 62838 114452 62902
rect 114240 62832 114452 62838
rect 114648 63038 114860 63044
rect 114648 62974 114790 63038
rect 114854 62974 114860 63038
rect 114648 62902 114860 62974
rect 114648 62838 114654 62902
rect 114718 62838 114860 62902
rect 114648 62832 114860 62838
rect 115056 62902 115268 63044
rect 115056 62838 115062 62902
rect 115126 62838 115268 62902
rect 115056 62832 115268 62838
rect 115464 62902 115676 63044
rect 115464 62838 115470 62902
rect 115534 62838 115676 62902
rect 115464 62832 115676 62838
rect 115872 63038 116084 63044
rect 115872 62974 116014 63038
rect 116078 62974 116084 63038
rect 115872 62902 116084 62974
rect 115872 62838 115878 62902
rect 115942 62838 116084 62902
rect 115872 62832 116084 62838
rect 132600 62772 132812 62908
rect 133280 62772 133492 62908
rect 132600 62696 134852 62772
rect 134776 62636 134852 62696
rect 109344 62566 109350 62630
rect 109414 62566 109556 62630
rect 109344 62424 109556 62566
rect 114240 62630 114452 62636
rect 114240 62566 114246 62630
rect 114310 62566 114452 62630
rect 114240 62494 114452 62566
rect 114240 62430 114382 62494
rect 114446 62430 114452 62494
rect 114240 62424 114452 62430
rect 114648 62630 114860 62636
rect 114648 62566 114654 62630
rect 114718 62566 114860 62630
rect 114648 62494 114860 62566
rect 114648 62430 114790 62494
rect 114854 62430 114860 62494
rect 114648 62424 114860 62430
rect 115056 62630 115268 62636
rect 115056 62566 115062 62630
rect 115126 62566 115268 62630
rect 115056 62494 115268 62566
rect 115056 62430 115198 62494
rect 115262 62430 115268 62494
rect 115056 62424 115268 62430
rect 115464 62630 115676 62636
rect 115464 62566 115470 62630
rect 115534 62566 115676 62630
rect 115464 62424 115676 62566
rect 115872 62630 116084 62636
rect 115872 62566 115878 62630
rect 115942 62566 116084 62630
rect 115872 62494 116084 62566
rect 115872 62430 115878 62494
rect 115942 62430 116084 62494
rect 115872 62424 116084 62430
rect 134776 62568 134988 62636
rect 134776 62512 134844 62568
rect 134900 62512 134988 62568
rect 134776 62500 134988 62512
rect 134776 62494 135396 62500
rect 134776 62430 135326 62494
rect 135390 62430 135396 62494
rect 134776 62424 135396 62430
rect 27472 62364 27548 62424
rect 109344 62364 109420 62424
rect 115464 62364 115540 62424
rect 20808 62222 21020 62228
rect 20808 62158 20814 62222
rect 20878 62158 21020 62222
rect 20808 62086 21020 62158
rect 20808 62022 20950 62086
rect 21014 62022 21020 62086
rect 20808 62016 21020 62022
rect 21216 62222 21428 62228
rect 21216 62158 21222 62222
rect 21286 62158 21428 62222
rect 21216 62086 21428 62158
rect 21216 62022 21358 62086
rect 21422 62022 21428 62086
rect 21216 62016 21428 62022
rect 21624 62222 21972 62228
rect 21624 62158 21630 62222
rect 21694 62158 21972 62222
rect 21624 62016 21972 62158
rect 22032 62222 22244 62228
rect 22032 62158 22038 62222
rect 22102 62158 22244 62222
rect 22032 62086 22244 62158
rect 22032 62022 22174 62086
rect 22238 62022 22244 62086
rect 22032 62016 22244 62022
rect 22440 62222 22652 62228
rect 22440 62158 22582 62222
rect 22646 62158 22652 62222
rect 22440 62086 22652 62158
rect 22440 62022 22446 62086
rect 22510 62022 22652 62086
rect 22440 62016 22652 62022
rect 27336 62152 27684 62364
rect 109344 62358 109556 62364
rect 109344 62294 109350 62358
rect 109414 62294 109556 62358
rect 109344 62152 109556 62294
rect 115192 62288 115540 62364
rect 115192 62228 115268 62288
rect 114240 62222 114452 62228
rect 114240 62158 114382 62222
rect 114446 62158 114452 62222
rect 27336 62092 27412 62152
rect 109344 62092 109420 62152
rect 21624 61956 21700 62016
rect 21352 61880 21700 61956
rect 27336 61880 27684 62092
rect 109344 61880 109556 62092
rect 114240 62086 114452 62158
rect 114240 62022 114246 62086
rect 114310 62022 114452 62086
rect 114240 62016 114452 62022
rect 114648 62222 114860 62228
rect 114648 62158 114790 62222
rect 114854 62158 114860 62222
rect 114648 62086 114860 62158
rect 114648 62022 114654 62086
rect 114718 62022 114860 62086
rect 114648 62016 114860 62022
rect 115056 62222 115676 62228
rect 115056 62158 115198 62222
rect 115262 62158 115676 62222
rect 115056 62152 115676 62158
rect 115056 62016 115268 62152
rect 115464 62086 115676 62152
rect 115464 62022 115470 62086
rect 115534 62022 115676 62086
rect 115464 62016 115676 62022
rect 115872 62222 116084 62228
rect 115872 62158 115878 62222
rect 115942 62158 116084 62222
rect 115872 62086 116084 62158
rect 134092 62123 134158 62124
rect 115872 62022 116014 62086
rect 116078 62022 116084 62086
rect 134050 62059 134093 62123
rect 134157 62059 134200 62123
rect 134092 62058 134158 62059
rect 115872 62016 116084 62022
rect 21352 61820 21428 61880
rect 27608 61820 27684 61880
rect 109480 61820 109556 61880
rect 20808 61814 21020 61820
rect 20808 61750 20950 61814
rect 21014 61750 21020 61814
rect 20808 61678 21020 61750
rect 20808 61614 20950 61678
rect 21014 61614 21020 61678
rect 20808 61608 21020 61614
rect 21216 61814 21972 61820
rect 21216 61750 21358 61814
rect 21422 61750 21972 61814
rect 21216 61744 21972 61750
rect 21216 61608 21428 61744
rect 21624 61678 21972 61744
rect 21624 61614 21766 61678
rect 21830 61614 21972 61678
rect 21624 61608 21972 61614
rect 22032 61814 22244 61820
rect 22032 61750 22174 61814
rect 22238 61750 22244 61814
rect 22032 61678 22244 61750
rect 22032 61614 22038 61678
rect 22102 61614 22244 61678
rect 22032 61608 22244 61614
rect 22440 61814 22652 61820
rect 22440 61750 22446 61814
rect 22510 61750 22652 61814
rect 22440 61678 22652 61750
rect 22440 61614 22446 61678
rect 22510 61614 22652 61678
rect 22440 61608 22652 61614
rect 27336 61608 27684 61820
rect 109344 61608 109556 61820
rect 114240 61814 114452 61820
rect 114240 61750 114246 61814
rect 114310 61750 114452 61814
rect 114240 61678 114452 61750
rect 114240 61614 114246 61678
rect 114310 61614 114452 61678
rect 114240 61608 114452 61614
rect 114648 61814 114860 61820
rect 114648 61750 114654 61814
rect 114718 61750 114860 61814
rect 114648 61678 114860 61750
rect 114648 61614 114654 61678
rect 114718 61614 114860 61678
rect 114648 61608 114860 61614
rect 115056 61678 115268 61820
rect 115056 61614 115062 61678
rect 115126 61614 115268 61678
rect 115056 61608 115268 61614
rect 115464 61814 115676 61820
rect 115464 61750 115470 61814
rect 115534 61750 115676 61814
rect 115464 61678 115676 61750
rect 115464 61614 115606 61678
rect 115670 61614 115676 61678
rect 115464 61608 115676 61614
rect 115872 61814 116084 61820
rect 115872 61750 116014 61814
rect 116078 61750 116084 61814
rect 115872 61678 116084 61750
rect 115872 61614 115878 61678
rect 115942 61614 116084 61678
rect 115872 61608 116084 61614
rect 27472 61548 27548 61608
rect 109344 61548 109420 61608
rect 20808 61406 21020 61412
rect 20808 61342 20950 61406
rect 21014 61342 21020 61406
rect 20808 61200 21020 61342
rect 21216 61270 21428 61412
rect 21216 61206 21358 61270
rect 21422 61206 21428 61270
rect 21216 61200 21428 61206
rect 21624 61406 21972 61412
rect 21624 61342 21766 61406
rect 21830 61342 21972 61406
rect 21624 61200 21972 61342
rect 22032 61406 22244 61412
rect 22032 61342 22038 61406
rect 22102 61342 22244 61406
rect 22032 61270 22244 61342
rect 22032 61206 22174 61270
rect 22238 61206 22244 61270
rect 22032 61200 22244 61206
rect 22440 61406 22652 61412
rect 22440 61342 22446 61406
rect 22510 61342 22652 61406
rect 22440 61270 22652 61342
rect 27336 61336 27684 61548
rect 27608 61276 27684 61336
rect 22440 61206 22446 61270
rect 22510 61206 22652 61270
rect 22440 61200 22652 61206
rect 20944 61140 21020 61200
rect 21624 61140 21700 61200
rect 1224 60998 1980 61004
rect 1224 60934 1230 60998
rect 1294 60934 1980 60998
rect 1224 60928 1980 60934
rect 1768 60888 1980 60928
rect 1768 60832 1794 60888
rect 1850 60832 1980 60888
rect 1768 60792 1980 60832
rect 20808 60792 21020 61140
rect 21352 61064 21700 61140
rect 27336 61064 27684 61276
rect 109344 61336 109556 61548
rect 132600 61412 132812 61548
rect 133280 61542 133492 61548
rect 133280 61478 133422 61542
rect 133486 61478 133492 61542
rect 133280 61412 133492 61478
rect 114240 61406 114452 61412
rect 114240 61342 114246 61406
rect 114310 61342 114452 61406
rect 109344 61276 109420 61336
rect 109344 61134 109556 61276
rect 114240 61270 114452 61342
rect 114240 61206 114246 61270
rect 114310 61206 114452 61270
rect 114240 61200 114452 61206
rect 114648 61406 114860 61412
rect 114648 61342 114654 61406
rect 114718 61342 114860 61406
rect 114648 61270 114860 61342
rect 114648 61206 114654 61270
rect 114718 61206 114860 61270
rect 114648 61200 114860 61206
rect 115056 61406 115676 61412
rect 115056 61342 115062 61406
rect 115126 61342 115606 61406
rect 115670 61342 115676 61406
rect 115056 61336 115676 61342
rect 115056 61276 115268 61336
rect 115056 61270 115404 61276
rect 115056 61206 115334 61270
rect 115398 61206 115404 61270
rect 115056 61200 115404 61206
rect 115464 61200 115676 61336
rect 115872 61406 116084 61412
rect 115872 61342 115878 61406
rect 115942 61342 116084 61406
rect 115872 61200 116084 61342
rect 132600 61336 133492 61412
rect 109344 61070 109486 61134
rect 109550 61070 109556 61134
rect 109344 61064 109556 61070
rect 115872 61140 115948 61200
rect 21352 61004 21428 61064
rect 27472 61004 27548 61064
rect 109344 61004 109420 61064
rect 21216 60998 21972 61004
rect 21216 60934 21358 60998
rect 21422 60934 21972 60998
rect 21216 60928 21972 60934
rect 21216 60868 21428 60928
rect 21216 60792 21564 60868
rect 21624 60792 21972 60928
rect 22032 60998 22244 61004
rect 22032 60934 22174 60998
rect 22238 60934 22244 60998
rect 22032 60862 22244 60934
rect 22032 60798 22174 60862
rect 22238 60798 22244 60862
rect 22032 60792 22244 60798
rect 22440 60998 22652 61004
rect 22440 60934 22446 60998
rect 22510 60934 22652 60998
rect 22440 60862 22652 60934
rect 22440 60798 22582 60862
rect 22646 60798 22652 60862
rect 22440 60792 22652 60798
rect 20808 60732 20884 60792
rect 21352 60732 21428 60792
rect 20808 60384 21020 60732
rect 21216 60384 21428 60732
rect 21488 60732 21564 60792
rect 21488 60656 21972 60732
rect 21624 60454 21972 60656
rect 21624 60390 21902 60454
rect 21966 60390 21972 60454
rect 21624 60384 21972 60390
rect 22032 60590 22244 60596
rect 22032 60526 22174 60590
rect 22238 60526 22244 60590
rect 22032 60454 22244 60526
rect 22032 60390 22038 60454
rect 22102 60390 22244 60454
rect 22032 60384 22244 60390
rect 22440 60590 22652 60596
rect 22440 60526 22582 60590
rect 22646 60526 22652 60590
rect 22440 60454 22652 60526
rect 27336 60520 27684 61004
rect 109344 60862 109556 61004
rect 109344 60798 109486 60862
rect 109550 60798 109556 60862
rect 109344 60520 109556 60798
rect 114240 60998 114452 61004
rect 114240 60934 114246 60998
rect 114310 60934 114452 60998
rect 114240 60862 114452 60934
rect 114240 60798 114246 60862
rect 114310 60798 114452 60862
rect 114240 60792 114452 60798
rect 114648 60998 114860 61004
rect 114648 60934 114654 60998
rect 114718 60934 114860 60998
rect 114648 60862 114860 60934
rect 114648 60798 114654 60862
rect 114718 60798 114860 60862
rect 114648 60792 114860 60798
rect 115056 60792 115268 61004
rect 115366 60998 115676 61004
rect 115328 60934 115334 60998
rect 115398 60934 115676 60998
rect 115366 60928 115676 60934
rect 115464 60792 115676 60928
rect 115872 60792 116084 61140
rect 134776 60888 134988 61004
rect 134776 60832 134844 60888
rect 134900 60868 134988 60888
rect 134900 60862 135396 60868
rect 134900 60832 135326 60862
rect 134776 60798 135326 60832
rect 135390 60798 135396 60862
rect 134776 60792 135396 60798
rect 115056 60732 115132 60792
rect 115464 60732 115540 60792
rect 116008 60732 116084 60792
rect 114240 60590 114452 60596
rect 114240 60526 114246 60590
rect 114310 60526 114452 60590
rect 27472 60460 27548 60520
rect 109344 60460 109420 60520
rect 22440 60390 22446 60454
rect 22510 60390 22652 60454
rect 22440 60384 22652 60390
rect 20808 60324 20884 60384
rect 20808 60182 21020 60324
rect 27336 60248 27684 60460
rect 109344 60248 109556 60460
rect 114240 60454 114452 60526
rect 114240 60390 114382 60454
rect 114446 60390 114452 60454
rect 114240 60384 114452 60390
rect 114648 60590 114860 60596
rect 114648 60526 114654 60590
rect 114718 60526 114860 60590
rect 114648 60454 114860 60526
rect 114648 60390 114654 60454
rect 114718 60390 114860 60454
rect 114648 60384 114860 60390
rect 115056 60454 115268 60732
rect 115464 60460 115676 60732
rect 115366 60454 115676 60460
rect 115056 60390 115198 60454
rect 115262 60390 115268 60454
rect 115328 60390 115334 60454
rect 115398 60390 115676 60454
rect 115056 60384 115268 60390
rect 115366 60384 115676 60390
rect 115872 60384 116084 60732
rect 115872 60324 115948 60384
rect 27472 60188 27548 60248
rect 109344 60188 109420 60248
rect 20808 60118 20814 60182
rect 20878 60118 21020 60182
rect 20808 60112 21020 60118
rect 21216 59976 21428 60188
rect 21624 60182 21972 60188
rect 21624 60118 21902 60182
rect 21966 60118 21972 60182
rect 21624 59976 21972 60118
rect 22032 60182 22244 60188
rect 22032 60118 22038 60182
rect 22102 60118 22244 60182
rect 22032 59976 22244 60118
rect 22440 60182 22652 60188
rect 22440 60118 22446 60182
rect 22510 60118 22652 60182
rect 22440 59976 22652 60118
rect 21216 59916 21292 59976
rect 21624 59916 21700 59976
rect 22032 59916 22108 59976
rect 22440 59916 22516 59976
rect 20808 59910 21020 59916
rect 20808 59846 20814 59910
rect 20878 59846 21020 59910
rect 20808 59774 21020 59846
rect 20808 59710 20814 59774
rect 20878 59710 21020 59774
rect 20808 59704 21020 59710
rect 21216 59840 21972 59916
rect 21216 59704 21428 59840
rect 21624 59774 21972 59840
rect 21624 59710 21766 59774
rect 21830 59710 21972 59774
rect 21624 59704 21972 59710
rect 22032 59568 22244 59916
rect 22440 59568 22652 59916
rect 27336 59910 27684 60188
rect 27336 59846 27342 59910
rect 27406 59846 27684 59910
rect 27336 59840 27684 59846
rect 109344 59910 109556 60188
rect 114240 60182 114452 60188
rect 114240 60118 114382 60182
rect 114446 60118 114452 60182
rect 114240 59976 114452 60118
rect 114376 59916 114452 59976
rect 109344 59846 109486 59910
rect 109550 59846 109556 59910
rect 109344 59840 109556 59846
rect 22168 59508 22244 59568
rect 22576 59508 22652 59568
rect 20808 59502 21020 59508
rect 20808 59438 20814 59502
rect 20878 59438 21020 59502
rect 20808 59366 21020 59438
rect 20808 59302 20814 59366
rect 20878 59302 21020 59366
rect 20808 59296 21020 59302
rect 1224 59230 1980 59236
rect 1224 59166 1230 59230
rect 1294 59208 1980 59230
rect 1294 59166 1794 59208
rect 1224 59160 1794 59166
rect 1768 59152 1794 59160
rect 1850 59152 1980 59208
rect 1768 59024 1980 59152
rect 21216 59160 21428 59508
rect 21624 59502 21972 59508
rect 21624 59438 21766 59502
rect 21830 59438 21972 59502
rect 21624 59160 21972 59438
rect 22032 59366 22244 59508
rect 22032 59302 22038 59366
rect 22102 59302 22244 59366
rect 22032 59296 22244 59302
rect 22440 59366 22652 59508
rect 22440 59302 22446 59366
rect 22510 59302 22652 59366
rect 22440 59296 22652 59302
rect 27336 59638 27684 59644
rect 27336 59574 27342 59638
rect 27406 59574 27684 59638
rect 27336 59296 27684 59574
rect 109344 59638 109556 59644
rect 109344 59574 109486 59638
rect 109550 59574 109556 59638
rect 109344 59296 109556 59574
rect 114240 59568 114452 59916
rect 114648 60182 114860 60188
rect 114648 60118 114654 60182
rect 114718 60118 114860 60182
rect 114648 59976 114860 60118
rect 115056 60182 115404 60188
rect 115056 60118 115198 60182
rect 115262 60118 115334 60182
rect 115398 60118 115404 60182
rect 115056 60112 115404 60118
rect 115056 60052 115268 60112
rect 115464 60052 115676 60188
rect 115872 60182 116084 60324
rect 115872 60118 116014 60182
rect 116078 60118 116084 60182
rect 115872 60112 116084 60118
rect 115056 59976 115676 60052
rect 114648 59916 114724 59976
rect 115192 59916 115268 59976
rect 114648 59568 114860 59916
rect 115056 59704 115268 59916
rect 115464 59916 115540 59976
rect 115464 59774 115676 59916
rect 115464 59710 115470 59774
rect 115534 59710 115676 59774
rect 115464 59704 115676 59710
rect 115872 59910 116084 59916
rect 115872 59846 116014 59910
rect 116078 59846 116084 59910
rect 115872 59774 116084 59846
rect 115872 59710 116014 59774
rect 116078 59710 116084 59774
rect 115872 59704 116084 59710
rect 114240 59508 114316 59568
rect 114648 59508 114724 59568
rect 114240 59366 114452 59508
rect 114240 59302 114382 59366
rect 114446 59302 114452 59366
rect 114240 59296 114452 59302
rect 114648 59366 114860 59508
rect 114648 59302 114790 59366
rect 114854 59302 114860 59366
rect 114648 59296 114860 59302
rect 115056 59372 115268 59508
rect 115464 59502 115676 59508
rect 115464 59438 115470 59502
rect 115534 59438 115676 59502
rect 115464 59372 115676 59438
rect 115056 59296 115676 59372
rect 115872 59502 116084 59508
rect 115872 59438 116014 59502
rect 116078 59438 116084 59502
rect 115872 59366 116084 59438
rect 115872 59302 115878 59366
rect 115942 59302 116084 59366
rect 115872 59296 116084 59302
rect 27472 59236 27548 59296
rect 109344 59236 109420 59296
rect 21216 59100 21292 59160
rect 21896 59100 21972 59160
rect 20808 59094 21020 59100
rect 20808 59030 20814 59094
rect 20878 59030 21020 59094
rect 20808 58958 21020 59030
rect 20808 58894 20814 58958
rect 20878 58894 21020 58958
rect 20808 58888 21020 58894
rect 21216 58958 21428 59100
rect 21216 58894 21222 58958
rect 21286 58894 21428 58958
rect 21216 58888 21428 58894
rect 21624 58888 21972 59100
rect 22032 59094 22244 59100
rect 22032 59030 22038 59094
rect 22102 59030 22244 59094
rect 22032 58958 22244 59030
rect 22032 58894 22174 58958
rect 22238 58894 22244 58958
rect 22032 58888 22244 58894
rect 22440 59094 22652 59100
rect 22440 59030 22446 59094
rect 22510 59030 22652 59094
rect 22440 58958 22652 59030
rect 22440 58894 22446 58958
rect 22510 58894 22652 58958
rect 22440 58888 22652 58894
rect 27336 59024 27684 59236
rect 109344 59024 109556 59236
rect 115056 59160 115268 59296
rect 115464 59160 115676 59296
rect 115192 59100 115268 59160
rect 115600 59100 115676 59160
rect 134776 59230 135396 59236
rect 134776 59208 135326 59230
rect 134776 59152 134844 59208
rect 134900 59166 135326 59208
rect 135390 59166 135396 59230
rect 134900 59160 135396 59166
rect 134900 59152 134988 59160
rect 114240 59094 114452 59100
rect 114240 59030 114382 59094
rect 114446 59030 114452 59094
rect 27336 58964 27412 59024
rect 109344 58964 109420 59024
rect 21624 58828 21700 58888
rect 21352 58752 21700 58828
rect 21352 58692 21428 58752
rect 20808 58686 21020 58692
rect 20808 58622 20814 58686
rect 20878 58622 21020 58686
rect 20808 58550 21020 58622
rect 20808 58486 20814 58550
rect 20878 58486 21020 58550
rect 20808 58480 21020 58486
rect 21216 58686 21972 58692
rect 21216 58622 21222 58686
rect 21286 58622 21972 58686
rect 21216 58616 21972 58622
rect 21216 58550 21428 58616
rect 21216 58486 21358 58550
rect 21422 58486 21428 58550
rect 21216 58480 21428 58486
rect 21624 58550 21972 58616
rect 21624 58486 21766 58550
rect 21830 58486 21972 58550
rect 21624 58480 21972 58486
rect 22032 58686 22244 58692
rect 22032 58622 22174 58686
rect 22238 58622 22244 58686
rect 22032 58550 22244 58622
rect 22032 58486 22174 58550
rect 22238 58486 22244 58550
rect 22032 58480 22244 58486
rect 22440 58686 22652 58692
rect 22440 58622 22446 58686
rect 22510 58622 22652 58686
rect 22440 58550 22652 58622
rect 22440 58486 22446 58550
rect 22510 58486 22652 58550
rect 22440 58480 22652 58486
rect 27336 58686 27684 58964
rect 27336 58622 27614 58686
rect 27678 58622 27684 58686
rect 27336 58480 27684 58622
rect 109344 58686 109556 58964
rect 114240 58958 114452 59030
rect 114240 58894 114382 58958
rect 114446 58894 114452 58958
rect 114240 58888 114452 58894
rect 114648 59094 114860 59100
rect 114648 59030 114790 59094
rect 114854 59030 114860 59094
rect 114648 58958 114860 59030
rect 114648 58894 114790 58958
rect 114854 58894 114860 58958
rect 114648 58888 114860 58894
rect 115056 58888 115268 59100
rect 115464 58958 115676 59100
rect 115464 58894 115470 58958
rect 115534 58894 115676 58958
rect 115464 58888 115676 58894
rect 115872 59094 116084 59100
rect 115872 59030 115878 59094
rect 115942 59030 116084 59094
rect 115872 58958 116084 59030
rect 134776 59024 134988 59152
rect 115872 58894 115878 58958
rect 115942 58894 116084 58958
rect 115872 58888 116084 58894
rect 109344 58622 109486 58686
rect 109550 58622 109556 58686
rect 109344 58480 109556 58622
rect 114240 58686 114452 58692
rect 114240 58622 114382 58686
rect 114446 58622 114452 58686
rect 114240 58550 114452 58622
rect 114240 58486 114246 58550
rect 114310 58486 114452 58550
rect 114240 58480 114452 58486
rect 114648 58686 114860 58692
rect 114648 58622 114790 58686
rect 114854 58622 114860 58686
rect 114648 58550 114860 58622
rect 114648 58486 114790 58550
rect 114854 58486 114860 58550
rect 114648 58480 114860 58486
rect 115056 58550 115268 58692
rect 115464 58686 115676 58692
rect 115464 58622 115470 58686
rect 115534 58622 115676 58686
rect 115464 58556 115676 58622
rect 115366 58550 115676 58556
rect 115056 58486 115062 58550
rect 115126 58486 115268 58550
rect 115328 58486 115334 58550
rect 115398 58486 115676 58550
rect 115056 58480 115268 58486
rect 115366 58480 115676 58486
rect 115872 58686 116084 58692
rect 115872 58622 115878 58686
rect 115942 58622 116084 58686
rect 115872 58550 116084 58622
rect 115872 58486 116014 58550
rect 116078 58486 116084 58550
rect 115872 58480 116084 58486
rect 27472 58420 27548 58480
rect 109480 58420 109556 58480
rect 27336 58414 27684 58420
rect 27336 58350 27614 58414
rect 27678 58350 27684 58414
rect 20808 58278 21020 58284
rect 20808 58214 20814 58278
rect 20878 58214 21020 58278
rect 20808 58142 21020 58214
rect 20808 58078 20950 58142
rect 21014 58078 21020 58142
rect 20808 58072 21020 58078
rect 21216 58278 21428 58284
rect 21216 58214 21358 58278
rect 21422 58214 21428 58278
rect 21216 58072 21428 58214
rect 21624 58278 21972 58284
rect 21624 58214 21766 58278
rect 21830 58214 21972 58278
rect 21624 58148 21972 58214
rect 21526 58142 21972 58148
rect 21488 58078 21494 58142
rect 21558 58078 21972 58142
rect 21526 58072 21972 58078
rect 22032 58278 22244 58284
rect 22032 58214 22174 58278
rect 22238 58214 22244 58278
rect 22032 58142 22244 58214
rect 22032 58078 22038 58142
rect 22102 58078 22244 58142
rect 22032 58072 22244 58078
rect 22440 58278 22652 58284
rect 22440 58214 22446 58278
rect 22510 58214 22652 58278
rect 22440 58142 22652 58214
rect 22440 58078 22446 58142
rect 22510 58078 22652 58142
rect 22440 58072 22652 58078
rect 27336 58208 27684 58350
rect 109344 58414 109556 58420
rect 109344 58350 109486 58414
rect 109550 58350 109556 58414
rect 109344 58208 109556 58350
rect 114240 58278 114452 58284
rect 114240 58214 114246 58278
rect 114310 58214 114452 58278
rect 27336 58148 27412 58208
rect 109344 58148 109420 58208
rect 27336 57936 27684 58148
rect 109344 57936 109556 58148
rect 114240 58142 114452 58214
rect 114240 58078 114382 58142
rect 114446 58078 114452 58142
rect 114240 58072 114452 58078
rect 114648 58278 114860 58284
rect 114648 58214 114790 58278
rect 114854 58214 114860 58278
rect 114648 58142 114860 58214
rect 114648 58078 114790 58142
rect 114854 58078 114860 58142
rect 114648 58072 114860 58078
rect 115056 58278 115404 58284
rect 115056 58214 115062 58278
rect 115126 58214 115334 58278
rect 115398 58214 115404 58278
rect 115056 58208 115404 58214
rect 115056 58142 115268 58208
rect 115464 58148 115676 58284
rect 115366 58142 115676 58148
rect 115056 58078 115198 58142
rect 115262 58078 115268 58142
rect 115328 58078 115334 58142
rect 115398 58078 115676 58142
rect 115056 58072 115268 58078
rect 115366 58072 115676 58078
rect 115872 58278 116084 58284
rect 115872 58214 116014 58278
rect 116078 58214 116084 58278
rect 115872 58142 116084 58214
rect 115872 58078 115878 58142
rect 115942 58078 116084 58142
rect 115872 58072 116084 58078
rect 27472 57876 27548 57936
rect 109344 57876 109420 57936
rect 20808 57870 21020 57876
rect 20808 57806 20950 57870
rect 21014 57806 21020 57870
rect 20808 57734 21020 57806
rect 20808 57670 20814 57734
rect 20878 57670 21020 57734
rect 20808 57664 21020 57670
rect 21216 57870 21564 57876
rect 21216 57806 21494 57870
rect 21558 57806 21564 57870
rect 21216 57800 21564 57806
rect 21216 57740 21428 57800
rect 21624 57740 21972 57876
rect 21216 57664 21972 57740
rect 22032 57870 22244 57876
rect 22032 57806 22038 57870
rect 22102 57806 22244 57870
rect 22032 57734 22244 57806
rect 22032 57670 22174 57734
rect 22238 57670 22244 57734
rect 22032 57664 22244 57670
rect 22440 57870 22652 57876
rect 22440 57806 22446 57870
rect 22510 57806 22652 57870
rect 22440 57734 22652 57806
rect 22440 57670 22582 57734
rect 22646 57670 22652 57734
rect 22440 57664 22652 57670
rect 27336 57664 27684 57876
rect 109344 57664 109556 57876
rect 114240 57870 114452 57876
rect 114240 57806 114382 57870
rect 114446 57806 114452 57870
rect 114240 57734 114452 57806
rect 114240 57670 114246 57734
rect 114310 57670 114452 57734
rect 114240 57664 114452 57670
rect 114648 57870 114860 57876
rect 114648 57806 114790 57870
rect 114854 57806 114860 57870
rect 114648 57734 114860 57806
rect 114648 57670 114654 57734
rect 114718 57670 114860 57734
rect 114648 57664 114860 57670
rect 115056 57870 115404 57876
rect 115056 57806 115198 57870
rect 115262 57806 115334 57870
rect 115398 57806 115404 57870
rect 115056 57800 115404 57806
rect 115056 57740 115268 57800
rect 115464 57740 115676 57876
rect 115056 57734 115676 57740
rect 115056 57670 115606 57734
rect 115670 57670 115676 57734
rect 115056 57664 115676 57670
rect 115872 57870 116084 57876
rect 115872 57806 115878 57870
rect 115942 57806 116084 57870
rect 115872 57734 116084 57806
rect 115872 57670 116014 57734
rect 116078 57670 116084 57734
rect 115872 57664 116084 57670
rect 21624 57604 21700 57664
rect 27608 57604 27684 57664
rect 109480 57604 109556 57664
rect 1224 57598 1980 57604
rect 1224 57534 1230 57598
rect 1294 57534 1980 57598
rect 1224 57528 1980 57534
rect 1768 57472 1794 57528
rect 1850 57472 1980 57528
rect 1768 57392 1980 57472
rect 21488 57528 21700 57604
rect 21488 57468 21564 57528
rect 20808 57462 21020 57468
rect 20808 57398 20814 57462
rect 20878 57398 21020 57462
rect 20808 57256 21020 57398
rect 21216 57392 21564 57468
rect 21216 57326 21428 57392
rect 21216 57262 21222 57326
rect 21286 57262 21428 57326
rect 21216 57256 21428 57262
rect 21624 57326 21972 57468
rect 21624 57262 21766 57326
rect 21830 57262 21972 57326
rect 21624 57256 21972 57262
rect 22032 57462 22244 57468
rect 22032 57398 22174 57462
rect 22238 57398 22244 57462
rect 22032 57326 22244 57398
rect 22032 57262 22038 57326
rect 22102 57262 22244 57326
rect 22032 57256 22244 57262
rect 22440 57462 22652 57468
rect 22440 57398 22582 57462
rect 22646 57398 22652 57462
rect 22440 57326 22652 57398
rect 27336 57392 27684 57604
rect 109344 57392 109556 57604
rect 134776 57598 135396 57604
rect 134776 57534 135326 57598
rect 135390 57534 135396 57598
rect 134776 57528 135396 57534
rect 134776 57472 134844 57528
rect 134900 57472 134988 57528
rect 27472 57332 27548 57392
rect 109480 57332 109556 57392
rect 22440 57262 22446 57326
rect 22510 57262 22652 57326
rect 22440 57256 22652 57262
rect 20944 57196 21020 57256
rect 20808 56848 21020 57196
rect 27336 57120 27684 57332
rect 109344 57120 109556 57332
rect 114240 57462 114452 57468
rect 114240 57398 114246 57462
rect 114310 57398 114452 57462
rect 114240 57326 114452 57398
rect 114240 57262 114246 57326
rect 114310 57262 114452 57326
rect 114240 57256 114452 57262
rect 114648 57462 114860 57468
rect 114648 57398 114654 57462
rect 114718 57398 114860 57462
rect 114648 57326 114860 57398
rect 114648 57262 114654 57326
rect 114718 57262 114860 57326
rect 114648 57256 114860 57262
rect 115056 57326 115268 57468
rect 115056 57262 115198 57326
rect 115262 57262 115268 57326
rect 115056 57256 115268 57262
rect 115464 57462 115676 57468
rect 115464 57398 115606 57462
rect 115670 57398 115676 57462
rect 115464 57326 115676 57398
rect 115464 57262 115606 57326
rect 115670 57262 115676 57326
rect 115464 57256 115676 57262
rect 115872 57462 116084 57468
rect 115872 57398 116014 57462
rect 116078 57398 116084 57462
rect 115872 57256 116084 57398
rect 134776 57392 134988 57472
rect 116008 57196 116084 57256
rect 27336 57060 27412 57120
rect 109344 57060 109420 57120
rect 20944 56788 21020 56848
rect 20808 56440 21020 56788
rect 21216 57054 21428 57060
rect 21216 56990 21222 57054
rect 21286 56990 21428 57054
rect 21216 56848 21428 56990
rect 21624 57054 21972 57060
rect 21624 56990 21766 57054
rect 21830 56990 21972 57054
rect 21624 56848 21972 56990
rect 22032 57054 22244 57060
rect 22032 56990 22038 57054
rect 22102 56990 22244 57054
rect 22032 56918 22244 56990
rect 22032 56854 22038 56918
rect 22102 56854 22244 56918
rect 22032 56848 22244 56854
rect 22440 57054 22652 57060
rect 22440 56990 22446 57054
rect 22510 56990 22652 57054
rect 22440 56918 22652 56990
rect 22440 56854 22446 56918
rect 22510 56854 22652 56918
rect 22440 56848 22652 56854
rect 27336 56848 27684 57060
rect 109344 56848 109556 57060
rect 114240 57054 114452 57060
rect 114240 56990 114246 57054
rect 114310 56990 114452 57054
rect 114240 56918 114452 56990
rect 114240 56854 114246 56918
rect 114310 56854 114452 56918
rect 114240 56848 114452 56854
rect 114648 57054 114860 57060
rect 114648 56990 114654 57054
rect 114718 56990 114860 57054
rect 114648 56918 114860 56990
rect 114648 56854 114790 56918
rect 114854 56854 114860 56918
rect 114648 56848 114860 56854
rect 115056 57054 115268 57060
rect 115056 56990 115198 57054
rect 115262 56990 115268 57054
rect 115056 56924 115268 56990
rect 115464 57054 115676 57060
rect 115464 56990 115606 57054
rect 115670 56990 115676 57054
rect 115464 56924 115676 56990
rect 115056 56848 115676 56924
rect 115872 56848 116084 57196
rect 21216 56788 21292 56848
rect 21896 56788 21972 56848
rect 21216 56516 21428 56788
rect 21624 56516 21972 56788
rect 27462 56652 27560 56848
rect 109344 56652 109448 56848
rect 115192 56788 115268 56848
rect 115600 56788 115676 56848
rect 116008 56788 116084 56848
rect 21216 56510 21972 56516
rect 21216 56446 21358 56510
rect 21422 56446 21630 56510
rect 21694 56446 21972 56510
rect 21216 56440 21972 56446
rect 22032 56646 22244 56652
rect 22032 56582 22038 56646
rect 22102 56582 22244 56646
rect 22032 56510 22244 56582
rect 22032 56446 22174 56510
rect 22238 56446 22244 56510
rect 22032 56440 22244 56446
rect 22440 56646 22652 56652
rect 22440 56582 22446 56646
rect 22510 56582 22652 56646
rect 22440 56510 22652 56582
rect 27336 56576 27684 56652
rect 109344 56576 109556 56652
rect 114240 56646 114452 56652
rect 114240 56582 114246 56646
rect 114310 56582 114452 56646
rect 27472 56516 27548 56576
rect 109344 56516 109420 56576
rect 22440 56446 22446 56510
rect 22510 56446 22652 56510
rect 22440 56440 22652 56446
rect 20808 56380 20884 56440
rect 20808 56238 21020 56380
rect 27336 56304 27684 56516
rect 109344 56304 109556 56516
rect 114240 56510 114452 56582
rect 114240 56446 114246 56510
rect 114310 56446 114452 56510
rect 114240 56440 114452 56446
rect 114648 56646 114860 56652
rect 114648 56582 114790 56646
rect 114854 56582 114860 56646
rect 114648 56510 114860 56582
rect 114648 56446 114654 56510
rect 114718 56446 114860 56510
rect 114648 56440 114860 56446
rect 115056 56510 115268 56788
rect 115056 56446 115062 56510
rect 115126 56446 115268 56510
rect 115056 56440 115268 56446
rect 115464 56440 115676 56788
rect 115872 56440 116084 56788
rect 116008 56380 116084 56440
rect 27608 56244 27684 56304
rect 109480 56244 109556 56304
rect 20808 56174 20950 56238
rect 21014 56174 21020 56238
rect 20808 56168 21020 56174
rect 21216 56238 21428 56244
rect 21216 56174 21358 56238
rect 21422 56174 21428 56238
rect 21216 56032 21428 56174
rect 21624 56238 21972 56244
rect 21624 56174 21630 56238
rect 21694 56174 21972 56238
rect 21624 56032 21972 56174
rect 21216 55972 21292 56032
rect 21896 55972 21972 56032
rect 1224 55966 1980 55972
rect 1224 55902 1230 55966
rect 1294 55902 1980 55966
rect 1224 55896 1980 55902
rect 1768 55848 1980 55896
rect 1768 55792 1794 55848
rect 1850 55792 1980 55848
rect 1768 55760 1980 55792
rect 20808 55966 21020 55972
rect 20808 55902 20950 55966
rect 21014 55902 21020 55966
rect 20808 55830 21020 55902
rect 20808 55766 20814 55830
rect 20878 55766 21020 55830
rect 20808 55760 21020 55766
rect 21216 55760 21428 55972
rect 21624 55836 21972 55972
rect 21526 55830 21972 55836
rect 21488 55766 21494 55830
rect 21558 55766 21972 55830
rect 21526 55760 21972 55766
rect 22032 56238 22244 56244
rect 22032 56174 22174 56238
rect 22238 56174 22244 56238
rect 22032 56032 22244 56174
rect 22440 56238 22652 56244
rect 22440 56174 22446 56238
rect 22510 56174 22652 56238
rect 22440 56032 22652 56174
rect 22032 55972 22108 56032
rect 22440 55972 22516 56032
rect 22032 55624 22244 55972
rect 22440 55624 22652 55972
rect 27336 55966 27684 56244
rect 27336 55902 27478 55966
rect 27542 55902 27684 55966
rect 27336 55896 27684 55902
rect 109344 56102 109556 56244
rect 109344 56038 109350 56102
rect 109414 56038 109556 56102
rect 109344 55966 109556 56038
rect 114240 56238 114452 56244
rect 114240 56174 114246 56238
rect 114310 56174 114452 56238
rect 114240 56032 114452 56174
rect 114648 56238 114860 56244
rect 114648 56174 114654 56238
rect 114718 56174 114860 56238
rect 114648 56032 114860 56174
rect 115056 56238 115268 56244
rect 115056 56174 115062 56238
rect 115126 56174 115268 56238
rect 115056 56032 115268 56174
rect 115464 56108 115676 56244
rect 115872 56238 116084 56380
rect 115872 56174 116014 56238
rect 116078 56174 116084 56238
rect 115872 56168 116084 56174
rect 115366 56102 115676 56108
rect 115328 56038 115334 56102
rect 115398 56038 115676 56102
rect 115366 56032 115676 56038
rect 114376 55972 114452 56032
rect 114784 55972 114860 56032
rect 115192 55972 115268 56032
rect 109344 55902 109486 55966
rect 109550 55902 109556 55966
rect 109344 55896 109556 55902
rect 22032 55564 22108 55624
rect 22440 55564 22516 55624
rect 20808 55558 21020 55564
rect 20808 55494 20814 55558
rect 20878 55494 21020 55558
rect 20808 55422 21020 55494
rect 20808 55358 20950 55422
rect 21014 55358 21020 55422
rect 20808 55352 21020 55358
rect 21216 55558 21564 55564
rect 21216 55494 21494 55558
rect 21558 55494 21564 55558
rect 21216 55488 21564 55494
rect 21216 55428 21428 55488
rect 21624 55428 21972 55564
rect 21216 55352 21972 55428
rect 21216 55216 21428 55352
rect 21624 55216 21972 55352
rect 22032 55216 22244 55564
rect 22440 55216 22652 55564
rect 27336 55558 27684 55700
rect 27336 55494 27478 55558
rect 27542 55494 27614 55558
rect 27678 55494 27684 55558
rect 27336 55286 27684 55494
rect 27336 55222 27614 55286
rect 27678 55222 27684 55286
rect 21216 55156 21292 55216
rect 21624 55156 21700 55216
rect 22032 55156 22108 55216
rect 22440 55156 22516 55216
rect 20808 55150 21020 55156
rect 20808 55086 20950 55150
rect 21014 55086 21020 55150
rect 20808 55014 21020 55086
rect 20808 54950 20814 55014
rect 20878 54950 21020 55014
rect 20808 54944 21020 54950
rect 21216 54944 21428 55156
rect 21624 55014 21972 55156
rect 21624 54950 21630 55014
rect 21694 54950 21972 55014
rect 21624 54944 21972 54950
rect 22032 55014 22244 55156
rect 22032 54950 22038 55014
rect 22102 54950 22244 55014
rect 22032 54944 22244 54950
rect 22440 55014 22652 55156
rect 27336 55080 27684 55222
rect 109344 55694 109556 55700
rect 109344 55630 109350 55694
rect 109414 55630 109486 55694
rect 109550 55630 109556 55694
rect 109344 55558 109556 55630
rect 114240 55624 114452 55972
rect 114376 55564 114452 55624
rect 109344 55494 109486 55558
rect 109550 55494 109556 55558
rect 109344 55286 109556 55494
rect 109344 55222 109486 55286
rect 109550 55222 109556 55286
rect 109344 55080 109556 55222
rect 27608 55020 27684 55080
rect 109480 55020 109556 55080
rect 22440 54950 22446 55014
rect 22510 54950 22652 55014
rect 22440 54944 22652 54950
rect 20808 54742 21020 54748
rect 20808 54678 20814 54742
rect 20878 54678 21020 54742
rect 20808 54606 21020 54678
rect 20808 54542 20950 54606
rect 21014 54542 21020 54606
rect 20808 54536 21020 54542
rect 21216 54606 21428 54748
rect 21624 54742 21972 54748
rect 21624 54678 21630 54742
rect 21694 54678 21972 54742
rect 21624 54612 21972 54678
rect 21526 54606 21972 54612
rect 21216 54542 21358 54606
rect 21422 54542 21428 54606
rect 21488 54542 21494 54606
rect 21558 54542 21972 54606
rect 21216 54536 21428 54542
rect 21526 54536 21972 54542
rect 22032 54742 22244 54748
rect 22032 54678 22038 54742
rect 22102 54678 22244 54742
rect 22032 54606 22244 54678
rect 22032 54542 22174 54606
rect 22238 54542 22244 54606
rect 22032 54536 22244 54542
rect 22440 54742 22652 54748
rect 22440 54678 22446 54742
rect 22510 54678 22652 54742
rect 22440 54606 22652 54678
rect 22440 54542 22582 54606
rect 22646 54542 22652 54606
rect 22440 54536 22652 54542
rect 27336 54536 27684 55020
rect 27608 54476 27684 54536
rect 20808 54334 21020 54340
rect 20808 54270 20950 54334
rect 21014 54270 21020 54334
rect 1224 54198 1980 54204
rect 1224 54134 1230 54198
rect 1294 54168 1980 54198
rect 1294 54134 1794 54168
rect 1224 54128 1794 54134
rect 1768 54112 1794 54128
rect 1850 54112 1980 54168
rect 20808 54198 21020 54270
rect 20808 54134 20814 54198
rect 20878 54134 21020 54198
rect 20808 54128 21020 54134
rect 21216 54334 21564 54340
rect 21216 54270 21358 54334
rect 21422 54270 21494 54334
rect 21558 54270 21564 54334
rect 21216 54264 21564 54270
rect 21216 54204 21428 54264
rect 21624 54204 21972 54340
rect 21216 54198 21972 54204
rect 21216 54134 21766 54198
rect 21830 54134 21972 54198
rect 21216 54128 21972 54134
rect 22032 54334 22244 54340
rect 22032 54270 22174 54334
rect 22238 54270 22244 54334
rect 22032 54198 22244 54270
rect 22032 54134 22174 54198
rect 22238 54134 22244 54198
rect 22032 54128 22244 54134
rect 22440 54334 22652 54340
rect 22440 54270 22582 54334
rect 22646 54270 22652 54334
rect 22440 54198 22652 54270
rect 27336 54264 27684 54476
rect 109344 54536 109556 55020
rect 114240 55216 114452 55564
rect 114648 55624 114860 55972
rect 115056 55966 115676 55972
rect 115056 55902 115198 55966
rect 115262 55902 115676 55966
rect 115056 55896 115676 55902
rect 115056 55836 115268 55896
rect 115056 55830 115404 55836
rect 115056 55766 115334 55830
rect 115398 55766 115404 55830
rect 115056 55760 115404 55766
rect 115464 55760 115676 55896
rect 115872 55966 116084 55972
rect 115872 55902 116014 55966
rect 116078 55902 116084 55966
rect 115872 55830 116084 55902
rect 115872 55766 116014 55830
rect 116078 55766 116084 55830
rect 115872 55760 116084 55766
rect 134776 55966 135396 55972
rect 134776 55902 135326 55966
rect 135390 55902 135396 55966
rect 134776 55896 135396 55902
rect 134776 55848 134988 55896
rect 134776 55792 134844 55848
rect 134900 55792 134988 55848
rect 134776 55760 134988 55792
rect 114648 55564 114724 55624
rect 114648 55216 114860 55564
rect 115056 55216 115268 55564
rect 115366 55558 115676 55564
rect 115328 55494 115334 55558
rect 115398 55494 115676 55558
rect 115366 55488 115676 55494
rect 115464 55216 115676 55488
rect 115872 55558 116084 55564
rect 115872 55494 116014 55558
rect 116078 55494 116084 55558
rect 115872 55422 116084 55494
rect 115872 55358 116014 55422
rect 116078 55358 116084 55422
rect 115872 55352 116084 55358
rect 114240 55156 114316 55216
rect 114648 55156 114724 55216
rect 115056 55156 115132 55216
rect 115600 55156 115676 55216
rect 114240 55014 114452 55156
rect 114240 54950 114382 55014
rect 114446 54950 114452 55014
rect 114240 54944 114452 54950
rect 114648 55014 114860 55156
rect 114648 54950 114790 55014
rect 114854 54950 114860 55014
rect 114648 54944 114860 54950
rect 115056 55014 115268 55156
rect 115464 55020 115676 55156
rect 115366 55014 115676 55020
rect 115056 54950 115198 55014
rect 115262 54950 115268 55014
rect 115328 54950 115334 55014
rect 115398 54950 115676 55014
rect 115056 54944 115268 54950
rect 115366 54944 115676 54950
rect 115872 55150 116084 55156
rect 115872 55086 116014 55150
rect 116078 55086 116084 55150
rect 115872 55014 116084 55086
rect 115872 54950 115878 55014
rect 115942 54950 116084 55014
rect 115872 54944 116084 54950
rect 114240 54742 114452 54748
rect 114240 54678 114382 54742
rect 114446 54678 114452 54742
rect 114240 54606 114452 54678
rect 114240 54542 114246 54606
rect 114310 54542 114452 54606
rect 114240 54536 114452 54542
rect 114648 54742 114860 54748
rect 114648 54678 114790 54742
rect 114854 54678 114860 54742
rect 114648 54606 114860 54678
rect 114648 54542 114790 54606
rect 114854 54542 114860 54606
rect 114648 54536 114860 54542
rect 115056 54742 115404 54748
rect 115056 54678 115198 54742
rect 115262 54678 115334 54742
rect 115398 54678 115404 54742
rect 115056 54672 115404 54678
rect 115056 54612 115268 54672
rect 115464 54612 115676 54748
rect 115056 54606 115676 54612
rect 115056 54542 115470 54606
rect 115534 54542 115676 54606
rect 115056 54536 115676 54542
rect 115872 54742 116084 54748
rect 115872 54678 115878 54742
rect 115942 54678 116084 54742
rect 115872 54606 116084 54678
rect 115872 54542 116014 54606
rect 116078 54542 116084 54606
rect 115872 54536 116084 54542
rect 109344 54476 109420 54536
rect 109344 54264 109556 54476
rect 27608 54204 27684 54264
rect 109480 54204 109556 54264
rect 22440 54134 22446 54198
rect 22510 54134 22652 54198
rect 22440 54128 22652 54134
rect 1768 53992 1980 54112
rect 27336 53992 27684 54204
rect 109344 53992 109556 54204
rect 114240 54334 114452 54340
rect 114240 54270 114246 54334
rect 114310 54270 114452 54334
rect 114240 54198 114452 54270
rect 114240 54134 114382 54198
rect 114446 54134 114452 54198
rect 114240 54128 114452 54134
rect 114648 54334 114860 54340
rect 114648 54270 114790 54334
rect 114854 54270 114860 54334
rect 114648 54198 114860 54270
rect 114648 54134 114790 54198
rect 114854 54134 114860 54198
rect 114648 54128 114860 54134
rect 115056 54198 115268 54340
rect 115464 54334 115676 54340
rect 115464 54270 115470 54334
rect 115534 54270 115676 54334
rect 115464 54204 115676 54270
rect 115366 54198 115676 54204
rect 115056 54134 115198 54198
rect 115262 54134 115268 54198
rect 115328 54134 115334 54198
rect 115398 54134 115676 54198
rect 115056 54128 115268 54134
rect 115366 54128 115676 54134
rect 115872 54334 116084 54340
rect 115872 54270 116014 54334
rect 116078 54270 116084 54334
rect 115872 54198 116084 54270
rect 115872 54134 116014 54198
rect 116078 54134 116084 54198
rect 115872 54128 116084 54134
rect 134776 54168 134988 54204
rect 134776 54112 134844 54168
rect 134900 54112 134988 54168
rect 134776 54068 134988 54112
rect 134776 54062 135396 54068
rect 134776 53998 135326 54062
rect 135390 53998 135396 54062
rect 134776 53992 135396 53998
rect 27336 53932 27412 53992
rect 109344 53932 109420 53992
rect 20808 53926 21020 53932
rect 20808 53862 20814 53926
rect 20878 53862 21020 53926
rect 20808 53790 21020 53862
rect 20808 53726 20814 53790
rect 20878 53726 21020 53790
rect 20808 53720 21020 53726
rect 21216 53926 21972 53932
rect 21216 53862 21766 53926
rect 21830 53862 21972 53926
rect 21216 53856 21972 53862
rect 21216 53720 21428 53856
rect 21624 53790 21972 53856
rect 21624 53726 21630 53790
rect 21694 53726 21972 53790
rect 21624 53720 21972 53726
rect 22032 53926 22244 53932
rect 22032 53862 22174 53926
rect 22238 53862 22244 53926
rect 22032 53790 22244 53862
rect 22032 53726 22038 53790
rect 22102 53726 22244 53790
rect 22032 53720 22244 53726
rect 22440 53926 22652 53932
rect 22440 53862 22446 53926
rect 22510 53862 22652 53926
rect 22440 53790 22652 53862
rect 22440 53726 22446 53790
rect 22510 53726 22652 53790
rect 22440 53720 22652 53726
rect 27336 53720 27684 53932
rect 109344 53720 109556 53932
rect 114240 53926 114452 53932
rect 114240 53862 114382 53926
rect 114446 53862 114452 53926
rect 114240 53790 114452 53862
rect 114240 53726 114382 53790
rect 114446 53726 114452 53790
rect 114240 53720 114452 53726
rect 114648 53926 114860 53932
rect 114648 53862 114790 53926
rect 114854 53862 114860 53926
rect 114648 53790 114860 53862
rect 114648 53726 114790 53790
rect 114854 53726 114860 53790
rect 114648 53720 114860 53726
rect 115056 53926 115404 53932
rect 115056 53862 115198 53926
rect 115262 53862 115334 53926
rect 115398 53862 115404 53926
rect 115056 53856 115404 53862
rect 115056 53796 115268 53856
rect 115464 53796 115676 53932
rect 115056 53720 115676 53796
rect 115872 53926 116084 53932
rect 115872 53862 116014 53926
rect 116078 53862 116084 53926
rect 115872 53790 116084 53862
rect 115872 53726 115878 53790
rect 115942 53726 116084 53790
rect 115872 53720 116084 53726
rect 27336 53660 27412 53720
rect 109344 53660 109420 53720
rect 115464 53660 115540 53720
rect 20808 53518 21020 53524
rect 20808 53454 20814 53518
rect 20878 53454 21020 53518
rect 20808 53312 21020 53454
rect 21216 53518 21972 53524
rect 21216 53454 21630 53518
rect 21694 53454 21972 53518
rect 21216 53448 21972 53454
rect 21216 53388 21428 53448
rect 21216 53382 21564 53388
rect 21216 53318 21358 53382
rect 21422 53318 21494 53382
rect 21558 53318 21564 53382
rect 21216 53312 21564 53318
rect 21624 53312 21972 53448
rect 22032 53518 22244 53524
rect 22032 53454 22038 53518
rect 22102 53454 22244 53518
rect 22032 53382 22244 53454
rect 22032 53318 22174 53382
rect 22238 53318 22244 53382
rect 22032 53312 22244 53318
rect 22440 53518 22652 53524
rect 22440 53454 22446 53518
rect 22510 53454 22652 53518
rect 22440 53382 22652 53454
rect 22440 53318 22446 53382
rect 22510 53318 22652 53382
rect 22440 53312 22652 53318
rect 27336 53448 27684 53660
rect 109344 53448 109556 53660
rect 115192 53584 115540 53660
rect 115192 53524 115268 53584
rect 27336 53388 27412 53448
rect 109480 53388 109556 53448
rect 20944 53252 21020 53312
rect 20808 52974 21020 53252
rect 27336 53176 27684 53388
rect 109344 53176 109556 53388
rect 114240 53518 114452 53524
rect 114240 53454 114382 53518
rect 114446 53454 114452 53518
rect 114240 53382 114452 53454
rect 114240 53318 114246 53382
rect 114310 53318 114452 53382
rect 114240 53312 114452 53318
rect 114648 53518 114860 53524
rect 114648 53454 114790 53518
rect 114854 53454 114860 53518
rect 114648 53382 114860 53454
rect 114648 53318 114654 53382
rect 114718 53318 114860 53382
rect 114648 53312 114860 53318
rect 115056 53448 115676 53524
rect 115056 53312 115268 53448
rect 115464 53382 115676 53448
rect 115464 53318 115470 53382
rect 115534 53318 115676 53382
rect 115464 53312 115676 53318
rect 115872 53518 116084 53524
rect 115872 53454 115878 53518
rect 115942 53454 116084 53518
rect 115872 53312 116084 53454
rect 116008 53252 116084 53312
rect 27608 53116 27684 53176
rect 109480 53116 109556 53176
rect 20808 52910 20950 52974
rect 21014 52910 21020 52974
rect 20808 52904 21020 52910
rect 21216 53110 21428 53116
rect 21526 53110 21972 53116
rect 21216 53046 21358 53110
rect 21422 53046 21428 53110
rect 21488 53046 21494 53110
rect 21558 53046 21972 53110
rect 21216 52974 21428 53046
rect 21526 53040 21972 53046
rect 21216 52910 21222 52974
rect 21286 52910 21428 52974
rect 21216 52904 21428 52910
rect 21624 52974 21972 53040
rect 21624 52910 21766 52974
rect 21830 52910 21972 52974
rect 21624 52904 21972 52910
rect 22032 53110 22244 53116
rect 22032 53046 22174 53110
rect 22238 53046 22244 53110
rect 22032 52974 22244 53046
rect 22032 52910 22174 52974
rect 22238 52910 22244 52974
rect 22032 52904 22244 52910
rect 22440 53110 22652 53116
rect 22440 53046 22446 53110
rect 22510 53046 22652 53110
rect 22440 52974 22652 53046
rect 22440 52910 22582 52974
rect 22646 52910 22652 52974
rect 22440 52904 22652 52910
rect 27336 52904 27684 53116
rect 109344 52904 109556 53116
rect 114240 53110 114452 53116
rect 114240 53046 114246 53110
rect 114310 53046 114452 53110
rect 114240 52974 114452 53046
rect 114240 52910 114246 52974
rect 114310 52910 114452 52974
rect 114240 52904 114452 52910
rect 114648 53110 114860 53116
rect 114648 53046 114654 53110
rect 114718 53046 114860 53110
rect 114648 52974 114860 53046
rect 114648 52910 114790 52974
rect 114854 52910 114860 52974
rect 114648 52904 114860 52910
rect 115056 52974 115268 53116
rect 115056 52910 115198 52974
rect 115262 52910 115268 52974
rect 115056 52904 115268 52910
rect 115464 53110 115676 53116
rect 115464 53046 115470 53110
rect 115534 53046 115676 53110
rect 115464 52974 115676 53046
rect 115464 52910 115606 52974
rect 115670 52910 115676 52974
rect 115464 52904 115676 52910
rect 115872 52974 116084 53252
rect 115872 52910 115878 52974
rect 115942 52910 116084 52974
rect 115872 52904 116084 52910
rect 27336 52844 27412 52904
rect 109480 52844 109556 52904
rect 20808 52702 21020 52708
rect 20808 52638 20950 52702
rect 21014 52638 21020 52702
rect 1224 52566 1980 52572
rect 1224 52502 1230 52566
rect 1294 52502 1980 52566
rect 1224 52496 1980 52502
rect 20808 52496 21020 52638
rect 21216 52702 21428 52708
rect 21216 52638 21222 52702
rect 21286 52638 21428 52702
rect 21216 52496 21428 52638
rect 21624 52702 21972 52708
rect 21624 52638 21766 52702
rect 21830 52638 21972 52702
rect 21624 52496 21972 52638
rect 22032 52702 22244 52708
rect 22032 52638 22174 52702
rect 22238 52638 22244 52702
rect 22032 52566 22244 52638
rect 22032 52502 22174 52566
rect 22238 52502 22244 52566
rect 22032 52496 22244 52502
rect 22440 52702 22652 52708
rect 22440 52638 22582 52702
rect 22646 52638 22652 52702
rect 22440 52566 22652 52638
rect 27336 52632 27684 52844
rect 27608 52572 27684 52632
rect 22440 52502 22446 52566
rect 22510 52502 22652 52566
rect 22440 52496 22652 52502
rect 1768 52488 1980 52496
rect 1768 52432 1794 52488
rect 1850 52432 1980 52488
rect 20944 52436 21020 52496
rect 21624 52436 21700 52496
rect 1768 52360 1980 52432
rect 20808 52294 21020 52436
rect 21352 52360 21700 52436
rect 27336 52430 27684 52572
rect 27336 52366 27478 52430
rect 27542 52366 27684 52430
rect 27336 52360 27684 52366
rect 109344 52632 109556 52844
rect 114240 52702 114452 52708
rect 114240 52638 114246 52702
rect 114310 52638 114452 52702
rect 109344 52572 109420 52632
rect 109344 52360 109556 52572
rect 114240 52566 114452 52638
rect 114240 52502 114382 52566
rect 114446 52502 114452 52566
rect 114240 52496 114452 52502
rect 114648 52702 114860 52708
rect 114648 52638 114790 52702
rect 114854 52638 114860 52702
rect 114648 52566 114860 52638
rect 114648 52502 114790 52566
rect 114854 52502 114860 52566
rect 114648 52496 114860 52502
rect 115056 52702 115268 52708
rect 115056 52638 115198 52702
rect 115262 52638 115268 52702
rect 115056 52572 115268 52638
rect 115464 52702 115676 52708
rect 115464 52638 115606 52702
rect 115670 52638 115676 52702
rect 115464 52572 115676 52638
rect 115056 52566 115676 52572
rect 115056 52502 115198 52566
rect 115262 52502 115676 52566
rect 115056 52496 115676 52502
rect 115872 52702 116084 52708
rect 115872 52638 115878 52702
rect 115942 52638 116084 52702
rect 115872 52496 116084 52638
rect 115192 52436 115268 52496
rect 115872 52436 115948 52496
rect 134776 52488 134988 52572
rect 115192 52360 115540 52436
rect 21352 52300 21428 52360
rect 27472 52300 27548 52360
rect 109480 52300 109556 52360
rect 115464 52300 115540 52360
rect 20808 52230 20814 52294
rect 20878 52230 21020 52294
rect 20808 52224 21020 52230
rect 21216 52224 21972 52300
rect 21216 52164 21428 52224
rect 21216 52088 21564 52164
rect 21624 52088 21972 52224
rect 22032 52294 22244 52300
rect 22032 52230 22174 52294
rect 22238 52230 22244 52294
rect 22032 52158 22244 52230
rect 22032 52094 22174 52158
rect 22238 52094 22244 52158
rect 22032 52088 22244 52094
rect 22440 52294 22652 52300
rect 22440 52230 22446 52294
rect 22510 52230 22652 52294
rect 22440 52158 22652 52230
rect 22440 52094 22582 52158
rect 22646 52094 22652 52158
rect 22440 52088 22652 52094
rect 27336 52158 27684 52300
rect 27336 52094 27478 52158
rect 27542 52094 27684 52158
rect 21352 52028 21428 52088
rect 20808 52022 21020 52028
rect 20808 51958 20814 52022
rect 20878 51958 21020 52022
rect 20808 51680 21020 51958
rect 21216 51680 21428 52028
rect 21488 52028 21564 52088
rect 21488 51952 21972 52028
rect 21624 51750 21972 51952
rect 21624 51686 21766 51750
rect 21830 51686 21972 51750
rect 21624 51680 21972 51686
rect 22032 51886 22244 51892
rect 22032 51822 22174 51886
rect 22238 51822 22244 51886
rect 22032 51680 22244 51822
rect 22440 51886 22652 51892
rect 22440 51822 22582 51886
rect 22646 51822 22652 51886
rect 22440 51680 22652 51822
rect 27336 51816 27684 52094
rect 27608 51756 27684 51816
rect 20808 51620 20884 51680
rect 22032 51620 22108 51680
rect 22576 51620 22652 51680
rect 20808 51478 21020 51620
rect 20808 51414 20814 51478
rect 20878 51414 21020 51478
rect 20808 51408 21020 51414
rect 21216 51272 21428 51484
rect 21624 51478 21972 51484
rect 21624 51414 21766 51478
rect 21830 51414 21972 51478
rect 21624 51348 21972 51414
rect 21488 51272 21972 51348
rect 22032 51272 22244 51620
rect 22440 51272 22652 51620
rect 27336 51342 27684 51756
rect 27336 51278 27342 51342
rect 27406 51278 27684 51342
rect 21216 51212 21292 51272
rect 21488 51212 21564 51272
rect 20808 51206 21020 51212
rect 20808 51142 20814 51206
rect 20878 51142 21020 51206
rect 20808 51070 21020 51142
rect 20808 51006 20814 51070
rect 20878 51006 21020 51070
rect 20808 51000 21020 51006
rect 21216 51136 21564 51212
rect 21624 51212 21700 51272
rect 22032 51212 22108 51272
rect 22440 51212 22516 51272
rect 21216 51070 21428 51136
rect 21216 51006 21358 51070
rect 21422 51006 21428 51070
rect 21216 51000 21428 51006
rect 21624 51070 21972 51212
rect 21624 51006 21902 51070
rect 21966 51006 21972 51070
rect 21624 51000 21972 51006
rect 22032 51070 22244 51212
rect 22032 51006 22174 51070
rect 22238 51006 22244 51070
rect 22032 51000 22244 51006
rect 22440 51070 22652 51212
rect 27336 51136 27684 51278
rect 27608 51076 27684 51136
rect 22440 51006 22582 51070
rect 22646 51006 22652 51070
rect 22440 51000 22652 51006
rect 27336 51070 27684 51076
rect 27336 51006 27342 51070
rect 27406 51006 27684 51070
rect 1224 50934 1980 50940
rect 1224 50870 1230 50934
rect 1294 50870 1980 50934
rect 1224 50864 1980 50870
rect 1768 50808 1980 50864
rect 1768 50752 1794 50808
rect 1850 50752 1980 50808
rect 1768 50728 1980 50752
rect 20808 50798 21020 50804
rect 20808 50734 20814 50798
rect 20878 50734 21020 50798
rect 20808 50662 21020 50734
rect 20808 50598 20814 50662
rect 20878 50598 21020 50662
rect 20808 50592 21020 50598
rect 21216 50798 21428 50804
rect 21216 50734 21358 50798
rect 21422 50734 21428 50798
rect 21216 50592 21428 50734
rect 21624 50798 21972 50804
rect 21624 50734 21902 50798
rect 21966 50734 21972 50798
rect 21624 50662 21972 50734
rect 21624 50598 21902 50662
rect 21966 50598 21972 50662
rect 21624 50592 21972 50598
rect 22032 50798 22244 50804
rect 22032 50734 22174 50798
rect 22238 50734 22244 50798
rect 22032 50662 22244 50734
rect 22032 50598 22038 50662
rect 22102 50598 22244 50662
rect 22032 50592 22244 50598
rect 22440 50798 22652 50804
rect 22440 50734 22582 50798
rect 22646 50734 22652 50798
rect 22440 50662 22652 50734
rect 22440 50598 22446 50662
rect 22510 50598 22652 50662
rect 22440 50592 22652 50598
rect 27336 50592 27684 51006
rect 109344 51816 109556 52300
rect 114240 52294 114452 52300
rect 114240 52230 114382 52294
rect 114446 52230 114452 52294
rect 114240 52158 114452 52230
rect 114240 52094 114246 52158
rect 114310 52094 114452 52158
rect 114240 52088 114452 52094
rect 114648 52294 114860 52300
rect 114648 52230 114790 52294
rect 114854 52230 114860 52294
rect 114648 52158 114860 52230
rect 114648 52094 114654 52158
rect 114718 52094 114860 52158
rect 114648 52088 114860 52094
rect 115056 52294 115268 52300
rect 115056 52230 115198 52294
rect 115262 52230 115268 52294
rect 115056 52088 115268 52230
rect 115464 52088 115676 52300
rect 115872 52294 116084 52436
rect 134776 52432 134844 52488
rect 134900 52436 134988 52488
rect 134900 52432 135396 52436
rect 134776 52430 135396 52432
rect 134776 52366 135326 52430
rect 135390 52366 135396 52430
rect 134776 52360 135396 52366
rect 115872 52230 116014 52294
rect 116078 52230 116084 52294
rect 115872 52224 116084 52230
rect 115056 52028 115132 52088
rect 114240 51886 114452 51892
rect 114240 51822 114246 51886
rect 114310 51822 114452 51886
rect 109344 51756 109420 51816
rect 109344 51136 109556 51756
rect 114240 51680 114452 51822
rect 114648 51886 114860 51892
rect 114648 51822 114654 51886
rect 114718 51822 114860 51886
rect 114648 51680 114860 51822
rect 115056 51750 115268 52028
rect 115056 51686 115198 51750
rect 115262 51686 115268 51750
rect 115056 51680 115268 51686
rect 115464 51680 115676 52028
rect 115872 52022 116084 52028
rect 115872 51958 116014 52022
rect 116078 51958 116084 52022
rect 115872 51680 116084 51958
rect 114376 51620 114452 51680
rect 114784 51620 114860 51680
rect 115464 51620 115540 51680
rect 114240 51272 114452 51620
rect 114648 51272 114860 51620
rect 115192 51544 115540 51620
rect 115872 51620 115948 51680
rect 115192 51484 115268 51544
rect 115056 51478 115676 51484
rect 115056 51414 115198 51478
rect 115262 51414 115676 51478
rect 115056 51408 115676 51414
rect 115872 51478 116084 51620
rect 115872 51414 115878 51478
rect 115942 51414 116084 51478
rect 115872 51408 116084 51414
rect 115056 51272 115268 51408
rect 114240 51212 114316 51272
rect 114784 51212 114860 51272
rect 115192 51212 115268 51272
rect 109344 51076 109420 51136
rect 109344 50592 109556 51076
rect 114240 51070 114452 51212
rect 114240 51006 114246 51070
rect 114310 51006 114452 51070
rect 114240 51000 114452 51006
rect 114648 51070 114860 51212
rect 114648 51006 114654 51070
rect 114718 51006 114860 51070
rect 114648 51000 114860 51006
rect 115056 51070 115268 51212
rect 115056 51006 115062 51070
rect 115126 51006 115268 51070
rect 115056 51000 115268 51006
rect 115464 51272 115676 51408
rect 115464 51212 115540 51272
rect 115464 51070 115676 51212
rect 115464 51006 115470 51070
rect 115534 51006 115676 51070
rect 115464 51000 115676 51006
rect 115872 51206 116084 51212
rect 115872 51142 115878 51206
rect 115942 51142 116084 51206
rect 115872 51070 116084 51142
rect 115872 51006 116014 51070
rect 116078 51006 116084 51070
rect 115872 51000 116084 51006
rect 134776 50808 134988 50940
rect 114240 50798 114452 50804
rect 114240 50734 114246 50798
rect 114310 50734 114452 50798
rect 114240 50662 114452 50734
rect 114240 50598 114382 50662
rect 114446 50598 114452 50662
rect 114240 50592 114452 50598
rect 114648 50798 114860 50804
rect 114648 50734 114654 50798
rect 114718 50734 114860 50798
rect 114648 50662 114860 50734
rect 114648 50598 114790 50662
rect 114854 50598 114860 50662
rect 114648 50592 114860 50598
rect 115056 50798 115268 50804
rect 115056 50734 115062 50798
rect 115126 50734 115268 50798
rect 115056 50592 115268 50734
rect 115464 50798 115676 50804
rect 115464 50734 115470 50798
rect 115534 50734 115676 50798
rect 115464 50592 115676 50734
rect 115872 50798 116084 50804
rect 115872 50734 116014 50798
rect 116078 50734 116084 50798
rect 115872 50662 116084 50734
rect 134776 50752 134844 50808
rect 134900 50804 134988 50808
rect 134900 50798 135396 50804
rect 134900 50752 135326 50798
rect 134776 50734 135326 50752
rect 135390 50734 135396 50798
rect 134776 50728 135396 50734
rect 115872 50598 115878 50662
rect 115942 50598 116084 50662
rect 115872 50592 116084 50598
rect 27472 50532 27548 50592
rect 109344 50532 109420 50592
rect 115464 50532 115540 50592
rect 20808 50390 21020 50396
rect 20808 50326 20814 50390
rect 20878 50326 21020 50390
rect 20808 50254 21020 50326
rect 20808 50190 20950 50254
rect 21014 50190 21020 50254
rect 20808 50184 21020 50190
rect 21216 50254 21428 50396
rect 21624 50390 21972 50396
rect 21624 50326 21902 50390
rect 21966 50326 21972 50390
rect 21624 50260 21972 50326
rect 21526 50254 21972 50260
rect 21216 50190 21222 50254
rect 21286 50190 21428 50254
rect 21488 50190 21494 50254
rect 21558 50190 21972 50254
rect 21216 50184 21428 50190
rect 21526 50184 21972 50190
rect 22032 50390 22244 50396
rect 22032 50326 22038 50390
rect 22102 50326 22244 50390
rect 22032 50254 22244 50326
rect 22032 50190 22174 50254
rect 22238 50190 22244 50254
rect 22032 50184 22244 50190
rect 22440 50390 22652 50396
rect 22440 50326 22446 50390
rect 22510 50326 22652 50390
rect 22440 50254 22652 50326
rect 22440 50190 22582 50254
rect 22646 50190 22652 50254
rect 22440 50184 22652 50190
rect 27336 50320 27684 50532
rect 109344 50320 109556 50532
rect 115192 50456 115540 50532
rect 115192 50396 115268 50456
rect 114240 50390 114452 50396
rect 114240 50326 114382 50390
rect 114446 50326 114452 50390
rect 27336 50260 27412 50320
rect 109344 50260 109420 50320
rect 27336 50048 27684 50260
rect 109344 50048 109556 50260
rect 114240 50254 114452 50326
rect 114240 50190 114246 50254
rect 114310 50190 114452 50254
rect 114240 50184 114452 50190
rect 114648 50390 114860 50396
rect 114648 50326 114790 50390
rect 114854 50326 114860 50390
rect 114648 50254 114860 50326
rect 114648 50190 114790 50254
rect 114854 50190 114860 50254
rect 114648 50184 114860 50190
rect 115056 50320 115676 50396
rect 115056 50184 115268 50320
rect 115464 50254 115676 50320
rect 115464 50190 115606 50254
rect 115670 50190 115676 50254
rect 115464 50184 115676 50190
rect 115872 50390 116084 50396
rect 115872 50326 115878 50390
rect 115942 50326 116084 50390
rect 115872 50254 116084 50326
rect 115872 50190 115878 50254
rect 115942 50190 116084 50254
rect 115872 50184 116084 50190
rect 27608 49988 27684 50048
rect 109480 49988 109556 50048
rect 20808 49982 21020 49988
rect 20808 49918 20950 49982
rect 21014 49918 21020 49982
rect 20808 49846 21020 49918
rect 20808 49782 20814 49846
rect 20878 49782 21020 49846
rect 20808 49776 21020 49782
rect 21216 49982 21564 49988
rect 21216 49918 21222 49982
rect 21286 49918 21494 49982
rect 21558 49918 21564 49982
rect 21216 49912 21564 49918
rect 21216 49852 21428 49912
rect 21624 49852 21972 49988
rect 21216 49846 21972 49852
rect 21216 49782 21766 49846
rect 21830 49782 21972 49846
rect 21216 49776 21972 49782
rect 22032 49982 22244 49988
rect 22032 49918 22174 49982
rect 22238 49918 22244 49982
rect 22032 49846 22244 49918
rect 22032 49782 22174 49846
rect 22238 49782 22244 49846
rect 22032 49776 22244 49782
rect 22440 49982 22652 49988
rect 22440 49918 22582 49982
rect 22646 49918 22652 49982
rect 22440 49846 22652 49918
rect 22440 49782 22446 49846
rect 22510 49782 22652 49846
rect 22440 49776 22652 49782
rect 27336 49776 27684 49988
rect 109344 49776 109556 49988
rect 114240 49982 114452 49988
rect 114240 49918 114246 49982
rect 114310 49918 114452 49982
rect 114240 49846 114452 49918
rect 114240 49782 114246 49846
rect 114310 49782 114452 49846
rect 114240 49776 114452 49782
rect 114648 49982 114860 49988
rect 114648 49918 114790 49982
rect 114854 49918 114860 49982
rect 114648 49846 114860 49918
rect 114648 49782 114654 49846
rect 114718 49782 114860 49846
rect 114648 49776 114860 49782
rect 115056 49846 115268 49988
rect 115464 49982 115676 49988
rect 115464 49918 115606 49982
rect 115670 49918 115676 49982
rect 115464 49852 115676 49918
rect 115366 49846 115676 49852
rect 115056 49782 115198 49846
rect 115262 49782 115268 49846
rect 115328 49782 115334 49846
rect 115398 49782 115676 49846
rect 115056 49776 115268 49782
rect 115366 49776 115676 49782
rect 115872 49982 116084 49988
rect 115872 49918 115878 49982
rect 115942 49918 116084 49982
rect 115872 49846 116084 49918
rect 115872 49782 115878 49846
rect 115942 49782 116084 49846
rect 115872 49776 116084 49782
rect 27472 49716 27548 49776
rect 109480 49716 109556 49776
rect 20808 49574 21020 49580
rect 20808 49510 20814 49574
rect 20878 49510 21020 49574
rect 20808 49438 21020 49510
rect 20808 49374 20950 49438
rect 21014 49374 21020 49438
rect 20808 49368 21020 49374
rect 21216 49438 21428 49580
rect 21216 49374 21222 49438
rect 21286 49374 21428 49438
rect 21216 49368 21428 49374
rect 21624 49574 21972 49580
rect 21624 49510 21766 49574
rect 21830 49510 21972 49574
rect 21624 49438 21972 49510
rect 21624 49374 21630 49438
rect 21694 49374 21972 49438
rect 21624 49368 21972 49374
rect 22032 49574 22244 49580
rect 22032 49510 22174 49574
rect 22238 49510 22244 49574
rect 22032 49438 22244 49510
rect 22032 49374 22038 49438
rect 22102 49374 22244 49438
rect 22032 49368 22244 49374
rect 22440 49574 22652 49580
rect 22440 49510 22446 49574
rect 22510 49510 22652 49574
rect 22440 49438 22652 49510
rect 22440 49374 22446 49438
rect 22510 49374 22652 49438
rect 22440 49368 22652 49374
rect 27336 49504 27684 49716
rect 109344 49504 109556 49716
rect 114240 49574 114452 49580
rect 114240 49510 114246 49574
rect 114310 49510 114452 49574
rect 27336 49444 27412 49504
rect 109344 49444 109420 49504
rect 27336 49232 27684 49444
rect 109344 49232 109556 49444
rect 114240 49438 114452 49510
rect 114240 49374 114382 49438
rect 114446 49374 114452 49438
rect 114240 49368 114452 49374
rect 114648 49574 114860 49580
rect 114648 49510 114654 49574
rect 114718 49510 114860 49574
rect 114648 49438 114860 49510
rect 114648 49374 114654 49438
rect 114718 49374 114860 49438
rect 114648 49368 114860 49374
rect 115056 49574 115404 49580
rect 115056 49510 115198 49574
rect 115262 49510 115334 49574
rect 115398 49510 115404 49574
rect 115056 49504 115404 49510
rect 115056 49444 115268 49504
rect 115464 49444 115676 49580
rect 115056 49368 115676 49444
rect 115872 49574 116084 49580
rect 115872 49510 115878 49574
rect 115942 49510 116084 49574
rect 115872 49438 116084 49510
rect 115872 49374 115878 49438
rect 115942 49374 116084 49438
rect 115872 49368 116084 49374
rect 115464 49308 115540 49368
rect 115192 49232 115540 49308
rect 27472 49172 27548 49232
rect 109344 49172 109420 49232
rect 115192 49172 115268 49232
rect 1768 49128 1980 49172
rect 1768 49072 1794 49128
rect 1850 49072 1980 49128
rect 1768 49036 1980 49072
rect 1224 49030 1980 49036
rect 1224 48966 1230 49030
rect 1294 48966 1980 49030
rect 1224 48960 1980 48966
rect 20808 49166 21020 49172
rect 20808 49102 20950 49166
rect 21014 49102 21020 49166
rect 20808 49030 21020 49102
rect 20808 48966 20814 49030
rect 20878 48966 21020 49030
rect 20808 48960 21020 48966
rect 21216 49166 21428 49172
rect 21216 49102 21222 49166
rect 21286 49102 21428 49166
rect 21216 49030 21428 49102
rect 21624 49166 21972 49172
rect 21624 49102 21630 49166
rect 21694 49102 21972 49166
rect 21624 49036 21972 49102
rect 21526 49030 21972 49036
rect 21216 48966 21358 49030
rect 21422 48966 21428 49030
rect 21488 48966 21494 49030
rect 21558 48966 21972 49030
rect 21216 48960 21428 48966
rect 21526 48960 21972 48966
rect 22032 49166 22244 49172
rect 22032 49102 22038 49166
rect 22102 49102 22244 49166
rect 22032 49030 22244 49102
rect 22032 48966 22174 49030
rect 22238 48966 22244 49030
rect 22032 48960 22244 48966
rect 22440 49166 22652 49172
rect 22440 49102 22446 49166
rect 22510 49102 22652 49166
rect 22440 49030 22652 49102
rect 22440 48966 22582 49030
rect 22646 48966 22652 49030
rect 22440 48960 22652 48966
rect 27336 48960 27684 49172
rect 109344 48960 109556 49172
rect 114240 49166 114452 49172
rect 114240 49102 114382 49166
rect 114446 49102 114452 49166
rect 114240 49030 114452 49102
rect 114240 48966 114246 49030
rect 114310 48966 114452 49030
rect 114240 48960 114452 48966
rect 114648 49166 114860 49172
rect 114648 49102 114654 49166
rect 114718 49102 114860 49166
rect 114648 49030 114860 49102
rect 114648 48966 114654 49030
rect 114718 48966 114860 49030
rect 114648 48960 114860 48966
rect 115056 49096 115676 49172
rect 115056 48960 115268 49096
rect 115464 49030 115676 49096
rect 115464 48966 115606 49030
rect 115670 48966 115676 49030
rect 115464 48960 115676 48966
rect 115872 49166 116084 49172
rect 115872 49102 115878 49166
rect 115942 49102 116084 49166
rect 115872 49030 116084 49102
rect 115872 48966 116014 49030
rect 116078 48966 116084 49030
rect 115872 48960 116084 48966
rect 134776 49128 134988 49172
rect 134776 49072 134844 49128
rect 134900 49072 134988 49128
rect 134776 49036 134988 49072
rect 134776 49030 135396 49036
rect 134776 48966 135326 49030
rect 135390 48966 135396 49030
rect 134776 48960 135396 48966
rect 27336 48900 27412 48960
rect 109480 48900 109556 48960
rect 20808 48758 21020 48764
rect 20808 48694 20814 48758
rect 20878 48694 21020 48758
rect 20808 48552 21020 48694
rect 21216 48758 21564 48764
rect 21216 48694 21358 48758
rect 21422 48694 21494 48758
rect 21558 48694 21564 48758
rect 21216 48688 21564 48694
rect 21216 48628 21428 48688
rect 21624 48628 21972 48764
rect 21216 48622 21972 48628
rect 21216 48558 21766 48622
rect 21830 48558 21972 48622
rect 21216 48552 21972 48558
rect 22032 48758 22244 48764
rect 22032 48694 22174 48758
rect 22238 48694 22244 48758
rect 22032 48622 22244 48694
rect 22032 48558 22174 48622
rect 22238 48558 22244 48622
rect 22032 48552 22244 48558
rect 22440 48758 22652 48764
rect 22440 48694 22582 48758
rect 22646 48694 22652 48758
rect 22440 48622 22652 48694
rect 27336 48688 27684 48900
rect 109344 48688 109556 48900
rect 27472 48628 27548 48688
rect 109480 48628 109556 48688
rect 22440 48558 22446 48622
rect 22510 48558 22652 48622
rect 22440 48552 22652 48558
rect 20808 48492 20884 48552
rect 20808 48350 21020 48492
rect 27336 48416 27684 48628
rect 109344 48416 109556 48628
rect 114240 48758 114452 48764
rect 114240 48694 114246 48758
rect 114310 48694 114452 48758
rect 114240 48622 114452 48694
rect 114240 48558 114382 48622
rect 114446 48558 114452 48622
rect 114240 48552 114452 48558
rect 114648 48758 114860 48764
rect 114648 48694 114654 48758
rect 114718 48694 114860 48758
rect 114648 48622 114860 48694
rect 114648 48558 114654 48622
rect 114718 48558 114860 48622
rect 114648 48552 114860 48558
rect 115056 48622 115268 48764
rect 115056 48558 115062 48622
rect 115126 48558 115268 48622
rect 115056 48552 115268 48558
rect 115464 48758 115676 48764
rect 115464 48694 115606 48758
rect 115670 48694 115676 48758
rect 115464 48622 115676 48694
rect 115464 48558 115470 48622
rect 115534 48558 115676 48622
rect 115464 48552 115676 48558
rect 115872 48758 116084 48764
rect 115872 48694 116014 48758
rect 116078 48694 116084 48758
rect 115872 48552 116084 48694
rect 115872 48492 115948 48552
rect 27336 48356 27412 48416
rect 109344 48356 109420 48416
rect 20808 48286 20814 48350
rect 20878 48286 21020 48350
rect 20808 48280 21020 48286
rect 21216 48144 21428 48356
rect 21624 48350 21972 48356
rect 21624 48286 21766 48350
rect 21830 48286 21972 48350
rect 21624 48144 21972 48286
rect 22032 48350 22244 48356
rect 22032 48286 22174 48350
rect 22238 48286 22244 48350
rect 22032 48214 22244 48286
rect 22032 48150 22174 48214
rect 22238 48150 22244 48214
rect 22032 48144 22244 48150
rect 22440 48350 22652 48356
rect 22440 48286 22446 48350
rect 22510 48286 22652 48350
rect 22440 48214 22652 48286
rect 22440 48150 22446 48214
rect 22510 48150 22652 48214
rect 22440 48144 22652 48150
rect 21216 48084 21292 48144
rect 21896 48084 21972 48144
rect 20808 48078 21020 48084
rect 20808 48014 20814 48078
rect 20878 48014 21020 48078
rect 20808 47736 21020 48014
rect 21216 47948 21428 48084
rect 21624 47948 21972 48084
rect 21216 47872 21972 47948
rect 21216 47812 21428 47872
rect 21216 47806 21564 47812
rect 21216 47742 21494 47806
rect 21558 47742 21564 47806
rect 21216 47736 21564 47742
rect 21624 47736 21972 47872
rect 22032 47942 22244 47948
rect 22032 47878 22174 47942
rect 22238 47878 22244 47942
rect 22032 47736 22244 47878
rect 20944 47676 21020 47736
rect 22168 47676 22244 47736
rect 1224 47534 1980 47540
rect 1224 47470 1230 47534
rect 1294 47470 1980 47534
rect 1224 47464 1980 47470
rect 20808 47534 21020 47676
rect 20808 47470 20814 47534
rect 20878 47470 21020 47534
rect 20808 47464 21020 47470
rect 1768 47448 1980 47464
rect 1768 47392 1794 47448
rect 1850 47392 1980 47448
rect 1768 47328 1980 47392
rect 21216 47328 21428 47540
rect 21526 47534 21972 47540
rect 21488 47470 21494 47534
rect 21558 47470 21972 47534
rect 21526 47464 21972 47470
rect 21624 47328 21972 47464
rect 22032 47328 22244 47676
rect 22440 47942 22652 47948
rect 22440 47878 22446 47942
rect 22510 47878 22652 47942
rect 22440 47736 22652 47878
rect 27336 47872 27684 48356
rect 109344 47872 109556 48356
rect 114240 48350 114452 48356
rect 114240 48286 114382 48350
rect 114446 48286 114452 48350
rect 114240 48214 114452 48286
rect 114240 48150 114246 48214
rect 114310 48150 114452 48214
rect 114240 48144 114452 48150
rect 114648 48350 114860 48356
rect 114648 48286 114654 48350
rect 114718 48286 114860 48350
rect 114648 48214 114860 48286
rect 114648 48150 114790 48214
rect 114854 48150 114860 48214
rect 114648 48144 114860 48150
rect 115056 48350 115404 48356
rect 115056 48286 115062 48350
rect 115126 48286 115334 48350
rect 115398 48286 115404 48350
rect 115056 48280 115404 48286
rect 115464 48350 115676 48356
rect 115464 48286 115470 48350
rect 115534 48286 115676 48350
rect 115056 48220 115268 48280
rect 115464 48220 115676 48286
rect 115872 48350 116084 48492
rect 115872 48286 115878 48350
rect 115942 48286 116084 48350
rect 115872 48280 116084 48286
rect 115056 48144 115676 48220
rect 115192 48084 115268 48144
rect 114240 47942 114452 47948
rect 114240 47878 114246 47942
rect 114310 47878 114452 47942
rect 27472 47812 27548 47872
rect 109344 47812 109420 47872
rect 22440 47676 22516 47736
rect 22440 47328 22652 47676
rect 21216 47268 21292 47328
rect 21624 47268 21700 47328
rect 22032 47268 22108 47328
rect 22576 47268 22652 47328
rect 20808 47262 21020 47268
rect 20808 47198 20814 47262
rect 20878 47198 21020 47262
rect 20808 47126 21020 47198
rect 20808 47062 20950 47126
rect 21014 47062 21020 47126
rect 20808 47056 21020 47062
rect 21216 47126 21428 47268
rect 21216 47062 21358 47126
rect 21422 47062 21428 47126
rect 21216 47056 21428 47062
rect 21624 47126 21972 47268
rect 21624 47062 21766 47126
rect 21830 47062 21972 47126
rect 21624 47056 21972 47062
rect 22032 46920 22244 47268
rect 22168 46860 22244 46920
rect 20808 46854 21020 46860
rect 20808 46790 20950 46854
rect 21014 46790 21020 46854
rect 20808 46718 21020 46790
rect 20808 46654 20814 46718
rect 20878 46654 21020 46718
rect 20808 46648 21020 46654
rect 21216 46854 21428 46860
rect 21216 46790 21358 46854
rect 21422 46790 21428 46854
rect 21216 46724 21428 46790
rect 21624 46854 21972 46860
rect 21624 46790 21766 46854
rect 21830 46790 21972 46854
rect 21624 46724 21972 46790
rect 21216 46648 21972 46724
rect 22032 46718 22244 46860
rect 22032 46654 22174 46718
rect 22238 46654 22244 46718
rect 22032 46648 22244 46654
rect 22440 46920 22652 47268
rect 27336 47262 27684 47812
rect 27336 47198 27342 47262
rect 27406 47198 27684 47262
rect 27336 47192 27684 47198
rect 109344 47262 109556 47812
rect 114240 47736 114452 47878
rect 114648 47942 114860 47948
rect 114648 47878 114790 47942
rect 114854 47878 114860 47942
rect 114648 47736 114860 47878
rect 115056 47806 115268 48084
rect 115366 48078 115676 48084
rect 115328 48014 115334 48078
rect 115398 48014 115676 48078
rect 115366 48008 115676 48014
rect 115056 47742 115062 47806
rect 115126 47742 115268 47806
rect 115056 47736 115268 47742
rect 115464 47736 115676 48008
rect 115872 48078 116084 48084
rect 115872 48014 115878 48078
rect 115942 48014 116084 48078
rect 115872 47736 116084 48014
rect 114240 47676 114316 47736
rect 114648 47676 114724 47736
rect 116008 47676 116084 47736
rect 114240 47328 114452 47676
rect 114648 47328 114860 47676
rect 115056 47534 115268 47540
rect 115056 47470 115062 47534
rect 115126 47470 115268 47534
rect 115056 47328 115268 47470
rect 114376 47268 114452 47328
rect 114784 47268 114860 47328
rect 115192 47268 115268 47328
rect 115464 47328 115676 47540
rect 115872 47534 116084 47676
rect 115872 47470 115878 47534
rect 115942 47470 116084 47534
rect 115872 47464 116084 47470
rect 134776 47534 135396 47540
rect 134776 47470 135326 47534
rect 135390 47470 135396 47534
rect 134776 47464 135396 47470
rect 134776 47448 134988 47464
rect 134776 47392 134844 47448
rect 134900 47392 134988 47448
rect 134776 47328 134988 47392
rect 115464 47268 115540 47328
rect 109344 47198 109350 47262
rect 109414 47198 109556 47262
rect 109344 47192 109556 47198
rect 27336 46990 27684 46996
rect 27336 46926 27342 46990
rect 27406 46926 27684 46990
rect 22440 46860 22516 46920
rect 22440 46718 22652 46860
rect 22440 46654 22582 46718
rect 22646 46654 22652 46718
rect 22440 46648 22652 46654
rect 27336 46854 27684 46926
rect 27336 46790 27342 46854
rect 27406 46790 27684 46854
rect 27336 46648 27684 46790
rect 109344 46990 109556 46996
rect 109344 46926 109350 46990
rect 109414 46926 109556 46990
rect 109344 46854 109556 46926
rect 109344 46790 109486 46854
rect 109550 46790 109556 46854
rect 109344 46648 109556 46790
rect 114240 46920 114452 47268
rect 114648 46920 114860 47268
rect 115056 47192 115676 47268
rect 115056 47132 115268 47192
rect 115056 47126 115404 47132
rect 115056 47062 115334 47126
rect 115398 47062 115404 47126
rect 115056 47056 115404 47062
rect 115464 47056 115676 47192
rect 115872 47262 116084 47268
rect 115872 47198 115878 47262
rect 115942 47198 116084 47262
rect 115872 47126 116084 47198
rect 115872 47062 115878 47126
rect 115942 47062 116084 47126
rect 115872 47056 116084 47062
rect 114240 46860 114316 46920
rect 114648 46860 114724 46920
rect 114240 46718 114452 46860
rect 114240 46654 114246 46718
rect 114310 46654 114452 46718
rect 114240 46648 114452 46654
rect 114648 46718 114860 46860
rect 114648 46654 114654 46718
rect 114718 46654 114860 46718
rect 114648 46648 114860 46654
rect 21216 46512 21428 46648
rect 21624 46512 21972 46648
rect 21352 46452 21428 46512
rect 21896 46452 21972 46512
rect 27336 46588 27412 46648
rect 109480 46588 109556 46648
rect 27336 46582 27684 46588
rect 27336 46518 27342 46582
rect 27406 46518 27684 46582
rect 20808 46446 21020 46452
rect 20808 46382 20814 46446
rect 20878 46382 21020 46446
rect 20808 46310 21020 46382
rect 20808 46246 20950 46310
rect 21014 46246 21020 46310
rect 20808 46240 21020 46246
rect 21216 46310 21428 46452
rect 21216 46246 21222 46310
rect 21286 46246 21428 46310
rect 21216 46240 21428 46246
rect 21624 46240 21972 46452
rect 22032 46446 22244 46452
rect 22032 46382 22174 46446
rect 22238 46382 22244 46446
rect 22032 46310 22244 46382
rect 22032 46246 22038 46310
rect 22102 46246 22244 46310
rect 22032 46240 22244 46246
rect 22440 46446 22652 46452
rect 22440 46382 22582 46446
rect 22646 46382 22652 46446
rect 22440 46310 22652 46382
rect 27336 46376 27684 46518
rect 109344 46582 109556 46588
rect 109344 46518 109486 46582
rect 109550 46518 109556 46582
rect 109344 46376 109556 46518
rect 115056 46512 115268 46860
rect 115366 46854 115676 46860
rect 115328 46790 115334 46854
rect 115398 46790 115676 46854
rect 115366 46784 115676 46790
rect 115464 46512 115676 46784
rect 115872 46854 116084 46860
rect 115872 46790 115878 46854
rect 115942 46790 116084 46854
rect 115872 46718 116084 46790
rect 115872 46654 116014 46718
rect 116078 46654 116084 46718
rect 115872 46648 116084 46654
rect 115056 46452 115132 46512
rect 115600 46452 115676 46512
rect 27608 46316 27684 46376
rect 109480 46316 109556 46376
rect 22440 46246 22582 46310
rect 22646 46246 22652 46310
rect 22440 46240 22652 46246
rect 27336 46240 27684 46316
rect 109344 46240 109556 46316
rect 114240 46446 114452 46452
rect 114240 46382 114246 46446
rect 114310 46382 114452 46446
rect 114240 46310 114452 46382
rect 114240 46246 114382 46310
rect 114446 46246 114452 46310
rect 114240 46240 114452 46246
rect 114648 46446 114860 46452
rect 114648 46382 114654 46446
rect 114718 46382 114860 46446
rect 114648 46310 114860 46382
rect 114648 46246 114790 46310
rect 114854 46246 114860 46310
rect 114648 46240 114860 46246
rect 115056 46310 115268 46452
rect 115464 46316 115676 46452
rect 115366 46310 115676 46316
rect 115056 46246 115198 46310
rect 115262 46246 115268 46310
rect 115328 46246 115334 46310
rect 115398 46246 115470 46310
rect 115534 46246 115676 46310
rect 115056 46240 115268 46246
rect 115366 46240 115676 46246
rect 115872 46446 116084 46452
rect 115872 46382 116014 46446
rect 116078 46382 116084 46446
rect 115872 46310 116084 46382
rect 115872 46246 115878 46310
rect 115942 46246 116084 46310
rect 115872 46240 116084 46246
rect 27462 46044 27560 46240
rect 109344 46044 109448 46240
rect 20808 46038 21020 46044
rect 20808 45974 20950 46038
rect 21014 45974 21020 46038
rect 1768 45768 1980 45908
rect 20808 45902 21020 45974
rect 20808 45838 20950 45902
rect 21014 45838 21020 45902
rect 20808 45832 21020 45838
rect 21216 46038 21428 46044
rect 21216 45974 21222 46038
rect 21286 45974 21428 46038
rect 21216 45902 21428 45974
rect 21216 45838 21358 45902
rect 21422 45838 21428 45902
rect 21216 45832 21428 45838
rect 21624 45832 21972 46044
rect 22032 46038 22244 46044
rect 22032 45974 22038 46038
rect 22102 45974 22244 46038
rect 22032 45902 22244 45974
rect 22032 45838 22038 45902
rect 22102 45838 22244 45902
rect 22032 45832 22244 45838
rect 22440 46038 22652 46044
rect 22440 45974 22582 46038
rect 22646 45974 22652 46038
rect 22440 45902 22652 45974
rect 22440 45838 22446 45902
rect 22510 45838 22652 45902
rect 22440 45832 22652 45838
rect 27336 45832 27684 46044
rect 109344 45832 109556 46044
rect 114240 46038 114452 46044
rect 114240 45974 114382 46038
rect 114446 45974 114452 46038
rect 114240 45902 114452 45974
rect 114240 45838 114382 45902
rect 114446 45838 114452 45902
rect 114240 45832 114452 45838
rect 114648 46038 114860 46044
rect 114648 45974 114790 46038
rect 114854 45974 114860 46038
rect 114648 45908 114860 45974
rect 115056 46038 115404 46044
rect 115056 45974 115198 46038
rect 115262 45974 115334 46038
rect 115398 45974 115404 46038
rect 115056 45968 115404 45974
rect 115464 46038 115676 46044
rect 115464 45974 115470 46038
rect 115534 45974 115676 46038
rect 114648 45902 114996 45908
rect 114648 45838 114654 45902
rect 114718 45838 114996 45902
rect 114648 45832 114996 45838
rect 115056 45832 115268 45968
rect 115464 45902 115676 45974
rect 115464 45838 115470 45902
rect 115534 45838 115676 45902
rect 115464 45832 115676 45838
rect 115872 46038 116084 46044
rect 115872 45974 115878 46038
rect 115942 45974 116084 46038
rect 115872 45902 116084 45974
rect 115872 45838 116014 45902
rect 116078 45838 116084 45902
rect 115872 45832 116084 45838
rect 21624 45772 21700 45832
rect 27608 45772 27684 45832
rect 109480 45772 109556 45832
rect 1768 45712 1794 45768
rect 1850 45712 1980 45768
rect 1768 45636 1980 45712
rect 21352 45696 21700 45772
rect 21352 45636 21428 45696
rect 1224 45630 1980 45636
rect 1224 45566 1230 45630
rect 1294 45566 1980 45630
rect 1224 45560 1980 45566
rect 20808 45630 21020 45636
rect 20808 45566 20950 45630
rect 21014 45566 21020 45630
rect 20808 45494 21020 45566
rect 20808 45430 20814 45494
rect 20878 45430 21020 45494
rect 20808 45424 21020 45430
rect 21216 45630 21972 45636
rect 21216 45566 21358 45630
rect 21422 45566 21972 45630
rect 21216 45560 21972 45566
rect 21216 45424 21428 45560
rect 21624 45494 21972 45560
rect 21624 45430 21766 45494
rect 21830 45430 21972 45494
rect 21624 45424 21972 45430
rect 22032 45630 22244 45636
rect 22032 45566 22038 45630
rect 22102 45566 22244 45630
rect 22032 45500 22244 45566
rect 22440 45630 22652 45636
rect 22440 45566 22446 45630
rect 22510 45566 22652 45630
rect 22032 45494 22380 45500
rect 22032 45430 22038 45494
rect 22102 45430 22380 45494
rect 22032 45424 22380 45430
rect 22440 45494 22652 45566
rect 27336 45560 27684 45772
rect 109344 45560 109556 45772
rect 114920 45772 114996 45832
rect 115872 45772 115948 45832
rect 114920 45696 115948 45772
rect 134776 45772 134988 45908
rect 134776 45768 135396 45772
rect 134776 45712 134844 45768
rect 134900 45766 135396 45768
rect 134900 45712 135326 45766
rect 134776 45702 135326 45712
rect 135390 45702 135396 45766
rect 134776 45696 135396 45702
rect 27472 45500 27548 45560
rect 109480 45500 109556 45560
rect 114240 45630 114452 45636
rect 114240 45566 114382 45630
rect 114446 45566 114452 45630
rect 114240 45500 114452 45566
rect 25878 45494 27684 45500
rect 22440 45430 22446 45494
rect 22510 45430 22652 45494
rect 25840 45430 25846 45494
rect 25910 45430 27684 45494
rect 22440 45424 22652 45430
rect 25878 45424 27684 45430
rect 22304 45364 22380 45424
rect 22304 45288 22924 45364
rect 22848 45228 22924 45288
rect 24208 45288 26052 45364
rect 27336 45288 27684 45424
rect 109344 45288 109556 45500
rect 113734 45494 114452 45500
rect 113696 45430 113702 45494
rect 113766 45430 114382 45494
rect 114446 45430 114452 45494
rect 113734 45424 114452 45430
rect 114648 45630 114860 45636
rect 114648 45566 114654 45630
rect 114718 45566 114860 45630
rect 114648 45494 114860 45566
rect 114648 45430 114790 45494
rect 114854 45430 114860 45494
rect 114648 45424 114860 45430
rect 115056 45494 115268 45636
rect 115464 45630 115676 45636
rect 115464 45566 115470 45630
rect 115534 45566 115676 45630
rect 115464 45500 115676 45566
rect 115366 45494 115676 45500
rect 115056 45430 115198 45494
rect 115262 45430 115268 45494
rect 115328 45430 115334 45494
rect 115398 45430 115676 45494
rect 115056 45424 115268 45430
rect 115366 45424 115676 45430
rect 115872 45630 116084 45636
rect 115872 45566 116014 45630
rect 116078 45566 116084 45630
rect 115872 45494 116084 45566
rect 134776 45560 134988 45696
rect 115872 45430 115878 45494
rect 115942 45430 116084 45494
rect 115872 45424 116084 45430
rect 114648 45364 114724 45424
rect 24208 45228 24284 45288
rect 25976 45228 26052 45288
rect 27472 45228 27548 45288
rect 109480 45228 109556 45288
rect 112200 45288 113500 45364
rect 112200 45228 112276 45288
rect 113424 45228 113500 45288
rect 114104 45288 114724 45364
rect 114104 45228 114180 45288
rect 20808 45222 21020 45228
rect 20808 45158 20814 45222
rect 20878 45158 21020 45222
rect 20808 45086 21020 45158
rect 20808 45022 20950 45086
rect 21014 45022 21020 45086
rect 20808 45016 21020 45022
rect 21216 45086 21428 45228
rect 21624 45222 21972 45228
rect 21624 45158 21766 45222
rect 21830 45158 21972 45222
rect 21624 45092 21972 45158
rect 21526 45086 21972 45092
rect 21216 45022 21222 45086
rect 21286 45022 21428 45086
rect 21488 45022 21494 45086
rect 21558 45022 21972 45086
rect 21216 45016 21428 45022
rect 21526 45016 21972 45022
rect 22032 45222 22244 45228
rect 22032 45158 22038 45222
rect 22102 45158 22244 45222
rect 22032 45086 22244 45158
rect 22032 45022 22038 45086
rect 22102 45022 22244 45086
rect 22032 45016 22244 45022
rect 22440 45222 22652 45228
rect 22440 45158 22446 45222
rect 22510 45158 22652 45222
rect 22440 45086 22652 45158
rect 22440 45022 22582 45086
rect 22646 45022 22652 45086
rect 22440 45016 22652 45022
rect 22848 45092 23060 45228
rect 23256 45152 24284 45228
rect 24344 45222 25916 45228
rect 24344 45158 25846 45222
rect 25910 45158 25916 45222
rect 24344 45152 25916 45158
rect 22848 45016 23196 45092
rect 23256 45086 23604 45152
rect 23256 45022 23262 45086
rect 23326 45022 23604 45086
rect 23256 45016 23604 45022
rect 24344 45016 24556 45152
rect 25976 45016 26188 45228
rect 27336 45016 27684 45228
rect 109344 45016 109556 45228
rect 110704 45152 112276 45228
rect 110704 45016 110916 45152
rect 112336 45092 112548 45228
rect 113424 45222 113772 45228
rect 113424 45158 113702 45222
rect 113766 45158 113772 45222
rect 113424 45152 113772 45158
rect 113832 45152 114180 45228
rect 114240 45222 114452 45228
rect 114240 45158 114382 45222
rect 114446 45158 114452 45222
rect 112336 45086 113364 45092
rect 112336 45022 112342 45086
rect 112406 45022 113364 45086
rect 112336 45016 113364 45022
rect 113424 45016 113636 45152
rect 113832 45016 114044 45152
rect 114240 45086 114452 45158
rect 114240 45022 114382 45086
rect 114446 45022 114452 45086
rect 114240 45016 114452 45022
rect 114648 45222 114860 45228
rect 114648 45158 114790 45222
rect 114854 45158 114860 45222
rect 114648 45086 114860 45158
rect 114648 45022 114654 45086
rect 114718 45022 114860 45086
rect 114648 45016 114860 45022
rect 115056 45222 115404 45228
rect 115056 45158 115198 45222
rect 115262 45158 115334 45222
rect 115398 45158 115404 45222
rect 115056 45152 115404 45158
rect 115056 45092 115268 45152
rect 115464 45092 115676 45228
rect 115056 45016 115676 45092
rect 115872 45222 116084 45228
rect 115872 45158 115878 45222
rect 115942 45158 116084 45222
rect 115872 45086 116084 45158
rect 115872 45022 115878 45086
rect 115942 45022 116084 45086
rect 115872 45016 116084 45022
rect 23120 44956 23196 45016
rect 24344 44956 24420 45016
rect 27472 44956 27548 45016
rect 109344 44956 109420 45016
rect 113288 44956 113364 45016
rect 113832 44956 113908 45016
rect 115464 44956 115540 45016
rect 23120 44880 24420 44956
rect 20808 44814 21020 44820
rect 20808 44750 20950 44814
rect 21014 44750 21020 44814
rect 20808 44608 21020 44750
rect 21216 44814 21564 44820
rect 21216 44750 21222 44814
rect 21286 44750 21494 44814
rect 21558 44750 21564 44814
rect 21216 44744 21564 44750
rect 21216 44684 21428 44744
rect 21624 44684 21972 44820
rect 21216 44678 21972 44684
rect 21216 44614 21358 44678
rect 21422 44614 21972 44678
rect 21216 44608 21972 44614
rect 22032 44814 22244 44820
rect 22032 44750 22038 44814
rect 22102 44750 22244 44814
rect 22032 44678 22244 44750
rect 22032 44614 22174 44678
rect 22238 44614 22244 44678
rect 22032 44608 22244 44614
rect 22440 44814 23332 44820
rect 22440 44750 22582 44814
rect 22646 44750 23262 44814
rect 23326 44750 23332 44814
rect 22440 44744 23332 44750
rect 27336 44744 27684 44956
rect 109344 44744 109556 44956
rect 113288 44880 113908 44956
rect 115192 44880 115540 44956
rect 115192 44820 115268 44880
rect 114240 44814 114452 44820
rect 114240 44750 114382 44814
rect 114446 44750 114452 44814
rect 22440 44678 22652 44744
rect 27472 44684 27548 44744
rect 109344 44684 109420 44744
rect 22440 44614 22446 44678
rect 22510 44614 22652 44678
rect 22440 44608 22652 44614
rect 20808 44548 20884 44608
rect 21352 44548 21428 44608
rect 20808 44200 21020 44548
rect 21352 44472 21700 44548
rect 27336 44472 27684 44684
rect 109344 44678 112412 44684
rect 109344 44614 112342 44678
rect 112406 44614 112412 44678
rect 109344 44608 112412 44614
rect 114240 44678 114452 44750
rect 114240 44614 114246 44678
rect 114310 44614 114452 44678
rect 114240 44608 114452 44614
rect 114648 44814 114860 44820
rect 114648 44750 114654 44814
rect 114718 44750 114860 44814
rect 114648 44678 114860 44750
rect 114648 44614 114654 44678
rect 114718 44614 114860 44678
rect 114648 44608 114860 44614
rect 115056 44744 115676 44820
rect 115056 44608 115268 44744
rect 115464 44678 115676 44744
rect 115464 44614 115470 44678
rect 115534 44614 115676 44678
rect 115464 44608 115676 44614
rect 115872 44814 116084 44820
rect 115872 44750 115878 44814
rect 115942 44750 116084 44814
rect 115872 44608 116084 44750
rect 109344 44472 109556 44608
rect 21624 44412 21700 44472
rect 27608 44412 27684 44472
rect 109480 44412 109556 44472
rect 115872 44548 115948 44608
rect 21216 44406 21428 44412
rect 21216 44342 21358 44406
rect 21422 44342 21428 44406
rect 21216 44200 21428 44342
rect 21624 44200 21972 44412
rect 22032 44406 22244 44412
rect 22032 44342 22174 44406
rect 22238 44342 22244 44406
rect 22032 44270 22244 44342
rect 22032 44206 22174 44270
rect 22238 44206 22244 44270
rect 22032 44200 22244 44206
rect 22440 44406 22652 44412
rect 22440 44342 22446 44406
rect 22510 44342 22652 44406
rect 22440 44270 22652 44342
rect 22440 44206 22582 44270
rect 22646 44206 22652 44270
rect 22440 44200 22652 44206
rect 20808 44140 20884 44200
rect 21352 44140 21428 44200
rect 21760 44140 21836 44200
rect 1224 44134 1980 44140
rect 1224 44070 1230 44134
rect 1294 44088 1980 44134
rect 1294 44070 1794 44088
rect 1224 44064 1794 44070
rect 1768 44032 1794 44064
rect 1850 44032 1980 44088
rect 1768 43928 1980 44032
rect 20808 43792 21020 44140
rect 21216 43792 21428 44140
rect 21624 43862 21972 44140
rect 21624 43798 21766 43862
rect 21830 43798 21972 43862
rect 21624 43792 21972 43798
rect 22032 43998 22244 44004
rect 22032 43934 22174 43998
rect 22238 43934 22244 43998
rect 22032 43862 22244 43934
rect 22032 43798 22038 43862
rect 22102 43798 22244 43862
rect 22032 43792 22244 43798
rect 22440 43998 22652 44004
rect 22440 43934 22582 43998
rect 22646 43934 22652 43998
rect 22440 43862 22652 43934
rect 27336 43928 27684 44412
rect 27608 43868 27684 43928
rect 22440 43798 22446 43862
rect 22510 43798 22652 43862
rect 22440 43792 22652 43798
rect 20808 43732 20884 43792
rect 20808 43590 21020 43732
rect 27336 43726 27684 43868
rect 27336 43662 27478 43726
rect 27542 43662 27684 43726
rect 27336 43656 27684 43662
rect 109344 43928 109556 44412
rect 114240 44406 114452 44412
rect 114240 44342 114246 44406
rect 114310 44342 114452 44406
rect 114240 44270 114452 44342
rect 114240 44206 114382 44270
rect 114446 44206 114452 44270
rect 114240 44200 114452 44206
rect 114648 44406 114860 44412
rect 114648 44342 114654 44406
rect 114718 44342 114860 44406
rect 114648 44270 114860 44342
rect 114648 44206 114790 44270
rect 114854 44206 114860 44270
rect 114648 44200 114860 44206
rect 115056 44406 115676 44412
rect 115056 44342 115470 44406
rect 115534 44342 115676 44406
rect 115056 44336 115676 44342
rect 115056 44276 115268 44336
rect 115056 44200 115404 44276
rect 115464 44200 115676 44336
rect 115872 44200 116084 44548
rect 115328 44140 115404 44200
rect 115872 44140 115948 44200
rect 114240 43998 114452 44004
rect 114240 43934 114382 43998
rect 114446 43934 114452 43998
rect 109344 43868 109420 43928
rect 109344 43726 109556 43868
rect 114240 43862 114452 43934
rect 114240 43798 114382 43862
rect 114446 43798 114452 43862
rect 114240 43792 114452 43798
rect 114648 43998 114860 44004
rect 114648 43934 114790 43998
rect 114854 43934 114860 43998
rect 114648 43862 114860 43934
rect 114648 43798 114790 43862
rect 114854 43798 114860 43862
rect 114648 43792 114860 43798
rect 115056 43868 115268 44140
rect 115328 44064 115676 44140
rect 115464 43868 115676 44064
rect 115056 43862 115676 43868
rect 115056 43798 115198 43862
rect 115262 43798 115676 43862
rect 115056 43792 115676 43798
rect 115872 43792 116084 44140
rect 134776 44088 134988 44140
rect 134776 44032 134844 44088
rect 134900 44032 134988 44088
rect 134776 44004 134988 44032
rect 134776 43998 135396 44004
rect 134776 43934 135326 43998
rect 135390 43934 135396 43998
rect 134776 43928 135396 43934
rect 109344 43662 109350 43726
rect 109414 43662 109556 43726
rect 109344 43656 109556 43662
rect 115192 43732 115268 43792
rect 115872 43732 115948 43792
rect 115192 43656 115540 43732
rect 27472 43596 27548 43656
rect 109344 43596 109420 43656
rect 115464 43596 115540 43656
rect 20808 43526 20814 43590
rect 20878 43526 21020 43590
rect 20808 43520 21020 43526
rect 21216 43460 21428 43596
rect 21624 43590 21972 43596
rect 21624 43526 21766 43590
rect 21830 43526 21972 43590
rect 21216 43384 21564 43460
rect 21624 43454 21972 43526
rect 21624 43390 21630 43454
rect 21694 43390 21972 43454
rect 21624 43384 21972 43390
rect 22032 43590 22244 43596
rect 22032 43526 22038 43590
rect 22102 43526 22244 43590
rect 22032 43384 22244 43526
rect 21488 43324 21564 43384
rect 21896 43324 21972 43384
rect 22168 43324 22244 43384
rect 20808 43318 21020 43324
rect 20808 43254 20814 43318
rect 20878 43254 21020 43318
rect 20808 43182 21020 43254
rect 20808 43118 20814 43182
rect 20878 43118 21020 43182
rect 20808 43112 21020 43118
rect 21216 43188 21428 43324
rect 21488 43248 21972 43324
rect 21216 43182 21564 43188
rect 21216 43118 21222 43182
rect 21286 43118 21494 43182
rect 21558 43118 21564 43182
rect 21216 43112 21564 43118
rect 21624 43112 21972 43248
rect 22032 42976 22244 43324
rect 22440 43590 22652 43596
rect 22440 43526 22446 43590
rect 22510 43526 22652 43590
rect 22440 43384 22652 43526
rect 27336 43454 27684 43596
rect 27336 43390 27478 43454
rect 27542 43390 27684 43454
rect 22440 43324 22516 43384
rect 22440 42976 22652 43324
rect 27336 43318 27684 43390
rect 27336 43254 27614 43318
rect 27678 43254 27684 43318
rect 27336 43248 27684 43254
rect 109344 43454 109556 43596
rect 109344 43390 109350 43454
rect 109414 43390 109556 43454
rect 109344 43318 109556 43390
rect 109344 43254 109350 43318
rect 109414 43254 109556 43318
rect 109344 43248 109556 43254
rect 114240 43590 114452 43596
rect 114240 43526 114382 43590
rect 114446 43526 114452 43590
rect 114240 43384 114452 43526
rect 114648 43590 114860 43596
rect 114648 43526 114790 43590
rect 114854 43526 114860 43590
rect 114648 43384 114860 43526
rect 115056 43590 115268 43596
rect 115056 43526 115198 43590
rect 115262 43526 115268 43590
rect 115056 43384 115268 43526
rect 115464 43384 115676 43596
rect 115872 43590 116084 43732
rect 115872 43526 116014 43590
rect 116078 43526 116084 43590
rect 115872 43520 116084 43526
rect 114240 43324 114316 43384
rect 114648 43324 114724 43384
rect 115056 43324 115132 43384
rect 115464 43324 115540 43384
rect 22168 42916 22244 42976
rect 22576 42916 22652 42976
rect 20808 42910 21020 42916
rect 20808 42846 20814 42910
rect 20878 42846 21020 42910
rect 20808 42774 21020 42846
rect 20808 42710 20814 42774
rect 20878 42710 21020 42774
rect 20808 42704 21020 42710
rect 21216 42910 21428 42916
rect 21216 42846 21222 42910
rect 21286 42846 21428 42910
rect 21216 42644 21428 42846
rect 21624 42644 21972 42916
rect 22032 42774 22244 42916
rect 22032 42710 22174 42774
rect 22238 42710 22244 42774
rect 22032 42704 22244 42710
rect 22440 42774 22652 42916
rect 22440 42710 22446 42774
rect 22510 42710 22652 42774
rect 22440 42704 22652 42710
rect 27336 43046 27684 43052
rect 27336 42982 27614 43046
rect 27678 42982 27684 43046
rect 27336 42704 27684 42982
rect 109344 43046 109556 43052
rect 109344 42982 109350 43046
rect 109414 42982 109556 43046
rect 109344 42910 109556 42982
rect 109344 42846 109350 42910
rect 109414 42846 109556 42910
rect 109344 42704 109556 42846
rect 114240 42976 114452 43324
rect 114648 42976 114860 43324
rect 115056 43182 115268 43324
rect 115056 43118 115062 43182
rect 115126 43118 115268 43182
rect 115056 43112 115268 43118
rect 115464 43112 115676 43324
rect 115872 43318 116084 43324
rect 115872 43254 116014 43318
rect 116078 43254 116084 43318
rect 115872 43182 116084 43254
rect 115872 43118 116014 43182
rect 116078 43118 116084 43182
rect 115872 43112 116084 43118
rect 114240 42916 114316 42976
rect 114784 42916 114860 42976
rect 114240 42774 114452 42916
rect 114240 42710 114246 42774
rect 114310 42710 114452 42774
rect 114240 42704 114452 42710
rect 114648 42774 114860 42916
rect 114648 42710 114790 42774
rect 114854 42710 114860 42774
rect 114648 42704 114860 42710
rect 115056 42910 115268 42916
rect 115056 42846 115062 42910
rect 115126 42846 115268 42910
rect 21216 42568 21972 42644
rect 27336 42644 27412 42704
rect 109344 42644 109420 42704
rect 115056 42644 115268 42846
rect 21624 42508 21700 42568
rect 1224 42502 1980 42508
rect 1224 42438 1230 42502
rect 1294 42438 1980 42502
rect 1224 42432 1980 42438
rect 1768 42408 1980 42432
rect 1768 42352 1794 42408
rect 1850 42352 1980 42408
rect 1768 42296 1980 42352
rect 20808 42502 21020 42508
rect 20808 42438 20814 42502
rect 20878 42438 21020 42502
rect 20808 42366 21020 42438
rect 20808 42302 20950 42366
rect 21014 42302 21020 42366
rect 20808 42296 21020 42302
rect 21216 42432 21972 42508
rect 21216 42296 21428 42432
rect 21624 42366 21972 42432
rect 21624 42302 21766 42366
rect 21830 42302 21972 42366
rect 21624 42296 21972 42302
rect 22032 42502 22244 42508
rect 22032 42438 22174 42502
rect 22238 42438 22244 42502
rect 22032 42366 22244 42438
rect 22032 42302 22174 42366
rect 22238 42302 22244 42366
rect 22032 42296 22244 42302
rect 22440 42502 22652 42508
rect 22440 42438 22446 42502
rect 22510 42438 22652 42502
rect 22440 42366 22652 42438
rect 27336 42432 27684 42644
rect 109344 42638 109556 42644
rect 109344 42574 109350 42638
rect 109414 42574 109556 42638
rect 109344 42432 109556 42574
rect 115056 42568 115404 42644
rect 115056 42508 115132 42568
rect 115328 42508 115404 42568
rect 115464 42568 115676 42916
rect 115872 42910 116084 42916
rect 115872 42846 116014 42910
rect 116078 42846 116084 42910
rect 115872 42774 116084 42846
rect 115872 42710 115878 42774
rect 115942 42710 116084 42774
rect 115872 42704 116084 42710
rect 115464 42508 115540 42568
rect 114240 42502 114452 42508
rect 114240 42438 114246 42502
rect 114310 42438 114452 42502
rect 27472 42372 27548 42432
rect 109344 42372 109420 42432
rect 22440 42302 22582 42366
rect 22646 42302 22652 42366
rect 22440 42296 22652 42302
rect 20808 42094 21020 42100
rect 20808 42030 20950 42094
rect 21014 42030 21020 42094
rect 20808 41958 21020 42030
rect 20808 41894 20814 41958
rect 20878 41894 21020 41958
rect 20808 41888 21020 41894
rect 21216 41958 21428 42100
rect 21216 41894 21222 41958
rect 21286 41894 21428 41958
rect 21216 41888 21428 41894
rect 21624 42094 21972 42100
rect 21624 42030 21766 42094
rect 21830 42030 21972 42094
rect 21624 41958 21972 42030
rect 21624 41894 21630 41958
rect 21694 41894 21972 41958
rect 21624 41888 21972 41894
rect 22032 42094 22244 42100
rect 22032 42030 22174 42094
rect 22238 42030 22244 42094
rect 22032 41958 22244 42030
rect 22032 41894 22038 41958
rect 22102 41894 22244 41958
rect 22032 41888 22244 41894
rect 22440 42094 22652 42100
rect 22440 42030 22582 42094
rect 22646 42030 22652 42094
rect 22440 41958 22652 42030
rect 22440 41894 22446 41958
rect 22510 41894 22652 41958
rect 22440 41888 22652 41894
rect 27336 41888 27684 42372
rect 27608 41828 27684 41888
rect 20808 41686 21020 41692
rect 20808 41622 20814 41686
rect 20878 41622 21020 41686
rect 20808 41550 21020 41622
rect 20808 41486 20814 41550
rect 20878 41486 21020 41550
rect 20808 41480 21020 41486
rect 21216 41686 21428 41692
rect 21216 41622 21222 41686
rect 21286 41622 21428 41686
rect 21216 41550 21428 41622
rect 21216 41486 21358 41550
rect 21422 41486 21428 41550
rect 21216 41480 21428 41486
rect 21624 41686 21972 41692
rect 21624 41622 21630 41686
rect 21694 41622 21972 41686
rect 21624 41480 21972 41622
rect 22032 41686 22244 41692
rect 22032 41622 22038 41686
rect 22102 41622 22244 41686
rect 22032 41550 22244 41622
rect 22032 41486 22038 41550
rect 22102 41486 22244 41550
rect 22032 41480 22244 41486
rect 22440 41686 22652 41692
rect 22440 41622 22446 41686
rect 22510 41622 22652 41686
rect 22440 41550 22652 41622
rect 27336 41616 27684 41828
rect 27608 41556 27684 41616
rect 22440 41486 22582 41550
rect 22646 41486 22652 41550
rect 22440 41480 22652 41486
rect 21624 41420 21700 41480
rect 21352 41344 21700 41420
rect 27336 41344 27684 41556
rect 109344 41888 109556 42372
rect 114240 42366 114452 42438
rect 114240 42302 114246 42366
rect 114310 42302 114452 42366
rect 114240 42296 114452 42302
rect 114648 42502 114860 42508
rect 114648 42438 114790 42502
rect 114854 42438 114860 42502
rect 114648 42366 114860 42438
rect 114648 42302 114654 42366
rect 114718 42302 114860 42366
rect 114648 42296 114860 42302
rect 115056 42366 115268 42508
rect 115328 42432 115676 42508
rect 115056 42302 115062 42366
rect 115126 42302 115268 42366
rect 115056 42296 115268 42302
rect 115464 42296 115676 42432
rect 115872 42502 116084 42508
rect 115872 42438 115878 42502
rect 115942 42438 116084 42502
rect 115872 42366 116084 42438
rect 115872 42302 116014 42366
rect 116078 42302 116084 42366
rect 115872 42296 116084 42302
rect 134776 42408 134988 42508
rect 134776 42352 134844 42408
rect 134900 42372 134988 42408
rect 134900 42366 135396 42372
rect 134900 42352 135326 42366
rect 134776 42302 135326 42352
rect 135390 42302 135396 42366
rect 134776 42296 135396 42302
rect 114240 42094 114452 42100
rect 114240 42030 114246 42094
rect 114310 42030 114452 42094
rect 114240 41958 114452 42030
rect 114240 41894 114382 41958
rect 114446 41894 114452 41958
rect 114240 41888 114452 41894
rect 114648 42094 114860 42100
rect 114648 42030 114654 42094
rect 114718 42030 114860 42094
rect 114648 41958 114860 42030
rect 114648 41894 114790 41958
rect 114854 41894 114860 41958
rect 114648 41888 114860 41894
rect 115056 42094 115268 42100
rect 115056 42030 115062 42094
rect 115126 42030 115268 42094
rect 115056 41958 115268 42030
rect 115464 41964 115676 42100
rect 115366 41958 115676 41964
rect 115056 41894 115198 41958
rect 115262 41894 115268 41958
rect 115328 41894 115334 41958
rect 115398 41894 115676 41958
rect 115056 41888 115268 41894
rect 115366 41888 115676 41894
rect 115872 42094 116084 42100
rect 115872 42030 116014 42094
rect 116078 42030 116084 42094
rect 115872 41958 116084 42030
rect 115872 41894 115878 41958
rect 115942 41894 116084 41958
rect 115872 41888 116084 41894
rect 109344 41828 109420 41888
rect 109344 41616 109556 41828
rect 114240 41686 114452 41692
rect 114240 41622 114382 41686
rect 114446 41622 114452 41686
rect 109344 41556 109420 41616
rect 109344 41344 109556 41556
rect 114240 41550 114452 41622
rect 114240 41486 114382 41550
rect 114446 41486 114452 41550
rect 114240 41480 114452 41486
rect 114648 41686 114860 41692
rect 114648 41622 114790 41686
rect 114854 41622 114860 41686
rect 114648 41550 114860 41622
rect 114648 41486 114790 41550
rect 114854 41486 114860 41550
rect 114648 41480 114860 41486
rect 115056 41686 115404 41692
rect 115056 41622 115198 41686
rect 115262 41622 115334 41686
rect 115398 41622 115404 41686
rect 115056 41616 115404 41622
rect 115056 41556 115268 41616
rect 115464 41556 115676 41692
rect 115056 41550 115676 41556
rect 115056 41486 115606 41550
rect 115670 41486 115676 41550
rect 115056 41480 115676 41486
rect 115872 41686 116084 41692
rect 115872 41622 115878 41686
rect 115942 41622 116084 41686
rect 115872 41550 116084 41622
rect 115872 41486 116014 41550
rect 116078 41486 116084 41550
rect 115872 41480 116084 41486
rect 21352 41284 21428 41344
rect 27608 41284 27684 41344
rect 109480 41284 109556 41344
rect 20808 41278 21020 41284
rect 20808 41214 20814 41278
rect 20878 41214 21020 41278
rect 20808 41142 21020 41214
rect 20808 41078 20814 41142
rect 20878 41078 21020 41142
rect 20808 41072 21020 41078
rect 21216 41278 21972 41284
rect 21216 41214 21358 41278
rect 21422 41214 21972 41278
rect 21216 41208 21972 41214
rect 21216 41072 21428 41208
rect 21624 41142 21972 41208
rect 21624 41078 21766 41142
rect 21830 41078 21972 41142
rect 21624 41072 21972 41078
rect 22032 41278 22244 41284
rect 22032 41214 22038 41278
rect 22102 41214 22244 41278
rect 22032 41142 22244 41214
rect 22032 41078 22038 41142
rect 22102 41078 22244 41142
rect 22032 41072 22244 41078
rect 22440 41278 22652 41284
rect 22440 41214 22582 41278
rect 22646 41214 22652 41278
rect 22440 41142 22652 41214
rect 22440 41078 22446 41142
rect 22510 41078 22652 41142
rect 22440 41072 22652 41078
rect 27336 41072 27684 41284
rect 109344 41072 109556 41284
rect 114240 41278 114452 41284
rect 114240 41214 114382 41278
rect 114446 41214 114452 41278
rect 114240 41142 114452 41214
rect 114240 41078 114382 41142
rect 114446 41078 114452 41142
rect 114240 41072 114452 41078
rect 114648 41278 114860 41284
rect 114648 41214 114790 41278
rect 114854 41214 114860 41278
rect 114648 41142 114860 41214
rect 114648 41078 114654 41142
rect 114718 41078 114860 41142
rect 114648 41072 114860 41078
rect 115056 41142 115268 41284
rect 115464 41278 115676 41284
rect 115464 41214 115606 41278
rect 115670 41214 115676 41278
rect 115464 41148 115676 41214
rect 115366 41142 115676 41148
rect 115056 41078 115198 41142
rect 115262 41078 115268 41142
rect 115328 41078 115334 41142
rect 115398 41078 115470 41142
rect 115534 41078 115676 41142
rect 115056 41072 115268 41078
rect 115366 41072 115676 41078
rect 115872 41278 116084 41284
rect 115872 41214 116014 41278
rect 116078 41214 116084 41278
rect 115872 41142 116084 41214
rect 115872 41078 116014 41142
rect 116078 41078 116084 41142
rect 115872 41072 116084 41078
rect 27472 41012 27548 41072
rect 109480 41012 109556 41072
rect 1224 40870 1980 40876
rect 1224 40806 1230 40870
rect 1294 40806 1980 40870
rect 1224 40800 1980 40806
rect 1768 40728 1980 40800
rect 1768 40672 1794 40728
rect 1850 40672 1980 40728
rect 1768 40528 1980 40672
rect 20808 40870 21020 40876
rect 20808 40806 20814 40870
rect 20878 40806 21020 40870
rect 20808 40664 21020 40806
rect 21216 40734 21428 40876
rect 21216 40670 21222 40734
rect 21286 40670 21428 40734
rect 21216 40664 21428 40670
rect 21624 40870 21972 40876
rect 21624 40806 21766 40870
rect 21830 40806 21972 40870
rect 21624 40734 21972 40806
rect 21624 40670 21630 40734
rect 21694 40670 21972 40734
rect 21624 40664 21972 40670
rect 22032 40870 22244 40876
rect 22032 40806 22038 40870
rect 22102 40806 22244 40870
rect 22032 40734 22244 40806
rect 22032 40670 22038 40734
rect 22102 40670 22244 40734
rect 22032 40664 22244 40670
rect 22440 40870 22652 40876
rect 22440 40806 22446 40870
rect 22510 40806 22652 40870
rect 22440 40734 22652 40806
rect 22440 40670 22582 40734
rect 22646 40670 22652 40734
rect 22440 40664 22652 40670
rect 27336 40800 27684 41012
rect 109344 40800 109556 41012
rect 114240 40870 114452 40876
rect 114240 40806 114382 40870
rect 114446 40806 114452 40870
rect 27336 40740 27412 40800
rect 109344 40740 109420 40800
rect 20808 40604 20884 40664
rect 20808 40256 21020 40604
rect 27336 40598 27684 40740
rect 27336 40534 27478 40598
rect 27542 40534 27684 40598
rect 27336 40528 27684 40534
rect 109344 40598 109556 40740
rect 114240 40734 114452 40806
rect 114240 40670 114382 40734
rect 114446 40670 114452 40734
rect 114240 40664 114452 40670
rect 114648 40870 114860 40876
rect 114648 40806 114654 40870
rect 114718 40806 114860 40870
rect 114648 40734 114860 40806
rect 114648 40670 114654 40734
rect 114718 40670 114860 40734
rect 114648 40664 114860 40670
rect 115056 40870 115404 40876
rect 115056 40806 115198 40870
rect 115262 40806 115334 40870
rect 115398 40806 115404 40870
rect 115056 40800 115404 40806
rect 115464 40870 115676 40876
rect 115464 40806 115470 40870
rect 115534 40806 115676 40870
rect 115056 40664 115268 40800
rect 115464 40740 115676 40806
rect 115366 40734 115676 40740
rect 115328 40670 115334 40734
rect 115398 40670 115676 40734
rect 115366 40664 115676 40670
rect 115872 40870 116084 40876
rect 115872 40806 116014 40870
rect 116078 40806 116084 40870
rect 115872 40664 116084 40806
rect 134776 40870 135396 40876
rect 134776 40806 135326 40870
rect 135390 40806 135396 40870
rect 134776 40800 135396 40806
rect 134776 40728 134988 40800
rect 134776 40672 134844 40728
rect 134900 40672 134988 40728
rect 109344 40534 109486 40598
rect 109550 40534 109556 40598
rect 109344 40528 109556 40534
rect 115872 40604 115948 40664
rect 27472 40468 27548 40528
rect 109344 40468 109420 40528
rect 21216 40462 21428 40468
rect 21216 40398 21222 40462
rect 21286 40398 21428 40462
rect 21216 40256 21428 40398
rect 21624 40462 21972 40468
rect 21624 40398 21630 40462
rect 21694 40398 21972 40462
rect 21624 40332 21972 40398
rect 21488 40256 21972 40332
rect 22032 40462 22244 40468
rect 22032 40398 22038 40462
rect 22102 40398 22244 40462
rect 22032 40326 22244 40398
rect 22032 40262 22174 40326
rect 22238 40262 22244 40326
rect 22032 40256 22244 40262
rect 22440 40462 22652 40468
rect 22440 40398 22582 40462
rect 22646 40398 22652 40462
rect 22440 40326 22652 40398
rect 22440 40262 22446 40326
rect 22510 40262 22652 40326
rect 22440 40256 22652 40262
rect 27336 40326 27684 40468
rect 27336 40262 27478 40326
rect 27542 40262 27684 40326
rect 20808 40196 20884 40256
rect 21216 40196 21292 40256
rect 21488 40196 21564 40256
rect 20808 39848 21020 40196
rect 21216 40120 21564 40196
rect 21216 39924 21428 40120
rect 21624 39924 21972 40196
rect 21216 39918 21972 39924
rect 21216 39854 21766 39918
rect 21830 39854 21972 39918
rect 21216 39848 21972 39854
rect 22032 40054 22244 40060
rect 22032 39990 22174 40054
rect 22238 39990 22244 40054
rect 22032 39918 22244 39990
rect 22032 39854 22038 39918
rect 22102 39854 22244 39918
rect 22032 39848 22244 39854
rect 22440 40054 22652 40060
rect 22440 39990 22446 40054
rect 22510 39990 22652 40054
rect 22440 39918 22652 39990
rect 27336 39984 27684 40262
rect 109344 40326 109556 40468
rect 109344 40262 109350 40326
rect 109414 40262 109486 40326
rect 109550 40262 109556 40326
rect 109344 39984 109556 40262
rect 114240 40462 114452 40468
rect 114240 40398 114382 40462
rect 114446 40398 114452 40462
rect 114240 40326 114452 40398
rect 114240 40262 114246 40326
rect 114310 40262 114452 40326
rect 114240 40256 114452 40262
rect 114648 40462 114860 40468
rect 114648 40398 114654 40462
rect 114718 40398 114860 40462
rect 114648 40326 114860 40398
rect 114648 40262 114654 40326
rect 114718 40262 114860 40326
rect 114648 40256 114860 40262
rect 115056 40462 115404 40468
rect 115056 40398 115334 40462
rect 115398 40398 115404 40462
rect 115056 40392 115404 40398
rect 115056 40332 115268 40392
rect 115464 40332 115676 40468
rect 115056 40326 115676 40332
rect 115056 40262 115198 40326
rect 115262 40262 115676 40326
rect 115056 40256 115676 40262
rect 115872 40256 116084 40604
rect 134776 40528 134988 40672
rect 115192 40196 115268 40256
rect 115872 40196 115948 40256
rect 114240 40054 114452 40060
rect 114240 39990 114246 40054
rect 114310 39990 114452 40054
rect 27608 39924 27684 39984
rect 22440 39854 22582 39918
rect 22646 39854 22652 39918
rect 22440 39848 22652 39854
rect 20808 39788 20884 39848
rect 20808 39646 21020 39788
rect 27336 39712 27684 39924
rect 27608 39652 27684 39712
rect 20808 39582 20814 39646
rect 20878 39582 21020 39646
rect 20808 39576 21020 39582
rect 21216 39440 21428 39652
rect 21624 39646 21972 39652
rect 21624 39582 21766 39646
rect 21830 39582 21972 39646
rect 21624 39516 21972 39582
rect 21488 39440 21972 39516
rect 21216 39380 21292 39440
rect 21488 39380 21564 39440
rect 21896 39380 21972 39440
rect 20808 39374 21020 39380
rect 20808 39310 20814 39374
rect 20878 39310 21020 39374
rect 20808 39238 21020 39310
rect 20808 39174 20814 39238
rect 20878 39174 21020 39238
rect 20808 39168 21020 39174
rect 21216 39304 21564 39380
rect 21216 39168 21428 39304
rect 21624 39244 21972 39380
rect 21526 39238 21972 39244
rect 21488 39174 21494 39238
rect 21558 39174 21972 39238
rect 21526 39168 21972 39174
rect 22032 39646 22244 39652
rect 22032 39582 22038 39646
rect 22102 39582 22244 39646
rect 22032 39440 22244 39582
rect 22440 39646 22652 39652
rect 22440 39582 22582 39646
rect 22646 39582 22652 39646
rect 22440 39440 22652 39582
rect 22032 39380 22108 39440
rect 22576 39380 22652 39440
rect 21352 39108 21428 39168
rect 1224 39102 1980 39108
rect 1224 39038 1230 39102
rect 1294 39048 1980 39102
rect 1294 39038 1794 39048
rect 1224 39032 1794 39038
rect 1768 38992 1794 39032
rect 1850 38992 1980 39048
rect 21352 39032 21700 39108
rect 1768 38896 1980 38992
rect 21624 38972 21700 39032
rect 22032 39032 22244 39380
rect 22440 39032 22652 39380
rect 27336 39374 27684 39652
rect 27336 39310 27478 39374
rect 27542 39310 27684 39374
rect 27336 39304 27684 39310
rect 109344 39918 109556 39924
rect 109344 39854 109350 39918
rect 109414 39854 109556 39918
rect 109344 39712 109556 39854
rect 114240 39918 114452 39990
rect 114240 39854 114246 39918
rect 114310 39854 114452 39918
rect 114240 39848 114452 39854
rect 114648 40054 114860 40060
rect 114648 39990 114654 40054
rect 114718 39990 114860 40054
rect 114648 39918 114860 39990
rect 114648 39854 114654 39918
rect 114718 39854 114860 39918
rect 114648 39848 114860 39854
rect 115056 39918 115268 40196
rect 115366 40190 115676 40196
rect 115328 40126 115334 40190
rect 115398 40126 115676 40190
rect 115366 40120 115676 40126
rect 115056 39854 115198 39918
rect 115262 39854 115268 39918
rect 115056 39848 115268 39854
rect 115464 39848 115676 40120
rect 115872 39848 116084 40196
rect 115872 39788 115948 39848
rect 109344 39652 109420 39712
rect 109344 39374 109556 39652
rect 114240 39646 114452 39652
rect 114240 39582 114246 39646
rect 114310 39582 114452 39646
rect 114240 39440 114452 39582
rect 114648 39646 114860 39652
rect 114648 39582 114654 39646
rect 114718 39582 114860 39646
rect 114648 39440 114860 39582
rect 115056 39646 115268 39652
rect 115056 39582 115198 39646
rect 115262 39582 115268 39646
rect 115056 39440 115268 39582
rect 115464 39516 115676 39652
rect 115872 39646 116084 39788
rect 115872 39582 115878 39646
rect 115942 39582 116084 39646
rect 115872 39576 116084 39582
rect 114376 39380 114452 39440
rect 114784 39380 114860 39440
rect 115192 39380 115268 39440
rect 115328 39440 115676 39516
rect 115328 39380 115404 39440
rect 115600 39380 115676 39440
rect 109344 39310 109486 39374
rect 109550 39310 109556 39374
rect 109344 39304 109556 39310
rect 27336 39102 27684 39108
rect 27336 39038 27478 39102
rect 27542 39038 27684 39102
rect 22032 38972 22108 39032
rect 22440 38972 22516 39032
rect 20808 38966 21020 38972
rect 20808 38902 20814 38966
rect 20878 38902 21020 38966
rect 20808 38830 21020 38902
rect 20808 38766 20814 38830
rect 20878 38766 21020 38830
rect 20808 38760 21020 38766
rect 21216 38966 21564 38972
rect 21216 38902 21494 38966
rect 21558 38902 21564 38966
rect 21216 38896 21564 38902
rect 21216 38624 21428 38896
rect 21624 38624 21972 38972
rect 21896 38564 21972 38624
rect 20808 38558 21020 38564
rect 20808 38494 20814 38558
rect 20878 38494 21020 38558
rect 20808 38422 21020 38494
rect 20808 38358 20814 38422
rect 20878 38358 21020 38422
rect 20808 38352 21020 38358
rect 21216 38422 21428 38564
rect 21216 38358 21358 38422
rect 21422 38358 21428 38422
rect 21216 38352 21428 38358
rect 21624 38352 21972 38564
rect 22032 38624 22244 38972
rect 22440 38624 22652 38972
rect 22032 38564 22108 38624
rect 22576 38564 22652 38624
rect 22032 38422 22244 38564
rect 22032 38358 22038 38422
rect 22102 38358 22244 38422
rect 22032 38352 22244 38358
rect 22440 38422 22652 38564
rect 27336 38488 27684 39038
rect 109344 39102 109556 39108
rect 109344 39038 109486 39102
rect 109550 39038 109556 39102
rect 109344 38488 109556 39038
rect 114240 39032 114452 39380
rect 114648 39032 114860 39380
rect 115056 39304 115404 39380
rect 115056 39168 115268 39304
rect 115464 39238 115676 39380
rect 115464 39174 115470 39238
rect 115534 39174 115676 39238
rect 115464 39168 115676 39174
rect 115872 39374 116084 39380
rect 115872 39310 115878 39374
rect 115942 39310 116084 39374
rect 115872 39238 116084 39310
rect 115872 39174 116014 39238
rect 116078 39174 116084 39238
rect 115872 39168 116084 39174
rect 134776 39102 135396 39108
rect 134776 39048 135326 39102
rect 114240 38972 114316 39032
rect 114648 38972 114724 39032
rect 134776 38992 134844 39048
rect 134900 39038 135326 39048
rect 135390 39038 135396 39102
rect 134900 39032 135396 39038
rect 134900 38992 134988 39032
rect 114240 38624 114452 38972
rect 114648 38624 114860 38972
rect 115056 38624 115268 38972
rect 114240 38564 114316 38624
rect 114784 38564 114860 38624
rect 115192 38564 115268 38624
rect 115464 38966 115676 38972
rect 115464 38902 115470 38966
rect 115534 38902 115676 38966
rect 115464 38624 115676 38902
rect 115872 38966 116084 38972
rect 115872 38902 116014 38966
rect 116078 38902 116084 38966
rect 115872 38830 116084 38902
rect 134776 38896 134988 38992
rect 115872 38766 116014 38830
rect 116078 38766 116084 38830
rect 115872 38760 116084 38766
rect 115464 38564 115540 38624
rect 27472 38428 27548 38488
rect 109344 38428 109420 38488
rect 22440 38358 22446 38422
rect 22510 38358 22652 38422
rect 22440 38352 22652 38358
rect 21624 38292 21700 38352
rect 21352 38216 21700 38292
rect 21352 38156 21428 38216
rect 20808 38150 21020 38156
rect 20808 38086 20814 38150
rect 20878 38086 21020 38150
rect 20808 38014 21020 38086
rect 20808 37950 20950 38014
rect 21014 37950 21020 38014
rect 20808 37944 21020 37950
rect 21216 38150 21972 38156
rect 21216 38086 21358 38150
rect 21422 38086 21972 38150
rect 21216 38080 21972 38086
rect 21216 37944 21428 38080
rect 21624 38014 21972 38080
rect 21624 37950 21766 38014
rect 21830 37950 21972 38014
rect 21624 37944 21972 37950
rect 22032 38150 22244 38156
rect 22032 38086 22038 38150
rect 22102 38086 22244 38150
rect 22032 38014 22244 38086
rect 22032 37950 22174 38014
rect 22238 37950 22244 38014
rect 22032 37944 22244 37950
rect 22440 38150 22652 38156
rect 22440 38086 22446 38150
rect 22510 38086 22652 38150
rect 22440 38014 22652 38086
rect 22440 37950 22446 38014
rect 22510 37950 22652 38014
rect 22440 37944 22652 37950
rect 27336 38150 27684 38428
rect 27336 38086 27342 38150
rect 27406 38086 27684 38150
rect 27336 37944 27684 38086
rect 109344 38150 109556 38428
rect 114240 38422 114452 38564
rect 114240 38358 114382 38422
rect 114446 38358 114452 38422
rect 114240 38352 114452 38358
rect 114648 38422 114860 38564
rect 114648 38358 114654 38422
rect 114718 38358 114860 38422
rect 114648 38352 114860 38358
rect 115056 38488 115676 38564
rect 115056 38428 115268 38488
rect 115056 38422 115404 38428
rect 115056 38358 115198 38422
rect 115262 38358 115334 38422
rect 115398 38358 115404 38422
rect 115056 38352 115404 38358
rect 115464 38352 115676 38488
rect 115872 38558 116084 38564
rect 115872 38494 116014 38558
rect 116078 38494 116084 38558
rect 115872 38422 116084 38494
rect 115872 38358 115878 38422
rect 115942 38358 116084 38422
rect 115872 38352 116084 38358
rect 109344 38086 109486 38150
rect 109550 38086 109556 38150
rect 109344 37944 109556 38086
rect 114240 38150 114452 38156
rect 114240 38086 114382 38150
rect 114446 38086 114452 38150
rect 114240 38014 114452 38086
rect 114240 37950 114246 38014
rect 114310 37950 114452 38014
rect 114240 37944 114452 37950
rect 114648 38150 114860 38156
rect 114648 38086 114654 38150
rect 114718 38086 114860 38150
rect 114648 38014 114860 38086
rect 114648 37950 114654 38014
rect 114718 37950 114860 38014
rect 114648 37944 114860 37950
rect 115056 38150 115268 38156
rect 115366 38150 115676 38156
rect 115056 38086 115198 38150
rect 115262 38086 115268 38150
rect 115328 38086 115334 38150
rect 115398 38086 115676 38150
rect 115056 38014 115268 38086
rect 115366 38080 115676 38086
rect 115056 37950 115062 38014
rect 115126 37950 115268 38014
rect 115056 37944 115268 37950
rect 115464 38014 115676 38080
rect 115464 37950 115470 38014
rect 115534 37950 115676 38014
rect 115464 37944 115676 37950
rect 115872 38150 116084 38156
rect 115872 38086 115878 38150
rect 115942 38086 116084 38150
rect 115872 38014 116084 38086
rect 115872 37950 116014 38014
rect 116078 37950 116084 38014
rect 115872 37944 116084 37950
rect 27336 37884 27412 37944
rect 109480 37884 109556 37944
rect 27336 37878 27684 37884
rect 27336 37814 27342 37878
rect 27406 37814 27684 37878
rect 14008 37606 14220 37748
rect 14008 37542 14150 37606
rect 14214 37542 14220 37606
rect 14008 37536 14220 37542
rect 20808 37742 21020 37748
rect 20808 37678 20950 37742
rect 21014 37678 21020 37742
rect 20808 37606 21020 37678
rect 20808 37542 20814 37606
rect 20878 37542 21020 37606
rect 20808 37536 21020 37542
rect 21216 37606 21428 37748
rect 21216 37542 21222 37606
rect 21286 37542 21428 37606
rect 21216 37536 21428 37542
rect 21624 37742 21972 37748
rect 21624 37678 21766 37742
rect 21830 37678 21972 37742
rect 21624 37606 21972 37678
rect 21624 37542 21630 37606
rect 21694 37542 21972 37606
rect 21624 37536 21972 37542
rect 22032 37742 22244 37748
rect 22032 37678 22174 37742
rect 22238 37678 22244 37742
rect 22032 37606 22244 37678
rect 22032 37542 22038 37606
rect 22102 37542 22244 37606
rect 22032 37536 22244 37542
rect 22440 37742 22652 37748
rect 22440 37678 22446 37742
rect 22510 37678 22652 37742
rect 22440 37606 22652 37678
rect 27336 37672 27684 37814
rect 27608 37612 27684 37672
rect 22440 37542 22582 37606
rect 22646 37542 22652 37606
rect 22440 37536 22652 37542
rect 1768 37368 1980 37476
rect 1768 37340 1794 37368
rect 1224 37334 1794 37340
rect 1224 37270 1230 37334
rect 1294 37312 1794 37334
rect 1850 37312 1980 37368
rect 27336 37400 27684 37612
rect 109344 37878 109556 37884
rect 109344 37814 109486 37878
rect 109550 37814 109556 37878
rect 109344 37672 109556 37814
rect 114240 37742 114452 37748
rect 114240 37678 114246 37742
rect 114310 37678 114452 37742
rect 109344 37612 109420 37672
rect 109344 37400 109556 37612
rect 114240 37606 114452 37678
rect 114240 37542 114382 37606
rect 114446 37542 114452 37606
rect 114240 37536 114452 37542
rect 114648 37742 114860 37748
rect 114648 37678 114654 37742
rect 114718 37678 114860 37742
rect 114648 37606 114860 37678
rect 114648 37542 114790 37606
rect 114854 37542 114860 37606
rect 114648 37536 114860 37542
rect 115056 37742 115268 37748
rect 115056 37678 115062 37742
rect 115126 37678 115268 37742
rect 115056 37536 115268 37678
rect 115464 37742 115676 37748
rect 115464 37678 115470 37742
rect 115534 37678 115676 37742
rect 115464 37536 115676 37678
rect 115872 37742 116084 37748
rect 115872 37678 116014 37742
rect 116078 37678 116084 37742
rect 115872 37606 116084 37678
rect 115872 37542 115878 37606
rect 115942 37542 116084 37606
rect 115872 37536 116084 37542
rect 115464 37476 115540 37536
rect 115192 37400 115540 37476
rect 134776 37470 135396 37476
rect 134776 37406 135326 37470
rect 135390 37406 135396 37470
rect 134776 37400 135396 37406
rect 27336 37340 27412 37400
rect 109344 37340 109420 37400
rect 115192 37340 115268 37400
rect 134776 37368 134988 37400
rect 1294 37270 1980 37312
rect 1224 37264 1980 37270
rect 20808 37334 21020 37340
rect 20808 37270 20814 37334
rect 20878 37270 21020 37334
rect 20808 37198 21020 37270
rect 20808 37134 20814 37198
rect 20878 37134 21020 37198
rect 20808 37128 21020 37134
rect 21216 37334 21428 37340
rect 21216 37270 21222 37334
rect 21286 37270 21428 37334
rect 21216 37198 21428 37270
rect 21624 37334 21972 37340
rect 21624 37270 21630 37334
rect 21694 37270 21972 37334
rect 21624 37204 21972 37270
rect 21526 37198 21972 37204
rect 21216 37134 21358 37198
rect 21422 37134 21428 37198
rect 21488 37134 21494 37198
rect 21558 37134 21972 37198
rect 21216 37128 21428 37134
rect 21526 37128 21972 37134
rect 22032 37334 22244 37340
rect 22032 37270 22038 37334
rect 22102 37270 22244 37334
rect 22032 37198 22244 37270
rect 22032 37134 22174 37198
rect 22238 37134 22244 37198
rect 22032 37128 22244 37134
rect 22440 37334 22652 37340
rect 22440 37270 22582 37334
rect 22646 37270 22652 37334
rect 22440 37198 22652 37270
rect 22440 37134 22582 37198
rect 22646 37134 22652 37198
rect 22440 37128 22652 37134
rect 27336 37128 27684 37340
rect 27608 37068 27684 37128
rect 0 36856 13812 36932
rect 20808 36926 21020 36932
rect 13600 36822 13812 36856
rect 14608 36895 14674 36898
rect 15342 36895 15408 36898
rect 14608 36893 15408 36895
rect 14608 36837 14613 36893
rect 14669 36837 15347 36893
rect 15403 36837 15408 36893
rect 14608 36835 15408 36837
rect 14608 36832 14674 36835
rect 15342 36832 15408 36835
rect 20808 36862 20814 36926
rect 20878 36862 21020 36926
rect 13600 36766 13668 36822
rect 13724 36766 13812 36822
rect 13600 36720 13812 36766
rect 20808 36720 21020 36862
rect 21216 36926 21564 36932
rect 21216 36862 21358 36926
rect 21422 36862 21494 36926
rect 21558 36862 21564 36926
rect 21216 36856 21564 36862
rect 21216 36796 21428 36856
rect 21624 36796 21972 36932
rect 21216 36790 21972 36796
rect 21216 36726 21766 36790
rect 21830 36726 21972 36790
rect 21216 36720 21972 36726
rect 22032 36926 22244 36932
rect 22032 36862 22174 36926
rect 22238 36862 22244 36926
rect 22032 36790 22244 36862
rect 22032 36726 22038 36790
rect 22102 36726 22244 36790
rect 22032 36720 22244 36726
rect 22440 36926 22652 36932
rect 22440 36862 22582 36926
rect 22646 36862 22652 36926
rect 22440 36790 22652 36862
rect 27336 36856 27684 37068
rect 109344 37128 109556 37340
rect 114240 37334 114452 37340
rect 114240 37270 114382 37334
rect 114446 37270 114452 37334
rect 114240 37198 114452 37270
rect 114240 37134 114246 37198
rect 114310 37134 114452 37198
rect 114240 37128 114452 37134
rect 114648 37334 114860 37340
rect 114648 37270 114790 37334
rect 114854 37270 114860 37334
rect 114648 37198 114860 37270
rect 114648 37134 114790 37198
rect 114854 37134 114860 37198
rect 114648 37128 114860 37134
rect 115056 37264 115676 37340
rect 115056 37128 115268 37264
rect 115464 37198 115676 37264
rect 115464 37134 115606 37198
rect 115670 37134 115676 37198
rect 115464 37128 115676 37134
rect 115872 37334 116084 37340
rect 115872 37270 115878 37334
rect 115942 37270 116084 37334
rect 115872 37198 116084 37270
rect 134776 37312 134844 37368
rect 134900 37312 134988 37368
rect 134776 37264 134988 37312
rect 115872 37134 115878 37198
rect 115942 37134 116084 37198
rect 115872 37128 116084 37134
rect 109344 37068 109420 37128
rect 109344 36856 109556 37068
rect 27608 36796 27684 36856
rect 109480 36796 109556 36856
rect 22440 36726 22446 36790
rect 22510 36726 22652 36790
rect 22440 36720 22652 36726
rect 20808 36660 20884 36720
rect 14008 36252 14220 36388
rect 20808 36382 21020 36660
rect 27336 36584 27684 36796
rect 109344 36584 109556 36796
rect 114240 36926 114452 36932
rect 114240 36862 114246 36926
rect 114310 36862 114452 36926
rect 114240 36790 114452 36862
rect 114240 36726 114246 36790
rect 114310 36726 114452 36790
rect 114240 36720 114452 36726
rect 114648 36926 114860 36932
rect 114648 36862 114790 36926
rect 114854 36862 114860 36926
rect 114648 36790 114860 36862
rect 114648 36726 114654 36790
rect 114718 36726 114860 36790
rect 114648 36720 114860 36726
rect 115056 36790 115268 36932
rect 115056 36726 115198 36790
rect 115262 36726 115268 36790
rect 115056 36720 115268 36726
rect 115464 36926 115676 36932
rect 115464 36862 115606 36926
rect 115670 36862 115676 36926
rect 115464 36790 115676 36862
rect 115464 36726 115470 36790
rect 115534 36726 115676 36790
rect 115464 36720 115676 36726
rect 115872 36926 116084 36932
rect 115872 36862 115878 36926
rect 115942 36862 116084 36926
rect 115872 36720 116084 36862
rect 116008 36660 116084 36720
rect 27336 36524 27412 36584
rect 109480 36524 109556 36584
rect 20808 36318 20950 36382
rect 21014 36318 21020 36382
rect 20808 36312 21020 36318
rect 21216 36388 21428 36524
rect 21624 36518 21972 36524
rect 21624 36454 21766 36518
rect 21830 36454 21972 36518
rect 21216 36382 21564 36388
rect 21216 36318 21494 36382
rect 21558 36318 21564 36382
rect 21216 36312 21564 36318
rect 21624 36382 21972 36454
rect 21624 36318 21630 36382
rect 21694 36318 21972 36382
rect 21624 36312 21972 36318
rect 22032 36518 22244 36524
rect 22032 36454 22038 36518
rect 22102 36454 22244 36518
rect 22032 36382 22244 36454
rect 22032 36318 22038 36382
rect 22102 36318 22244 36382
rect 22032 36312 22244 36318
rect 22440 36518 22652 36524
rect 22440 36454 22446 36518
rect 22510 36454 22652 36518
rect 22440 36382 22652 36454
rect 22440 36318 22446 36382
rect 22510 36318 22652 36382
rect 22440 36312 22652 36318
rect 27336 36312 27684 36524
rect 109344 36312 109556 36524
rect 114240 36518 114452 36524
rect 114240 36454 114246 36518
rect 114310 36454 114452 36518
rect 114240 36382 114452 36454
rect 114240 36318 114382 36382
rect 114446 36318 114452 36382
rect 114240 36312 114452 36318
rect 114648 36518 114860 36524
rect 114648 36454 114654 36518
rect 114718 36454 114860 36518
rect 114648 36382 114860 36454
rect 114648 36318 114790 36382
rect 114854 36318 114860 36382
rect 114648 36312 114860 36318
rect 115056 36518 115268 36524
rect 115056 36454 115198 36518
rect 115262 36454 115268 36518
rect 115056 36382 115268 36454
rect 115464 36518 115676 36524
rect 115464 36454 115470 36518
rect 115534 36454 115676 36518
rect 115464 36388 115676 36454
rect 115366 36382 115676 36388
rect 115056 36318 115198 36382
rect 115262 36318 115268 36382
rect 115328 36318 115334 36382
rect 115398 36318 115676 36382
rect 115056 36312 115268 36318
rect 115366 36312 115676 36318
rect 115872 36382 116084 36660
rect 115872 36318 116014 36382
rect 116078 36318 116084 36382
rect 115872 36312 116084 36318
rect 27472 36252 27548 36312
rect 109344 36252 109420 36312
rect 14008 36246 14318 36252
rect 14008 36182 14286 36246
rect 14350 36182 14356 36246
rect 14008 36176 14318 36182
rect 20808 36110 21020 36116
rect 20808 36046 20950 36110
rect 21014 36046 21020 36110
rect 0 35904 2116 35980
rect 2040 35844 2116 35904
rect 20808 35904 21020 36046
rect 21216 35980 21428 36116
rect 21526 36110 21972 36116
rect 21488 36046 21494 36110
rect 21558 36046 21630 36110
rect 21694 36046 21972 36110
rect 21526 36040 21972 36046
rect 21216 35974 21564 35980
rect 21216 35910 21494 35974
rect 21558 35910 21564 35974
rect 21216 35904 21564 35910
rect 21624 35904 21972 36040
rect 22032 36110 22244 36116
rect 22032 36046 22038 36110
rect 22102 36046 22244 36110
rect 22032 35974 22244 36046
rect 22032 35910 22174 35974
rect 22238 35910 22244 35974
rect 22032 35904 22244 35910
rect 22440 36110 22652 36116
rect 22440 36046 22446 36110
rect 22510 36046 22652 36110
rect 22440 35974 22652 36046
rect 27336 36040 27684 36252
rect 109344 36040 109556 36252
rect 27472 35980 27548 36040
rect 109480 35980 109556 36040
rect 22440 35910 22446 35974
rect 22510 35910 22652 35974
rect 22440 35904 22652 35910
rect 20808 35844 20884 35904
rect 21624 35844 21700 35904
rect 2040 35768 13812 35844
rect 1773 35708 1871 35709
rect 1224 35702 1980 35708
rect 1224 35638 1230 35702
rect 1294 35688 1980 35702
rect 1294 35638 1794 35688
rect 1224 35632 1794 35638
rect 1850 35632 1980 35688
rect 1768 35496 1980 35632
rect 13600 35694 13812 35768
rect 13600 35638 13668 35694
rect 13724 35638 13812 35694
rect 13600 35496 13812 35638
rect 20808 35702 21020 35844
rect 21352 35768 21700 35844
rect 27336 35768 27684 35980
rect 109344 35768 109556 35980
rect 114240 36110 114452 36116
rect 114240 36046 114382 36110
rect 114446 36046 114452 36110
rect 114240 35974 114452 36046
rect 114240 35910 114246 35974
rect 114310 35910 114452 35974
rect 114240 35904 114452 35910
rect 114648 36110 114860 36116
rect 114648 36046 114790 36110
rect 114854 36046 114860 36110
rect 114648 35974 114860 36046
rect 114648 35910 114654 35974
rect 114718 35910 114860 35974
rect 114648 35904 114860 35910
rect 115056 36110 115404 36116
rect 115056 36046 115198 36110
rect 115262 36046 115334 36110
rect 115398 36046 115404 36110
rect 115056 36040 115404 36046
rect 115056 35980 115268 36040
rect 115464 35980 115676 36116
rect 115056 35974 115676 35980
rect 115056 35910 115470 35974
rect 115534 35910 115676 35974
rect 115056 35904 115676 35910
rect 115872 36110 116084 36116
rect 115872 36046 116014 36110
rect 116078 36046 116084 36110
rect 115872 35904 116084 36046
rect 116008 35844 116084 35904
rect 21352 35708 21428 35768
rect 27608 35708 27684 35768
rect 109480 35708 109556 35768
rect 20808 35638 20814 35702
rect 20878 35638 21020 35702
rect 20808 35632 21020 35638
rect 14608 35625 14674 35628
rect 15262 35625 15328 35628
rect 14608 35623 15328 35625
rect 14608 35567 14613 35623
rect 14669 35567 15267 35623
rect 15323 35567 15328 35623
rect 14608 35565 15328 35567
rect 14608 35562 14674 35565
rect 15262 35562 15328 35565
rect 21216 35572 21428 35708
rect 21526 35702 21972 35708
rect 21488 35638 21494 35702
rect 21558 35638 21972 35702
rect 21526 35632 21972 35638
rect 21216 35566 21564 35572
rect 21216 35502 21358 35566
rect 21422 35502 21564 35566
rect 21216 35496 21564 35502
rect 21624 35566 21972 35632
rect 21624 35502 21630 35566
rect 21694 35502 21972 35566
rect 21624 35496 21972 35502
rect 22032 35702 22244 35708
rect 22032 35638 22174 35702
rect 22238 35638 22244 35702
rect 22032 35496 22244 35638
rect 22440 35702 22652 35708
rect 22440 35638 22446 35702
rect 22510 35638 22652 35702
rect 22440 35496 22652 35638
rect 27336 35496 27684 35708
rect 109344 35496 109556 35708
rect 114240 35702 114452 35708
rect 114240 35638 114246 35702
rect 114310 35638 114452 35702
rect 114240 35496 114452 35638
rect 21216 35436 21292 35496
rect 21488 35436 21564 35496
rect 22032 35436 22108 35496
rect 22576 35436 22652 35496
rect 20808 35430 21020 35436
rect 20808 35366 20814 35430
rect 20878 35366 21020 35430
rect 20808 35294 21020 35366
rect 20808 35230 20950 35294
rect 21014 35230 21020 35294
rect 20808 35224 21020 35230
rect 21216 35224 21428 35436
rect 21488 35360 21972 35436
rect 21624 35294 21972 35360
rect 21624 35230 21902 35294
rect 21966 35230 21972 35294
rect 21624 35224 21972 35230
rect 22032 35088 22244 35436
rect 22440 35088 22652 35436
rect 27462 35300 27560 35496
rect 109344 35300 109448 35496
rect 114376 35436 114452 35496
rect 27336 35294 27684 35300
rect 27336 35230 27478 35294
rect 27542 35230 27684 35294
rect 27336 35224 27684 35230
rect 27608 35164 27684 35224
rect 22032 35028 22108 35088
rect 22576 35028 22652 35088
rect 20808 35022 21020 35028
rect 20808 34958 20950 35022
rect 21014 34958 21020 35022
rect 14008 34886 14220 34892
rect 14008 34822 14150 34886
rect 14214 34822 14220 34886
rect 14008 34750 14220 34822
rect 20808 34886 21020 34958
rect 20808 34822 20814 34886
rect 20878 34822 21020 34886
rect 20808 34816 21020 34822
rect 21216 34886 21972 34892
rect 21216 34822 21902 34886
rect 21966 34822 21972 34886
rect 21216 34816 21972 34822
rect 14008 34686 14014 34750
rect 14078 34686 14220 34750
rect 14008 34680 14220 34686
rect 21216 34680 21428 34816
rect 21624 34680 21972 34816
rect 22032 34680 22244 35028
rect 22440 34680 22652 35028
rect 21352 34620 21428 34680
rect 21760 34620 21836 34680
rect 22168 34620 22244 34680
rect 22576 34620 22652 34680
rect 20808 34614 21020 34620
rect 20808 34550 20814 34614
rect 20878 34550 21020 34614
rect 20808 34478 21020 34550
rect 20808 34414 20814 34478
rect 20878 34414 21020 34478
rect 20808 34408 21020 34414
rect 21216 34478 21428 34620
rect 21216 34414 21222 34478
rect 21286 34414 21428 34478
rect 21216 34408 21428 34414
rect 21624 34408 21972 34620
rect 22032 34478 22244 34620
rect 22032 34414 22038 34478
rect 22102 34414 22244 34478
rect 22032 34408 22244 34414
rect 22440 34478 22652 34620
rect 27336 35022 27684 35164
rect 27336 34958 27478 35022
rect 27542 34958 27684 35022
rect 27336 34544 27684 34958
rect 109344 35224 109556 35300
rect 109344 35164 109420 35224
rect 109344 35022 109556 35164
rect 109344 34958 109350 35022
rect 109414 34958 109556 35022
rect 109344 34750 109556 34958
rect 109344 34686 109350 34750
rect 109414 34686 109486 34750
rect 109550 34686 109556 34750
rect 109344 34544 109556 34686
rect 114240 35088 114452 35436
rect 114648 35702 114860 35708
rect 114648 35638 114654 35702
rect 114718 35638 114860 35702
rect 114648 35496 114860 35638
rect 115056 35496 115268 35708
rect 115464 35702 115676 35708
rect 115464 35638 115470 35702
rect 115534 35638 115676 35702
rect 115464 35496 115676 35638
rect 115872 35702 116084 35844
rect 115872 35638 115878 35702
rect 115942 35638 116084 35702
rect 115872 35632 116084 35638
rect 134776 35688 134988 35844
rect 134776 35632 134844 35688
rect 134900 35632 134988 35688
rect 134776 35572 134988 35632
rect 134776 35566 135396 35572
rect 134776 35502 135326 35566
rect 135390 35502 135396 35566
rect 134776 35496 135396 35502
rect 114648 35436 114724 35496
rect 115056 35436 115132 35496
rect 115464 35436 115540 35496
rect 114648 35088 114860 35436
rect 115056 35360 115676 35436
rect 115056 35224 115268 35360
rect 115464 35294 115676 35360
rect 115464 35230 115470 35294
rect 115534 35230 115676 35294
rect 115464 35224 115676 35230
rect 115872 35430 116084 35436
rect 115872 35366 115878 35430
rect 115942 35366 116084 35430
rect 115872 35294 116084 35366
rect 115872 35230 115878 35294
rect 115942 35230 116084 35294
rect 115872 35224 116084 35230
rect 114240 35028 114316 35088
rect 114784 35028 114860 35088
rect 114240 34680 114452 35028
rect 114648 34680 114860 35028
rect 115872 35022 116084 35028
rect 115872 34958 115878 35022
rect 115942 34958 116084 35022
rect 114240 34620 114316 34680
rect 114784 34620 114860 34680
rect 27608 34484 27684 34544
rect 22440 34414 22446 34478
rect 22510 34414 22652 34478
rect 22440 34408 22652 34414
rect 20808 34206 21020 34212
rect 20808 34142 20814 34206
rect 20878 34142 21020 34206
rect 1224 34070 1844 34076
rect 1224 34006 1230 34070
rect 1294 34029 1844 34070
rect 1294 34008 1871 34029
rect 1294 34006 1794 34008
rect 1224 34000 1794 34006
rect 1773 33952 1794 34000
rect 1850 33952 1871 34008
rect 1773 33931 1871 33952
rect 13600 33994 13812 34076
rect 20808 34070 21020 34142
rect 14608 34067 14674 34070
rect 15182 34067 15248 34070
rect 14608 34065 15248 34067
rect 14608 34009 14613 34065
rect 14669 34009 15187 34065
rect 15243 34009 15248 34065
rect 14608 34007 15248 34009
rect 14608 34004 14674 34007
rect 15182 34004 15248 34007
rect 20808 34006 20814 34070
rect 20878 34006 21020 34070
rect 20808 34000 21020 34006
rect 21216 34206 21428 34212
rect 21216 34142 21222 34206
rect 21286 34142 21428 34206
rect 21216 34070 21428 34142
rect 21216 34006 21358 34070
rect 21422 34006 21428 34070
rect 21216 34000 21428 34006
rect 21624 34000 21972 34212
rect 22032 34206 22244 34212
rect 22032 34142 22038 34206
rect 22102 34142 22244 34206
rect 22032 34070 22244 34142
rect 22032 34006 22038 34070
rect 22102 34006 22244 34070
rect 22032 34000 22244 34006
rect 22440 34206 22652 34212
rect 22440 34142 22446 34206
rect 22510 34142 22652 34206
rect 22440 34070 22652 34142
rect 22440 34006 22446 34070
rect 22510 34006 22652 34070
rect 22440 34000 22652 34006
rect 27336 34000 27684 34484
rect 109344 34478 109556 34484
rect 109344 34414 109486 34478
rect 109550 34414 109556 34478
rect 109344 34206 109556 34414
rect 114240 34478 114452 34620
rect 114240 34414 114246 34478
rect 114310 34414 114452 34478
rect 114240 34408 114452 34414
rect 114648 34478 114860 34620
rect 114648 34414 114654 34478
rect 114718 34414 114860 34478
rect 114648 34408 114860 34414
rect 115056 34680 115268 34892
rect 115464 34886 115676 34892
rect 115464 34822 115470 34886
rect 115534 34822 115676 34886
rect 115464 34680 115676 34822
rect 115872 34886 116084 34958
rect 115872 34822 116014 34886
rect 116078 34822 116084 34886
rect 115872 34816 116084 34822
rect 115056 34620 115132 34680
rect 115600 34620 115676 34680
rect 115056 34478 115268 34620
rect 115056 34414 115198 34478
rect 115262 34414 115268 34478
rect 115056 34408 115268 34414
rect 115464 34478 115676 34620
rect 115464 34414 115606 34478
rect 115670 34414 115676 34478
rect 115464 34408 115676 34414
rect 115872 34614 116084 34620
rect 115872 34550 116014 34614
rect 116078 34550 116084 34614
rect 115872 34478 116084 34550
rect 115872 34414 116014 34478
rect 116078 34414 116084 34478
rect 115872 34408 116084 34414
rect 109344 34142 109486 34206
rect 109550 34142 109556 34206
rect 109344 34000 109556 34142
rect 114240 34206 114452 34212
rect 114240 34142 114246 34206
rect 114310 34142 114452 34206
rect 114240 34070 114452 34142
rect 114240 34006 114246 34070
rect 114310 34006 114452 34070
rect 114240 34000 114452 34006
rect 114648 34206 114860 34212
rect 114648 34142 114654 34206
rect 114718 34142 114860 34206
rect 114648 34070 114860 34142
rect 114648 34006 114790 34070
rect 114854 34006 114860 34070
rect 114648 34000 114860 34006
rect 115056 34206 115268 34212
rect 115056 34142 115198 34206
rect 115262 34142 115268 34206
rect 115056 34076 115268 34142
rect 115464 34206 115676 34212
rect 115464 34142 115606 34206
rect 115670 34142 115676 34206
rect 115056 34070 115404 34076
rect 115056 34006 115334 34070
rect 115398 34006 115404 34070
rect 115056 34000 115404 34006
rect 115464 34070 115676 34142
rect 115464 34006 115606 34070
rect 115670 34006 115676 34070
rect 115464 34000 115676 34006
rect 115872 34206 116084 34212
rect 115872 34142 116014 34206
rect 116078 34142 116084 34206
rect 115872 34070 116084 34142
rect 115872 34006 116014 34070
rect 116078 34006 116084 34070
rect 115872 34000 116084 34006
rect 134776 34008 134988 34076
rect 13600 33940 13668 33994
rect 2040 33938 13668 33940
rect 13724 33938 13812 33994
rect 21624 33940 21700 34000
rect 2040 33864 13812 33938
rect 21352 33864 21700 33940
rect 27336 33940 27412 34000
rect 109344 33940 109420 34000
rect 134776 33952 134844 34008
rect 134900 33952 134988 34008
rect 134776 33940 134988 33952
rect 2040 33804 2116 33864
rect 21352 33804 21428 33864
rect 0 33728 2116 33804
rect 20808 33798 21020 33804
rect 20808 33734 20814 33798
rect 20878 33734 21020 33798
rect 20808 33662 21020 33734
rect 20808 33598 20814 33662
rect 20878 33598 21020 33662
rect 20808 33592 21020 33598
rect 21216 33798 21972 33804
rect 21216 33734 21358 33798
rect 21422 33734 21972 33798
rect 21216 33728 21972 33734
rect 21216 33662 21428 33728
rect 21216 33598 21358 33662
rect 21422 33598 21428 33662
rect 21216 33592 21428 33598
rect 21624 33662 21972 33728
rect 21624 33598 21766 33662
rect 21830 33598 21972 33662
rect 21624 33592 21972 33598
rect 22032 33798 22244 33804
rect 22032 33734 22038 33798
rect 22102 33734 22244 33798
rect 22032 33662 22244 33734
rect 22032 33598 22174 33662
rect 22238 33598 22244 33662
rect 22032 33592 22244 33598
rect 22440 33798 22652 33804
rect 22440 33734 22446 33798
rect 22510 33734 22652 33798
rect 22440 33662 22652 33734
rect 27336 33728 27684 33940
rect 109344 33934 109556 33940
rect 109344 33870 109486 33934
rect 109550 33870 109556 33934
rect 109344 33728 109556 33870
rect 134776 33934 135396 33940
rect 134776 33870 135326 33934
rect 135390 33870 135396 33934
rect 134776 33864 135396 33870
rect 27472 33668 27548 33728
rect 109480 33668 109556 33728
rect 22440 33598 22446 33662
rect 22510 33598 22652 33662
rect 22440 33592 22652 33598
rect 14008 33526 14356 33532
rect 14008 33462 14286 33526
rect 14350 33462 14356 33526
rect 14008 33456 14356 33462
rect 27336 33456 27684 33668
rect 109344 33456 109556 33668
rect 114240 33798 114452 33804
rect 114240 33734 114246 33798
rect 114310 33734 114452 33798
rect 114240 33662 114452 33734
rect 114240 33598 114246 33662
rect 114310 33598 114452 33662
rect 114240 33592 114452 33598
rect 114648 33798 114860 33804
rect 114648 33734 114790 33798
rect 114854 33734 114860 33798
rect 114648 33662 114860 33734
rect 114648 33598 114654 33662
rect 114718 33598 114860 33662
rect 114648 33592 114860 33598
rect 115056 33662 115268 33804
rect 115366 33798 115676 33804
rect 115328 33734 115334 33798
rect 115398 33734 115606 33798
rect 115670 33734 115676 33798
rect 115366 33728 115676 33734
rect 115056 33598 115062 33662
rect 115126 33598 115268 33662
rect 115056 33592 115268 33598
rect 115464 33662 115676 33728
rect 115464 33598 115606 33662
rect 115670 33598 115676 33662
rect 115464 33592 115676 33598
rect 115872 33798 116084 33804
rect 115872 33734 116014 33798
rect 116078 33734 116084 33798
rect 115872 33662 116084 33734
rect 115872 33598 116014 33662
rect 116078 33598 116084 33662
rect 115872 33592 116084 33598
rect 14008 33390 14220 33456
rect 27608 33396 27684 33456
rect 109480 33396 109556 33456
rect 14008 33326 14150 33390
rect 14214 33326 14220 33390
rect 14008 33320 14220 33326
rect 20808 33390 21020 33396
rect 20808 33326 20814 33390
rect 20878 33326 21020 33390
rect 20808 33254 21020 33326
rect 20808 33190 20814 33254
rect 20878 33190 21020 33254
rect 20808 33184 21020 33190
rect 21216 33390 21428 33396
rect 21216 33326 21358 33390
rect 21422 33326 21428 33390
rect 21216 33184 21428 33326
rect 21624 33390 21972 33396
rect 21624 33326 21766 33390
rect 21830 33326 21972 33390
rect 21624 33254 21972 33326
rect 21624 33190 21630 33254
rect 21694 33190 21972 33254
rect 21624 33184 21972 33190
rect 22032 33390 22244 33396
rect 22032 33326 22174 33390
rect 22238 33326 22244 33390
rect 22032 33254 22244 33326
rect 22032 33190 22038 33254
rect 22102 33190 22244 33254
rect 22032 33184 22244 33190
rect 22440 33390 22652 33396
rect 22440 33326 22446 33390
rect 22510 33326 22652 33390
rect 22440 33254 22652 33326
rect 22440 33190 22446 33254
rect 22510 33190 22652 33254
rect 22440 33184 22652 33190
rect 27336 33184 27684 33396
rect 109344 33184 109556 33396
rect 114240 33390 114452 33396
rect 114240 33326 114246 33390
rect 114310 33326 114452 33390
rect 114240 33254 114452 33326
rect 114240 33190 114382 33254
rect 114446 33190 114452 33254
rect 114240 33184 114452 33190
rect 114648 33390 114860 33396
rect 114648 33326 114654 33390
rect 114718 33326 114860 33390
rect 114648 33254 114860 33326
rect 114648 33190 114790 33254
rect 114854 33190 114860 33254
rect 114648 33184 114860 33190
rect 115056 33390 115268 33396
rect 115056 33326 115062 33390
rect 115126 33326 115268 33390
rect 115056 33254 115268 33326
rect 115056 33190 115198 33254
rect 115262 33190 115268 33254
rect 115056 33184 115268 33190
rect 115464 33390 115676 33396
rect 115464 33326 115606 33390
rect 115670 33326 115676 33390
rect 115464 33184 115676 33326
rect 115872 33390 116084 33396
rect 115872 33326 116014 33390
rect 116078 33326 116084 33390
rect 115872 33254 116084 33326
rect 115872 33190 115878 33254
rect 115942 33190 116084 33254
rect 115872 33184 116084 33190
rect 27472 33124 27548 33184
rect 109344 33124 109420 33184
rect 115464 33124 115540 33184
rect 13600 32866 13812 32988
rect 13600 32852 13668 32866
rect 0 32810 13668 32852
rect 13724 32810 13812 32866
rect 0 32776 13812 32810
rect 20808 32982 21020 32988
rect 20808 32918 20814 32982
rect 20878 32918 21020 32982
rect 20808 32846 21020 32918
rect 14608 32797 14674 32800
rect 15102 32797 15168 32800
rect 14608 32795 15168 32797
rect 14608 32739 14613 32795
rect 14669 32739 15107 32795
rect 15163 32739 15168 32795
rect 20808 32782 20950 32846
rect 21014 32782 21020 32846
rect 20808 32776 21020 32782
rect 21216 32846 21428 32988
rect 21216 32782 21222 32846
rect 21286 32782 21428 32846
rect 21216 32776 21428 32782
rect 21624 32982 21972 32988
rect 21624 32918 21630 32982
rect 21694 32918 21972 32982
rect 21624 32776 21972 32918
rect 22032 32982 22244 32988
rect 22032 32918 22038 32982
rect 22102 32918 22244 32982
rect 22032 32846 22244 32918
rect 22032 32782 22038 32846
rect 22102 32782 22244 32846
rect 22032 32776 22244 32782
rect 22440 32982 22652 32988
rect 22440 32918 22446 32982
rect 22510 32918 22652 32982
rect 22440 32846 22652 32918
rect 22440 32782 22582 32846
rect 22646 32782 22652 32846
rect 22440 32776 22652 32782
rect 27336 32912 27684 33124
rect 109344 32912 109556 33124
rect 115192 33048 115540 33124
rect 115192 32988 115268 33048
rect 114240 32982 114452 32988
rect 114240 32918 114382 32982
rect 114446 32918 114452 32982
rect 27336 32852 27412 32912
rect 109344 32852 109420 32912
rect 14608 32737 15168 32739
rect 14608 32734 14674 32737
rect 15102 32734 15168 32737
rect 21624 32716 21700 32776
rect 21352 32640 21700 32716
rect 27336 32640 27684 32852
rect 109344 32640 109556 32852
rect 114240 32846 114452 32918
rect 114240 32782 114382 32846
rect 114446 32782 114452 32846
rect 114240 32776 114452 32782
rect 114648 32982 114860 32988
rect 114648 32918 114790 32982
rect 114854 32918 114860 32982
rect 114648 32846 114860 32918
rect 114648 32782 114790 32846
rect 114854 32782 114860 32846
rect 114648 32776 114860 32782
rect 115056 32982 115676 32988
rect 115056 32918 115198 32982
rect 115262 32918 115676 32982
rect 115056 32912 115676 32918
rect 115056 32776 115268 32912
rect 115464 32846 115676 32912
rect 115464 32782 115606 32846
rect 115670 32782 115676 32846
rect 115464 32776 115676 32782
rect 115872 32982 116084 32988
rect 115872 32918 115878 32982
rect 115942 32918 116084 32982
rect 115872 32846 116084 32918
rect 115872 32782 115878 32846
rect 115942 32782 116084 32846
rect 115872 32776 116084 32782
rect 21352 32580 21428 32640
rect 27608 32580 27684 32640
rect 109480 32580 109556 32640
rect 20808 32574 21020 32580
rect 20808 32510 20950 32574
rect 21014 32510 21020 32574
rect 1224 32438 1980 32444
rect 1224 32374 1230 32438
rect 1294 32374 1980 32438
rect 1224 32368 1980 32374
rect 20808 32438 21020 32510
rect 20808 32374 20950 32438
rect 21014 32374 21020 32438
rect 20808 32368 21020 32374
rect 21216 32574 21972 32580
rect 21216 32510 21222 32574
rect 21286 32510 21972 32574
rect 21216 32504 21972 32510
rect 21216 32368 21428 32504
rect 21624 32438 21972 32504
rect 21624 32374 21766 32438
rect 21830 32374 21972 32438
rect 21624 32368 21972 32374
rect 22032 32574 22244 32580
rect 22032 32510 22038 32574
rect 22102 32510 22244 32574
rect 22032 32438 22244 32510
rect 22032 32374 22038 32438
rect 22102 32374 22244 32438
rect 22032 32368 22244 32374
rect 22440 32574 22652 32580
rect 22440 32510 22582 32574
rect 22646 32510 22652 32574
rect 22440 32438 22652 32510
rect 22440 32374 22446 32438
rect 22510 32374 22652 32438
rect 22440 32368 22652 32374
rect 27336 32368 27684 32580
rect 109344 32368 109556 32580
rect 114240 32574 114452 32580
rect 114240 32510 114382 32574
rect 114446 32510 114452 32574
rect 114240 32438 114452 32510
rect 114240 32374 114246 32438
rect 114310 32374 114452 32438
rect 114240 32368 114452 32374
rect 114648 32574 114860 32580
rect 114648 32510 114790 32574
rect 114854 32510 114860 32574
rect 114648 32438 114860 32510
rect 114648 32374 114654 32438
rect 114718 32374 114860 32438
rect 114648 32368 114860 32374
rect 115056 32438 115268 32580
rect 115464 32574 115676 32580
rect 115464 32510 115606 32574
rect 115670 32510 115676 32574
rect 115464 32444 115676 32510
rect 115366 32438 115676 32444
rect 115056 32374 115198 32438
rect 115262 32374 115268 32438
rect 115328 32374 115334 32438
rect 115398 32374 115676 32438
rect 115056 32368 115268 32374
rect 115366 32368 115676 32374
rect 115872 32574 116084 32580
rect 115872 32510 115878 32574
rect 115942 32510 116084 32574
rect 115872 32438 116084 32510
rect 115872 32374 115878 32438
rect 115942 32374 116084 32438
rect 115872 32368 116084 32374
rect 1768 32328 1980 32368
rect 1768 32272 1794 32328
rect 1850 32272 1980 32328
rect 27472 32308 27548 32368
rect 109480 32308 109556 32368
rect 1768 32232 1980 32272
rect 14008 32166 14220 32172
rect 14008 32102 14014 32166
rect 14078 32102 14220 32166
rect 14008 31894 14220 32102
rect 20808 32166 21020 32172
rect 20808 32102 20950 32166
rect 21014 32102 21020 32166
rect 20808 31960 21020 32102
rect 21216 32030 21428 32172
rect 21216 31966 21222 32030
rect 21286 31966 21428 32030
rect 21216 31960 21428 31966
rect 21624 32166 21972 32172
rect 21624 32102 21766 32166
rect 21830 32102 21972 32166
rect 21624 32030 21972 32102
rect 21624 31966 21630 32030
rect 21694 31966 21972 32030
rect 21624 31960 21972 31966
rect 22032 32166 22244 32172
rect 22032 32102 22038 32166
rect 22102 32102 22244 32166
rect 22032 32030 22244 32102
rect 22032 31966 22038 32030
rect 22102 31966 22244 32030
rect 22032 31960 22244 31966
rect 22440 32166 22652 32172
rect 22440 32102 22446 32166
rect 22510 32102 22652 32166
rect 22440 32030 22652 32102
rect 22440 31966 22582 32030
rect 22646 31966 22652 32030
rect 22440 31960 22652 31966
rect 27336 32096 27684 32308
rect 109344 32096 109556 32308
rect 134776 32328 134988 32444
rect 134776 32272 134844 32328
rect 134900 32308 134988 32328
rect 134900 32302 135396 32308
rect 134900 32272 135326 32302
rect 134776 32238 135326 32272
rect 135390 32238 135396 32302
rect 134776 32232 135396 32238
rect 114240 32166 114452 32172
rect 114240 32102 114246 32166
rect 114310 32102 114452 32166
rect 27336 32036 27412 32096
rect 109344 32036 109420 32096
rect 20944 31900 21020 31960
rect 14008 31830 14150 31894
rect 14214 31830 14220 31894
rect 14008 31824 14220 31830
rect 20808 31758 21020 31900
rect 27336 31824 27684 32036
rect 109344 31894 109556 32036
rect 114240 32030 114452 32102
rect 114240 31966 114382 32030
rect 114446 31966 114452 32030
rect 114240 31960 114452 31966
rect 114648 32166 114860 32172
rect 114648 32102 114654 32166
rect 114718 32102 114860 32166
rect 114648 32030 114860 32102
rect 114648 31966 114790 32030
rect 114854 31966 114860 32030
rect 114648 31960 114860 31966
rect 115056 32166 115404 32172
rect 115056 32102 115198 32166
rect 115262 32102 115334 32166
rect 115398 32102 115404 32166
rect 115056 32096 115404 32102
rect 115056 32036 115268 32096
rect 115464 32036 115676 32172
rect 115056 31960 115676 32036
rect 115872 32166 116084 32172
rect 115872 32102 115878 32166
rect 115942 32102 116084 32166
rect 115872 31960 116084 32102
rect 115464 31900 115540 31960
rect 109344 31830 109486 31894
rect 109550 31830 109556 31894
rect 109344 31824 109556 31830
rect 115192 31824 115540 31900
rect 115872 31900 115948 31960
rect 27472 31764 27548 31824
rect 109344 31764 109420 31824
rect 115192 31764 115268 31824
rect 20808 31694 20950 31758
rect 21014 31694 21020 31758
rect 20808 31688 21020 31694
rect 21216 31758 21972 31764
rect 21216 31694 21222 31758
rect 21286 31694 21630 31758
rect 21694 31694 21972 31758
rect 21216 31688 21972 31694
rect 21216 31628 21428 31688
rect 21216 31552 21564 31628
rect 21624 31552 21972 31688
rect 22032 31758 22244 31764
rect 22032 31694 22038 31758
rect 22102 31694 22244 31758
rect 22032 31622 22244 31694
rect 22032 31558 22174 31622
rect 22238 31558 22244 31622
rect 22032 31552 22244 31558
rect 22440 31758 22652 31764
rect 22440 31694 22582 31758
rect 22646 31694 22652 31758
rect 22440 31622 22652 31694
rect 22440 31558 22446 31622
rect 22510 31558 22652 31622
rect 22440 31552 22652 31558
rect 21216 31492 21292 31552
rect 21488 31492 21564 31552
rect 20808 31486 21020 31492
rect 20808 31422 20950 31486
rect 21014 31422 21020 31486
rect 14608 31239 14674 31242
rect 15022 31239 15088 31242
rect 14608 31237 15088 31239
rect 13600 31166 13812 31220
rect 14608 31181 14613 31237
rect 14669 31181 15027 31237
rect 15083 31181 15088 31237
rect 14608 31179 15088 31181
rect 14608 31176 14674 31179
rect 15022 31176 15088 31179
rect 13600 31110 13668 31166
rect 13724 31110 13812 31166
rect 13600 31084 13812 31110
rect 0 31008 13812 31084
rect 20808 31144 21020 31422
rect 21216 31144 21428 31492
rect 21488 31416 21972 31492
rect 21624 31214 21972 31416
rect 21624 31150 21766 31214
rect 21830 31150 21972 31214
rect 21624 31144 21972 31150
rect 22032 31350 22244 31356
rect 22032 31286 22174 31350
rect 22238 31286 22244 31350
rect 22032 31144 22244 31286
rect 22440 31350 22652 31356
rect 22440 31286 22446 31350
rect 22510 31286 22652 31350
rect 22440 31144 22652 31286
rect 27336 31280 27684 31764
rect 109344 31622 109556 31764
rect 109344 31558 109350 31622
rect 109414 31558 109486 31622
rect 109550 31558 109556 31622
rect 109344 31280 109556 31558
rect 114240 31758 114452 31764
rect 114240 31694 114382 31758
rect 114446 31694 114452 31758
rect 114240 31622 114452 31694
rect 114240 31558 114246 31622
rect 114310 31558 114452 31622
rect 114240 31552 114452 31558
rect 114648 31758 114860 31764
rect 114648 31694 114790 31758
rect 114854 31694 114860 31758
rect 114648 31622 114860 31694
rect 114648 31558 114654 31622
rect 114718 31558 114860 31622
rect 114648 31552 114860 31558
rect 115056 31688 115676 31764
rect 115872 31758 116084 31900
rect 115872 31694 115878 31758
rect 115942 31694 116084 31758
rect 115872 31688 116084 31694
rect 115056 31628 115268 31688
rect 115056 31552 115404 31628
rect 115464 31552 115676 31688
rect 115192 31492 115268 31552
rect 114240 31350 114452 31356
rect 114240 31286 114246 31350
rect 114310 31286 114452 31350
rect 27608 31220 27684 31280
rect 20808 31084 20884 31144
rect 22032 31084 22108 31144
rect 22440 31084 22516 31144
rect 20808 30942 21020 31084
rect 20808 30878 20814 30942
rect 20878 30878 21020 30942
rect 20808 30872 21020 30878
rect 21216 30736 21428 30948
rect 21624 30942 21972 30948
rect 21624 30878 21766 30942
rect 21830 30878 21972 30942
rect 21624 30812 21972 30878
rect 21488 30736 21972 30812
rect 22032 30736 22244 31084
rect 22440 30736 22652 31084
rect 21216 30676 21292 30736
rect 21488 30676 21564 30736
rect 22168 30676 22244 30736
rect 22576 30676 22652 30736
rect 1768 30648 1980 30676
rect 1768 30592 1794 30648
rect 1850 30592 1980 30648
rect 1768 30540 1980 30592
rect 1224 30534 1980 30540
rect 1224 30470 1230 30534
rect 1294 30470 1980 30534
rect 1224 30464 1980 30470
rect 14008 30670 14220 30676
rect 14008 30606 14014 30670
rect 14078 30606 14220 30670
rect 14008 30534 14220 30606
rect 14008 30470 14014 30534
rect 14078 30470 14220 30534
rect 14008 30464 14220 30470
rect 20808 30670 21020 30676
rect 20808 30606 20814 30670
rect 20878 30606 21020 30670
rect 20808 30534 21020 30606
rect 20808 30470 20814 30534
rect 20878 30470 21020 30534
rect 20808 30464 21020 30470
rect 21216 30600 21564 30676
rect 21216 30540 21428 30600
rect 21624 30540 21972 30676
rect 21216 30534 21972 30540
rect 21216 30470 21358 30534
rect 21422 30470 21972 30534
rect 21216 30464 21972 30470
rect 21352 30404 21428 30464
rect 21352 30328 21700 30404
rect 22032 30328 22244 30676
rect 22440 30328 22652 30676
rect 27336 31078 27684 31220
rect 27336 31014 27342 31078
rect 27406 31014 27684 31078
rect 27336 30806 27684 31014
rect 27336 30742 27342 30806
rect 27406 30742 27684 30806
rect 27336 30670 27684 30742
rect 27336 30606 27478 30670
rect 27542 30606 27684 30670
rect 27336 30600 27684 30606
rect 109344 31214 109556 31220
rect 109344 31150 109350 31214
rect 109414 31150 109556 31214
rect 109344 30670 109556 31150
rect 114240 31144 114452 31286
rect 114648 31350 114860 31356
rect 114648 31286 114654 31350
rect 114718 31286 114860 31350
rect 114648 31144 114860 31286
rect 115056 31144 115268 31492
rect 115328 31492 115404 31552
rect 115328 31416 115676 31492
rect 115464 31214 115676 31416
rect 115464 31150 115470 31214
rect 115534 31150 115676 31214
rect 115464 31144 115676 31150
rect 115872 31486 116084 31492
rect 115872 31422 115878 31486
rect 115942 31422 116084 31486
rect 115872 31144 116084 31422
rect 114376 31084 114452 31144
rect 114784 31084 114860 31144
rect 109344 30606 109350 30670
rect 109414 30606 109556 30670
rect 109344 30600 109556 30606
rect 114240 30736 114452 31084
rect 114648 30736 114860 31084
rect 115872 31084 115948 31144
rect 115056 30812 115268 30948
rect 115464 30942 115676 30948
rect 115464 30878 115470 30942
rect 115534 30878 115676 30942
rect 115056 30736 115404 30812
rect 115464 30736 115676 30878
rect 115872 30942 116084 31084
rect 115872 30878 115878 30942
rect 115942 30878 116084 30942
rect 115872 30872 116084 30878
rect 114240 30676 114316 30736
rect 114648 30676 114724 30736
rect 115192 30676 115268 30736
rect 21624 30268 21700 30328
rect 22168 30268 22244 30328
rect 22576 30268 22652 30328
rect 20808 30262 21020 30268
rect 20808 30198 20814 30262
rect 20878 30198 21020 30262
rect 13600 30038 13812 30132
rect 20808 30126 21020 30198
rect 20808 30062 20950 30126
rect 21014 30062 21020 30126
rect 20808 30056 21020 30062
rect 21216 30262 21428 30268
rect 21216 30198 21358 30262
rect 21422 30198 21428 30262
rect 13600 29996 13668 30038
rect 0 29982 13668 29996
rect 13724 29982 13812 30038
rect 0 29920 13812 29982
rect 14608 29969 14674 29972
rect 14942 29969 15008 29972
rect 14608 29967 15008 29969
rect 14608 29911 14613 29967
rect 14669 29911 14947 29967
rect 15003 29911 15008 29967
rect 21216 29920 21428 30198
rect 14608 29909 15008 29911
rect 14608 29906 14674 29909
rect 14942 29906 15008 29909
rect 21352 29860 21428 29920
rect 20808 29854 21020 29860
rect 20808 29790 20950 29854
rect 21014 29790 21020 29854
rect 20808 29718 21020 29790
rect 20808 29654 20814 29718
rect 20878 29654 21020 29718
rect 20808 29648 21020 29654
rect 21216 29648 21428 29860
rect 21624 29920 21972 30268
rect 22032 30126 22244 30268
rect 22032 30062 22174 30126
rect 22238 30062 22244 30126
rect 22032 30056 22244 30062
rect 22440 30126 22652 30268
rect 22440 30062 22582 30126
rect 22646 30062 22652 30126
rect 22440 30056 22652 30062
rect 27336 30398 27684 30404
rect 27336 30334 27478 30398
rect 27542 30334 27684 30398
rect 27336 30056 27684 30334
rect 109344 30398 109556 30404
rect 109344 30334 109350 30398
rect 109414 30334 109556 30398
rect 109344 30262 109556 30334
rect 109344 30198 109350 30262
rect 109414 30198 109556 30262
rect 109344 30056 109556 30198
rect 114240 30328 114452 30676
rect 114648 30328 114860 30676
rect 115056 30464 115268 30676
rect 115328 30676 115404 30736
rect 115600 30676 115676 30736
rect 115328 30600 115676 30676
rect 115464 30534 115676 30600
rect 115464 30470 115470 30534
rect 115534 30470 115676 30534
rect 115464 30464 115676 30470
rect 115872 30670 116084 30676
rect 115872 30606 115878 30670
rect 115942 30606 116084 30670
rect 115872 30534 116084 30606
rect 115872 30470 116014 30534
rect 116078 30470 116084 30534
rect 115872 30464 116084 30470
rect 134776 30648 134988 30676
rect 134776 30592 134844 30648
rect 134900 30592 134988 30648
rect 134776 30540 134988 30592
rect 134776 30534 135396 30540
rect 134776 30470 135326 30534
rect 135390 30470 135396 30534
rect 134776 30464 135396 30470
rect 114240 30268 114316 30328
rect 114784 30268 114860 30328
rect 114240 30126 114452 30268
rect 114240 30062 114246 30126
rect 114310 30062 114452 30126
rect 114240 30056 114452 30062
rect 114648 30126 114860 30268
rect 114648 30062 114654 30126
rect 114718 30062 114860 30126
rect 114648 30056 114860 30062
rect 27472 29996 27548 30056
rect 109480 29996 109556 30056
rect 21624 29860 21700 29920
rect 21624 29724 21972 29860
rect 21526 29718 21972 29724
rect 21488 29654 21494 29718
rect 21558 29654 21766 29718
rect 21830 29654 21972 29718
rect 21526 29648 21972 29654
rect 22032 29854 22244 29860
rect 22032 29790 22174 29854
rect 22238 29790 22244 29854
rect 22032 29718 22244 29790
rect 22032 29654 22038 29718
rect 22102 29654 22244 29718
rect 22032 29648 22244 29654
rect 22440 29854 22652 29860
rect 22440 29790 22582 29854
rect 22646 29790 22652 29854
rect 22440 29718 22652 29790
rect 22440 29654 22446 29718
rect 22510 29654 22652 29718
rect 22440 29648 22652 29654
rect 27336 29784 27684 29996
rect 109344 29990 109556 29996
rect 109344 29926 109350 29990
rect 109414 29926 109556 29990
rect 109344 29784 109556 29926
rect 115056 29920 115268 30268
rect 115192 29860 115268 29920
rect 114240 29854 114452 29860
rect 114240 29790 114246 29854
rect 114310 29790 114452 29854
rect 27336 29724 27412 29784
rect 109344 29724 109420 29784
rect 21896 29588 21972 29648
rect 22440 29588 22516 29648
rect 21896 29512 22516 29588
rect 27336 29512 27684 29724
rect 109344 29512 109556 29724
rect 114240 29718 114452 29790
rect 114240 29654 114246 29718
rect 114310 29654 114452 29718
rect 114240 29648 114452 29654
rect 114648 29854 114860 29860
rect 114648 29790 114654 29854
rect 114718 29790 114860 29854
rect 114648 29718 114860 29790
rect 114648 29654 114654 29718
rect 114718 29654 114860 29718
rect 114648 29648 114860 29654
rect 115056 29724 115268 29860
rect 115464 30262 115676 30268
rect 115464 30198 115470 30262
rect 115534 30198 115676 30262
rect 115464 29920 115676 30198
rect 115872 30262 116084 30268
rect 115872 30198 116014 30262
rect 116078 30198 116084 30262
rect 115872 30126 116084 30198
rect 115872 30062 115878 30126
rect 115942 30062 116084 30126
rect 115872 30056 116084 30062
rect 115464 29860 115540 29920
rect 115056 29718 115404 29724
rect 115056 29654 115334 29718
rect 115398 29654 115404 29718
rect 115056 29648 115404 29654
rect 115464 29718 115676 29860
rect 115464 29654 115470 29718
rect 115534 29654 115676 29718
rect 115464 29648 115676 29654
rect 115872 29854 116084 29860
rect 115872 29790 115878 29854
rect 115942 29790 116084 29854
rect 115872 29718 116084 29790
rect 115872 29654 115878 29718
rect 115942 29654 116084 29718
rect 115872 29648 116084 29654
rect 27336 29452 27412 29512
rect 109480 29452 109556 29512
rect 20808 29446 21020 29452
rect 20808 29382 20814 29446
rect 20878 29382 21020 29446
rect 14008 29310 14220 29316
rect 14008 29246 14150 29310
rect 14214 29246 14220 29310
rect 14008 29180 14220 29246
rect 20808 29310 21020 29382
rect 20808 29246 20814 29310
rect 20878 29246 21020 29310
rect 20808 29240 21020 29246
rect 21216 29446 21564 29452
rect 21216 29382 21494 29446
rect 21558 29382 21564 29446
rect 21216 29376 21564 29382
rect 21624 29446 21972 29452
rect 21624 29382 21766 29446
rect 21830 29382 21972 29446
rect 21216 29240 21428 29376
rect 21624 29310 21972 29382
rect 21624 29246 21766 29310
rect 21830 29246 21972 29310
rect 21624 29240 21972 29246
rect 22032 29446 22244 29452
rect 22032 29382 22038 29446
rect 22102 29382 22244 29446
rect 22032 29310 22244 29382
rect 22032 29246 22174 29310
rect 22238 29246 22244 29310
rect 22032 29240 22244 29246
rect 22440 29446 22652 29452
rect 22440 29382 22446 29446
rect 22510 29382 22652 29446
rect 22440 29310 22652 29382
rect 22440 29246 22582 29310
rect 22646 29246 22652 29310
rect 22440 29240 22652 29246
rect 27336 29240 27684 29452
rect 109344 29240 109556 29452
rect 114240 29446 114452 29452
rect 114240 29382 114246 29446
rect 114310 29382 114452 29446
rect 114240 29310 114452 29382
rect 114240 29246 114246 29310
rect 114310 29246 114452 29310
rect 114240 29240 114452 29246
rect 114648 29446 114860 29452
rect 114648 29382 114654 29446
rect 114718 29382 114860 29446
rect 114648 29310 114860 29382
rect 114648 29246 114654 29310
rect 114718 29246 114860 29310
rect 114648 29240 114860 29246
rect 115056 29310 115268 29452
rect 115366 29446 115676 29452
rect 115328 29382 115334 29446
rect 115398 29382 115470 29446
rect 115534 29382 115676 29446
rect 115366 29376 115676 29382
rect 115464 29316 115676 29376
rect 115366 29310 115676 29316
rect 115056 29246 115062 29310
rect 115126 29246 115268 29310
rect 115328 29246 115334 29310
rect 115398 29246 115676 29310
rect 115056 29240 115268 29246
rect 115366 29240 115676 29246
rect 115872 29446 116084 29452
rect 115872 29382 115878 29446
rect 115942 29382 116084 29446
rect 115872 29310 116084 29382
rect 115872 29246 116014 29310
rect 116078 29246 116084 29310
rect 115872 29240 116084 29246
rect 27472 29180 27548 29240
rect 109480 29180 109556 29240
rect 14008 29174 17892 29180
rect 14008 29110 17822 29174
rect 17886 29110 17892 29174
rect 14008 29104 17892 29110
rect 1224 29038 1980 29044
rect 1224 28974 1230 29038
rect 1294 28974 1980 29038
rect 1224 28968 1980 28974
rect 1768 28912 1794 28968
rect 1850 28912 1980 28968
rect 1768 28832 1980 28912
rect 20808 29038 21020 29044
rect 20808 28974 20814 29038
rect 20878 28974 21020 29038
rect 20808 28902 21020 28974
rect 20808 28838 20950 28902
rect 21014 28838 21020 28902
rect 20808 28832 21020 28838
rect 21216 28902 21428 29044
rect 21216 28838 21222 28902
rect 21286 28838 21428 28902
rect 21216 28832 21428 28838
rect 21624 29038 21972 29044
rect 21624 28974 21766 29038
rect 21830 28974 21972 29038
rect 21624 28902 21972 28974
rect 21624 28838 21630 28902
rect 21694 28838 21972 28902
rect 21624 28832 21972 28838
rect 22032 29038 22244 29044
rect 22032 28974 22174 29038
rect 22238 28974 22244 29038
rect 22032 28902 22244 28974
rect 22032 28838 22038 28902
rect 22102 28838 22244 28902
rect 22032 28832 22244 28838
rect 22440 29038 22652 29044
rect 22440 28974 22582 29038
rect 22646 28974 22652 29038
rect 22440 28902 22652 28974
rect 27336 28968 27684 29180
rect 109344 28968 109556 29180
rect 27608 28908 27684 28968
rect 109480 28908 109556 28968
rect 22440 28838 22582 28902
rect 22646 28838 22652 28902
rect 22440 28832 22652 28838
rect 27336 28696 27684 28908
rect 109344 28696 109556 28908
rect 114240 29038 114452 29044
rect 114240 28974 114246 29038
rect 114310 28974 114452 29038
rect 114240 28902 114452 28974
rect 114240 28838 114382 28902
rect 114446 28838 114452 28902
rect 114240 28832 114452 28838
rect 114648 29038 114860 29044
rect 114648 28974 114654 29038
rect 114718 28974 114860 29038
rect 114648 28902 114860 28974
rect 114648 28838 114790 28902
rect 114854 28838 114860 28902
rect 114648 28832 114860 28838
rect 115056 29038 115404 29044
rect 115056 28974 115062 29038
rect 115126 28974 115334 29038
rect 115398 28974 115404 29038
rect 115056 28968 115404 28974
rect 115056 28902 115268 28968
rect 115056 28838 115198 28902
rect 115262 28838 115268 28902
rect 115056 28832 115268 28838
rect 115464 28832 115676 29044
rect 115872 29038 116084 29044
rect 115872 28974 116014 29038
rect 116078 28974 116084 29038
rect 115872 28902 116084 28974
rect 115872 28838 115878 28902
rect 115942 28838 116084 28902
rect 115872 28832 116084 28838
rect 134776 29038 135396 29044
rect 134776 28974 135326 29038
rect 135390 28974 135396 29038
rect 134776 28968 135396 28974
rect 134776 28912 134844 28968
rect 134900 28912 134988 28968
rect 134776 28832 134988 28912
rect 115464 28772 115540 28832
rect 115192 28696 115540 28772
rect 27472 28636 27548 28696
rect 109344 28636 109420 28696
rect 115192 28636 115268 28696
rect 20808 28630 21020 28636
rect 20808 28566 20950 28630
rect 21014 28566 21020 28630
rect 20808 28494 21020 28566
rect 20808 28430 20950 28494
rect 21014 28430 21020 28494
rect 20808 28424 21020 28430
rect 21216 28630 21428 28636
rect 21216 28566 21222 28630
rect 21286 28566 21428 28630
rect 21216 28494 21428 28566
rect 21624 28630 21972 28636
rect 21624 28566 21630 28630
rect 21694 28566 21972 28630
rect 21624 28500 21972 28566
rect 21526 28494 21972 28500
rect 21216 28430 21358 28494
rect 21422 28430 21428 28494
rect 21488 28430 21494 28494
rect 21558 28430 21972 28494
rect 21216 28424 21428 28430
rect 21526 28424 21972 28430
rect 22032 28630 22244 28636
rect 22032 28566 22038 28630
rect 22102 28566 22244 28630
rect 22032 28494 22244 28566
rect 22032 28430 22174 28494
rect 22238 28430 22244 28494
rect 22032 28424 22244 28430
rect 22440 28630 22652 28636
rect 22440 28566 22582 28630
rect 22646 28566 22652 28630
rect 22440 28494 22652 28566
rect 22440 28430 22446 28494
rect 22510 28430 22652 28494
rect 22440 28424 22652 28430
rect 27336 28424 27684 28636
rect 109344 28424 109556 28636
rect 114240 28630 114452 28636
rect 114240 28566 114382 28630
rect 114446 28566 114452 28630
rect 114240 28494 114452 28566
rect 114240 28430 114382 28494
rect 114446 28430 114452 28494
rect 114240 28424 114452 28430
rect 114648 28630 114860 28636
rect 114648 28566 114790 28630
rect 114854 28566 114860 28630
rect 114648 28494 114860 28566
rect 114648 28430 114790 28494
rect 114854 28430 114860 28494
rect 114648 28424 114860 28430
rect 115056 28630 115676 28636
rect 115056 28566 115198 28630
rect 115262 28566 115676 28630
rect 115056 28560 115676 28566
rect 115056 28424 115268 28560
rect 115464 28494 115676 28560
rect 115464 28430 115606 28494
rect 115670 28430 115676 28494
rect 115464 28424 115676 28430
rect 115872 28630 116084 28636
rect 115872 28566 115878 28630
rect 115942 28566 116084 28630
rect 115872 28494 116084 28566
rect 115872 28430 115878 28494
rect 115942 28430 116084 28494
rect 115872 28424 116084 28430
rect 14608 28411 14674 28414
rect 14862 28411 14928 28414
rect 14608 28409 14928 28411
rect 13600 28338 13812 28364
rect 14608 28353 14613 28409
rect 14669 28353 14867 28409
rect 14923 28353 14928 28409
rect 27608 28364 27684 28424
rect 109480 28364 109556 28424
rect 14608 28351 14928 28353
rect 14608 28348 14674 28351
rect 14862 28348 14928 28351
rect 13600 28282 13668 28338
rect 13724 28282 13812 28338
rect 13600 28228 13812 28282
rect 0 28152 13812 28228
rect 20808 28222 21020 28228
rect 20808 28158 20950 28222
rect 21014 28158 21020 28222
rect 20808 28092 21020 28158
rect 14694 28087 14778 28091
rect 14694 28082 14811 28087
rect 18942 28086 21020 28092
rect 14694 28026 14750 28082
rect 14806 28026 14811 28082
rect 14694 28021 14811 28026
rect 18904 28022 18910 28086
rect 18974 28022 21020 28086
rect 14694 28017 14778 28021
rect 18942 28016 21020 28022
rect 21216 28222 21564 28228
rect 21216 28158 21358 28222
rect 21422 28158 21494 28222
rect 21558 28158 21564 28222
rect 21216 28152 21564 28158
rect 21216 28092 21428 28152
rect 21624 28092 21972 28228
rect 21216 28086 21972 28092
rect 21216 28022 21766 28086
rect 21830 28022 21972 28086
rect 21216 28016 21972 28022
rect 22032 28222 22244 28228
rect 22032 28158 22174 28222
rect 22238 28158 22244 28222
rect 22032 28086 22244 28158
rect 22032 28022 22038 28086
rect 22102 28022 22244 28086
rect 22032 28016 22244 28022
rect 22440 28222 22652 28228
rect 22440 28158 22446 28222
rect 22510 28158 22652 28222
rect 22440 28086 22652 28158
rect 27336 28152 27684 28364
rect 109344 28152 109556 28364
rect 27472 28092 27548 28152
rect 109480 28092 109556 28152
rect 22440 28022 22446 28086
rect 22510 28022 22652 28086
rect 22440 28016 22652 28022
rect 20808 27956 20884 28016
rect 14008 27814 14220 27820
rect 14008 27750 14014 27814
rect 14078 27750 14220 27814
rect 14008 27684 14220 27750
rect 14008 27678 15988 27684
rect 14008 27614 15918 27678
rect 15982 27614 15988 27678
rect 14008 27608 15988 27614
rect 20808 27608 21020 27956
rect 27336 27880 27684 28092
rect 109344 27880 109556 28092
rect 114240 28222 114452 28228
rect 114240 28158 114382 28222
rect 114446 28158 114452 28222
rect 114240 28086 114452 28158
rect 114240 28022 114382 28086
rect 114446 28022 114452 28086
rect 114240 28016 114452 28022
rect 114648 28222 114860 28228
rect 114648 28158 114790 28222
rect 114854 28158 114860 28222
rect 114648 28086 114860 28158
rect 114648 28022 114790 28086
rect 114854 28022 114860 28086
rect 114648 28016 114860 28022
rect 115056 28086 115268 28228
rect 115056 28022 115198 28086
rect 115262 28022 115268 28086
rect 115056 28016 115268 28022
rect 115464 28222 115676 28228
rect 115464 28158 115606 28222
rect 115670 28158 115676 28222
rect 115464 28016 115676 28158
rect 115872 28222 116084 28228
rect 115872 28158 115878 28222
rect 115942 28158 116084 28222
rect 115872 28016 116084 28158
rect 115464 27956 115540 28016
rect 116008 27956 116084 28016
rect 27472 27820 27548 27880
rect 109480 27820 109556 27880
rect 115192 27880 115540 27956
rect 115192 27820 115268 27880
rect 20944 27548 21020 27608
rect 1768 27288 1980 27412
rect 1768 27276 1794 27288
rect 1224 27270 1794 27276
rect 1224 27206 1230 27270
rect 1294 27232 1794 27270
rect 1850 27232 1980 27288
rect 1294 27206 1980 27232
rect 1224 27200 1980 27206
rect 17408 27270 17620 27548
rect 17408 27206 17414 27270
rect 17478 27206 17620 27270
rect 17408 27200 17620 27206
rect 17816 27542 18436 27548
rect 17816 27478 17822 27542
rect 17886 27478 18436 27542
rect 17816 27472 18436 27478
rect 17816 27200 18028 27472
rect 18224 27270 18436 27472
rect 18224 27206 18366 27270
rect 18430 27206 18436 27270
rect 18224 27200 18436 27206
rect 18632 27406 18980 27412
rect 18632 27342 18910 27406
rect 18974 27342 18980 27406
rect 18632 27336 18980 27342
rect 18632 27270 18844 27336
rect 18632 27206 18638 27270
rect 18702 27206 18844 27270
rect 18632 27200 18844 27206
rect 19040 27276 19252 27412
rect 19040 27270 20748 27276
rect 19040 27206 19046 27270
rect 19110 27206 20678 27270
rect 20742 27206 20748 27270
rect 19040 27200 20748 27206
rect 20808 27200 21020 27548
rect 21216 27608 21428 27820
rect 21624 27814 21972 27820
rect 21624 27750 21766 27814
rect 21830 27750 21972 27814
rect 21624 27608 21972 27750
rect 22032 27814 22244 27820
rect 22032 27750 22038 27814
rect 22102 27750 22244 27814
rect 22032 27678 22244 27750
rect 22032 27614 22038 27678
rect 22102 27614 22244 27678
rect 22032 27608 22244 27614
rect 22440 27814 22652 27820
rect 22440 27750 22446 27814
rect 22510 27750 22652 27814
rect 22440 27678 22652 27750
rect 22440 27614 22582 27678
rect 22646 27614 22652 27678
rect 22440 27608 22652 27614
rect 21216 27548 21292 27608
rect 21624 27548 21700 27608
rect 21216 27270 21428 27548
rect 21624 27276 21972 27548
rect 21526 27270 21972 27276
rect 21216 27206 21358 27270
rect 21422 27206 21428 27270
rect 21488 27206 21494 27270
rect 21558 27206 21972 27270
rect 21216 27200 21428 27206
rect 21526 27200 21972 27206
rect 22032 27406 22244 27412
rect 22032 27342 22038 27406
rect 22102 27342 22244 27406
rect 22032 27200 22244 27342
rect 20808 27140 20884 27200
rect 22168 27140 22244 27200
rect 20808 26998 21020 27140
rect 20808 26934 20814 26998
rect 20878 26934 21020 26998
rect 20808 26928 21020 26934
rect 21216 26998 21564 27004
rect 21216 26934 21358 26998
rect 21422 26934 21494 26998
rect 21558 26934 21564 26998
rect 21216 26928 21564 26934
rect 21216 26868 21428 26928
rect 18496 26792 19116 26868
rect 20710 26862 21428 26868
rect 20672 26798 20678 26862
rect 20742 26798 21428 26862
rect 20710 26792 21428 26798
rect 21624 26792 21972 27004
rect 22032 26792 22244 27140
rect 22440 27406 22652 27412
rect 22440 27342 22582 27406
rect 22646 27342 22652 27406
rect 22440 27200 22652 27342
rect 27336 27336 27684 27820
rect 109344 27336 109556 27820
rect 114240 27814 114452 27820
rect 114240 27750 114382 27814
rect 114446 27750 114452 27814
rect 114240 27678 114452 27750
rect 114240 27614 114382 27678
rect 114446 27614 114452 27678
rect 114240 27608 114452 27614
rect 114648 27814 114860 27820
rect 114648 27750 114790 27814
rect 114854 27750 114860 27814
rect 114648 27678 114860 27750
rect 114648 27614 114790 27678
rect 114854 27614 114860 27678
rect 114648 27608 114860 27614
rect 115056 27814 115676 27820
rect 115056 27750 115198 27814
rect 115262 27750 115676 27814
rect 115056 27744 115676 27750
rect 115056 27684 115268 27744
rect 115056 27608 115404 27684
rect 115464 27608 115676 27744
rect 115872 27608 116084 27956
rect 115192 27548 115268 27608
rect 27472 27276 27548 27336
rect 109480 27276 109556 27336
rect 22440 27140 22516 27200
rect 22440 26792 22652 27140
rect 18496 26732 18572 26792
rect 19040 26732 19116 26792
rect 21216 26732 21292 26792
rect 21760 26732 21836 26792
rect 22168 26732 22244 26792
rect 22576 26732 22652 26792
rect 17408 26726 17620 26732
rect 17408 26662 17414 26726
rect 17478 26662 17620 26726
rect 17408 26596 17620 26662
rect 17816 26596 18028 26732
rect 18224 26726 18572 26732
rect 18224 26662 18366 26726
rect 18430 26662 18572 26726
rect 18224 26656 18572 26662
rect 18632 26726 18844 26732
rect 18632 26662 18638 26726
rect 18702 26662 18844 26726
rect 18224 26596 18436 26656
rect 17408 26590 17756 26596
rect 17408 26526 17550 26590
rect 17614 26526 17686 26590
rect 17750 26526 17756 26590
rect 17408 26520 17756 26526
rect 17816 26520 18436 26596
rect 17952 26460 18028 26520
rect 17952 26454 18300 26460
rect 17952 26390 18230 26454
rect 18294 26390 18300 26454
rect 17952 26384 18300 26390
rect 18632 26454 18844 26662
rect 18632 26390 18638 26454
rect 18702 26390 18844 26454
rect 18632 26384 18844 26390
rect 19040 26726 19252 26732
rect 19040 26662 19046 26726
rect 19110 26662 19252 26726
rect 19040 26384 19252 26662
rect 20808 26726 21020 26732
rect 20808 26662 20814 26726
rect 20878 26662 21020 26726
rect 20808 26590 21020 26662
rect 20808 26526 20814 26590
rect 20878 26526 21020 26590
rect 20808 26520 21020 26526
rect 21216 26590 21428 26732
rect 21216 26526 21222 26590
rect 21286 26526 21428 26590
rect 21216 26520 21428 26526
rect 21624 26590 21972 26732
rect 21624 26526 21902 26590
rect 21966 26526 21972 26590
rect 21624 26520 21972 26526
rect 22032 26384 22244 26732
rect 22440 26384 22652 26732
rect 27336 26726 27684 27276
rect 27336 26662 27342 26726
rect 27406 26662 27684 26726
rect 27336 26656 27684 26662
rect 109344 26726 109556 27276
rect 114240 27406 114452 27412
rect 114240 27342 114382 27406
rect 114446 27342 114452 27406
rect 114240 27200 114452 27342
rect 114648 27406 114860 27412
rect 114648 27342 114790 27406
rect 114854 27342 114860 27406
rect 114648 27200 114860 27342
rect 115056 27200 115268 27548
rect 115328 27548 115404 27608
rect 115872 27548 115948 27608
rect 115328 27472 115676 27548
rect 115464 27276 115676 27472
rect 115464 27270 115812 27276
rect 115464 27206 115606 27270
rect 115670 27206 115742 27270
rect 115806 27206 115812 27270
rect 115464 27200 115812 27206
rect 115872 27200 116084 27548
rect 117912 27472 118668 27548
rect 117912 27412 117988 27472
rect 117640 27336 117988 27412
rect 117640 27270 117852 27336
rect 117640 27206 117646 27270
rect 117710 27206 117782 27270
rect 117846 27206 117852 27270
rect 117640 27200 117852 27206
rect 118048 27270 118260 27412
rect 118048 27206 118190 27270
rect 118254 27206 118260 27270
rect 118048 27200 118260 27206
rect 118456 27276 118668 27472
rect 118864 27276 119076 27548
rect 118456 27270 119076 27276
rect 118456 27206 118870 27270
rect 118934 27206 119076 27270
rect 118456 27200 119076 27206
rect 119272 27270 119484 27548
rect 119272 27206 119278 27270
rect 119342 27206 119484 27270
rect 119272 27200 119484 27206
rect 134776 27288 134988 27412
rect 134776 27232 134844 27288
rect 134900 27276 134988 27288
rect 134900 27270 135396 27276
rect 134900 27232 135326 27270
rect 134776 27206 135326 27232
rect 135390 27206 135396 27270
rect 134776 27200 135396 27206
rect 114240 27140 114316 27200
rect 114648 27140 114724 27200
rect 116008 27140 116084 27200
rect 114240 26792 114452 27140
rect 114648 26792 114860 27140
rect 115056 26792 115268 27004
rect 115464 26998 115676 27004
rect 115464 26934 115606 26998
rect 115670 26934 115676 26998
rect 115464 26868 115676 26934
rect 115872 26998 116084 27140
rect 115872 26934 115878 26998
rect 115942 26934 116084 26998
rect 115872 26928 116084 26934
rect 114376 26732 114452 26792
rect 114784 26732 114860 26792
rect 115192 26732 115268 26792
rect 115328 26792 115676 26868
rect 115774 26862 117716 26868
rect 115736 26798 115742 26862
rect 115806 26798 117646 26862
rect 117710 26798 117716 26862
rect 115774 26792 117716 26798
rect 115328 26732 115404 26792
rect 109344 26662 109350 26726
rect 109414 26662 109556 26726
rect 109344 26656 109556 26662
rect 27336 26454 27684 26460
rect 27336 26390 27342 26454
rect 27406 26390 27684 26454
rect 18632 26324 18708 26384
rect 22032 26324 22108 26384
rect 22440 26324 22516 26384
rect 17718 26318 18708 26324
rect 17680 26254 17686 26318
rect 17750 26254 18708 26318
rect 17718 26248 18708 26254
rect 20808 26318 21020 26324
rect 20808 26254 20814 26318
rect 20878 26254 21020 26318
rect 20808 26182 21020 26254
rect 20808 26118 20814 26182
rect 20878 26118 21020 26182
rect 20808 26112 21020 26118
rect 21216 26318 21428 26324
rect 21216 26254 21222 26318
rect 21286 26254 21428 26318
rect 3128 25976 4156 26052
rect 3128 25840 3340 25976
rect 3944 25916 4156 25976
rect 18496 25976 19116 26052
rect 21216 25976 21428 26254
rect 21624 26318 21972 26324
rect 21624 26254 21902 26318
rect 21966 26254 21972 26318
rect 21624 26052 21972 26254
rect 22032 26182 22244 26324
rect 22032 26118 22174 26182
rect 22238 26118 22244 26182
rect 22032 26112 22244 26118
rect 22440 26182 22652 26324
rect 22440 26118 22582 26182
rect 22646 26118 22652 26182
rect 22440 26112 22652 26118
rect 27336 26318 27684 26390
rect 27336 26254 27478 26318
rect 27542 26254 27684 26318
rect 27336 26112 27684 26254
rect 109344 26454 109556 26460
rect 109344 26390 109350 26454
rect 109414 26390 109556 26454
rect 109344 26318 109556 26390
rect 114240 26384 114452 26732
rect 114376 26324 114452 26384
rect 109344 26254 109350 26318
rect 109414 26254 109556 26318
rect 109344 26112 109556 26254
rect 114240 26182 114452 26324
rect 114240 26118 114246 26182
rect 114310 26118 114452 26182
rect 114240 26112 114452 26118
rect 114648 26384 114860 26732
rect 115056 26656 115404 26732
rect 115464 26732 115540 26792
rect 115056 26520 115268 26656
rect 115464 26590 115676 26732
rect 115464 26526 115470 26590
rect 115534 26526 115676 26590
rect 115464 26520 115676 26526
rect 115872 26726 116084 26732
rect 115872 26662 115878 26726
rect 115942 26662 116084 26726
rect 115872 26590 116084 26662
rect 115872 26526 115878 26590
rect 115942 26526 116084 26590
rect 115872 26520 116084 26526
rect 117640 26726 117852 26732
rect 117640 26662 117782 26726
rect 117846 26662 117852 26726
rect 117640 26454 117852 26662
rect 117640 26390 117646 26454
rect 117710 26390 117852 26454
rect 117640 26384 117852 26390
rect 118048 26726 118260 26732
rect 118048 26662 118190 26726
rect 118254 26662 118260 26726
rect 118048 26454 118260 26662
rect 118456 26726 118804 26732
rect 118456 26662 118734 26726
rect 118798 26662 118804 26726
rect 118456 26656 118804 26662
rect 118456 26596 118668 26656
rect 118864 26596 119076 26732
rect 118456 26590 119076 26596
rect 118456 26526 119006 26590
rect 119070 26526 119076 26590
rect 118456 26520 119076 26526
rect 119272 26726 119484 26732
rect 119272 26662 119278 26726
rect 119342 26662 119484 26726
rect 119272 26590 119484 26662
rect 119272 26526 119278 26590
rect 119342 26526 119484 26590
rect 119272 26520 119484 26526
rect 118048 26390 118190 26454
rect 118254 26390 118260 26454
rect 118048 26384 118260 26390
rect 114648 26324 114724 26384
rect 114648 26182 114860 26324
rect 114648 26118 114654 26182
rect 114718 26118 114860 26182
rect 114648 26112 114860 26118
rect 27472 26052 27548 26112
rect 109480 26052 109556 26112
rect 18496 25916 18572 25976
rect 19040 25916 19116 25976
rect 21352 25916 21428 25976
rect 21488 25976 21972 26052
rect 27336 26046 27684 26052
rect 27336 25982 27478 26046
rect 27542 25982 27684 26046
rect 21488 25916 21564 25976
rect 3846 25910 4156 25916
rect 3808 25846 3814 25910
rect 3878 25846 4156 25910
rect 3846 25840 4156 25846
rect 17408 25910 17620 25916
rect 17408 25846 17550 25910
rect 17614 25846 17620 25910
rect 17408 25774 17620 25846
rect 17408 25710 17414 25774
rect 17478 25710 17620 25774
rect 17408 25704 17620 25710
rect 17816 25780 18028 25916
rect 18224 25910 18572 25916
rect 18224 25846 18230 25910
rect 18294 25846 18572 25910
rect 18224 25840 18572 25846
rect 18632 25910 18844 25916
rect 18632 25846 18638 25910
rect 18702 25846 18844 25910
rect 18224 25780 18436 25840
rect 17816 25774 18436 25780
rect 17816 25710 18230 25774
rect 18294 25710 18436 25774
rect 17816 25704 18436 25710
rect 18632 25774 18844 25846
rect 18632 25710 18774 25774
rect 18838 25710 18844 25774
rect 18632 25704 18844 25710
rect 19040 25774 19252 25916
rect 19040 25710 19182 25774
rect 19246 25710 19252 25774
rect 19040 25704 19252 25710
rect 20808 25910 21020 25916
rect 20808 25846 20814 25910
rect 20878 25846 21020 25910
rect 20808 25774 21020 25846
rect 20808 25710 20814 25774
rect 20878 25710 21020 25774
rect 20808 25704 21020 25710
rect 21216 25840 21564 25916
rect 21216 25780 21428 25840
rect 21624 25780 21972 25916
rect 21216 25704 21972 25780
rect 22032 25910 22244 25916
rect 22032 25846 22174 25910
rect 22238 25846 22244 25910
rect 22032 25774 22244 25846
rect 22032 25710 22174 25774
rect 22238 25710 22244 25774
rect 22032 25704 22244 25710
rect 22440 25910 22652 25916
rect 22440 25846 22582 25910
rect 22646 25846 22652 25910
rect 22440 25774 22652 25846
rect 27336 25840 27684 25982
rect 109344 26046 109556 26052
rect 109344 25982 109350 26046
rect 109414 25982 109556 26046
rect 109344 25840 109556 25982
rect 115056 25976 115268 26324
rect 115464 26318 115676 26324
rect 115464 26254 115470 26318
rect 115534 26254 115676 26318
rect 115464 25976 115676 26254
rect 115872 26318 116084 26324
rect 115872 26254 115878 26318
rect 115942 26254 116084 26318
rect 115872 26182 116084 26254
rect 115872 26118 116014 26182
rect 116078 26118 116084 26182
rect 115872 26112 116084 26118
rect 115056 25916 115132 25976
rect 115600 25916 115676 25976
rect 118320 25976 119348 26052
rect 118320 25916 118396 25976
rect 119272 25916 119348 25976
rect 27608 25780 27684 25840
rect 109480 25780 109556 25840
rect 22440 25710 22582 25774
rect 22646 25710 22652 25774
rect 22440 25704 22652 25710
rect 21624 25644 21700 25704
rect 1224 25638 1980 25644
rect 1224 25574 1230 25638
rect 1294 25608 1980 25638
rect 1294 25574 1794 25608
rect 1224 25568 1794 25574
rect 1768 25552 1794 25568
rect 1850 25552 1980 25608
rect 1768 25432 1980 25552
rect 21488 25568 21700 25644
rect 21488 25508 21564 25568
rect 20808 25502 21020 25508
rect 20808 25438 20814 25502
rect 20878 25438 21020 25502
rect 20808 25366 21020 25438
rect 2536 25365 2602 25366
rect 2494 25301 2537 25365
rect 2601 25301 2644 25365
rect 20808 25302 20814 25366
rect 20878 25302 21020 25366
rect 2536 25300 2602 25301
rect 20808 25296 21020 25302
rect 21216 25432 21564 25508
rect 21216 25366 21428 25432
rect 21624 25372 21972 25508
rect 21526 25366 21972 25372
rect 21216 25302 21358 25366
rect 21422 25302 21428 25366
rect 21488 25302 21494 25366
rect 21558 25302 21766 25366
rect 21830 25302 21972 25366
rect 21216 25296 21428 25302
rect 21526 25296 21972 25302
rect 22032 25502 22244 25508
rect 22032 25438 22174 25502
rect 22238 25438 22244 25502
rect 22032 25366 22244 25438
rect 22032 25302 22174 25366
rect 22238 25302 22244 25366
rect 22032 25296 22244 25302
rect 22440 25502 22652 25508
rect 22440 25438 22582 25502
rect 22646 25438 22652 25502
rect 22440 25366 22652 25438
rect 22440 25302 22446 25366
rect 22510 25302 22652 25366
rect 22440 25296 22652 25302
rect 27336 25296 27684 25780
rect 109344 25296 109556 25780
rect 114240 25910 114452 25916
rect 114240 25846 114246 25910
rect 114310 25846 114452 25910
rect 114240 25774 114452 25846
rect 114240 25710 114246 25774
rect 114310 25710 114452 25774
rect 114240 25704 114452 25710
rect 114648 25910 114860 25916
rect 114648 25846 114654 25910
rect 114718 25846 114860 25910
rect 114648 25774 114860 25846
rect 114648 25710 114790 25774
rect 114854 25710 114860 25774
rect 114648 25704 114860 25710
rect 115056 25774 115268 25916
rect 115056 25710 115062 25774
rect 115126 25710 115268 25774
rect 115056 25704 115268 25710
rect 115464 25774 115676 25916
rect 115464 25710 115606 25774
rect 115670 25710 115676 25774
rect 115464 25704 115676 25710
rect 115872 25910 116084 25916
rect 115872 25846 116014 25910
rect 116078 25846 116084 25910
rect 115872 25774 116084 25846
rect 115872 25710 116014 25774
rect 116078 25710 116084 25774
rect 115872 25704 116084 25710
rect 117640 25910 117852 25916
rect 117640 25846 117646 25910
rect 117710 25846 117852 25910
rect 117640 25774 117852 25846
rect 117640 25710 117646 25774
rect 117710 25710 117852 25774
rect 117640 25704 117852 25710
rect 118048 25910 118396 25916
rect 118048 25846 118190 25910
rect 118254 25846 118396 25910
rect 118048 25840 118396 25846
rect 118048 25774 118260 25840
rect 118048 25710 118190 25774
rect 118254 25710 118260 25774
rect 118048 25704 118260 25710
rect 118456 25780 118668 25916
rect 118864 25910 119076 25916
rect 118864 25846 119006 25910
rect 119070 25846 119076 25910
rect 118864 25780 119076 25846
rect 118456 25774 119076 25780
rect 118456 25710 119006 25774
rect 119070 25710 119076 25774
rect 118456 25704 119076 25710
rect 119272 25910 119484 25916
rect 119272 25846 119278 25910
rect 119342 25846 119484 25910
rect 119272 25780 119484 25846
rect 119272 25774 120844 25780
rect 119272 25710 119414 25774
rect 119478 25710 120774 25774
rect 120838 25710 120844 25774
rect 119272 25704 120844 25710
rect 134776 25608 134988 25644
rect 134776 25552 134844 25608
rect 134900 25552 134988 25608
rect 134776 25508 134988 25552
rect 114240 25502 114452 25508
rect 114240 25438 114246 25502
rect 114310 25438 114452 25502
rect 114240 25366 114452 25438
rect 114240 25302 114246 25366
rect 114310 25302 114452 25366
rect 114240 25296 114452 25302
rect 114648 25502 114860 25508
rect 114648 25438 114790 25502
rect 114854 25438 114860 25502
rect 114648 25366 114860 25438
rect 114648 25302 114654 25366
rect 114718 25302 114860 25366
rect 114648 25296 114860 25302
rect 115056 25502 115268 25508
rect 115056 25438 115062 25502
rect 115126 25438 115268 25502
rect 115056 25372 115268 25438
rect 115464 25502 115676 25508
rect 115464 25438 115606 25502
rect 115670 25438 115676 25502
rect 115464 25372 115676 25438
rect 115056 25366 115676 25372
rect 115056 25302 115198 25366
rect 115262 25302 115470 25366
rect 115534 25302 115676 25366
rect 115056 25296 115676 25302
rect 115872 25502 116084 25508
rect 115872 25438 116014 25502
rect 116078 25438 116084 25502
rect 115872 25366 116084 25438
rect 134776 25502 135396 25508
rect 134776 25438 135326 25502
rect 135390 25438 135396 25502
rect 134776 25432 135396 25438
rect 115872 25302 115878 25366
rect 115942 25302 116084 25366
rect 115872 25296 116084 25302
rect 27336 25236 27412 25296
rect 109344 25236 109420 25296
rect 17272 25160 17892 25236
rect 17272 25100 17348 25160
rect 17816 25100 17892 25160
rect 15912 25094 16124 25100
rect 15912 25030 15918 25094
rect 15982 25030 16124 25094
rect 15912 24964 16124 25030
rect 16320 25024 17348 25100
rect 17408 25094 17620 25100
rect 17408 25030 17414 25094
rect 17478 25030 17620 25094
rect 15912 24888 16260 24964
rect 16320 24888 16532 25024
rect 17408 24964 17620 25030
rect 17816 24964 18028 25100
rect 18224 25094 18436 25100
rect 18224 25030 18230 25094
rect 18294 25030 18436 25094
rect 18224 24964 18436 25030
rect 17408 24958 17756 24964
rect 17408 24894 17686 24958
rect 17750 24894 17756 24958
rect 17408 24888 17756 24894
rect 17816 24958 18436 24964
rect 17816 24894 18230 24958
rect 18294 24894 18436 24958
rect 17816 24888 18436 24894
rect 18632 25094 18844 25100
rect 18632 25030 18774 25094
rect 18838 25030 18844 25094
rect 18632 24888 18844 25030
rect 19040 25094 19252 25100
rect 19040 25030 19182 25094
rect 19246 25030 19252 25094
rect 19040 24888 19252 25030
rect 20808 25094 21020 25100
rect 20808 25030 20814 25094
rect 20878 25030 21020 25094
rect 20808 24958 21020 25030
rect 20808 24894 20814 24958
rect 20878 24894 21020 24958
rect 20808 24888 21020 24894
rect 21216 25094 21564 25100
rect 21216 25030 21358 25094
rect 21422 25030 21494 25094
rect 21558 25030 21564 25094
rect 21216 25024 21564 25030
rect 21624 25094 21972 25100
rect 21624 25030 21766 25094
rect 21830 25030 21972 25094
rect 21216 24888 21428 25024
rect 21624 24958 21972 25030
rect 21624 24894 21902 24958
rect 21966 24894 21972 24958
rect 21624 24888 21972 24894
rect 22032 25094 22244 25100
rect 22032 25030 22174 25094
rect 22238 25030 22244 25094
rect 22032 24958 22244 25030
rect 22032 24894 22174 24958
rect 22238 24894 22244 24958
rect 22032 24888 22244 24894
rect 22440 25094 22652 25100
rect 22440 25030 22446 25094
rect 22510 25030 22652 25094
rect 22440 24958 22652 25030
rect 27336 25024 27684 25236
rect 109344 25024 109556 25236
rect 119136 25160 120436 25236
rect 119136 25100 119212 25160
rect 120360 25100 120436 25160
rect 27472 24964 27548 25024
rect 109480 24964 109556 25024
rect 22440 24894 22582 24958
rect 22646 24894 22652 24958
rect 22440 24888 22652 24894
rect 16184 24828 16260 24888
rect 17408 24828 17484 24888
rect 16184 24752 17484 24828
rect 27336 24752 27684 24964
rect 109344 24752 109556 24964
rect 114240 25094 114452 25100
rect 114240 25030 114246 25094
rect 114310 25030 114452 25094
rect 114240 24958 114452 25030
rect 114240 24894 114246 24958
rect 114310 24894 114452 24958
rect 114240 24888 114452 24894
rect 114648 25094 114860 25100
rect 114648 25030 114654 25094
rect 114718 25030 114860 25094
rect 114648 24958 114860 25030
rect 114648 24894 114654 24958
rect 114718 24894 114860 24958
rect 114648 24888 114860 24894
rect 115056 25094 115268 25100
rect 115056 25030 115198 25094
rect 115262 25030 115268 25094
rect 115056 24958 115268 25030
rect 115056 24894 115062 24958
rect 115126 24894 115268 24958
rect 115056 24888 115268 24894
rect 115464 25094 115676 25100
rect 115464 25030 115470 25094
rect 115534 25030 115676 25094
rect 115464 24958 115676 25030
rect 115464 24894 115470 24958
rect 115534 24894 115676 24958
rect 115464 24888 115676 24894
rect 115872 25094 116084 25100
rect 115872 25030 115878 25094
rect 115942 25030 116084 25094
rect 115872 24958 116084 25030
rect 115872 24894 116014 24958
rect 116078 24894 116084 24958
rect 115872 24888 116084 24894
rect 117640 25094 117852 25100
rect 117640 25030 117646 25094
rect 117710 25030 117852 25094
rect 117640 24958 117852 25030
rect 117640 24894 117646 24958
rect 117710 24894 117852 24958
rect 117640 24888 117852 24894
rect 118048 25094 118260 25100
rect 118048 25030 118190 25094
rect 118254 25030 118260 25094
rect 118048 24958 118260 25030
rect 118048 24894 118190 24958
rect 118254 24894 118260 24958
rect 118048 24888 118260 24894
rect 118456 24964 118668 25100
rect 118864 25094 119212 25100
rect 118864 25030 119006 25094
rect 119070 25030 119212 25094
rect 118864 25024 119212 25030
rect 119272 25094 119484 25100
rect 119272 25030 119414 25094
rect 119478 25030 119484 25094
rect 118864 24964 119076 25024
rect 118456 24888 119076 24964
rect 119272 24888 119484 25030
rect 120360 24888 120572 25100
rect 120768 25094 120980 25100
rect 120768 25030 120774 25094
rect 120838 25030 120980 25094
rect 120768 24888 120980 25030
rect 27608 24692 27684 24752
rect 109480 24692 109556 24752
rect 3128 24556 3340 24692
rect 3944 24556 4156 24692
rect 2350 24550 4156 24556
rect 2312 24486 2318 24550
rect 2382 24486 4156 24550
rect 2350 24480 4156 24486
rect 20808 24686 21020 24692
rect 20808 24622 20814 24686
rect 20878 24622 21020 24686
rect 20808 24550 21020 24622
rect 20808 24486 20950 24550
rect 21014 24486 21020 24550
rect 20808 24480 21020 24486
rect 21216 24686 21972 24692
rect 21216 24622 21902 24686
rect 21966 24622 21972 24686
rect 21216 24616 21972 24622
rect 21216 24480 21428 24616
rect 21624 24550 21972 24616
rect 21624 24486 21630 24550
rect 21694 24486 21972 24550
rect 21624 24480 21972 24486
rect 22032 24686 22244 24692
rect 22032 24622 22174 24686
rect 22238 24622 22244 24686
rect 22032 24550 22244 24622
rect 22032 24486 22038 24550
rect 22102 24486 22244 24550
rect 22032 24480 22244 24486
rect 22440 24686 22652 24692
rect 22440 24622 22582 24686
rect 22646 24622 22652 24686
rect 22440 24550 22652 24622
rect 22440 24486 22446 24550
rect 22510 24486 22652 24550
rect 22440 24480 22652 24486
rect 27336 24480 27684 24692
rect 27608 24420 27684 24480
rect 20808 24278 21020 24284
rect 20808 24214 20950 24278
rect 21014 24214 21020 24278
rect 20808 24072 21020 24214
rect 21216 24142 21428 24284
rect 21624 24278 21972 24284
rect 21624 24214 21630 24278
rect 21694 24214 21972 24278
rect 21624 24148 21972 24214
rect 21526 24142 21972 24148
rect 21216 24078 21222 24142
rect 21286 24078 21428 24142
rect 21488 24078 21494 24142
rect 21558 24078 21972 24142
rect 21216 24072 21428 24078
rect 21526 24072 21972 24078
rect 22032 24278 22244 24284
rect 22032 24214 22038 24278
rect 22102 24214 22244 24278
rect 22032 24142 22244 24214
rect 22032 24078 22038 24142
rect 22102 24078 22244 24142
rect 22032 24072 22244 24078
rect 22440 24278 22652 24284
rect 22440 24214 22446 24278
rect 22510 24214 22652 24278
rect 22440 24142 22652 24214
rect 22440 24078 22446 24142
rect 22510 24078 22652 24142
rect 22440 24072 22652 24078
rect 27336 24208 27684 24420
rect 109344 24480 109556 24692
rect 114240 24686 114452 24692
rect 114240 24622 114246 24686
rect 114310 24622 114452 24686
rect 114240 24550 114452 24622
rect 114240 24486 114382 24550
rect 114446 24486 114452 24550
rect 114240 24480 114452 24486
rect 114648 24686 114860 24692
rect 114648 24622 114654 24686
rect 114718 24622 114860 24686
rect 114648 24550 114860 24622
rect 114648 24486 114790 24550
rect 114854 24486 114860 24550
rect 114648 24480 114860 24486
rect 115056 24686 115268 24692
rect 115056 24622 115062 24686
rect 115126 24622 115268 24686
rect 115056 24480 115268 24622
rect 115464 24686 115676 24692
rect 115464 24622 115470 24686
rect 115534 24622 115676 24686
rect 115464 24480 115676 24622
rect 115872 24686 116084 24692
rect 115872 24622 116014 24686
rect 116078 24622 116084 24686
rect 115872 24550 116084 24622
rect 115872 24486 115878 24550
rect 115942 24486 116084 24550
rect 115872 24480 116084 24486
rect 109344 24420 109420 24480
rect 115464 24420 115540 24480
rect 109344 24208 109556 24420
rect 115192 24344 115540 24420
rect 115192 24284 115268 24344
rect 114240 24278 114452 24284
rect 114240 24214 114382 24278
rect 114446 24214 114452 24278
rect 27336 24148 27412 24208
rect 109344 24148 109420 24208
rect 20944 24012 21020 24072
rect 1224 24006 2388 24012
rect 1224 23942 1230 24006
rect 1294 23942 2318 24006
rect 2382 23942 2388 24006
rect 1224 23936 2388 23942
rect 1768 23928 1980 23936
rect 1768 23872 1794 23928
rect 1850 23872 1980 23928
rect 1768 23800 1980 23872
rect 20808 23664 21020 24012
rect 21352 23936 21700 24012
rect 27336 24006 27684 24148
rect 27336 23942 27614 24006
rect 27678 23942 27684 24006
rect 27336 23936 27684 23942
rect 109344 23936 109556 24148
rect 114240 24142 114452 24214
rect 114240 24078 114246 24142
rect 114310 24078 114452 24142
rect 114240 24072 114452 24078
rect 114648 24278 114860 24284
rect 114648 24214 114790 24278
rect 114854 24214 114860 24278
rect 114648 24142 114860 24214
rect 114648 24078 114790 24142
rect 114854 24078 114860 24142
rect 114648 24072 114860 24078
rect 115056 24208 115676 24284
rect 115056 24142 115268 24208
rect 115056 24078 115198 24142
rect 115262 24078 115268 24142
rect 115056 24072 115268 24078
rect 115464 24142 115676 24208
rect 115464 24078 115606 24142
rect 115670 24078 115676 24142
rect 115464 24072 115676 24078
rect 115872 24278 116084 24284
rect 115872 24214 115878 24278
rect 115942 24214 116084 24278
rect 115872 24072 116084 24214
rect 21352 23876 21428 23936
rect 21624 23876 21700 23936
rect 27608 23876 27684 23936
rect 109480 23876 109556 23936
rect 115872 24012 115948 24072
rect 21216 23870 21564 23876
rect 21216 23806 21222 23870
rect 21286 23806 21494 23870
rect 21558 23806 21564 23870
rect 21216 23800 21564 23806
rect 21216 23740 21428 23800
rect 21216 23664 21564 23740
rect 21624 23664 21972 23876
rect 22032 23870 22244 23876
rect 22032 23806 22038 23870
rect 22102 23806 22244 23870
rect 22032 23734 22244 23806
rect 22032 23670 22174 23734
rect 22238 23670 22244 23734
rect 22032 23664 22244 23670
rect 22440 23870 22652 23876
rect 22440 23806 22446 23870
rect 22510 23806 22652 23870
rect 22440 23734 22652 23806
rect 22440 23670 22446 23734
rect 22510 23670 22652 23734
rect 22440 23664 22652 23670
rect 27336 23734 27684 23876
rect 27336 23670 27478 23734
rect 27542 23670 27614 23734
rect 27678 23670 27684 23734
rect 20808 23604 20884 23664
rect 21488 23604 21564 23664
rect 18496 23528 19116 23604
rect 18496 23468 18572 23528
rect 19040 23468 19116 23528
rect 3264 23392 4020 23468
rect 17718 23462 18028 23468
rect 17680 23398 17686 23462
rect 17750 23398 18028 23462
rect 17718 23392 18028 23398
rect 3264 23332 3340 23392
rect 3944 23332 4020 23392
rect 17816 23332 18028 23392
rect 18224 23462 18572 23468
rect 18224 23398 18230 23462
rect 18294 23398 18572 23462
rect 18224 23392 18572 23398
rect 3128 23326 3884 23332
rect 3128 23262 3814 23326
rect 3878 23262 3884 23326
rect 3128 23256 3884 23262
rect 3128 23196 3340 23256
rect 544 23190 3884 23196
rect 544 23126 550 23190
rect 614 23126 3814 23190
rect 3878 23126 3884 23190
rect 544 23120 3884 23126
rect 3944 23120 4156 23332
rect 17816 23256 18164 23332
rect 18224 23326 18436 23392
rect 18224 23262 18230 23326
rect 18294 23262 18436 23326
rect 18224 23256 18436 23262
rect 18632 23326 18844 23468
rect 18632 23262 18638 23326
rect 18702 23262 18844 23326
rect 18632 23256 18844 23262
rect 19040 23326 19252 23468
rect 19040 23262 19046 23326
rect 19110 23262 19252 23326
rect 19040 23256 19252 23262
rect 20808 23256 21020 23604
rect 21216 23326 21428 23604
rect 21488 23528 21972 23604
rect 21216 23262 21358 23326
rect 21422 23262 21428 23326
rect 21216 23256 21428 23262
rect 21624 23326 21972 23528
rect 21624 23262 21630 23326
rect 21694 23262 21972 23326
rect 21624 23256 21972 23262
rect 22032 23462 22244 23468
rect 22032 23398 22174 23462
rect 22238 23398 22244 23462
rect 22032 23326 22244 23398
rect 22032 23262 22038 23326
rect 22102 23262 22244 23326
rect 22032 23256 22244 23262
rect 22440 23462 22652 23468
rect 22440 23398 22446 23462
rect 22510 23398 22652 23462
rect 22440 23326 22652 23398
rect 27336 23392 27684 23670
rect 109344 23392 109556 23876
rect 114240 23870 114452 23876
rect 114240 23806 114246 23870
rect 114310 23806 114452 23870
rect 114240 23734 114452 23806
rect 114240 23670 114246 23734
rect 114310 23670 114452 23734
rect 114240 23664 114452 23670
rect 114648 23870 114860 23876
rect 114648 23806 114790 23870
rect 114854 23806 114860 23870
rect 114648 23734 114860 23806
rect 114648 23670 114790 23734
rect 114854 23670 114860 23734
rect 114648 23664 114860 23670
rect 115056 23870 115268 23876
rect 115056 23806 115198 23870
rect 115262 23806 115268 23870
rect 115056 23664 115268 23806
rect 115464 23870 115676 23876
rect 115464 23806 115606 23870
rect 115670 23806 115676 23870
rect 115464 23664 115676 23806
rect 115872 23664 116084 24012
rect 134776 23928 134988 24012
rect 134776 23872 134844 23928
rect 134900 23876 134988 23928
rect 134900 23872 135396 23876
rect 134776 23870 135396 23872
rect 134776 23806 135326 23870
rect 135390 23806 135396 23870
rect 134776 23800 135396 23806
rect 115056 23604 115132 23664
rect 115600 23604 115676 23664
rect 116008 23604 116084 23664
rect 114240 23462 114452 23468
rect 114240 23398 114246 23462
rect 114310 23398 114452 23462
rect 109344 23332 109420 23392
rect 22440 23262 22582 23326
rect 22646 23262 22652 23326
rect 22440 23256 22652 23262
rect 27336 23326 27684 23332
rect 27336 23262 27478 23326
rect 27542 23262 27684 23326
rect 18088 23196 18164 23256
rect 18632 23196 18708 23256
rect 20944 23196 21020 23256
rect 18088 23120 18708 23196
rect 20808 23054 21020 23196
rect 27336 23190 27684 23262
rect 27336 23126 27342 23190
rect 27406 23126 27684 23190
rect 27336 23120 27684 23126
rect 109344 23190 109556 23332
rect 114240 23326 114452 23398
rect 114240 23262 114382 23326
rect 114446 23262 114452 23326
rect 114240 23256 114452 23262
rect 114648 23462 114860 23468
rect 114648 23398 114790 23462
rect 114854 23398 114860 23462
rect 114648 23326 114860 23398
rect 114648 23262 114790 23326
rect 114854 23262 114860 23326
rect 114648 23256 114860 23262
rect 115056 23256 115268 23604
rect 115464 23256 115676 23604
rect 115872 23256 116084 23604
rect 117640 23462 117852 23468
rect 117640 23398 117646 23462
rect 117710 23398 117852 23462
rect 117640 23326 117852 23398
rect 117640 23262 117646 23326
rect 117710 23262 117852 23326
rect 117640 23256 117852 23262
rect 118048 23462 118260 23468
rect 118048 23398 118190 23462
rect 118254 23398 118260 23462
rect 118048 23326 118260 23398
rect 118048 23262 118054 23326
rect 118118 23262 118260 23326
rect 118048 23256 118260 23262
rect 118456 23326 118668 23468
rect 118456 23262 118598 23326
rect 118662 23262 118668 23326
rect 118456 23256 118668 23262
rect 118864 23326 119076 23468
rect 118864 23262 119006 23326
rect 119070 23262 119076 23326
rect 118864 23256 119076 23262
rect 115464 23196 115540 23256
rect 109344 23126 109350 23190
rect 109414 23126 109556 23190
rect 109344 23120 109556 23126
rect 115192 23120 115540 23196
rect 115872 23196 115948 23256
rect 27472 23060 27548 23120
rect 109344 23060 109420 23120
rect 115192 23060 115268 23120
rect 20808 22990 20950 23054
rect 21014 22990 21020 23054
rect 20808 22984 21020 22990
rect 21216 23054 21564 23060
rect 21216 22990 21358 23054
rect 21422 22990 21494 23054
rect 21558 22990 21564 23054
rect 21216 22984 21564 22990
rect 21624 23054 21972 23060
rect 21624 22990 21630 23054
rect 21694 22990 21972 23054
rect 21216 22924 21428 22984
rect 21624 22924 21972 22990
rect 17680 22848 18300 22924
rect 21216 22848 21972 22924
rect 22032 23054 22244 23060
rect 22032 22990 22038 23054
rect 22102 22990 22244 23054
rect 22032 22848 22244 22990
rect 17680 22788 17756 22848
rect 18224 22788 18300 22848
rect 21352 22788 21428 22848
rect 22168 22788 22244 22848
rect 16592 22516 16804 22788
rect 17000 22712 17756 22788
rect 16592 22440 16940 22516
rect 17000 22440 17212 22712
rect 17816 22516 18028 22788
rect 18224 22782 18436 22788
rect 18224 22718 18230 22782
rect 18294 22718 18436 22782
rect 17816 22440 18164 22516
rect 18224 22510 18436 22718
rect 18224 22446 18366 22510
rect 18430 22446 18436 22510
rect 18224 22440 18436 22446
rect 18632 22782 18844 22788
rect 18632 22718 18638 22782
rect 18702 22718 18844 22782
rect 18632 22510 18844 22718
rect 18632 22446 18638 22510
rect 18702 22446 18844 22510
rect 18632 22440 18844 22446
rect 19040 22782 19252 22788
rect 19040 22718 19046 22782
rect 19110 22718 19252 22782
rect 19040 22440 19252 22718
rect 20808 22782 21020 22788
rect 20808 22718 20950 22782
rect 21014 22718 21020 22782
rect 20808 22646 21020 22718
rect 20808 22582 20814 22646
rect 20878 22582 21020 22646
rect 20808 22576 21020 22582
rect 21216 22576 21428 22788
rect 21526 22782 21972 22788
rect 21488 22718 21494 22782
rect 21558 22718 21972 22782
rect 21526 22712 21972 22718
rect 21624 22646 21972 22712
rect 21624 22582 21630 22646
rect 21694 22582 21972 22646
rect 21624 22576 21972 22582
rect 22032 22440 22244 22788
rect 22440 23054 22652 23060
rect 22440 22990 22582 23054
rect 22646 22990 22652 23054
rect 22440 22848 22652 22990
rect 27336 22918 27684 23060
rect 27336 22854 27342 22918
rect 27406 22854 27684 22918
rect 22440 22788 22516 22848
rect 22440 22440 22652 22788
rect 27336 22782 27684 22854
rect 27336 22718 27478 22782
rect 27542 22718 27684 22782
rect 27336 22712 27684 22718
rect 109344 22918 109556 23060
rect 109344 22854 109350 22918
rect 109414 22854 109556 22918
rect 109344 22782 109556 22854
rect 109344 22718 109486 22782
rect 109550 22718 109556 22782
rect 109344 22712 109556 22718
rect 114240 23054 114452 23060
rect 114240 22990 114382 23054
rect 114446 22990 114452 23054
rect 114240 22848 114452 22990
rect 114648 23054 114860 23060
rect 114648 22990 114790 23054
rect 114854 22990 114860 23054
rect 114648 22848 114860 22990
rect 115056 22984 115676 23060
rect 115872 23054 116084 23196
rect 118358 23054 118940 23060
rect 115872 22990 116014 23054
rect 116078 22990 116084 23054
rect 118320 22990 118326 23054
rect 118390 22990 118870 23054
rect 118934 22990 118940 23054
rect 115872 22984 116084 22990
rect 118358 22984 118940 22990
rect 115056 22924 115268 22984
rect 115056 22848 115404 22924
rect 115464 22848 115676 22984
rect 118728 22848 119756 22924
rect 114240 22788 114316 22848
rect 114648 22788 114724 22848
rect 115056 22788 115132 22848
rect 115328 22788 115404 22848
rect 118728 22788 118804 22848
rect 119680 22788 119756 22848
rect 16864 22380 16940 22440
rect 17816 22380 17892 22440
rect 1224 22374 1980 22380
rect 1224 22310 1230 22374
rect 1294 22310 1980 22374
rect 1224 22304 1980 22310
rect 16864 22304 17892 22380
rect 18088 22380 18164 22440
rect 18632 22380 18708 22440
rect 22032 22380 22108 22440
rect 22576 22380 22652 22440
rect 18088 22304 18708 22380
rect 20808 22374 21020 22380
rect 20808 22310 20814 22374
rect 20878 22310 21020 22374
rect 1768 22248 1980 22304
rect 1768 22192 1794 22248
rect 1850 22244 1980 22248
rect 1850 22238 3204 22244
rect 1850 22192 3134 22238
rect 1768 22174 3134 22192
rect 3198 22174 3204 22238
rect 1768 22168 3204 22174
rect 20808 22238 21020 22310
rect 20808 22174 20950 22238
rect 21014 22174 21020 22238
rect 20808 22168 21020 22174
rect 21216 22032 21428 22380
rect 21624 22374 21972 22380
rect 21624 22310 21630 22374
rect 21694 22310 21972 22374
rect 21624 22108 21972 22310
rect 21488 22032 21972 22108
rect 22032 22032 22244 22380
rect 22440 22032 22652 22380
rect 21216 21972 21292 22032
rect 21488 21972 21564 22032
rect 22032 21972 22108 22032
rect 22576 21972 22652 22032
rect 20808 21966 21020 21972
rect 20808 21902 20950 21966
rect 21014 21902 21020 21966
rect 3128 21830 3340 21836
rect 3128 21766 3134 21830
rect 3198 21766 3340 21830
rect 3128 21700 3340 21766
rect 3944 21700 4156 21836
rect 20808 21830 21020 21902
rect 20808 21766 20950 21830
rect 21014 21766 21020 21830
rect 20808 21760 21020 21766
rect 21216 21896 21564 21972
rect 21216 21830 21428 21896
rect 21624 21836 21972 21972
rect 21526 21830 21972 21836
rect 21216 21766 21358 21830
rect 21422 21766 21428 21830
rect 21488 21766 21494 21830
rect 21558 21766 21766 21830
rect 21830 21766 21972 21830
rect 21216 21760 21428 21766
rect 21526 21760 21972 21766
rect 22032 21830 22244 21972
rect 22032 21766 22174 21830
rect 22238 21766 22244 21830
rect 22032 21760 22244 21766
rect 22440 21830 22652 21972
rect 27336 22510 27684 22516
rect 27336 22446 27478 22510
rect 27542 22446 27684 22510
rect 27336 22374 27684 22446
rect 27336 22310 27342 22374
rect 27406 22310 27684 22374
rect 27336 22102 27684 22310
rect 27336 22038 27342 22102
rect 27406 22038 27684 22102
rect 27336 21896 27684 22038
rect 109344 22510 109556 22516
rect 109344 22446 109486 22510
rect 109550 22446 109556 22510
rect 109344 22374 109556 22446
rect 114240 22440 114452 22788
rect 114648 22440 114860 22788
rect 115056 22646 115268 22788
rect 115328 22712 115676 22788
rect 115056 22582 115062 22646
rect 115126 22582 115268 22646
rect 115056 22576 115268 22582
rect 115464 22576 115676 22712
rect 115872 22782 116084 22788
rect 115872 22718 116014 22782
rect 116078 22718 116084 22782
rect 115872 22646 116084 22718
rect 115872 22582 115878 22646
rect 115942 22582 116084 22646
rect 115872 22576 116084 22582
rect 117640 22782 117852 22788
rect 117640 22718 117646 22782
rect 117710 22718 117852 22782
rect 117640 22516 117852 22718
rect 118048 22782 118396 22788
rect 118048 22718 118054 22782
rect 118118 22718 118326 22782
rect 118390 22718 118396 22782
rect 118048 22712 118396 22718
rect 118456 22782 118804 22788
rect 118456 22718 118598 22782
rect 118662 22718 118804 22782
rect 118456 22712 118804 22718
rect 118864 22782 119076 22788
rect 118864 22718 118870 22782
rect 118934 22718 119006 22782
rect 119070 22718 119076 22782
rect 117640 22440 117988 22516
rect 118048 22440 118260 22712
rect 118456 22510 118668 22712
rect 118456 22446 118462 22510
rect 118526 22446 118668 22510
rect 118456 22440 118668 22446
rect 118864 22516 119076 22718
rect 118864 22510 119620 22516
rect 118864 22446 118870 22510
rect 118934 22446 119620 22510
rect 118864 22440 119620 22446
rect 119680 22440 120028 22788
rect 120088 22440 120300 22788
rect 114376 22380 114452 22440
rect 114784 22380 114860 22440
rect 117912 22380 117988 22440
rect 118456 22380 118532 22440
rect 109344 22310 109350 22374
rect 109414 22310 109556 22374
rect 109344 22102 109556 22310
rect 109344 22038 109350 22102
rect 109414 22038 109556 22102
rect 109344 21896 109556 22038
rect 114240 22032 114452 22380
rect 114648 22032 114860 22380
rect 115056 22374 115268 22380
rect 115056 22310 115062 22374
rect 115126 22310 115268 22374
rect 115056 22032 115268 22310
rect 115464 22108 115676 22380
rect 115872 22374 116084 22380
rect 115872 22310 115878 22374
rect 115942 22310 116084 22374
rect 115872 22238 116084 22310
rect 117912 22304 118532 22380
rect 119544 22380 119620 22440
rect 120088 22380 120164 22440
rect 119544 22304 120164 22380
rect 134776 22248 134988 22380
rect 118358 22238 118940 22244
rect 115872 22174 115878 22238
rect 115942 22174 116084 22238
rect 118320 22174 118326 22238
rect 118390 22174 118870 22238
rect 118934 22174 118940 22238
rect 115872 22168 116084 22174
rect 118358 22168 118940 22174
rect 134776 22192 134844 22248
rect 134900 22244 134988 22248
rect 134900 22238 135396 22244
rect 134900 22192 135326 22238
rect 134776 22174 135326 22192
rect 135390 22174 135396 22238
rect 134776 22168 135396 22174
rect 114240 21972 114316 22032
rect 114648 21972 114724 22032
rect 115192 21972 115268 22032
rect 115328 22032 115676 22108
rect 115328 21972 115404 22032
rect 27472 21836 27548 21896
rect 109344 21836 109420 21896
rect 22440 21766 22446 21830
rect 22510 21766 22652 21830
rect 22440 21760 22652 21766
rect 3128 21624 4156 21700
rect 20808 21558 21020 21564
rect 20808 21494 20950 21558
rect 21014 21494 21020 21558
rect 20808 21422 21020 21494
rect 20808 21358 20950 21422
rect 21014 21358 21020 21422
rect 20808 21352 21020 21358
rect 21216 21558 21564 21564
rect 21216 21494 21358 21558
rect 21422 21494 21494 21558
rect 21558 21494 21564 21558
rect 21216 21488 21564 21494
rect 21624 21558 21972 21564
rect 21624 21494 21766 21558
rect 21830 21494 21972 21558
rect 21216 21352 21428 21488
rect 21624 21422 21972 21494
rect 21624 21358 21630 21422
rect 21694 21358 21972 21422
rect 21624 21352 21972 21358
rect 22032 21558 22244 21564
rect 22032 21494 22174 21558
rect 22238 21494 22244 21558
rect 22032 21422 22244 21494
rect 22032 21358 22174 21422
rect 22238 21358 22244 21422
rect 22032 21352 22244 21358
rect 22440 21558 22652 21564
rect 22440 21494 22446 21558
rect 22510 21494 22652 21558
rect 22440 21422 22652 21494
rect 22440 21358 22446 21422
rect 22510 21358 22652 21422
rect 22440 21352 22652 21358
rect 27336 21352 27684 21836
rect 27608 21292 27684 21352
rect 18088 21216 18708 21292
rect 18088 21156 18164 21216
rect 18632 21156 18708 21216
rect 17816 21080 18164 21156
rect 18224 21150 18436 21156
rect 18224 21086 18366 21150
rect 18430 21086 18436 21150
rect 17816 21014 18028 21080
rect 17816 20950 17822 21014
rect 17886 20950 18028 21014
rect 17816 20944 18028 20950
rect 18224 21020 18436 21086
rect 18632 21150 18844 21156
rect 18632 21086 18638 21150
rect 18702 21086 18844 21150
rect 18224 21014 18572 21020
rect 18224 20950 18366 21014
rect 18430 20950 18572 21014
rect 18224 20944 18572 20950
rect 18632 21014 18844 21086
rect 18632 20950 18638 21014
rect 18702 20950 18844 21014
rect 18632 20944 18844 20950
rect 19040 21014 19252 21156
rect 19040 20950 19182 21014
rect 19246 20950 19252 21014
rect 19040 20944 19252 20950
rect 20808 21150 21020 21156
rect 20808 21086 20950 21150
rect 21014 21086 21020 21150
rect 20808 21014 21020 21086
rect 20808 20950 20814 21014
rect 20878 20950 21020 21014
rect 20808 20944 21020 20950
rect 21216 21014 21428 21156
rect 21216 20950 21358 21014
rect 21422 20950 21428 21014
rect 21216 20944 21428 20950
rect 21624 21150 21972 21156
rect 21624 21086 21630 21150
rect 21694 21086 21972 21150
rect 21624 21014 21972 21086
rect 21624 20950 21766 21014
rect 21830 20950 21972 21014
rect 21624 20944 21972 20950
rect 22032 21150 22244 21156
rect 22032 21086 22174 21150
rect 22238 21086 22244 21150
rect 22032 21014 22244 21086
rect 22032 20950 22038 21014
rect 22102 20950 22244 21014
rect 22032 20944 22244 20950
rect 22440 21150 22652 21156
rect 22440 21086 22446 21150
rect 22510 21086 22652 21150
rect 22440 21014 22652 21086
rect 22440 20950 22446 21014
rect 22510 20950 22652 21014
rect 22440 20944 22652 20950
rect 27336 21080 27684 21292
rect 109344 21558 109556 21836
rect 114240 21830 114452 21972
rect 114240 21766 114246 21830
rect 114310 21766 114452 21830
rect 114240 21760 114452 21766
rect 114648 21830 114860 21972
rect 114648 21766 114654 21830
rect 114718 21766 114860 21830
rect 114648 21760 114860 21766
rect 115056 21896 115404 21972
rect 115056 21836 115268 21896
rect 115464 21836 115676 21972
rect 115056 21830 115676 21836
rect 115056 21766 115062 21830
rect 115126 21766 115606 21830
rect 115670 21766 115676 21830
rect 115056 21760 115676 21766
rect 115872 21966 116084 21972
rect 115872 21902 115878 21966
rect 115942 21902 116084 21966
rect 115872 21830 116084 21902
rect 115872 21766 116014 21830
rect 116078 21766 116084 21830
rect 115872 21760 116084 21766
rect 109344 21494 109350 21558
rect 109414 21494 109556 21558
rect 109344 21352 109556 21494
rect 114240 21558 114452 21564
rect 114240 21494 114246 21558
rect 114310 21494 114452 21558
rect 114240 21422 114452 21494
rect 114240 21358 114246 21422
rect 114310 21358 114452 21422
rect 114240 21352 114452 21358
rect 114648 21558 114860 21564
rect 114648 21494 114654 21558
rect 114718 21494 114860 21558
rect 114648 21422 114860 21494
rect 114648 21358 114654 21422
rect 114718 21358 114860 21422
rect 114648 21352 114860 21358
rect 115056 21558 115268 21564
rect 115056 21494 115062 21558
rect 115126 21494 115268 21558
rect 115056 21352 115268 21494
rect 115464 21558 115676 21564
rect 115464 21494 115606 21558
rect 115670 21494 115676 21558
rect 115464 21422 115676 21494
rect 115464 21358 115606 21422
rect 115670 21358 115676 21422
rect 115464 21352 115676 21358
rect 115872 21558 116084 21564
rect 115872 21494 116014 21558
rect 116078 21494 116084 21558
rect 115872 21428 116084 21494
rect 115872 21422 118124 21428
rect 115872 21358 115878 21422
rect 115942 21358 118054 21422
rect 118118 21358 118124 21422
rect 115872 21352 118124 21358
rect 109344 21292 109420 21352
rect 109344 21286 109556 21292
rect 109344 21222 109350 21286
rect 109414 21222 109556 21286
rect 109344 21080 109556 21222
rect 117912 21286 118532 21292
rect 117912 21222 118462 21286
rect 118526 21222 118532 21286
rect 117912 21216 118532 21222
rect 117912 21156 117988 21216
rect 114240 21150 114452 21156
rect 114240 21086 114246 21150
rect 114310 21086 114452 21150
rect 27336 21020 27412 21080
rect 109344 21020 109420 21080
rect 18496 20884 18572 20944
rect 19040 20884 19116 20944
rect 18496 20808 19116 20884
rect 27336 20808 27684 21020
rect 109344 20808 109556 21020
rect 114240 21014 114452 21086
rect 114240 20950 114246 21014
rect 114310 20950 114452 21014
rect 114240 20944 114452 20950
rect 114648 21150 114860 21156
rect 114648 21086 114654 21150
rect 114718 21086 114860 21150
rect 114648 21014 114860 21086
rect 114648 20950 114654 21014
rect 114718 20950 114860 21014
rect 114648 20944 114860 20950
rect 115056 21150 115676 21156
rect 115056 21086 115606 21150
rect 115670 21086 115676 21150
rect 115056 21080 115676 21086
rect 115056 21020 115268 21080
rect 115056 21014 115404 21020
rect 115056 20950 115198 21014
rect 115262 20950 115334 21014
rect 115398 20950 115404 21014
rect 115056 20944 115404 20950
rect 115464 20944 115676 21080
rect 115872 21150 116084 21156
rect 115872 21086 115878 21150
rect 115942 21086 116084 21150
rect 115872 21014 116084 21086
rect 115872 20950 116014 21014
rect 116078 20950 116084 21014
rect 115872 20944 116084 20950
rect 117640 21080 117988 21156
rect 118048 21150 118396 21156
rect 118048 21086 118054 21150
rect 118118 21086 118326 21150
rect 118390 21086 118396 21150
rect 118048 21080 118396 21086
rect 117640 21020 117852 21080
rect 117640 21014 117988 21020
rect 117640 20950 117646 21014
rect 117710 20950 117988 21014
rect 117640 20944 117988 20950
rect 118048 21014 118260 21080
rect 118048 20950 118190 21014
rect 118254 20950 118260 21014
rect 118048 20944 118260 20950
rect 118456 21014 118668 21156
rect 118456 20950 118598 21014
rect 118662 20950 118668 21014
rect 118456 20944 118668 20950
rect 118864 21014 119076 21156
rect 118864 20950 119006 21014
rect 119070 20950 119076 21014
rect 118864 20944 119076 20950
rect 117912 20884 117988 20944
rect 118456 20884 118532 20944
rect 117912 20808 118532 20884
rect 27336 20748 27412 20808
rect 109344 20748 109420 20808
rect 20808 20742 21020 20748
rect 20808 20678 20814 20742
rect 20878 20678 21020 20742
rect 1224 20606 1980 20612
rect 1224 20542 1230 20606
rect 1294 20568 1980 20606
rect 1294 20542 1794 20568
rect 1224 20536 1794 20542
rect 1768 20512 1794 20536
rect 1850 20512 1980 20568
rect 20808 20606 21020 20678
rect 20808 20542 20950 20606
rect 21014 20542 21020 20606
rect 20808 20536 21020 20542
rect 21216 20742 21972 20748
rect 21216 20678 21358 20742
rect 21422 20678 21766 20742
rect 21830 20678 21972 20742
rect 21216 20672 21972 20678
rect 21216 20606 21428 20672
rect 21216 20542 21358 20606
rect 21422 20542 21428 20606
rect 21216 20536 21428 20542
rect 21624 20606 21972 20672
rect 21624 20542 21766 20606
rect 21830 20542 21972 20606
rect 21624 20536 21972 20542
rect 22032 20742 22244 20748
rect 22032 20678 22038 20742
rect 22102 20678 22244 20742
rect 22032 20606 22244 20678
rect 22032 20542 22174 20606
rect 22238 20542 22244 20606
rect 22032 20536 22244 20542
rect 22440 20742 22652 20748
rect 22440 20678 22446 20742
rect 22510 20678 22652 20742
rect 22440 20606 22652 20678
rect 22440 20542 22446 20606
rect 22510 20542 22652 20606
rect 22440 20536 22652 20542
rect 27336 20536 27684 20748
rect 109344 20536 109556 20748
rect 114240 20742 114452 20748
rect 114240 20678 114246 20742
rect 114310 20678 114452 20742
rect 114240 20606 114452 20678
rect 114240 20542 114246 20606
rect 114310 20542 114452 20606
rect 114240 20536 114452 20542
rect 114648 20742 114860 20748
rect 114648 20678 114654 20742
rect 114718 20678 114860 20742
rect 114648 20606 114860 20678
rect 114648 20542 114654 20606
rect 114718 20542 114860 20606
rect 114648 20536 114860 20542
rect 115056 20742 115268 20748
rect 115366 20742 115676 20748
rect 115056 20678 115198 20742
rect 115262 20678 115268 20742
rect 115328 20678 115334 20742
rect 115398 20678 115676 20742
rect 115056 20606 115268 20678
rect 115366 20672 115676 20678
rect 115056 20542 115062 20606
rect 115126 20542 115268 20606
rect 115056 20536 115268 20542
rect 115464 20606 115676 20672
rect 115464 20542 115470 20606
rect 115534 20542 115676 20606
rect 115464 20536 115676 20542
rect 115872 20742 116084 20748
rect 115872 20678 116014 20742
rect 116078 20678 116084 20742
rect 115872 20606 116084 20678
rect 115872 20542 116014 20606
rect 116078 20542 116084 20606
rect 115872 20536 116084 20542
rect 134776 20606 135396 20612
rect 134776 20568 135326 20606
rect 1768 20400 1980 20512
rect 27472 20476 27548 20536
rect 109480 20476 109556 20536
rect 134776 20512 134844 20568
rect 134900 20542 135326 20568
rect 135390 20542 135396 20606
rect 134900 20536 135396 20542
rect 134900 20512 134988 20536
rect 3128 20470 3748 20476
rect 3846 20470 4156 20476
rect 3128 20406 3678 20470
rect 3742 20406 3748 20470
rect 3808 20406 3814 20470
rect 3878 20406 4156 20470
rect 3128 20400 3748 20406
rect 3846 20400 4156 20406
rect 3128 20340 3340 20400
rect 3944 20340 4156 20400
rect 17680 20400 18300 20476
rect 17680 20340 17756 20400
rect 18224 20340 18300 20400
rect 3128 20264 4156 20340
rect 16592 20204 16804 20340
rect 17000 20264 17756 20340
rect 17816 20334 18028 20340
rect 17816 20270 17822 20334
rect 17886 20270 18028 20334
rect 16592 20198 16940 20204
rect 16592 20134 16598 20198
rect 16662 20134 16940 20198
rect 16592 20128 16940 20134
rect 17000 20198 17212 20264
rect 17000 20134 17006 20198
rect 17070 20134 17212 20198
rect 17000 20128 17212 20134
rect 17816 20128 18028 20270
rect 18224 20334 18436 20340
rect 18224 20270 18366 20334
rect 18430 20270 18436 20334
rect 18224 20128 18436 20270
rect 18632 20334 18844 20340
rect 18632 20270 18638 20334
rect 18702 20270 18844 20334
rect 18632 20128 18844 20270
rect 19040 20334 19252 20340
rect 19040 20270 19182 20334
rect 19246 20270 19252 20334
rect 19040 20128 19252 20270
rect 20808 20334 21020 20340
rect 20808 20270 20950 20334
rect 21014 20270 21020 20334
rect 20808 20204 21020 20270
rect 21216 20334 21428 20340
rect 21216 20270 21358 20334
rect 21422 20270 21428 20334
rect 20808 20198 21156 20204
rect 20808 20134 21086 20198
rect 21150 20134 21156 20198
rect 20808 20128 21156 20134
rect 21216 20128 21428 20270
rect 21624 20334 21972 20340
rect 21624 20270 21766 20334
rect 21830 20270 21972 20334
rect 21624 20128 21972 20270
rect 22032 20334 22244 20340
rect 22032 20270 22174 20334
rect 22238 20270 22244 20334
rect 22032 20128 22244 20270
rect 22440 20334 22652 20340
rect 22440 20270 22446 20334
rect 22510 20270 22652 20334
rect 22440 20198 22652 20270
rect 27336 20264 27684 20476
rect 109344 20264 109556 20476
rect 118728 20400 119756 20476
rect 134776 20400 134988 20512
rect 118728 20340 118804 20400
rect 119680 20340 119756 20400
rect 27608 20204 27684 20264
rect 109480 20204 109556 20264
rect 22440 20134 22446 20198
rect 22510 20134 22652 20198
rect 22440 20128 22652 20134
rect 16864 20068 16940 20128
rect 17816 20068 17892 20128
rect 16864 19992 17892 20068
rect 27336 19992 27684 20204
rect 109344 20068 109556 20204
rect 114240 20334 114452 20340
rect 114240 20270 114246 20334
rect 114310 20270 114452 20334
rect 114240 20128 114452 20270
rect 114648 20334 114860 20340
rect 114648 20270 114654 20334
rect 114718 20270 114860 20334
rect 114648 20128 114860 20270
rect 115056 20334 115268 20340
rect 115056 20270 115062 20334
rect 115126 20270 115268 20334
rect 115056 20128 115268 20270
rect 115464 20334 115676 20340
rect 115464 20270 115470 20334
rect 115534 20270 115676 20334
rect 115464 20128 115676 20270
rect 115872 20334 116084 20340
rect 115872 20270 116014 20334
rect 116078 20270 116084 20334
rect 115872 20128 116084 20270
rect 117640 20334 117852 20340
rect 117640 20270 117646 20334
rect 117710 20270 117852 20334
rect 117640 20128 117852 20270
rect 118048 20334 118260 20340
rect 118048 20270 118190 20334
rect 118254 20270 118260 20334
rect 118048 20204 118260 20270
rect 118456 20334 118804 20340
rect 118456 20270 118598 20334
rect 118662 20270 118804 20334
rect 118456 20264 118804 20270
rect 118864 20334 119076 20340
rect 118864 20270 119006 20334
rect 119070 20270 119076 20334
rect 118048 20128 118396 20204
rect 118456 20128 118668 20264
rect 118864 20204 119076 20270
rect 118864 20128 119620 20204
rect 119680 20198 120028 20340
rect 119680 20134 119958 20198
rect 120022 20134 120028 20198
rect 119680 20128 120028 20134
rect 120088 20204 120300 20340
rect 120088 20198 122884 20204
rect 120088 20134 122814 20198
rect 122878 20134 122884 20198
rect 120088 20128 122884 20134
rect 118320 20068 118396 20128
rect 118864 20068 118940 20128
rect 109344 20062 109692 20068
rect 109344 19998 109622 20062
rect 109686 19998 109692 20062
rect 109344 19992 109692 19998
rect 118320 19992 118940 20068
rect 119544 20068 119620 20128
rect 120088 20068 120164 20128
rect 119544 19992 120164 20068
rect 27472 19932 27548 19992
rect 109344 19932 109420 19992
rect 27336 19796 27684 19932
rect 22440 19790 22652 19796
rect 22440 19726 22446 19790
rect 22510 19726 22652 19790
rect 22440 19660 22652 19726
rect 23256 19660 23604 19796
rect 25976 19660 26188 19796
rect 27064 19790 29044 19796
rect 27064 19726 28974 19790
rect 29038 19726 29044 19790
rect 27064 19720 29044 19726
rect 109344 19720 109556 19932
rect 122808 19926 123020 19932
rect 122808 19862 122814 19926
rect 122878 19862 123020 19926
rect 109616 19790 109828 19796
rect 109616 19726 109622 19790
rect 109686 19726 109828 19790
rect 22440 19654 27004 19660
rect 22440 19590 22446 19654
rect 22510 19590 26934 19654
rect 26998 19590 27004 19654
rect 22440 19584 27004 19590
rect 27064 19584 27276 19720
rect 109616 19584 109828 19726
rect 122808 19790 123020 19862
rect 122808 19726 122814 19790
rect 122878 19726 123020 19790
rect 122808 19720 123020 19726
rect 122216 19571 122300 19575
rect 122183 19566 122300 19571
rect 122183 19510 122188 19566
rect 122244 19510 122300 19566
rect 122183 19505 122300 19510
rect 122216 19501 122300 19505
rect 26966 19382 28908 19388
rect 26928 19318 26934 19382
rect 26998 19318 28908 19382
rect 26966 19312 28908 19318
rect 28152 19252 28364 19312
rect 28696 19252 28908 19312
rect 29376 19312 30812 19388
rect 29376 19252 29588 19312
rect 28152 19246 28636 19252
rect 28152 19182 28294 19246
rect 28358 19182 28566 19246
rect 28630 19182 28636 19246
rect 28152 19176 28636 19182
rect 28696 19246 29588 19252
rect 28696 19182 29518 19246
rect 29582 19182 29588 19246
rect 28696 19176 29588 19182
rect 29920 19176 30132 19312
rect 30600 19252 30812 19312
rect 31144 19312 32716 19388
rect 31144 19252 31492 19312
rect 30600 19246 31492 19252
rect 30600 19182 30742 19246
rect 30806 19182 31492 19246
rect 30600 19176 31492 19182
rect 31824 19176 32036 19312
rect 32504 19252 32716 19312
rect 33048 19252 33260 19388
rect 32504 19246 33260 19252
rect 32504 19182 32510 19246
rect 32574 19182 33190 19246
rect 33254 19182 33260 19246
rect 32504 19176 33260 19182
rect 33728 19312 34620 19388
rect 33728 19246 33940 19312
rect 33728 19182 33734 19246
rect 33798 19182 33940 19246
rect 33728 19176 33940 19182
rect 34272 19252 34620 19312
rect 34952 19252 35164 19388
rect 35632 19312 37748 19388
rect 35632 19252 35844 19312
rect 34272 19246 35844 19252
rect 34272 19182 34550 19246
rect 34614 19182 35638 19246
rect 35702 19182 35844 19246
rect 34272 19176 35844 19182
rect 36176 19176 36388 19312
rect 36856 19252 37068 19312
rect 37400 19252 37748 19312
rect 38080 19252 38292 19388
rect 36856 19246 37340 19252
rect 36856 19182 37270 19246
rect 37334 19182 37340 19246
rect 36856 19176 37340 19182
rect 37400 19246 38292 19252
rect 37400 19182 38222 19246
rect 38286 19182 38292 19246
rect 37400 19176 38292 19182
rect 38760 19252 38972 19388
rect 39304 19252 39516 19388
rect 38760 19246 39516 19252
rect 38760 19182 38766 19246
rect 38830 19182 39446 19246
rect 39510 19182 39516 19246
rect 38760 19176 39516 19182
rect 39984 19312 40740 19388
rect 39984 19246 40196 19312
rect 39984 19182 39990 19246
rect 40054 19182 40196 19246
rect 39984 19176 40196 19182
rect 40528 19246 40740 19312
rect 40528 19182 40670 19246
rect 40734 19182 40740 19246
rect 40528 19176 40740 19182
rect 41208 19252 41420 19388
rect 41752 19252 42100 19388
rect 41208 19246 42100 19252
rect 41208 19182 41214 19246
rect 41278 19182 42030 19246
rect 42094 19182 42100 19246
rect 41208 19176 42100 19182
rect 42432 19312 43324 19388
rect 42432 19246 42644 19312
rect 42432 19182 42438 19246
rect 42502 19182 42644 19246
rect 42432 19176 42644 19182
rect 43112 19246 43324 19312
rect 43656 19252 43868 19388
rect 44336 19312 45228 19388
rect 44336 19252 44548 19312
rect 43422 19246 44548 19252
rect 43112 19182 43254 19246
rect 43318 19182 43324 19246
rect 43384 19182 43390 19246
rect 43454 19182 44478 19246
rect 44542 19182 44548 19246
rect 43112 19176 43324 19182
rect 43422 19176 44548 19182
rect 44880 19252 45228 19312
rect 45560 19252 45772 19388
rect 46240 19312 46996 19388
rect 46240 19252 46452 19312
rect 44880 19246 46452 19252
rect 44880 19182 45702 19246
rect 45766 19182 46452 19246
rect 44880 19176 46452 19182
rect 46784 19246 46996 19312
rect 46784 19182 46926 19246
rect 46990 19182 46996 19246
rect 46784 19176 46996 19182
rect 47464 19252 47676 19388
rect 48008 19252 48356 19388
rect 48688 19312 49580 19388
rect 48688 19252 48900 19312
rect 47464 19246 48900 19252
rect 47464 19182 47470 19246
rect 47534 19182 48150 19246
rect 48214 19182 48900 19246
rect 47464 19176 48900 19182
rect 49368 19252 49580 19312
rect 49912 19252 50124 19388
rect 50592 19312 52028 19388
rect 50592 19252 50804 19312
rect 49368 19246 50804 19252
rect 49368 19182 49918 19246
rect 49982 19182 50804 19246
rect 49368 19176 50804 19182
rect 51136 19246 51348 19312
rect 51136 19182 51278 19246
rect 51342 19182 51348 19246
rect 51136 19176 51348 19182
rect 51816 19252 52028 19312
rect 52360 19252 52708 19388
rect 53040 19252 53252 19388
rect 51816 19246 53252 19252
rect 51816 19182 51958 19246
rect 52022 19182 53182 19246
rect 53246 19182 53252 19246
rect 51816 19176 53252 19182
rect 53720 19252 53932 19388
rect 54264 19252 54476 19388
rect 53720 19246 54476 19252
rect 53720 19182 53726 19246
rect 53790 19182 54406 19246
rect 54470 19182 54476 19246
rect 53720 19176 54476 19182
rect 54944 19312 55836 19388
rect 54944 19246 55156 19312
rect 54944 19182 54950 19246
rect 55014 19182 55156 19246
rect 54944 19176 55156 19182
rect 55488 19246 55836 19312
rect 55488 19182 55630 19246
rect 55694 19182 55836 19246
rect 55488 19176 55836 19182
rect 56168 19252 56380 19388
rect 56848 19312 58284 19388
rect 56848 19252 57060 19312
rect 56168 19246 57060 19252
rect 56168 19182 56174 19246
rect 56238 19182 57060 19246
rect 56168 19176 57060 19182
rect 57392 19246 57604 19312
rect 57392 19182 57398 19246
rect 57462 19182 57604 19246
rect 57392 19176 57604 19182
rect 58072 19252 58284 19312
rect 58616 19312 59508 19388
rect 58616 19252 58964 19312
rect 58072 19246 58964 19252
rect 58072 19182 58214 19246
rect 58278 19182 58964 19246
rect 58072 19176 58964 19182
rect 59296 19246 59508 19312
rect 59296 19182 59438 19246
rect 59502 19182 59508 19246
rect 59296 19176 59508 19182
rect 59976 19252 60188 19388
rect 60520 19252 60732 19388
rect 61200 19312 61956 19388
rect 61200 19252 61412 19312
rect 59976 19246 60732 19252
rect 60830 19246 61412 19252
rect 59976 19182 59982 19246
rect 60046 19182 60662 19246
rect 60726 19182 60732 19246
rect 60792 19182 60798 19246
rect 60862 19182 61412 19246
rect 59976 19176 60732 19182
rect 60830 19176 61412 19182
rect 61744 19246 61956 19312
rect 61744 19182 61886 19246
rect 61950 19182 61956 19246
rect 61744 19176 61956 19182
rect 62424 19252 62636 19388
rect 62968 19312 64540 19388
rect 62968 19252 63316 19312
rect 62424 19246 63316 19252
rect 62424 19182 62430 19246
rect 62494 19182 63110 19246
rect 63174 19182 63316 19246
rect 62424 19176 63316 19182
rect 63648 19176 63860 19312
rect 64328 19252 64540 19312
rect 64872 19252 65084 19388
rect 65552 19312 66444 19388
rect 65552 19252 65764 19312
rect 64328 19246 65764 19252
rect 64328 19182 64470 19246
rect 64534 19182 65764 19246
rect 64328 19176 65764 19182
rect 66096 19246 66444 19312
rect 66096 19182 66238 19246
rect 66302 19182 66444 19246
rect 66096 19176 66444 19182
rect 66776 19246 66988 19388
rect 66776 19182 66918 19246
rect 66982 19182 66988 19246
rect 66776 19176 66988 19182
rect 67456 19312 68892 19388
rect 67456 19246 67668 19312
rect 67456 19182 67462 19246
rect 67526 19182 67668 19246
rect 67456 19176 67668 19182
rect 68000 19176 68212 19312
rect 68680 19252 68892 19312
rect 69224 19252 69572 19388
rect 69904 19312 71340 19388
rect 69904 19252 70116 19312
rect 68680 19246 70116 19252
rect 68680 19182 68686 19246
rect 68750 19182 69366 19246
rect 69430 19182 70116 19246
rect 68680 19176 70116 19182
rect 70584 19252 70796 19312
rect 71128 19252 71340 19312
rect 71808 19252 72020 19388
rect 70584 19246 71068 19252
rect 70584 19182 70998 19246
rect 71062 19182 71068 19246
rect 70584 19176 71068 19182
rect 71128 19246 72020 19252
rect 71128 19182 71950 19246
rect 72014 19182 72020 19246
rect 71128 19176 72020 19182
rect 72352 19312 73244 19388
rect 72352 19246 72564 19312
rect 72352 19182 72358 19246
rect 72422 19182 72564 19246
rect 72352 19176 72564 19182
rect 73032 19252 73244 19312
rect 73576 19252 73924 19388
rect 74256 19312 75148 19388
rect 74256 19252 74468 19312
rect 73032 19246 74468 19252
rect 73032 19182 73174 19246
rect 73238 19182 74468 19246
rect 73032 19176 74468 19182
rect 74936 19252 75148 19312
rect 75480 19252 75692 19388
rect 74936 19246 75692 19252
rect 74936 19182 74942 19246
rect 75006 19182 75622 19246
rect 75686 19182 75692 19246
rect 74936 19176 75692 19182
rect 76160 19312 77596 19388
rect 76160 19246 76372 19312
rect 76160 19182 76166 19246
rect 76230 19182 76372 19246
rect 76160 19176 76372 19182
rect 76704 19176 77052 19312
rect 77384 19252 77596 19312
rect 78064 19312 80724 19388
rect 78064 19252 78276 19312
rect 77384 19246 78276 19252
rect 77384 19182 77390 19246
rect 77454 19182 78070 19246
rect 78134 19182 78276 19246
rect 77384 19176 78276 19182
rect 78608 19176 78820 19312
rect 79288 19252 79500 19312
rect 79288 19246 79772 19252
rect 79288 19182 79702 19246
rect 79766 19182 79772 19246
rect 79288 19176 79772 19182
rect 79832 19176 80180 19312
rect 80512 19246 80724 19312
rect 80512 19182 80654 19246
rect 80718 19182 80724 19246
rect 80512 19176 80724 19182
rect 81192 19252 81404 19388
rect 81736 19252 81948 19388
rect 82416 19312 83852 19388
rect 82416 19252 82628 19312
rect 81192 19246 82628 19252
rect 81192 19182 81198 19246
rect 81262 19182 81878 19246
rect 81942 19182 82628 19246
rect 81192 19176 82628 19182
rect 82960 19176 83172 19312
rect 83640 19252 83852 19312
rect 84184 19252 84532 19388
rect 83640 19246 84532 19252
rect 83640 19182 83646 19246
rect 83710 19182 84326 19246
rect 84390 19182 84532 19246
rect 83640 19176 84532 19182
rect 84864 19312 85756 19388
rect 84864 19246 85076 19312
rect 84864 19182 84870 19246
rect 84934 19182 85076 19246
rect 84864 19176 85076 19182
rect 85544 19252 85756 19312
rect 86088 19252 86300 19388
rect 86768 19252 86980 19388
rect 85544 19246 86980 19252
rect 85544 19182 86094 19246
rect 86158 19182 86910 19246
rect 86974 19182 86980 19246
rect 85544 19176 86980 19182
rect 87312 19312 88204 19388
rect 87312 19246 87660 19312
rect 87312 19182 87318 19246
rect 87382 19182 87660 19246
rect 87312 19176 87660 19182
rect 87992 19246 88204 19312
rect 88672 19312 89428 19388
rect 88672 19252 88884 19312
rect 88302 19246 88884 19252
rect 87992 19182 88134 19246
rect 88198 19182 88204 19246
rect 88264 19182 88270 19246
rect 88334 19182 88884 19246
rect 87992 19176 88204 19182
rect 88302 19176 88884 19182
rect 89216 19246 89428 19312
rect 89216 19182 89358 19246
rect 89422 19182 89428 19246
rect 89216 19176 89428 19182
rect 89896 19252 90108 19388
rect 90440 19252 90788 19388
rect 91120 19312 92012 19388
rect 91120 19252 91332 19312
rect 89896 19246 91332 19252
rect 89896 19182 89902 19246
rect 89966 19182 90718 19246
rect 90782 19182 91332 19246
rect 89896 19176 91332 19182
rect 91800 19246 92012 19312
rect 91800 19182 91806 19246
rect 91870 19182 92012 19246
rect 91800 19176 92012 19182
rect 92344 19252 92556 19388
rect 93024 19312 94460 19388
rect 94558 19382 95140 19388
rect 94520 19318 94526 19382
rect 94590 19318 95140 19382
rect 94558 19312 95140 19318
rect 93024 19252 93236 19312
rect 92344 19246 93508 19252
rect 92344 19182 92350 19246
rect 92414 19182 93438 19246
rect 93502 19182 93508 19246
rect 92344 19176 93508 19182
rect 93568 19176 93780 19312
rect 94248 19252 94460 19312
rect 94792 19252 95140 19312
rect 95472 19252 95684 19388
rect 94248 19246 95684 19252
rect 94248 19182 95614 19246
rect 95678 19182 95684 19246
rect 94248 19176 95684 19182
rect 96152 19252 96364 19388
rect 96696 19252 96908 19388
rect 97376 19312 98268 19388
rect 97376 19252 97588 19312
rect 96152 19246 97588 19252
rect 96152 19182 96158 19246
rect 96222 19182 96838 19246
rect 96902 19182 97588 19246
rect 96152 19176 97588 19182
rect 97920 19246 98268 19312
rect 97920 19182 98198 19246
rect 98262 19182 98268 19246
rect 97920 19176 98268 19182
rect 98600 19252 98812 19388
rect 99280 19312 100716 19388
rect 99280 19252 99492 19312
rect 98600 19246 99492 19252
rect 98600 19182 98606 19246
rect 98670 19182 99492 19246
rect 98600 19176 99492 19182
rect 99824 19246 100036 19312
rect 99824 19182 99830 19246
rect 99894 19182 100036 19246
rect 99824 19176 100036 19182
rect 100504 19252 100716 19312
rect 101048 19252 101396 19388
rect 101728 19252 101940 19388
rect 100504 19246 101940 19252
rect 100504 19182 101190 19246
rect 101254 19182 101870 19246
rect 101934 19182 101940 19246
rect 100504 19176 101940 19182
rect 102408 19252 102620 19388
rect 102952 19252 103164 19388
rect 103632 19312 104388 19388
rect 103632 19252 103844 19312
rect 102408 19246 103844 19252
rect 102408 19182 102414 19246
rect 102478 19182 103094 19246
rect 103158 19182 103844 19246
rect 102408 19176 103844 19182
rect 104176 19246 104388 19312
rect 104176 19182 104318 19246
rect 104382 19182 104388 19246
rect 104176 19176 104388 19182
rect 104856 19252 105068 19388
rect 105400 19252 105748 19388
rect 106080 19312 106972 19388
rect 106080 19252 106292 19312
rect 104856 19246 105748 19252
rect 105846 19246 106292 19252
rect 104856 19182 104862 19246
rect 104926 19182 105542 19246
rect 105606 19182 105748 19246
rect 105808 19182 105814 19246
rect 105878 19182 106292 19246
rect 104856 19176 105748 19182
rect 105846 19176 106292 19182
rect 106760 19252 106972 19312
rect 107304 19252 107516 19388
rect 107984 19312 108876 19388
rect 107984 19252 108196 19312
rect 106760 19246 107244 19252
rect 106760 19182 107174 19246
rect 107238 19182 107244 19246
rect 106760 19176 107244 19182
rect 107304 19246 108196 19252
rect 107304 19182 107310 19246
rect 107374 19182 108196 19246
rect 107304 19176 108196 19182
rect 108528 19246 108876 19312
rect 108528 19182 108534 19246
rect 108598 19182 108876 19246
rect 123216 19312 136620 19388
rect 123216 19310 123428 19312
rect 123216 19254 123270 19310
rect 123326 19254 123428 19310
rect 108528 19176 108876 19182
rect 121982 19241 122048 19244
rect 122320 19241 122386 19244
rect 121982 19239 122386 19241
rect 121982 19183 121987 19239
rect 122043 19183 122325 19239
rect 122381 19183 122386 19239
rect 121982 19181 122386 19183
rect 121982 19178 122048 19181
rect 122320 19178 122386 19181
rect 123216 19176 123428 19254
rect 3128 19040 4156 19116
rect 1768 18888 1980 18980
rect 1768 18844 1794 18888
rect 1224 18838 1794 18844
rect 1224 18774 1230 18838
rect 1294 18832 1794 18838
rect 1850 18844 1980 18888
rect 3128 18844 3340 19040
rect 1850 18832 3340 18844
rect 1294 18774 3340 18832
rect 1224 18768 3340 18774
rect 3944 18768 4156 19040
rect 14552 19110 16668 19116
rect 14552 19046 16598 19110
rect 16662 19046 16668 19110
rect 14552 19040 16668 19046
rect 14552 18838 14764 19040
rect 134776 18974 135396 18980
rect 134776 18910 135326 18974
rect 135390 18910 135396 18974
rect 134776 18904 135396 18910
rect 134776 18888 134988 18904
rect 14552 18774 14694 18838
rect 14758 18774 14764 18838
rect 14552 18768 14764 18774
rect 28152 18838 28500 18844
rect 28152 18774 28294 18838
rect 28358 18774 28500 18838
rect 28152 18632 28500 18774
rect 28560 18838 28772 18844
rect 28560 18774 28566 18838
rect 28630 18774 28772 18838
rect 28560 18632 28772 18774
rect 29512 18838 29724 18844
rect 29512 18774 29518 18838
rect 29582 18774 29724 18838
rect 29512 18708 29724 18774
rect 29784 18708 30132 18844
rect 29512 18632 30132 18708
rect 30736 18838 31356 18844
rect 30736 18774 30742 18838
rect 30806 18774 31356 18838
rect 30736 18768 31356 18774
rect 30736 18632 30948 18768
rect 31144 18632 31356 18768
rect 31960 18708 32172 18844
rect 32368 18838 32580 18844
rect 32368 18774 32510 18838
rect 32574 18774 32580 18838
rect 32368 18708 32580 18774
rect 31960 18632 32580 18708
rect 33184 18838 33804 18844
rect 33184 18774 33190 18838
rect 33254 18774 33734 18838
rect 33798 18774 33804 18838
rect 33184 18768 33804 18774
rect 33184 18632 33396 18768
rect 33592 18632 33804 18768
rect 34408 18838 34620 18844
rect 34408 18774 34550 18838
rect 34614 18774 34620 18838
rect 34408 18708 34620 18774
rect 34816 18708 35028 18844
rect 34408 18632 35028 18708
rect 35632 18838 36252 18844
rect 35632 18774 35638 18838
rect 35702 18774 36252 18838
rect 35632 18768 36252 18774
rect 35632 18632 35980 18768
rect 36040 18632 36252 18768
rect 36992 18838 37612 18844
rect 36992 18774 37270 18838
rect 37334 18774 37612 18838
rect 36992 18768 37612 18774
rect 36992 18632 37204 18768
rect 37264 18632 37612 18768
rect 38216 18838 38428 18844
rect 38216 18774 38222 18838
rect 38286 18774 38428 18838
rect 38216 18708 38428 18774
rect 38624 18838 38836 18844
rect 38624 18774 38766 18838
rect 38830 18774 38836 18838
rect 38624 18708 38836 18774
rect 38216 18632 38836 18708
rect 39440 18838 40060 18844
rect 39440 18774 39446 18838
rect 39510 18774 39990 18838
rect 40054 18774 40060 18838
rect 39440 18768 40060 18774
rect 39440 18632 39652 18768
rect 39848 18632 40060 18768
rect 40664 18838 40876 18844
rect 40664 18774 40670 18838
rect 40734 18774 40876 18838
rect 40664 18708 40876 18774
rect 41072 18838 41284 18844
rect 41072 18774 41214 18838
rect 41278 18774 41284 18838
rect 41072 18708 41284 18774
rect 40664 18632 41284 18708
rect 41888 18838 42508 18844
rect 41888 18774 42030 18838
rect 42094 18774 42438 18838
rect 42502 18774 42508 18838
rect 41888 18768 42508 18774
rect 41888 18632 42236 18768
rect 42296 18632 42508 18768
rect 43248 18838 43868 18844
rect 43248 18774 43254 18838
rect 43318 18774 43390 18838
rect 43454 18774 43868 18838
rect 43248 18768 43868 18774
rect 43248 18632 43460 18768
rect 43520 18632 43868 18768
rect 44472 18838 44684 18844
rect 44472 18774 44478 18838
rect 44542 18774 44684 18838
rect 44472 18708 44684 18774
rect 44880 18708 45092 18844
rect 44472 18632 45092 18708
rect 45696 18838 46316 18844
rect 45696 18774 45702 18838
rect 45766 18774 46316 18838
rect 45696 18768 46316 18774
rect 45696 18632 45908 18768
rect 46104 18632 46316 18768
rect 46920 18838 47132 18844
rect 46920 18774 46926 18838
rect 46990 18774 47132 18838
rect 46920 18708 47132 18774
rect 47328 18838 47540 18844
rect 47328 18774 47470 18838
rect 47534 18774 47540 18838
rect 47328 18708 47540 18774
rect 46920 18632 47540 18708
rect 48144 18838 48764 18844
rect 48144 18774 48150 18838
rect 48214 18774 48764 18838
rect 48144 18768 48764 18774
rect 48144 18632 48356 18768
rect 48552 18632 48764 18768
rect 49368 18708 49716 18844
rect 49776 18838 49988 18844
rect 49776 18774 49918 18838
rect 49982 18774 49988 18838
rect 49776 18708 49988 18774
rect 49368 18632 49988 18708
rect 50728 18708 50940 18844
rect 51000 18838 51348 18844
rect 51000 18774 51278 18838
rect 51342 18774 51348 18838
rect 51000 18708 51348 18774
rect 50728 18632 51348 18708
rect 51952 18838 52572 18844
rect 51952 18774 51958 18838
rect 52022 18774 52572 18838
rect 51952 18768 52572 18774
rect 51952 18632 52164 18768
rect 52360 18632 52572 18768
rect 53176 18838 53388 18844
rect 53176 18774 53182 18838
rect 53246 18774 53388 18838
rect 53176 18708 53388 18774
rect 53584 18838 53796 18844
rect 53584 18774 53726 18838
rect 53790 18774 53796 18838
rect 53584 18708 53796 18774
rect 53176 18632 53796 18708
rect 54400 18838 55020 18844
rect 54400 18774 54406 18838
rect 54470 18774 54950 18838
rect 55014 18774 55020 18838
rect 54400 18768 55020 18774
rect 54400 18632 54612 18768
rect 54808 18632 55020 18768
rect 55624 18838 55836 18844
rect 55624 18774 55630 18838
rect 55694 18774 55836 18838
rect 55624 18708 55836 18774
rect 56032 18838 56244 18844
rect 56032 18774 56174 18838
rect 56238 18774 56244 18838
rect 56032 18708 56244 18774
rect 55624 18632 56244 18708
rect 56848 18838 57468 18844
rect 56848 18774 57398 18838
rect 57462 18774 57468 18838
rect 56848 18768 57468 18774
rect 56848 18632 57196 18768
rect 57256 18632 57468 18768
rect 58208 18838 58828 18844
rect 58208 18774 58214 18838
rect 58278 18774 58828 18838
rect 58208 18768 58828 18774
rect 58208 18702 58420 18768
rect 58208 18638 58350 18702
rect 58414 18638 58420 18702
rect 58208 18632 58420 18638
rect 58480 18632 58828 18768
rect 59432 18838 59644 18844
rect 59432 18774 59438 18838
rect 59502 18774 59644 18838
rect 59432 18708 59644 18774
rect 59840 18838 60052 18844
rect 59840 18774 59982 18838
rect 60046 18774 60052 18838
rect 59840 18708 60052 18774
rect 59432 18632 60052 18708
rect 60656 18838 61276 18844
rect 60656 18774 60662 18838
rect 60726 18774 60798 18838
rect 60862 18774 61276 18838
rect 60656 18768 61276 18774
rect 60656 18632 60868 18768
rect 61064 18632 61276 18768
rect 61880 18838 62092 18844
rect 61880 18774 61886 18838
rect 61950 18774 62092 18838
rect 61880 18708 62092 18774
rect 62288 18838 62500 18844
rect 62288 18774 62430 18838
rect 62494 18774 62500 18838
rect 62288 18708 62500 18774
rect 61880 18632 62500 18708
rect 63104 18838 63452 18844
rect 63104 18774 63110 18838
rect 63174 18774 63452 18838
rect 63104 18708 63452 18774
rect 63512 18708 63724 18844
rect 63104 18632 63724 18708
rect 64464 18838 65084 18844
rect 64464 18774 64470 18838
rect 64534 18774 65084 18838
rect 64464 18768 65084 18774
rect 64464 18632 64676 18768
rect 64736 18632 65084 18768
rect 65688 18708 65900 18844
rect 66096 18838 67532 18844
rect 66096 18774 66238 18838
rect 66302 18774 66918 18838
rect 66982 18774 67462 18838
rect 67526 18774 67532 18838
rect 66096 18768 67532 18774
rect 66096 18708 66308 18768
rect 65688 18632 66308 18708
rect 66912 18632 67124 18768
rect 67320 18632 67532 18768
rect 68136 18708 68348 18844
rect 68544 18838 68756 18844
rect 68544 18774 68686 18838
rect 68750 18774 68756 18838
rect 68544 18708 68756 18774
rect 68136 18632 68756 18708
rect 69360 18838 69980 18844
rect 69360 18774 69366 18838
rect 69430 18774 69980 18838
rect 69360 18768 69980 18774
rect 69360 18632 69572 18768
rect 69768 18632 69980 18768
rect 70584 18708 70932 18844
rect 70992 18838 71204 18844
rect 70992 18774 70998 18838
rect 71062 18774 71204 18838
rect 70992 18708 71204 18774
rect 70584 18632 71204 18708
rect 71944 18838 72156 18844
rect 71944 18774 71950 18838
rect 72014 18774 72156 18838
rect 71944 18708 72156 18774
rect 72216 18838 72564 18844
rect 72216 18774 72358 18838
rect 72422 18774 72564 18838
rect 72216 18708 72564 18774
rect 71944 18632 72564 18708
rect 73168 18838 73788 18844
rect 73168 18774 73174 18838
rect 73238 18774 73788 18838
rect 73168 18768 73788 18774
rect 73168 18632 73380 18768
rect 73576 18632 73788 18768
rect 74392 18708 74604 18844
rect 74800 18838 75012 18844
rect 74800 18774 74942 18838
rect 75006 18774 75012 18838
rect 74800 18708 75012 18774
rect 74392 18632 75012 18708
rect 75616 18838 76236 18844
rect 75616 18774 75622 18838
rect 75686 18774 76166 18838
rect 76230 18774 76236 18838
rect 75616 18768 76236 18774
rect 75616 18632 75828 18768
rect 76024 18632 76236 18768
rect 76840 18708 77052 18844
rect 77248 18838 77460 18844
rect 77248 18774 77390 18838
rect 77454 18774 77460 18838
rect 77248 18708 77460 18774
rect 76840 18632 77460 18708
rect 78064 18838 78684 18844
rect 78064 18774 78070 18838
rect 78134 18774 78684 18838
rect 78064 18768 78684 18774
rect 78064 18632 78412 18768
rect 78472 18632 78684 18768
rect 79424 18838 80044 18844
rect 79424 18774 79702 18838
rect 79766 18774 80044 18838
rect 79424 18768 80044 18774
rect 79424 18632 79636 18768
rect 79696 18632 80044 18768
rect 80648 18838 80860 18844
rect 80648 18774 80654 18838
rect 80718 18774 80860 18838
rect 80648 18708 80860 18774
rect 81056 18838 81268 18844
rect 81056 18774 81198 18838
rect 81262 18774 81268 18838
rect 81056 18708 81268 18774
rect 80648 18632 81268 18708
rect 81872 18838 82492 18844
rect 81872 18774 81878 18838
rect 81942 18774 82492 18838
rect 81872 18768 82492 18774
rect 81872 18632 82084 18768
rect 82280 18632 82492 18768
rect 83096 18708 83308 18844
rect 83504 18838 83716 18844
rect 83504 18774 83646 18838
rect 83710 18774 83716 18838
rect 83504 18708 83716 18774
rect 83096 18632 83716 18708
rect 84320 18838 84668 18844
rect 84320 18774 84326 18838
rect 84390 18774 84668 18838
rect 84320 18708 84668 18774
rect 84728 18838 84940 18844
rect 84728 18774 84870 18838
rect 84934 18774 84940 18838
rect 84728 18708 84940 18774
rect 84320 18632 84940 18708
rect 85680 18838 86300 18844
rect 85680 18774 86094 18838
rect 86158 18774 86300 18838
rect 85680 18768 86300 18774
rect 85680 18632 85892 18768
rect 85952 18632 86300 18768
rect 86904 18838 87116 18844
rect 86904 18774 86910 18838
rect 86974 18774 87116 18838
rect 86904 18708 87116 18774
rect 87312 18838 87524 18844
rect 87312 18774 87318 18838
rect 87382 18774 87524 18838
rect 87312 18708 87524 18774
rect 86904 18632 87524 18708
rect 88128 18838 88748 18844
rect 88128 18774 88134 18838
rect 88198 18774 88270 18838
rect 88334 18774 88748 18838
rect 88128 18768 88748 18774
rect 88128 18632 88340 18768
rect 88536 18632 88748 18768
rect 89352 18838 89564 18844
rect 89352 18774 89358 18838
rect 89422 18774 89564 18838
rect 89352 18708 89564 18774
rect 89760 18838 89972 18844
rect 89760 18774 89902 18838
rect 89966 18774 89972 18838
rect 89760 18708 89972 18774
rect 89352 18632 89972 18708
rect 90576 18838 91196 18844
rect 90576 18774 90718 18838
rect 90782 18774 91196 18838
rect 90576 18768 91196 18774
rect 90576 18632 90788 18768
rect 90984 18632 91196 18768
rect 91800 18838 92148 18844
rect 91800 18774 91806 18838
rect 91870 18774 92148 18838
rect 91800 18708 92148 18774
rect 92208 18838 92420 18844
rect 92208 18774 92350 18838
rect 92414 18774 92420 18838
rect 92208 18708 92420 18774
rect 91800 18632 92420 18708
rect 93160 18708 93372 18844
rect 93432 18838 93780 18844
rect 93432 18774 93438 18838
rect 93502 18774 93780 18838
rect 93432 18708 93780 18774
rect 93160 18632 93780 18708
rect 94384 18838 95004 18844
rect 94384 18774 94526 18838
rect 94590 18774 95004 18838
rect 94384 18768 95004 18774
rect 94384 18632 94596 18768
rect 94792 18632 95004 18768
rect 95608 18838 95820 18844
rect 95608 18774 95614 18838
rect 95678 18774 95820 18838
rect 95608 18708 95820 18774
rect 96016 18838 96228 18844
rect 96016 18774 96158 18838
rect 96222 18774 96228 18838
rect 96016 18708 96228 18774
rect 95608 18632 96228 18708
rect 96832 18838 97452 18844
rect 96832 18774 96838 18838
rect 96902 18774 97452 18838
rect 96832 18768 97452 18774
rect 96832 18632 97044 18768
rect 97240 18632 97452 18768
rect 98056 18838 98268 18844
rect 98056 18774 98198 18838
rect 98262 18774 98268 18838
rect 98056 18708 98268 18774
rect 98464 18838 98676 18844
rect 98464 18774 98606 18838
rect 98670 18774 98676 18838
rect 98464 18708 98676 18774
rect 98056 18632 98676 18708
rect 99280 18708 99628 18844
rect 99688 18838 99900 18844
rect 99688 18774 99830 18838
rect 99894 18774 99900 18838
rect 99688 18708 99900 18774
rect 99280 18632 99900 18708
rect 100640 18838 101260 18844
rect 100640 18774 101190 18838
rect 101254 18774 101260 18838
rect 100640 18768 101260 18774
rect 100640 18632 100852 18768
rect 100912 18632 101260 18768
rect 101864 18838 102076 18844
rect 101864 18774 101870 18838
rect 101934 18774 102076 18838
rect 101864 18708 102076 18774
rect 102272 18838 102484 18844
rect 102272 18774 102414 18838
rect 102478 18774 102484 18838
rect 102272 18708 102484 18774
rect 101864 18632 102484 18708
rect 103088 18838 103708 18844
rect 103088 18774 103094 18838
rect 103158 18774 103708 18838
rect 103088 18768 103708 18774
rect 103088 18632 103300 18768
rect 103496 18632 103708 18768
rect 104312 18838 104524 18844
rect 104312 18774 104318 18838
rect 104382 18774 104524 18838
rect 104312 18708 104524 18774
rect 104720 18838 104932 18844
rect 104720 18774 104862 18838
rect 104926 18774 104932 18838
rect 104720 18708 104932 18774
rect 104312 18632 104932 18708
rect 105536 18838 106156 18844
rect 105536 18774 105542 18838
rect 105606 18774 105814 18838
rect 105878 18774 106156 18838
rect 105536 18768 106156 18774
rect 105536 18632 105884 18768
rect 105944 18632 106156 18768
rect 106896 18838 107516 18844
rect 106896 18774 107174 18838
rect 107238 18774 107310 18838
rect 107374 18774 107516 18838
rect 106896 18768 107516 18774
rect 106896 18632 107108 18768
rect 107168 18632 107516 18768
rect 108120 18838 108604 18844
rect 108120 18774 108534 18838
rect 108598 18774 108604 18838
rect 108120 18768 108604 18774
rect 134776 18832 134844 18888
rect 134900 18832 134988 18888
rect 134776 18768 134988 18832
rect 108120 18632 108332 18768
rect 119990 18566 123020 18572
rect 119952 18502 119958 18566
rect 120022 18502 123020 18566
rect 119990 18496 123020 18502
rect 122808 18430 123020 18496
rect 122808 18366 122950 18430
rect 123014 18366 123020 18430
rect 122808 18360 123020 18366
rect 14661 18255 14727 18258
rect 22803 18255 22869 18258
rect 14661 18253 22869 18255
rect 14661 18197 14666 18253
rect 14722 18197 22808 18253
rect 22864 18197 22869 18253
rect 14661 18195 22869 18197
rect 14661 18192 14727 18195
rect 22803 18192 22869 18195
rect 2531 17894 2537 17958
rect 2601 17956 2607 17958
rect 2601 17896 28439 17956
rect 2601 17894 2607 17896
rect 121902 17683 121968 17686
rect 122320 17683 122386 17686
rect 121902 17681 122386 17683
rect 121902 17625 121907 17681
rect 121963 17625 122325 17681
rect 122381 17625 122386 17681
rect 121902 17623 122386 17625
rect 121902 17620 121968 17623
rect 122320 17620 122386 17623
rect 123216 17680 136620 17756
rect 3128 17484 3340 17620
rect 3710 17614 4156 17620
rect 3672 17550 3678 17614
rect 3742 17550 4156 17614
rect 3710 17544 4156 17550
rect 3944 17484 4156 17544
rect 3128 17408 4156 17484
rect 14552 17614 17076 17620
rect 14552 17550 17006 17614
rect 17070 17550 17076 17614
rect 14552 17544 17076 17550
rect 123216 17610 123428 17680
rect 123216 17554 123270 17610
rect 123326 17554 123428 17610
rect 14552 17478 14764 17544
rect 14552 17414 14558 17478
rect 14622 17414 14764 17478
rect 14552 17408 14764 17414
rect 123216 17408 123428 17554
rect 1768 17208 1980 17348
rect 1768 17152 1794 17208
rect 1850 17152 1980 17208
rect 1768 17076 1980 17152
rect 20128 17342 21564 17348
rect 20128 17278 21222 17342
rect 21286 17278 21564 17342
rect 20128 17272 21564 17278
rect 20128 17136 20340 17272
rect 21216 17206 21564 17272
rect 134776 17212 134988 17348
rect 21216 17142 21358 17206
rect 21422 17142 21564 17206
rect 21216 17136 21564 17142
rect 28968 17206 30540 17212
rect 28968 17142 28974 17206
rect 29038 17142 30540 17206
rect 28968 17136 30540 17142
rect 1224 17070 1980 17076
rect 1224 17006 1230 17070
rect 1294 17006 1980 17070
rect 1224 17000 1980 17006
rect 28968 17070 29316 17136
rect 28968 17006 28974 17070
rect 29038 17006 29316 17070
rect 28968 17000 29316 17006
rect 30328 17076 30540 17136
rect 31552 17136 32988 17212
rect 31552 17076 31764 17136
rect 30328 17070 31764 17076
rect 30328 17006 31694 17070
rect 31758 17006 31764 17070
rect 30328 17000 31764 17006
rect 32776 17076 32988 17136
rect 34000 17136 35436 17212
rect 34000 17076 34212 17136
rect 32776 17070 34212 17076
rect 32776 17006 34006 17070
rect 34070 17006 34212 17070
rect 32776 17000 34212 17006
rect 35224 17076 35436 17136
rect 36448 17076 36796 17212
rect 37808 17136 39244 17212
rect 37808 17076 38020 17136
rect 35224 17070 38020 17076
rect 35224 17006 36454 17070
rect 36518 17006 38020 17070
rect 35224 17000 38020 17006
rect 39032 17076 39244 17136
rect 40256 17136 41692 17212
rect 40256 17076 40468 17136
rect 39032 17070 40468 17076
rect 39032 17006 39174 17070
rect 39238 17006 40468 17070
rect 39032 17000 40468 17006
rect 41480 17076 41692 17136
rect 42704 17076 43052 17212
rect 44064 17136 45500 17212
rect 44064 17076 44276 17136
rect 41480 17070 44276 17076
rect 41480 17006 41622 17070
rect 41686 17006 44070 17070
rect 44134 17006 44276 17070
rect 41480 17000 44276 17006
rect 45288 17076 45500 17136
rect 46512 17136 47948 17212
rect 46512 17076 46724 17136
rect 45288 17070 46724 17076
rect 45288 17006 46654 17070
rect 46718 17006 46724 17070
rect 45288 17000 46724 17006
rect 47736 17076 47948 17136
rect 48960 17136 50532 17212
rect 48960 17076 49172 17136
rect 47736 17070 49172 17076
rect 47736 17006 48966 17070
rect 49030 17006 49172 17070
rect 47736 17000 49172 17006
rect 50184 17076 50532 17136
rect 51544 17076 51756 17212
rect 52768 17136 54204 17212
rect 52768 17076 52980 17136
rect 50184 17070 52980 17076
rect 50184 17006 51550 17070
rect 51614 17006 52980 17070
rect 50184 17000 52980 17006
rect 53992 17076 54204 17136
rect 55216 17136 56652 17212
rect 55216 17076 55428 17136
rect 53992 17070 55428 17076
rect 53992 17006 54134 17070
rect 54198 17006 55428 17070
rect 53992 17000 55428 17006
rect 56440 17076 56652 17136
rect 57664 17136 60460 17212
rect 57664 17076 58012 17136
rect 56440 17070 58012 17076
rect 56440 17006 56446 17070
rect 56510 17006 58012 17070
rect 56440 17000 58012 17006
rect 59024 17070 59236 17136
rect 59024 17006 59166 17070
rect 59230 17006 59236 17070
rect 59024 17000 59236 17006
rect 60248 17076 60460 17136
rect 61472 17136 62908 17212
rect 61472 17076 61684 17136
rect 60248 17070 61684 17076
rect 60248 17006 61614 17070
rect 61678 17006 61684 17070
rect 60248 17000 61684 17006
rect 62696 17076 62908 17136
rect 63920 17076 64268 17212
rect 65280 17136 66716 17212
rect 65280 17076 65492 17136
rect 62696 17070 65492 17076
rect 62696 17006 63926 17070
rect 63990 17006 65492 17070
rect 62696 17000 65492 17006
rect 66504 17076 66716 17136
rect 67728 17136 69164 17212
rect 67728 17076 67940 17136
rect 66504 17070 67940 17076
rect 66504 17006 66646 17070
rect 66710 17006 67940 17070
rect 66504 17000 67940 17006
rect 68952 17076 69164 17136
rect 70176 17136 71748 17212
rect 70176 17076 70388 17136
rect 68952 17070 70388 17076
rect 68952 17006 69094 17070
rect 69158 17006 70388 17070
rect 68952 17000 70388 17006
rect 71400 17076 71748 17136
rect 72760 17076 72972 17212
rect 73984 17136 75420 17212
rect 73984 17076 74196 17136
rect 71400 17070 74196 17076
rect 71400 17006 71406 17070
rect 71470 17006 74126 17070
rect 74190 17006 74196 17070
rect 71400 17000 74196 17006
rect 75208 17076 75420 17136
rect 76432 17136 77868 17212
rect 76432 17076 76644 17136
rect 75208 17070 76644 17076
rect 75208 17006 76438 17070
rect 76502 17006 76644 17070
rect 75208 17000 76644 17006
rect 77656 17076 77868 17136
rect 78880 17136 81676 17212
rect 78880 17076 79228 17136
rect 77656 17070 79228 17076
rect 77656 17006 78886 17070
rect 78950 17006 79228 17070
rect 77656 17000 79228 17006
rect 80240 17000 80452 17136
rect 81464 17076 81676 17136
rect 82688 17136 84124 17212
rect 82688 17076 82900 17136
rect 81464 17070 82900 17076
rect 81464 17006 81606 17070
rect 81670 17006 82900 17070
rect 81464 17000 82900 17006
rect 83912 17076 84124 17136
rect 85136 17136 87932 17212
rect 85136 17076 85484 17136
rect 86496 17076 86708 17136
rect 83912 17070 85484 17076
rect 86398 17070 86708 17076
rect 83912 17006 83918 17070
rect 83982 17006 85484 17070
rect 86360 17006 86366 17070
rect 86430 17006 86708 17070
rect 83912 17000 85484 17006
rect 86398 17000 86708 17006
rect 87720 17076 87932 17136
rect 88944 17136 90380 17212
rect 88944 17076 89156 17136
rect 87720 17070 89156 17076
rect 87720 17006 89086 17070
rect 89150 17006 89156 17070
rect 87720 17000 89156 17006
rect 90168 17076 90380 17136
rect 91392 17136 92964 17212
rect 91392 17076 91604 17136
rect 90168 17070 91604 17076
rect 90168 17006 91398 17070
rect 91462 17006 91604 17070
rect 90168 17000 91604 17006
rect 92616 17076 92964 17136
rect 93976 17076 94188 17212
rect 95200 17136 96636 17212
rect 95200 17076 95412 17136
rect 92616 17070 95412 17076
rect 92616 17006 93982 17070
rect 94046 17006 95412 17070
rect 92616 17000 95412 17006
rect 96424 17076 96636 17136
rect 97648 17136 99084 17212
rect 97648 17076 97860 17136
rect 96424 17070 97860 17076
rect 96424 17006 96566 17070
rect 96630 17006 97860 17070
rect 96424 17000 97860 17006
rect 98872 17076 99084 17136
rect 100096 17136 102892 17212
rect 100096 17076 100444 17136
rect 98872 17070 100444 17076
rect 98872 17006 98878 17070
rect 98942 17006 100444 17070
rect 98872 17000 100444 17006
rect 101456 17070 101668 17136
rect 101456 17006 101598 17070
rect 101662 17006 101668 17070
rect 101456 17000 101668 17006
rect 102680 17076 102892 17136
rect 103904 17136 105340 17212
rect 103904 17076 104116 17136
rect 102680 17070 104116 17076
rect 102680 17006 104046 17070
rect 104110 17006 104116 17070
rect 102680 17000 104116 17006
rect 105128 17076 105340 17136
rect 106352 17136 107924 17212
rect 106352 17076 106700 17136
rect 105128 17070 106700 17076
rect 105128 17006 106358 17070
rect 106422 17006 106700 17070
rect 105128 17000 106700 17006
rect 107712 17000 107924 17136
rect 134776 17208 135396 17212
rect 134776 17152 134844 17208
rect 134900 17206 135396 17208
rect 134900 17152 135326 17206
rect 134776 17142 135326 17152
rect 135390 17142 135396 17206
rect 134776 17136 135396 17142
rect 122808 17070 123020 17076
rect 122808 17006 122814 17070
rect 122878 17006 123020 17070
rect 122808 16934 123020 17006
rect 134776 17000 134988 17136
rect 122808 16870 122814 16934
rect 122878 16870 123020 16934
rect 122808 16864 123020 16870
rect 123216 16482 123428 16532
rect 123216 16426 123270 16482
rect 123326 16426 123428 16482
rect 121822 16413 121888 16416
rect 122320 16413 122386 16416
rect 121822 16411 122386 16413
rect 121822 16355 121827 16411
rect 121883 16355 122325 16411
rect 122381 16355 122386 16411
rect 121822 16353 122386 16355
rect 121822 16350 121888 16353
rect 122320 16350 122386 16353
rect 123216 16396 123428 16426
rect 123216 16320 136620 16396
rect 3128 16184 4156 16260
rect 3128 16118 3340 16184
rect 3128 16054 3134 16118
rect 3198 16054 3340 16118
rect 3128 16048 3340 16054
rect 3944 16048 4156 16184
rect 14552 16254 14764 16260
rect 14552 16190 14694 16254
rect 14758 16190 14764 16254
rect 14552 16118 14764 16190
rect 14552 16054 14694 16118
rect 14758 16054 14764 16118
rect 14552 16048 14764 16054
rect 20128 15912 21564 15988
rect 20128 15776 20340 15912
rect 21216 15852 21564 15912
rect 21216 15846 22516 15852
rect 21216 15782 21222 15846
rect 21286 15782 22446 15846
rect 22510 15782 22516 15846
rect 21216 15776 22516 15782
rect 122808 15710 123020 15716
rect 122808 15646 122950 15710
rect 123014 15646 123020 15710
rect 1224 15574 3204 15580
rect 1224 15510 1230 15574
rect 1294 15528 3134 15574
rect 1294 15510 1794 15528
rect 1224 15504 1794 15510
rect 1768 15472 1794 15504
rect 1850 15510 3134 15528
rect 3198 15510 3204 15574
rect 1850 15504 3204 15510
rect 122808 15574 123020 15646
rect 122808 15510 122950 15574
rect 123014 15510 123020 15574
rect 122808 15504 123020 15510
rect 134776 15528 134988 15580
rect 1850 15472 1980 15504
rect 1768 15368 1980 15472
rect 134776 15472 134844 15528
rect 134900 15472 134988 15528
rect 134776 15444 134988 15472
rect 134776 15438 135396 15444
rect 14661 15427 14727 15430
rect 26506 15427 26572 15430
rect 14661 15425 26572 15427
rect 14661 15369 14666 15425
rect 14722 15369 26511 15425
rect 26567 15369 26572 15425
rect 14661 15367 26572 15369
rect 134776 15374 135326 15438
rect 135390 15374 135396 15438
rect 134776 15368 135396 15374
rect 14661 15364 14727 15367
rect 26506 15364 26572 15367
rect 28921 15172 29019 15197
rect 31417 15172 31515 15197
rect 33913 15172 34011 15197
rect 36409 15172 36507 15197
rect 38905 15172 39003 15197
rect 41401 15172 41499 15197
rect 43897 15172 43995 15197
rect 46393 15172 46491 15197
rect 48889 15172 48987 15197
rect 51385 15172 51483 15197
rect 53881 15172 53979 15197
rect 56377 15172 56475 15197
rect 58873 15172 58971 15197
rect 61369 15172 61467 15197
rect 63865 15172 63963 15197
rect 66361 15172 66459 15197
rect 68857 15172 68955 15197
rect 71353 15172 71451 15197
rect 73849 15172 73947 15197
rect 76345 15172 76443 15197
rect 78841 15172 78939 15197
rect 81337 15172 81435 15197
rect 83833 15172 83931 15197
rect 86329 15172 86427 15197
rect 88825 15172 88923 15197
rect 91321 15172 91419 15197
rect 93817 15172 93915 15197
rect 96313 15172 96411 15197
rect 98809 15172 98907 15197
rect 101305 15172 101403 15197
rect 103801 15172 103899 15197
rect 106297 15172 106395 15197
rect 28832 15166 29142 15172
rect 31416 15166 31764 15172
rect 28832 15102 28974 15166
rect 29038 15102 29110 15166
rect 29174 15102 29180 15166
rect 31416 15102 31558 15166
rect 31622 15102 31694 15166
rect 31758 15102 31764 15166
rect 28832 15096 29142 15102
rect 31416 15096 31764 15102
rect 33864 15166 34174 15172
rect 36312 15166 36622 15172
rect 38896 15166 39244 15172
rect 33864 15102 34006 15166
rect 34070 15102 34142 15166
rect 34206 15102 34212 15166
rect 36312 15102 36454 15166
rect 36518 15102 36590 15166
rect 36654 15102 36660 15166
rect 38896 15102 39038 15166
rect 39102 15102 39174 15166
rect 39238 15102 39244 15166
rect 33864 15096 34174 15102
rect 36312 15096 36622 15102
rect 38896 15096 39244 15102
rect 41344 15166 41692 15172
rect 41344 15102 41486 15166
rect 41550 15102 41622 15166
rect 41686 15102 41692 15166
rect 41344 15096 41692 15102
rect 43792 15166 44102 15172
rect 46376 15166 46724 15172
rect 43792 15102 43934 15166
rect 43998 15102 44070 15166
rect 44134 15102 44140 15166
rect 46376 15102 46518 15166
rect 46582 15102 46654 15166
rect 46718 15102 46724 15166
rect 43792 15096 44102 15102
rect 46376 15096 46724 15102
rect 48824 15166 49134 15172
rect 51272 15166 51582 15172
rect 53856 15166 54204 15172
rect 48824 15102 48966 15166
rect 49030 15102 49102 15166
rect 49166 15102 49172 15166
rect 51272 15102 51414 15166
rect 51478 15102 51550 15166
rect 51614 15102 51620 15166
rect 53856 15102 53998 15166
rect 54062 15102 54134 15166
rect 54198 15102 54204 15166
rect 48824 15096 49134 15102
rect 51272 15096 51582 15102
rect 53856 15096 54204 15102
rect 56304 15166 56614 15172
rect 58752 15166 59236 15172
rect 56304 15102 56446 15166
rect 56510 15102 56582 15166
rect 56646 15102 56652 15166
rect 58752 15102 59030 15166
rect 59094 15102 59166 15166
rect 59230 15102 59236 15166
rect 56304 15096 56614 15102
rect 58752 15096 59236 15102
rect 61336 15166 61684 15172
rect 61336 15102 61478 15166
rect 61542 15102 61614 15166
rect 61678 15102 61684 15166
rect 61336 15096 61684 15102
rect 63784 15166 64094 15172
rect 66232 15166 66716 15172
rect 63784 15102 63926 15166
rect 63990 15102 64062 15166
rect 64126 15102 64132 15166
rect 66232 15102 66510 15166
rect 66574 15102 66646 15166
rect 66710 15102 66716 15166
rect 63784 15096 64094 15102
rect 66232 15096 66716 15102
rect 68816 15166 69164 15172
rect 68816 15102 68958 15166
rect 69022 15102 69094 15166
rect 69158 15102 69164 15166
rect 68816 15096 69164 15102
rect 71264 15166 71574 15172
rect 73848 15166 74196 15172
rect 71264 15102 71406 15166
rect 71470 15102 71542 15166
rect 71606 15102 71612 15166
rect 73848 15102 73990 15166
rect 74054 15102 74126 15166
rect 74190 15102 74196 15166
rect 71264 15096 71574 15102
rect 73848 15096 74196 15102
rect 76296 15166 76606 15172
rect 78744 15166 79054 15172
rect 81328 15166 81676 15172
rect 76296 15102 76438 15166
rect 76502 15102 76574 15166
rect 76638 15102 76644 15166
rect 78744 15102 78886 15166
rect 78950 15102 79022 15166
rect 79086 15102 79092 15166
rect 81328 15102 81470 15166
rect 81534 15102 81606 15166
rect 81670 15102 81676 15166
rect 76296 15096 76606 15102
rect 78744 15096 79054 15102
rect 81328 15096 81676 15102
rect 83776 15166 84086 15172
rect 86224 15166 86534 15172
rect 88808 15166 89156 15172
rect 83776 15102 83918 15166
rect 83982 15102 84054 15166
rect 84118 15102 84124 15166
rect 86224 15102 86366 15166
rect 86430 15102 86502 15166
rect 86566 15102 86572 15166
rect 88808 15102 88950 15166
rect 89014 15102 89086 15166
rect 89150 15102 89156 15166
rect 83776 15096 84086 15102
rect 86224 15096 86534 15102
rect 88808 15096 89156 15102
rect 91256 15166 91566 15172
rect 93704 15166 94014 15172
rect 96288 15166 96636 15172
rect 91256 15102 91398 15166
rect 91462 15102 91534 15166
rect 91598 15102 91604 15166
rect 93704 15102 93846 15166
rect 93910 15102 93982 15166
rect 94046 15102 94052 15166
rect 96288 15102 96430 15166
rect 96494 15102 96566 15166
rect 96630 15102 96636 15166
rect 91256 15096 91566 15102
rect 93704 15096 94014 15102
rect 96288 15096 96636 15102
rect 98736 15166 99046 15172
rect 101184 15166 101668 15172
rect 98736 15102 98878 15166
rect 98942 15102 99014 15166
rect 99078 15102 99084 15166
rect 101184 15102 101462 15166
rect 101526 15102 101598 15166
rect 101662 15102 101668 15166
rect 98736 15096 99046 15102
rect 101184 15096 101668 15102
rect 103768 15166 104116 15172
rect 103768 15102 103910 15166
rect 103974 15102 104046 15166
rect 104110 15102 104116 15166
rect 103768 15096 104116 15102
rect 106216 15166 106526 15172
rect 106216 15102 106358 15166
rect 106422 15102 106494 15166
rect 106558 15102 106564 15166
rect 106216 15096 106526 15102
rect 121742 14855 121808 14858
rect 122320 14855 122386 14858
rect 121742 14853 122386 14855
rect 121742 14797 121747 14853
rect 121803 14797 122325 14853
rect 122381 14797 122386 14853
rect 121742 14795 122386 14797
rect 121742 14792 121808 14795
rect 122320 14792 122386 14795
rect 123216 14824 136620 14900
rect 123216 14782 123428 14824
rect 544 14758 3340 14764
rect 544 14694 550 14758
rect 614 14694 3340 14758
rect 544 14688 3340 14694
rect 3128 14628 3340 14688
rect 3944 14628 4156 14764
rect 3128 14552 4156 14628
rect 14552 14758 14764 14764
rect 14552 14694 14558 14758
rect 14622 14694 14764 14758
rect 14552 14622 14764 14694
rect 123216 14726 123270 14782
rect 123326 14726 123428 14782
rect 123216 14688 123428 14726
rect 14552 14558 14558 14622
rect 14622 14558 14764 14622
rect 14552 14552 14764 14558
rect 20128 14356 20340 14628
rect 21216 14622 21564 14628
rect 21216 14558 21358 14622
rect 21422 14558 21564 14622
rect 21216 14356 21564 14558
rect 20128 14350 21564 14356
rect 20128 14286 20270 14350
rect 20334 14286 21564 14350
rect 20128 14280 21564 14286
rect 28832 14350 29044 14492
rect 28832 14286 28838 14350
rect 28902 14286 29044 14350
rect 28832 14280 29044 14286
rect 31280 14350 31492 14492
rect 33728 14356 33940 14492
rect 33630 14350 33940 14356
rect 31280 14286 31422 14350
rect 31486 14286 31492 14350
rect 33592 14286 33598 14350
rect 33662 14286 33870 14350
rect 33934 14286 33940 14350
rect 31280 14280 31492 14286
rect 33630 14280 33940 14286
rect 36312 14350 36524 14492
rect 36312 14286 36454 14350
rect 36518 14286 36524 14350
rect 36312 14280 36524 14286
rect 38760 14356 38972 14492
rect 38760 14350 41148 14356
rect 38760 14286 38902 14350
rect 38966 14286 41078 14350
rect 41142 14286 41148 14350
rect 38760 14280 41148 14286
rect 41208 14350 41420 14492
rect 41208 14286 41214 14350
rect 41278 14286 41420 14350
rect 41208 14280 41420 14286
rect 43792 14350 44004 14492
rect 43792 14286 43798 14350
rect 43862 14286 44004 14350
rect 43792 14280 44004 14286
rect 46240 14350 46452 14492
rect 46240 14286 46246 14350
rect 46310 14286 46452 14350
rect 46240 14280 46452 14286
rect 48688 14350 49036 14492
rect 48688 14286 48830 14350
rect 48894 14286 49036 14350
rect 48688 14280 49036 14286
rect 51272 14350 51484 14492
rect 51272 14286 51414 14350
rect 51478 14286 51484 14350
rect 51272 14280 51484 14286
rect 53720 14356 53932 14492
rect 56168 14356 56516 14492
rect 58382 14486 58964 14492
rect 58344 14422 58350 14486
rect 58414 14422 58964 14486
rect 58382 14416 58964 14422
rect 58752 14356 58964 14416
rect 61200 14356 61412 14492
rect 53720 14350 56516 14356
rect 58654 14350 58964 14356
rect 61102 14350 61412 14356
rect 53720 14286 53862 14350
rect 53926 14286 56446 14350
rect 56510 14286 56516 14350
rect 58616 14286 58622 14350
rect 58686 14286 58894 14350
rect 58958 14286 58964 14350
rect 61064 14286 61070 14350
rect 61134 14286 61342 14350
rect 61406 14286 61412 14350
rect 53720 14280 56516 14286
rect 58654 14280 58964 14286
rect 61102 14280 61412 14286
rect 63648 14350 63996 14492
rect 63648 14286 63654 14350
rect 63718 14286 63790 14350
rect 63854 14286 63996 14350
rect 63648 14280 63996 14286
rect 66232 14350 66444 14492
rect 66232 14286 66238 14350
rect 66302 14286 66444 14350
rect 66232 14280 66444 14286
rect 68680 14350 68892 14492
rect 68680 14286 68822 14350
rect 68886 14286 68892 14350
rect 68680 14280 68892 14286
rect 71264 14350 71476 14492
rect 71264 14286 71270 14350
rect 71334 14286 71476 14350
rect 71264 14280 71476 14286
rect 73712 14350 73924 14492
rect 76160 14356 76372 14492
rect 76062 14350 76372 14356
rect 73712 14286 73854 14350
rect 73918 14286 73924 14350
rect 76024 14286 76030 14350
rect 76094 14286 76302 14350
rect 76366 14286 76372 14350
rect 73712 14280 73924 14286
rect 76062 14280 76372 14286
rect 78744 14350 78956 14492
rect 78744 14286 78886 14350
rect 78950 14286 78956 14350
rect 78744 14280 78956 14286
rect 81192 14350 81404 14492
rect 81192 14286 81334 14350
rect 81398 14286 81404 14350
rect 81192 14280 81404 14286
rect 83640 14350 83852 14492
rect 86224 14356 86436 14492
rect 86126 14350 86436 14356
rect 83640 14286 83646 14350
rect 83710 14286 83852 14350
rect 86088 14286 86094 14350
rect 86158 14286 86230 14350
rect 86294 14286 86436 14350
rect 83640 14280 83852 14286
rect 86126 14280 86436 14286
rect 88672 14350 88884 14492
rect 88672 14286 88678 14350
rect 88742 14286 88884 14350
rect 88672 14280 88884 14286
rect 91120 14350 91468 14492
rect 91120 14286 91262 14350
rect 91326 14286 91468 14350
rect 91120 14280 91468 14286
rect 93704 14350 93916 14492
rect 93704 14286 93846 14350
rect 93910 14286 93916 14350
rect 93704 14280 93916 14286
rect 96152 14356 96364 14492
rect 98600 14416 101396 14492
rect 98600 14356 98948 14416
rect 96152 14350 98948 14356
rect 96152 14286 96294 14350
rect 96358 14286 98878 14350
rect 98942 14286 98948 14350
rect 96152 14280 98948 14286
rect 101184 14350 101396 14416
rect 103632 14416 106428 14492
rect 103632 14356 103844 14416
rect 103534 14350 103844 14356
rect 101184 14286 101326 14350
rect 101390 14286 101396 14350
rect 103496 14286 103502 14350
rect 103566 14286 103774 14350
rect 103838 14286 103844 14350
rect 101184 14280 101396 14286
rect 103534 14280 103844 14286
rect 106080 14350 106428 14416
rect 106080 14286 106358 14350
rect 106422 14286 106428 14350
rect 106080 14280 106428 14286
rect 122808 14350 123020 14356
rect 122808 14286 122814 14350
rect 122878 14286 123020 14350
rect 122808 14078 123020 14286
rect 14661 14013 14727 14016
rect 26754 14013 26820 14016
rect 14661 14011 26820 14013
rect 14661 13955 14666 14011
rect 14722 13955 26759 14011
rect 26815 13955 26820 14011
rect 122808 14014 122814 14078
rect 122878 14014 123020 14078
rect 122808 14008 123020 14014
rect 14661 13953 26820 13955
rect 14661 13950 14727 13953
rect 26754 13950 26820 13953
rect 1224 13942 1980 13948
rect 1224 13878 1230 13942
rect 1294 13878 1980 13942
rect 1224 13872 1980 13878
rect 134776 13942 135396 13948
rect 134776 13878 135326 13942
rect 135390 13878 135396 13942
rect 134776 13872 135396 13878
rect 1768 13848 1980 13872
rect 1768 13792 1794 13848
rect 1850 13812 1980 13848
rect 134823 13848 134921 13872
rect 1850 13806 3204 13812
rect 1850 13792 3134 13806
rect 1768 13742 3134 13792
rect 3198 13742 3204 13806
rect 134823 13792 134844 13848
rect 134900 13792 134921 13848
rect 134823 13771 134921 13792
rect 1768 13736 3204 13742
rect 28832 13670 29044 13676
rect 28832 13606 28838 13670
rect 28902 13606 29044 13670
rect 28832 13600 29044 13606
rect 28851 13534 29044 13600
rect 28851 13487 28974 13534
rect 28968 13470 28974 13487
rect 29038 13470 29044 13534
rect 28968 13464 29044 13470
rect 31280 13670 33668 13676
rect 31280 13606 31422 13670
rect 31486 13606 33598 13670
rect 33662 13606 33668 13670
rect 31280 13600 33668 13606
rect 33728 13670 34076 13676
rect 33728 13606 33870 13670
rect 33934 13606 34076 13670
rect 33728 13600 34076 13606
rect 36312 13670 36524 13676
rect 36312 13606 36454 13670
rect 36518 13606 36524 13670
rect 36312 13600 36524 13606
rect 38760 13670 38972 13676
rect 41110 13670 41556 13676
rect 38760 13606 38902 13670
rect 38966 13606 38972 13670
rect 41072 13606 41078 13670
rect 41142 13606 41214 13670
rect 41278 13606 41556 13670
rect 38760 13600 38972 13606
rect 41110 13600 41556 13606
rect 43792 13670 44004 13676
rect 43792 13606 43798 13670
rect 43862 13606 44004 13670
rect 43792 13600 44004 13606
rect 46240 13670 49036 13676
rect 46240 13606 46246 13670
rect 46310 13606 48830 13670
rect 48894 13606 49036 13670
rect 46240 13600 49036 13606
rect 51272 13670 51484 13676
rect 51272 13606 51414 13670
rect 51478 13606 51484 13670
rect 51272 13600 51484 13606
rect 53720 13670 53932 13676
rect 53720 13606 53862 13670
rect 53926 13606 53932 13670
rect 53720 13600 53932 13606
rect 31280 13534 31492 13600
rect 31280 13470 31286 13534
rect 31350 13470 31492 13534
rect 33843 13534 34076 13600
rect 33843 13487 34006 13534
rect 31280 13464 31492 13470
rect 34000 13470 34006 13487
rect 34070 13470 34076 13534
rect 36339 13534 36524 13600
rect 36339 13487 36454 13534
rect 34000 13464 34076 13470
rect 36448 13470 36454 13487
rect 36518 13470 36524 13534
rect 38835 13534 38972 13600
rect 38835 13487 38902 13534
rect 36448 13464 36524 13470
rect 38896 13470 38902 13487
rect 38966 13470 38972 13534
rect 41331 13534 41556 13600
rect 41331 13487 41350 13534
rect 38896 13464 38972 13470
rect 41344 13470 41350 13487
rect 41414 13470 41556 13534
rect 43827 13534 44004 13600
rect 43827 13487 43934 13534
rect 41344 13464 41556 13470
rect 43928 13470 43934 13487
rect 43998 13470 44004 13534
rect 46323 13534 46452 13600
rect 46323 13487 46382 13534
rect 43928 13464 44004 13470
rect 46376 13470 46382 13487
rect 46446 13470 46452 13534
rect 48819 13534 49036 13600
rect 48819 13487 48966 13534
rect 46376 13464 46452 13470
rect 48960 13470 48966 13487
rect 49030 13470 49036 13534
rect 51315 13534 51484 13600
rect 51315 13487 51414 13534
rect 48960 13464 49036 13470
rect 51408 13470 51414 13487
rect 51478 13470 51484 13534
rect 53811 13534 53932 13600
rect 53811 13487 53862 13534
rect 51408 13464 51484 13470
rect 53856 13470 53862 13487
rect 53926 13470 53932 13534
rect 53856 13464 53932 13470
rect 56304 13670 58692 13676
rect 56304 13606 56446 13670
rect 56510 13606 58622 13670
rect 58686 13606 58692 13670
rect 56304 13600 58692 13606
rect 58752 13670 61140 13676
rect 58752 13606 58894 13670
rect 58958 13606 61070 13670
rect 61134 13606 61140 13670
rect 58752 13600 61140 13606
rect 61200 13670 63724 13676
rect 61200 13606 61206 13670
rect 61270 13606 61342 13670
rect 61406 13606 63654 13670
rect 63718 13606 63724 13670
rect 61200 13600 63724 13606
rect 63784 13670 63996 13676
rect 63784 13606 63790 13670
rect 63854 13606 63996 13670
rect 63784 13600 63996 13606
rect 66232 13670 66444 13676
rect 66232 13606 66238 13670
rect 66302 13606 66444 13670
rect 66232 13600 66444 13606
rect 68680 13670 68892 13676
rect 68680 13606 68686 13670
rect 68750 13606 68822 13670
rect 68886 13606 68892 13670
rect 68680 13600 68892 13606
rect 71264 13670 71476 13676
rect 71264 13606 71270 13670
rect 71334 13606 71476 13670
rect 71264 13600 71476 13606
rect 73712 13670 76100 13676
rect 73712 13606 73854 13670
rect 73918 13606 76030 13670
rect 76094 13606 76100 13670
rect 73712 13600 76100 13606
rect 76160 13670 76508 13676
rect 76160 13606 76302 13670
rect 76366 13606 76508 13670
rect 76160 13600 76508 13606
rect 78744 13670 78956 13676
rect 78744 13606 78886 13670
rect 78950 13606 78956 13670
rect 78744 13600 78956 13606
rect 81192 13670 81404 13676
rect 81192 13606 81334 13670
rect 81398 13606 81404 13670
rect 81192 13600 81404 13606
rect 83640 13670 86164 13676
rect 83640 13606 83646 13670
rect 83710 13606 86094 13670
rect 86158 13606 86164 13670
rect 83640 13600 86164 13606
rect 86224 13670 86436 13676
rect 86224 13606 86230 13670
rect 86294 13606 86436 13670
rect 86224 13600 86436 13606
rect 88672 13670 88884 13676
rect 88672 13606 88678 13670
rect 88742 13606 88884 13670
rect 88672 13600 88884 13606
rect 91120 13670 91468 13676
rect 91120 13606 91262 13670
rect 91326 13606 91468 13670
rect 91120 13600 91468 13606
rect 93704 13670 93916 13676
rect 93704 13606 93846 13670
rect 93910 13606 93916 13670
rect 93704 13600 93916 13606
rect 96152 13670 96364 13676
rect 96152 13606 96294 13670
rect 96358 13606 96364 13670
rect 96152 13600 96364 13606
rect 98736 13670 98948 13676
rect 98736 13606 98878 13670
rect 98942 13606 98948 13670
rect 98736 13600 98948 13606
rect 101184 13670 103572 13676
rect 101184 13606 101326 13670
rect 101390 13606 103502 13670
rect 103566 13606 103572 13670
rect 101184 13600 103572 13606
rect 103632 13670 103844 13676
rect 103632 13606 103638 13670
rect 103702 13606 103774 13670
rect 103838 13606 103844 13670
rect 103632 13600 103844 13606
rect 106216 13670 106428 13676
rect 106216 13606 106358 13670
rect 106422 13606 106428 13670
rect 106216 13600 106428 13606
rect 56304 13534 56516 13600
rect 56304 13470 56310 13534
rect 56374 13470 56516 13534
rect 58803 13534 58964 13600
rect 58803 13487 58894 13534
rect 56304 13464 56516 13470
rect 58888 13470 58894 13487
rect 58958 13470 58964 13534
rect 61299 13487 61397 13600
rect 63795 13534 63996 13600
rect 63795 13487 63926 13534
rect 58888 13464 58964 13470
rect 63920 13470 63926 13487
rect 63990 13470 63996 13534
rect 66291 13534 66444 13600
rect 66291 13487 66374 13534
rect 63920 13464 63996 13470
rect 66368 13470 66374 13487
rect 66438 13470 66444 13534
rect 68787 13487 68885 13600
rect 71283 13534 71476 13600
rect 71283 13487 71406 13534
rect 66368 13464 66444 13470
rect 71400 13470 71406 13487
rect 71470 13470 71476 13534
rect 73779 13534 73924 13600
rect 73779 13487 73854 13534
rect 71400 13464 71476 13470
rect 73848 13470 73854 13487
rect 73918 13470 73924 13534
rect 76275 13534 76508 13600
rect 76275 13487 76438 13534
rect 73848 13464 73924 13470
rect 76432 13470 76438 13487
rect 76502 13470 76508 13534
rect 78771 13534 78956 13600
rect 78771 13487 78886 13534
rect 76432 13464 76508 13470
rect 78880 13470 78886 13487
rect 78950 13470 78956 13534
rect 81267 13534 81404 13600
rect 81267 13487 81334 13534
rect 78880 13464 78956 13470
rect 81328 13470 81334 13487
rect 81398 13470 81404 13534
rect 83763 13534 83988 13600
rect 83763 13487 83918 13534
rect 81328 13464 81404 13470
rect 83912 13470 83918 13487
rect 83982 13470 83988 13534
rect 86259 13534 86436 13600
rect 86259 13487 86366 13534
rect 83912 13464 83988 13470
rect 86360 13470 86366 13487
rect 86430 13470 86436 13534
rect 88755 13534 88884 13600
rect 88755 13487 88814 13534
rect 86360 13464 86436 13470
rect 88808 13470 88814 13487
rect 88878 13470 88884 13534
rect 91251 13534 91468 13600
rect 91251 13487 91398 13534
rect 88808 13464 88884 13470
rect 91392 13470 91398 13487
rect 91462 13470 91468 13534
rect 93747 13534 93916 13600
rect 93747 13487 93846 13534
rect 91392 13464 91468 13470
rect 93840 13470 93846 13487
rect 93910 13470 93916 13534
rect 96243 13534 96364 13600
rect 96243 13487 96294 13534
rect 93840 13464 93916 13470
rect 96288 13470 96294 13487
rect 96358 13470 96364 13534
rect 98739 13534 98948 13600
rect 98739 13487 98878 13534
rect 96288 13464 96364 13470
rect 98872 13470 98878 13487
rect 98942 13470 98948 13534
rect 101235 13534 101396 13600
rect 101235 13487 101326 13534
rect 98872 13464 98948 13470
rect 101320 13470 101326 13487
rect 101390 13470 101396 13534
rect 103731 13487 103829 13600
rect 106227 13534 106428 13600
rect 123216 13654 136620 13676
rect 123216 13598 123270 13654
rect 123326 13600 136620 13654
rect 123326 13598 123428 13600
rect 106227 13487 106358 13534
rect 101320 13464 101396 13470
rect 106352 13470 106358 13487
rect 106422 13470 106428 13534
rect 121662 13585 121728 13588
rect 122320 13585 122386 13588
rect 121662 13583 122386 13585
rect 121662 13527 121667 13583
rect 121723 13527 122325 13583
rect 122381 13527 122386 13583
rect 121662 13525 122386 13527
rect 121662 13522 121728 13525
rect 122320 13522 122386 13525
rect 106352 13464 106428 13470
rect 123216 13464 123428 13598
rect 3128 13398 3340 13404
rect 3128 13334 3134 13398
rect 3198 13334 3340 13398
rect 3128 13268 3340 13334
rect 3944 13268 4156 13404
rect 3128 13192 4156 13268
rect 14552 13398 14764 13404
rect 14552 13334 14694 13398
rect 14758 13334 14764 13398
rect 14552 13262 14764 13334
rect 14552 13198 14694 13262
rect 14758 13198 14764 13262
rect 14552 13192 14764 13198
rect 28560 13261 28772 13404
rect 28968 13263 29180 13268
rect 28560 13205 28618 13261
rect 28674 13205 28772 13261
rect 28560 13132 28772 13205
rect 28851 13262 29180 13263
rect 28851 13198 29110 13262
rect 29174 13198 29180 13262
rect 28851 13192 29180 13198
rect 31008 13261 31220 13404
rect 33456 13328 33804 13404
rect 31008 13205 31114 13261
rect 31170 13205 31220 13261
rect 28851 13165 29044 13192
rect 20128 13126 21564 13132
rect 20128 13062 21222 13126
rect 21286 13062 21564 13126
rect 20128 13056 21564 13062
rect 28288 13126 28772 13132
rect 28288 13062 28294 13126
rect 28358 13062 28772 13126
rect 28288 13056 28772 13062
rect 28968 13132 29044 13165
rect 31008 13132 31220 13205
rect 28968 13126 29142 13132
rect 30736 13126 31220 13132
rect 28968 13062 29110 13126
rect 29174 13062 29180 13126
rect 30736 13062 30742 13126
rect 30806 13062 31220 13126
rect 28968 13056 29142 13062
rect 30736 13056 31220 13062
rect 31280 13262 31628 13268
rect 31280 13198 31558 13262
rect 31622 13198 31628 13262
rect 31280 13192 31628 13198
rect 33456 13261 33687 13328
rect 34000 13263 34212 13268
rect 33456 13205 33610 13261
rect 33666 13205 33687 13261
rect 31280 13126 31492 13192
rect 31280 13062 31422 13126
rect 31486 13062 31492 13126
rect 31280 13056 31492 13062
rect 33456 13184 33687 13205
rect 33843 13262 34212 13263
rect 33843 13198 34142 13262
rect 34206 13198 34212 13262
rect 33843 13192 34212 13198
rect 36040 13261 36252 13404
rect 36448 13263 36660 13268
rect 36040 13205 36106 13261
rect 36162 13205 36252 13261
rect 33456 13126 33668 13184
rect 33843 13165 34076 13192
rect 33456 13062 33598 13126
rect 33662 13062 33668 13126
rect 33456 13056 33668 13062
rect 33864 13126 34076 13165
rect 33864 13062 33870 13126
rect 33934 13062 34076 13126
rect 33864 13056 34076 13062
rect 36040 13126 36252 13205
rect 36339 13262 36660 13263
rect 36339 13198 36590 13262
rect 36654 13198 36660 13262
rect 36339 13192 36660 13198
rect 38488 13261 38700 13404
rect 41072 13328 41284 13404
rect 38896 13263 39108 13268
rect 38488 13205 38602 13261
rect 38658 13205 38700 13261
rect 36339 13165 36524 13192
rect 36040 13062 36046 13126
rect 36110 13062 36252 13126
rect 36040 13056 36252 13062
rect 36448 13132 36524 13165
rect 36448 13126 36622 13132
rect 38488 13126 38700 13205
rect 38835 13262 39108 13263
rect 38835 13198 39038 13262
rect 39102 13198 39108 13262
rect 38835 13192 39108 13198
rect 41072 13261 41175 13328
rect 41344 13263 41556 13268
rect 41072 13205 41098 13261
rect 41154 13205 41175 13261
rect 38835 13165 38972 13192
rect 36448 13062 36590 13126
rect 36654 13062 36660 13126
rect 38488 13062 38494 13126
rect 38558 13062 38700 13126
rect 36448 13056 36622 13062
rect 38488 13056 38700 13062
rect 38896 13132 38972 13165
rect 41072 13184 41175 13205
rect 41331 13262 41556 13263
rect 41331 13198 41486 13262
rect 41550 13198 41556 13262
rect 38896 13126 39070 13132
rect 41072 13126 41148 13184
rect 41331 13165 41556 13198
rect 38896 13062 39038 13126
rect 39102 13062 39108 13126
rect 41072 13062 41078 13126
rect 41142 13062 41148 13126
rect 38896 13056 39070 13062
rect 41072 13056 41148 13062
rect 41344 13126 41556 13165
rect 41344 13062 41486 13126
rect 41550 13062 41556 13126
rect 41344 13056 41556 13062
rect 43520 13261 43732 13404
rect 43928 13263 44140 13268
rect 43520 13205 43594 13261
rect 43650 13205 43732 13261
rect 43520 13126 43732 13205
rect 43827 13262 44140 13263
rect 43827 13198 44070 13262
rect 44134 13198 44140 13262
rect 43827 13192 44140 13198
rect 45968 13261 46180 13404
rect 48552 13328 48764 13404
rect 46376 13263 46588 13268
rect 45968 13205 46090 13261
rect 46146 13205 46180 13261
rect 43827 13165 44004 13192
rect 43520 13062 43526 13126
rect 43590 13062 43732 13126
rect 43520 13056 43732 13062
rect 43928 13132 44004 13165
rect 43928 13126 44102 13132
rect 45968 13126 46180 13205
rect 46323 13262 46588 13263
rect 46323 13198 46518 13262
rect 46582 13198 46588 13262
rect 46323 13192 46588 13198
rect 48552 13261 48663 13328
rect 48960 13263 49172 13268
rect 48552 13205 48586 13261
rect 48642 13205 48663 13261
rect 46323 13165 46452 13192
rect 43928 13062 44070 13126
rect 44134 13062 44140 13126
rect 45968 13062 45974 13126
rect 46038 13062 46180 13126
rect 43928 13056 44102 13062
rect 45968 13056 46180 13062
rect 46376 13132 46452 13165
rect 48552 13184 48663 13205
rect 48819 13262 49172 13263
rect 48819 13198 49102 13262
rect 49166 13198 49172 13262
rect 48819 13192 49172 13198
rect 51000 13261 51212 13404
rect 51408 13263 51620 13268
rect 51000 13205 51082 13261
rect 51138 13205 51212 13261
rect 48552 13132 48628 13184
rect 48819 13165 49036 13192
rect 46376 13126 46550 13132
rect 48280 13126 48628 13132
rect 46376 13062 46518 13126
rect 46582 13062 46588 13126
rect 48280 13062 48286 13126
rect 48350 13062 48628 13126
rect 46376 13056 46550 13062
rect 48280 13056 48628 13062
rect 48824 13126 49036 13165
rect 48824 13062 48830 13126
rect 48894 13062 49036 13126
rect 48824 13056 49036 13062
rect 51000 13126 51212 13205
rect 51315 13262 51620 13263
rect 51315 13198 51550 13262
rect 51614 13198 51620 13262
rect 51315 13192 51620 13198
rect 53448 13261 53660 13404
rect 53856 13263 54068 13268
rect 53448 13205 53578 13261
rect 53634 13205 53660 13261
rect 51315 13165 51484 13192
rect 51000 13062 51006 13126
rect 51070 13062 51212 13126
rect 51000 13056 51212 13062
rect 51408 13132 51484 13165
rect 51408 13126 51582 13132
rect 53448 13126 53660 13205
rect 53811 13262 54068 13263
rect 53811 13198 53998 13262
rect 54062 13198 54068 13262
rect 53811 13192 54068 13198
rect 56032 13261 56244 13404
rect 56032 13205 56074 13261
rect 56130 13205 56244 13261
rect 53811 13165 53932 13192
rect 51408 13062 51550 13126
rect 51614 13062 51620 13126
rect 53448 13062 53590 13126
rect 53654 13062 53660 13126
rect 51408 13056 51582 13062
rect 53448 13056 53660 13062
rect 53856 13132 53932 13165
rect 53856 13126 54030 13132
rect 56032 13126 56244 13205
rect 53856 13062 53998 13126
rect 54062 13062 54068 13126
rect 56032 13062 56038 13126
rect 56102 13062 56244 13126
rect 53856 13056 54030 13062
rect 56032 13056 56244 13062
rect 56304 13262 56652 13268
rect 56304 13198 56582 13262
rect 56646 13198 56652 13262
rect 56304 13192 56652 13198
rect 58480 13261 58692 13404
rect 60928 13328 61276 13404
rect 58888 13263 59100 13268
rect 58480 13205 58570 13261
rect 58626 13205 58692 13261
rect 56304 13126 56516 13192
rect 56304 13062 56446 13126
rect 56510 13062 56516 13126
rect 56304 13056 56516 13062
rect 58480 13126 58692 13205
rect 58803 13262 59100 13263
rect 58803 13198 59030 13262
rect 59094 13198 59100 13262
rect 58803 13192 59100 13198
rect 60928 13261 61143 13328
rect 60928 13205 61066 13261
rect 61122 13205 61143 13261
rect 58803 13165 58964 13192
rect 58480 13062 58486 13126
rect 58550 13062 58692 13126
rect 58480 13056 58692 13062
rect 58888 13132 58964 13165
rect 60928 13184 61143 13205
rect 58888 13126 59062 13132
rect 60928 13126 61140 13184
rect 58888 13062 59030 13126
rect 59094 13062 59100 13126
rect 60928 13062 60934 13126
rect 60998 13062 61140 13126
rect 61299 13132 61397 13263
rect 63512 13261 63724 13404
rect 63920 13263 64132 13268
rect 63512 13205 63562 13261
rect 63618 13205 63724 13261
rect 61299 13126 61548 13132
rect 61299 13094 61342 13126
rect 58888 13056 59062 13062
rect 60928 13056 61140 13062
rect 61336 13062 61342 13094
rect 61406 13062 61478 13126
rect 61542 13062 61548 13126
rect 61336 13056 61548 13062
rect 63512 13126 63724 13205
rect 63795 13262 64132 13263
rect 63795 13198 64062 13262
rect 64126 13198 64132 13262
rect 63795 13192 64132 13198
rect 65960 13261 66172 13404
rect 68408 13328 68756 13404
rect 66368 13263 66580 13268
rect 65960 13205 66058 13261
rect 66114 13205 66172 13261
rect 63795 13165 63996 13192
rect 63512 13062 63518 13126
rect 63582 13062 63724 13126
rect 63512 13056 63724 13062
rect 63920 13132 63996 13165
rect 63920 13126 64094 13132
rect 65960 13126 66172 13205
rect 66291 13262 66580 13263
rect 66291 13198 66510 13262
rect 66574 13198 66580 13262
rect 66291 13192 66580 13198
rect 68408 13261 68631 13328
rect 68408 13205 68554 13261
rect 68610 13205 68631 13261
rect 66291 13165 66444 13192
rect 63920 13062 64062 13126
rect 64126 13062 64132 13126
rect 65960 13062 65966 13126
rect 66030 13062 66172 13126
rect 63920 13056 64094 13062
rect 65960 13056 66172 13062
rect 66368 13132 66444 13165
rect 68408 13184 68631 13205
rect 68408 13132 68620 13184
rect 66368 13126 66542 13132
rect 68272 13126 68620 13132
rect 66368 13062 66510 13126
rect 66574 13062 66580 13126
rect 68272 13062 68278 13126
rect 68342 13062 68620 13126
rect 68787 13132 68885 13263
rect 70992 13261 71204 13404
rect 71400 13263 71612 13268
rect 70992 13205 71050 13261
rect 71106 13205 71204 13261
rect 68787 13126 69028 13132
rect 68787 13094 68822 13126
rect 66368 13056 66542 13062
rect 68272 13056 68620 13062
rect 68816 13062 68822 13094
rect 68886 13062 68958 13126
rect 69022 13062 69028 13126
rect 68816 13056 69028 13062
rect 70992 13126 71204 13205
rect 71283 13262 71612 13263
rect 71283 13198 71542 13262
rect 71606 13198 71612 13262
rect 71283 13192 71612 13198
rect 73440 13261 73652 13404
rect 75888 13328 76236 13404
rect 73848 13263 74060 13268
rect 73440 13205 73546 13261
rect 73602 13205 73652 13261
rect 71283 13165 71476 13192
rect 70992 13062 70998 13126
rect 71062 13062 71204 13126
rect 70992 13056 71204 13062
rect 71400 13132 71476 13165
rect 71400 13126 71574 13132
rect 73440 13126 73652 13205
rect 73779 13262 74060 13263
rect 73779 13198 73990 13262
rect 74054 13198 74060 13262
rect 73779 13192 74060 13198
rect 75888 13261 76119 13328
rect 76432 13263 76644 13268
rect 75888 13205 76042 13261
rect 76098 13205 76119 13261
rect 73779 13165 73924 13192
rect 71400 13062 71542 13126
rect 71606 13062 71612 13126
rect 73440 13062 73446 13126
rect 73510 13062 73652 13126
rect 71400 13056 71574 13062
rect 73440 13056 73652 13062
rect 73848 13132 73924 13165
rect 75888 13184 76119 13205
rect 76275 13262 76644 13263
rect 76275 13198 76574 13262
rect 76638 13198 76644 13262
rect 76275 13192 76644 13198
rect 78472 13261 78684 13404
rect 78880 13263 79092 13268
rect 78472 13205 78538 13261
rect 78594 13205 78684 13261
rect 73848 13126 74022 13132
rect 75888 13126 76100 13184
rect 76275 13165 76508 13192
rect 73848 13062 73990 13126
rect 74054 13062 74060 13126
rect 75888 13062 75894 13126
rect 75958 13062 76100 13126
rect 73848 13056 74022 13062
rect 75888 13056 76100 13062
rect 76296 13126 76508 13165
rect 76296 13062 76302 13126
rect 76366 13062 76508 13126
rect 76296 13056 76508 13062
rect 78472 13126 78684 13205
rect 78771 13262 79092 13263
rect 78771 13198 79022 13262
rect 79086 13198 79092 13262
rect 78771 13192 79092 13198
rect 80920 13261 81132 13404
rect 83504 13328 83716 13404
rect 81328 13263 81540 13268
rect 80920 13205 81034 13261
rect 81090 13205 81132 13261
rect 78771 13165 78956 13192
rect 78472 13062 78478 13126
rect 78542 13062 78684 13126
rect 78472 13056 78684 13062
rect 78880 13132 78956 13165
rect 78880 13126 79054 13132
rect 80920 13126 81132 13205
rect 81267 13262 81540 13263
rect 81267 13198 81470 13262
rect 81534 13198 81540 13262
rect 81267 13192 81540 13198
rect 83504 13261 83607 13328
rect 83912 13263 84124 13268
rect 83504 13205 83530 13261
rect 83586 13205 83607 13261
rect 81267 13165 81404 13192
rect 78880 13062 79022 13126
rect 79086 13062 79092 13126
rect 80920 13062 80926 13126
rect 80990 13062 81132 13126
rect 78880 13056 79054 13062
rect 80920 13056 81132 13062
rect 81328 13132 81404 13165
rect 83504 13184 83607 13205
rect 83763 13262 84124 13263
rect 83763 13198 84054 13262
rect 84118 13198 84124 13262
rect 83763 13192 84124 13198
rect 85952 13261 86164 13404
rect 86360 13263 86572 13268
rect 85952 13205 86026 13261
rect 86082 13205 86164 13261
rect 81328 13126 81502 13132
rect 83504 13126 83580 13184
rect 83763 13165 83988 13192
rect 81328 13062 81470 13126
rect 81534 13062 81540 13126
rect 83504 13062 83510 13126
rect 83574 13062 83580 13126
rect 81328 13056 81502 13062
rect 83504 13056 83580 13062
rect 83776 13126 83988 13165
rect 83776 13062 83782 13126
rect 83846 13062 83988 13126
rect 83776 13056 83988 13062
rect 85952 13126 86164 13205
rect 86259 13262 86572 13263
rect 86259 13198 86502 13262
rect 86566 13198 86572 13262
rect 86259 13192 86572 13198
rect 88400 13261 88612 13404
rect 90984 13328 91196 13404
rect 88808 13263 89020 13268
rect 88400 13205 88522 13261
rect 88578 13205 88612 13261
rect 86259 13165 86436 13192
rect 85952 13062 85958 13126
rect 86022 13062 86164 13126
rect 85952 13056 86164 13062
rect 86360 13132 86436 13165
rect 86360 13126 86534 13132
rect 88400 13126 88612 13205
rect 88755 13262 89020 13263
rect 88755 13198 88950 13262
rect 89014 13198 89020 13262
rect 88755 13192 89020 13198
rect 90984 13261 91095 13328
rect 91392 13263 91604 13268
rect 90984 13205 91018 13261
rect 91074 13205 91095 13261
rect 88755 13165 88884 13192
rect 86360 13062 86502 13126
rect 86566 13062 86572 13126
rect 88400 13062 88542 13126
rect 88606 13062 88612 13126
rect 86360 13056 86534 13062
rect 88400 13056 88612 13062
rect 88808 13132 88884 13165
rect 90984 13184 91095 13205
rect 91251 13262 91604 13263
rect 91251 13198 91534 13262
rect 91598 13198 91604 13262
rect 91251 13192 91604 13198
rect 93432 13261 93644 13404
rect 93840 13263 94052 13268
rect 93432 13205 93514 13261
rect 93570 13205 93644 13261
rect 88808 13126 88982 13132
rect 90984 13126 91060 13184
rect 91251 13165 91468 13192
rect 88808 13062 88950 13126
rect 89014 13062 89020 13126
rect 90984 13062 90990 13126
rect 91054 13062 91060 13126
rect 88808 13056 88982 13062
rect 90984 13056 91060 13062
rect 91256 13126 91468 13165
rect 91256 13062 91262 13126
rect 91326 13062 91468 13126
rect 91256 13056 91468 13062
rect 93432 13126 93644 13205
rect 93747 13262 94052 13263
rect 93747 13198 93982 13262
rect 94046 13198 94052 13262
rect 93747 13192 94052 13198
rect 95880 13261 96092 13404
rect 96288 13263 96500 13268
rect 95880 13205 96010 13261
rect 96066 13205 96092 13261
rect 93747 13165 93916 13192
rect 93432 13062 93438 13126
rect 93502 13062 93644 13126
rect 93432 13056 93644 13062
rect 93840 13132 93916 13165
rect 93840 13126 94014 13132
rect 95880 13126 96092 13205
rect 96243 13262 96500 13263
rect 96243 13198 96430 13262
rect 96494 13198 96500 13262
rect 96243 13192 96500 13198
rect 98464 13261 98676 13404
rect 98872 13263 99084 13268
rect 98464 13205 98506 13261
rect 98562 13205 98676 13261
rect 96243 13165 96364 13192
rect 93840 13062 93982 13126
rect 94046 13062 94052 13126
rect 95880 13062 95886 13126
rect 95950 13062 96092 13126
rect 93840 13056 94014 13062
rect 95880 13056 96092 13062
rect 96288 13132 96364 13165
rect 96288 13126 96462 13132
rect 98464 13126 98676 13205
rect 98739 13262 99084 13263
rect 98739 13198 99014 13262
rect 99078 13198 99084 13262
rect 98739 13192 99084 13198
rect 100912 13261 101124 13404
rect 103360 13328 103708 13404
rect 101320 13263 101532 13268
rect 100912 13205 101002 13261
rect 101058 13205 101124 13261
rect 98739 13165 98948 13192
rect 96288 13062 96430 13126
rect 96494 13062 96500 13126
rect 98464 13062 98470 13126
rect 98534 13062 98676 13126
rect 96288 13056 96462 13062
rect 98464 13056 98676 13062
rect 98872 13132 98948 13165
rect 98872 13126 99046 13132
rect 100912 13126 101124 13205
rect 101235 13262 101532 13263
rect 101235 13198 101462 13262
rect 101526 13198 101532 13262
rect 101235 13192 101532 13198
rect 103360 13261 103575 13328
rect 103360 13205 103498 13261
rect 103554 13205 103575 13261
rect 101235 13165 101396 13192
rect 98872 13062 99014 13126
rect 99078 13062 99084 13126
rect 100912 13062 100918 13126
rect 100982 13062 101124 13126
rect 98872 13056 99046 13062
rect 100912 13056 101124 13062
rect 101320 13132 101396 13165
rect 103360 13184 103575 13205
rect 101320 13126 101494 13132
rect 103360 13126 103572 13184
rect 101320 13062 101462 13126
rect 101526 13062 101532 13126
rect 103360 13062 103366 13126
rect 103430 13062 103572 13126
rect 103731 13132 103829 13263
rect 105944 13261 106156 13404
rect 106352 13263 106564 13268
rect 105944 13205 105994 13261
rect 106050 13205 106156 13261
rect 103731 13126 103980 13132
rect 103731 13094 103774 13126
rect 101320 13056 101494 13062
rect 103360 13056 103572 13062
rect 103768 13062 103774 13094
rect 103838 13062 103910 13126
rect 103974 13062 103980 13126
rect 103768 13056 103980 13062
rect 105944 13126 106156 13205
rect 106227 13262 106564 13263
rect 106227 13198 106494 13262
rect 106558 13198 106564 13262
rect 106227 13192 106564 13198
rect 106227 13165 106428 13192
rect 105944 13062 105950 13126
rect 106014 13062 106156 13126
rect 105944 13056 106156 13062
rect 106352 13132 106428 13165
rect 106352 13126 106526 13132
rect 106352 13062 106494 13126
rect 106558 13062 106564 13126
rect 106352 13056 106526 13062
rect 20128 12920 20340 13056
rect 21216 12920 21564 13056
rect 122808 12854 123020 12860
rect 122808 12790 122950 12854
rect 123014 12790 123020 12854
rect 122808 12718 123020 12790
rect 122808 12654 122950 12718
rect 123014 12654 123020 12718
rect 122808 12648 123020 12654
rect 14661 12599 14727 12602
rect 26630 12599 26696 12602
rect 14661 12597 26696 12599
rect 14661 12541 14666 12597
rect 14722 12541 26635 12597
rect 26691 12541 26696 12597
rect 14661 12539 26696 12541
rect 14661 12536 14727 12539
rect 26630 12536 26696 12539
rect 28696 12582 29180 12588
rect 28696 12518 29110 12582
rect 29174 12518 29180 12582
rect 28696 12512 29180 12518
rect 31144 12582 31492 12588
rect 31144 12518 31422 12582
rect 31486 12518 31492 12582
rect 31144 12512 31492 12518
rect 33728 12582 33940 12588
rect 33728 12518 33870 12582
rect 33934 12518 33940 12582
rect 1224 12310 1980 12316
rect 1224 12246 1230 12310
rect 1294 12246 1980 12310
rect 1224 12240 1980 12246
rect 28696 12310 28908 12512
rect 28696 12246 28838 12310
rect 28902 12246 28908 12310
rect 28696 12240 28908 12246
rect 31144 12316 31356 12512
rect 33728 12316 33940 12518
rect 31144 12310 31492 12316
rect 31144 12246 31422 12310
rect 31486 12246 31492 12310
rect 31144 12240 31492 12246
rect 33456 12310 33940 12316
rect 33456 12246 33462 12310
rect 33526 12246 33940 12310
rect 33456 12240 33940 12246
rect 36176 12582 36660 12588
rect 36176 12518 36590 12582
rect 36654 12518 36660 12582
rect 36176 12512 36660 12518
rect 38624 12582 39108 12588
rect 38624 12518 39038 12582
rect 39102 12518 39108 12582
rect 38624 12512 39108 12518
rect 41208 12582 41556 12588
rect 41208 12518 41486 12582
rect 41550 12518 41556 12582
rect 41208 12512 41556 12518
rect 43656 12582 44140 12588
rect 43656 12518 44070 12582
rect 44134 12518 44140 12582
rect 43656 12512 44140 12518
rect 46104 12582 46588 12588
rect 46104 12518 46518 12582
rect 46582 12518 46588 12582
rect 46104 12512 46588 12518
rect 48688 12582 48900 12588
rect 48688 12518 48830 12582
rect 48894 12518 48900 12582
rect 36176 12310 36388 12512
rect 36176 12246 36182 12310
rect 36246 12246 36388 12310
rect 36176 12240 36388 12246
rect 38624 12310 38836 12512
rect 38624 12246 38630 12310
rect 38694 12246 38836 12310
rect 38624 12240 38836 12246
rect 41208 12316 41420 12512
rect 43656 12316 43868 12512
rect 41208 12310 41556 12316
rect 43422 12310 43868 12316
rect 41208 12246 41486 12310
rect 41550 12246 41556 12310
rect 43384 12246 43390 12310
rect 43454 12246 43868 12310
rect 41208 12240 41556 12246
rect 43422 12240 43868 12246
rect 46104 12316 46316 12512
rect 46104 12310 46588 12316
rect 46104 12246 46518 12310
rect 46582 12246 46588 12310
rect 46104 12240 46588 12246
rect 48688 12310 48900 12518
rect 48688 12246 48830 12310
rect 48894 12246 48900 12310
rect 48688 12240 48900 12246
rect 51136 12582 51620 12588
rect 51136 12518 51550 12582
rect 51614 12518 51620 12582
rect 51136 12512 51620 12518
rect 53584 12582 54068 12588
rect 53584 12518 53998 12582
rect 54062 12518 54068 12582
rect 53584 12512 54068 12518
rect 56168 12582 56516 12588
rect 56168 12518 56446 12582
rect 56510 12518 56516 12582
rect 56168 12512 56516 12518
rect 58616 12582 59100 12588
rect 58616 12518 59030 12582
rect 59094 12518 59100 12582
rect 58616 12512 59100 12518
rect 61064 12582 61412 12588
rect 61064 12518 61342 12582
rect 61406 12518 61412 12582
rect 51136 12310 51348 12512
rect 51136 12246 51278 12310
rect 51342 12246 51348 12310
rect 51136 12240 51348 12246
rect 53584 12316 53796 12512
rect 56168 12316 56380 12512
rect 58616 12316 58828 12512
rect 53584 12310 54068 12316
rect 53584 12246 53998 12310
rect 54062 12246 54068 12310
rect 53584 12240 54068 12246
rect 56168 12310 56516 12316
rect 56168 12246 56446 12310
rect 56510 12246 56516 12310
rect 56168 12240 56516 12246
rect 58616 12310 59100 12316
rect 58616 12246 59030 12310
rect 59094 12246 59100 12310
rect 58616 12240 59100 12246
rect 61064 12310 61412 12518
rect 61064 12246 61342 12310
rect 61406 12246 61412 12310
rect 61064 12240 61412 12246
rect 63648 12582 64132 12588
rect 63648 12518 64062 12582
rect 64126 12518 64132 12582
rect 63648 12512 64132 12518
rect 66096 12582 66580 12588
rect 66096 12518 66510 12582
rect 66574 12518 66580 12582
rect 66096 12512 66580 12518
rect 68544 12582 68892 12588
rect 68544 12518 68822 12582
rect 68886 12518 68892 12582
rect 63648 12310 63860 12512
rect 63648 12246 63654 12310
rect 63718 12246 63860 12310
rect 63648 12240 63860 12246
rect 66096 12310 66308 12512
rect 66096 12246 66238 12310
rect 66302 12246 66308 12310
rect 66096 12240 66308 12246
rect 68544 12310 68892 12518
rect 68544 12246 68550 12310
rect 68614 12246 68892 12310
rect 68544 12240 68892 12246
rect 71128 12582 71612 12588
rect 71128 12518 71542 12582
rect 71606 12518 71612 12582
rect 71128 12512 71612 12518
rect 73576 12582 74060 12588
rect 73576 12518 73990 12582
rect 74054 12518 74060 12582
rect 73576 12512 74060 12518
rect 76160 12582 76372 12588
rect 76160 12518 76302 12582
rect 76366 12518 76372 12582
rect 71128 12316 71340 12512
rect 73576 12316 73788 12512
rect 71128 12310 71612 12316
rect 73342 12310 73788 12316
rect 71128 12246 71542 12310
rect 71606 12246 71612 12310
rect 73304 12246 73310 12310
rect 73374 12246 73788 12310
rect 71128 12240 71612 12246
rect 73342 12240 73788 12246
rect 76160 12310 76372 12518
rect 76160 12246 76166 12310
rect 76230 12246 76372 12310
rect 76160 12240 76372 12246
rect 78608 12582 79092 12588
rect 78608 12518 79022 12582
rect 79086 12518 79092 12582
rect 78608 12512 79092 12518
rect 81056 12582 81540 12588
rect 81056 12518 81470 12582
rect 81534 12518 81540 12582
rect 81056 12512 81540 12518
rect 83640 12582 83852 12588
rect 83640 12518 83782 12582
rect 83846 12518 83852 12582
rect 78608 12310 78820 12512
rect 78608 12246 78614 12310
rect 78678 12246 78820 12310
rect 78608 12240 78820 12246
rect 81056 12310 81268 12512
rect 81056 12246 81062 12310
rect 81126 12246 81268 12310
rect 81056 12240 81268 12246
rect 83640 12316 83852 12518
rect 86088 12582 86572 12588
rect 86088 12518 86502 12582
rect 86566 12518 86572 12582
rect 86088 12512 86572 12518
rect 88536 12582 89020 12588
rect 88536 12518 88950 12582
rect 89014 12518 89020 12582
rect 88536 12512 89020 12518
rect 91120 12582 91332 12588
rect 91120 12518 91262 12582
rect 91326 12518 91332 12582
rect 86088 12316 86300 12512
rect 88536 12316 88748 12512
rect 83640 12310 84124 12316
rect 83640 12246 84054 12310
rect 84118 12246 84124 12310
rect 83640 12240 84124 12246
rect 86088 12310 86572 12316
rect 86088 12246 86502 12310
rect 86566 12246 86572 12310
rect 86088 12240 86572 12246
rect 88536 12310 89020 12316
rect 88536 12246 88950 12310
rect 89014 12246 89020 12310
rect 88536 12240 89020 12246
rect 91120 12310 91332 12518
rect 91120 12246 91262 12310
rect 91326 12246 91332 12310
rect 91120 12240 91332 12246
rect 93568 12582 94052 12588
rect 93568 12518 93982 12582
rect 94046 12518 94052 12582
rect 93568 12512 94052 12518
rect 96016 12582 96500 12588
rect 96016 12518 96430 12582
rect 96494 12518 96500 12582
rect 96016 12512 96500 12518
rect 98600 12582 99084 12588
rect 98600 12518 99014 12582
rect 99078 12518 99084 12582
rect 98600 12512 99084 12518
rect 101048 12582 101532 12588
rect 101048 12518 101462 12582
rect 101526 12518 101532 12582
rect 101048 12512 101532 12518
rect 103496 12582 103844 12588
rect 103496 12518 103774 12582
rect 103838 12518 103844 12582
rect 93568 12310 93780 12512
rect 93568 12246 93710 12310
rect 93774 12246 93780 12310
rect 93568 12240 93780 12246
rect 96016 12310 96228 12512
rect 96016 12246 96022 12310
rect 96086 12246 96228 12310
rect 96016 12240 96228 12246
rect 98600 12316 98812 12512
rect 101048 12316 101260 12512
rect 98600 12310 99084 12316
rect 98600 12246 99014 12310
rect 99078 12246 99084 12310
rect 98600 12240 99084 12246
rect 101048 12310 101532 12316
rect 101048 12246 101462 12310
rect 101526 12246 101532 12310
rect 101048 12240 101532 12246
rect 103496 12310 103844 12518
rect 103496 12246 103774 12310
rect 103838 12246 103844 12310
rect 103496 12240 103844 12246
rect 106080 12582 106564 12588
rect 106080 12518 106494 12582
rect 106558 12518 106564 12582
rect 106080 12512 106564 12518
rect 106080 12310 106292 12512
rect 106080 12246 106086 12310
rect 106150 12246 106292 12310
rect 106080 12240 106292 12246
rect 134776 12310 135396 12316
rect 134776 12246 135326 12310
rect 135390 12246 135396 12310
rect 134776 12240 135396 12246
rect 1768 12168 1980 12240
rect 1768 12112 1794 12168
rect 1850 12112 1980 12168
rect 1768 11968 1980 12112
rect 134776 12168 134988 12240
rect 134776 12112 134844 12168
rect 134900 12112 134988 12168
rect 14552 12038 14764 12044
rect 14552 11974 14558 12038
rect 14622 11974 14764 12038
rect 14552 11766 14764 11974
rect 28696 12038 29044 12044
rect 28696 11974 28974 12038
rect 29038 11974 29044 12038
rect 28696 11968 29044 11974
rect 31144 12038 31356 12044
rect 31144 11974 31286 12038
rect 31350 11974 31356 12038
rect 28696 11902 28908 11968
rect 28696 11838 28702 11902
rect 28766 11838 28908 11902
rect 28696 11832 28908 11838
rect 31144 11902 31356 11974
rect 31144 11838 31150 11902
rect 31214 11838 31356 11902
rect 31144 11832 31356 11838
rect 33592 12038 34076 12044
rect 33592 11974 34006 12038
rect 34070 11974 34076 12038
rect 33592 11968 34076 11974
rect 36176 12038 36524 12044
rect 36176 11974 36454 12038
rect 36518 11974 36524 12038
rect 36176 11968 36524 11974
rect 38624 12038 38972 12044
rect 38624 11974 38902 12038
rect 38966 11974 38972 12038
rect 38624 11968 38972 11974
rect 41072 12038 44004 12044
rect 41072 11974 41350 12038
rect 41414 11974 43934 12038
rect 43998 11974 44004 12038
rect 41072 11968 44004 11974
rect 46104 12038 46452 12044
rect 46104 11974 46382 12038
rect 46446 11974 46452 12038
rect 46104 11968 46452 11974
rect 48688 12038 49036 12044
rect 48688 11974 48966 12038
rect 49030 11974 49036 12038
rect 48688 11968 49036 11974
rect 51136 12038 51484 12044
rect 51136 11974 51414 12038
rect 51478 11974 51484 12038
rect 51136 11968 51484 11974
rect 53584 12038 53932 12044
rect 53584 11974 53862 12038
rect 53926 11974 53932 12038
rect 53584 11968 53932 11974
rect 56168 12038 56380 12044
rect 56168 11974 56310 12038
rect 56374 11974 56380 12038
rect 33592 11902 33940 11968
rect 33592 11838 33870 11902
rect 33934 11838 33940 11902
rect 33592 11832 33940 11838
rect 36176 11908 36388 11968
rect 38624 11908 38836 11968
rect 36176 11902 38836 11908
rect 36176 11838 36318 11902
rect 36382 11838 38766 11902
rect 38830 11838 38836 11902
rect 36176 11832 38836 11838
rect 41072 11902 41420 11968
rect 41072 11838 41350 11902
rect 41414 11838 41420 11902
rect 41072 11832 41420 11838
rect 43656 11902 43868 11968
rect 43656 11838 43798 11902
rect 43862 11838 43868 11902
rect 43656 11832 43868 11838
rect 46104 11902 46316 11968
rect 46104 11838 46246 11902
rect 46310 11838 46316 11902
rect 46104 11832 46316 11838
rect 48688 11902 48900 11968
rect 48688 11838 48694 11902
rect 48758 11838 48900 11902
rect 48688 11832 48900 11838
rect 51136 11902 51348 11968
rect 51136 11838 51142 11902
rect 51206 11838 51348 11902
rect 51136 11832 51348 11838
rect 53584 11908 53796 11968
rect 53584 11902 53932 11908
rect 53584 11838 53862 11902
rect 53926 11838 53932 11902
rect 53584 11832 53932 11838
rect 56168 11902 56380 11974
rect 56168 11838 56310 11902
rect 56374 11838 56380 11902
rect 56168 11832 56380 11838
rect 58616 12038 58964 12044
rect 58616 11974 58894 12038
rect 58958 11974 58964 12038
rect 58616 11968 58964 11974
rect 61064 12038 61276 12044
rect 61064 11974 61206 12038
rect 61270 11974 61276 12038
rect 58616 11902 58828 11968
rect 58616 11838 58758 11902
rect 58822 11838 58828 11902
rect 58616 11832 58828 11838
rect 61064 11902 61276 11974
rect 61064 11838 61206 11902
rect 61270 11838 61276 11902
rect 61064 11832 61276 11838
rect 63648 12038 63996 12044
rect 63648 11974 63926 12038
rect 63990 11974 63996 12038
rect 63648 11968 63996 11974
rect 66096 12038 66444 12044
rect 66096 11974 66374 12038
rect 66438 11974 66444 12038
rect 66096 11968 66444 11974
rect 68544 12038 68892 12044
rect 68544 11974 68686 12038
rect 68750 11974 68892 12038
rect 63648 11908 63860 11968
rect 66096 11908 66308 11968
rect 63648 11902 66308 11908
rect 63648 11838 63790 11902
rect 63854 11838 66102 11902
rect 66166 11838 66308 11902
rect 63648 11832 66308 11838
rect 68544 11902 68892 11974
rect 68544 11838 68822 11902
rect 68886 11838 68892 11902
rect 68544 11832 68892 11838
rect 71128 12038 71476 12044
rect 71128 11974 71406 12038
rect 71470 11974 71476 12038
rect 71128 11968 71476 11974
rect 73576 12038 73924 12044
rect 73576 11974 73854 12038
rect 73918 11974 73924 12038
rect 73576 11968 73924 11974
rect 76024 12038 76508 12044
rect 76024 11974 76438 12038
rect 76502 11974 76508 12038
rect 76024 11968 76508 11974
rect 78608 12038 78956 12044
rect 78608 11974 78886 12038
rect 78950 11974 78956 12038
rect 78608 11968 78956 11974
rect 81056 12038 81404 12044
rect 81056 11974 81334 12038
rect 81398 11974 81404 12038
rect 81056 11968 81404 11974
rect 83504 12038 83988 12044
rect 83504 11974 83918 12038
rect 83982 11974 83988 12038
rect 83504 11968 83988 11974
rect 86088 12038 86436 12044
rect 86088 11974 86366 12038
rect 86430 11974 86436 12038
rect 86088 11968 86436 11974
rect 88536 12038 88884 12044
rect 88536 11974 88814 12038
rect 88878 11974 88884 12038
rect 88536 11968 88884 11974
rect 91120 12038 91468 12044
rect 91120 11974 91398 12038
rect 91462 11974 91468 12038
rect 91120 11968 91468 11974
rect 93568 12038 93916 12044
rect 93568 11974 93846 12038
rect 93910 11974 93916 12038
rect 93568 11968 93916 11974
rect 96016 12038 96364 12044
rect 96016 11974 96294 12038
rect 96358 11974 96364 12038
rect 96016 11968 96364 11974
rect 98600 12038 98948 12044
rect 98600 11974 98878 12038
rect 98942 11974 98948 12038
rect 98600 11968 98948 11974
rect 101048 12038 101396 12044
rect 101048 11974 101326 12038
rect 101390 11974 101396 12038
rect 101048 11968 101396 11974
rect 103496 12038 103708 12044
rect 103496 11974 103638 12038
rect 103702 11974 103708 12038
rect 71128 11902 71340 11968
rect 71128 11838 71270 11902
rect 71334 11838 71340 11902
rect 71128 11832 71340 11838
rect 73576 11902 73788 11968
rect 73576 11838 73718 11902
rect 73782 11838 73788 11902
rect 73576 11832 73788 11838
rect 76024 11902 76372 11968
rect 76024 11838 76302 11902
rect 76366 11838 76372 11902
rect 76024 11832 76372 11838
rect 78608 11908 78820 11968
rect 81056 11908 81268 11968
rect 83504 11908 83852 11968
rect 78608 11902 83852 11908
rect 78608 11838 78750 11902
rect 78814 11838 81198 11902
rect 81262 11838 83782 11902
rect 83846 11838 83852 11902
rect 78608 11832 83852 11838
rect 86088 11902 86300 11968
rect 86088 11838 86230 11902
rect 86294 11838 86300 11902
rect 86088 11832 86300 11838
rect 88536 11908 88748 11968
rect 88536 11902 88884 11908
rect 88536 11838 88814 11902
rect 88878 11838 88884 11902
rect 88536 11832 88884 11838
rect 91120 11902 91332 11968
rect 91120 11838 91126 11902
rect 91190 11838 91332 11902
rect 91120 11832 91332 11838
rect 93568 11902 93780 11968
rect 93568 11838 93574 11902
rect 93638 11838 93780 11902
rect 93568 11832 93780 11838
rect 96016 11902 96228 11968
rect 96016 11838 96158 11902
rect 96222 11838 96228 11902
rect 96016 11832 96228 11838
rect 98600 11902 98812 11968
rect 98600 11838 98742 11902
rect 98806 11838 98812 11902
rect 98600 11832 98812 11838
rect 101048 11902 101260 11968
rect 101048 11838 101190 11902
rect 101254 11838 101260 11902
rect 101048 11832 101260 11838
rect 103496 11902 103708 11974
rect 103496 11838 103638 11902
rect 103702 11838 103708 11902
rect 103496 11832 103708 11838
rect 106080 12038 106428 12044
rect 106080 11974 106358 12038
rect 106422 11974 106428 12038
rect 106080 11968 106428 11974
rect 121582 12027 121648 12030
rect 122320 12027 122386 12030
rect 121582 12025 122386 12027
rect 121582 11969 121587 12025
rect 121643 11969 122325 12025
rect 122381 11969 122386 12025
rect 106080 11902 106292 11968
rect 121582 11967 122386 11969
rect 121582 11964 121648 11967
rect 122320 11964 122386 11967
rect 106080 11838 106222 11902
rect 106286 11838 106292 11902
rect 106080 11832 106292 11838
rect 123216 11954 123428 12044
rect 134776 11968 134988 12112
rect 123216 11902 123270 11954
rect 123216 11838 123222 11902
rect 123326 11898 123428 11954
rect 123286 11838 123428 11898
rect 123216 11832 123428 11838
rect 14552 11702 14558 11766
rect 14622 11702 14764 11766
rect 14552 11696 14764 11702
rect 20128 11766 21564 11772
rect 20128 11702 20270 11766
rect 20334 11702 21564 11766
rect 20128 11696 21564 11702
rect 20128 11560 20340 11696
rect 21216 11560 21564 11696
rect 28832 11766 29044 11772
rect 28832 11702 28838 11766
rect 28902 11702 29044 11766
rect 28832 11560 29044 11702
rect 31280 11766 31492 11772
rect 33494 11766 33940 11772
rect 36214 11766 36524 11772
rect 38662 11766 38972 11772
rect 31280 11702 31422 11766
rect 31486 11702 31492 11766
rect 33456 11702 33462 11766
rect 33526 11702 33940 11766
rect 36176 11702 36182 11766
rect 36246 11702 36524 11766
rect 38624 11702 38630 11766
rect 38694 11702 38972 11766
rect 31280 11560 31492 11702
rect 33494 11696 33940 11702
rect 36214 11696 36524 11702
rect 38662 11696 38972 11702
rect 33728 11560 33940 11696
rect 28832 11500 28908 11560
rect 31280 11500 31356 11560
rect 33864 11500 33940 11560
rect 36312 11560 36524 11696
rect 38760 11560 38972 11696
rect 41208 11766 41556 11772
rect 41208 11702 41486 11766
rect 41550 11702 41556 11766
rect 41208 11560 41556 11702
rect 43792 11560 44004 11772
rect 46240 11766 46550 11772
rect 48688 11766 49036 11772
rect 46240 11702 46518 11766
rect 46582 11702 46588 11766
rect 48688 11702 48830 11766
rect 48894 11702 49036 11766
rect 46240 11696 46550 11702
rect 46240 11560 46452 11696
rect 48688 11560 49036 11702
rect 51272 11766 51484 11772
rect 51272 11702 51278 11766
rect 51342 11702 51484 11766
rect 51272 11560 51484 11702
rect 53720 11766 54030 11772
rect 56168 11766 56516 11772
rect 53720 11702 53998 11766
rect 54062 11702 54068 11766
rect 56168 11702 56446 11766
rect 56510 11702 56516 11766
rect 53720 11696 54030 11702
rect 53720 11560 53932 11696
rect 56168 11560 56516 11702
rect 58752 11766 59062 11772
rect 61200 11766 61412 11772
rect 63686 11766 63996 11772
rect 58752 11702 59030 11766
rect 59094 11702 59100 11766
rect 61200 11702 61342 11766
rect 61406 11702 61412 11766
rect 63648 11702 63654 11766
rect 63718 11702 63996 11766
rect 58752 11696 59062 11702
rect 58752 11560 58964 11696
rect 61200 11560 61412 11702
rect 63686 11696 63996 11702
rect 63784 11560 63996 11696
rect 66232 11766 66444 11772
rect 68582 11766 68892 11772
rect 66232 11702 66238 11766
rect 66302 11702 66444 11766
rect 68544 11702 68550 11766
rect 68614 11702 68892 11766
rect 66232 11560 66444 11702
rect 68582 11696 68892 11702
rect 68680 11560 68892 11696
rect 71264 11766 71574 11772
rect 71264 11702 71542 11766
rect 71606 11702 71612 11766
rect 71264 11696 71574 11702
rect 71264 11560 71476 11696
rect 73712 11560 73924 11772
rect 76160 11766 76372 11772
rect 78646 11766 78956 11772
rect 81094 11766 81404 11772
rect 76160 11702 76166 11766
rect 76230 11702 76372 11766
rect 78608 11702 78614 11766
rect 78678 11702 78956 11766
rect 81056 11702 81062 11766
rect 81126 11702 81404 11766
rect 76160 11560 76372 11702
rect 78646 11696 78956 11702
rect 81094 11696 81404 11702
rect 78744 11560 78956 11696
rect 81192 11560 81404 11696
rect 83640 11766 84086 11772
rect 86224 11766 86534 11772
rect 88672 11766 88982 11772
rect 91120 11766 91468 11772
rect 83640 11702 84054 11766
rect 84118 11702 84124 11766
rect 86224 11702 86502 11766
rect 86566 11702 86572 11766
rect 88672 11702 88950 11766
rect 89014 11702 89020 11766
rect 91120 11702 91262 11766
rect 91326 11702 91468 11766
rect 83640 11696 84086 11702
rect 86224 11696 86534 11702
rect 88672 11696 88982 11702
rect 83640 11560 83988 11696
rect 86224 11560 86436 11696
rect 88672 11560 88884 11696
rect 91120 11560 91468 11702
rect 93704 11560 93916 11772
rect 96054 11766 96364 11772
rect 96016 11702 96022 11766
rect 96086 11702 96364 11766
rect 96054 11696 96364 11702
rect 96152 11560 96364 11696
rect 98600 11766 99046 11772
rect 101184 11766 101494 11772
rect 103632 11766 103844 11772
rect 106118 11766 106428 11772
rect 98600 11702 99014 11766
rect 99078 11702 99084 11766
rect 101184 11702 101462 11766
rect 101526 11702 101532 11766
rect 103632 11702 103774 11766
rect 103838 11702 103844 11766
rect 106080 11702 106086 11766
rect 106150 11702 106428 11766
rect 98600 11696 99046 11702
rect 101184 11696 101494 11702
rect 98600 11560 98948 11696
rect 101184 11560 101396 11696
rect 103632 11560 103844 11702
rect 106118 11696 106428 11702
rect 106216 11560 106428 11696
rect 36312 11500 36388 11560
rect 38760 11500 38836 11560
rect 28696 11364 28908 11500
rect 28190 11358 28908 11364
rect 28152 11294 28158 11358
rect 28222 11294 28908 11358
rect 28190 11288 28908 11294
rect 31144 11288 31356 11500
rect 33592 11288 33940 11500
rect 36176 11288 36388 11500
rect 38624 11288 38836 11500
rect 41208 11500 41284 11560
rect 43792 11500 43868 11560
rect 46240 11500 46316 11560
rect 48824 11500 48900 11560
rect 51272 11500 51348 11560
rect 53720 11500 53796 11560
rect 41208 11288 41420 11500
rect 43384 11494 43868 11500
rect 43384 11430 43390 11494
rect 43454 11430 43868 11494
rect 43384 11424 43868 11430
rect 43656 11288 43868 11424
rect 46104 11288 46316 11500
rect 48688 11288 48900 11500
rect 51136 11288 51348 11500
rect 53584 11288 53796 11500
rect 56168 11500 56244 11560
rect 58752 11500 58828 11560
rect 61200 11500 61276 11560
rect 63784 11500 63860 11560
rect 66232 11500 66308 11560
rect 68680 11500 68756 11560
rect 71264 11500 71340 11560
rect 73712 11500 73788 11560
rect 76160 11500 76236 11560
rect 78744 11500 78820 11560
rect 81192 11500 81268 11560
rect 56168 11288 56380 11500
rect 58616 11288 58828 11500
rect 61064 11288 61412 11500
rect 63648 11288 63860 11500
rect 66096 11288 66308 11500
rect 68544 11288 68892 11500
rect 71128 11288 71340 11500
rect 73304 11494 73788 11500
rect 73304 11430 73310 11494
rect 73374 11430 73788 11494
rect 73304 11424 73788 11430
rect 73576 11288 73788 11424
rect 76024 11288 76372 11500
rect 78608 11288 78820 11500
rect 81056 11288 81268 11500
rect 83640 11500 83716 11560
rect 86224 11500 86300 11560
rect 88672 11500 88748 11560
rect 91256 11500 91332 11560
rect 93704 11500 93780 11560
rect 96152 11500 96228 11560
rect 83640 11288 83852 11500
rect 86088 11288 86300 11500
rect 88536 11288 88748 11500
rect 91120 11288 91332 11500
rect 93568 11494 93780 11500
rect 93568 11430 93710 11494
rect 93774 11430 93780 11494
rect 93568 11288 93780 11430
rect 96016 11288 96228 11500
rect 98600 11500 98676 11560
rect 101184 11500 101260 11560
rect 103632 11500 103708 11560
rect 106216 11500 106292 11560
rect 98600 11288 98812 11500
rect 101048 11288 101260 11500
rect 103496 11288 103844 11500
rect 106080 11364 106292 11500
rect 122808 11494 123020 11500
rect 122808 11430 122814 11494
rect 122878 11430 123020 11494
rect 106080 11358 108468 11364
rect 106080 11294 108398 11358
rect 108462 11294 108468 11358
rect 106080 11288 108468 11294
rect 122808 11288 123020 11430
rect 28598 11086 31356 11092
rect 28560 11022 28566 11086
rect 28630 11022 28702 11086
rect 28766 11022 31150 11086
rect 31214 11022 31356 11086
rect 28598 11016 31356 11022
rect 33728 11086 36388 11092
rect 33728 11022 33870 11086
rect 33934 11022 36318 11086
rect 36382 11022 36388 11086
rect 33728 11016 36388 11022
rect 38624 11086 38836 11092
rect 38624 11022 38766 11086
rect 38830 11022 38836 11086
rect 38624 11016 38836 11022
rect 41208 11086 41420 11092
rect 41208 11022 41350 11086
rect 41414 11022 41420 11086
rect 41208 11016 41420 11022
rect 43656 11086 46452 11092
rect 43656 11022 43798 11086
rect 43862 11022 46246 11086
rect 46310 11022 46452 11086
rect 43656 11016 46452 11022
rect 48688 11086 53932 11092
rect 48688 11022 48694 11086
rect 48758 11022 51142 11086
rect 51206 11022 53862 11086
rect 53926 11022 53932 11086
rect 48688 11016 53932 11022
rect 56168 11086 56380 11092
rect 56168 11022 56310 11086
rect 56374 11022 56380 11086
rect 56168 11016 56380 11022
rect 58616 11086 58828 11092
rect 58616 11022 58758 11086
rect 58822 11022 58828 11086
rect 58616 11016 58828 11022
rect 61064 11086 61412 11092
rect 61064 11022 61206 11086
rect 61270 11022 61412 11086
rect 61064 11016 61412 11022
rect 63648 11086 63860 11092
rect 63648 11022 63790 11086
rect 63854 11022 63860 11086
rect 63648 11016 63860 11022
rect 66096 11086 73788 11092
rect 66096 11022 66102 11086
rect 66166 11022 68822 11086
rect 68886 11022 71270 11086
rect 71334 11022 73718 11086
rect 73782 11022 73788 11086
rect 66096 11016 73788 11022
rect 76160 11086 78820 11092
rect 76160 11022 76302 11086
rect 76366 11022 78750 11086
rect 78814 11022 78820 11086
rect 76160 11016 78820 11022
rect 81056 11086 81268 11092
rect 81056 11022 81198 11086
rect 81262 11022 81268 11086
rect 81056 11016 81268 11022
rect 83640 11086 83852 11092
rect 83640 11022 83782 11086
rect 83846 11022 83852 11086
rect 83640 11016 83852 11022
rect 86088 11086 96364 11092
rect 86088 11022 86230 11086
rect 86294 11022 88814 11086
rect 88878 11022 91126 11086
rect 91190 11022 93574 11086
rect 93638 11022 96158 11086
rect 96222 11022 96364 11086
rect 86088 11016 96364 11022
rect 98600 11086 98812 11092
rect 98600 11022 98742 11086
rect 98806 11022 98812 11086
rect 98600 11016 98812 11022
rect 101048 11086 101260 11092
rect 101048 11022 101190 11086
rect 101254 11022 101260 11086
rect 101048 11016 101260 11022
rect 103496 11086 103844 11092
rect 103496 11022 103638 11086
rect 103702 11022 103844 11086
rect 103496 11016 103844 11022
rect 106080 11086 108332 11092
rect 106080 11022 106222 11086
rect 106286 11022 108262 11086
rect 108326 11022 108332 11086
rect 106080 11016 108332 11022
rect 28746 10985 28844 11016
rect 31242 10985 31340 11016
rect 33738 10985 33836 11016
rect 36234 10985 36332 11016
rect 38730 10985 38828 11016
rect 41226 10985 41324 11016
rect 43722 10985 43820 11016
rect 46218 10985 46316 11016
rect 48714 10985 48812 11016
rect 51210 10985 51308 11016
rect 53706 10985 53804 11016
rect 56202 10985 56300 11016
rect 58698 10985 58796 11016
rect 61194 10985 61292 11016
rect 63690 10985 63788 11016
rect 66186 10985 66284 11016
rect 68682 10985 68780 11016
rect 71178 10985 71276 11016
rect 73674 10985 73772 11016
rect 76170 10985 76268 11016
rect 78666 10985 78764 11016
rect 81162 10985 81260 11016
rect 83658 10985 83756 11016
rect 86154 10985 86252 11016
rect 88650 10985 88748 11016
rect 91146 10985 91244 11016
rect 93642 10985 93740 11016
rect 96138 10985 96236 11016
rect 98634 10985 98732 11016
rect 101130 10985 101228 11016
rect 103626 10985 103724 11016
rect 106122 10985 106220 11016
rect 123216 10826 123428 10956
rect 123216 10770 123270 10826
rect 123326 10814 123428 10826
rect 123326 10770 123358 10814
rect 121502 10757 121568 10760
rect 122320 10757 122386 10760
rect 121502 10755 122386 10757
rect 121502 10699 121507 10755
rect 121563 10699 122325 10755
rect 122381 10699 122386 10755
rect 123216 10750 123358 10770
rect 123422 10750 123428 10814
rect 123216 10744 123428 10750
rect 121502 10697 122386 10699
rect 121502 10694 121568 10697
rect 122320 10694 122386 10697
rect 27064 10678 28636 10684
rect 27064 10614 28566 10678
rect 28630 10614 28636 10678
rect 27064 10608 28636 10614
rect 108256 10678 108468 10684
rect 108256 10614 108262 10678
rect 108326 10614 108468 10678
rect 1224 10542 1980 10548
rect 1224 10478 1230 10542
rect 1294 10488 1980 10542
rect 1294 10478 1794 10488
rect 1224 10472 1794 10478
rect 1768 10432 1794 10472
rect 1850 10432 1980 10488
rect 1768 10336 1980 10432
rect 2448 10412 2796 10548
rect 2040 10336 2796 10412
rect 14552 10542 14764 10548
rect 14552 10478 14694 10542
rect 14758 10478 14764 10542
rect 14552 10406 14764 10478
rect 27064 10472 27276 10608
rect 108256 10472 108468 10614
rect 134776 10488 134988 10548
rect 14552 10342 14694 10406
rect 14758 10342 14764 10406
rect 14552 10336 14764 10342
rect 134776 10432 134844 10488
rect 134900 10432 134988 10488
rect 134776 10412 134988 10432
rect 134776 10406 135396 10412
rect 134776 10342 135326 10406
rect 135390 10342 135396 10406
rect 134776 10336 135396 10342
rect 2040 10276 2116 10336
rect 544 10270 2116 10276
rect 544 10206 550 10270
rect 614 10206 2116 10270
rect 544 10200 2116 10206
rect 0 9928 2932 10004
rect 2720 9912 2932 9928
rect 2720 9856 2754 9912
rect 2810 9856 2932 9912
rect 2720 9792 2932 9856
rect 122808 9998 123020 10004
rect 122808 9934 122950 9998
rect 123014 9934 123020 9998
rect 122808 9792 123020 9934
rect 27064 9590 28228 9596
rect 27064 9526 28158 9590
rect 28222 9526 28228 9590
rect 27064 9520 28228 9526
rect 108256 9590 108468 9596
rect 108256 9526 108398 9590
rect 108462 9526 108468 9590
rect 27064 9384 27276 9520
rect 108256 9384 108468 9526
rect 2448 8976 2796 9188
rect 14552 9182 14764 9188
rect 14552 9118 14558 9182
rect 14622 9118 14764 9182
rect 14552 9052 14764 9118
rect 14552 9046 16396 9052
rect 14552 8982 16326 9046
rect 16390 8982 16396 9046
rect 14552 8976 16396 8982
rect 2448 8916 2524 8976
rect 1768 8840 2524 8916
rect 1768 8808 1980 8840
rect 1768 8780 1794 8808
rect 1224 8774 1794 8780
rect 1224 8710 1230 8774
rect 1294 8752 1794 8774
rect 1850 8752 1980 8808
rect 1294 8710 1980 8752
rect 1224 8704 1980 8710
rect 134776 8808 134988 8916
rect 134776 8752 134844 8808
rect 134900 8780 134988 8808
rect 134900 8774 135396 8780
rect 134900 8752 135326 8774
rect 134776 8710 135326 8752
rect 135390 8710 135396 8774
rect 134776 8704 135396 8710
rect 0 8317 6060 8372
rect 0 8296 5975 8317
rect 5848 8261 5975 8296
rect 6031 8261 6060 8317
rect 2720 8212 2932 8236
rect 2720 8156 2754 8212
rect 2810 8156 2932 8212
rect 5848 8160 6060 8261
rect 2720 8100 2932 8156
rect 0 8024 2932 8100
rect 544 7686 2796 7692
rect 544 7622 550 7686
rect 614 7622 2796 7686
rect 544 7616 2796 7622
rect 2448 7480 2796 7616
rect 14552 7686 14764 7692
rect 14552 7622 14694 7686
rect 14758 7622 14764 7686
rect 14552 7480 14764 7622
rect 1224 7278 1980 7284
rect 1224 7214 1230 7278
rect 1294 7214 1980 7278
rect 1224 7208 1980 7214
rect 1768 7128 1980 7208
rect 1768 7072 1794 7128
rect 1850 7072 1980 7128
rect 1768 6936 1980 7072
rect 134776 7148 134988 7284
rect 134776 7142 135396 7148
rect 134776 7128 135326 7142
rect 134776 7072 134844 7128
rect 134900 7078 135326 7128
rect 135390 7078 135396 7142
rect 134900 7072 135396 7078
rect 134776 6936 134988 7072
rect 1224 5510 1980 5516
rect 1224 5446 1230 5510
rect 1294 5448 1980 5510
rect 1294 5446 1794 5448
rect 1224 5440 1794 5446
rect 1768 5392 1794 5440
rect 1850 5392 1980 5448
rect 1768 5304 1980 5392
rect 134776 5448 134988 5516
rect 134776 5392 134844 5448
rect 134900 5392 134988 5448
rect 134776 5380 134988 5392
rect 134776 5374 135396 5380
rect 134776 5310 135326 5374
rect 135390 5310 135396 5374
rect 134776 5304 135396 5310
rect 1224 3878 1980 3884
rect 1224 3814 1230 3878
rect 1294 3814 1980 3878
rect 1224 3808 1980 3814
rect 1768 3768 1980 3808
rect 1768 3712 1794 3768
rect 1850 3712 1980 3768
rect 1768 3672 1980 3712
rect 16320 3878 17756 3884
rect 16320 3814 16326 3878
rect 16390 3814 17756 3878
rect 16320 3808 17756 3814
rect 16320 3672 16532 3808
rect 17544 3748 17756 3808
rect 18632 3748 18844 3884
rect 19856 3808 21292 3884
rect 19856 3748 20068 3808
rect 20944 3748 21292 3808
rect 22168 3748 22380 3884
rect 23392 3808 25916 3884
rect 23392 3748 23604 3808
rect 17544 3742 20340 3748
rect 17544 3678 20270 3742
rect 20334 3678 20340 3742
rect 17544 3672 20340 3678
rect 20944 3672 23604 3748
rect 24480 3672 24692 3808
rect 25704 3748 25916 3808
rect 26792 3748 27140 3884
rect 28016 3808 29452 3884
rect 28016 3748 28228 3808
rect 25704 3672 28228 3748
rect 29240 3748 29452 3808
rect 30328 3748 30540 3884
rect 31552 3808 34076 3884
rect 31552 3748 31764 3808
rect 29240 3672 31764 3748
rect 32640 3672 32852 3808
rect 33864 3748 34076 3808
rect 34952 3808 37612 3884
rect 34952 3748 35300 3808
rect 33864 3672 35300 3748
rect 36176 3672 36388 3808
rect 37400 3748 37612 3808
rect 38488 3748 38700 3884
rect 39712 3808 41148 3884
rect 39712 3748 39924 3808
rect 37400 3672 39924 3748
rect 40800 3748 41148 3808
rect 42024 3748 42236 3884
rect 43248 3808 45772 3884
rect 43248 3748 43460 3808
rect 40800 3672 43460 3748
rect 44336 3672 44548 3808
rect 45560 3748 45772 3808
rect 46648 3748 46996 3884
rect 47872 3808 49308 3884
rect 47872 3748 48084 3808
rect 45560 3672 48084 3748
rect 49096 3748 49308 3808
rect 50184 3748 50396 3884
rect 51408 3808 53932 3884
rect 51408 3748 51620 3808
rect 49096 3672 51620 3748
rect 52496 3672 52708 3808
rect 53720 3748 53932 3808
rect 54808 3748 55156 3884
rect 56032 3808 57468 3884
rect 56032 3748 56244 3808
rect 53720 3672 56244 3748
rect 57256 3748 57468 3808
rect 58344 3748 58556 3884
rect 59568 3748 59780 3884
rect 57256 3672 59780 3748
rect 134776 3768 134988 3884
rect 134776 3712 134844 3768
rect 134900 3748 134988 3768
rect 134900 3742 135396 3748
rect 134900 3712 135326 3742
rect 134776 3678 135326 3712
rect 135390 3678 135396 3742
rect 134776 3672 135396 3678
rect 15912 2988 16124 3068
rect 15912 2932 16004 2988
rect 16060 2932 16124 2988
rect 15912 2926 16124 2932
rect 15912 2862 16054 2926
rect 16118 2862 16124 2926
rect 15912 2856 16124 2862
rect 17136 2988 17348 3068
rect 17136 2932 17172 2988
rect 17228 2932 17348 2988
rect 17136 2926 17348 2932
rect 17136 2862 17142 2926
rect 17206 2862 17348 2926
rect 17136 2856 17348 2862
rect 18224 2988 18436 3068
rect 19584 3009 19660 3068
rect 20672 3009 20884 3068
rect 21896 3009 21972 3068
rect 18224 2932 18340 2988
rect 18396 2932 18436 2988
rect 19487 2988 19660 3009
rect 19487 2932 19508 2988
rect 19564 2932 19660 2988
rect 20655 2988 20884 3009
rect 20655 2932 20676 2988
rect 20732 2932 20884 2988
rect 21823 2988 21972 3009
rect 21823 2932 21844 2988
rect 21900 2932 21972 2988
rect 18224 2926 18436 2932
rect 18224 2862 18230 2926
rect 18294 2862 18436 2926
rect 18224 2856 18436 2862
rect 19448 2926 19660 2932
rect 19448 2862 19590 2926
rect 19654 2862 19660 2926
rect 19448 2856 19660 2862
rect 20536 2926 20884 2932
rect 20536 2862 20542 2926
rect 20606 2862 20884 2926
rect 20536 2856 20884 2862
rect 21760 2926 21972 2932
rect 21760 2862 21766 2926
rect 21830 2862 21972 2926
rect 21760 2856 21972 2862
rect 22984 2988 23196 3068
rect 24208 3009 24284 3068
rect 22984 2932 23012 2988
rect 23068 2932 23196 2988
rect 24159 2988 24284 3009
rect 24159 2932 24180 2988
rect 24236 2932 24284 2988
rect 22984 2926 23196 2932
rect 22984 2862 23126 2926
rect 23190 2862 23196 2926
rect 22984 2856 23196 2862
rect 24072 2926 24284 2932
rect 24072 2862 24214 2926
rect 24278 2862 24284 2926
rect 24072 2856 24284 2862
rect 25296 2988 25508 3068
rect 26520 3009 26596 3068
rect 27744 3009 27820 3068
rect 28832 3009 29044 3068
rect 30056 3009 30132 3068
rect 25296 2932 25348 2988
rect 25404 2932 25508 2988
rect 26495 2988 26596 3009
rect 26495 2932 26516 2988
rect 26572 2932 26596 2988
rect 27663 2988 27820 3009
rect 27663 2932 27684 2988
rect 27740 2932 27820 2988
rect 28831 2988 29044 3009
rect 28831 2932 28852 2988
rect 28908 2932 29044 2988
rect 29999 2988 30132 3009
rect 29999 2932 30020 2988
rect 30076 2932 30132 2988
rect 25296 2926 25508 2932
rect 25296 2862 25438 2926
rect 25502 2862 25508 2926
rect 25296 2856 25508 2862
rect 26384 2926 26596 2932
rect 26384 2862 26526 2926
rect 26590 2862 26596 2926
rect 26384 2856 26596 2862
rect 27608 2926 27820 2932
rect 27608 2862 27614 2926
rect 27678 2862 27820 2926
rect 27608 2856 27820 2862
rect 28696 2926 29044 2932
rect 28696 2862 28702 2926
rect 28766 2862 29044 2926
rect 28696 2856 29044 2862
rect 29920 2926 30132 2932
rect 29920 2862 30062 2926
rect 30126 2862 30132 2926
rect 29920 2856 30132 2862
rect 31144 2988 31356 3068
rect 32368 3009 32444 3068
rect 33592 3009 33668 3068
rect 34680 3009 34892 3068
rect 35904 3009 35980 3068
rect 31144 2932 31188 2988
rect 31244 2932 31356 2988
rect 32335 2988 32444 3009
rect 32335 2932 32356 2988
rect 32412 2932 32444 2988
rect 33503 2988 33668 3009
rect 33503 2932 33524 2988
rect 33580 2932 33668 2988
rect 34671 2988 34892 3009
rect 34671 2932 34692 2988
rect 34748 2932 34892 2988
rect 35839 2988 35980 3009
rect 35839 2932 35860 2988
rect 35916 2932 35980 2988
rect 31144 2926 31356 2932
rect 31144 2862 31286 2926
rect 31350 2862 31356 2926
rect 31144 2856 31356 2862
rect 32232 2926 32444 2932
rect 32232 2862 32374 2926
rect 32438 2862 32444 2926
rect 32232 2856 32444 2862
rect 33456 2926 33668 2932
rect 33456 2862 33462 2926
rect 33526 2862 33668 2926
rect 33456 2856 33668 2862
rect 34544 2926 34892 2932
rect 34544 2862 34550 2926
rect 34614 2862 34892 2926
rect 34544 2856 34892 2862
rect 35768 2926 35980 2932
rect 35768 2862 35910 2926
rect 35974 2862 35980 2926
rect 35768 2856 35980 2862
rect 36992 2988 37204 3068
rect 38216 3009 38292 3068
rect 39440 3009 39516 3068
rect 40528 3009 40740 3068
rect 41752 3009 41828 3068
rect 36992 2932 37028 2988
rect 37084 2932 37204 2988
rect 38175 2988 38292 3009
rect 38175 2932 38196 2988
rect 38252 2932 38292 2988
rect 39343 2988 39516 3009
rect 39343 2932 39364 2988
rect 39420 2932 39516 2988
rect 40511 2988 40740 3009
rect 40511 2932 40532 2988
rect 40588 2932 40740 2988
rect 41679 2988 41828 3009
rect 41679 2932 41700 2988
rect 41756 2932 41828 2988
rect 36992 2926 37204 2932
rect 36992 2862 36998 2926
rect 37062 2862 37204 2926
rect 36992 2856 37204 2862
rect 38080 2926 38292 2932
rect 38080 2862 38086 2926
rect 38150 2862 38292 2926
rect 38080 2856 38292 2862
rect 39304 2926 39516 2932
rect 39304 2862 39446 2926
rect 39510 2862 39516 2926
rect 39304 2856 39516 2862
rect 40392 2926 40740 2932
rect 40392 2862 40670 2926
rect 40734 2862 40740 2926
rect 40392 2856 40740 2862
rect 41616 2926 41828 2932
rect 41616 2862 41758 2926
rect 41822 2862 41828 2926
rect 41616 2856 41828 2862
rect 42840 2988 43052 3068
rect 44064 3009 44140 3068
rect 42840 2932 42868 2988
rect 42924 2932 43052 2988
rect 44015 2988 44140 3009
rect 44015 2932 44036 2988
rect 44092 2932 44140 2988
rect 42840 2926 43052 2932
rect 42840 2862 42846 2926
rect 42910 2862 43052 2926
rect 42840 2856 43052 2862
rect 43928 2926 44140 2932
rect 43928 2862 43934 2926
rect 43998 2862 44140 2926
rect 43928 2856 44140 2862
rect 45152 2988 45364 3068
rect 46376 3009 46452 3068
rect 47600 3009 47676 3068
rect 48688 3009 48900 3068
rect 49912 3009 49988 3068
rect 45152 2932 45204 2988
rect 45260 2932 45364 2988
rect 46351 2988 46452 3009
rect 46351 2932 46372 2988
rect 46428 2932 46452 2988
rect 47519 2988 47676 3009
rect 47519 2932 47540 2988
rect 47596 2932 47676 2988
rect 48687 2988 48900 3009
rect 48687 2932 48708 2988
rect 48764 2932 48900 2988
rect 49855 2988 49988 3009
rect 49855 2932 49876 2988
rect 49932 2932 49988 2988
rect 45152 2926 45364 2932
rect 45152 2862 45294 2926
rect 45358 2862 45364 2926
rect 45152 2856 45364 2862
rect 46240 2926 46452 2932
rect 46240 2862 46382 2926
rect 46446 2862 46452 2926
rect 46240 2856 46452 2862
rect 47464 2926 47676 2932
rect 47464 2862 47606 2926
rect 47670 2862 47676 2926
rect 47464 2856 47676 2862
rect 48552 2926 48900 2932
rect 48552 2862 48694 2926
rect 48758 2862 48900 2926
rect 48552 2856 48900 2862
rect 49776 2926 49988 2932
rect 49776 2862 49782 2926
rect 49846 2862 49988 2926
rect 49776 2856 49988 2862
rect 51000 2988 51212 3068
rect 52224 3009 52300 3068
rect 53448 3009 53524 3068
rect 54536 3009 54748 3068
rect 55760 3009 55836 3068
rect 51000 2932 51044 2988
rect 51100 2932 51212 2988
rect 52191 2988 52300 3009
rect 52191 2932 52212 2988
rect 52268 2932 52300 2988
rect 53359 2988 53524 3009
rect 53359 2932 53380 2988
rect 53436 2932 53524 2988
rect 54527 2988 54748 3009
rect 54527 2932 54548 2988
rect 54604 2932 54748 2988
rect 55695 2988 55836 3009
rect 55695 2932 55716 2988
rect 55772 2932 55836 2988
rect 51000 2926 51212 2932
rect 51000 2862 51142 2926
rect 51206 2862 51212 2926
rect 51000 2856 51212 2862
rect 52088 2926 52300 2932
rect 52088 2862 52230 2926
rect 52294 2862 52300 2926
rect 52088 2856 52300 2862
rect 53312 2926 53524 2932
rect 53312 2862 53318 2926
rect 53382 2862 53524 2926
rect 53312 2856 53524 2862
rect 54400 2926 54748 2932
rect 54400 2862 54406 2926
rect 54470 2862 54748 2926
rect 54400 2856 54748 2862
rect 55624 2926 55836 2932
rect 55624 2862 55766 2926
rect 55830 2862 55836 2926
rect 55624 2856 55836 2862
rect 56848 2988 57060 3068
rect 58072 3009 58148 3068
rect 59296 3009 59372 3068
rect 56848 2932 56884 2988
rect 56940 2932 57060 2988
rect 58031 2988 58148 3009
rect 58031 2932 58052 2988
rect 58108 2932 58148 2988
rect 59199 2988 59372 3009
rect 59199 2932 59220 2988
rect 59276 2932 59372 2988
rect 56848 2926 57060 2932
rect 56848 2862 56990 2926
rect 57054 2862 57060 2926
rect 56848 2856 57060 2862
rect 57936 2926 58148 2932
rect 57936 2862 58078 2926
rect 58142 2862 58148 2926
rect 57936 2856 58148 2862
rect 59160 2926 59372 2932
rect 59160 2862 59166 2926
rect 59230 2862 59372 2926
rect 59160 2856 59372 2862
rect 14745 2734 14811 2737
rect 14745 2732 17030 2734
rect 14745 2676 14750 2732
rect 14806 2676 17030 2732
rect 14745 2674 17030 2676
rect 14745 2671 14811 2674
rect 16320 2448 17756 2524
rect 16320 2312 16532 2448
rect 17544 2388 17756 2448
rect 18632 2388 18844 2524
rect 19856 2448 22380 2524
rect 19856 2388 20068 2448
rect 17544 2312 20068 2388
rect 20944 2312 21292 2448
rect 22168 2388 22380 2448
rect 23392 2448 25916 2524
rect 23392 2388 23604 2448
rect 22168 2312 23604 2388
rect 24480 2312 24692 2448
rect 25704 2388 25916 2448
rect 26792 2388 27140 2524
rect 28016 2448 29452 2524
rect 28016 2388 28228 2448
rect 25704 2312 28228 2388
rect 29240 2388 29452 2448
rect 30328 2388 30540 2524
rect 31552 2448 34076 2524
rect 31552 2388 31764 2448
rect 29240 2312 31764 2388
rect 32640 2312 32852 2448
rect 33864 2388 34076 2448
rect 34952 2388 35300 2524
rect 36176 2448 37612 2524
rect 36176 2388 36388 2448
rect 33864 2312 36388 2388
rect 37400 2388 37612 2448
rect 38488 2388 38700 2524
rect 39712 2448 42236 2524
rect 39712 2388 39924 2448
rect 37400 2382 39924 2388
rect 37400 2318 39718 2382
rect 39782 2318 39924 2382
rect 37400 2312 39924 2318
rect 40800 2312 41148 2448
rect 42024 2388 42236 2448
rect 43248 2448 45772 2524
rect 43248 2388 43460 2448
rect 42024 2312 43460 2388
rect 44336 2312 44548 2448
rect 45560 2388 45772 2448
rect 46648 2388 46996 2524
rect 47872 2448 49308 2524
rect 47872 2388 48084 2448
rect 45560 2312 48084 2388
rect 49096 2388 49308 2448
rect 50184 2388 50396 2524
rect 51408 2448 53932 2524
rect 51408 2388 51620 2448
rect 49096 2312 51620 2388
rect 52496 2312 52708 2448
rect 53720 2388 53932 2448
rect 54808 2448 57468 2524
rect 54808 2388 55156 2448
rect 53720 2312 55156 2388
rect 56032 2312 56244 2448
rect 57256 2388 57468 2448
rect 58344 2388 58556 2524
rect 59568 2388 59780 2524
rect 57256 2312 59780 2388
rect 1768 2088 1980 2116
rect 1768 2032 1794 2088
rect 1850 2032 1980 2088
rect 1768 1980 1980 2032
rect 134776 2110 135396 2116
rect 134776 2088 135326 2110
rect 134776 2032 134844 2088
rect 134900 2046 135326 2088
rect 135390 2046 135396 2110
rect 134900 2040 135396 2046
rect 134900 2032 134988 2040
rect 1768 1904 2116 1980
rect 134776 1904 134988 2032
rect 2040 1844 2116 1904
rect 2040 1752 2252 1844
rect 2040 1702 2130 1752
rect 2040 1638 2046 1702
rect 2110 1696 2130 1702
rect 2186 1696 2252 1752
rect 2110 1638 2252 1696
rect 2040 1632 2252 1638
rect 3672 1752 4020 1844
rect 3672 1696 3810 1752
rect 3866 1702 4020 1752
rect 3672 1638 3814 1696
rect 3878 1638 4020 1702
rect 3672 1632 4020 1638
rect 5440 1752 5652 1844
rect 5440 1696 5490 1752
rect 5546 1702 5652 1752
rect 5546 1696 5582 1702
rect 5440 1638 5582 1696
rect 5646 1638 5652 1702
rect 5440 1632 5652 1638
rect 7072 1752 7284 1844
rect 7072 1702 7170 1752
rect 7072 1638 7078 1702
rect 7142 1696 7170 1702
rect 7226 1696 7284 1752
rect 7142 1638 7284 1696
rect 7072 1632 7284 1638
rect 8704 1752 9052 1844
rect 8704 1702 8850 1752
rect 8704 1638 8710 1702
rect 8774 1696 8850 1702
rect 8906 1696 9052 1752
rect 8774 1638 9052 1696
rect 8704 1632 9052 1638
rect 10472 1752 10684 1844
rect 10472 1702 10530 1752
rect 10472 1638 10478 1702
rect 10586 1696 10684 1752
rect 10542 1638 10684 1696
rect 10472 1632 10684 1638
rect 12104 1752 12316 1844
rect 12104 1702 12210 1752
rect 12104 1638 12110 1702
rect 12174 1696 12210 1702
rect 12266 1696 12316 1752
rect 12174 1638 12316 1696
rect 12104 1632 12316 1638
rect 13736 1752 14084 1844
rect 13736 1696 13890 1752
rect 13946 1702 14084 1752
rect 13946 1696 14014 1702
rect 13736 1638 14014 1696
rect 14078 1638 14084 1702
rect 13736 1632 14084 1638
rect 15504 1752 15716 1844
rect 15504 1702 15570 1752
rect 15504 1638 15510 1702
rect 15626 1696 15716 1752
rect 15574 1638 15716 1696
rect 15504 1632 15716 1638
rect 17136 1752 17348 1844
rect 17136 1696 17250 1752
rect 17306 1708 17348 1752
rect 18904 1752 19116 1844
rect 20302 1838 20748 1844
rect 20264 1774 20270 1838
rect 20334 1774 20748 1838
rect 20302 1768 20748 1774
rect 17306 1702 17484 1708
rect 17306 1696 17414 1702
rect 17136 1638 17414 1696
rect 17478 1638 17484 1702
rect 17136 1632 17484 1638
rect 18904 1696 18930 1752
rect 18986 1702 19116 1752
rect 18986 1696 19046 1702
rect 18904 1638 19046 1696
rect 19110 1638 19116 1702
rect 18904 1632 19116 1638
rect 20536 1752 20748 1768
rect 20536 1696 20610 1752
rect 20666 1708 20748 1752
rect 22168 1752 22380 1844
rect 20666 1702 20884 1708
rect 20666 1696 20814 1702
rect 20536 1638 20814 1696
rect 20878 1638 20884 1702
rect 20536 1632 20884 1638
rect 22168 1702 22290 1752
rect 22168 1638 22174 1702
rect 22238 1696 22290 1702
rect 22346 1696 22380 1752
rect 22238 1638 22380 1696
rect 22168 1632 22380 1638
rect 23936 1752 24148 1844
rect 23936 1702 23970 1752
rect 23936 1638 23942 1702
rect 24026 1696 24148 1752
rect 24006 1638 24148 1696
rect 23936 1632 24148 1638
rect 25568 1752 25780 1844
rect 25568 1696 25650 1752
rect 25706 1702 25780 1752
rect 25706 1696 25710 1702
rect 25568 1638 25710 1696
rect 25774 1638 25780 1702
rect 25568 1632 25780 1638
rect 27200 1752 27412 1844
rect 27200 1696 27330 1752
rect 27386 1702 27412 1752
rect 27200 1638 27342 1696
rect 27406 1638 27412 1702
rect 27200 1632 27412 1638
rect 28968 1752 29180 1844
rect 28968 1702 29010 1752
rect 28968 1638 28974 1702
rect 29066 1696 29180 1752
rect 30600 1752 30812 1844
rect 30600 1708 30690 1752
rect 29038 1638 29180 1696
rect 28968 1632 29180 1638
rect 30464 1702 30690 1708
rect 30464 1638 30470 1702
rect 30534 1696 30690 1702
rect 30746 1696 30812 1752
rect 32232 1752 32580 1844
rect 32232 1708 32370 1752
rect 30534 1638 30812 1696
rect 30464 1632 30812 1638
rect 32096 1702 32370 1708
rect 32096 1638 32102 1702
rect 32166 1696 32370 1702
rect 32426 1696 32580 1752
rect 32166 1638 32580 1696
rect 32096 1632 32580 1638
rect 34000 1752 34212 1844
rect 34000 1702 34050 1752
rect 34000 1638 34006 1702
rect 34106 1696 34212 1752
rect 34070 1638 34212 1696
rect 34000 1632 34212 1638
rect 35632 1752 35844 1844
rect 35632 1696 35730 1752
rect 35786 1702 35844 1752
rect 35632 1638 35774 1696
rect 35838 1638 35844 1702
rect 35632 1632 35844 1638
rect 37264 1752 37612 1844
rect 37264 1702 37410 1752
rect 37466 1702 37612 1752
rect 37264 1638 37406 1702
rect 37470 1638 37612 1702
rect 37264 1632 37612 1638
rect 39032 1752 39244 1844
rect 39032 1696 39090 1752
rect 39146 1702 39244 1752
rect 39146 1696 39174 1702
rect 39032 1638 39174 1696
rect 39238 1638 39244 1702
rect 39032 1632 39244 1638
rect 40664 1752 40876 1844
rect 40664 1696 40770 1752
rect 40826 1702 40876 1752
rect 40664 1638 40806 1696
rect 40870 1638 40876 1702
rect 40664 1632 40876 1638
rect 42296 1752 42644 1844
rect 42296 1702 42450 1752
rect 42296 1638 42438 1702
rect 42506 1696 42644 1752
rect 42502 1638 42644 1696
rect 42296 1632 42644 1638
rect 44064 1752 44276 1844
rect 44064 1696 44130 1752
rect 44186 1702 44276 1752
rect 44186 1696 44206 1702
rect 44064 1638 44206 1696
rect 44270 1638 44276 1702
rect 44064 1632 44276 1638
rect 45696 1752 45908 1844
rect 45696 1702 45810 1752
rect 45696 1638 45702 1702
rect 45766 1696 45810 1702
rect 45866 1696 45908 1752
rect 47464 1752 47676 1844
rect 47464 1708 47490 1752
rect 45766 1638 45908 1696
rect 45696 1632 45908 1638
rect 47328 1702 47490 1708
rect 47328 1638 47334 1702
rect 47398 1696 47490 1702
rect 47546 1696 47676 1752
rect 47398 1638 47676 1696
rect 47328 1632 47676 1638
rect 49096 1752 49308 1844
rect 49096 1702 49170 1752
rect 49096 1638 49102 1702
rect 49166 1696 49170 1702
rect 49226 1696 49308 1752
rect 49166 1638 49308 1696
rect 49096 1632 49308 1638
rect 50728 1752 50940 1844
rect 50728 1702 50850 1752
rect 50728 1638 50734 1702
rect 50798 1696 50850 1702
rect 50906 1696 50940 1752
rect 50798 1638 50940 1696
rect 50728 1632 50940 1638
rect 52496 1752 52708 1844
rect 52496 1702 52530 1752
rect 52496 1638 52502 1702
rect 52586 1696 52708 1752
rect 52566 1638 52708 1696
rect 52496 1632 52708 1638
rect 54128 1752 54340 1844
rect 54128 1702 54210 1752
rect 54128 1638 54134 1702
rect 54198 1696 54210 1702
rect 54266 1696 54340 1752
rect 55760 1752 55972 1844
rect 55760 1708 55890 1752
rect 54198 1638 54340 1696
rect 54128 1632 54340 1638
rect 55488 1702 55890 1708
rect 55488 1638 55494 1702
rect 55558 1696 55890 1702
rect 55946 1696 55972 1752
rect 55558 1638 55972 1696
rect 55488 1632 55972 1638
rect 57528 1752 57740 1844
rect 57528 1702 57570 1752
rect 57528 1638 57534 1702
rect 57626 1696 57740 1752
rect 57598 1638 57740 1696
rect 57528 1632 57740 1638
rect 59160 1752 59372 1844
rect 59160 1696 59250 1752
rect 59306 1708 59372 1752
rect 60792 1752 61140 1844
rect 59306 1702 59508 1708
rect 59306 1696 59438 1702
rect 59160 1638 59438 1696
rect 59502 1638 59508 1702
rect 59160 1632 59508 1638
rect 60792 1702 60930 1752
rect 60792 1638 60798 1702
rect 60862 1696 60930 1702
rect 60986 1696 61140 1752
rect 60862 1638 61140 1696
rect 60792 1632 61140 1638
rect 62560 1752 62772 1844
rect 62560 1702 62610 1752
rect 62560 1638 62566 1702
rect 62666 1696 62772 1752
rect 62630 1638 62772 1696
rect 62560 1632 62772 1638
rect 64192 1752 64404 1844
rect 64192 1696 64290 1752
rect 64346 1702 64404 1752
rect 64192 1638 64334 1696
rect 64398 1638 64404 1702
rect 64192 1632 64404 1638
rect 65824 1752 66172 1844
rect 65824 1702 65970 1752
rect 65824 1638 65830 1702
rect 65894 1696 65970 1702
rect 66026 1696 66172 1752
rect 65894 1638 66172 1696
rect 65824 1632 66172 1638
rect 67592 1752 67804 1844
rect 67592 1702 67650 1752
rect 67592 1638 67598 1702
rect 67706 1696 67804 1752
rect 67662 1638 67804 1696
rect 67592 1632 67804 1638
rect 69224 1752 69436 1844
rect 69224 1702 69330 1752
rect 69224 1638 69230 1702
rect 69294 1696 69330 1702
rect 69386 1696 69436 1752
rect 69294 1638 69436 1696
rect 69224 1632 69436 1638
rect 70856 1752 71204 1844
rect 70856 1702 71010 1752
rect 70856 1638 70862 1702
rect 70926 1696 71010 1702
rect 71066 1696 71204 1752
rect 70926 1638 71204 1696
rect 70856 1632 71204 1638
rect 72624 1752 72836 1844
rect 72624 1696 72690 1752
rect 72746 1702 72836 1752
rect 72746 1696 72766 1702
rect 72624 1638 72766 1696
rect 72830 1638 72836 1702
rect 72624 1632 72836 1638
rect 74256 1752 74468 1844
rect 74256 1702 74370 1752
rect 74256 1638 74262 1702
rect 74326 1696 74370 1702
rect 74426 1696 74468 1752
rect 74326 1638 74468 1696
rect 74256 1632 74468 1638
rect 76024 1752 76236 1844
rect 76024 1696 76050 1752
rect 76106 1702 76236 1752
rect 76106 1696 76166 1702
rect 76024 1638 76166 1696
rect 76230 1638 76236 1702
rect 76024 1632 76236 1638
rect 77656 1752 77868 1844
rect 77656 1702 77730 1752
rect 77656 1638 77662 1702
rect 77726 1696 77730 1702
rect 77786 1696 77868 1752
rect 77726 1638 77868 1696
rect 77656 1632 77868 1638
rect 79288 1752 79500 1844
rect 79288 1702 79410 1752
rect 79288 1638 79294 1702
rect 79358 1696 79410 1702
rect 79466 1696 79500 1752
rect 79358 1638 79500 1696
rect 79288 1632 79500 1638
rect 81056 1752 81268 1844
rect 81056 1702 81090 1752
rect 81056 1638 81062 1702
rect 81146 1696 81268 1752
rect 81126 1638 81268 1696
rect 81056 1632 81268 1638
rect 82688 1752 82900 1844
rect 82688 1696 82770 1752
rect 82826 1702 82900 1752
rect 82826 1696 82830 1702
rect 82688 1638 82830 1696
rect 82894 1638 82900 1702
rect 82688 1632 82900 1638
rect 84320 1752 84532 1844
rect 84320 1702 84450 1752
rect 84320 1638 84326 1702
rect 84390 1696 84450 1702
rect 84506 1696 84532 1752
rect 84390 1638 84532 1696
rect 84320 1632 84532 1638
rect 86088 1752 86300 1844
rect 86088 1696 86130 1752
rect 86186 1702 86300 1752
rect 86186 1696 86230 1702
rect 86088 1638 86230 1696
rect 86294 1638 86300 1702
rect 86088 1632 86300 1638
rect 87720 1752 87932 1844
rect 87720 1702 87810 1752
rect 87720 1638 87726 1702
rect 87790 1696 87810 1702
rect 87866 1696 87932 1752
rect 87790 1638 87932 1696
rect 87720 1632 87932 1638
rect 89352 1752 89700 1844
rect 89352 1702 89490 1752
rect 89352 1638 89358 1702
rect 89422 1696 89490 1702
rect 89546 1696 89700 1752
rect 89422 1638 89700 1696
rect 89352 1632 89700 1638
rect 91120 1752 91332 1844
rect 91120 1696 91170 1752
rect 91226 1702 91332 1752
rect 91226 1696 91262 1702
rect 91120 1638 91262 1696
rect 91326 1638 91332 1702
rect 91120 1632 91332 1638
rect 92752 1752 92964 1844
rect 92752 1702 92850 1752
rect 92752 1638 92758 1702
rect 92822 1696 92850 1702
rect 92906 1696 92964 1752
rect 92822 1638 92964 1696
rect 92752 1632 92964 1638
rect 94384 1752 94732 1844
rect 94384 1702 94530 1752
rect 94384 1638 94390 1702
rect 94454 1696 94530 1702
rect 94586 1696 94732 1752
rect 94454 1638 94732 1696
rect 94384 1632 94732 1638
rect 96152 1752 96364 1844
rect 96152 1702 96210 1752
rect 96152 1638 96158 1702
rect 96266 1696 96364 1752
rect 96222 1638 96364 1696
rect 96152 1632 96364 1638
rect 97784 1752 97996 1844
rect 97784 1702 97890 1752
rect 97784 1638 97790 1702
rect 97854 1696 97890 1702
rect 97946 1696 97996 1752
rect 97854 1638 97996 1696
rect 97784 1632 97996 1638
rect 99416 1752 99764 1844
rect 99416 1702 99570 1752
rect 99416 1638 99558 1702
rect 99626 1696 99764 1752
rect 99622 1638 99764 1696
rect 99416 1632 99764 1638
rect 101184 1752 101396 1844
rect 101184 1696 101250 1752
rect 101306 1702 101396 1752
rect 101306 1696 101326 1702
rect 101184 1638 101326 1696
rect 101390 1638 101396 1702
rect 101184 1632 101396 1638
rect 102816 1752 103028 1844
rect 102816 1702 102930 1752
rect 102816 1638 102822 1702
rect 102886 1696 102930 1702
rect 102986 1696 103028 1752
rect 102886 1638 103028 1696
rect 102816 1632 103028 1638
rect 104584 1752 104796 1844
rect 104584 1702 104610 1752
rect 104584 1638 104590 1702
rect 104666 1696 104796 1752
rect 104654 1638 104796 1696
rect 104584 1632 104796 1638
rect 106216 1752 106428 1844
rect 106216 1702 106290 1752
rect 106216 1638 106222 1702
rect 106286 1696 106290 1702
rect 106346 1696 106428 1752
rect 106286 1638 106428 1696
rect 106216 1632 106428 1638
rect 107848 1752 108060 1844
rect 107848 1702 107970 1752
rect 107848 1638 107854 1702
rect 107918 1696 107970 1702
rect 108026 1696 108060 1752
rect 107918 1638 108060 1696
rect 107848 1632 108060 1638
rect 109616 1752 109828 1844
rect 109616 1696 109650 1752
rect 109706 1702 109828 1752
rect 109706 1696 109758 1702
rect 109616 1638 109758 1696
rect 109822 1638 109828 1702
rect 109616 1632 109828 1638
rect 111248 1752 111460 1844
rect 111248 1702 111330 1752
rect 111248 1638 111254 1702
rect 111318 1696 111330 1702
rect 111386 1696 111460 1752
rect 111318 1638 111460 1696
rect 111248 1632 111460 1638
rect 112880 1752 113092 1844
rect 112880 1696 113010 1752
rect 113066 1702 113092 1752
rect 112880 1638 113022 1696
rect 113086 1638 113092 1702
rect 112880 1632 113092 1638
rect 114648 1752 114860 1844
rect 114648 1696 114690 1752
rect 114746 1702 114860 1752
rect 114746 1696 114790 1702
rect 114648 1638 114790 1696
rect 114854 1638 114860 1702
rect 114648 1632 114860 1638
rect 116280 1752 116492 1844
rect 116280 1702 116370 1752
rect 116280 1638 116286 1702
rect 116350 1696 116370 1702
rect 116426 1696 116492 1752
rect 116350 1638 116492 1696
rect 116280 1632 116492 1638
rect 117912 1752 118260 1844
rect 117912 1696 118050 1752
rect 118106 1702 118260 1752
rect 117912 1638 118054 1696
rect 118118 1638 118260 1702
rect 117912 1632 118260 1638
rect 119680 1752 119892 1844
rect 119680 1696 119730 1752
rect 119786 1702 119892 1752
rect 119786 1696 119822 1702
rect 119680 1638 119822 1696
rect 119886 1638 119892 1702
rect 119680 1632 119892 1638
rect 121312 1752 121524 1844
rect 121312 1702 121410 1752
rect 121312 1638 121318 1702
rect 121382 1696 121410 1702
rect 121466 1696 121524 1752
rect 121382 1638 121524 1696
rect 121312 1632 121524 1638
rect 122944 1752 123292 1844
rect 122944 1702 123090 1752
rect 123146 1702 123292 1752
rect 122944 1638 123086 1702
rect 123150 1638 123292 1702
rect 122944 1632 123292 1638
rect 124712 1752 124924 1844
rect 124712 1702 124770 1752
rect 124712 1638 124718 1702
rect 124826 1696 124924 1752
rect 124782 1638 124924 1696
rect 124712 1632 124924 1638
rect 126344 1752 126556 1844
rect 126344 1702 126450 1752
rect 126344 1638 126350 1702
rect 126414 1696 126450 1702
rect 126506 1696 126556 1752
rect 126414 1638 126556 1696
rect 126344 1632 126556 1638
rect 127976 1752 128324 1844
rect 127976 1702 128130 1752
rect 127976 1638 127982 1702
rect 128046 1696 128130 1702
rect 128186 1696 128324 1752
rect 128046 1638 128324 1696
rect 127976 1632 128324 1638
rect 129744 1752 129956 1844
rect 129744 1702 129810 1752
rect 129744 1638 129750 1702
rect 129866 1696 129956 1752
rect 129814 1638 129956 1696
rect 129744 1632 129956 1638
rect 131376 1752 131588 1844
rect 131376 1696 131490 1752
rect 131546 1702 131588 1752
rect 131376 1638 131518 1696
rect 131582 1638 131588 1702
rect 131376 1632 131588 1638
rect 133144 1752 133356 1844
rect 133144 1702 133170 1752
rect 133144 1638 133150 1702
rect 133226 1696 133356 1752
rect 133214 1638 133356 1696
rect 133144 1632 133356 1638
rect 952 1294 135668 1300
rect 952 1230 958 1294
rect 1022 1230 1094 1294
rect 1158 1230 1230 1294
rect 1294 1230 2046 1294
rect 2110 1230 3814 1294
rect 3878 1230 5582 1294
rect 5646 1230 7078 1294
rect 7142 1230 8710 1294
rect 8774 1230 10478 1294
rect 10542 1230 12110 1294
rect 12174 1230 14014 1294
rect 14078 1230 15510 1294
rect 15574 1230 17414 1294
rect 17478 1230 19046 1294
rect 19110 1230 20814 1294
rect 20878 1230 22174 1294
rect 22238 1230 23942 1294
rect 24006 1230 25710 1294
rect 25774 1230 27342 1294
rect 27406 1230 28974 1294
rect 29038 1230 30470 1294
rect 30534 1230 32102 1294
rect 32166 1230 34006 1294
rect 34070 1230 35774 1294
rect 35838 1230 37406 1294
rect 37470 1230 39174 1294
rect 39238 1230 40806 1294
rect 40870 1230 42438 1294
rect 42502 1230 44206 1294
rect 44270 1230 45702 1294
rect 45766 1230 47334 1294
rect 47398 1230 49102 1294
rect 49166 1230 50734 1294
rect 50798 1230 52502 1294
rect 52566 1230 54134 1294
rect 54198 1230 55494 1294
rect 55558 1230 57534 1294
rect 57598 1230 59438 1294
rect 59502 1230 60798 1294
rect 60862 1230 62566 1294
rect 62630 1230 64334 1294
rect 64398 1230 65830 1294
rect 65894 1230 67598 1294
rect 67662 1230 69230 1294
rect 69294 1230 70862 1294
rect 70926 1230 72766 1294
rect 72830 1230 74262 1294
rect 74326 1230 76166 1294
rect 76230 1230 77662 1294
rect 77726 1230 79294 1294
rect 79358 1230 81062 1294
rect 81126 1230 82830 1294
rect 82894 1230 84326 1294
rect 84390 1230 86230 1294
rect 86294 1230 87726 1294
rect 87790 1230 89358 1294
rect 89422 1230 91262 1294
rect 91326 1230 92758 1294
rect 92822 1230 94390 1294
rect 94454 1230 96158 1294
rect 96222 1230 97790 1294
rect 97854 1230 99558 1294
rect 99622 1230 101326 1294
rect 101390 1230 102822 1294
rect 102886 1230 104590 1294
rect 104654 1230 106222 1294
rect 106286 1230 107854 1294
rect 107918 1230 109758 1294
rect 109822 1230 111254 1294
rect 111318 1230 113022 1294
rect 113086 1230 114790 1294
rect 114854 1230 116286 1294
rect 116350 1230 118054 1294
rect 118118 1230 119822 1294
rect 119886 1230 121318 1294
rect 121382 1230 123086 1294
rect 123150 1230 124718 1294
rect 124782 1230 126350 1294
rect 126414 1230 127982 1294
rect 128046 1230 129750 1294
rect 129814 1230 131518 1294
rect 131582 1230 133150 1294
rect 133214 1230 135326 1294
rect 135390 1230 135462 1294
rect 135526 1230 135598 1294
rect 135662 1230 135668 1294
rect 952 1158 135668 1230
rect 952 1094 958 1158
rect 1022 1094 1094 1158
rect 1158 1094 1230 1158
rect 1294 1094 135326 1158
rect 135390 1094 135462 1158
rect 135526 1094 135598 1158
rect 135662 1094 135668 1158
rect 952 1022 135668 1094
rect 952 958 958 1022
rect 1022 958 1094 1022
rect 1158 958 1230 1022
rect 1294 958 135326 1022
rect 135390 958 135462 1022
rect 135526 958 135598 1022
rect 135662 958 135668 1022
rect 952 952 135668 958
rect 272 614 136348 620
rect 272 550 278 614
rect 342 550 414 614
rect 478 550 550 614
rect 614 550 39718 614
rect 39782 550 136006 614
rect 136070 550 136142 614
rect 136206 550 136278 614
rect 136342 550 136348 614
rect 272 478 136348 550
rect 272 414 278 478
rect 342 414 414 478
rect 478 414 550 478
rect 614 414 136006 478
rect 136070 414 136142 478
rect 136206 414 136278 478
rect 136342 414 136348 478
rect 272 342 136348 414
rect 272 278 278 342
rect 342 278 414 342
rect 478 278 550 342
rect 614 278 136006 342
rect 136070 278 136142 342
rect 136206 278 136278 342
rect 136342 278 136348 342
rect 272 272 136348 278
<< via3 >>
rect 278 82966 342 83030
rect 414 82966 478 83030
rect 550 82966 614 83030
rect 136006 82966 136070 83030
rect 136142 82966 136206 83030
rect 136278 82966 136342 83030
rect 278 82830 342 82894
rect 414 82830 478 82894
rect 550 82830 614 82894
rect 136006 82830 136070 82894
rect 136142 82830 136206 82894
rect 136278 82830 136342 82894
rect 278 82694 342 82758
rect 414 82694 478 82758
rect 550 82694 614 82758
rect 118054 82694 118118 82758
rect 136006 82694 136070 82758
rect 136142 82694 136206 82758
rect 136278 82694 136342 82758
rect 958 82286 1022 82350
rect 1094 82286 1158 82350
rect 1230 82286 1294 82350
rect 135326 82286 135390 82350
rect 135462 82286 135526 82350
rect 135598 82286 135662 82350
rect 958 82150 1022 82214
rect 1094 82150 1158 82214
rect 1230 82150 1294 82214
rect 135326 82150 135390 82214
rect 135462 82150 135526 82214
rect 135598 82150 135662 82214
rect 958 82014 1022 82078
rect 1094 82014 1158 82078
rect 1230 82014 1294 82078
rect 2182 82014 2246 82078
rect 3950 82014 4014 82078
rect 5446 82014 5510 82078
rect 7214 82014 7278 82078
rect 8710 82014 8774 82078
rect 10478 82014 10542 82078
rect 12110 82014 12174 82078
rect 14014 82014 14078 82078
rect 15646 82014 15710 82078
rect 17142 82014 17206 82078
rect 18910 82014 18974 82078
rect 20678 82014 20742 82078
rect 22174 82014 22238 82078
rect 23942 82014 24006 82078
rect 25710 82014 25774 82078
rect 27206 82014 27270 82078
rect 28974 82014 29038 82078
rect 30606 82014 30670 82078
rect 32374 82014 32438 82078
rect 34142 82014 34206 82078
rect 35638 82014 35702 82078
rect 37542 82014 37606 82078
rect 39174 82014 39238 82078
rect 40670 82014 40734 82078
rect 42438 82014 42502 82078
rect 44206 82014 44270 82078
rect 45702 82014 45766 82078
rect 47470 82014 47534 82078
rect 49238 82014 49302 82078
rect 50734 82014 50798 82078
rect 52638 82014 52702 82078
rect 54134 82014 54198 82078
rect 55902 82014 55966 82078
rect 57670 82014 57734 82078
rect 59166 82014 59230 82078
rect 60798 82014 60862 82078
rect 62702 82014 62766 82078
rect 64198 82014 64262 82078
rect 65830 82014 65894 82078
rect 67598 82014 67662 82078
rect 69230 82014 69294 82078
rect 70862 82014 70926 82078
rect 72630 82014 72694 82078
rect 74398 82014 74462 82078
rect 76166 82014 76230 82078
rect 77662 82014 77726 82078
rect 79430 82014 79494 82078
rect 81334 82014 81398 82078
rect 82694 82014 82758 82078
rect 84462 82014 84526 82078
rect 86230 82014 86294 82078
rect 87726 82014 87790 82078
rect 89358 82014 89422 82078
rect 91126 82014 91190 82078
rect 92894 82014 92958 82078
rect 94390 82014 94454 82078
rect 96294 82014 96358 82078
rect 97926 82014 97990 82078
rect 99694 82014 99758 82078
rect 101326 82014 101390 82078
rect 102958 82014 103022 82078
rect 104590 82014 104654 82078
rect 106358 82014 106422 82078
rect 107854 82014 107918 82078
rect 109622 82014 109686 82078
rect 111390 82014 111454 82078
rect 112886 82014 112950 82078
rect 114654 82014 114718 82078
rect 116422 82014 116486 82078
rect 117918 82014 117982 82078
rect 119550 82014 119614 82078
rect 121454 82014 121518 82078
rect 123222 82014 123286 82078
rect 124718 82014 124782 82078
rect 126350 82014 126414 82078
rect 128118 82014 128182 82078
rect 129886 82014 129950 82078
rect 131382 82014 131446 82078
rect 133150 82014 133214 82078
rect 135326 82014 135390 82078
rect 135462 82014 135526 82078
rect 135598 82014 135662 82078
rect 2182 81501 2246 81534
rect 2182 81470 2186 81501
rect 2186 81470 2246 81501
rect 2046 81334 2110 81398
rect 3950 81470 4014 81534
rect 5446 81501 5510 81534
rect 5446 81470 5490 81501
rect 5490 81470 5510 81501
rect 7214 81501 7278 81534
rect 7214 81470 7226 81501
rect 7226 81470 7278 81501
rect 8710 81470 8774 81534
rect 10478 81501 10542 81534
rect 10478 81470 10530 81501
rect 10530 81470 10542 81501
rect 12110 81470 12174 81534
rect 14014 81470 14078 81534
rect 15646 81470 15710 81534
rect 17142 81470 17206 81534
rect 18910 81501 18974 81534
rect 18910 81470 18930 81501
rect 18930 81470 18974 81501
rect 20678 81470 20742 81534
rect 22174 81470 22238 81534
rect 23942 81501 24006 81534
rect 23942 81470 23970 81501
rect 23970 81470 24006 81501
rect 25710 81470 25774 81534
rect 27206 81470 27270 81534
rect 28974 81501 29038 81534
rect 28974 81470 29010 81501
rect 29010 81470 29038 81501
rect 30606 81470 30670 81534
rect 32374 81501 32438 81534
rect 32374 81470 32426 81501
rect 32426 81470 32438 81501
rect 34142 81470 34206 81534
rect 35638 81470 35702 81534
rect 37542 81470 37606 81534
rect 39174 81470 39238 81534
rect 40670 81470 40734 81534
rect 42438 81501 42502 81534
rect 42438 81470 42450 81501
rect 42450 81470 42502 81501
rect 44206 81470 44270 81534
rect 45702 81470 45766 81534
rect 47470 81501 47534 81534
rect 47470 81470 47490 81501
rect 47490 81470 47534 81501
rect 49238 81470 49302 81534
rect 50734 81470 50798 81534
rect 52638 81470 52702 81534
rect 54134 81470 54198 81534
rect 55902 81501 55966 81534
rect 55902 81470 55946 81501
rect 55946 81470 55966 81501
rect 57670 81470 57734 81534
rect 59166 81470 59230 81534
rect 60798 81470 60862 81534
rect 62702 81470 62766 81534
rect 64198 81470 64262 81534
rect 65830 81470 65894 81534
rect 67598 81501 67662 81534
rect 67598 81470 67650 81501
rect 67650 81470 67662 81501
rect 69230 81470 69294 81534
rect 70862 81470 70926 81534
rect 72630 81501 72694 81534
rect 72630 81470 72690 81501
rect 72690 81470 72694 81501
rect 74398 81501 74462 81534
rect 74398 81470 74426 81501
rect 74426 81470 74462 81501
rect 76166 81470 76230 81534
rect 77662 81470 77726 81534
rect 79430 81501 79494 81534
rect 79430 81470 79466 81501
rect 79466 81470 79494 81501
rect 81334 81470 81398 81534
rect 82694 81470 82758 81534
rect 84462 81501 84526 81534
rect 84462 81470 84506 81501
rect 84506 81470 84526 81501
rect 86230 81470 86294 81534
rect 87726 81470 87790 81534
rect 89358 81470 89422 81534
rect 91126 81501 91190 81534
rect 91126 81470 91170 81501
rect 91170 81470 91190 81501
rect 92894 81501 92958 81534
rect 92894 81470 92906 81501
rect 92906 81470 92958 81501
rect 94390 81470 94454 81534
rect 96294 81470 96358 81534
rect 97926 81501 97990 81534
rect 97926 81470 97946 81501
rect 97946 81470 97990 81501
rect 99694 81470 99758 81534
rect 101326 81470 101390 81534
rect 102958 81501 103022 81534
rect 102958 81470 102986 81501
rect 102986 81470 103022 81501
rect 104590 81501 104654 81534
rect 104590 81470 104610 81501
rect 104610 81470 104654 81501
rect 106358 81470 106422 81534
rect 107854 81470 107918 81534
rect 109622 81501 109686 81534
rect 109622 81470 109650 81501
rect 109650 81470 109686 81501
rect 111390 81470 111454 81534
rect 112886 81470 112950 81534
rect 114654 81501 114718 81534
rect 114654 81470 114690 81501
rect 114690 81470 114718 81501
rect 116422 81501 116486 81534
rect 116422 81470 116426 81501
rect 116426 81470 116486 81501
rect 117918 81470 117982 81534
rect 119550 81470 119614 81534
rect 118190 81334 118254 81398
rect 121454 81501 121518 81534
rect 121454 81470 121466 81501
rect 121466 81470 121518 81501
rect 123222 81470 123286 81534
rect 122950 81334 123014 81398
rect 124718 81501 124782 81534
rect 124718 81470 124770 81501
rect 124770 81470 124782 81501
rect 126350 81470 126414 81534
rect 128118 81501 128182 81534
rect 128118 81470 128130 81501
rect 128130 81470 128182 81501
rect 129886 81470 129950 81534
rect 131382 81470 131446 81534
rect 133150 81501 133214 81534
rect 133150 81470 133170 81501
rect 133170 81470 133214 81501
rect 2046 81062 2110 81126
rect 135326 80926 135390 80990
rect 118054 80790 118118 80854
rect 117918 80654 117982 80718
rect 122270 80654 122334 80718
rect 118462 80246 118526 80310
rect 119686 80246 119750 80310
rect 122270 79838 122334 79902
rect 122406 79702 122470 79766
rect 136006 79838 136070 79902
rect 1230 79430 1294 79494
rect 118190 79430 118254 79494
rect 135326 79430 135390 79494
rect 118054 79294 118118 79358
rect 130838 79158 130902 79222
rect 117918 78614 117982 78678
rect 116558 78478 116622 78542
rect 122950 78478 123014 78542
rect 122270 78342 122334 78406
rect 134782 78342 134846 78406
rect 1230 77526 1294 77590
rect 134782 77688 134846 77726
rect 134782 77662 134844 77688
rect 134844 77662 134846 77688
rect 135326 77662 135390 77726
rect 118054 77254 118118 77318
rect 28702 77118 28766 77182
rect 28974 76982 29038 77046
rect 31014 77118 31078 77182
rect 31422 76982 31486 77046
rect 33462 77118 33526 77182
rect 34006 76982 34070 77046
rect 36182 77118 36246 77182
rect 36454 76982 36518 77046
rect 38494 77118 38558 77182
rect 41078 77118 41142 77182
rect 39038 76982 39102 77046
rect 41486 76982 41550 77046
rect 43526 77118 43590 77182
rect 43934 76982 43998 77046
rect 46110 77118 46174 77182
rect 48558 77118 48622 77182
rect 46518 76982 46582 77046
rect 48966 76982 49030 77046
rect 51142 77118 51206 77182
rect 51414 76982 51478 77046
rect 53590 77118 53654 77182
rect 53862 76982 53926 77046
rect 56174 77118 56238 77182
rect 56446 76982 56510 77046
rect 58486 77118 58550 77182
rect 58894 76982 58958 77046
rect 60934 77118 60998 77182
rect 61478 77118 61542 77182
rect 63654 77118 63718 77182
rect 63926 76982 63990 77046
rect 66102 77118 66166 77182
rect 68550 77118 68614 77182
rect 68958 77118 69022 77182
rect 70998 77118 71062 77182
rect 66510 76982 66574 77046
rect 71406 76982 71470 77046
rect 73582 77118 73646 77182
rect 73854 76982 73918 77046
rect 75894 77118 75958 77182
rect 76438 76982 76502 77046
rect 78614 77118 78678 77182
rect 78886 76982 78950 77046
rect 81062 77118 81126 77182
rect 83510 77118 83574 77182
rect 81470 76982 81534 77046
rect 83918 76982 83982 77046
rect 85958 77118 86022 77182
rect 86366 76982 86430 77046
rect 88406 77118 88470 77182
rect 90990 77118 91054 77182
rect 91262 77118 91326 77182
rect 88950 76982 89014 77046
rect 93574 77118 93638 77182
rect 93846 76982 93910 77046
rect 96022 77118 96086 77182
rect 96294 76982 96358 77046
rect 98470 77118 98534 77182
rect 98878 76982 98942 77046
rect 101054 77118 101118 77182
rect 101326 76982 101390 77046
rect 103366 77118 103430 77182
rect 103910 77118 103974 77182
rect 106086 77118 106150 77182
rect 115334 77118 115398 77182
rect 106358 76982 106422 77046
rect 122406 76982 122470 77046
rect 122406 76846 122470 76910
rect 28974 76574 29038 76638
rect 31286 76574 31350 76638
rect 33734 76574 33798 76638
rect 36318 76574 36382 76638
rect 38630 76574 38694 76638
rect 38902 76574 38966 76638
rect 41350 76574 41414 76638
rect 43662 76574 43726 76638
rect 43934 76574 43998 76638
rect 46382 76574 46446 76638
rect 48694 76574 48758 76638
rect 51414 76574 51478 76638
rect 53726 76574 53790 76638
rect 56174 76574 56238 76638
rect 56310 76574 56374 76638
rect 58758 76574 58822 76638
rect 61342 76574 61406 76638
rect 63790 76574 63854 76638
rect 66374 76574 66438 76638
rect 68822 76574 68886 76638
rect 71134 76574 71198 76638
rect 71406 76574 71470 76638
rect 73718 76574 73782 76638
rect 76166 76574 76230 76638
rect 78614 76574 78678 76638
rect 78750 76574 78814 76638
rect 81334 76574 81398 76638
rect 83782 76574 83846 76638
rect 86366 76574 86430 76638
rect 88542 76574 88606 76638
rect 88814 76574 88878 76638
rect 91398 76574 91462 76638
rect 93574 76574 93638 76638
rect 93846 76574 93910 76638
rect 96158 76574 96222 76638
rect 98606 76574 98670 76638
rect 98742 76574 98806 76638
rect 101190 76574 101254 76638
rect 103774 76574 103838 76638
rect 106222 76574 106286 76638
rect 1230 76030 1294 76094
rect 135326 76030 135390 76094
rect 28974 75894 29038 75958
rect 31286 75894 31350 75958
rect 33734 75894 33798 75958
rect 36318 75894 36382 75958
rect 38630 75894 38694 75958
rect 38902 75894 38966 75958
rect 41350 75894 41414 75958
rect 43662 75894 43726 75958
rect 43934 75894 43998 75958
rect 46382 75894 46446 75958
rect 48694 75894 48758 75958
rect 51414 75894 51478 75958
rect 53726 75894 53790 75958
rect 56174 75894 56238 75958
rect 56310 75894 56374 75958
rect 58758 75894 58822 75958
rect 61342 75894 61406 75958
rect 63790 75894 63854 75958
rect 66374 75894 66438 75958
rect 59438 75758 59502 75822
rect 68822 75894 68886 75958
rect 71134 75894 71198 75958
rect 71406 75894 71470 75958
rect 73718 75894 73782 75958
rect 76166 75894 76230 75958
rect 78614 75894 78678 75958
rect 78750 75894 78814 75958
rect 81334 75894 81398 75958
rect 83782 75894 83846 75958
rect 86366 75894 86430 75958
rect 88542 75894 88606 75958
rect 88814 75894 88878 75958
rect 91398 75894 91462 75958
rect 93574 75894 93638 75958
rect 93846 75894 93910 75958
rect 96158 75894 96222 75958
rect 98606 75894 98670 75958
rect 98742 75894 98806 75958
rect 101190 75894 101254 75958
rect 103774 75894 103838 75958
rect 106222 75894 106286 75958
rect 116558 75894 116622 75958
rect 115470 75622 115534 75686
rect 122270 75622 122334 75686
rect 122270 75486 122334 75550
rect 28838 75214 28902 75278
rect 28974 75078 29038 75142
rect 31422 75214 31486 75278
rect 31558 75078 31622 75142
rect 34006 75214 34070 75278
rect 34006 75078 34070 75142
rect 36454 75214 36518 75278
rect 36454 75078 36518 75142
rect 39038 75214 39102 75278
rect 39038 75078 39102 75142
rect 41486 75214 41550 75278
rect 41486 75078 41550 75142
rect 43798 75214 43862 75278
rect 46518 75214 46582 75278
rect 44070 75078 44134 75142
rect 46518 75078 46582 75142
rect 48966 75214 49030 75278
rect 48966 75078 49030 75142
rect 51278 75214 51342 75278
rect 53862 75214 53926 75278
rect 51550 75078 51614 75142
rect 53998 75078 54062 75142
rect 56446 75214 56510 75278
rect 56310 75078 56374 75142
rect 58894 75214 58958 75278
rect 59030 75078 59094 75142
rect 61478 75214 61542 75278
rect 61478 75078 61542 75142
rect 63926 75214 63990 75278
rect 63926 75078 63990 75142
rect 66510 75214 66574 75278
rect 66510 75078 66574 75142
rect 68958 75214 69022 75278
rect 68958 75078 69022 75142
rect 71270 75214 71334 75278
rect 71406 75078 71470 75142
rect 73854 75214 73918 75278
rect 73990 75078 74054 75142
rect 76438 75214 76502 75278
rect 76438 75078 76502 75142
rect 78886 75214 78950 75278
rect 78886 75078 78950 75142
rect 81470 75214 81534 75278
rect 81470 75078 81534 75142
rect 83918 75214 83982 75278
rect 83918 75078 83982 75142
rect 86230 75214 86294 75278
rect 88950 75214 89014 75278
rect 86502 75078 86566 75142
rect 88950 75078 89014 75142
rect 91262 75214 91326 75278
rect 91398 75078 91462 75142
rect 93710 75214 93774 75278
rect 93710 75078 93774 75142
rect 96294 75214 96358 75278
rect 96430 75078 96494 75142
rect 98878 75214 98942 75278
rect 98878 75078 98942 75142
rect 101326 75214 101390 75278
rect 101462 75078 101526 75142
rect 103910 75214 103974 75278
rect 103910 75078 103974 75142
rect 106358 75214 106422 75278
rect 106358 75078 106422 75142
rect 115334 74398 115398 74462
rect 115334 74262 115398 74326
rect 122406 74262 122470 74326
rect 1230 74126 1294 74190
rect 122406 73990 122470 74054
rect 135326 74126 135390 74190
rect 28974 73174 29038 73238
rect 31558 73174 31622 73238
rect 28974 73038 29038 73102
rect 34006 73174 34070 73238
rect 36454 73174 36518 73238
rect 39038 73174 39102 73238
rect 41486 73174 41550 73238
rect 44070 73174 44134 73238
rect 46518 73174 46582 73238
rect 48966 73174 49030 73238
rect 51550 73174 51614 73238
rect 53998 73174 54062 73238
rect 56310 73174 56374 73238
rect 59030 73174 59094 73238
rect 61478 73174 61542 73238
rect 63926 73174 63990 73238
rect 66510 73174 66574 73238
rect 68958 73174 69022 73238
rect 71406 73174 71470 73238
rect 73990 73174 74054 73238
rect 76438 73174 76502 73238
rect 78886 73174 78950 73238
rect 81470 73174 81534 73238
rect 83918 73174 83982 73238
rect 86502 73174 86566 73238
rect 88950 73174 89014 73238
rect 91398 73174 91462 73238
rect 93710 73174 93774 73238
rect 96430 73174 96494 73238
rect 98878 73174 98942 73238
rect 101462 73174 101526 73238
rect 103910 73174 103974 73238
rect 106358 73174 106422 73238
rect 109622 73038 109686 73102
rect 115470 73038 115534 73102
rect 115878 72902 115942 72966
rect 122270 72766 122334 72830
rect 1230 72630 1294 72694
rect 136006 72766 136070 72830
rect 135326 72494 135390 72558
rect 134093 72294 134157 72358
rect 28566 71406 28630 71470
rect 28702 71406 28766 71470
rect 29790 71406 29854 71470
rect 31286 71406 31350 71470
rect 31966 71406 32030 71470
rect 32510 71406 32574 71470
rect 33734 71406 33798 71470
rect 34414 71406 34478 71470
rect 34958 71406 35022 71470
rect 35774 71406 35838 71470
rect 36182 71406 36246 71470
rect 36998 71406 37062 71470
rect 37542 71406 37606 71470
rect 38222 71406 38286 71470
rect 39990 71406 40054 71470
rect 40670 71406 40734 71470
rect 41214 71406 41278 71470
rect 41894 71406 41958 71470
rect 42438 71406 42502 71470
rect 43254 71406 43318 71470
rect 44614 71406 44678 71470
rect 45702 71406 45766 71470
rect 46246 71406 46310 71470
rect 46926 71406 46990 71470
rect 48694 71406 48758 71470
rect 49918 71406 49982 71470
rect 50734 71406 50798 71470
rect 51278 71406 51342 71470
rect 52502 71406 52566 71470
rect 53182 71406 53246 71470
rect 53318 71406 53382 71470
rect 54406 71406 54470 71470
rect 54950 71406 55014 71470
rect 56038 71406 56102 71470
rect 57398 71406 57462 71470
rect 58622 71406 58686 71470
rect 59438 71542 59502 71606
rect 59438 71406 59502 71470
rect 59982 71406 60046 71470
rect 61206 71406 61270 71470
rect 61886 71406 61950 71470
rect 62430 71406 62494 71470
rect 63110 71406 63174 71470
rect 63654 71406 63718 71470
rect 65014 71406 65078 71470
rect 66102 71406 66166 71470
rect 66918 71406 66982 71470
rect 67462 71406 67526 71470
rect 68142 71406 68206 71470
rect 68686 71406 68750 71470
rect 69910 71406 69974 71470
rect 70590 71406 70654 71470
rect 72086 71406 72150 71470
rect 72222 71406 72286 71470
rect 73718 71406 73782 71470
rect 74398 71406 74462 71470
rect 74942 71406 75006 71470
rect 75622 71406 75686 71470
rect 76166 71406 76230 71470
rect 76846 71406 76910 71470
rect 77390 71406 77454 71470
rect 78206 71406 78270 71470
rect 78478 71406 78542 71470
rect 79430 71406 79494 71470
rect 79974 71406 80038 71470
rect 80654 71406 80718 71470
rect 81878 71406 81942 71470
rect 82422 71406 82486 71470
rect 83102 71406 83166 71470
rect 83646 71406 83710 71470
rect 84598 71406 84662 71470
rect 86094 71406 86158 71470
rect 86910 71406 86974 71470
rect 88134 71406 88198 71470
rect 88678 71406 88742 71470
rect 89358 71406 89422 71470
rect 89902 71406 89966 71470
rect 90718 71406 90782 71470
rect 91126 71406 91190 71470
rect 92350 71406 92414 71470
rect 93302 71406 93366 71470
rect 94934 71406 94998 71470
rect 95614 71406 95678 71470
rect 96838 71406 96902 71470
rect 97382 71406 97446 71470
rect 99830 71406 99894 71470
rect 100918 71406 100982 71470
rect 101870 71406 101934 71470
rect 102414 71406 102478 71470
rect 103094 71406 103158 71470
rect 103638 71406 103702 71470
rect 104318 71406 104382 71470
rect 104862 71406 104926 71470
rect 105542 71406 105606 71470
rect 106086 71406 106150 71470
rect 107310 71406 107374 71470
rect 108534 71406 108598 71470
rect 122406 71406 122470 71470
rect 98606 71270 98670 71334
rect 134782 71270 134846 71334
rect 1230 70998 1294 71062
rect 28566 70998 28630 71062
rect 28702 70998 28766 71062
rect 29790 70998 29854 71062
rect 31286 70998 31350 71062
rect 31966 70998 32030 71062
rect 32510 70998 32574 71062
rect 33734 70998 33798 71062
rect 34414 70998 34478 71062
rect 34958 70998 35022 71062
rect 35774 70998 35838 71062
rect 36182 70998 36246 71062
rect 36998 70998 37062 71062
rect 37542 70998 37606 71062
rect 38222 70998 38286 71062
rect 39990 70998 40054 71062
rect 40670 70998 40734 71062
rect 41214 70998 41278 71062
rect 41894 70998 41958 71062
rect 42438 70998 42502 71062
rect 43254 70998 43318 71062
rect 44614 70862 44678 70926
rect 45702 70998 45766 71062
rect 46246 70998 46310 71062
rect 46926 70998 46990 71062
rect 48694 70998 48758 71062
rect 49918 70998 49982 71062
rect 50734 70998 50798 71062
rect 51278 70998 51342 71062
rect 52502 70998 52566 71062
rect 53182 70998 53246 71062
rect 53318 70998 53382 71062
rect 54406 70998 54470 71062
rect 54950 70998 55014 71062
rect 56038 70998 56102 71062
rect 57398 70998 57462 71062
rect 58622 70998 58686 71062
rect 59438 70998 59502 71062
rect 59982 70998 60046 71062
rect 61206 70998 61270 71062
rect 61886 70998 61950 71062
rect 62430 70998 62494 71062
rect 63110 70998 63174 71062
rect 63654 70998 63718 71062
rect 65014 70998 65078 71062
rect 66102 70998 66166 71062
rect 66918 70998 66982 71062
rect 67462 70998 67526 71062
rect 68142 70998 68206 71062
rect 68686 70998 68750 71062
rect 69910 70998 69974 71062
rect 70590 70998 70654 71062
rect 72222 70998 72286 71062
rect 72086 70862 72150 70926
rect 73718 70998 73782 71062
rect 74398 70998 74462 71062
rect 74942 70998 75006 71062
rect 75622 70998 75686 71062
rect 76166 70998 76230 71062
rect 76846 70998 76910 71062
rect 77390 70998 77454 71062
rect 78206 70998 78270 71062
rect 78478 70998 78542 71062
rect 79430 70998 79494 71062
rect 79974 70998 80038 71062
rect 80654 70998 80718 71062
rect 81878 70998 81942 71062
rect 82422 70998 82486 71062
rect 83102 70998 83166 71062
rect 83646 70998 83710 71062
rect 84598 70998 84662 71062
rect 86094 70998 86158 71062
rect 86910 70998 86974 71062
rect 88134 70998 88198 71062
rect 88678 70998 88742 71062
rect 89358 70998 89422 71062
rect 89902 70998 89966 71062
rect 90718 70998 90782 71062
rect 91126 70998 91190 71062
rect 92350 70998 92414 71062
rect 93302 70862 93366 70926
rect 94934 70998 94998 71062
rect 95614 70998 95678 71062
rect 96838 70998 96902 71062
rect 97382 70998 97446 71062
rect 98606 70998 98670 71062
rect 99830 70998 99894 71062
rect 100918 70998 100982 71062
rect 101870 70998 101934 71062
rect 102414 70998 102478 71062
rect 103094 70998 103158 71062
rect 103638 70998 103702 71062
rect 104318 70998 104382 71062
rect 104862 70998 104926 71062
rect 105542 70998 105606 71062
rect 106086 70998 106150 71062
rect 107310 70998 107374 71062
rect 108534 70998 108598 71062
rect 110710 70998 110774 71062
rect 134782 70998 134846 71062
rect 109622 70862 109686 70926
rect 28974 70726 29038 70790
rect 135326 70862 135390 70926
rect 110710 70590 110774 70654
rect 115334 70590 115398 70654
rect 114246 70454 114310 70518
rect 22174 69910 22238 69974
rect 22446 69910 22510 69974
rect 114246 70046 114310 70110
rect 114382 69910 114446 69974
rect 114654 69910 114718 69974
rect 115334 69910 115398 69974
rect 115470 69910 115534 69974
rect 115878 70046 115942 70110
rect 20814 69502 20878 69566
rect 21358 69502 21422 69566
rect 21630 69502 21694 69566
rect 22174 69638 22238 69702
rect 22174 69502 22238 69566
rect 22446 69638 22510 69702
rect 22446 69502 22510 69566
rect 114382 69638 114446 69702
rect 114246 69502 114310 69566
rect 114654 69638 114718 69702
rect 114654 69502 114718 69566
rect 115334 69638 115398 69702
rect 115470 69638 115534 69702
rect 115062 69502 115126 69566
rect 115606 69502 115670 69566
rect 133150 69774 133214 69838
rect 116014 69502 116078 69566
rect 1230 69230 1294 69294
rect 20814 69230 20878 69294
rect 21358 69230 21422 69294
rect 21630 69230 21694 69294
rect 21766 69094 21830 69158
rect 22174 69230 22238 69294
rect 22038 69094 22102 69158
rect 22446 69230 22510 69294
rect 135326 69366 135390 69430
rect 22446 69094 22510 69158
rect 114246 69230 114310 69294
rect 114382 69094 114446 69158
rect 114654 69230 114718 69294
rect 114790 69094 114854 69158
rect 115062 69230 115126 69294
rect 115198 69094 115262 69158
rect 115606 69230 115670 69294
rect 116014 69230 116078 69294
rect 134782 69094 134846 69158
rect 20814 68822 20878 68886
rect 21766 68822 21830 68886
rect 22038 68822 22102 68886
rect 22038 68686 22102 68750
rect 22446 68822 22510 68886
rect 22446 68686 22510 68750
rect 20814 68550 20878 68614
rect 21902 68278 21966 68342
rect 22038 68414 22102 68478
rect 22446 68414 22510 68478
rect 114382 68822 114446 68886
rect 114790 68822 114854 68886
rect 114382 68686 114446 68750
rect 114654 68686 114718 68750
rect 115198 68822 115262 68886
rect 116014 68822 116078 68886
rect 20814 68006 20878 68070
rect 21902 68006 21966 68070
rect 20814 67734 20878 67798
rect 20814 67598 20878 67662
rect 21222 67598 21286 67662
rect 21630 67598 21694 67662
rect 27478 68142 27542 68206
rect 27342 67870 27406 67934
rect 27478 67870 27542 67934
rect 1230 67462 1294 67526
rect 20814 67326 20878 67390
rect 20814 67190 20878 67254
rect 21222 67326 21286 67390
rect 21630 67326 21694 67390
rect 21494 67190 21558 67254
rect 22038 67190 22102 67254
rect 109486 68142 109550 68206
rect 109486 67870 109550 67934
rect 114382 68414 114446 68478
rect 114654 68414 114718 68478
rect 115334 68278 115398 68342
rect 116014 68550 116078 68614
rect 134782 68550 134846 68614
rect 115334 68006 115398 68070
rect 115878 68006 115942 68070
rect 109350 67734 109414 67798
rect 27342 67598 27406 67662
rect 115606 67598 115670 67662
rect 115878 67734 115942 67798
rect 116014 67598 116078 67662
rect 135326 67598 135390 67662
rect 22446 67190 22510 67254
rect 109350 67326 109414 67390
rect 109486 67326 109550 67390
rect 114382 67190 114446 67254
rect 114654 67190 114718 67254
rect 20814 66918 20878 66982
rect 20814 66782 20878 66846
rect 21494 66918 21558 66982
rect 21630 66782 21694 66846
rect 22038 66918 22102 66982
rect 22038 66782 22102 66846
rect 22446 66918 22510 66982
rect 22446 66782 22510 66846
rect 109486 67054 109550 67118
rect 115606 67326 115670 67390
rect 116014 67326 116078 67390
rect 115878 67190 115942 67254
rect 133150 67054 133214 67118
rect 114382 66918 114446 66982
rect 114382 66782 114446 66846
rect 114654 66918 114718 66982
rect 114790 66782 114854 66846
rect 115606 66782 115670 66846
rect 115878 66918 115942 66982
rect 132606 66918 132670 66982
rect 115878 66782 115942 66846
rect 20814 66510 20878 66574
rect 20950 66374 21014 66438
rect 21630 66510 21694 66574
rect 21358 66374 21422 66438
rect 21494 66374 21558 66438
rect 22038 66510 22102 66574
rect 22174 66374 22238 66438
rect 22446 66510 22510 66574
rect 22582 66374 22646 66438
rect 114382 66510 114446 66574
rect 114246 66374 114310 66438
rect 114790 66510 114854 66574
rect 114654 66374 114718 66438
rect 115606 66510 115670 66574
rect 115062 66374 115126 66438
rect 115334 66374 115398 66438
rect 115878 66510 115942 66574
rect 116014 66374 116078 66438
rect 20950 66102 21014 66166
rect 1230 65966 1294 66030
rect 20814 65966 20878 66030
rect 21358 66102 21422 66166
rect 21494 66102 21558 66166
rect 21766 65966 21830 66030
rect 22174 66102 22238 66166
rect 22038 65966 22102 66030
rect 22582 66102 22646 66166
rect 22582 65966 22646 66030
rect 20814 65694 20878 65758
rect 20950 65558 21014 65622
rect 21766 65694 21830 65758
rect 21358 65558 21422 65622
rect 21494 65558 21558 65622
rect 22038 65694 22102 65758
rect 22038 65558 22102 65622
rect 22582 65694 22646 65758
rect 22446 65558 22510 65622
rect 20950 65286 21014 65350
rect 21358 65286 21422 65350
rect 21494 65286 21558 65350
rect 21902 65150 21966 65214
rect 22038 65286 22102 65350
rect 22174 65150 22238 65214
rect 22446 65286 22510 65350
rect 114246 66102 114310 66166
rect 114382 65966 114446 66030
rect 114654 66102 114718 66166
rect 114654 65966 114718 66030
rect 115062 66102 115126 66166
rect 115334 66102 115398 66166
rect 115606 65966 115670 66030
rect 116014 66102 116078 66166
rect 116014 65966 116078 66030
rect 135326 65830 135390 65894
rect 114382 65694 114446 65758
rect 114382 65558 114446 65622
rect 114654 65694 114718 65758
rect 114654 65558 114718 65622
rect 115606 65694 115670 65758
rect 115198 65558 115262 65622
rect 115334 65558 115398 65622
rect 116014 65694 116078 65758
rect 115878 65558 115942 65622
rect 22446 65150 22510 65214
rect 22038 65014 22102 65078
rect 27614 65014 27678 65078
rect 114382 65286 114446 65350
rect 114246 65150 114310 65214
rect 114654 65286 114718 65350
rect 114654 65150 114718 65214
rect 115198 65286 115262 65350
rect 115334 65286 115398 65350
rect 115062 65150 115126 65214
rect 115470 65150 115534 65214
rect 115878 65286 115942 65350
rect 21902 64878 21966 64942
rect 22174 64878 22238 64942
rect 22174 64742 22238 64806
rect 22446 64878 22510 64942
rect 22582 64742 22646 64806
rect 27614 64742 27678 64806
rect 1230 64062 1294 64126
rect 21766 64334 21830 64398
rect 22038 64470 22102 64534
rect 22174 64470 22238 64534
rect 22582 64470 22646 64534
rect 27342 64470 27406 64534
rect 109350 64742 109414 64806
rect 114246 64878 114310 64942
rect 114382 64742 114446 64806
rect 114654 64878 114718 64942
rect 114654 64742 114718 64806
rect 115062 64878 115126 64942
rect 115470 64878 115534 64942
rect 114382 64470 114446 64534
rect 20814 64062 20878 64126
rect 21766 64062 21830 64126
rect 20814 63790 20878 63854
rect 20814 63654 20878 63718
rect 21902 63654 21966 63718
rect 27342 64198 27406 64262
rect 27614 64198 27678 64262
rect 109350 64334 109414 64398
rect 109486 64198 109550 64262
rect 27614 63926 27678 63990
rect 109214 63926 109278 63990
rect 109486 63926 109550 63990
rect 27478 63790 27542 63854
rect 109350 63790 109414 63854
rect 114654 64470 114718 64534
rect 115334 64334 115398 64398
rect 136006 64470 136070 64534
rect 115334 64062 115398 64126
rect 132606 64334 132670 64398
rect 133422 64198 133486 64262
rect 116014 64062 116078 64126
rect 135326 64062 135390 64126
rect 20814 63382 20878 63446
rect 20814 63246 20878 63310
rect 21902 63382 21966 63446
rect 22038 63246 22102 63310
rect 22582 63246 22646 63310
rect 27478 63518 27542 63582
rect 109214 63518 109278 63582
rect 109350 63518 109414 63582
rect 115470 63654 115534 63718
rect 116014 63790 116078 63854
rect 115878 63654 115942 63718
rect 114246 63246 114310 63310
rect 114790 63246 114854 63310
rect 20814 62974 20878 63038
rect 20814 62838 20878 62902
rect 21766 62838 21830 62902
rect 22038 62974 22102 63038
rect 22038 62838 22102 62902
rect 22582 62974 22646 63038
rect 115470 63382 115534 63446
rect 115878 63382 115942 63446
rect 116014 63246 116078 63310
rect 22446 62838 22510 62902
rect 1230 62566 1294 62630
rect 20814 62566 20878 62630
rect 20814 62430 20878 62494
rect 21222 62430 21286 62494
rect 21766 62566 21830 62630
rect 21630 62430 21694 62494
rect 22038 62566 22102 62630
rect 22038 62430 22102 62494
rect 22446 62566 22510 62630
rect 22582 62430 22646 62494
rect 114246 62974 114310 63038
rect 114246 62838 114310 62902
rect 114790 62974 114854 63038
rect 114654 62838 114718 62902
rect 115062 62838 115126 62902
rect 115470 62838 115534 62902
rect 116014 62974 116078 63038
rect 115878 62838 115942 62902
rect 109350 62566 109414 62630
rect 114246 62566 114310 62630
rect 114382 62430 114446 62494
rect 114654 62566 114718 62630
rect 114790 62430 114854 62494
rect 115062 62566 115126 62630
rect 115198 62430 115262 62494
rect 115470 62566 115534 62630
rect 115878 62566 115942 62630
rect 115878 62430 115942 62494
rect 135326 62430 135390 62494
rect 20814 62158 20878 62222
rect 20950 62022 21014 62086
rect 21222 62158 21286 62222
rect 21358 62022 21422 62086
rect 21630 62158 21694 62222
rect 22038 62158 22102 62222
rect 22174 62022 22238 62086
rect 22582 62158 22646 62222
rect 22446 62022 22510 62086
rect 109350 62294 109414 62358
rect 114382 62158 114446 62222
rect 114246 62022 114310 62086
rect 114790 62158 114854 62222
rect 114654 62022 114718 62086
rect 115198 62158 115262 62222
rect 115470 62022 115534 62086
rect 115878 62158 115942 62222
rect 116014 62022 116078 62086
rect 134093 62119 134157 62123
rect 134093 62063 134097 62119
rect 134097 62063 134153 62119
rect 134153 62063 134157 62119
rect 134093 62059 134157 62063
rect 20950 61750 21014 61814
rect 20950 61614 21014 61678
rect 21358 61750 21422 61814
rect 21766 61614 21830 61678
rect 22174 61750 22238 61814
rect 22038 61614 22102 61678
rect 22446 61750 22510 61814
rect 22446 61614 22510 61678
rect 114246 61750 114310 61814
rect 114246 61614 114310 61678
rect 114654 61750 114718 61814
rect 114654 61614 114718 61678
rect 115062 61614 115126 61678
rect 115470 61750 115534 61814
rect 115606 61614 115670 61678
rect 116014 61750 116078 61814
rect 115878 61614 115942 61678
rect 20950 61342 21014 61406
rect 21358 61206 21422 61270
rect 21766 61342 21830 61406
rect 22038 61342 22102 61406
rect 22174 61206 22238 61270
rect 22446 61342 22510 61406
rect 22446 61206 22510 61270
rect 1230 60934 1294 60998
rect 133422 61478 133486 61542
rect 114246 61342 114310 61406
rect 114246 61206 114310 61270
rect 114654 61342 114718 61406
rect 114654 61206 114718 61270
rect 115062 61342 115126 61406
rect 115606 61342 115670 61406
rect 115334 61206 115398 61270
rect 115878 61342 115942 61406
rect 109486 61070 109550 61134
rect 21358 60934 21422 60998
rect 22174 60934 22238 60998
rect 22174 60798 22238 60862
rect 22446 60934 22510 60998
rect 22582 60798 22646 60862
rect 21902 60390 21966 60454
rect 22174 60526 22238 60590
rect 22038 60390 22102 60454
rect 22582 60526 22646 60590
rect 109486 60798 109550 60862
rect 114246 60934 114310 60998
rect 114246 60798 114310 60862
rect 114654 60934 114718 60998
rect 114654 60798 114718 60862
rect 115334 60934 115398 60998
rect 135326 60798 135390 60862
rect 114246 60526 114310 60590
rect 22446 60390 22510 60454
rect 114382 60390 114446 60454
rect 114654 60526 114718 60590
rect 114654 60390 114718 60454
rect 115198 60390 115262 60454
rect 115334 60390 115398 60454
rect 20814 60118 20878 60182
rect 21902 60118 21966 60182
rect 22038 60118 22102 60182
rect 22446 60118 22510 60182
rect 20814 59846 20878 59910
rect 20814 59710 20878 59774
rect 21766 59710 21830 59774
rect 27342 59846 27406 59910
rect 114382 60118 114446 60182
rect 109486 59846 109550 59910
rect 20814 59438 20878 59502
rect 20814 59302 20878 59366
rect 1230 59166 1294 59230
rect 21766 59438 21830 59502
rect 22038 59302 22102 59366
rect 22446 59302 22510 59366
rect 27342 59574 27406 59638
rect 109486 59574 109550 59638
rect 114654 60118 114718 60182
rect 115198 60118 115262 60182
rect 115334 60118 115398 60182
rect 116014 60118 116078 60182
rect 115470 59710 115534 59774
rect 116014 59846 116078 59910
rect 116014 59710 116078 59774
rect 114382 59302 114446 59366
rect 114790 59302 114854 59366
rect 115470 59438 115534 59502
rect 116014 59438 116078 59502
rect 115878 59302 115942 59366
rect 20814 59030 20878 59094
rect 20814 58894 20878 58958
rect 21222 58894 21286 58958
rect 22038 59030 22102 59094
rect 22174 58894 22238 58958
rect 22446 59030 22510 59094
rect 22446 58894 22510 58958
rect 135326 59166 135390 59230
rect 114382 59030 114446 59094
rect 20814 58622 20878 58686
rect 20814 58486 20878 58550
rect 21222 58622 21286 58686
rect 21358 58486 21422 58550
rect 21766 58486 21830 58550
rect 22174 58622 22238 58686
rect 22174 58486 22238 58550
rect 22446 58622 22510 58686
rect 22446 58486 22510 58550
rect 27614 58622 27678 58686
rect 114382 58894 114446 58958
rect 114790 59030 114854 59094
rect 114790 58894 114854 58958
rect 115470 58894 115534 58958
rect 115878 59030 115942 59094
rect 115878 58894 115942 58958
rect 109486 58622 109550 58686
rect 114382 58622 114446 58686
rect 114246 58486 114310 58550
rect 114790 58622 114854 58686
rect 114790 58486 114854 58550
rect 115470 58622 115534 58686
rect 115062 58486 115126 58550
rect 115334 58486 115398 58550
rect 115878 58622 115942 58686
rect 116014 58486 116078 58550
rect 27614 58350 27678 58414
rect 20814 58214 20878 58278
rect 20950 58078 21014 58142
rect 21358 58214 21422 58278
rect 21766 58214 21830 58278
rect 21494 58078 21558 58142
rect 22174 58214 22238 58278
rect 22038 58078 22102 58142
rect 22446 58214 22510 58278
rect 22446 58078 22510 58142
rect 109486 58350 109550 58414
rect 114246 58214 114310 58278
rect 114382 58078 114446 58142
rect 114790 58214 114854 58278
rect 114790 58078 114854 58142
rect 115062 58214 115126 58278
rect 115334 58214 115398 58278
rect 115198 58078 115262 58142
rect 115334 58078 115398 58142
rect 116014 58214 116078 58278
rect 115878 58078 115942 58142
rect 20950 57806 21014 57870
rect 20814 57670 20878 57734
rect 21494 57806 21558 57870
rect 22038 57806 22102 57870
rect 22174 57670 22238 57734
rect 22446 57806 22510 57870
rect 22582 57670 22646 57734
rect 114382 57806 114446 57870
rect 114246 57670 114310 57734
rect 114790 57806 114854 57870
rect 114654 57670 114718 57734
rect 115198 57806 115262 57870
rect 115334 57806 115398 57870
rect 115606 57670 115670 57734
rect 115878 57806 115942 57870
rect 116014 57670 116078 57734
rect 1230 57534 1294 57598
rect 20814 57398 20878 57462
rect 21222 57262 21286 57326
rect 21766 57262 21830 57326
rect 22174 57398 22238 57462
rect 22038 57262 22102 57326
rect 22582 57398 22646 57462
rect 135326 57534 135390 57598
rect 22446 57262 22510 57326
rect 114246 57398 114310 57462
rect 114246 57262 114310 57326
rect 114654 57398 114718 57462
rect 114654 57262 114718 57326
rect 115198 57262 115262 57326
rect 115606 57398 115670 57462
rect 115606 57262 115670 57326
rect 116014 57398 116078 57462
rect 21222 56990 21286 57054
rect 21766 56990 21830 57054
rect 22038 56990 22102 57054
rect 22038 56854 22102 56918
rect 22446 56990 22510 57054
rect 22446 56854 22510 56918
rect 114246 56990 114310 57054
rect 114246 56854 114310 56918
rect 114654 56990 114718 57054
rect 114790 56854 114854 56918
rect 115198 56990 115262 57054
rect 115606 56990 115670 57054
rect 21358 56446 21422 56510
rect 21630 56446 21694 56510
rect 22038 56582 22102 56646
rect 22174 56446 22238 56510
rect 22446 56582 22510 56646
rect 114246 56582 114310 56646
rect 22446 56446 22510 56510
rect 114246 56446 114310 56510
rect 114790 56582 114854 56646
rect 114654 56446 114718 56510
rect 115062 56446 115126 56510
rect 20950 56174 21014 56238
rect 21358 56174 21422 56238
rect 21630 56174 21694 56238
rect 1230 55902 1294 55966
rect 20950 55902 21014 55966
rect 20814 55766 20878 55830
rect 21494 55766 21558 55830
rect 22174 56174 22238 56238
rect 22446 56174 22510 56238
rect 27478 55902 27542 55966
rect 109350 56038 109414 56102
rect 114246 56174 114310 56238
rect 114654 56174 114718 56238
rect 115062 56174 115126 56238
rect 116014 56174 116078 56238
rect 115334 56038 115398 56102
rect 109486 55902 109550 55966
rect 20814 55494 20878 55558
rect 20950 55358 21014 55422
rect 21494 55494 21558 55558
rect 27478 55494 27542 55558
rect 27614 55494 27678 55558
rect 27614 55222 27678 55286
rect 20950 55086 21014 55150
rect 20814 54950 20878 55014
rect 21630 54950 21694 55014
rect 22038 54950 22102 55014
rect 109350 55630 109414 55694
rect 109486 55630 109550 55694
rect 109486 55494 109550 55558
rect 109486 55222 109550 55286
rect 22446 54950 22510 55014
rect 20814 54678 20878 54742
rect 20950 54542 21014 54606
rect 21630 54678 21694 54742
rect 21358 54542 21422 54606
rect 21494 54542 21558 54606
rect 22038 54678 22102 54742
rect 22174 54542 22238 54606
rect 22446 54678 22510 54742
rect 22582 54542 22646 54606
rect 20950 54270 21014 54334
rect 1230 54134 1294 54198
rect 20814 54134 20878 54198
rect 21358 54270 21422 54334
rect 21494 54270 21558 54334
rect 21766 54134 21830 54198
rect 22174 54270 22238 54334
rect 22174 54134 22238 54198
rect 22582 54270 22646 54334
rect 115198 55902 115262 55966
rect 115334 55766 115398 55830
rect 116014 55902 116078 55966
rect 116014 55766 116078 55830
rect 135326 55902 135390 55966
rect 115334 55494 115398 55558
rect 116014 55494 116078 55558
rect 116014 55358 116078 55422
rect 114382 54950 114446 55014
rect 114790 54950 114854 55014
rect 115198 54950 115262 55014
rect 115334 54950 115398 55014
rect 116014 55086 116078 55150
rect 115878 54950 115942 55014
rect 114382 54678 114446 54742
rect 114246 54542 114310 54606
rect 114790 54678 114854 54742
rect 114790 54542 114854 54606
rect 115198 54678 115262 54742
rect 115334 54678 115398 54742
rect 115470 54542 115534 54606
rect 115878 54678 115942 54742
rect 116014 54542 116078 54606
rect 22446 54134 22510 54198
rect 114246 54270 114310 54334
rect 114382 54134 114446 54198
rect 114790 54270 114854 54334
rect 114790 54134 114854 54198
rect 115470 54270 115534 54334
rect 115198 54134 115262 54198
rect 115334 54134 115398 54198
rect 116014 54270 116078 54334
rect 116014 54134 116078 54198
rect 135326 53998 135390 54062
rect 20814 53862 20878 53926
rect 20814 53726 20878 53790
rect 21766 53862 21830 53926
rect 21630 53726 21694 53790
rect 22174 53862 22238 53926
rect 22038 53726 22102 53790
rect 22446 53862 22510 53926
rect 22446 53726 22510 53790
rect 114382 53862 114446 53926
rect 114382 53726 114446 53790
rect 114790 53862 114854 53926
rect 114790 53726 114854 53790
rect 115198 53862 115262 53926
rect 115334 53862 115398 53926
rect 116014 53862 116078 53926
rect 115878 53726 115942 53790
rect 20814 53454 20878 53518
rect 21630 53454 21694 53518
rect 21358 53318 21422 53382
rect 21494 53318 21558 53382
rect 22038 53454 22102 53518
rect 22174 53318 22238 53382
rect 22446 53454 22510 53518
rect 22446 53318 22510 53382
rect 114382 53454 114446 53518
rect 114246 53318 114310 53382
rect 114790 53454 114854 53518
rect 114654 53318 114718 53382
rect 115470 53318 115534 53382
rect 115878 53454 115942 53518
rect 20950 52910 21014 52974
rect 21358 53046 21422 53110
rect 21494 53046 21558 53110
rect 21222 52910 21286 52974
rect 21766 52910 21830 52974
rect 22174 53046 22238 53110
rect 22174 52910 22238 52974
rect 22446 53046 22510 53110
rect 22582 52910 22646 52974
rect 114246 53046 114310 53110
rect 114246 52910 114310 52974
rect 114654 53046 114718 53110
rect 114790 52910 114854 52974
rect 115198 52910 115262 52974
rect 115470 53046 115534 53110
rect 115606 52910 115670 52974
rect 115878 52910 115942 52974
rect 20950 52638 21014 52702
rect 1230 52502 1294 52566
rect 21222 52638 21286 52702
rect 21766 52638 21830 52702
rect 22174 52638 22238 52702
rect 22174 52502 22238 52566
rect 22582 52638 22646 52702
rect 22446 52502 22510 52566
rect 27478 52366 27542 52430
rect 114246 52638 114310 52702
rect 114382 52502 114446 52566
rect 114790 52638 114854 52702
rect 114790 52502 114854 52566
rect 115198 52638 115262 52702
rect 115606 52638 115670 52702
rect 115198 52502 115262 52566
rect 115878 52638 115942 52702
rect 20814 52230 20878 52294
rect 22174 52230 22238 52294
rect 22174 52094 22238 52158
rect 22446 52230 22510 52294
rect 22582 52094 22646 52158
rect 27478 52094 27542 52158
rect 20814 51958 20878 52022
rect 21766 51686 21830 51750
rect 22174 51822 22238 51886
rect 22582 51822 22646 51886
rect 20814 51414 20878 51478
rect 21766 51414 21830 51478
rect 27342 51278 27406 51342
rect 20814 51142 20878 51206
rect 20814 51006 20878 51070
rect 21358 51006 21422 51070
rect 21902 51006 21966 51070
rect 22174 51006 22238 51070
rect 22582 51006 22646 51070
rect 27342 51006 27406 51070
rect 1230 50870 1294 50934
rect 20814 50734 20878 50798
rect 20814 50598 20878 50662
rect 21358 50734 21422 50798
rect 21902 50734 21966 50798
rect 21902 50598 21966 50662
rect 22174 50734 22238 50798
rect 22038 50598 22102 50662
rect 22582 50734 22646 50798
rect 22446 50598 22510 50662
rect 114382 52230 114446 52294
rect 114246 52094 114310 52158
rect 114790 52230 114854 52294
rect 114654 52094 114718 52158
rect 115198 52230 115262 52294
rect 135326 52366 135390 52430
rect 116014 52230 116078 52294
rect 114246 51822 114310 51886
rect 114654 51822 114718 51886
rect 115198 51686 115262 51750
rect 116014 51958 116078 52022
rect 115198 51414 115262 51478
rect 115878 51414 115942 51478
rect 114246 51006 114310 51070
rect 114654 51006 114718 51070
rect 115062 51006 115126 51070
rect 115470 51006 115534 51070
rect 115878 51142 115942 51206
rect 116014 51006 116078 51070
rect 114246 50734 114310 50798
rect 114382 50598 114446 50662
rect 114654 50734 114718 50798
rect 114790 50598 114854 50662
rect 115062 50734 115126 50798
rect 115470 50734 115534 50798
rect 116014 50734 116078 50798
rect 135326 50734 135390 50798
rect 115878 50598 115942 50662
rect 20814 50326 20878 50390
rect 20950 50190 21014 50254
rect 21902 50326 21966 50390
rect 21222 50190 21286 50254
rect 21494 50190 21558 50254
rect 22038 50326 22102 50390
rect 22174 50190 22238 50254
rect 22446 50326 22510 50390
rect 22582 50190 22646 50254
rect 114382 50326 114446 50390
rect 114246 50190 114310 50254
rect 114790 50326 114854 50390
rect 114790 50190 114854 50254
rect 115606 50190 115670 50254
rect 115878 50326 115942 50390
rect 115878 50190 115942 50254
rect 20950 49918 21014 49982
rect 20814 49782 20878 49846
rect 21222 49918 21286 49982
rect 21494 49918 21558 49982
rect 21766 49782 21830 49846
rect 22174 49918 22238 49982
rect 22174 49782 22238 49846
rect 22582 49918 22646 49982
rect 22446 49782 22510 49846
rect 114246 49918 114310 49982
rect 114246 49782 114310 49846
rect 114790 49918 114854 49982
rect 114654 49782 114718 49846
rect 115606 49918 115670 49982
rect 115198 49782 115262 49846
rect 115334 49782 115398 49846
rect 115878 49918 115942 49982
rect 115878 49782 115942 49846
rect 20814 49510 20878 49574
rect 20950 49374 21014 49438
rect 21222 49374 21286 49438
rect 21766 49510 21830 49574
rect 21630 49374 21694 49438
rect 22174 49510 22238 49574
rect 22038 49374 22102 49438
rect 22446 49510 22510 49574
rect 22446 49374 22510 49438
rect 114246 49510 114310 49574
rect 114382 49374 114446 49438
rect 114654 49510 114718 49574
rect 114654 49374 114718 49438
rect 115198 49510 115262 49574
rect 115334 49510 115398 49574
rect 115878 49510 115942 49574
rect 115878 49374 115942 49438
rect 1230 48966 1294 49030
rect 20950 49102 21014 49166
rect 20814 48966 20878 49030
rect 21222 49102 21286 49166
rect 21630 49102 21694 49166
rect 21358 48966 21422 49030
rect 21494 48966 21558 49030
rect 22038 49102 22102 49166
rect 22174 48966 22238 49030
rect 22446 49102 22510 49166
rect 22582 48966 22646 49030
rect 114382 49102 114446 49166
rect 114246 48966 114310 49030
rect 114654 49102 114718 49166
rect 114654 48966 114718 49030
rect 115606 48966 115670 49030
rect 115878 49102 115942 49166
rect 116014 48966 116078 49030
rect 135326 48966 135390 49030
rect 20814 48694 20878 48758
rect 21358 48694 21422 48758
rect 21494 48694 21558 48758
rect 21766 48558 21830 48622
rect 22174 48694 22238 48758
rect 22174 48558 22238 48622
rect 22582 48694 22646 48758
rect 22446 48558 22510 48622
rect 114246 48694 114310 48758
rect 114382 48558 114446 48622
rect 114654 48694 114718 48758
rect 114654 48558 114718 48622
rect 115062 48558 115126 48622
rect 115606 48694 115670 48758
rect 115470 48558 115534 48622
rect 116014 48694 116078 48758
rect 20814 48286 20878 48350
rect 21766 48286 21830 48350
rect 22174 48286 22238 48350
rect 22174 48150 22238 48214
rect 22446 48286 22510 48350
rect 22446 48150 22510 48214
rect 20814 48014 20878 48078
rect 21494 47742 21558 47806
rect 22174 47878 22238 47942
rect 1230 47470 1294 47534
rect 20814 47470 20878 47534
rect 21494 47470 21558 47534
rect 22446 47878 22510 47942
rect 114382 48286 114446 48350
rect 114246 48150 114310 48214
rect 114654 48286 114718 48350
rect 114790 48150 114854 48214
rect 115062 48286 115126 48350
rect 115334 48286 115398 48350
rect 115470 48286 115534 48350
rect 115878 48286 115942 48350
rect 114246 47878 114310 47942
rect 20814 47198 20878 47262
rect 20950 47062 21014 47126
rect 21358 47062 21422 47126
rect 21766 47062 21830 47126
rect 20950 46790 21014 46854
rect 20814 46654 20878 46718
rect 21358 46790 21422 46854
rect 21766 46790 21830 46854
rect 22174 46654 22238 46718
rect 27342 47198 27406 47262
rect 114790 47878 114854 47942
rect 115334 48014 115398 48078
rect 115062 47742 115126 47806
rect 115878 48014 115942 48078
rect 115062 47470 115126 47534
rect 115878 47470 115942 47534
rect 135326 47470 135390 47534
rect 109350 47198 109414 47262
rect 27342 46926 27406 46990
rect 22582 46654 22646 46718
rect 27342 46790 27406 46854
rect 109350 46926 109414 46990
rect 109486 46790 109550 46854
rect 115334 47062 115398 47126
rect 115878 47198 115942 47262
rect 115878 47062 115942 47126
rect 114246 46654 114310 46718
rect 114654 46654 114718 46718
rect 27342 46518 27406 46582
rect 20814 46382 20878 46446
rect 20950 46246 21014 46310
rect 21222 46246 21286 46310
rect 22174 46382 22238 46446
rect 22038 46246 22102 46310
rect 22582 46382 22646 46446
rect 109486 46518 109550 46582
rect 115334 46790 115398 46854
rect 115878 46790 115942 46854
rect 116014 46654 116078 46718
rect 22582 46246 22646 46310
rect 114246 46382 114310 46446
rect 114382 46246 114446 46310
rect 114654 46382 114718 46446
rect 114790 46246 114854 46310
rect 115198 46246 115262 46310
rect 115334 46246 115398 46310
rect 115470 46246 115534 46310
rect 116014 46382 116078 46446
rect 115878 46246 115942 46310
rect 20950 45974 21014 46038
rect 20950 45838 21014 45902
rect 21222 45974 21286 46038
rect 21358 45838 21422 45902
rect 22038 45974 22102 46038
rect 22038 45838 22102 45902
rect 22582 45974 22646 46038
rect 22446 45838 22510 45902
rect 114382 45974 114446 46038
rect 114382 45838 114446 45902
rect 114790 45974 114854 46038
rect 115198 45974 115262 46038
rect 115334 45974 115398 46038
rect 115470 45974 115534 46038
rect 114654 45838 114718 45902
rect 115470 45838 115534 45902
rect 115878 45974 115942 46038
rect 116014 45838 116078 45902
rect 1230 45566 1294 45630
rect 20950 45566 21014 45630
rect 20814 45430 20878 45494
rect 21358 45566 21422 45630
rect 21766 45430 21830 45494
rect 22038 45566 22102 45630
rect 22446 45566 22510 45630
rect 22038 45430 22102 45494
rect 135326 45702 135390 45766
rect 114382 45566 114446 45630
rect 22446 45430 22510 45494
rect 25846 45430 25910 45494
rect 113702 45430 113766 45494
rect 114382 45430 114446 45494
rect 114654 45566 114718 45630
rect 114790 45430 114854 45494
rect 115470 45566 115534 45630
rect 115198 45430 115262 45494
rect 115334 45430 115398 45494
rect 116014 45566 116078 45630
rect 115878 45430 115942 45494
rect 20814 45158 20878 45222
rect 20950 45022 21014 45086
rect 21766 45158 21830 45222
rect 21222 45022 21286 45086
rect 21494 45022 21558 45086
rect 22038 45158 22102 45222
rect 22038 45022 22102 45086
rect 22446 45158 22510 45222
rect 22582 45022 22646 45086
rect 25846 45158 25910 45222
rect 23262 45022 23326 45086
rect 113702 45158 113766 45222
rect 114382 45158 114446 45222
rect 112342 45022 112406 45086
rect 114382 45022 114446 45086
rect 114790 45158 114854 45222
rect 114654 45022 114718 45086
rect 115198 45158 115262 45222
rect 115334 45158 115398 45222
rect 115878 45158 115942 45222
rect 115878 45022 115942 45086
rect 20950 44750 21014 44814
rect 21222 44750 21286 44814
rect 21494 44750 21558 44814
rect 21358 44614 21422 44678
rect 22038 44750 22102 44814
rect 22174 44614 22238 44678
rect 22582 44750 22646 44814
rect 23262 44750 23326 44814
rect 114382 44750 114446 44814
rect 22446 44614 22510 44678
rect 112342 44614 112406 44678
rect 114246 44614 114310 44678
rect 114654 44750 114718 44814
rect 114654 44614 114718 44678
rect 115470 44614 115534 44678
rect 115878 44750 115942 44814
rect 21358 44342 21422 44406
rect 22174 44342 22238 44406
rect 22174 44206 22238 44270
rect 22446 44342 22510 44406
rect 22582 44206 22646 44270
rect 1230 44070 1294 44134
rect 21766 43798 21830 43862
rect 22174 43934 22238 43998
rect 22038 43798 22102 43862
rect 22582 43934 22646 43998
rect 22446 43798 22510 43862
rect 27478 43662 27542 43726
rect 114246 44342 114310 44406
rect 114382 44206 114446 44270
rect 114654 44342 114718 44406
rect 114790 44206 114854 44270
rect 115470 44342 115534 44406
rect 114382 43934 114446 43998
rect 114382 43798 114446 43862
rect 114790 43934 114854 43998
rect 114790 43798 114854 43862
rect 115198 43798 115262 43862
rect 135326 43934 135390 43998
rect 109350 43662 109414 43726
rect 20814 43526 20878 43590
rect 21766 43526 21830 43590
rect 21630 43390 21694 43454
rect 22038 43526 22102 43590
rect 20814 43254 20878 43318
rect 20814 43118 20878 43182
rect 21222 43118 21286 43182
rect 21494 43118 21558 43182
rect 22446 43526 22510 43590
rect 27478 43390 27542 43454
rect 27614 43254 27678 43318
rect 109350 43390 109414 43454
rect 109350 43254 109414 43318
rect 114382 43526 114446 43590
rect 114790 43526 114854 43590
rect 115198 43526 115262 43590
rect 116014 43526 116078 43590
rect 20814 42846 20878 42910
rect 20814 42710 20878 42774
rect 21222 42846 21286 42910
rect 22174 42710 22238 42774
rect 22446 42710 22510 42774
rect 27614 42982 27678 43046
rect 109350 42982 109414 43046
rect 109350 42846 109414 42910
rect 115062 43118 115126 43182
rect 116014 43254 116078 43318
rect 116014 43118 116078 43182
rect 114246 42710 114310 42774
rect 114790 42710 114854 42774
rect 115062 42846 115126 42910
rect 1230 42438 1294 42502
rect 20814 42438 20878 42502
rect 20950 42302 21014 42366
rect 21766 42302 21830 42366
rect 22174 42438 22238 42502
rect 22174 42302 22238 42366
rect 22446 42438 22510 42502
rect 109350 42574 109414 42638
rect 116014 42846 116078 42910
rect 115878 42710 115942 42774
rect 114246 42438 114310 42502
rect 22582 42302 22646 42366
rect 20950 42030 21014 42094
rect 20814 41894 20878 41958
rect 21222 41894 21286 41958
rect 21766 42030 21830 42094
rect 21630 41894 21694 41958
rect 22174 42030 22238 42094
rect 22038 41894 22102 41958
rect 22582 42030 22646 42094
rect 22446 41894 22510 41958
rect 20814 41622 20878 41686
rect 20814 41486 20878 41550
rect 21222 41622 21286 41686
rect 21358 41486 21422 41550
rect 21630 41622 21694 41686
rect 22038 41622 22102 41686
rect 22038 41486 22102 41550
rect 22446 41622 22510 41686
rect 22582 41486 22646 41550
rect 114246 42302 114310 42366
rect 114790 42438 114854 42502
rect 114654 42302 114718 42366
rect 115062 42302 115126 42366
rect 115878 42438 115942 42502
rect 116014 42302 116078 42366
rect 135326 42302 135390 42366
rect 114246 42030 114310 42094
rect 114382 41894 114446 41958
rect 114654 42030 114718 42094
rect 114790 41894 114854 41958
rect 115062 42030 115126 42094
rect 115198 41894 115262 41958
rect 115334 41894 115398 41958
rect 116014 42030 116078 42094
rect 115878 41894 115942 41958
rect 114382 41622 114446 41686
rect 114382 41486 114446 41550
rect 114790 41622 114854 41686
rect 114790 41486 114854 41550
rect 115198 41622 115262 41686
rect 115334 41622 115398 41686
rect 115606 41486 115670 41550
rect 115878 41622 115942 41686
rect 116014 41486 116078 41550
rect 20814 41214 20878 41278
rect 20814 41078 20878 41142
rect 21358 41214 21422 41278
rect 21766 41078 21830 41142
rect 22038 41214 22102 41278
rect 22038 41078 22102 41142
rect 22582 41214 22646 41278
rect 22446 41078 22510 41142
rect 114382 41214 114446 41278
rect 114382 41078 114446 41142
rect 114790 41214 114854 41278
rect 114654 41078 114718 41142
rect 115606 41214 115670 41278
rect 115198 41078 115262 41142
rect 115334 41078 115398 41142
rect 115470 41078 115534 41142
rect 116014 41214 116078 41278
rect 116014 41078 116078 41142
rect 1230 40806 1294 40870
rect 20814 40806 20878 40870
rect 21222 40670 21286 40734
rect 21766 40806 21830 40870
rect 21630 40670 21694 40734
rect 22038 40806 22102 40870
rect 22038 40670 22102 40734
rect 22446 40806 22510 40870
rect 22582 40670 22646 40734
rect 114382 40806 114446 40870
rect 27478 40534 27542 40598
rect 114382 40670 114446 40734
rect 114654 40806 114718 40870
rect 114654 40670 114718 40734
rect 115198 40806 115262 40870
rect 115334 40806 115398 40870
rect 115470 40806 115534 40870
rect 115334 40670 115398 40734
rect 116014 40806 116078 40870
rect 135326 40806 135390 40870
rect 109486 40534 109550 40598
rect 21222 40398 21286 40462
rect 21630 40398 21694 40462
rect 22038 40398 22102 40462
rect 22174 40262 22238 40326
rect 22582 40398 22646 40462
rect 22446 40262 22510 40326
rect 27478 40262 27542 40326
rect 21766 39854 21830 39918
rect 22174 39990 22238 40054
rect 22038 39854 22102 39918
rect 22446 39990 22510 40054
rect 109350 40262 109414 40326
rect 109486 40262 109550 40326
rect 114382 40398 114446 40462
rect 114246 40262 114310 40326
rect 114654 40398 114718 40462
rect 114654 40262 114718 40326
rect 115334 40398 115398 40462
rect 115198 40262 115262 40326
rect 114246 39990 114310 40054
rect 22582 39854 22646 39918
rect 20814 39582 20878 39646
rect 21766 39582 21830 39646
rect 20814 39310 20878 39374
rect 20814 39174 20878 39238
rect 21494 39174 21558 39238
rect 22038 39582 22102 39646
rect 22582 39582 22646 39646
rect 1230 39038 1294 39102
rect 27478 39310 27542 39374
rect 109350 39854 109414 39918
rect 114246 39854 114310 39918
rect 114654 39990 114718 40054
rect 114654 39854 114718 39918
rect 115334 40126 115398 40190
rect 115198 39854 115262 39918
rect 114246 39582 114310 39646
rect 114654 39582 114718 39646
rect 115198 39582 115262 39646
rect 115878 39582 115942 39646
rect 109486 39310 109550 39374
rect 27478 39038 27542 39102
rect 20814 38902 20878 38966
rect 20814 38766 20878 38830
rect 21494 38902 21558 38966
rect 20814 38494 20878 38558
rect 20814 38358 20878 38422
rect 21358 38358 21422 38422
rect 22038 38358 22102 38422
rect 109486 39038 109550 39102
rect 115470 39174 115534 39238
rect 115878 39310 115942 39374
rect 116014 39174 116078 39238
rect 135326 39038 135390 39102
rect 115470 38902 115534 38966
rect 116014 38902 116078 38966
rect 116014 38766 116078 38830
rect 22446 38358 22510 38422
rect 20814 38086 20878 38150
rect 20950 37950 21014 38014
rect 21358 38086 21422 38150
rect 21766 37950 21830 38014
rect 22038 38086 22102 38150
rect 22174 37950 22238 38014
rect 22446 38086 22510 38150
rect 22446 37950 22510 38014
rect 27342 38086 27406 38150
rect 114382 38358 114446 38422
rect 114654 38358 114718 38422
rect 115198 38358 115262 38422
rect 115334 38358 115398 38422
rect 116014 38494 116078 38558
rect 115878 38358 115942 38422
rect 109486 38086 109550 38150
rect 114382 38086 114446 38150
rect 114246 37950 114310 38014
rect 114654 38086 114718 38150
rect 114654 37950 114718 38014
rect 115198 38086 115262 38150
rect 115334 38086 115398 38150
rect 115062 37950 115126 38014
rect 115470 37950 115534 38014
rect 115878 38086 115942 38150
rect 116014 37950 116078 38014
rect 27342 37814 27406 37878
rect 14150 37542 14214 37606
rect 20950 37678 21014 37742
rect 20814 37542 20878 37606
rect 21222 37542 21286 37606
rect 21766 37678 21830 37742
rect 21630 37542 21694 37606
rect 22174 37678 22238 37742
rect 22038 37542 22102 37606
rect 22446 37678 22510 37742
rect 22582 37542 22646 37606
rect 1230 37270 1294 37334
rect 109486 37814 109550 37878
rect 114246 37678 114310 37742
rect 114382 37542 114446 37606
rect 114654 37678 114718 37742
rect 114790 37542 114854 37606
rect 115062 37678 115126 37742
rect 115470 37678 115534 37742
rect 116014 37678 116078 37742
rect 115878 37542 115942 37606
rect 135326 37406 135390 37470
rect 20814 37270 20878 37334
rect 20814 37134 20878 37198
rect 21222 37270 21286 37334
rect 21630 37270 21694 37334
rect 21358 37134 21422 37198
rect 21494 37134 21558 37198
rect 22038 37270 22102 37334
rect 22174 37134 22238 37198
rect 22582 37270 22646 37334
rect 22582 37134 22646 37198
rect 20814 36862 20878 36926
rect 21358 36862 21422 36926
rect 21494 36862 21558 36926
rect 21766 36726 21830 36790
rect 22174 36862 22238 36926
rect 22038 36726 22102 36790
rect 22582 36862 22646 36926
rect 114382 37270 114446 37334
rect 114246 37134 114310 37198
rect 114790 37270 114854 37334
rect 114790 37134 114854 37198
rect 115606 37134 115670 37198
rect 115878 37270 115942 37334
rect 115878 37134 115942 37198
rect 22446 36726 22510 36790
rect 114246 36862 114310 36926
rect 114246 36726 114310 36790
rect 114790 36862 114854 36926
rect 114654 36726 114718 36790
rect 115198 36726 115262 36790
rect 115606 36862 115670 36926
rect 115470 36726 115534 36790
rect 115878 36862 115942 36926
rect 20950 36318 21014 36382
rect 21766 36454 21830 36518
rect 21494 36318 21558 36382
rect 21630 36318 21694 36382
rect 22038 36454 22102 36518
rect 22038 36318 22102 36382
rect 22446 36454 22510 36518
rect 22446 36318 22510 36382
rect 114246 36454 114310 36518
rect 114382 36318 114446 36382
rect 114654 36454 114718 36518
rect 114790 36318 114854 36382
rect 115198 36454 115262 36518
rect 115470 36454 115534 36518
rect 115198 36318 115262 36382
rect 115334 36318 115398 36382
rect 116014 36318 116078 36382
rect 14286 36182 14350 36246
rect 20950 36046 21014 36110
rect 21494 36046 21558 36110
rect 21630 36046 21694 36110
rect 21494 35910 21558 35974
rect 22038 36046 22102 36110
rect 22174 35910 22238 35974
rect 22446 36046 22510 36110
rect 22446 35910 22510 35974
rect 1230 35638 1294 35702
rect 114382 36046 114446 36110
rect 114246 35910 114310 35974
rect 114790 36046 114854 36110
rect 114654 35910 114718 35974
rect 115198 36046 115262 36110
rect 115334 36046 115398 36110
rect 115470 35910 115534 35974
rect 116014 36046 116078 36110
rect 20814 35638 20878 35702
rect 21494 35638 21558 35702
rect 21358 35502 21422 35566
rect 21630 35502 21694 35566
rect 22174 35638 22238 35702
rect 22446 35638 22510 35702
rect 114246 35638 114310 35702
rect 20814 35366 20878 35430
rect 20950 35230 21014 35294
rect 21902 35230 21966 35294
rect 27478 35230 27542 35294
rect 20950 34958 21014 35022
rect 14150 34822 14214 34886
rect 20814 34822 20878 34886
rect 21902 34822 21966 34886
rect 14014 34686 14078 34750
rect 20814 34550 20878 34614
rect 20814 34414 20878 34478
rect 21222 34414 21286 34478
rect 22038 34414 22102 34478
rect 27478 34958 27542 35022
rect 109350 34958 109414 35022
rect 109350 34686 109414 34750
rect 109486 34686 109550 34750
rect 114654 35638 114718 35702
rect 115470 35638 115534 35702
rect 115878 35638 115942 35702
rect 135326 35502 135390 35566
rect 115470 35230 115534 35294
rect 115878 35366 115942 35430
rect 115878 35230 115942 35294
rect 115878 34958 115942 35022
rect 22446 34414 22510 34478
rect 20814 34142 20878 34206
rect 1230 34006 1294 34070
rect 20814 34006 20878 34070
rect 21222 34142 21286 34206
rect 21358 34006 21422 34070
rect 22038 34142 22102 34206
rect 22038 34006 22102 34070
rect 22446 34142 22510 34206
rect 22446 34006 22510 34070
rect 109486 34414 109550 34478
rect 114246 34414 114310 34478
rect 114654 34414 114718 34478
rect 115470 34822 115534 34886
rect 116014 34822 116078 34886
rect 115198 34414 115262 34478
rect 115606 34414 115670 34478
rect 116014 34550 116078 34614
rect 116014 34414 116078 34478
rect 109486 34142 109550 34206
rect 114246 34142 114310 34206
rect 114246 34006 114310 34070
rect 114654 34142 114718 34206
rect 114790 34006 114854 34070
rect 115198 34142 115262 34206
rect 115606 34142 115670 34206
rect 115334 34006 115398 34070
rect 115606 34006 115670 34070
rect 116014 34142 116078 34206
rect 116014 34006 116078 34070
rect 20814 33734 20878 33798
rect 20814 33598 20878 33662
rect 21358 33734 21422 33798
rect 21358 33598 21422 33662
rect 21766 33598 21830 33662
rect 22038 33734 22102 33798
rect 22174 33598 22238 33662
rect 22446 33734 22510 33798
rect 109486 33870 109550 33934
rect 135326 33870 135390 33934
rect 22446 33598 22510 33662
rect 14286 33462 14350 33526
rect 114246 33734 114310 33798
rect 114246 33598 114310 33662
rect 114790 33734 114854 33798
rect 114654 33598 114718 33662
rect 115334 33734 115398 33798
rect 115606 33734 115670 33798
rect 115062 33598 115126 33662
rect 115606 33598 115670 33662
rect 116014 33734 116078 33798
rect 116014 33598 116078 33662
rect 14150 33326 14214 33390
rect 20814 33326 20878 33390
rect 20814 33190 20878 33254
rect 21358 33326 21422 33390
rect 21766 33326 21830 33390
rect 21630 33190 21694 33254
rect 22174 33326 22238 33390
rect 22038 33190 22102 33254
rect 22446 33326 22510 33390
rect 22446 33190 22510 33254
rect 114246 33326 114310 33390
rect 114382 33190 114446 33254
rect 114654 33326 114718 33390
rect 114790 33190 114854 33254
rect 115062 33326 115126 33390
rect 115198 33190 115262 33254
rect 115606 33326 115670 33390
rect 116014 33326 116078 33390
rect 115878 33190 115942 33254
rect 20814 32918 20878 32982
rect 20950 32782 21014 32846
rect 21222 32782 21286 32846
rect 21630 32918 21694 32982
rect 22038 32918 22102 32982
rect 22038 32782 22102 32846
rect 22446 32918 22510 32982
rect 22582 32782 22646 32846
rect 114382 32918 114446 32982
rect 114382 32782 114446 32846
rect 114790 32918 114854 32982
rect 114790 32782 114854 32846
rect 115198 32918 115262 32982
rect 115606 32782 115670 32846
rect 115878 32918 115942 32982
rect 115878 32782 115942 32846
rect 20950 32510 21014 32574
rect 1230 32374 1294 32438
rect 20950 32374 21014 32438
rect 21222 32510 21286 32574
rect 21766 32374 21830 32438
rect 22038 32510 22102 32574
rect 22038 32374 22102 32438
rect 22582 32510 22646 32574
rect 22446 32374 22510 32438
rect 114382 32510 114446 32574
rect 114246 32374 114310 32438
rect 114790 32510 114854 32574
rect 114654 32374 114718 32438
rect 115606 32510 115670 32574
rect 115198 32374 115262 32438
rect 115334 32374 115398 32438
rect 115878 32510 115942 32574
rect 115878 32374 115942 32438
rect 14014 32102 14078 32166
rect 20950 32102 21014 32166
rect 21222 31966 21286 32030
rect 21766 32102 21830 32166
rect 21630 31966 21694 32030
rect 22038 32102 22102 32166
rect 22038 31966 22102 32030
rect 22446 32102 22510 32166
rect 22582 31966 22646 32030
rect 135326 32238 135390 32302
rect 114246 32102 114310 32166
rect 14150 31830 14214 31894
rect 114382 31966 114446 32030
rect 114654 32102 114718 32166
rect 114790 31966 114854 32030
rect 115198 32102 115262 32166
rect 115334 32102 115398 32166
rect 115878 32102 115942 32166
rect 109486 31830 109550 31894
rect 20950 31694 21014 31758
rect 21222 31694 21286 31758
rect 21630 31694 21694 31758
rect 22038 31694 22102 31758
rect 22174 31558 22238 31622
rect 22582 31694 22646 31758
rect 22446 31558 22510 31622
rect 20950 31422 21014 31486
rect 21766 31150 21830 31214
rect 22174 31286 22238 31350
rect 22446 31286 22510 31350
rect 109350 31558 109414 31622
rect 109486 31558 109550 31622
rect 114382 31694 114446 31758
rect 114246 31558 114310 31622
rect 114790 31694 114854 31758
rect 114654 31558 114718 31622
rect 115878 31694 115942 31758
rect 114246 31286 114310 31350
rect 20814 30878 20878 30942
rect 21766 30878 21830 30942
rect 1230 30470 1294 30534
rect 14014 30606 14078 30670
rect 14014 30470 14078 30534
rect 20814 30606 20878 30670
rect 20814 30470 20878 30534
rect 21358 30470 21422 30534
rect 27342 31014 27406 31078
rect 27342 30742 27406 30806
rect 27478 30606 27542 30670
rect 109350 31150 109414 31214
rect 114654 31286 114718 31350
rect 115470 31150 115534 31214
rect 115878 31422 115942 31486
rect 109350 30606 109414 30670
rect 115470 30878 115534 30942
rect 115878 30878 115942 30942
rect 20814 30198 20878 30262
rect 20950 30062 21014 30126
rect 21358 30198 21422 30262
rect 20950 29790 21014 29854
rect 20814 29654 20878 29718
rect 22174 30062 22238 30126
rect 22582 30062 22646 30126
rect 27478 30334 27542 30398
rect 109350 30334 109414 30398
rect 109350 30198 109414 30262
rect 115470 30470 115534 30534
rect 115878 30606 115942 30670
rect 116014 30470 116078 30534
rect 135326 30470 135390 30534
rect 114246 30062 114310 30126
rect 114654 30062 114718 30126
rect 21494 29654 21558 29718
rect 21766 29654 21830 29718
rect 22174 29790 22238 29854
rect 22038 29654 22102 29718
rect 22582 29790 22646 29854
rect 22446 29654 22510 29718
rect 109350 29926 109414 29990
rect 114246 29790 114310 29854
rect 114246 29654 114310 29718
rect 114654 29790 114718 29854
rect 114654 29654 114718 29718
rect 115470 30198 115534 30262
rect 116014 30198 116078 30262
rect 115878 30062 115942 30126
rect 115334 29654 115398 29718
rect 115470 29654 115534 29718
rect 115878 29790 115942 29854
rect 115878 29654 115942 29718
rect 20814 29382 20878 29446
rect 14150 29246 14214 29310
rect 20814 29246 20878 29310
rect 21494 29382 21558 29446
rect 21766 29382 21830 29446
rect 21766 29246 21830 29310
rect 22038 29382 22102 29446
rect 22174 29246 22238 29310
rect 22446 29382 22510 29446
rect 22582 29246 22646 29310
rect 114246 29382 114310 29446
rect 114246 29246 114310 29310
rect 114654 29382 114718 29446
rect 114654 29246 114718 29310
rect 115334 29382 115398 29446
rect 115470 29382 115534 29446
rect 115062 29246 115126 29310
rect 115334 29246 115398 29310
rect 115878 29382 115942 29446
rect 116014 29246 116078 29310
rect 17822 29110 17886 29174
rect 1230 28974 1294 29038
rect 20814 28974 20878 29038
rect 20950 28838 21014 28902
rect 21222 28838 21286 28902
rect 21766 28974 21830 29038
rect 21630 28838 21694 28902
rect 22174 28974 22238 29038
rect 22038 28838 22102 28902
rect 22582 28974 22646 29038
rect 22582 28838 22646 28902
rect 114246 28974 114310 29038
rect 114382 28838 114446 28902
rect 114654 28974 114718 29038
rect 114790 28838 114854 28902
rect 115062 28974 115126 29038
rect 115334 28974 115398 29038
rect 115198 28838 115262 28902
rect 116014 28974 116078 29038
rect 115878 28838 115942 28902
rect 135326 28974 135390 29038
rect 20950 28566 21014 28630
rect 20950 28430 21014 28494
rect 21222 28566 21286 28630
rect 21630 28566 21694 28630
rect 21358 28430 21422 28494
rect 21494 28430 21558 28494
rect 22038 28566 22102 28630
rect 22174 28430 22238 28494
rect 22582 28566 22646 28630
rect 22446 28430 22510 28494
rect 114382 28566 114446 28630
rect 114382 28430 114446 28494
rect 114790 28566 114854 28630
rect 114790 28430 114854 28494
rect 115198 28566 115262 28630
rect 115606 28430 115670 28494
rect 115878 28566 115942 28630
rect 115878 28430 115942 28494
rect 20950 28158 21014 28222
rect 18910 28022 18974 28086
rect 21358 28158 21422 28222
rect 21494 28158 21558 28222
rect 21766 28022 21830 28086
rect 22174 28158 22238 28222
rect 22038 28022 22102 28086
rect 22446 28158 22510 28222
rect 22446 28022 22510 28086
rect 14014 27750 14078 27814
rect 15918 27614 15982 27678
rect 114382 28158 114446 28222
rect 114382 28022 114446 28086
rect 114790 28158 114854 28222
rect 114790 28022 114854 28086
rect 115198 28022 115262 28086
rect 115606 28158 115670 28222
rect 115878 28158 115942 28222
rect 1230 27206 1294 27270
rect 17414 27206 17478 27270
rect 17822 27478 17886 27542
rect 18366 27206 18430 27270
rect 18910 27342 18974 27406
rect 18638 27206 18702 27270
rect 19046 27206 19110 27270
rect 20678 27206 20742 27270
rect 21766 27750 21830 27814
rect 22038 27750 22102 27814
rect 22038 27614 22102 27678
rect 22446 27750 22510 27814
rect 22582 27614 22646 27678
rect 21358 27206 21422 27270
rect 21494 27206 21558 27270
rect 22038 27342 22102 27406
rect 20814 26934 20878 26998
rect 21358 26934 21422 26998
rect 21494 26934 21558 26998
rect 20678 26798 20742 26862
rect 22582 27342 22646 27406
rect 114382 27750 114446 27814
rect 114382 27614 114446 27678
rect 114790 27750 114854 27814
rect 114790 27614 114854 27678
rect 115198 27750 115262 27814
rect 17414 26662 17478 26726
rect 18366 26662 18430 26726
rect 18638 26662 18702 26726
rect 17550 26526 17614 26590
rect 17686 26526 17750 26590
rect 18230 26390 18294 26454
rect 18638 26390 18702 26454
rect 19046 26662 19110 26726
rect 20814 26662 20878 26726
rect 20814 26526 20878 26590
rect 21222 26526 21286 26590
rect 21902 26526 21966 26590
rect 27342 26662 27406 26726
rect 114382 27342 114446 27406
rect 114790 27342 114854 27406
rect 115606 27206 115670 27270
rect 115742 27206 115806 27270
rect 117646 27206 117710 27270
rect 117782 27206 117846 27270
rect 118190 27206 118254 27270
rect 118870 27206 118934 27270
rect 119278 27206 119342 27270
rect 135326 27206 135390 27270
rect 115606 26934 115670 26998
rect 115878 26934 115942 26998
rect 115742 26798 115806 26862
rect 117646 26798 117710 26862
rect 109350 26662 109414 26726
rect 27342 26390 27406 26454
rect 17686 26254 17750 26318
rect 20814 26254 20878 26318
rect 20814 26118 20878 26182
rect 21222 26254 21286 26318
rect 21902 26254 21966 26318
rect 22174 26118 22238 26182
rect 22582 26118 22646 26182
rect 27478 26254 27542 26318
rect 109350 26390 109414 26454
rect 109350 26254 109414 26318
rect 114246 26118 114310 26182
rect 115470 26526 115534 26590
rect 115878 26662 115942 26726
rect 115878 26526 115942 26590
rect 117782 26662 117846 26726
rect 117646 26390 117710 26454
rect 118190 26662 118254 26726
rect 118734 26662 118798 26726
rect 119006 26526 119070 26590
rect 119278 26662 119342 26726
rect 119278 26526 119342 26590
rect 118190 26390 118254 26454
rect 114654 26118 114718 26182
rect 27478 25982 27542 26046
rect 3814 25846 3878 25910
rect 17550 25846 17614 25910
rect 17414 25710 17478 25774
rect 18230 25846 18294 25910
rect 18638 25846 18702 25910
rect 18230 25710 18294 25774
rect 18774 25710 18838 25774
rect 19182 25710 19246 25774
rect 20814 25846 20878 25910
rect 20814 25710 20878 25774
rect 22174 25846 22238 25910
rect 22174 25710 22238 25774
rect 22582 25846 22646 25910
rect 109350 25982 109414 26046
rect 115470 26254 115534 26318
rect 115878 26254 115942 26318
rect 116014 26118 116078 26182
rect 22582 25710 22646 25774
rect 1230 25574 1294 25638
rect 20814 25438 20878 25502
rect 2537 25361 2601 25365
rect 2537 25305 2541 25361
rect 2541 25305 2597 25361
rect 2597 25305 2601 25361
rect 2537 25301 2601 25305
rect 20814 25302 20878 25366
rect 21358 25302 21422 25366
rect 21494 25302 21558 25366
rect 21766 25302 21830 25366
rect 22174 25438 22238 25502
rect 22174 25302 22238 25366
rect 22582 25438 22646 25502
rect 22446 25302 22510 25366
rect 114246 25846 114310 25910
rect 114246 25710 114310 25774
rect 114654 25846 114718 25910
rect 114790 25710 114854 25774
rect 115062 25710 115126 25774
rect 115606 25710 115670 25774
rect 116014 25846 116078 25910
rect 116014 25710 116078 25774
rect 117646 25846 117710 25910
rect 117646 25710 117710 25774
rect 118190 25846 118254 25910
rect 118190 25710 118254 25774
rect 119006 25846 119070 25910
rect 119006 25710 119070 25774
rect 119278 25846 119342 25910
rect 119414 25710 119478 25774
rect 120774 25710 120838 25774
rect 114246 25438 114310 25502
rect 114246 25302 114310 25366
rect 114790 25438 114854 25502
rect 114654 25302 114718 25366
rect 115062 25438 115126 25502
rect 115606 25438 115670 25502
rect 115198 25302 115262 25366
rect 115470 25302 115534 25366
rect 116014 25438 116078 25502
rect 135326 25438 135390 25502
rect 115878 25302 115942 25366
rect 15918 25030 15982 25094
rect 17414 25030 17478 25094
rect 18230 25030 18294 25094
rect 17686 24894 17750 24958
rect 18230 24894 18294 24958
rect 18774 25030 18838 25094
rect 19182 25030 19246 25094
rect 20814 25030 20878 25094
rect 20814 24894 20878 24958
rect 21358 25030 21422 25094
rect 21494 25030 21558 25094
rect 21766 25030 21830 25094
rect 21902 24894 21966 24958
rect 22174 25030 22238 25094
rect 22174 24894 22238 24958
rect 22446 25030 22510 25094
rect 22582 24894 22646 24958
rect 114246 25030 114310 25094
rect 114246 24894 114310 24958
rect 114654 25030 114718 25094
rect 114654 24894 114718 24958
rect 115198 25030 115262 25094
rect 115062 24894 115126 24958
rect 115470 25030 115534 25094
rect 115470 24894 115534 24958
rect 115878 25030 115942 25094
rect 116014 24894 116078 24958
rect 117646 25030 117710 25094
rect 117646 24894 117710 24958
rect 118190 25030 118254 25094
rect 118190 24894 118254 24958
rect 119006 25030 119070 25094
rect 119414 25030 119478 25094
rect 120774 25030 120838 25094
rect 2318 24486 2382 24550
rect 20814 24622 20878 24686
rect 20950 24486 21014 24550
rect 21902 24622 21966 24686
rect 21630 24486 21694 24550
rect 22174 24622 22238 24686
rect 22038 24486 22102 24550
rect 22582 24622 22646 24686
rect 22446 24486 22510 24550
rect 20950 24214 21014 24278
rect 21630 24214 21694 24278
rect 21222 24078 21286 24142
rect 21494 24078 21558 24142
rect 22038 24214 22102 24278
rect 22038 24078 22102 24142
rect 22446 24214 22510 24278
rect 22446 24078 22510 24142
rect 114246 24622 114310 24686
rect 114382 24486 114446 24550
rect 114654 24622 114718 24686
rect 114790 24486 114854 24550
rect 115062 24622 115126 24686
rect 115470 24622 115534 24686
rect 116014 24622 116078 24686
rect 115878 24486 115942 24550
rect 114382 24214 114446 24278
rect 1230 23942 1294 24006
rect 2318 23942 2382 24006
rect 27614 23942 27678 24006
rect 114246 24078 114310 24142
rect 114790 24214 114854 24278
rect 114790 24078 114854 24142
rect 115198 24078 115262 24142
rect 115606 24078 115670 24142
rect 115878 24214 115942 24278
rect 21222 23806 21286 23870
rect 21494 23806 21558 23870
rect 22038 23806 22102 23870
rect 22174 23670 22238 23734
rect 22446 23806 22510 23870
rect 22446 23670 22510 23734
rect 27478 23670 27542 23734
rect 27614 23670 27678 23734
rect 17686 23398 17750 23462
rect 18230 23398 18294 23462
rect 3814 23262 3878 23326
rect 550 23126 614 23190
rect 3814 23126 3878 23190
rect 18230 23262 18294 23326
rect 18638 23262 18702 23326
rect 19046 23262 19110 23326
rect 21358 23262 21422 23326
rect 21630 23262 21694 23326
rect 22174 23398 22238 23462
rect 22038 23262 22102 23326
rect 22446 23398 22510 23462
rect 114246 23806 114310 23870
rect 114246 23670 114310 23734
rect 114790 23806 114854 23870
rect 114790 23670 114854 23734
rect 115198 23806 115262 23870
rect 115606 23806 115670 23870
rect 135326 23806 135390 23870
rect 114246 23398 114310 23462
rect 22582 23262 22646 23326
rect 27478 23262 27542 23326
rect 27342 23126 27406 23190
rect 114382 23262 114446 23326
rect 114790 23398 114854 23462
rect 114790 23262 114854 23326
rect 117646 23398 117710 23462
rect 117646 23262 117710 23326
rect 118190 23398 118254 23462
rect 118054 23262 118118 23326
rect 118598 23262 118662 23326
rect 119006 23262 119070 23326
rect 109350 23126 109414 23190
rect 20950 22990 21014 23054
rect 21358 22990 21422 23054
rect 21494 22990 21558 23054
rect 21630 22990 21694 23054
rect 22038 22990 22102 23054
rect 18230 22718 18294 22782
rect 18366 22446 18430 22510
rect 18638 22718 18702 22782
rect 18638 22446 18702 22510
rect 19046 22718 19110 22782
rect 20950 22718 21014 22782
rect 20814 22582 20878 22646
rect 21494 22718 21558 22782
rect 21630 22582 21694 22646
rect 22582 22990 22646 23054
rect 27342 22854 27406 22918
rect 27478 22718 27542 22782
rect 109350 22854 109414 22918
rect 109486 22718 109550 22782
rect 114382 22990 114446 23054
rect 114790 22990 114854 23054
rect 116014 22990 116078 23054
rect 118326 22990 118390 23054
rect 118870 22990 118934 23054
rect 1230 22310 1294 22374
rect 20814 22310 20878 22374
rect 3134 22174 3198 22238
rect 20950 22174 21014 22238
rect 21630 22310 21694 22374
rect 20950 21902 21014 21966
rect 3134 21766 3198 21830
rect 20950 21766 21014 21830
rect 21358 21766 21422 21830
rect 21494 21766 21558 21830
rect 21766 21766 21830 21830
rect 22174 21766 22238 21830
rect 27478 22446 27542 22510
rect 27342 22310 27406 22374
rect 27342 22038 27406 22102
rect 109486 22446 109550 22510
rect 115062 22582 115126 22646
rect 116014 22718 116078 22782
rect 115878 22582 115942 22646
rect 117646 22718 117710 22782
rect 118054 22718 118118 22782
rect 118326 22718 118390 22782
rect 118598 22718 118662 22782
rect 118870 22718 118934 22782
rect 119006 22718 119070 22782
rect 118462 22446 118526 22510
rect 118870 22446 118934 22510
rect 109350 22310 109414 22374
rect 109350 22038 109414 22102
rect 115062 22310 115126 22374
rect 115878 22310 115942 22374
rect 115878 22174 115942 22238
rect 118326 22174 118390 22238
rect 118870 22174 118934 22238
rect 135326 22174 135390 22238
rect 22446 21766 22510 21830
rect 20950 21494 21014 21558
rect 20950 21358 21014 21422
rect 21358 21494 21422 21558
rect 21494 21494 21558 21558
rect 21766 21494 21830 21558
rect 21630 21358 21694 21422
rect 22174 21494 22238 21558
rect 22174 21358 22238 21422
rect 22446 21494 22510 21558
rect 22446 21358 22510 21422
rect 18366 21086 18430 21150
rect 17822 20950 17886 21014
rect 18638 21086 18702 21150
rect 18366 20950 18430 21014
rect 18638 20950 18702 21014
rect 19182 20950 19246 21014
rect 20950 21086 21014 21150
rect 20814 20950 20878 21014
rect 21358 20950 21422 21014
rect 21630 21086 21694 21150
rect 21766 20950 21830 21014
rect 22174 21086 22238 21150
rect 22038 20950 22102 21014
rect 22446 21086 22510 21150
rect 22446 20950 22510 21014
rect 114246 21766 114310 21830
rect 114654 21766 114718 21830
rect 115062 21766 115126 21830
rect 115606 21766 115670 21830
rect 115878 21902 115942 21966
rect 116014 21766 116078 21830
rect 109350 21494 109414 21558
rect 114246 21494 114310 21558
rect 114246 21358 114310 21422
rect 114654 21494 114718 21558
rect 114654 21358 114718 21422
rect 115062 21494 115126 21558
rect 115606 21494 115670 21558
rect 115606 21358 115670 21422
rect 116014 21494 116078 21558
rect 115878 21358 115942 21422
rect 118054 21358 118118 21422
rect 109350 21222 109414 21286
rect 118462 21222 118526 21286
rect 114246 21086 114310 21150
rect 114246 20950 114310 21014
rect 114654 21086 114718 21150
rect 114654 20950 114718 21014
rect 115606 21086 115670 21150
rect 115198 20950 115262 21014
rect 115334 20950 115398 21014
rect 115878 21086 115942 21150
rect 116014 20950 116078 21014
rect 118054 21086 118118 21150
rect 118326 21086 118390 21150
rect 117646 20950 117710 21014
rect 118190 20950 118254 21014
rect 118598 20950 118662 21014
rect 119006 20950 119070 21014
rect 20814 20678 20878 20742
rect 1230 20542 1294 20606
rect 20950 20542 21014 20606
rect 21358 20678 21422 20742
rect 21766 20678 21830 20742
rect 21358 20542 21422 20606
rect 21766 20542 21830 20606
rect 22038 20678 22102 20742
rect 22174 20542 22238 20606
rect 22446 20678 22510 20742
rect 22446 20542 22510 20606
rect 114246 20678 114310 20742
rect 114246 20542 114310 20606
rect 114654 20678 114718 20742
rect 114654 20542 114718 20606
rect 115198 20678 115262 20742
rect 115334 20678 115398 20742
rect 115062 20542 115126 20606
rect 115470 20542 115534 20606
rect 116014 20678 116078 20742
rect 116014 20542 116078 20606
rect 135326 20542 135390 20606
rect 3678 20406 3742 20470
rect 3814 20406 3878 20470
rect 17822 20270 17886 20334
rect 16598 20134 16662 20198
rect 17006 20134 17070 20198
rect 18366 20270 18430 20334
rect 18638 20270 18702 20334
rect 19182 20270 19246 20334
rect 20950 20270 21014 20334
rect 21358 20270 21422 20334
rect 21086 20134 21150 20198
rect 21766 20270 21830 20334
rect 22174 20270 22238 20334
rect 22446 20270 22510 20334
rect 22446 20134 22510 20198
rect 114246 20270 114310 20334
rect 114654 20270 114718 20334
rect 115062 20270 115126 20334
rect 115470 20270 115534 20334
rect 116014 20270 116078 20334
rect 117646 20270 117710 20334
rect 118190 20270 118254 20334
rect 118598 20270 118662 20334
rect 119006 20270 119070 20334
rect 119958 20134 120022 20198
rect 122814 20134 122878 20198
rect 109622 19998 109686 20062
rect 22446 19726 22510 19790
rect 28974 19726 29038 19790
rect 122814 19862 122878 19926
rect 109622 19726 109686 19790
rect 22446 19590 22510 19654
rect 26934 19590 26998 19654
rect 122814 19726 122878 19790
rect 26934 19318 26998 19382
rect 28294 19182 28358 19246
rect 28566 19182 28630 19246
rect 29518 19182 29582 19246
rect 30742 19182 30806 19246
rect 32510 19182 32574 19246
rect 33190 19182 33254 19246
rect 33734 19182 33798 19246
rect 34550 19182 34614 19246
rect 35638 19182 35702 19246
rect 37270 19182 37334 19246
rect 38222 19182 38286 19246
rect 38766 19182 38830 19246
rect 39446 19182 39510 19246
rect 39990 19182 40054 19246
rect 40670 19182 40734 19246
rect 41214 19182 41278 19246
rect 42030 19182 42094 19246
rect 42438 19182 42502 19246
rect 43254 19182 43318 19246
rect 43390 19182 43454 19246
rect 44478 19182 44542 19246
rect 45702 19182 45766 19246
rect 46926 19182 46990 19246
rect 47470 19182 47534 19246
rect 48150 19182 48214 19246
rect 49918 19182 49982 19246
rect 51278 19182 51342 19246
rect 51958 19182 52022 19246
rect 53182 19182 53246 19246
rect 53726 19182 53790 19246
rect 54406 19182 54470 19246
rect 54950 19182 55014 19246
rect 55630 19182 55694 19246
rect 56174 19182 56238 19246
rect 57398 19182 57462 19246
rect 58214 19182 58278 19246
rect 59438 19182 59502 19246
rect 59982 19182 60046 19246
rect 60662 19182 60726 19246
rect 60798 19182 60862 19246
rect 61886 19182 61950 19246
rect 62430 19182 62494 19246
rect 63110 19182 63174 19246
rect 64470 19182 64534 19246
rect 66238 19182 66302 19246
rect 66918 19182 66982 19246
rect 67462 19182 67526 19246
rect 68686 19182 68750 19246
rect 69366 19182 69430 19246
rect 70998 19182 71062 19246
rect 71950 19182 72014 19246
rect 72358 19182 72422 19246
rect 73174 19182 73238 19246
rect 74942 19182 75006 19246
rect 75622 19182 75686 19246
rect 76166 19182 76230 19246
rect 77390 19182 77454 19246
rect 78070 19182 78134 19246
rect 79702 19182 79766 19246
rect 80654 19182 80718 19246
rect 81198 19182 81262 19246
rect 81878 19182 81942 19246
rect 83646 19182 83710 19246
rect 84326 19182 84390 19246
rect 84870 19182 84934 19246
rect 86094 19182 86158 19246
rect 86910 19182 86974 19246
rect 87318 19182 87382 19246
rect 88134 19182 88198 19246
rect 88270 19182 88334 19246
rect 89358 19182 89422 19246
rect 89902 19182 89966 19246
rect 90718 19182 90782 19246
rect 91806 19182 91870 19246
rect 94526 19318 94590 19382
rect 92350 19182 92414 19246
rect 93438 19182 93502 19246
rect 95614 19182 95678 19246
rect 96158 19182 96222 19246
rect 96838 19182 96902 19246
rect 98198 19182 98262 19246
rect 98606 19182 98670 19246
rect 99830 19182 99894 19246
rect 101190 19182 101254 19246
rect 101870 19182 101934 19246
rect 102414 19182 102478 19246
rect 103094 19182 103158 19246
rect 104318 19182 104382 19246
rect 104862 19182 104926 19246
rect 105542 19182 105606 19246
rect 105814 19182 105878 19246
rect 107174 19182 107238 19246
rect 107310 19182 107374 19246
rect 108534 19182 108598 19246
rect 1230 18774 1294 18838
rect 16598 19046 16662 19110
rect 135326 18910 135390 18974
rect 14694 18774 14758 18838
rect 28294 18774 28358 18838
rect 28566 18774 28630 18838
rect 29518 18774 29582 18838
rect 30742 18774 30806 18838
rect 32510 18774 32574 18838
rect 33190 18774 33254 18838
rect 33734 18774 33798 18838
rect 34550 18774 34614 18838
rect 35638 18774 35702 18838
rect 37270 18774 37334 18838
rect 38222 18774 38286 18838
rect 38766 18774 38830 18838
rect 39446 18774 39510 18838
rect 39990 18774 40054 18838
rect 40670 18774 40734 18838
rect 41214 18774 41278 18838
rect 42030 18774 42094 18838
rect 42438 18774 42502 18838
rect 43254 18774 43318 18838
rect 43390 18774 43454 18838
rect 44478 18774 44542 18838
rect 45702 18774 45766 18838
rect 46926 18774 46990 18838
rect 47470 18774 47534 18838
rect 48150 18774 48214 18838
rect 49918 18774 49982 18838
rect 51278 18774 51342 18838
rect 51958 18774 52022 18838
rect 53182 18774 53246 18838
rect 53726 18774 53790 18838
rect 54406 18774 54470 18838
rect 54950 18774 55014 18838
rect 55630 18774 55694 18838
rect 56174 18774 56238 18838
rect 57398 18774 57462 18838
rect 58214 18774 58278 18838
rect 58350 18638 58414 18702
rect 59438 18774 59502 18838
rect 59982 18774 60046 18838
rect 60662 18774 60726 18838
rect 60798 18774 60862 18838
rect 61886 18774 61950 18838
rect 62430 18774 62494 18838
rect 63110 18774 63174 18838
rect 64470 18774 64534 18838
rect 66238 18774 66302 18838
rect 66918 18774 66982 18838
rect 67462 18774 67526 18838
rect 68686 18774 68750 18838
rect 69366 18774 69430 18838
rect 70998 18774 71062 18838
rect 71950 18774 72014 18838
rect 72358 18774 72422 18838
rect 73174 18774 73238 18838
rect 74942 18774 75006 18838
rect 75622 18774 75686 18838
rect 76166 18774 76230 18838
rect 77390 18774 77454 18838
rect 78070 18774 78134 18838
rect 79702 18774 79766 18838
rect 80654 18774 80718 18838
rect 81198 18774 81262 18838
rect 81878 18774 81942 18838
rect 83646 18774 83710 18838
rect 84326 18774 84390 18838
rect 84870 18774 84934 18838
rect 86094 18774 86158 18838
rect 86910 18774 86974 18838
rect 87318 18774 87382 18838
rect 88134 18774 88198 18838
rect 88270 18774 88334 18838
rect 89358 18774 89422 18838
rect 89902 18774 89966 18838
rect 90718 18774 90782 18838
rect 91806 18774 91870 18838
rect 92350 18774 92414 18838
rect 93438 18774 93502 18838
rect 94526 18774 94590 18838
rect 95614 18774 95678 18838
rect 96158 18774 96222 18838
rect 96838 18774 96902 18838
rect 98198 18774 98262 18838
rect 98606 18774 98670 18838
rect 99830 18774 99894 18838
rect 101190 18774 101254 18838
rect 101870 18774 101934 18838
rect 102414 18774 102478 18838
rect 103094 18774 103158 18838
rect 104318 18774 104382 18838
rect 104862 18774 104926 18838
rect 105542 18774 105606 18838
rect 105814 18774 105878 18838
rect 107174 18774 107238 18838
rect 107310 18774 107374 18838
rect 108534 18774 108598 18838
rect 119958 18502 120022 18566
rect 122950 18366 123014 18430
rect 2537 17894 2601 17958
rect 3678 17550 3742 17614
rect 17006 17550 17070 17614
rect 14558 17414 14622 17478
rect 21222 17278 21286 17342
rect 21358 17142 21422 17206
rect 28974 17142 29038 17206
rect 1230 17006 1294 17070
rect 28974 17006 29038 17070
rect 31694 17006 31758 17070
rect 34006 17006 34070 17070
rect 36454 17006 36518 17070
rect 39174 17006 39238 17070
rect 41622 17006 41686 17070
rect 44070 17006 44134 17070
rect 46654 17006 46718 17070
rect 48966 17006 49030 17070
rect 51550 17006 51614 17070
rect 54134 17006 54198 17070
rect 56446 17006 56510 17070
rect 59166 17006 59230 17070
rect 61614 17006 61678 17070
rect 63926 17006 63990 17070
rect 66646 17006 66710 17070
rect 69094 17006 69158 17070
rect 71406 17006 71470 17070
rect 74126 17006 74190 17070
rect 76438 17006 76502 17070
rect 78886 17006 78950 17070
rect 81606 17006 81670 17070
rect 83918 17006 83982 17070
rect 86366 17006 86430 17070
rect 89086 17006 89150 17070
rect 91398 17006 91462 17070
rect 93982 17006 94046 17070
rect 96566 17006 96630 17070
rect 98878 17006 98942 17070
rect 101598 17006 101662 17070
rect 104046 17006 104110 17070
rect 106358 17006 106422 17070
rect 135326 17142 135390 17206
rect 122814 17006 122878 17070
rect 122814 16870 122878 16934
rect 3134 16054 3198 16118
rect 14694 16190 14758 16254
rect 14694 16054 14758 16118
rect 21222 15782 21286 15846
rect 22446 15782 22510 15846
rect 122950 15646 123014 15710
rect 1230 15510 1294 15574
rect 3134 15510 3198 15574
rect 122950 15510 123014 15574
rect 135326 15374 135390 15438
rect 28974 15102 29038 15166
rect 29110 15102 29174 15166
rect 31558 15102 31622 15166
rect 31694 15102 31758 15166
rect 34006 15102 34070 15166
rect 34142 15102 34206 15166
rect 36454 15102 36518 15166
rect 36590 15102 36654 15166
rect 39038 15102 39102 15166
rect 39174 15102 39238 15166
rect 41486 15102 41550 15166
rect 41622 15102 41686 15166
rect 43934 15102 43998 15166
rect 44070 15102 44134 15166
rect 46518 15102 46582 15166
rect 46654 15102 46718 15166
rect 48966 15102 49030 15166
rect 49102 15102 49166 15166
rect 51414 15102 51478 15166
rect 51550 15102 51614 15166
rect 53998 15102 54062 15166
rect 54134 15102 54198 15166
rect 56446 15102 56510 15166
rect 56582 15102 56646 15166
rect 59030 15102 59094 15166
rect 59166 15102 59230 15166
rect 61478 15102 61542 15166
rect 61614 15102 61678 15166
rect 63926 15102 63990 15166
rect 64062 15102 64126 15166
rect 66510 15102 66574 15166
rect 66646 15102 66710 15166
rect 68958 15102 69022 15166
rect 69094 15102 69158 15166
rect 71406 15102 71470 15166
rect 71542 15102 71606 15166
rect 73990 15102 74054 15166
rect 74126 15102 74190 15166
rect 76438 15102 76502 15166
rect 76574 15102 76638 15166
rect 78886 15102 78950 15166
rect 79022 15102 79086 15166
rect 81470 15102 81534 15166
rect 81606 15102 81670 15166
rect 83918 15102 83982 15166
rect 84054 15102 84118 15166
rect 86366 15102 86430 15166
rect 86502 15102 86566 15166
rect 88950 15102 89014 15166
rect 89086 15102 89150 15166
rect 91398 15102 91462 15166
rect 91534 15102 91598 15166
rect 93846 15102 93910 15166
rect 93982 15102 94046 15166
rect 96430 15102 96494 15166
rect 96566 15102 96630 15166
rect 98878 15102 98942 15166
rect 99014 15102 99078 15166
rect 101462 15102 101526 15166
rect 101598 15102 101662 15166
rect 103910 15102 103974 15166
rect 104046 15102 104110 15166
rect 106358 15102 106422 15166
rect 106494 15102 106558 15166
rect 550 14694 614 14758
rect 14558 14694 14622 14758
rect 14558 14558 14622 14622
rect 21358 14558 21422 14622
rect 20270 14286 20334 14350
rect 28838 14286 28902 14350
rect 31422 14286 31486 14350
rect 33598 14286 33662 14350
rect 33870 14286 33934 14350
rect 36454 14286 36518 14350
rect 38902 14286 38966 14350
rect 41078 14286 41142 14350
rect 41214 14286 41278 14350
rect 43798 14286 43862 14350
rect 46246 14286 46310 14350
rect 48830 14286 48894 14350
rect 51414 14286 51478 14350
rect 58350 14422 58414 14486
rect 53862 14286 53926 14350
rect 56446 14286 56510 14350
rect 58622 14286 58686 14350
rect 58894 14286 58958 14350
rect 61070 14286 61134 14350
rect 61342 14286 61406 14350
rect 63654 14286 63718 14350
rect 63790 14286 63854 14350
rect 66238 14286 66302 14350
rect 68822 14286 68886 14350
rect 71270 14286 71334 14350
rect 73854 14286 73918 14350
rect 76030 14286 76094 14350
rect 76302 14286 76366 14350
rect 78886 14286 78950 14350
rect 81334 14286 81398 14350
rect 83646 14286 83710 14350
rect 86094 14286 86158 14350
rect 86230 14286 86294 14350
rect 88678 14286 88742 14350
rect 91262 14286 91326 14350
rect 93846 14286 93910 14350
rect 96294 14286 96358 14350
rect 98878 14286 98942 14350
rect 101326 14286 101390 14350
rect 103502 14286 103566 14350
rect 103774 14286 103838 14350
rect 106358 14286 106422 14350
rect 122814 14286 122878 14350
rect 122814 14014 122878 14078
rect 1230 13878 1294 13942
rect 135326 13878 135390 13942
rect 3134 13742 3198 13806
rect 28838 13606 28902 13670
rect 28974 13470 29038 13534
rect 31422 13606 31486 13670
rect 33598 13606 33662 13670
rect 33870 13606 33934 13670
rect 36454 13606 36518 13670
rect 38902 13606 38966 13670
rect 41078 13606 41142 13670
rect 41214 13606 41278 13670
rect 43798 13606 43862 13670
rect 46246 13606 46310 13670
rect 48830 13606 48894 13670
rect 51414 13606 51478 13670
rect 53862 13606 53926 13670
rect 31286 13470 31350 13534
rect 34006 13470 34070 13534
rect 36454 13470 36518 13534
rect 38902 13470 38966 13534
rect 41350 13470 41414 13534
rect 43934 13470 43998 13534
rect 46382 13470 46446 13534
rect 48966 13470 49030 13534
rect 51414 13470 51478 13534
rect 53862 13470 53926 13534
rect 56446 13606 56510 13670
rect 58622 13606 58686 13670
rect 58894 13606 58958 13670
rect 61070 13606 61134 13670
rect 61206 13606 61270 13670
rect 61342 13606 61406 13670
rect 63654 13606 63718 13670
rect 63790 13606 63854 13670
rect 66238 13606 66302 13670
rect 68686 13606 68750 13670
rect 68822 13606 68886 13670
rect 71270 13606 71334 13670
rect 73854 13606 73918 13670
rect 76030 13606 76094 13670
rect 76302 13606 76366 13670
rect 78886 13606 78950 13670
rect 81334 13606 81398 13670
rect 83646 13606 83710 13670
rect 86094 13606 86158 13670
rect 86230 13606 86294 13670
rect 88678 13606 88742 13670
rect 91262 13606 91326 13670
rect 93846 13606 93910 13670
rect 96294 13606 96358 13670
rect 98878 13606 98942 13670
rect 101326 13606 101390 13670
rect 103502 13606 103566 13670
rect 103638 13606 103702 13670
rect 103774 13606 103838 13670
rect 106358 13606 106422 13670
rect 56310 13470 56374 13534
rect 58894 13470 58958 13534
rect 63926 13470 63990 13534
rect 66374 13470 66438 13534
rect 71406 13470 71470 13534
rect 73854 13470 73918 13534
rect 76438 13470 76502 13534
rect 78886 13470 78950 13534
rect 81334 13470 81398 13534
rect 83918 13470 83982 13534
rect 86366 13470 86430 13534
rect 88814 13470 88878 13534
rect 91398 13470 91462 13534
rect 93846 13470 93910 13534
rect 96294 13470 96358 13534
rect 98878 13470 98942 13534
rect 101326 13470 101390 13534
rect 106358 13470 106422 13534
rect 3134 13334 3198 13398
rect 14694 13334 14758 13398
rect 14694 13198 14758 13262
rect 29110 13198 29174 13262
rect 21222 13062 21286 13126
rect 28294 13062 28358 13126
rect 29110 13062 29174 13126
rect 30742 13062 30806 13126
rect 31558 13198 31622 13262
rect 31422 13062 31486 13126
rect 34142 13198 34206 13262
rect 33598 13062 33662 13126
rect 33870 13062 33934 13126
rect 36590 13198 36654 13262
rect 36046 13062 36110 13126
rect 39038 13198 39102 13262
rect 36590 13062 36654 13126
rect 38494 13062 38558 13126
rect 41486 13198 41550 13262
rect 39038 13062 39102 13126
rect 41078 13062 41142 13126
rect 41486 13062 41550 13126
rect 44070 13198 44134 13262
rect 43526 13062 43590 13126
rect 46518 13198 46582 13262
rect 44070 13062 44134 13126
rect 45974 13062 46038 13126
rect 49102 13198 49166 13262
rect 46518 13062 46582 13126
rect 48286 13062 48350 13126
rect 48830 13062 48894 13126
rect 51550 13198 51614 13262
rect 51006 13062 51070 13126
rect 53998 13198 54062 13262
rect 51550 13062 51614 13126
rect 53590 13062 53654 13126
rect 53998 13062 54062 13126
rect 56038 13062 56102 13126
rect 56582 13198 56646 13262
rect 56446 13062 56510 13126
rect 59030 13198 59094 13262
rect 58486 13062 58550 13126
rect 59030 13062 59094 13126
rect 60934 13062 60998 13126
rect 61342 13062 61406 13126
rect 61478 13062 61542 13126
rect 64062 13198 64126 13262
rect 63518 13062 63582 13126
rect 66510 13198 66574 13262
rect 64062 13062 64126 13126
rect 65966 13062 66030 13126
rect 66510 13062 66574 13126
rect 68278 13062 68342 13126
rect 68822 13062 68886 13126
rect 68958 13062 69022 13126
rect 71542 13198 71606 13262
rect 70998 13062 71062 13126
rect 73990 13198 74054 13262
rect 71542 13062 71606 13126
rect 73446 13062 73510 13126
rect 76574 13198 76638 13262
rect 73990 13062 74054 13126
rect 75894 13062 75958 13126
rect 76302 13062 76366 13126
rect 79022 13198 79086 13262
rect 78478 13062 78542 13126
rect 81470 13198 81534 13262
rect 79022 13062 79086 13126
rect 80926 13062 80990 13126
rect 84054 13198 84118 13262
rect 81470 13062 81534 13126
rect 83510 13062 83574 13126
rect 83782 13062 83846 13126
rect 86502 13198 86566 13262
rect 85958 13062 86022 13126
rect 88950 13198 89014 13262
rect 86502 13062 86566 13126
rect 88542 13062 88606 13126
rect 91534 13198 91598 13262
rect 88950 13062 89014 13126
rect 90990 13062 91054 13126
rect 91262 13062 91326 13126
rect 93982 13198 94046 13262
rect 93438 13062 93502 13126
rect 96430 13198 96494 13262
rect 93982 13062 94046 13126
rect 95886 13062 95950 13126
rect 99014 13198 99078 13262
rect 96430 13062 96494 13126
rect 98470 13062 98534 13126
rect 101462 13198 101526 13262
rect 99014 13062 99078 13126
rect 100918 13062 100982 13126
rect 101462 13062 101526 13126
rect 103366 13062 103430 13126
rect 103774 13062 103838 13126
rect 103910 13062 103974 13126
rect 106494 13198 106558 13262
rect 105950 13062 106014 13126
rect 106494 13062 106558 13126
rect 122950 12790 123014 12854
rect 122950 12654 123014 12718
rect 29110 12518 29174 12582
rect 31422 12518 31486 12582
rect 33870 12518 33934 12582
rect 1230 12246 1294 12310
rect 28838 12246 28902 12310
rect 31422 12246 31486 12310
rect 33462 12246 33526 12310
rect 36590 12518 36654 12582
rect 39038 12518 39102 12582
rect 41486 12518 41550 12582
rect 44070 12518 44134 12582
rect 46518 12518 46582 12582
rect 48830 12518 48894 12582
rect 36182 12246 36246 12310
rect 38630 12246 38694 12310
rect 41486 12246 41550 12310
rect 43390 12246 43454 12310
rect 46518 12246 46582 12310
rect 48830 12246 48894 12310
rect 51550 12518 51614 12582
rect 53998 12518 54062 12582
rect 56446 12518 56510 12582
rect 59030 12518 59094 12582
rect 61342 12518 61406 12582
rect 51278 12246 51342 12310
rect 53998 12246 54062 12310
rect 56446 12246 56510 12310
rect 59030 12246 59094 12310
rect 61342 12246 61406 12310
rect 64062 12518 64126 12582
rect 66510 12518 66574 12582
rect 68822 12518 68886 12582
rect 63654 12246 63718 12310
rect 66238 12246 66302 12310
rect 68550 12246 68614 12310
rect 71542 12518 71606 12582
rect 73990 12518 74054 12582
rect 76302 12518 76366 12582
rect 71542 12246 71606 12310
rect 73310 12246 73374 12310
rect 76166 12246 76230 12310
rect 79022 12518 79086 12582
rect 81470 12518 81534 12582
rect 83782 12518 83846 12582
rect 78614 12246 78678 12310
rect 81062 12246 81126 12310
rect 86502 12518 86566 12582
rect 88950 12518 89014 12582
rect 91262 12518 91326 12582
rect 84054 12246 84118 12310
rect 86502 12246 86566 12310
rect 88950 12246 89014 12310
rect 91262 12246 91326 12310
rect 93982 12518 94046 12582
rect 96430 12518 96494 12582
rect 99014 12518 99078 12582
rect 101462 12518 101526 12582
rect 103774 12518 103838 12582
rect 93710 12246 93774 12310
rect 96022 12246 96086 12310
rect 99014 12246 99078 12310
rect 101462 12246 101526 12310
rect 103774 12246 103838 12310
rect 106494 12518 106558 12582
rect 106086 12246 106150 12310
rect 135326 12246 135390 12310
rect 14558 11974 14622 12038
rect 28974 11974 29038 12038
rect 31286 11974 31350 12038
rect 28702 11838 28766 11902
rect 31150 11838 31214 11902
rect 34006 11974 34070 12038
rect 36454 11974 36518 12038
rect 38902 11974 38966 12038
rect 41350 11974 41414 12038
rect 43934 11974 43998 12038
rect 46382 11974 46446 12038
rect 48966 11974 49030 12038
rect 51414 11974 51478 12038
rect 53862 11974 53926 12038
rect 56310 11974 56374 12038
rect 33870 11838 33934 11902
rect 36318 11838 36382 11902
rect 38766 11838 38830 11902
rect 41350 11838 41414 11902
rect 43798 11838 43862 11902
rect 46246 11838 46310 11902
rect 48694 11838 48758 11902
rect 51142 11838 51206 11902
rect 53862 11838 53926 11902
rect 56310 11838 56374 11902
rect 58894 11974 58958 12038
rect 61206 11974 61270 12038
rect 58758 11838 58822 11902
rect 61206 11838 61270 11902
rect 63926 11974 63990 12038
rect 66374 11974 66438 12038
rect 68686 11974 68750 12038
rect 63790 11838 63854 11902
rect 66102 11838 66166 11902
rect 68822 11838 68886 11902
rect 71406 11974 71470 12038
rect 73854 11974 73918 12038
rect 76438 11974 76502 12038
rect 78886 11974 78950 12038
rect 81334 11974 81398 12038
rect 83918 11974 83982 12038
rect 86366 11974 86430 12038
rect 88814 11974 88878 12038
rect 91398 11974 91462 12038
rect 93846 11974 93910 12038
rect 96294 11974 96358 12038
rect 98878 11974 98942 12038
rect 101326 11974 101390 12038
rect 103638 11974 103702 12038
rect 71270 11838 71334 11902
rect 73718 11838 73782 11902
rect 76302 11838 76366 11902
rect 78750 11838 78814 11902
rect 81198 11838 81262 11902
rect 83782 11838 83846 11902
rect 86230 11838 86294 11902
rect 88814 11838 88878 11902
rect 91126 11838 91190 11902
rect 93574 11838 93638 11902
rect 96158 11838 96222 11902
rect 98742 11838 98806 11902
rect 101190 11838 101254 11902
rect 103638 11838 103702 11902
rect 106358 11974 106422 12038
rect 106222 11838 106286 11902
rect 123222 11898 123270 11902
rect 123270 11898 123286 11902
rect 123222 11838 123286 11898
rect 14558 11702 14622 11766
rect 20270 11702 20334 11766
rect 28838 11702 28902 11766
rect 31422 11702 31486 11766
rect 33462 11702 33526 11766
rect 36182 11702 36246 11766
rect 38630 11702 38694 11766
rect 41486 11702 41550 11766
rect 46518 11702 46582 11766
rect 48830 11702 48894 11766
rect 51278 11702 51342 11766
rect 53998 11702 54062 11766
rect 56446 11702 56510 11766
rect 59030 11702 59094 11766
rect 61342 11702 61406 11766
rect 63654 11702 63718 11766
rect 66238 11702 66302 11766
rect 68550 11702 68614 11766
rect 71542 11702 71606 11766
rect 76166 11702 76230 11766
rect 78614 11702 78678 11766
rect 81062 11702 81126 11766
rect 84054 11702 84118 11766
rect 86502 11702 86566 11766
rect 88950 11702 89014 11766
rect 91262 11702 91326 11766
rect 96022 11702 96086 11766
rect 99014 11702 99078 11766
rect 101462 11702 101526 11766
rect 103774 11702 103838 11766
rect 106086 11702 106150 11766
rect 28158 11294 28222 11358
rect 43390 11430 43454 11494
rect 73310 11430 73374 11494
rect 93710 11430 93774 11494
rect 122814 11430 122878 11494
rect 108398 11294 108462 11358
rect 28566 11022 28630 11086
rect 28702 11022 28766 11086
rect 31150 11022 31214 11086
rect 33870 11022 33934 11086
rect 36318 11022 36382 11086
rect 38766 11022 38830 11086
rect 41350 11022 41414 11086
rect 43798 11022 43862 11086
rect 46246 11022 46310 11086
rect 48694 11022 48758 11086
rect 51142 11022 51206 11086
rect 53862 11022 53926 11086
rect 56310 11022 56374 11086
rect 58758 11022 58822 11086
rect 61206 11022 61270 11086
rect 63790 11022 63854 11086
rect 66102 11022 66166 11086
rect 68822 11022 68886 11086
rect 71270 11022 71334 11086
rect 73718 11022 73782 11086
rect 76302 11022 76366 11086
rect 78750 11022 78814 11086
rect 81198 11022 81262 11086
rect 83782 11022 83846 11086
rect 86230 11022 86294 11086
rect 88814 11022 88878 11086
rect 91126 11022 91190 11086
rect 93574 11022 93638 11086
rect 96158 11022 96222 11086
rect 98742 11022 98806 11086
rect 101190 11022 101254 11086
rect 103638 11022 103702 11086
rect 106222 11022 106286 11086
rect 108262 11022 108326 11086
rect 123358 10750 123422 10814
rect 28566 10614 28630 10678
rect 108262 10614 108326 10678
rect 1230 10478 1294 10542
rect 14694 10478 14758 10542
rect 14694 10342 14758 10406
rect 135326 10342 135390 10406
rect 550 10206 614 10270
rect 122950 9934 123014 9998
rect 28158 9526 28222 9590
rect 108398 9526 108462 9590
rect 14558 9118 14622 9182
rect 16326 8982 16390 9046
rect 1230 8710 1294 8774
rect 135326 8710 135390 8774
rect 550 7622 614 7686
rect 14694 7622 14758 7686
rect 1230 7214 1294 7278
rect 135326 7078 135390 7142
rect 1230 5446 1294 5510
rect 135326 5310 135390 5374
rect 1230 3814 1294 3878
rect 16326 3814 16390 3878
rect 20270 3678 20334 3742
rect 135326 3678 135390 3742
rect 16054 2862 16118 2926
rect 17142 2862 17206 2926
rect 18230 2862 18294 2926
rect 19590 2862 19654 2926
rect 20542 2862 20606 2926
rect 21766 2862 21830 2926
rect 23126 2862 23190 2926
rect 24214 2862 24278 2926
rect 25438 2862 25502 2926
rect 26526 2862 26590 2926
rect 27614 2862 27678 2926
rect 28702 2862 28766 2926
rect 30062 2862 30126 2926
rect 31286 2862 31350 2926
rect 32374 2862 32438 2926
rect 33462 2862 33526 2926
rect 34550 2862 34614 2926
rect 35910 2862 35974 2926
rect 36998 2862 37062 2926
rect 38086 2862 38150 2926
rect 39446 2862 39510 2926
rect 40670 2862 40734 2926
rect 41758 2862 41822 2926
rect 42846 2862 42910 2926
rect 43934 2862 43998 2926
rect 45294 2862 45358 2926
rect 46382 2862 46446 2926
rect 47606 2862 47670 2926
rect 48694 2862 48758 2926
rect 49782 2862 49846 2926
rect 51142 2862 51206 2926
rect 52230 2862 52294 2926
rect 53318 2862 53382 2926
rect 54406 2862 54470 2926
rect 55766 2862 55830 2926
rect 56990 2862 57054 2926
rect 58078 2862 58142 2926
rect 59166 2862 59230 2926
rect 39718 2318 39782 2382
rect 135326 2046 135390 2110
rect 2046 1638 2110 1702
rect 3814 1696 3866 1702
rect 3866 1696 3878 1702
rect 3814 1638 3878 1696
rect 5582 1638 5646 1702
rect 7078 1638 7142 1702
rect 8710 1638 8774 1702
rect 10478 1696 10530 1702
rect 10530 1696 10542 1702
rect 10478 1638 10542 1696
rect 12110 1638 12174 1702
rect 14014 1638 14078 1702
rect 15510 1696 15570 1702
rect 15570 1696 15574 1702
rect 15510 1638 15574 1696
rect 20270 1774 20334 1838
rect 17414 1638 17478 1702
rect 19046 1638 19110 1702
rect 20814 1638 20878 1702
rect 22174 1638 22238 1702
rect 23942 1696 23970 1702
rect 23970 1696 24006 1702
rect 23942 1638 24006 1696
rect 25710 1638 25774 1702
rect 27342 1696 27386 1702
rect 27386 1696 27406 1702
rect 27342 1638 27406 1696
rect 28974 1696 29010 1702
rect 29010 1696 29038 1702
rect 28974 1638 29038 1696
rect 30470 1638 30534 1702
rect 32102 1638 32166 1702
rect 34006 1696 34050 1702
rect 34050 1696 34070 1702
rect 34006 1638 34070 1696
rect 35774 1696 35786 1702
rect 35786 1696 35838 1702
rect 35774 1638 35838 1696
rect 37406 1696 37410 1702
rect 37410 1696 37466 1702
rect 37466 1696 37470 1702
rect 37406 1638 37470 1696
rect 39174 1638 39238 1702
rect 40806 1696 40826 1702
rect 40826 1696 40870 1702
rect 40806 1638 40870 1696
rect 42438 1696 42450 1702
rect 42450 1696 42502 1702
rect 42438 1638 42502 1696
rect 44206 1638 44270 1702
rect 45702 1638 45766 1702
rect 47334 1638 47398 1702
rect 49102 1638 49166 1702
rect 50734 1638 50798 1702
rect 52502 1696 52530 1702
rect 52530 1696 52566 1702
rect 52502 1638 52566 1696
rect 54134 1638 54198 1702
rect 55494 1638 55558 1702
rect 57534 1696 57570 1702
rect 57570 1696 57598 1702
rect 57534 1638 57598 1696
rect 59438 1638 59502 1702
rect 60798 1638 60862 1702
rect 62566 1696 62610 1702
rect 62610 1696 62630 1702
rect 62566 1638 62630 1696
rect 64334 1696 64346 1702
rect 64346 1696 64398 1702
rect 64334 1638 64398 1696
rect 65830 1638 65894 1702
rect 67598 1696 67650 1702
rect 67650 1696 67662 1702
rect 67598 1638 67662 1696
rect 69230 1638 69294 1702
rect 70862 1638 70926 1702
rect 72766 1638 72830 1702
rect 74262 1638 74326 1702
rect 76166 1638 76230 1702
rect 77662 1638 77726 1702
rect 79294 1638 79358 1702
rect 81062 1696 81090 1702
rect 81090 1696 81126 1702
rect 81062 1638 81126 1696
rect 82830 1638 82894 1702
rect 84326 1638 84390 1702
rect 86230 1638 86294 1702
rect 87726 1638 87790 1702
rect 89358 1638 89422 1702
rect 91262 1638 91326 1702
rect 92758 1638 92822 1702
rect 94390 1638 94454 1702
rect 96158 1696 96210 1702
rect 96210 1696 96222 1702
rect 96158 1638 96222 1696
rect 97790 1638 97854 1702
rect 99558 1696 99570 1702
rect 99570 1696 99622 1702
rect 99558 1638 99622 1696
rect 101326 1638 101390 1702
rect 102822 1638 102886 1702
rect 104590 1696 104610 1702
rect 104610 1696 104654 1702
rect 104590 1638 104654 1696
rect 106222 1638 106286 1702
rect 107854 1638 107918 1702
rect 109758 1638 109822 1702
rect 111254 1638 111318 1702
rect 113022 1696 113066 1702
rect 113066 1696 113086 1702
rect 113022 1638 113086 1696
rect 114790 1638 114854 1702
rect 116286 1638 116350 1702
rect 118054 1696 118106 1702
rect 118106 1696 118118 1702
rect 118054 1638 118118 1696
rect 119822 1638 119886 1702
rect 121318 1638 121382 1702
rect 123086 1696 123090 1702
rect 123090 1696 123146 1702
rect 123146 1696 123150 1702
rect 123086 1638 123150 1696
rect 124718 1696 124770 1702
rect 124770 1696 124782 1702
rect 124718 1638 124782 1696
rect 126350 1638 126414 1702
rect 127982 1638 128046 1702
rect 129750 1696 129810 1702
rect 129810 1696 129814 1702
rect 129750 1638 129814 1696
rect 131518 1696 131546 1702
rect 131546 1696 131582 1702
rect 131518 1638 131582 1696
rect 133150 1696 133170 1702
rect 133170 1696 133214 1702
rect 133150 1638 133214 1696
rect 958 1230 1022 1294
rect 1094 1230 1158 1294
rect 1230 1230 1294 1294
rect 2046 1230 2110 1294
rect 3814 1230 3878 1294
rect 5582 1230 5646 1294
rect 7078 1230 7142 1294
rect 8710 1230 8774 1294
rect 10478 1230 10542 1294
rect 12110 1230 12174 1294
rect 14014 1230 14078 1294
rect 15510 1230 15574 1294
rect 17414 1230 17478 1294
rect 19046 1230 19110 1294
rect 20814 1230 20878 1294
rect 22174 1230 22238 1294
rect 23942 1230 24006 1294
rect 25710 1230 25774 1294
rect 27342 1230 27406 1294
rect 28974 1230 29038 1294
rect 30470 1230 30534 1294
rect 32102 1230 32166 1294
rect 34006 1230 34070 1294
rect 35774 1230 35838 1294
rect 37406 1230 37470 1294
rect 39174 1230 39238 1294
rect 40806 1230 40870 1294
rect 42438 1230 42502 1294
rect 44206 1230 44270 1294
rect 45702 1230 45766 1294
rect 47334 1230 47398 1294
rect 49102 1230 49166 1294
rect 50734 1230 50798 1294
rect 52502 1230 52566 1294
rect 54134 1230 54198 1294
rect 55494 1230 55558 1294
rect 57534 1230 57598 1294
rect 59438 1230 59502 1294
rect 60798 1230 60862 1294
rect 62566 1230 62630 1294
rect 64334 1230 64398 1294
rect 65830 1230 65894 1294
rect 67598 1230 67662 1294
rect 69230 1230 69294 1294
rect 70862 1230 70926 1294
rect 72766 1230 72830 1294
rect 74262 1230 74326 1294
rect 76166 1230 76230 1294
rect 77662 1230 77726 1294
rect 79294 1230 79358 1294
rect 81062 1230 81126 1294
rect 82830 1230 82894 1294
rect 84326 1230 84390 1294
rect 86230 1230 86294 1294
rect 87726 1230 87790 1294
rect 89358 1230 89422 1294
rect 91262 1230 91326 1294
rect 92758 1230 92822 1294
rect 94390 1230 94454 1294
rect 96158 1230 96222 1294
rect 97790 1230 97854 1294
rect 99558 1230 99622 1294
rect 101326 1230 101390 1294
rect 102822 1230 102886 1294
rect 104590 1230 104654 1294
rect 106222 1230 106286 1294
rect 107854 1230 107918 1294
rect 109758 1230 109822 1294
rect 111254 1230 111318 1294
rect 113022 1230 113086 1294
rect 114790 1230 114854 1294
rect 116286 1230 116350 1294
rect 118054 1230 118118 1294
rect 119822 1230 119886 1294
rect 121318 1230 121382 1294
rect 123086 1230 123150 1294
rect 124718 1230 124782 1294
rect 126350 1230 126414 1294
rect 127982 1230 128046 1294
rect 129750 1230 129814 1294
rect 131518 1230 131582 1294
rect 133150 1230 133214 1294
rect 135326 1230 135390 1294
rect 135462 1230 135526 1294
rect 135598 1230 135662 1294
rect 958 1094 1022 1158
rect 1094 1094 1158 1158
rect 1230 1094 1294 1158
rect 135326 1094 135390 1158
rect 135462 1094 135526 1158
rect 135598 1094 135662 1158
rect 958 958 1022 1022
rect 1094 958 1158 1022
rect 1230 958 1294 1022
rect 135326 958 135390 1022
rect 135462 958 135526 1022
rect 135598 958 135662 1022
rect 278 550 342 614
rect 414 550 478 614
rect 550 550 614 614
rect 39718 550 39782 614
rect 136006 550 136070 614
rect 136142 550 136206 614
rect 136278 550 136342 614
rect 278 414 342 478
rect 414 414 478 478
rect 550 414 614 478
rect 136006 414 136070 478
rect 136142 414 136206 478
rect 136278 414 136342 478
rect 278 278 342 342
rect 414 278 478 342
rect 550 278 614 342
rect 136006 278 136070 342
rect 136142 278 136206 342
rect 136278 278 136342 342
<< metal4 >>
rect 272 83030 620 83036
rect 272 82966 278 83030
rect 342 82966 414 83030
rect 478 82966 550 83030
rect 614 82966 620 83030
rect 272 82894 620 82966
rect 272 82830 278 82894
rect 342 82830 414 82894
rect 478 82830 550 82894
rect 614 82830 620 82894
rect 272 82758 620 82830
rect 272 82694 278 82758
rect 342 82694 414 82758
rect 478 82694 550 82758
rect 614 82694 620 82758
rect 272 23190 620 82694
rect 272 23126 550 23190
rect 614 23126 620 23190
rect 272 14758 620 23126
rect 272 14694 550 14758
rect 614 14694 620 14758
rect 272 10270 620 14694
rect 272 10206 550 10270
rect 614 10206 620 10270
rect 272 7686 620 10206
rect 272 7622 550 7686
rect 614 7622 620 7686
rect 272 614 620 7622
rect 952 82350 1300 82356
rect 952 82286 958 82350
rect 1022 82286 1094 82350
rect 1158 82286 1230 82350
rect 1294 82286 1300 82350
rect 952 82214 1300 82286
rect 952 82150 958 82214
rect 1022 82150 1094 82214
rect 1158 82150 1230 82214
rect 1294 82150 1300 82214
rect 952 82078 1300 82150
rect 952 82014 958 82078
rect 1022 82014 1094 82078
rect 1158 82014 1230 82078
rect 1294 82014 1300 82078
rect 952 79494 1300 82014
rect 2176 82078 2252 82084
rect 2176 82014 2182 82078
rect 2246 82014 2252 82078
rect 2176 81534 2252 82014
rect 2176 81502 2182 81534
rect 2181 81470 2182 81502
rect 2246 81502 2252 81534
rect 3944 82078 4020 82084
rect 3944 82014 3950 82078
rect 4014 82014 4020 82078
rect 3944 81534 4020 82014
rect 3944 81502 3950 81534
rect 2246 81470 2247 81502
rect 2181 81469 2247 81470
rect 3949 81470 3950 81502
rect 4014 81502 4020 81534
rect 5440 82078 5516 82084
rect 5440 82014 5446 82078
rect 5510 82014 5516 82078
rect 5440 81534 5516 82014
rect 5440 81502 5446 81534
rect 4014 81470 4015 81502
rect 3949 81469 4015 81470
rect 5445 81470 5446 81502
rect 5510 81502 5516 81534
rect 7208 82078 7284 82084
rect 7208 82014 7214 82078
rect 7278 82014 7284 82078
rect 7208 81534 7284 82014
rect 7208 81502 7214 81534
rect 5510 81470 5511 81502
rect 5445 81469 5511 81470
rect 7213 81470 7214 81502
rect 7278 81502 7284 81534
rect 8704 82078 8780 82084
rect 8704 82014 8710 82078
rect 8774 82014 8780 82078
rect 8704 81534 8780 82014
rect 8704 81502 8710 81534
rect 7278 81470 7279 81502
rect 7213 81469 7279 81470
rect 8709 81470 8710 81502
rect 8774 81502 8780 81534
rect 10472 82078 10548 82084
rect 10472 82014 10478 82078
rect 10542 82014 10548 82078
rect 10472 81534 10548 82014
rect 10472 81502 10478 81534
rect 8774 81470 8775 81502
rect 8709 81469 8775 81470
rect 10477 81470 10478 81502
rect 10542 81502 10548 81534
rect 12104 82078 12180 82084
rect 12104 82014 12110 82078
rect 12174 82014 12180 82078
rect 12104 81534 12180 82014
rect 12104 81502 12110 81534
rect 10542 81470 10543 81502
rect 10477 81469 10543 81470
rect 12109 81470 12110 81502
rect 12174 81502 12180 81534
rect 14008 82078 14084 82084
rect 14008 82014 14014 82078
rect 14078 82014 14084 82078
rect 14008 81534 14084 82014
rect 14008 81502 14014 81534
rect 12174 81470 12175 81502
rect 12109 81469 12175 81470
rect 14013 81470 14014 81502
rect 14078 81502 14084 81534
rect 15640 82078 15716 82084
rect 15640 82014 15646 82078
rect 15710 82014 15716 82078
rect 15640 81534 15716 82014
rect 15640 81502 15646 81534
rect 14078 81470 14079 81502
rect 14013 81469 14079 81470
rect 15645 81470 15646 81502
rect 15710 81502 15716 81534
rect 17136 82078 17212 82084
rect 17136 82014 17142 82078
rect 17206 82014 17212 82078
rect 17136 81534 17212 82014
rect 17136 81502 17142 81534
rect 15710 81470 15711 81502
rect 15645 81469 15711 81470
rect 17141 81470 17142 81502
rect 17206 81502 17212 81534
rect 18904 82078 18980 82084
rect 18904 82014 18910 82078
rect 18974 82014 18980 82078
rect 18904 81534 18980 82014
rect 18904 81502 18910 81534
rect 17206 81470 17207 81502
rect 17141 81469 17207 81470
rect 18909 81470 18910 81502
rect 18974 81502 18980 81534
rect 20672 82078 20748 82084
rect 20672 82014 20678 82078
rect 20742 82014 20748 82078
rect 20672 81534 20748 82014
rect 20672 81502 20678 81534
rect 18974 81470 18975 81502
rect 18909 81469 18975 81470
rect 20677 81470 20678 81502
rect 20742 81502 20748 81534
rect 22168 82078 22244 82084
rect 22168 82014 22174 82078
rect 22238 82014 22244 82078
rect 22168 81534 22244 82014
rect 22168 81502 22174 81534
rect 20742 81470 20743 81502
rect 20677 81469 20743 81470
rect 22173 81470 22174 81502
rect 22238 81502 22244 81534
rect 23936 82078 24012 82084
rect 23936 82014 23942 82078
rect 24006 82014 24012 82078
rect 23936 81534 24012 82014
rect 23936 81502 23942 81534
rect 22238 81470 22239 81502
rect 22173 81469 22239 81470
rect 23941 81470 23942 81502
rect 24006 81502 24012 81534
rect 25704 82078 25780 82084
rect 25704 82014 25710 82078
rect 25774 82014 25780 82078
rect 25704 81534 25780 82014
rect 25704 81502 25710 81534
rect 24006 81470 24007 81502
rect 23941 81469 24007 81470
rect 25709 81470 25710 81502
rect 25774 81502 25780 81534
rect 27200 82078 27276 82084
rect 27200 82014 27206 82078
rect 27270 82014 27276 82078
rect 27200 81534 27276 82014
rect 27200 81502 27206 81534
rect 25774 81470 25775 81502
rect 25709 81469 25775 81470
rect 27205 81470 27206 81502
rect 27270 81502 27276 81534
rect 27270 81470 27271 81502
rect 27205 81469 27271 81470
rect 2040 81398 2116 81404
rect 2040 81334 2046 81398
rect 2110 81334 2116 81398
rect 2040 81126 2116 81334
rect 2040 81094 2046 81126
rect 2045 81062 2046 81094
rect 2110 81094 2116 81126
rect 2110 81062 2111 81094
rect 2045 81061 2111 81062
rect 952 79430 1230 79494
rect 1294 79430 1300 79494
rect 952 77590 1300 79430
rect 952 77526 1230 77590
rect 1294 77526 1300 77590
rect 952 76094 1300 77526
rect 28696 77182 28772 83308
rect 28968 82078 29044 82084
rect 28968 82014 28974 82078
rect 29038 82014 29044 82078
rect 28968 81534 29044 82014
rect 28968 81502 28974 81534
rect 28973 81470 28974 81502
rect 29038 81502 29044 81534
rect 30600 82078 30676 82084
rect 30600 82014 30606 82078
rect 30670 82014 30676 82078
rect 30600 81534 30676 82014
rect 30600 81502 30606 81534
rect 29038 81470 29039 81502
rect 28973 81469 29039 81470
rect 30605 81470 30606 81502
rect 30670 81502 30676 81534
rect 30670 81470 30671 81502
rect 30605 81469 30671 81470
rect 28696 77150 28702 77182
rect 28701 77118 28702 77150
rect 28766 77150 28772 77182
rect 31008 77182 31084 83308
rect 32368 82078 32444 82084
rect 32368 82014 32374 82078
rect 32438 82014 32444 82078
rect 32368 81534 32444 82014
rect 32368 81502 32374 81534
rect 32373 81470 32374 81502
rect 32438 81502 32444 81534
rect 32438 81470 32439 81502
rect 32373 81469 32439 81470
rect 31008 77150 31014 77182
rect 28766 77118 28767 77150
rect 28701 77117 28767 77118
rect 31013 77118 31014 77150
rect 31078 77150 31084 77182
rect 33456 77182 33532 83308
rect 34136 82078 34212 82084
rect 34136 82014 34142 82078
rect 34206 82014 34212 82078
rect 34136 81534 34212 82014
rect 34136 81502 34142 81534
rect 34141 81470 34142 81502
rect 34206 81502 34212 81534
rect 35632 82078 35708 82084
rect 35632 82014 35638 82078
rect 35702 82014 35708 82078
rect 35632 81534 35708 82014
rect 35632 81502 35638 81534
rect 34206 81470 34207 81502
rect 34141 81469 34207 81470
rect 35637 81470 35638 81502
rect 35702 81502 35708 81534
rect 35702 81470 35703 81502
rect 35637 81469 35703 81470
rect 33456 77150 33462 77182
rect 31078 77118 31079 77150
rect 31013 77117 31079 77118
rect 33461 77118 33462 77150
rect 33526 77150 33532 77182
rect 36176 77182 36252 83308
rect 37536 82078 37612 82084
rect 37536 82014 37542 82078
rect 37606 82014 37612 82078
rect 37536 81534 37612 82014
rect 37536 81502 37542 81534
rect 37541 81470 37542 81502
rect 37606 81502 37612 81534
rect 37606 81470 37607 81502
rect 37541 81469 37607 81470
rect 36176 77150 36182 77182
rect 33526 77118 33527 77150
rect 33461 77117 33527 77118
rect 36181 77118 36182 77150
rect 36246 77150 36252 77182
rect 38488 77182 38564 83308
rect 39168 82078 39244 82084
rect 39168 82014 39174 82078
rect 39238 82014 39244 82078
rect 39168 81534 39244 82014
rect 39168 81502 39174 81534
rect 39173 81470 39174 81502
rect 39238 81502 39244 81534
rect 40664 82078 40740 82084
rect 40664 82014 40670 82078
rect 40734 82014 40740 82078
rect 40664 81534 40740 82014
rect 40664 81502 40670 81534
rect 39238 81470 39239 81502
rect 39173 81469 39239 81470
rect 40669 81470 40670 81502
rect 40734 81502 40740 81534
rect 40734 81470 40735 81502
rect 40669 81469 40735 81470
rect 38488 77150 38494 77182
rect 36246 77118 36247 77150
rect 36181 77117 36247 77118
rect 38493 77118 38494 77150
rect 38558 77150 38564 77182
rect 41072 77182 41148 83308
rect 42432 82078 42508 82084
rect 42432 82014 42438 82078
rect 42502 82014 42508 82078
rect 42432 81534 42508 82014
rect 42432 81502 42438 81534
rect 42437 81470 42438 81502
rect 42502 81502 42508 81534
rect 42502 81470 42503 81502
rect 42437 81469 42503 81470
rect 41072 77150 41078 77182
rect 38558 77118 38559 77150
rect 38493 77117 38559 77118
rect 41077 77118 41078 77150
rect 41142 77150 41148 77182
rect 43520 77182 43596 83308
rect 44200 82078 44276 82084
rect 44200 82014 44206 82078
rect 44270 82014 44276 82078
rect 44200 81534 44276 82014
rect 44200 81502 44206 81534
rect 44205 81470 44206 81502
rect 44270 81502 44276 81534
rect 45696 82078 45772 82084
rect 45696 82014 45702 82078
rect 45766 82014 45772 82078
rect 45696 81534 45772 82014
rect 45696 81502 45702 81534
rect 44270 81470 44271 81502
rect 44205 81469 44271 81470
rect 45701 81470 45702 81502
rect 45766 81502 45772 81534
rect 45766 81470 45767 81502
rect 45701 81469 45767 81470
rect 43520 77150 43526 77182
rect 41142 77118 41143 77150
rect 41077 77117 41143 77118
rect 43525 77118 43526 77150
rect 43590 77150 43596 77182
rect 46104 77182 46180 83308
rect 47464 82078 47540 82084
rect 47464 82014 47470 82078
rect 47534 82014 47540 82078
rect 47464 81534 47540 82014
rect 47464 81502 47470 81534
rect 47469 81470 47470 81502
rect 47534 81502 47540 81534
rect 47534 81470 47535 81502
rect 47469 81469 47535 81470
rect 46104 77150 46110 77182
rect 43590 77118 43591 77150
rect 43525 77117 43591 77118
rect 46109 77118 46110 77150
rect 46174 77150 46180 77182
rect 48552 77182 48628 83308
rect 49232 82078 49308 82084
rect 49232 82014 49238 82078
rect 49302 82014 49308 82078
rect 49232 81534 49308 82014
rect 49232 81502 49238 81534
rect 49237 81470 49238 81502
rect 49302 81502 49308 81534
rect 50728 82078 50804 82084
rect 50728 82014 50734 82078
rect 50798 82014 50804 82078
rect 50728 81534 50804 82014
rect 50728 81502 50734 81534
rect 49302 81470 49303 81502
rect 49237 81469 49303 81470
rect 50733 81470 50734 81502
rect 50798 81502 50804 81534
rect 50798 81470 50799 81502
rect 50733 81469 50799 81470
rect 48552 77150 48558 77182
rect 46174 77118 46175 77150
rect 46109 77117 46175 77118
rect 48557 77118 48558 77150
rect 48622 77150 48628 77182
rect 51136 77182 51212 83308
rect 52632 82078 52708 82084
rect 52632 82014 52638 82078
rect 52702 82014 52708 82078
rect 52632 81534 52708 82014
rect 52632 81502 52638 81534
rect 52637 81470 52638 81502
rect 52702 81502 52708 81534
rect 52702 81470 52703 81502
rect 52637 81469 52703 81470
rect 51136 77150 51142 77182
rect 48622 77118 48623 77150
rect 48557 77117 48623 77118
rect 51141 77118 51142 77150
rect 51206 77150 51212 77182
rect 53584 77182 53660 83308
rect 54128 82078 54204 82084
rect 54128 82014 54134 82078
rect 54198 82014 54204 82078
rect 54128 81534 54204 82014
rect 54128 81502 54134 81534
rect 54133 81470 54134 81502
rect 54198 81502 54204 81534
rect 55896 82078 55972 82084
rect 55896 82014 55902 82078
rect 55966 82014 55972 82078
rect 55896 81534 55972 82014
rect 55896 81502 55902 81534
rect 54198 81470 54199 81502
rect 54133 81469 54199 81470
rect 55901 81470 55902 81502
rect 55966 81502 55972 81534
rect 55966 81470 55967 81502
rect 55901 81469 55967 81470
rect 53584 77150 53590 77182
rect 51206 77118 51207 77150
rect 51141 77117 51207 77118
rect 53589 77118 53590 77150
rect 53654 77150 53660 77182
rect 56168 77182 56244 83308
rect 57664 82078 57740 82084
rect 57664 82014 57670 82078
rect 57734 82014 57740 82078
rect 57664 81534 57740 82014
rect 57664 81502 57670 81534
rect 57669 81470 57670 81502
rect 57734 81502 57740 81534
rect 57734 81470 57735 81502
rect 57669 81469 57735 81470
rect 56168 77150 56174 77182
rect 53654 77118 53655 77150
rect 53589 77117 53655 77118
rect 56173 77118 56174 77150
rect 56238 77150 56244 77182
rect 58480 77182 58556 83308
rect 59160 82078 59236 82084
rect 59160 82014 59166 82078
rect 59230 82014 59236 82078
rect 59160 81534 59236 82014
rect 59160 81502 59166 81534
rect 59165 81470 59166 81502
rect 59230 81502 59236 81534
rect 60792 82078 60868 82084
rect 60792 82014 60798 82078
rect 60862 82014 60868 82078
rect 60792 81534 60868 82014
rect 60792 81502 60798 81534
rect 59230 81470 59231 81502
rect 59165 81469 59231 81470
rect 60797 81470 60798 81502
rect 60862 81502 60868 81534
rect 60862 81470 60863 81502
rect 60797 81469 60863 81470
rect 58480 77150 58486 77182
rect 56238 77118 56239 77150
rect 56173 77117 56239 77118
rect 58485 77118 58486 77150
rect 58550 77150 58556 77182
rect 60928 77182 61004 83308
rect 62696 82078 62772 82084
rect 62696 82014 62702 82078
rect 62766 82014 62772 82078
rect 62696 81534 62772 82014
rect 62696 81502 62702 81534
rect 62701 81470 62702 81502
rect 62766 81502 62772 81534
rect 62766 81470 62767 81502
rect 62701 81469 62767 81470
rect 60928 77150 60934 77182
rect 58550 77118 58551 77150
rect 58485 77117 58551 77118
rect 60933 77118 60934 77150
rect 60998 77150 61004 77182
rect 61477 77182 61543 77183
rect 61477 77150 61478 77182
rect 60998 77118 60999 77150
rect 60933 77117 60999 77118
rect 61472 77118 61478 77150
rect 61542 77150 61543 77182
rect 63648 77182 63724 83308
rect 64192 82078 64268 82084
rect 64192 82014 64198 82078
rect 64262 82014 64268 82078
rect 64192 81534 64268 82014
rect 64192 81502 64198 81534
rect 64197 81470 64198 81502
rect 64262 81502 64268 81534
rect 65824 82078 65900 82084
rect 65824 82014 65830 82078
rect 65894 82014 65900 82078
rect 65824 81534 65900 82014
rect 65824 81502 65830 81534
rect 64262 81470 64263 81502
rect 64197 81469 64263 81470
rect 65829 81470 65830 81502
rect 65894 81502 65900 81534
rect 65894 81470 65895 81502
rect 65829 81469 65895 81470
rect 63648 77150 63654 77182
rect 61542 77118 61548 77150
rect 28973 77046 29039 77047
rect 28973 77014 28974 77046
rect 28968 76982 28974 77014
rect 29038 77014 29039 77046
rect 31421 77046 31487 77047
rect 31421 77014 31422 77046
rect 29038 76982 29044 77014
rect 28968 76780 29044 76982
rect 952 76030 1230 76094
rect 1294 76030 1300 76094
rect 952 74190 1300 76030
rect 28832 76704 29044 76780
rect 31416 76982 31422 77014
rect 31486 77014 31487 77046
rect 34005 77046 34071 77047
rect 34005 77014 34006 77046
rect 31486 76982 31492 77014
rect 28832 75278 28908 76704
rect 28968 76638 29044 76644
rect 28968 76574 28974 76638
rect 29038 76574 29044 76638
rect 28968 75958 29044 76574
rect 28968 75926 28974 75958
rect 28973 75894 28974 75926
rect 29038 75926 29044 75958
rect 31280 76638 31356 76644
rect 31280 76574 31286 76638
rect 31350 76574 31356 76638
rect 31280 75958 31356 76574
rect 31280 75926 31286 75958
rect 29038 75894 29039 75926
rect 28973 75893 29039 75894
rect 31285 75894 31286 75926
rect 31350 75926 31356 75958
rect 31350 75894 31351 75926
rect 31285 75893 31351 75894
rect 28832 75214 28838 75278
rect 28902 75214 28908 75278
rect 28832 75208 28908 75214
rect 31416 75278 31492 76982
rect 34000 76982 34006 77014
rect 34070 77014 34071 77046
rect 36453 77046 36519 77047
rect 36453 77014 36454 77046
rect 34070 76982 34076 77014
rect 33728 76638 33804 76644
rect 33728 76574 33734 76638
rect 33798 76574 33804 76638
rect 33728 75958 33804 76574
rect 33728 75926 33734 75958
rect 33733 75894 33734 75926
rect 33798 75926 33804 75958
rect 33798 75894 33799 75926
rect 33733 75893 33799 75894
rect 31416 75214 31422 75278
rect 31486 75214 31492 75278
rect 31416 75208 31492 75214
rect 34000 75278 34076 76982
rect 36448 76982 36454 77014
rect 36518 77014 36519 77046
rect 39037 77046 39103 77047
rect 39037 77014 39038 77046
rect 36518 76982 36524 77014
rect 36312 76638 36388 76644
rect 36312 76574 36318 76638
rect 36382 76574 36388 76638
rect 36312 75958 36388 76574
rect 36312 75926 36318 75958
rect 36317 75894 36318 75926
rect 36382 75926 36388 75958
rect 36382 75894 36383 75926
rect 36317 75893 36383 75894
rect 34000 75214 34006 75278
rect 34070 75214 34076 75278
rect 34000 75208 34076 75214
rect 36448 75278 36524 76982
rect 39032 76982 39038 77014
rect 39102 77014 39103 77046
rect 41485 77046 41551 77047
rect 41485 77014 41486 77046
rect 39102 76982 39108 77014
rect 38629 76638 38695 76639
rect 38629 76606 38630 76638
rect 38624 76574 38630 76606
rect 38694 76606 38695 76638
rect 38896 76638 38972 76644
rect 38694 76574 38700 76606
rect 38624 75958 38700 76574
rect 38624 75894 38630 75958
rect 38694 75894 38700 75958
rect 38896 76574 38902 76638
rect 38966 76574 38972 76638
rect 38896 75958 38972 76574
rect 38896 75926 38902 75958
rect 38624 75888 38700 75894
rect 38901 75894 38902 75926
rect 38966 75926 38972 75958
rect 38966 75894 38967 75926
rect 38901 75893 38967 75894
rect 36448 75214 36454 75278
rect 36518 75214 36524 75278
rect 36448 75208 36524 75214
rect 39032 75278 39108 76982
rect 41480 76982 41486 77014
rect 41550 77014 41551 77046
rect 43933 77046 43999 77047
rect 43933 77014 43934 77046
rect 41550 76982 41556 77014
rect 41344 76638 41420 76644
rect 41344 76574 41350 76638
rect 41414 76574 41420 76638
rect 41344 75958 41420 76574
rect 41344 75926 41350 75958
rect 41349 75894 41350 75926
rect 41414 75926 41420 75958
rect 41414 75894 41415 75926
rect 41349 75893 41415 75894
rect 39032 75214 39038 75278
rect 39102 75214 39108 75278
rect 39032 75208 39108 75214
rect 41480 75278 41556 76982
rect 43928 76982 43934 77014
rect 43998 77014 43999 77046
rect 46517 77046 46583 77047
rect 46517 77014 46518 77046
rect 43998 76982 44004 77014
rect 43928 76780 44004 76982
rect 43792 76704 44004 76780
rect 46512 76982 46518 77014
rect 46582 77014 46583 77046
rect 48965 77046 49031 77047
rect 48965 77014 48966 77046
rect 46582 76982 46588 77014
rect 43661 76638 43727 76639
rect 43661 76606 43662 76638
rect 43656 76574 43662 76606
rect 43726 76606 43727 76638
rect 43726 76574 43732 76606
rect 43656 75958 43732 76574
rect 43656 75894 43662 75958
rect 43726 75894 43732 75958
rect 43656 75888 43732 75894
rect 41480 75214 41486 75278
rect 41550 75214 41556 75278
rect 41480 75208 41556 75214
rect 43792 75278 43868 76704
rect 43928 76638 44004 76644
rect 43928 76574 43934 76638
rect 43998 76574 44004 76638
rect 43928 75958 44004 76574
rect 43928 75926 43934 75958
rect 43933 75894 43934 75926
rect 43998 75926 44004 75958
rect 46376 76638 46452 76644
rect 46376 76574 46382 76638
rect 46446 76574 46452 76638
rect 46376 75958 46452 76574
rect 46376 75926 46382 75958
rect 43998 75894 43999 75926
rect 43933 75893 43999 75894
rect 46381 75894 46382 75926
rect 46446 75926 46452 75958
rect 46446 75894 46447 75926
rect 46381 75893 46447 75894
rect 43792 75214 43798 75278
rect 43862 75214 43868 75278
rect 43792 75208 43868 75214
rect 46512 75278 46588 76982
rect 48960 76982 48966 77014
rect 49030 77014 49031 77046
rect 51413 77046 51479 77047
rect 51413 77014 51414 77046
rect 49030 76982 49036 77014
rect 48688 76638 48764 76644
rect 48688 76574 48694 76638
rect 48758 76574 48764 76638
rect 48688 75958 48764 76574
rect 48688 75926 48694 75958
rect 48693 75894 48694 75926
rect 48758 75926 48764 75958
rect 48758 75894 48759 75926
rect 48693 75893 48759 75894
rect 46512 75214 46518 75278
rect 46582 75214 46588 75278
rect 46512 75208 46588 75214
rect 48960 75278 49036 76982
rect 51408 76982 51414 77014
rect 51478 77014 51479 77046
rect 53861 77046 53927 77047
rect 53861 77014 53862 77046
rect 51478 76982 51484 77014
rect 51408 76780 51484 76982
rect 48960 75214 48966 75278
rect 49030 75214 49036 75278
rect 48960 75208 49036 75214
rect 51272 76704 51484 76780
rect 53856 76982 53862 77014
rect 53926 77014 53927 77046
rect 56445 77046 56511 77047
rect 56445 77014 56446 77046
rect 53926 76982 53932 77014
rect 51272 75278 51348 76704
rect 51408 76638 51484 76644
rect 51408 76574 51414 76638
rect 51478 76574 51484 76638
rect 51408 75958 51484 76574
rect 51408 75926 51414 75958
rect 51413 75894 51414 75926
rect 51478 75926 51484 75958
rect 53720 76638 53796 76644
rect 53720 76574 53726 76638
rect 53790 76574 53796 76638
rect 53720 75958 53796 76574
rect 53720 75926 53726 75958
rect 51478 75894 51479 75926
rect 51413 75893 51479 75894
rect 53725 75894 53726 75926
rect 53790 75926 53796 75958
rect 53790 75894 53791 75926
rect 53725 75893 53791 75894
rect 51272 75214 51278 75278
rect 51342 75214 51348 75278
rect 51272 75208 51348 75214
rect 53856 75278 53932 76982
rect 56440 76982 56446 77014
rect 56510 77014 56511 77046
rect 58893 77046 58959 77047
rect 58893 77014 58894 77046
rect 56510 76982 56516 77014
rect 56173 76638 56239 76639
rect 56173 76606 56174 76638
rect 56168 76574 56174 76606
rect 56238 76606 56239 76638
rect 56304 76638 56380 76644
rect 56238 76574 56244 76606
rect 56168 75958 56244 76574
rect 56168 75894 56174 75958
rect 56238 75894 56244 75958
rect 56304 76574 56310 76638
rect 56374 76574 56380 76638
rect 56304 75958 56380 76574
rect 56304 75926 56310 75958
rect 56168 75888 56244 75894
rect 56309 75894 56310 75926
rect 56374 75926 56380 75958
rect 56374 75894 56375 75926
rect 56309 75893 56375 75894
rect 53856 75214 53862 75278
rect 53926 75214 53932 75278
rect 53856 75208 53932 75214
rect 56440 75278 56516 76982
rect 58888 76982 58894 77014
rect 58958 77014 58959 77046
rect 58958 76982 58964 77014
rect 58752 76638 58828 76644
rect 58752 76574 58758 76638
rect 58822 76574 58828 76638
rect 58752 75958 58828 76574
rect 58752 75926 58758 75958
rect 58757 75894 58758 75926
rect 58822 75926 58828 75958
rect 58822 75894 58823 75926
rect 58757 75893 58823 75894
rect 56440 75214 56446 75278
rect 56510 75214 56516 75278
rect 56440 75208 56516 75214
rect 58888 75278 58964 76982
rect 61336 76638 61412 76644
rect 61336 76574 61342 76638
rect 61406 76574 61412 76638
rect 61336 75958 61412 76574
rect 61336 75926 61342 75958
rect 61341 75894 61342 75926
rect 61406 75926 61412 75958
rect 61406 75894 61407 75926
rect 61341 75893 61407 75894
rect 59437 75822 59503 75823
rect 59437 75790 59438 75822
rect 58888 75214 58894 75278
rect 58958 75214 58964 75278
rect 58888 75208 58964 75214
rect 59432 75758 59438 75790
rect 59502 75790 59503 75822
rect 59502 75758 59508 75790
rect 28973 75142 29039 75143
rect 28973 75110 28974 75142
rect 952 74126 1230 74190
rect 1294 74126 1300 74190
rect 952 72694 1300 74126
rect 28968 75078 28974 75110
rect 29038 75110 29039 75142
rect 31557 75142 31623 75143
rect 31557 75110 31558 75142
rect 29038 75078 29044 75110
rect 28968 73238 29044 75078
rect 28968 73174 28974 73238
rect 29038 73174 29044 73238
rect 28968 73168 29044 73174
rect 31552 75078 31558 75110
rect 31622 75110 31623 75142
rect 34005 75142 34071 75143
rect 34005 75110 34006 75142
rect 31622 75078 31628 75110
rect 31552 73238 31628 75078
rect 31552 73174 31558 73238
rect 31622 73174 31628 73238
rect 31552 73168 31628 73174
rect 34000 75078 34006 75110
rect 34070 75110 34071 75142
rect 36453 75142 36519 75143
rect 36453 75110 36454 75142
rect 34070 75078 34076 75110
rect 34000 73238 34076 75078
rect 34000 73174 34006 73238
rect 34070 73174 34076 73238
rect 34000 73168 34076 73174
rect 36448 75078 36454 75110
rect 36518 75110 36519 75142
rect 39037 75142 39103 75143
rect 39037 75110 39038 75142
rect 36518 75078 36524 75110
rect 36448 73238 36524 75078
rect 36448 73174 36454 73238
rect 36518 73174 36524 73238
rect 36448 73168 36524 73174
rect 39032 75078 39038 75110
rect 39102 75110 39103 75142
rect 41485 75142 41551 75143
rect 41485 75110 41486 75142
rect 39102 75078 39108 75110
rect 39032 73238 39108 75078
rect 39032 73174 39038 73238
rect 39102 73174 39108 73238
rect 39032 73168 39108 73174
rect 41480 75078 41486 75110
rect 41550 75110 41551 75142
rect 44069 75142 44135 75143
rect 44069 75110 44070 75142
rect 41550 75078 41556 75110
rect 41480 73238 41556 75078
rect 41480 73174 41486 73238
rect 41550 73174 41556 73238
rect 41480 73168 41556 73174
rect 44064 75078 44070 75110
rect 44134 75110 44135 75142
rect 46517 75142 46583 75143
rect 46517 75110 46518 75142
rect 44134 75078 44140 75110
rect 44064 73238 44140 75078
rect 44064 73174 44070 73238
rect 44134 73174 44140 73238
rect 44064 73168 44140 73174
rect 46512 75078 46518 75110
rect 46582 75110 46583 75142
rect 48965 75142 49031 75143
rect 48965 75110 48966 75142
rect 46582 75078 46588 75110
rect 46512 73238 46588 75078
rect 46512 73174 46518 73238
rect 46582 73174 46588 73238
rect 46512 73168 46588 73174
rect 48960 75078 48966 75110
rect 49030 75110 49031 75142
rect 51549 75142 51615 75143
rect 51549 75110 51550 75142
rect 49030 75078 49036 75110
rect 48960 73238 49036 75078
rect 48960 73174 48966 73238
rect 49030 73174 49036 73238
rect 48960 73168 49036 73174
rect 51544 75078 51550 75110
rect 51614 75110 51615 75142
rect 53997 75142 54063 75143
rect 53997 75110 53998 75142
rect 51614 75078 51620 75110
rect 51544 73238 51620 75078
rect 51544 73174 51550 73238
rect 51614 73174 51620 73238
rect 51544 73168 51620 73174
rect 53992 75078 53998 75110
rect 54062 75110 54063 75142
rect 56304 75142 56380 75148
rect 54062 75078 54068 75110
rect 53992 73238 54068 75078
rect 53992 73174 53998 73238
rect 54062 73174 54068 73238
rect 56304 75078 56310 75142
rect 56374 75078 56380 75142
rect 59029 75142 59095 75143
rect 59029 75110 59030 75142
rect 56304 73238 56380 75078
rect 56304 73206 56310 73238
rect 53992 73168 54068 73174
rect 56309 73174 56310 73206
rect 56374 73206 56380 73238
rect 59024 75078 59030 75110
rect 59094 75110 59095 75142
rect 59094 75078 59100 75110
rect 59024 73238 59100 75078
rect 56374 73174 56375 73206
rect 56309 73173 56375 73174
rect 59024 73174 59030 73238
rect 59094 73174 59100 73238
rect 59024 73168 59100 73174
rect 952 72630 1230 72694
rect 1294 72630 1300 72694
rect 952 71062 1300 72630
rect 28968 73102 29044 73108
rect 28968 73038 28974 73102
rect 29038 73038 29044 73102
rect 952 70998 1230 71062
rect 1294 70998 1300 71062
rect 28560 71470 28636 71476
rect 28560 71406 28566 71470
rect 28630 71406 28636 71470
rect 28701 71470 28767 71471
rect 28701 71438 28702 71470
rect 28560 71062 28636 71406
rect 28560 71030 28566 71062
rect 952 69294 1300 70998
rect 28565 70998 28566 71030
rect 28630 71030 28636 71062
rect 28696 71406 28702 71438
rect 28766 71438 28767 71470
rect 28766 71406 28772 71438
rect 28696 71062 28772 71406
rect 28630 70998 28631 71030
rect 28565 70997 28631 70998
rect 28696 70998 28702 71062
rect 28766 70998 28772 71062
rect 28696 70992 28772 70998
rect 28968 70790 29044 73038
rect 59432 71606 59508 75758
rect 61472 75278 61548 77118
rect 63653 77118 63654 77150
rect 63718 77150 63724 77182
rect 66096 77182 66172 83308
rect 67592 82078 67668 82084
rect 67592 82014 67598 82078
rect 67662 82014 67668 82078
rect 67592 81534 67668 82014
rect 67592 81502 67598 81534
rect 67597 81470 67598 81502
rect 67662 81502 67668 81534
rect 67662 81470 67663 81502
rect 67597 81469 67663 81470
rect 66096 77150 66102 77182
rect 63718 77118 63719 77150
rect 63653 77117 63719 77118
rect 66101 77118 66102 77150
rect 66166 77150 66172 77182
rect 68544 77182 68620 83308
rect 69224 82078 69300 82084
rect 69224 82014 69230 82078
rect 69294 82014 69300 82078
rect 69224 81534 69300 82014
rect 69224 81502 69230 81534
rect 69229 81470 69230 81502
rect 69294 81502 69300 81534
rect 70856 82078 70932 82084
rect 70856 82014 70862 82078
rect 70926 82014 70932 82078
rect 70856 81534 70932 82014
rect 70856 81502 70862 81534
rect 69294 81470 69295 81502
rect 69229 81469 69295 81470
rect 70861 81470 70862 81502
rect 70926 81502 70932 81534
rect 70926 81470 70927 81502
rect 70861 81469 70927 81470
rect 68544 77150 68550 77182
rect 66166 77118 66167 77150
rect 66101 77117 66167 77118
rect 68549 77118 68550 77150
rect 68614 77150 68620 77182
rect 68957 77182 69023 77183
rect 68957 77150 68958 77182
rect 68614 77118 68615 77150
rect 68549 77117 68615 77118
rect 68952 77118 68958 77150
rect 69022 77150 69023 77182
rect 70992 77182 71068 83308
rect 72624 82078 72700 82084
rect 72624 82014 72630 82078
rect 72694 82014 72700 82078
rect 72624 81534 72700 82014
rect 72624 81502 72630 81534
rect 72629 81470 72630 81502
rect 72694 81502 72700 81534
rect 72694 81470 72695 81502
rect 72629 81469 72695 81470
rect 70992 77150 70998 77182
rect 69022 77118 69028 77150
rect 63925 77046 63991 77047
rect 63925 77014 63926 77046
rect 63920 76982 63926 77014
rect 63990 77014 63991 77046
rect 66509 77046 66575 77047
rect 66509 77014 66510 77046
rect 63990 76982 63996 77014
rect 63784 76638 63860 76644
rect 63784 76574 63790 76638
rect 63854 76574 63860 76638
rect 63784 75958 63860 76574
rect 63784 75926 63790 75958
rect 63789 75894 63790 75926
rect 63854 75926 63860 75958
rect 63854 75894 63855 75926
rect 63789 75893 63855 75894
rect 61472 75214 61478 75278
rect 61542 75214 61548 75278
rect 61472 75208 61548 75214
rect 63920 75278 63996 76982
rect 66504 76982 66510 77014
rect 66574 77014 66575 77046
rect 66574 76982 66580 77014
rect 66368 76638 66444 76644
rect 66368 76574 66374 76638
rect 66438 76574 66444 76638
rect 66368 75958 66444 76574
rect 66368 75926 66374 75958
rect 66373 75894 66374 75926
rect 66438 75926 66444 75958
rect 66438 75894 66439 75926
rect 66373 75893 66439 75894
rect 63920 75214 63926 75278
rect 63990 75214 63996 75278
rect 63920 75208 63996 75214
rect 66504 75278 66580 76982
rect 68816 76638 68892 76644
rect 68816 76574 68822 76638
rect 68886 76574 68892 76638
rect 68816 75958 68892 76574
rect 68816 75926 68822 75958
rect 68821 75894 68822 75926
rect 68886 75926 68892 75958
rect 68886 75894 68887 75926
rect 68821 75893 68887 75894
rect 66504 75214 66510 75278
rect 66574 75214 66580 75278
rect 66504 75208 66580 75214
rect 68952 75278 69028 77118
rect 70997 77118 70998 77150
rect 71062 77150 71068 77182
rect 73576 77182 73652 83308
rect 74392 82078 74468 82084
rect 74392 82014 74398 82078
rect 74462 82014 74468 82078
rect 74392 81534 74468 82014
rect 74392 81502 74398 81534
rect 74397 81470 74398 81502
rect 74462 81502 74468 81534
rect 74462 81470 74463 81502
rect 74397 81469 74463 81470
rect 73576 77150 73582 77182
rect 71062 77118 71063 77150
rect 70997 77117 71063 77118
rect 73581 77118 73582 77150
rect 73646 77150 73652 77182
rect 75888 77182 75964 83308
rect 76160 82078 76236 82084
rect 76160 82014 76166 82078
rect 76230 82014 76236 82078
rect 76160 81534 76236 82014
rect 76160 81502 76166 81534
rect 76165 81470 76166 81502
rect 76230 81502 76236 81534
rect 77656 82078 77732 82084
rect 77656 82014 77662 82078
rect 77726 82014 77732 82078
rect 77656 81534 77732 82014
rect 77656 81502 77662 81534
rect 76230 81470 76231 81502
rect 76165 81469 76231 81470
rect 77661 81470 77662 81502
rect 77726 81502 77732 81534
rect 77726 81470 77727 81502
rect 77661 81469 77727 81470
rect 75888 77150 75894 77182
rect 73646 77118 73647 77150
rect 73581 77117 73647 77118
rect 75893 77118 75894 77150
rect 75958 77150 75964 77182
rect 78608 77182 78684 83308
rect 79424 82078 79500 82084
rect 79424 82014 79430 82078
rect 79494 82014 79500 82078
rect 79424 81534 79500 82014
rect 79424 81502 79430 81534
rect 79429 81470 79430 81502
rect 79494 81502 79500 81534
rect 79494 81470 79495 81502
rect 79429 81469 79495 81470
rect 78608 77150 78614 77182
rect 75958 77118 75959 77150
rect 75893 77117 75959 77118
rect 78613 77118 78614 77150
rect 78678 77150 78684 77182
rect 81056 77182 81132 83308
rect 81328 82078 81404 82084
rect 81328 82014 81334 82078
rect 81398 82014 81404 82078
rect 81328 81534 81404 82014
rect 81328 81502 81334 81534
rect 81333 81470 81334 81502
rect 81398 81502 81404 81534
rect 82688 82078 82764 82084
rect 82688 82014 82694 82078
rect 82758 82014 82764 82078
rect 82688 81534 82764 82014
rect 82688 81502 82694 81534
rect 81398 81470 81399 81502
rect 81333 81469 81399 81470
rect 82693 81470 82694 81502
rect 82758 81502 82764 81534
rect 82758 81470 82759 81502
rect 82693 81469 82759 81470
rect 81056 77150 81062 77182
rect 78678 77118 78679 77150
rect 78613 77117 78679 77118
rect 81061 77118 81062 77150
rect 81126 77150 81132 77182
rect 83504 77182 83580 83308
rect 84456 82078 84532 82084
rect 84456 82014 84462 82078
rect 84526 82014 84532 82078
rect 84456 81534 84532 82014
rect 84456 81502 84462 81534
rect 84461 81470 84462 81502
rect 84526 81502 84532 81534
rect 84526 81470 84527 81502
rect 84461 81469 84527 81470
rect 83504 77150 83510 77182
rect 81126 77118 81127 77150
rect 81061 77117 81127 77118
rect 83509 77118 83510 77150
rect 83574 77150 83580 77182
rect 85952 77182 86028 83308
rect 86224 82078 86300 82084
rect 86224 82014 86230 82078
rect 86294 82014 86300 82078
rect 86224 81534 86300 82014
rect 86224 81502 86230 81534
rect 86229 81470 86230 81502
rect 86294 81502 86300 81534
rect 87720 82078 87796 82084
rect 87720 82014 87726 82078
rect 87790 82014 87796 82078
rect 87720 81534 87796 82014
rect 87720 81502 87726 81534
rect 86294 81470 86295 81502
rect 86229 81469 86295 81470
rect 87725 81470 87726 81502
rect 87790 81502 87796 81534
rect 87790 81470 87791 81502
rect 87725 81469 87791 81470
rect 85952 77150 85958 77182
rect 83574 77118 83575 77150
rect 83509 77117 83575 77118
rect 85957 77118 85958 77150
rect 86022 77150 86028 77182
rect 88400 77182 88476 83308
rect 89352 82078 89428 82084
rect 89352 82014 89358 82078
rect 89422 82014 89428 82078
rect 89352 81534 89428 82014
rect 89352 81502 89358 81534
rect 89357 81470 89358 81502
rect 89422 81502 89428 81534
rect 89422 81470 89423 81502
rect 89357 81469 89423 81470
rect 88400 77150 88406 77182
rect 86022 77118 86023 77150
rect 85957 77117 86023 77118
rect 88405 77118 88406 77150
rect 88470 77150 88476 77182
rect 90984 77182 91060 83308
rect 91120 82078 91196 82084
rect 91120 82014 91126 82078
rect 91190 82014 91196 82078
rect 91120 81534 91196 82014
rect 91120 81502 91126 81534
rect 91125 81470 91126 81502
rect 91190 81502 91196 81534
rect 92888 82078 92964 82084
rect 92888 82014 92894 82078
rect 92958 82014 92964 82078
rect 92888 81534 92964 82014
rect 92888 81502 92894 81534
rect 91190 81470 91191 81502
rect 91125 81469 91191 81470
rect 92893 81470 92894 81502
rect 92958 81502 92964 81534
rect 92958 81470 92959 81502
rect 92893 81469 92959 81470
rect 90984 77150 90990 77182
rect 88470 77118 88471 77150
rect 88405 77117 88471 77118
rect 90989 77118 90990 77150
rect 91054 77150 91060 77182
rect 91261 77182 91327 77183
rect 91261 77150 91262 77182
rect 91054 77118 91055 77150
rect 90989 77117 91055 77118
rect 91256 77118 91262 77150
rect 91326 77150 91327 77182
rect 93568 77182 93644 83308
rect 94384 82078 94460 82084
rect 94384 82014 94390 82078
rect 94454 82014 94460 82078
rect 94384 81534 94460 82014
rect 94384 81502 94390 81534
rect 94389 81470 94390 81502
rect 94454 81502 94460 81534
rect 94454 81470 94455 81502
rect 94389 81469 94455 81470
rect 93568 77150 93574 77182
rect 91326 77118 91332 77150
rect 71405 77046 71471 77047
rect 71405 77014 71406 77046
rect 71400 76982 71406 77014
rect 71470 77014 71471 77046
rect 73853 77046 73919 77047
rect 73853 77014 73854 77046
rect 71470 76982 71476 77014
rect 71400 76780 71476 76982
rect 71264 76704 71476 76780
rect 73848 76982 73854 77014
rect 73918 77014 73919 77046
rect 76437 77046 76503 77047
rect 76437 77014 76438 77046
rect 73918 76982 73924 77014
rect 71128 76638 71204 76644
rect 71128 76574 71134 76638
rect 71198 76574 71204 76638
rect 71128 75958 71204 76574
rect 71128 75926 71134 75958
rect 71133 75894 71134 75926
rect 71198 75926 71204 75958
rect 71198 75894 71199 75926
rect 71133 75893 71199 75894
rect 68952 75214 68958 75278
rect 69022 75214 69028 75278
rect 68952 75208 69028 75214
rect 71264 75278 71340 76704
rect 71400 76638 71476 76644
rect 71400 76574 71406 76638
rect 71470 76574 71476 76638
rect 71400 75958 71476 76574
rect 71400 75926 71406 75958
rect 71405 75894 71406 75926
rect 71470 75926 71476 75958
rect 73712 76638 73788 76644
rect 73712 76574 73718 76638
rect 73782 76574 73788 76638
rect 73712 75958 73788 76574
rect 73712 75926 73718 75958
rect 71470 75894 71471 75926
rect 71405 75893 71471 75894
rect 73717 75894 73718 75926
rect 73782 75926 73788 75958
rect 73782 75894 73783 75926
rect 73717 75893 73783 75894
rect 71264 75214 71270 75278
rect 71334 75214 71340 75278
rect 71264 75208 71340 75214
rect 73848 75278 73924 76982
rect 76432 76982 76438 77014
rect 76502 77014 76503 77046
rect 78885 77046 78951 77047
rect 78885 77014 78886 77046
rect 76502 76982 76508 77014
rect 76160 76638 76236 76644
rect 76160 76574 76166 76638
rect 76230 76574 76236 76638
rect 76160 75958 76236 76574
rect 76160 75926 76166 75958
rect 76165 75894 76166 75926
rect 76230 75926 76236 75958
rect 76230 75894 76231 75926
rect 76165 75893 76231 75894
rect 73848 75214 73854 75278
rect 73918 75214 73924 75278
rect 73848 75208 73924 75214
rect 76432 75278 76508 76982
rect 78880 76982 78886 77014
rect 78950 77014 78951 77046
rect 81469 77046 81535 77047
rect 81469 77014 81470 77046
rect 78950 76982 78956 77014
rect 78613 76638 78679 76639
rect 78613 76606 78614 76638
rect 78608 76574 78614 76606
rect 78678 76606 78679 76638
rect 78744 76638 78820 76644
rect 78678 76574 78684 76606
rect 78608 75958 78684 76574
rect 78608 75894 78614 75958
rect 78678 75894 78684 75958
rect 78744 76574 78750 76638
rect 78814 76574 78820 76638
rect 78744 75958 78820 76574
rect 78744 75926 78750 75958
rect 78608 75888 78684 75894
rect 78749 75894 78750 75926
rect 78814 75926 78820 75958
rect 78814 75894 78815 75926
rect 78749 75893 78815 75894
rect 76432 75214 76438 75278
rect 76502 75214 76508 75278
rect 76432 75208 76508 75214
rect 78880 75278 78956 76982
rect 81464 76982 81470 77014
rect 81534 77014 81535 77046
rect 83917 77046 83983 77047
rect 83917 77014 83918 77046
rect 81534 76982 81540 77014
rect 81328 76638 81404 76644
rect 81328 76574 81334 76638
rect 81398 76574 81404 76638
rect 81328 75958 81404 76574
rect 81328 75926 81334 75958
rect 81333 75894 81334 75926
rect 81398 75926 81404 75958
rect 81398 75894 81399 75926
rect 81333 75893 81399 75894
rect 78880 75214 78886 75278
rect 78950 75214 78956 75278
rect 78880 75208 78956 75214
rect 81464 75278 81540 76982
rect 83912 76982 83918 77014
rect 83982 77014 83983 77046
rect 86365 77046 86431 77047
rect 86365 77014 86366 77046
rect 83982 76982 83988 77014
rect 83776 76638 83852 76644
rect 83776 76574 83782 76638
rect 83846 76574 83852 76638
rect 83776 75958 83852 76574
rect 83776 75926 83782 75958
rect 83781 75894 83782 75926
rect 83846 75926 83852 75958
rect 83846 75894 83847 75926
rect 83781 75893 83847 75894
rect 81464 75214 81470 75278
rect 81534 75214 81540 75278
rect 81464 75208 81540 75214
rect 83912 75278 83988 76982
rect 86360 76982 86366 77014
rect 86430 77014 86431 77046
rect 88949 77046 89015 77047
rect 88949 77014 88950 77046
rect 86430 76982 86436 77014
rect 86360 76780 86436 76982
rect 83912 75214 83918 75278
rect 83982 75214 83988 75278
rect 83912 75208 83988 75214
rect 86224 76704 86436 76780
rect 88944 76982 88950 77014
rect 89014 77014 89015 77046
rect 89014 76982 89020 77014
rect 86224 75278 86300 76704
rect 86360 76638 86436 76644
rect 86360 76574 86366 76638
rect 86430 76574 86436 76638
rect 86360 75958 86436 76574
rect 86360 75926 86366 75958
rect 86365 75894 86366 75926
rect 86430 75926 86436 75958
rect 88536 76638 88612 76644
rect 88536 76574 88542 76638
rect 88606 76574 88612 76638
rect 88536 75958 88612 76574
rect 88536 75926 88542 75958
rect 86430 75894 86431 75926
rect 86365 75893 86431 75894
rect 88541 75894 88542 75926
rect 88606 75926 88612 75958
rect 88808 76638 88884 76644
rect 88808 76574 88814 76638
rect 88878 76574 88884 76638
rect 88808 75958 88884 76574
rect 88808 75926 88814 75958
rect 88606 75894 88607 75926
rect 88541 75893 88607 75894
rect 88813 75894 88814 75926
rect 88878 75926 88884 75958
rect 88878 75894 88879 75926
rect 88813 75893 88879 75894
rect 86224 75214 86230 75278
rect 86294 75214 86300 75278
rect 86224 75208 86300 75214
rect 88944 75278 89020 76982
rect 88944 75214 88950 75278
rect 89014 75214 89020 75278
rect 88944 75208 89020 75214
rect 91256 75278 91332 77118
rect 93573 77118 93574 77150
rect 93638 77150 93644 77182
rect 96016 77182 96092 83308
rect 96288 82078 96364 82084
rect 96288 82014 96294 82078
rect 96358 82014 96364 82078
rect 96288 81534 96364 82014
rect 96288 81502 96294 81534
rect 96293 81470 96294 81502
rect 96358 81502 96364 81534
rect 97920 82078 97996 82084
rect 97920 82014 97926 82078
rect 97990 82014 97996 82078
rect 97920 81534 97996 82014
rect 97920 81502 97926 81534
rect 96358 81470 96359 81502
rect 96293 81469 96359 81470
rect 97925 81470 97926 81502
rect 97990 81502 97996 81534
rect 97990 81470 97991 81502
rect 97925 81469 97991 81470
rect 96016 77150 96022 77182
rect 93638 77118 93639 77150
rect 93573 77117 93639 77118
rect 96021 77118 96022 77150
rect 96086 77150 96092 77182
rect 98464 77182 98540 83308
rect 99688 82078 99764 82084
rect 99688 82014 99694 82078
rect 99758 82014 99764 82078
rect 99688 81534 99764 82014
rect 99688 81502 99694 81534
rect 99693 81470 99694 81502
rect 99758 81502 99764 81534
rect 99758 81470 99759 81502
rect 99693 81469 99759 81470
rect 98464 77150 98470 77182
rect 96086 77118 96087 77150
rect 96021 77117 96087 77118
rect 98469 77118 98470 77150
rect 98534 77150 98540 77182
rect 101048 77182 101124 83308
rect 101320 82078 101396 82084
rect 101320 82014 101326 82078
rect 101390 82014 101396 82078
rect 101320 81534 101396 82014
rect 101320 81502 101326 81534
rect 101325 81470 101326 81502
rect 101390 81502 101396 81534
rect 102952 82078 103028 82084
rect 102952 82014 102958 82078
rect 103022 82014 103028 82078
rect 102952 81534 103028 82014
rect 102952 81502 102958 81534
rect 101390 81470 101391 81502
rect 101325 81469 101391 81470
rect 102957 81470 102958 81502
rect 103022 81502 103028 81534
rect 103022 81470 103023 81502
rect 102957 81469 103023 81470
rect 101048 77150 101054 77182
rect 98534 77118 98535 77150
rect 98469 77117 98535 77118
rect 101053 77118 101054 77150
rect 101118 77150 101124 77182
rect 103360 77182 103436 83308
rect 104584 82078 104660 82084
rect 104584 82014 104590 82078
rect 104654 82014 104660 82078
rect 104584 81534 104660 82014
rect 104584 81502 104590 81534
rect 104589 81470 104590 81502
rect 104654 81502 104660 81534
rect 104654 81470 104655 81502
rect 104589 81469 104655 81470
rect 103360 77150 103366 77182
rect 101118 77118 101119 77150
rect 101053 77117 101119 77118
rect 103365 77118 103366 77150
rect 103430 77150 103436 77182
rect 103909 77182 103975 77183
rect 103909 77150 103910 77182
rect 103430 77118 103431 77150
rect 103365 77117 103431 77118
rect 103904 77118 103910 77150
rect 103974 77150 103975 77182
rect 106080 77182 106156 83308
rect 118048 82758 118124 82764
rect 118048 82694 118054 82758
rect 118118 82694 118124 82758
rect 106352 82078 106428 82084
rect 106352 82014 106358 82078
rect 106422 82014 106428 82078
rect 106352 81534 106428 82014
rect 106352 81502 106358 81534
rect 106357 81470 106358 81502
rect 106422 81502 106428 81534
rect 107848 82078 107924 82084
rect 107848 82014 107854 82078
rect 107918 82014 107924 82078
rect 107848 81534 107924 82014
rect 107848 81502 107854 81534
rect 106422 81470 106423 81502
rect 106357 81469 106423 81470
rect 107853 81470 107854 81502
rect 107918 81502 107924 81534
rect 109616 82078 109692 82084
rect 109616 82014 109622 82078
rect 109686 82014 109692 82078
rect 109616 81534 109692 82014
rect 109616 81502 109622 81534
rect 107918 81470 107919 81502
rect 107853 81469 107919 81470
rect 109621 81470 109622 81502
rect 109686 81502 109692 81534
rect 111384 82078 111460 82084
rect 111384 82014 111390 82078
rect 111454 82014 111460 82078
rect 111384 81534 111460 82014
rect 111384 81502 111390 81534
rect 109686 81470 109687 81502
rect 109621 81469 109687 81470
rect 111389 81470 111390 81502
rect 111454 81502 111460 81534
rect 112880 82078 112956 82084
rect 112880 82014 112886 82078
rect 112950 82014 112956 82078
rect 112880 81534 112956 82014
rect 112880 81502 112886 81534
rect 111454 81470 111455 81502
rect 111389 81469 111455 81470
rect 112885 81470 112886 81502
rect 112950 81502 112956 81534
rect 114648 82078 114724 82084
rect 114648 82014 114654 82078
rect 114718 82014 114724 82078
rect 114648 81534 114724 82014
rect 114648 81502 114654 81534
rect 112950 81470 112951 81502
rect 112885 81469 112951 81470
rect 114653 81470 114654 81502
rect 114718 81502 114724 81534
rect 116416 82078 116492 82084
rect 116416 82014 116422 82078
rect 116486 82014 116492 82078
rect 116416 81534 116492 82014
rect 116416 81502 116422 81534
rect 114718 81470 114719 81502
rect 114653 81469 114719 81470
rect 116421 81470 116422 81502
rect 116486 81502 116492 81534
rect 117912 82078 117988 82084
rect 117912 82014 117918 82078
rect 117982 82014 117988 82078
rect 117912 81534 117988 82014
rect 117912 81502 117918 81534
rect 116486 81470 116487 81502
rect 116421 81469 116487 81470
rect 117917 81470 117918 81502
rect 117982 81502 117988 81534
rect 117982 81470 117983 81502
rect 117917 81469 117983 81470
rect 118048 80854 118124 82694
rect 118189 81398 118255 81399
rect 118189 81366 118190 81398
rect 118048 80822 118054 80854
rect 118053 80790 118054 80822
rect 118118 80822 118124 80854
rect 118184 81334 118190 81366
rect 118254 81366 118255 81398
rect 118254 81334 118260 81366
rect 118118 80790 118119 80822
rect 118053 80789 118119 80790
rect 117912 80718 117988 80724
rect 117912 80654 117918 80718
rect 117982 80654 117988 80718
rect 117912 78678 117988 80654
rect 118184 79494 118260 81334
rect 118456 80310 118532 83308
rect 119544 82078 119620 82084
rect 119544 82014 119550 82078
rect 119614 82014 119620 82078
rect 119544 81534 119620 82014
rect 119544 81502 119550 81534
rect 119549 81470 119550 81502
rect 119614 81502 119620 81534
rect 119614 81470 119615 81502
rect 119549 81469 119615 81470
rect 118456 80278 118462 80310
rect 118461 80246 118462 80278
rect 118526 80278 118532 80310
rect 119680 80310 119756 83308
rect 121448 82078 121524 82084
rect 121448 82014 121454 82078
rect 121518 82014 121524 82078
rect 121448 81534 121524 82014
rect 121448 81502 121454 81534
rect 121453 81470 121454 81502
rect 121518 81502 121524 81534
rect 123216 82078 123292 82084
rect 123216 82014 123222 82078
rect 123286 82014 123292 82078
rect 123216 81534 123292 82014
rect 123216 81502 123222 81534
rect 121518 81470 121519 81502
rect 121453 81469 121519 81470
rect 123221 81470 123222 81502
rect 123286 81502 123292 81534
rect 124712 82078 124788 82084
rect 124712 82014 124718 82078
rect 124782 82014 124788 82078
rect 124712 81534 124788 82014
rect 124712 81502 124718 81534
rect 123286 81470 123287 81502
rect 123221 81469 123287 81470
rect 124717 81470 124718 81502
rect 124782 81502 124788 81534
rect 126344 82078 126420 82084
rect 126344 82014 126350 82078
rect 126414 82014 126420 82078
rect 126344 81534 126420 82014
rect 126344 81502 126350 81534
rect 124782 81470 124783 81502
rect 124717 81469 124783 81470
rect 126349 81470 126350 81502
rect 126414 81502 126420 81534
rect 128112 82078 128188 82084
rect 128112 82014 128118 82078
rect 128182 82014 128188 82078
rect 128112 81534 128188 82014
rect 128112 81502 128118 81534
rect 126414 81470 126415 81502
rect 126349 81469 126415 81470
rect 128117 81470 128118 81502
rect 128182 81502 128188 81534
rect 129880 82078 129956 82084
rect 129880 82014 129886 82078
rect 129950 82014 129956 82078
rect 129880 81534 129956 82014
rect 129880 81502 129886 81534
rect 128182 81470 128183 81502
rect 128117 81469 128183 81470
rect 129885 81470 129886 81502
rect 129950 81502 129956 81534
rect 129950 81470 129951 81502
rect 129885 81469 129951 81470
rect 122944 81398 123020 81404
rect 122944 81334 122950 81398
rect 123014 81334 123020 81398
rect 122269 80718 122335 80719
rect 122269 80686 122270 80718
rect 119680 80278 119686 80310
rect 118526 80246 118527 80278
rect 118461 80245 118527 80246
rect 119685 80246 119686 80278
rect 119750 80278 119756 80310
rect 122264 80654 122270 80686
rect 122334 80686 122335 80718
rect 122334 80654 122340 80686
rect 119750 80246 119751 80278
rect 119685 80245 119751 80246
rect 122264 79902 122340 80654
rect 122264 79838 122270 79902
rect 122334 79838 122340 79902
rect 122264 79832 122340 79838
rect 122405 79766 122471 79767
rect 122405 79734 122406 79766
rect 118184 79430 118190 79494
rect 118254 79430 118260 79494
rect 118184 79424 118260 79430
rect 122400 79702 122406 79734
rect 122470 79734 122471 79766
rect 122470 79702 122476 79734
rect 117912 78646 117918 78678
rect 117917 78614 117918 78646
rect 117982 78646 117988 78678
rect 118048 79358 118124 79364
rect 118048 79294 118054 79358
rect 118118 79294 118124 79358
rect 117982 78614 117983 78646
rect 117917 78613 117983 78614
rect 116557 78542 116623 78543
rect 116557 78510 116558 78542
rect 116552 78478 116558 78510
rect 116622 78510 116623 78542
rect 116622 78478 116628 78510
rect 106080 77150 106086 77182
rect 103974 77118 103980 77150
rect 93845 77046 93911 77047
rect 93845 77014 93846 77046
rect 93840 76982 93846 77014
rect 93910 77014 93911 77046
rect 96293 77046 96359 77047
rect 96293 77014 96294 77046
rect 93910 76982 93916 77014
rect 93840 76780 93916 76982
rect 93704 76704 93916 76780
rect 96288 76982 96294 77014
rect 96358 77014 96359 77046
rect 98877 77046 98943 77047
rect 98877 77014 98878 77046
rect 96358 76982 96364 77014
rect 91392 76638 91468 76644
rect 91392 76574 91398 76638
rect 91462 76574 91468 76638
rect 93573 76638 93639 76639
rect 93573 76606 93574 76638
rect 91392 75958 91468 76574
rect 91392 75926 91398 75958
rect 91397 75894 91398 75926
rect 91462 75926 91468 75958
rect 93568 76574 93574 76606
rect 93638 76606 93639 76638
rect 93638 76574 93644 76606
rect 93568 75958 93644 76574
rect 91462 75894 91463 75926
rect 91397 75893 91463 75894
rect 93568 75894 93574 75958
rect 93638 75894 93644 75958
rect 93568 75888 93644 75894
rect 91256 75214 91262 75278
rect 91326 75214 91332 75278
rect 91256 75208 91332 75214
rect 93704 75278 93780 76704
rect 93840 76638 93916 76644
rect 93840 76574 93846 76638
rect 93910 76574 93916 76638
rect 93840 75958 93916 76574
rect 93840 75926 93846 75958
rect 93845 75894 93846 75926
rect 93910 75926 93916 75958
rect 96152 76638 96228 76644
rect 96152 76574 96158 76638
rect 96222 76574 96228 76638
rect 96152 75958 96228 76574
rect 96152 75926 96158 75958
rect 93910 75894 93911 75926
rect 93845 75893 93911 75894
rect 96157 75894 96158 75926
rect 96222 75926 96228 75958
rect 96222 75894 96223 75926
rect 96157 75893 96223 75894
rect 93704 75214 93710 75278
rect 93774 75214 93780 75278
rect 93704 75208 93780 75214
rect 96288 75278 96364 76982
rect 98872 76982 98878 77014
rect 98942 77014 98943 77046
rect 101325 77046 101391 77047
rect 101325 77014 101326 77046
rect 98942 76982 98948 77014
rect 98605 76638 98671 76639
rect 98605 76606 98606 76638
rect 98600 76574 98606 76606
rect 98670 76606 98671 76638
rect 98736 76638 98812 76644
rect 98670 76574 98676 76606
rect 98600 75958 98676 76574
rect 98600 75894 98606 75958
rect 98670 75894 98676 75958
rect 98736 76574 98742 76638
rect 98806 76574 98812 76638
rect 98736 75958 98812 76574
rect 98736 75926 98742 75958
rect 98600 75888 98676 75894
rect 98741 75894 98742 75926
rect 98806 75926 98812 75958
rect 98806 75894 98807 75926
rect 98741 75893 98807 75894
rect 96288 75214 96294 75278
rect 96358 75214 96364 75278
rect 96288 75208 96364 75214
rect 98872 75278 98948 76982
rect 101320 76982 101326 77014
rect 101390 77014 101391 77046
rect 101390 76982 101396 77014
rect 101184 76638 101260 76644
rect 101184 76574 101190 76638
rect 101254 76574 101260 76638
rect 101184 75958 101260 76574
rect 101184 75926 101190 75958
rect 101189 75894 101190 75926
rect 101254 75926 101260 75958
rect 101254 75894 101255 75926
rect 101189 75893 101255 75894
rect 98872 75214 98878 75278
rect 98942 75214 98948 75278
rect 98872 75208 98948 75214
rect 101320 75278 101396 76982
rect 103768 76638 103844 76644
rect 103768 76574 103774 76638
rect 103838 76574 103844 76638
rect 103768 75958 103844 76574
rect 103768 75926 103774 75958
rect 103773 75894 103774 75926
rect 103838 75926 103844 75958
rect 103838 75894 103839 75926
rect 103773 75893 103839 75894
rect 101320 75214 101326 75278
rect 101390 75214 101396 75278
rect 101320 75208 101396 75214
rect 103904 75278 103980 77118
rect 106085 77118 106086 77150
rect 106150 77150 106156 77182
rect 115333 77182 115399 77183
rect 115333 77150 115334 77182
rect 106150 77118 106151 77150
rect 106085 77117 106151 77118
rect 115328 77118 115334 77150
rect 115398 77150 115399 77182
rect 115398 77118 115404 77150
rect 106357 77046 106423 77047
rect 106357 77014 106358 77046
rect 106352 76982 106358 77014
rect 106422 77014 106423 77046
rect 106422 76982 106428 77014
rect 106216 76638 106292 76644
rect 106216 76574 106222 76638
rect 106286 76574 106292 76638
rect 106216 75958 106292 76574
rect 106216 75926 106222 75958
rect 106221 75894 106222 75926
rect 106286 75926 106292 75958
rect 106286 75894 106287 75926
rect 106221 75893 106287 75894
rect 103904 75214 103910 75278
rect 103974 75214 103980 75278
rect 103904 75208 103980 75214
rect 106352 75278 106428 76982
rect 106352 75214 106358 75278
rect 106422 75214 106428 75278
rect 106352 75208 106428 75214
rect 61477 75142 61543 75143
rect 61477 75110 61478 75142
rect 61472 75078 61478 75110
rect 61542 75110 61543 75142
rect 63925 75142 63991 75143
rect 63925 75110 63926 75142
rect 61542 75078 61548 75110
rect 61472 73238 61548 75078
rect 61472 73174 61478 73238
rect 61542 73174 61548 73238
rect 61472 73168 61548 73174
rect 63920 75078 63926 75110
rect 63990 75110 63991 75142
rect 66509 75142 66575 75143
rect 66509 75110 66510 75142
rect 63990 75078 63996 75110
rect 63920 73238 63996 75078
rect 63920 73174 63926 73238
rect 63990 73174 63996 73238
rect 63920 73168 63996 73174
rect 66504 75078 66510 75110
rect 66574 75110 66575 75142
rect 68957 75142 69023 75143
rect 68957 75110 68958 75142
rect 66574 75078 66580 75110
rect 66504 73238 66580 75078
rect 66504 73174 66510 73238
rect 66574 73174 66580 73238
rect 66504 73168 66580 73174
rect 68952 75078 68958 75110
rect 69022 75110 69023 75142
rect 71405 75142 71471 75143
rect 71405 75110 71406 75142
rect 69022 75078 69028 75110
rect 68952 73238 69028 75078
rect 68952 73174 68958 73238
rect 69022 73174 69028 73238
rect 68952 73168 69028 73174
rect 71400 75078 71406 75110
rect 71470 75110 71471 75142
rect 73989 75142 74055 75143
rect 73989 75110 73990 75142
rect 71470 75078 71476 75110
rect 71400 73238 71476 75078
rect 71400 73174 71406 73238
rect 71470 73174 71476 73238
rect 71400 73168 71476 73174
rect 73984 75078 73990 75110
rect 74054 75110 74055 75142
rect 76437 75142 76503 75143
rect 76437 75110 76438 75142
rect 74054 75078 74060 75110
rect 73984 73238 74060 75078
rect 73984 73174 73990 73238
rect 74054 73174 74060 73238
rect 73984 73168 74060 73174
rect 76432 75078 76438 75110
rect 76502 75110 76503 75142
rect 78885 75142 78951 75143
rect 78885 75110 78886 75142
rect 76502 75078 76508 75110
rect 76432 73238 76508 75078
rect 76432 73174 76438 73238
rect 76502 73174 76508 73238
rect 76432 73168 76508 73174
rect 78880 75078 78886 75110
rect 78950 75110 78951 75142
rect 81469 75142 81535 75143
rect 81469 75110 81470 75142
rect 78950 75078 78956 75110
rect 78880 73238 78956 75078
rect 78880 73174 78886 73238
rect 78950 73174 78956 73238
rect 78880 73168 78956 73174
rect 81464 75078 81470 75110
rect 81534 75110 81535 75142
rect 83917 75142 83983 75143
rect 83917 75110 83918 75142
rect 81534 75078 81540 75110
rect 81464 73238 81540 75078
rect 81464 73174 81470 73238
rect 81534 73174 81540 73238
rect 81464 73168 81540 73174
rect 83912 75078 83918 75110
rect 83982 75110 83983 75142
rect 86501 75142 86567 75143
rect 86501 75110 86502 75142
rect 83982 75078 83988 75110
rect 83912 73238 83988 75078
rect 83912 73174 83918 73238
rect 83982 73174 83988 73238
rect 83912 73168 83988 73174
rect 86496 75078 86502 75110
rect 86566 75110 86567 75142
rect 88949 75142 89015 75143
rect 88949 75110 88950 75142
rect 86566 75078 86572 75110
rect 86496 73238 86572 75078
rect 86496 73174 86502 73238
rect 86566 73174 86572 73238
rect 86496 73168 86572 73174
rect 88944 75078 88950 75110
rect 89014 75110 89015 75142
rect 91397 75142 91463 75143
rect 91397 75110 91398 75142
rect 89014 75078 89020 75110
rect 88944 73238 89020 75078
rect 88944 73174 88950 73238
rect 89014 73174 89020 73238
rect 88944 73168 89020 73174
rect 91392 75078 91398 75110
rect 91462 75110 91463 75142
rect 93704 75142 93780 75148
rect 91462 75078 91468 75110
rect 91392 73238 91468 75078
rect 91392 73174 91398 73238
rect 91462 73174 91468 73238
rect 93704 75078 93710 75142
rect 93774 75078 93780 75142
rect 96429 75142 96495 75143
rect 96429 75110 96430 75142
rect 93704 73238 93780 75078
rect 93704 73206 93710 73238
rect 91392 73168 91468 73174
rect 93709 73174 93710 73206
rect 93774 73206 93780 73238
rect 96424 75078 96430 75110
rect 96494 75110 96495 75142
rect 98877 75142 98943 75143
rect 98877 75110 98878 75142
rect 96494 75078 96500 75110
rect 96424 73238 96500 75078
rect 93774 73174 93775 73206
rect 93709 73173 93775 73174
rect 96424 73174 96430 73238
rect 96494 73174 96500 73238
rect 96424 73168 96500 73174
rect 98872 75078 98878 75110
rect 98942 75110 98943 75142
rect 101461 75142 101527 75143
rect 101461 75110 101462 75142
rect 98942 75078 98948 75110
rect 98872 73238 98948 75078
rect 98872 73174 98878 73238
rect 98942 73174 98948 73238
rect 98872 73168 98948 73174
rect 101456 75078 101462 75110
rect 101526 75110 101527 75142
rect 103909 75142 103975 75143
rect 103909 75110 103910 75142
rect 101526 75078 101532 75110
rect 101456 73238 101532 75078
rect 101456 73174 101462 73238
rect 101526 73174 101532 73238
rect 101456 73168 101532 73174
rect 103904 75078 103910 75110
rect 103974 75110 103975 75142
rect 106357 75142 106423 75143
rect 106357 75110 106358 75142
rect 103974 75078 103980 75110
rect 103904 73238 103980 75078
rect 103904 73174 103910 73238
rect 103974 73174 103980 73238
rect 103904 73168 103980 73174
rect 106352 75078 106358 75110
rect 106422 75110 106423 75142
rect 106422 75078 106428 75110
rect 106352 73238 106428 75078
rect 115328 74462 115404 77118
rect 116552 75958 116628 78478
rect 118048 77318 118124 79294
rect 122269 78406 122335 78407
rect 122269 78374 122270 78406
rect 118048 77286 118054 77318
rect 118053 77254 118054 77286
rect 118118 77286 118124 77318
rect 122264 78342 122270 78374
rect 122334 78374 122335 78406
rect 122334 78342 122340 78374
rect 118118 77254 118119 77286
rect 118053 77253 118119 77254
rect 116552 75894 116558 75958
rect 116622 75894 116628 75958
rect 116552 75888 116628 75894
rect 115469 75686 115535 75687
rect 115469 75654 115470 75686
rect 115328 74398 115334 74462
rect 115398 74398 115404 74462
rect 115328 74392 115404 74398
rect 115464 75622 115470 75654
rect 115534 75654 115535 75686
rect 122264 75686 122340 78342
rect 122400 77046 122476 79702
rect 122944 78542 123020 81334
rect 130832 79222 130908 83308
rect 136000 83030 136348 83036
rect 136000 82966 136006 83030
rect 136070 82966 136142 83030
rect 136206 82966 136278 83030
rect 136342 82966 136348 83030
rect 136000 82894 136348 82966
rect 136000 82830 136006 82894
rect 136070 82830 136142 82894
rect 136206 82830 136278 82894
rect 136342 82830 136348 82894
rect 136000 82758 136348 82830
rect 136000 82694 136006 82758
rect 136070 82694 136142 82758
rect 136206 82694 136278 82758
rect 136342 82694 136348 82758
rect 135320 82350 135668 82356
rect 135320 82286 135326 82350
rect 135390 82286 135462 82350
rect 135526 82286 135598 82350
rect 135662 82286 135668 82350
rect 135320 82214 135668 82286
rect 135320 82150 135326 82214
rect 135390 82150 135462 82214
rect 135526 82150 135598 82214
rect 135662 82150 135668 82214
rect 131376 82078 131452 82084
rect 131376 82014 131382 82078
rect 131446 82014 131452 82078
rect 131376 81534 131452 82014
rect 131376 81502 131382 81534
rect 131381 81470 131382 81502
rect 131446 81502 131452 81534
rect 133144 82078 133220 82084
rect 133144 82014 133150 82078
rect 133214 82014 133220 82078
rect 133144 81534 133220 82014
rect 133144 81502 133150 81534
rect 131446 81470 131447 81502
rect 131381 81469 131447 81470
rect 133149 81470 133150 81502
rect 133214 81502 133220 81534
rect 135320 82078 135668 82150
rect 135320 82014 135326 82078
rect 135390 82014 135462 82078
rect 135526 82014 135598 82078
rect 135662 82014 135668 82078
rect 133214 81470 133215 81502
rect 133149 81469 133215 81470
rect 130832 79190 130838 79222
rect 130837 79158 130838 79190
rect 130902 79190 130908 79222
rect 135320 80990 135668 82014
rect 135320 80926 135326 80990
rect 135390 80926 135668 80990
rect 135320 79494 135668 80926
rect 135320 79430 135326 79494
rect 135390 79430 135668 79494
rect 130902 79158 130903 79190
rect 130837 79157 130903 79158
rect 122944 78510 122950 78542
rect 122949 78478 122950 78510
rect 123014 78510 123020 78542
rect 123014 78478 123015 78510
rect 122949 78477 123015 78478
rect 134781 78406 134847 78407
rect 134781 78374 134782 78406
rect 134776 78342 134782 78374
rect 134846 78374 134847 78406
rect 134846 78342 134852 78374
rect 134776 77726 134852 78342
rect 134776 77662 134782 77726
rect 134846 77662 134852 77726
rect 134776 77656 134852 77662
rect 135320 77726 135668 79430
rect 135320 77662 135326 77726
rect 135390 77662 135668 77726
rect 122400 76982 122406 77046
rect 122470 76982 122476 77046
rect 122400 76976 122476 76982
rect 115534 75622 115540 75654
rect 106352 73174 106358 73238
rect 106422 73174 106428 73238
rect 106352 73168 106428 73174
rect 115328 74326 115404 74332
rect 115328 74262 115334 74326
rect 115398 74262 115404 74326
rect 109621 73102 109687 73103
rect 109621 73070 109622 73102
rect 59432 71542 59438 71606
rect 59502 71542 59508 71606
rect 59432 71536 59508 71542
rect 109616 73038 109622 73070
rect 109686 73070 109687 73102
rect 109686 73038 109692 73070
rect 29784 71470 29860 71476
rect 29784 71406 29790 71470
rect 29854 71406 29860 71470
rect 31285 71470 31351 71471
rect 31285 71438 31286 71470
rect 29784 71062 29860 71406
rect 29784 71030 29790 71062
rect 29789 70998 29790 71030
rect 29854 71030 29860 71062
rect 31280 71406 31286 71438
rect 31350 71438 31351 71470
rect 31960 71470 32036 71476
rect 31350 71406 31356 71438
rect 31280 71062 31356 71406
rect 29854 70998 29855 71030
rect 29789 70997 29855 70998
rect 31280 70998 31286 71062
rect 31350 70998 31356 71062
rect 31960 71406 31966 71470
rect 32030 71406 32036 71470
rect 32509 71470 32575 71471
rect 32509 71438 32510 71470
rect 31960 71062 32036 71406
rect 31960 71030 31966 71062
rect 31280 70992 31356 70998
rect 31965 70998 31966 71030
rect 32030 71030 32036 71062
rect 32504 71406 32510 71438
rect 32574 71438 32575 71470
rect 33733 71470 33799 71471
rect 33733 71438 33734 71470
rect 32574 71406 32580 71438
rect 32504 71062 32580 71406
rect 32030 70998 32031 71030
rect 31965 70997 32031 70998
rect 32504 70998 32510 71062
rect 32574 70998 32580 71062
rect 32504 70992 32580 70998
rect 33728 71406 33734 71438
rect 33798 71438 33799 71470
rect 34408 71470 34484 71476
rect 33798 71406 33804 71438
rect 33728 71062 33804 71406
rect 33728 70998 33734 71062
rect 33798 70998 33804 71062
rect 34408 71406 34414 71470
rect 34478 71406 34484 71470
rect 34957 71470 35023 71471
rect 34957 71438 34958 71470
rect 34408 71062 34484 71406
rect 34408 71030 34414 71062
rect 33728 70992 33804 70998
rect 34413 70998 34414 71030
rect 34478 71030 34484 71062
rect 34952 71406 34958 71438
rect 35022 71438 35023 71470
rect 35768 71470 35844 71476
rect 35022 71406 35028 71438
rect 34952 71062 35028 71406
rect 34478 70998 34479 71030
rect 34413 70997 34479 70998
rect 34952 70998 34958 71062
rect 35022 70998 35028 71062
rect 35768 71406 35774 71470
rect 35838 71406 35844 71470
rect 36181 71470 36247 71471
rect 36181 71438 36182 71470
rect 35768 71062 35844 71406
rect 35768 71030 35774 71062
rect 34952 70992 35028 70998
rect 35773 70998 35774 71030
rect 35838 71030 35844 71062
rect 36176 71406 36182 71438
rect 36246 71438 36247 71470
rect 36992 71470 37068 71476
rect 36246 71406 36252 71438
rect 36176 71062 36252 71406
rect 35838 70998 35839 71030
rect 35773 70997 35839 70998
rect 36176 70998 36182 71062
rect 36246 70998 36252 71062
rect 36992 71406 36998 71470
rect 37062 71406 37068 71470
rect 37541 71470 37607 71471
rect 37541 71438 37542 71470
rect 36992 71062 37068 71406
rect 36992 71030 36998 71062
rect 36176 70992 36252 70998
rect 36997 70998 36998 71030
rect 37062 71030 37068 71062
rect 37536 71406 37542 71438
rect 37606 71438 37607 71470
rect 38216 71470 38292 71476
rect 37606 71406 37612 71438
rect 37536 71062 37612 71406
rect 37062 70998 37063 71030
rect 36997 70997 37063 70998
rect 37536 70998 37542 71062
rect 37606 70998 37612 71062
rect 38216 71406 38222 71470
rect 38286 71406 38292 71470
rect 39989 71470 40055 71471
rect 39989 71438 39990 71470
rect 38216 71062 38292 71406
rect 38216 71030 38222 71062
rect 37536 70992 37612 70998
rect 38221 70998 38222 71030
rect 38286 71030 38292 71062
rect 39984 71406 39990 71438
rect 40054 71438 40055 71470
rect 40664 71470 40740 71476
rect 40054 71406 40060 71438
rect 39984 71062 40060 71406
rect 38286 70998 38287 71030
rect 38221 70997 38287 70998
rect 39984 70998 39990 71062
rect 40054 70998 40060 71062
rect 40664 71406 40670 71470
rect 40734 71406 40740 71470
rect 41213 71470 41279 71471
rect 41213 71438 41214 71470
rect 40664 71062 40740 71406
rect 40664 71030 40670 71062
rect 39984 70992 40060 70998
rect 40669 70998 40670 71030
rect 40734 71030 40740 71062
rect 41208 71406 41214 71438
rect 41278 71438 41279 71470
rect 41888 71470 41964 71476
rect 41278 71406 41284 71438
rect 41208 71062 41284 71406
rect 40734 70998 40735 71030
rect 40669 70997 40735 70998
rect 41208 70998 41214 71062
rect 41278 70998 41284 71062
rect 41888 71406 41894 71470
rect 41958 71406 41964 71470
rect 42437 71470 42503 71471
rect 42437 71438 42438 71470
rect 41888 71062 41964 71406
rect 41888 71030 41894 71062
rect 41208 70992 41284 70998
rect 41893 70998 41894 71030
rect 41958 71030 41964 71062
rect 42432 71406 42438 71438
rect 42502 71438 42503 71470
rect 43248 71470 43324 71476
rect 42502 71406 42508 71438
rect 42432 71062 42508 71406
rect 41958 70998 41959 71030
rect 41893 70997 41959 70998
rect 42432 70998 42438 71062
rect 42502 70998 42508 71062
rect 43248 71406 43254 71470
rect 43318 71406 43324 71470
rect 44613 71470 44679 71471
rect 44613 71438 44614 71470
rect 43248 71062 43324 71406
rect 43248 71030 43254 71062
rect 42432 70992 42508 70998
rect 43253 70998 43254 71030
rect 43318 71030 43324 71062
rect 44608 71406 44614 71438
rect 44678 71438 44679 71470
rect 45696 71470 45772 71476
rect 44678 71406 44684 71438
rect 43318 70998 43319 71030
rect 43253 70997 43319 70998
rect 44608 70926 44684 71406
rect 45696 71406 45702 71470
rect 45766 71406 45772 71470
rect 46245 71470 46311 71471
rect 46245 71438 46246 71470
rect 45696 71062 45772 71406
rect 45696 71030 45702 71062
rect 45701 70998 45702 71030
rect 45766 71030 45772 71062
rect 46240 71406 46246 71438
rect 46310 71438 46311 71470
rect 46920 71470 46996 71476
rect 46310 71406 46316 71438
rect 46240 71062 46316 71406
rect 45766 70998 45767 71030
rect 45701 70997 45767 70998
rect 46240 70998 46246 71062
rect 46310 70998 46316 71062
rect 46920 71406 46926 71470
rect 46990 71406 46996 71470
rect 48693 71470 48759 71471
rect 48693 71438 48694 71470
rect 46920 71062 46996 71406
rect 46920 71030 46926 71062
rect 46240 70992 46316 70998
rect 46925 70998 46926 71030
rect 46990 71030 46996 71062
rect 48688 71406 48694 71438
rect 48758 71438 48759 71470
rect 49917 71470 49983 71471
rect 49917 71438 49918 71470
rect 48758 71406 48764 71438
rect 48688 71062 48764 71406
rect 46990 70998 46991 71030
rect 46925 70997 46991 70998
rect 48688 70998 48694 71062
rect 48758 70998 48764 71062
rect 48688 70992 48764 70998
rect 49912 71406 49918 71438
rect 49982 71438 49983 71470
rect 50728 71470 50804 71476
rect 49982 71406 49988 71438
rect 49912 71062 49988 71406
rect 49912 70998 49918 71062
rect 49982 70998 49988 71062
rect 50728 71406 50734 71470
rect 50798 71406 50804 71470
rect 51277 71470 51343 71471
rect 51277 71438 51278 71470
rect 50728 71062 50804 71406
rect 50728 71030 50734 71062
rect 49912 70992 49988 70998
rect 50733 70998 50734 71030
rect 50798 71030 50804 71062
rect 51272 71406 51278 71438
rect 51342 71438 51343 71470
rect 52501 71470 52567 71471
rect 52501 71438 52502 71470
rect 51342 71406 51348 71438
rect 51272 71062 51348 71406
rect 50798 70998 50799 71030
rect 50733 70997 50799 70998
rect 51272 70998 51278 71062
rect 51342 70998 51348 71062
rect 51272 70992 51348 70998
rect 52496 71406 52502 71438
rect 52566 71438 52567 71470
rect 53176 71470 53252 71476
rect 52566 71406 52572 71438
rect 52496 71062 52572 71406
rect 52496 70998 52502 71062
rect 52566 70998 52572 71062
rect 53176 71406 53182 71470
rect 53246 71406 53252 71470
rect 53317 71470 53383 71471
rect 53317 71438 53318 71470
rect 53176 71062 53252 71406
rect 53176 71030 53182 71062
rect 52496 70992 52572 70998
rect 53181 70998 53182 71030
rect 53246 71030 53252 71062
rect 53312 71406 53318 71438
rect 53382 71438 53383 71470
rect 54400 71470 54476 71476
rect 53382 71406 53388 71438
rect 53312 71062 53388 71406
rect 53246 70998 53247 71030
rect 53181 70997 53247 70998
rect 53312 70998 53318 71062
rect 53382 70998 53388 71062
rect 54400 71406 54406 71470
rect 54470 71406 54476 71470
rect 54949 71470 55015 71471
rect 54949 71438 54950 71470
rect 54400 71062 54476 71406
rect 54400 71030 54406 71062
rect 53312 70992 53388 70998
rect 54405 70998 54406 71030
rect 54470 71030 54476 71062
rect 54944 71406 54950 71438
rect 55014 71438 55015 71470
rect 56032 71470 56108 71476
rect 55014 71406 55020 71438
rect 54944 71062 55020 71406
rect 54470 70998 54471 71030
rect 54405 70997 54471 70998
rect 54944 70998 54950 71062
rect 55014 70998 55020 71062
rect 56032 71406 56038 71470
rect 56102 71406 56108 71470
rect 57397 71470 57463 71471
rect 57397 71438 57398 71470
rect 56032 71062 56108 71406
rect 56032 71030 56038 71062
rect 54944 70992 55020 70998
rect 56037 70998 56038 71030
rect 56102 71030 56108 71062
rect 57392 71406 57398 71438
rect 57462 71438 57463 71470
rect 58621 71470 58687 71471
rect 58621 71438 58622 71470
rect 57462 71406 57468 71438
rect 57392 71062 57468 71406
rect 56102 70998 56103 71030
rect 56037 70997 56103 70998
rect 57392 70998 57398 71062
rect 57462 70998 57468 71062
rect 57392 70992 57468 70998
rect 58616 71406 58622 71438
rect 58686 71438 58687 71470
rect 59432 71470 59508 71476
rect 58686 71406 58692 71438
rect 58616 71062 58692 71406
rect 58616 70998 58622 71062
rect 58686 70998 58692 71062
rect 59432 71406 59438 71470
rect 59502 71406 59508 71470
rect 59981 71470 60047 71471
rect 59981 71438 59982 71470
rect 59432 71062 59508 71406
rect 59432 71030 59438 71062
rect 58616 70992 58692 70998
rect 59437 70998 59438 71030
rect 59502 71030 59508 71062
rect 59976 71406 59982 71438
rect 60046 71438 60047 71470
rect 61205 71470 61271 71471
rect 61205 71438 61206 71470
rect 60046 71406 60052 71438
rect 59976 71062 60052 71406
rect 59502 70998 59503 71030
rect 59437 70997 59503 70998
rect 59976 70998 59982 71062
rect 60046 70998 60052 71062
rect 59976 70992 60052 70998
rect 61200 71406 61206 71438
rect 61270 71438 61271 71470
rect 61880 71470 61956 71476
rect 61270 71406 61276 71438
rect 61200 71062 61276 71406
rect 61200 70998 61206 71062
rect 61270 70998 61276 71062
rect 61880 71406 61886 71470
rect 61950 71406 61956 71470
rect 62429 71470 62495 71471
rect 62429 71438 62430 71470
rect 61880 71062 61956 71406
rect 61880 71030 61886 71062
rect 61200 70992 61276 70998
rect 61885 70998 61886 71030
rect 61950 71030 61956 71062
rect 62424 71406 62430 71438
rect 62494 71438 62495 71470
rect 63104 71470 63180 71476
rect 62494 71406 62500 71438
rect 62424 71062 62500 71406
rect 61950 70998 61951 71030
rect 61885 70997 61951 70998
rect 62424 70998 62430 71062
rect 62494 70998 62500 71062
rect 63104 71406 63110 71470
rect 63174 71406 63180 71470
rect 63653 71470 63719 71471
rect 63653 71438 63654 71470
rect 63104 71062 63180 71406
rect 63104 71030 63110 71062
rect 62424 70992 62500 70998
rect 63109 70998 63110 71030
rect 63174 71030 63180 71062
rect 63648 71406 63654 71438
rect 63718 71438 63719 71470
rect 65013 71470 65079 71471
rect 65013 71438 65014 71470
rect 63718 71406 63724 71438
rect 63648 71062 63724 71406
rect 63174 70998 63175 71030
rect 63109 70997 63175 70998
rect 63648 70998 63654 71062
rect 63718 70998 63724 71062
rect 63648 70992 63724 70998
rect 65008 71406 65014 71438
rect 65078 71438 65079 71470
rect 66101 71470 66167 71471
rect 66101 71438 66102 71470
rect 65078 71406 65084 71438
rect 65008 71062 65084 71406
rect 65008 70998 65014 71062
rect 65078 70998 65084 71062
rect 65008 70992 65084 70998
rect 66096 71406 66102 71438
rect 66166 71438 66167 71470
rect 66912 71470 66988 71476
rect 66166 71406 66172 71438
rect 66096 71062 66172 71406
rect 66096 70998 66102 71062
rect 66166 70998 66172 71062
rect 66912 71406 66918 71470
rect 66982 71406 66988 71470
rect 67461 71470 67527 71471
rect 67461 71438 67462 71470
rect 66912 71062 66988 71406
rect 66912 71030 66918 71062
rect 66096 70992 66172 70998
rect 66917 70998 66918 71030
rect 66982 71030 66988 71062
rect 67456 71406 67462 71438
rect 67526 71438 67527 71470
rect 68136 71470 68212 71476
rect 67526 71406 67532 71438
rect 67456 71062 67532 71406
rect 66982 70998 66983 71030
rect 66917 70997 66983 70998
rect 67456 70998 67462 71062
rect 67526 70998 67532 71062
rect 68136 71406 68142 71470
rect 68206 71406 68212 71470
rect 68685 71470 68751 71471
rect 68685 71438 68686 71470
rect 68136 71062 68212 71406
rect 68136 71030 68142 71062
rect 67456 70992 67532 70998
rect 68141 70998 68142 71030
rect 68206 71030 68212 71062
rect 68680 71406 68686 71438
rect 68750 71438 68751 71470
rect 69909 71470 69975 71471
rect 69909 71438 69910 71470
rect 68750 71406 68756 71438
rect 68680 71062 68756 71406
rect 68206 70998 68207 71030
rect 68141 70997 68207 70998
rect 68680 70998 68686 71062
rect 68750 70998 68756 71062
rect 68680 70992 68756 70998
rect 69904 71406 69910 71438
rect 69974 71438 69975 71470
rect 70584 71470 70660 71476
rect 69974 71406 69980 71438
rect 69904 71062 69980 71406
rect 69904 70998 69910 71062
rect 69974 70998 69980 71062
rect 70584 71406 70590 71470
rect 70654 71406 70660 71470
rect 72085 71470 72151 71471
rect 72085 71438 72086 71470
rect 70584 71062 70660 71406
rect 70584 71030 70590 71062
rect 69904 70992 69980 70998
rect 70589 70998 70590 71030
rect 70654 71030 70660 71062
rect 72080 71406 72086 71438
rect 72150 71438 72151 71470
rect 72216 71470 72292 71476
rect 72150 71406 72156 71438
rect 70654 70998 70655 71030
rect 70589 70997 70655 70998
rect 44608 70862 44614 70926
rect 44678 70862 44684 70926
rect 44608 70856 44684 70862
rect 72080 70926 72156 71406
rect 72216 71406 72222 71470
rect 72286 71406 72292 71470
rect 73717 71470 73783 71471
rect 73717 71438 73718 71470
rect 72216 71062 72292 71406
rect 72216 71030 72222 71062
rect 72221 70998 72222 71030
rect 72286 71030 72292 71062
rect 73712 71406 73718 71438
rect 73782 71438 73783 71470
rect 74392 71470 74468 71476
rect 73782 71406 73788 71438
rect 73712 71062 73788 71406
rect 72286 70998 72287 71030
rect 72221 70997 72287 70998
rect 73712 70998 73718 71062
rect 73782 70998 73788 71062
rect 74392 71406 74398 71470
rect 74462 71406 74468 71470
rect 74941 71470 75007 71471
rect 74941 71438 74942 71470
rect 74392 71062 74468 71406
rect 74392 71030 74398 71062
rect 73712 70992 73788 70998
rect 74397 70998 74398 71030
rect 74462 71030 74468 71062
rect 74936 71406 74942 71438
rect 75006 71438 75007 71470
rect 75616 71470 75692 71476
rect 75006 71406 75012 71438
rect 74936 71062 75012 71406
rect 74462 70998 74463 71030
rect 74397 70997 74463 70998
rect 74936 70998 74942 71062
rect 75006 70998 75012 71062
rect 75616 71406 75622 71470
rect 75686 71406 75692 71470
rect 76165 71470 76231 71471
rect 76165 71438 76166 71470
rect 75616 71062 75692 71406
rect 75616 71030 75622 71062
rect 74936 70992 75012 70998
rect 75621 70998 75622 71030
rect 75686 71030 75692 71062
rect 76160 71406 76166 71438
rect 76230 71438 76231 71470
rect 76840 71470 76916 71476
rect 76230 71406 76236 71438
rect 76160 71062 76236 71406
rect 75686 70998 75687 71030
rect 75621 70997 75687 70998
rect 76160 70998 76166 71062
rect 76230 70998 76236 71062
rect 76840 71406 76846 71470
rect 76910 71406 76916 71470
rect 77389 71470 77455 71471
rect 77389 71438 77390 71470
rect 76840 71062 76916 71406
rect 76840 71030 76846 71062
rect 76160 70992 76236 70998
rect 76845 70998 76846 71030
rect 76910 71030 76916 71062
rect 77384 71406 77390 71438
rect 77454 71438 77455 71470
rect 78200 71470 78276 71476
rect 77454 71406 77460 71438
rect 77384 71062 77460 71406
rect 76910 70998 76911 71030
rect 76845 70997 76911 70998
rect 77384 70998 77390 71062
rect 77454 70998 77460 71062
rect 78200 71406 78206 71470
rect 78270 71406 78276 71470
rect 78200 71062 78276 71406
rect 78200 71030 78206 71062
rect 77384 70992 77460 70998
rect 78205 70998 78206 71030
rect 78270 71030 78276 71062
rect 78472 71470 78548 71476
rect 78472 71406 78478 71470
rect 78542 71406 78548 71470
rect 78472 71062 78548 71406
rect 78472 71030 78478 71062
rect 78270 70998 78271 71030
rect 78205 70997 78271 70998
rect 78477 70998 78478 71030
rect 78542 71030 78548 71062
rect 79424 71470 79500 71476
rect 79424 71406 79430 71470
rect 79494 71406 79500 71470
rect 79973 71470 80039 71471
rect 79973 71438 79974 71470
rect 79424 71062 79500 71406
rect 79424 71030 79430 71062
rect 78542 70998 78543 71030
rect 78477 70997 78543 70998
rect 79429 70998 79430 71030
rect 79494 71030 79500 71062
rect 79968 71406 79974 71438
rect 80038 71438 80039 71470
rect 80648 71470 80724 71476
rect 80038 71406 80044 71438
rect 79968 71062 80044 71406
rect 79494 70998 79495 71030
rect 79429 70997 79495 70998
rect 79968 70998 79974 71062
rect 80038 70998 80044 71062
rect 80648 71406 80654 71470
rect 80718 71406 80724 71470
rect 80648 71062 80724 71406
rect 80648 71030 80654 71062
rect 79968 70992 80044 70998
rect 80653 70998 80654 71030
rect 80718 71030 80724 71062
rect 81872 71470 81948 71476
rect 81872 71406 81878 71470
rect 81942 71406 81948 71470
rect 82421 71470 82487 71471
rect 82421 71438 82422 71470
rect 81872 71062 81948 71406
rect 81872 71030 81878 71062
rect 80718 70998 80719 71030
rect 80653 70997 80719 70998
rect 81877 70998 81878 71030
rect 81942 71030 81948 71062
rect 82416 71406 82422 71438
rect 82486 71438 82487 71470
rect 83096 71470 83172 71476
rect 82486 71406 82492 71438
rect 82416 71062 82492 71406
rect 81942 70998 81943 71030
rect 81877 70997 81943 70998
rect 82416 70998 82422 71062
rect 82486 70998 82492 71062
rect 83096 71406 83102 71470
rect 83166 71406 83172 71470
rect 83645 71470 83711 71471
rect 83645 71438 83646 71470
rect 83096 71062 83172 71406
rect 83096 71030 83102 71062
rect 82416 70992 82492 70998
rect 83101 70998 83102 71030
rect 83166 71030 83172 71062
rect 83640 71406 83646 71438
rect 83710 71438 83711 71470
rect 84597 71470 84663 71471
rect 84597 71438 84598 71470
rect 83710 71406 83716 71438
rect 83640 71062 83716 71406
rect 83166 70998 83167 71030
rect 83101 70997 83167 70998
rect 83640 70998 83646 71062
rect 83710 70998 83716 71062
rect 83640 70992 83716 70998
rect 84592 71406 84598 71438
rect 84662 71438 84663 71470
rect 86093 71470 86159 71471
rect 86093 71438 86094 71470
rect 84662 71406 84668 71438
rect 84592 71062 84668 71406
rect 84592 70998 84598 71062
rect 84662 70998 84668 71062
rect 84592 70992 84668 70998
rect 86088 71406 86094 71438
rect 86158 71438 86159 71470
rect 86904 71470 86980 71476
rect 86158 71406 86164 71438
rect 86088 71062 86164 71406
rect 86088 70998 86094 71062
rect 86158 70998 86164 71062
rect 86904 71406 86910 71470
rect 86974 71406 86980 71470
rect 86904 71062 86980 71406
rect 86904 71030 86910 71062
rect 86088 70992 86164 70998
rect 86909 70998 86910 71030
rect 86974 71030 86980 71062
rect 88128 71470 88204 71476
rect 88128 71406 88134 71470
rect 88198 71406 88204 71470
rect 88677 71470 88743 71471
rect 88677 71438 88678 71470
rect 88128 71062 88204 71406
rect 88128 71030 88134 71062
rect 86974 70998 86975 71030
rect 86909 70997 86975 70998
rect 88133 70998 88134 71030
rect 88198 71030 88204 71062
rect 88672 71406 88678 71438
rect 88742 71438 88743 71470
rect 89352 71470 89428 71476
rect 88742 71406 88748 71438
rect 88672 71062 88748 71406
rect 88198 70998 88199 71030
rect 88133 70997 88199 70998
rect 88672 70998 88678 71062
rect 88742 70998 88748 71062
rect 89352 71406 89358 71470
rect 89422 71406 89428 71470
rect 89901 71470 89967 71471
rect 89901 71438 89902 71470
rect 89352 71062 89428 71406
rect 89352 71030 89358 71062
rect 88672 70992 88748 70998
rect 89357 70998 89358 71030
rect 89422 71030 89428 71062
rect 89896 71406 89902 71438
rect 89966 71438 89967 71470
rect 90712 71470 90788 71476
rect 89966 71406 89972 71438
rect 89896 71062 89972 71406
rect 89422 70998 89423 71030
rect 89357 70997 89423 70998
rect 89896 70998 89902 71062
rect 89966 70998 89972 71062
rect 90712 71406 90718 71470
rect 90782 71406 90788 71470
rect 91125 71470 91191 71471
rect 91125 71438 91126 71470
rect 90712 71062 90788 71406
rect 90712 71030 90718 71062
rect 89896 70992 89972 70998
rect 90717 70998 90718 71030
rect 90782 71030 90788 71062
rect 91120 71406 91126 71438
rect 91190 71438 91191 71470
rect 92349 71470 92415 71471
rect 92349 71438 92350 71470
rect 91190 71406 91196 71438
rect 91120 71062 91196 71406
rect 90782 70998 90783 71030
rect 90717 70997 90783 70998
rect 91120 70998 91126 71062
rect 91190 70998 91196 71062
rect 91120 70992 91196 70998
rect 92344 71406 92350 71438
rect 92414 71438 92415 71470
rect 93301 71470 93367 71471
rect 93301 71438 93302 71470
rect 92414 71406 92420 71438
rect 92344 71062 92420 71406
rect 92344 70998 92350 71062
rect 92414 70998 92420 71062
rect 92344 70992 92420 70998
rect 93296 71406 93302 71438
rect 93366 71438 93367 71470
rect 94933 71470 94999 71471
rect 94933 71438 94934 71470
rect 93366 71406 93372 71438
rect 72080 70862 72086 70926
rect 72150 70862 72156 70926
rect 72080 70856 72156 70862
rect 93296 70926 93372 71406
rect 94928 71406 94934 71438
rect 94998 71438 94999 71470
rect 95608 71470 95684 71476
rect 94998 71406 95004 71438
rect 94928 71062 95004 71406
rect 94928 70998 94934 71062
rect 94998 70998 95004 71062
rect 95608 71406 95614 71470
rect 95678 71406 95684 71470
rect 95608 71062 95684 71406
rect 95608 71030 95614 71062
rect 94928 70992 95004 70998
rect 95613 70998 95614 71030
rect 95678 71030 95684 71062
rect 96832 71470 96908 71476
rect 96832 71406 96838 71470
rect 96902 71406 96908 71470
rect 97381 71470 97447 71471
rect 97381 71438 97382 71470
rect 96832 71062 96908 71406
rect 96832 71030 96838 71062
rect 95678 70998 95679 71030
rect 95613 70997 95679 70998
rect 96837 70998 96838 71030
rect 96902 71030 96908 71062
rect 97376 71406 97382 71438
rect 97446 71438 97447 71470
rect 99829 71470 99895 71471
rect 99829 71438 99830 71470
rect 97446 71406 97452 71438
rect 97376 71062 97452 71406
rect 99824 71406 99830 71438
rect 99894 71438 99895 71470
rect 100912 71470 100988 71476
rect 99894 71406 99900 71438
rect 98605 71334 98671 71335
rect 98605 71302 98606 71334
rect 96902 70998 96903 71030
rect 96837 70997 96903 70998
rect 97376 70998 97382 71062
rect 97446 70998 97452 71062
rect 97376 70992 97452 70998
rect 98600 71270 98606 71302
rect 98670 71302 98671 71334
rect 98670 71270 98676 71302
rect 98600 71062 98676 71270
rect 98600 70998 98606 71062
rect 98670 70998 98676 71062
rect 98600 70992 98676 70998
rect 99824 71062 99900 71406
rect 99824 70998 99830 71062
rect 99894 70998 99900 71062
rect 100912 71406 100918 71470
rect 100982 71406 100988 71470
rect 100912 71062 100988 71406
rect 100912 71030 100918 71062
rect 99824 70992 99900 70998
rect 100917 70998 100918 71030
rect 100982 71030 100988 71062
rect 101864 71470 101940 71476
rect 101864 71406 101870 71470
rect 101934 71406 101940 71470
rect 102413 71470 102479 71471
rect 102413 71438 102414 71470
rect 101864 71062 101940 71406
rect 101864 71030 101870 71062
rect 100982 70998 100983 71030
rect 100917 70997 100983 70998
rect 101869 70998 101870 71030
rect 101934 71030 101940 71062
rect 102408 71406 102414 71438
rect 102478 71438 102479 71470
rect 103088 71470 103164 71476
rect 102478 71406 102484 71438
rect 102408 71062 102484 71406
rect 101934 70998 101935 71030
rect 101869 70997 101935 70998
rect 102408 70998 102414 71062
rect 102478 70998 102484 71062
rect 103088 71406 103094 71470
rect 103158 71406 103164 71470
rect 103637 71470 103703 71471
rect 103637 71438 103638 71470
rect 103088 71062 103164 71406
rect 103088 71030 103094 71062
rect 102408 70992 102484 70998
rect 103093 70998 103094 71030
rect 103158 71030 103164 71062
rect 103632 71406 103638 71438
rect 103702 71438 103703 71470
rect 104312 71470 104388 71476
rect 103702 71406 103708 71438
rect 103632 71062 103708 71406
rect 103158 70998 103159 71030
rect 103093 70997 103159 70998
rect 103632 70998 103638 71062
rect 103702 70998 103708 71062
rect 104312 71406 104318 71470
rect 104382 71406 104388 71470
rect 104861 71470 104927 71471
rect 104861 71438 104862 71470
rect 104312 71062 104388 71406
rect 104312 71030 104318 71062
rect 103632 70992 103708 70998
rect 104317 70998 104318 71030
rect 104382 71030 104388 71062
rect 104856 71406 104862 71438
rect 104926 71438 104927 71470
rect 105536 71470 105612 71476
rect 104926 71406 104932 71438
rect 104856 71062 104932 71406
rect 104382 70998 104383 71030
rect 104317 70997 104383 70998
rect 104856 70998 104862 71062
rect 104926 70998 104932 71062
rect 105536 71406 105542 71470
rect 105606 71406 105612 71470
rect 106085 71470 106151 71471
rect 106085 71438 106086 71470
rect 105536 71062 105612 71406
rect 105536 71030 105542 71062
rect 104856 70992 104932 70998
rect 105541 70998 105542 71030
rect 105606 71030 105612 71062
rect 106080 71406 106086 71438
rect 106150 71438 106151 71470
rect 107309 71470 107375 71471
rect 107309 71438 107310 71470
rect 106150 71406 106156 71438
rect 106080 71062 106156 71406
rect 105606 70998 105607 71030
rect 105541 70997 105607 70998
rect 106080 70998 106086 71062
rect 106150 70998 106156 71062
rect 106080 70992 106156 70998
rect 107304 71406 107310 71438
rect 107374 71438 107375 71470
rect 108533 71470 108599 71471
rect 108533 71438 108534 71470
rect 107374 71406 107380 71438
rect 107304 71062 107380 71406
rect 107304 70998 107310 71062
rect 107374 70998 107380 71062
rect 107304 70992 107380 70998
rect 108528 71406 108534 71438
rect 108598 71438 108599 71470
rect 108598 71406 108604 71438
rect 108528 71062 108604 71406
rect 108528 70998 108534 71062
rect 108598 70998 108604 71062
rect 108528 70992 108604 70998
rect 93296 70862 93302 70926
rect 93366 70862 93372 70926
rect 93296 70856 93372 70862
rect 109616 70926 109692 73038
rect 110709 71062 110775 71063
rect 110709 71030 110710 71062
rect 109616 70862 109622 70926
rect 109686 70862 109692 70926
rect 109616 70856 109692 70862
rect 110704 70998 110710 71030
rect 110774 71030 110775 71062
rect 110774 70998 110780 71030
rect 28968 70758 28974 70790
rect 28973 70726 28974 70758
rect 29038 70758 29044 70790
rect 29038 70726 29039 70758
rect 28973 70725 29039 70726
rect 110704 70654 110780 70998
rect 110704 70590 110710 70654
rect 110774 70590 110780 70654
rect 115328 70654 115404 74262
rect 115464 73102 115540 75622
rect 122264 75622 122270 75686
rect 122334 75622 122340 75686
rect 122264 75616 122340 75622
rect 122400 76910 122476 76916
rect 122400 76846 122406 76910
rect 122470 76846 122476 76910
rect 115464 73038 115470 73102
rect 115534 73038 115540 73102
rect 115464 73032 115540 73038
rect 122264 75550 122340 75556
rect 122264 75486 122270 75550
rect 122334 75486 122340 75550
rect 115877 72966 115943 72967
rect 115877 72934 115878 72966
rect 115328 70622 115334 70654
rect 110704 70584 110780 70590
rect 115333 70590 115334 70622
rect 115398 70622 115404 70654
rect 115872 72902 115878 72934
rect 115942 72934 115943 72966
rect 115942 72902 115948 72934
rect 115398 70590 115399 70622
rect 115333 70589 115399 70590
rect 114245 70518 114311 70519
rect 114245 70486 114246 70518
rect 114240 70454 114246 70486
rect 114310 70486 114311 70518
rect 114310 70454 114316 70486
rect 114240 70110 114316 70454
rect 114240 70046 114246 70110
rect 114310 70046 114316 70110
rect 114240 70040 114316 70046
rect 115872 70110 115948 72902
rect 122264 72830 122340 75486
rect 122400 74326 122476 76846
rect 122400 74294 122406 74326
rect 122405 74262 122406 74294
rect 122470 74294 122476 74326
rect 135320 76094 135668 77662
rect 135320 76030 135326 76094
rect 135390 76030 135668 76094
rect 122470 74262 122471 74294
rect 122405 74261 122471 74262
rect 135320 74190 135668 76030
rect 135320 74126 135326 74190
rect 135390 74126 135668 74190
rect 122405 74054 122471 74055
rect 122405 74022 122406 74054
rect 122264 72798 122270 72830
rect 122269 72766 122270 72798
rect 122334 72798 122340 72830
rect 122400 73990 122406 74022
rect 122470 74022 122471 74054
rect 122470 73990 122476 74022
rect 122334 72766 122335 72798
rect 122269 72765 122335 72766
rect 122400 71470 122476 73990
rect 135320 72558 135668 74126
rect 135320 72494 135326 72558
rect 135390 72494 135668 72558
rect 134092 72358 134158 72359
rect 134092 72294 134093 72358
rect 134157 72294 134158 72358
rect 134092 72293 134158 72294
rect 122400 71406 122406 71470
rect 122470 71406 122476 71470
rect 122400 71400 122476 71406
rect 115872 70046 115878 70110
rect 115942 70046 115948 70110
rect 115872 70040 115948 70046
rect 22168 69974 22244 69980
rect 22168 69910 22174 69974
rect 22238 69910 22244 69974
rect 22168 69702 22244 69910
rect 22168 69670 22174 69702
rect 22173 69638 22174 69670
rect 22238 69670 22244 69702
rect 22440 69974 22516 69980
rect 22440 69910 22446 69974
rect 22510 69910 22516 69974
rect 114381 69974 114447 69975
rect 114381 69942 114382 69974
rect 22440 69702 22516 69910
rect 22440 69670 22446 69702
rect 22238 69638 22239 69670
rect 22173 69637 22239 69638
rect 22445 69638 22446 69670
rect 22510 69670 22516 69702
rect 114376 69910 114382 69942
rect 114446 69942 114447 69974
rect 114648 69974 114724 69980
rect 114446 69910 114452 69942
rect 114376 69702 114452 69910
rect 22510 69638 22511 69670
rect 22445 69637 22511 69638
rect 114376 69638 114382 69702
rect 114446 69638 114452 69702
rect 114648 69910 114654 69974
rect 114718 69910 114724 69974
rect 115333 69974 115399 69975
rect 115333 69942 115334 69974
rect 114648 69702 114724 69910
rect 114648 69670 114654 69702
rect 114376 69632 114452 69638
rect 114653 69638 114654 69670
rect 114718 69670 114724 69702
rect 115328 69910 115334 69942
rect 115398 69942 115399 69974
rect 115464 69974 115540 69980
rect 115398 69910 115404 69942
rect 115328 69702 115404 69910
rect 114718 69638 114719 69670
rect 114653 69637 114719 69638
rect 115328 69638 115334 69702
rect 115398 69638 115404 69702
rect 115464 69910 115470 69974
rect 115534 69910 115540 69974
rect 115464 69702 115540 69910
rect 115464 69670 115470 69702
rect 115328 69632 115404 69638
rect 115469 69638 115470 69670
rect 115534 69670 115540 69702
rect 133144 69838 133220 69844
rect 133144 69774 133150 69838
rect 133214 69774 133220 69838
rect 115534 69638 115535 69670
rect 115469 69637 115535 69638
rect 20813 69566 20879 69567
rect 20813 69534 20814 69566
rect 952 69230 1230 69294
rect 1294 69230 1300 69294
rect 952 67526 1300 69230
rect 20808 69502 20814 69534
rect 20878 69534 20879 69566
rect 21357 69566 21423 69567
rect 21357 69534 21358 69566
rect 20878 69502 20884 69534
rect 20808 69294 20884 69502
rect 20808 69230 20814 69294
rect 20878 69230 20884 69294
rect 20808 69224 20884 69230
rect 21352 69502 21358 69534
rect 21422 69534 21423 69566
rect 21624 69566 21700 69572
rect 21422 69502 21428 69534
rect 21352 69294 21428 69502
rect 21352 69230 21358 69294
rect 21422 69230 21428 69294
rect 21624 69502 21630 69566
rect 21694 69502 21700 69566
rect 21624 69294 21700 69502
rect 21624 69262 21630 69294
rect 21352 69224 21428 69230
rect 21629 69230 21630 69262
rect 21694 69262 21700 69294
rect 22168 69566 22244 69572
rect 22168 69502 22174 69566
rect 22238 69502 22244 69566
rect 22445 69566 22511 69567
rect 22445 69534 22446 69566
rect 22168 69294 22244 69502
rect 22168 69262 22174 69294
rect 21694 69230 21695 69262
rect 21629 69229 21695 69230
rect 22173 69230 22174 69262
rect 22238 69262 22244 69294
rect 22440 69502 22446 69534
rect 22510 69534 22511 69566
rect 114240 69566 114316 69572
rect 22510 69502 22516 69534
rect 22440 69294 22516 69502
rect 22238 69230 22239 69262
rect 22173 69229 22239 69230
rect 22440 69230 22446 69294
rect 22510 69230 22516 69294
rect 114240 69502 114246 69566
rect 114310 69502 114316 69566
rect 114653 69566 114719 69567
rect 114653 69534 114654 69566
rect 114240 69294 114316 69502
rect 114240 69262 114246 69294
rect 22440 69224 22516 69230
rect 114245 69230 114246 69262
rect 114310 69262 114316 69294
rect 114648 69502 114654 69534
rect 114718 69534 114719 69566
rect 115056 69566 115132 69572
rect 114718 69502 114724 69534
rect 114648 69294 114724 69502
rect 114310 69230 114311 69262
rect 114245 69229 114311 69230
rect 114648 69230 114654 69294
rect 114718 69230 114724 69294
rect 115056 69502 115062 69566
rect 115126 69502 115132 69566
rect 115056 69294 115132 69502
rect 115056 69262 115062 69294
rect 114648 69224 114724 69230
rect 115061 69230 115062 69262
rect 115126 69262 115132 69294
rect 115600 69566 115676 69572
rect 115600 69502 115606 69566
rect 115670 69502 115676 69566
rect 115600 69294 115676 69502
rect 115600 69262 115606 69294
rect 115126 69230 115127 69262
rect 115061 69229 115127 69230
rect 115605 69230 115606 69262
rect 115670 69262 115676 69294
rect 116008 69566 116084 69572
rect 116008 69502 116014 69566
rect 116078 69502 116084 69566
rect 116008 69294 116084 69502
rect 116008 69262 116014 69294
rect 115670 69230 115671 69262
rect 115605 69229 115671 69230
rect 116013 69230 116014 69262
rect 116078 69262 116084 69294
rect 116078 69230 116079 69262
rect 116013 69229 116079 69230
rect 21760 69158 21836 69164
rect 21760 69094 21766 69158
rect 21830 69094 21836 69158
rect 22037 69158 22103 69159
rect 22037 69126 22038 69158
rect 20813 68886 20879 68887
rect 20813 68854 20814 68886
rect 20808 68822 20814 68854
rect 20878 68854 20879 68886
rect 21760 68886 21836 69094
rect 21760 68854 21766 68886
rect 20878 68822 20884 68854
rect 20808 68614 20884 68822
rect 21765 68822 21766 68854
rect 21830 68854 21836 68886
rect 22032 69094 22038 69126
rect 22102 69126 22103 69158
rect 22445 69158 22511 69159
rect 22445 69126 22446 69158
rect 22102 69094 22108 69126
rect 22032 68886 22108 69094
rect 21830 68822 21831 68854
rect 21765 68821 21831 68822
rect 22032 68822 22038 68886
rect 22102 68822 22108 68886
rect 22032 68816 22108 68822
rect 22440 69094 22446 69126
rect 22510 69126 22511 69158
rect 114381 69158 114447 69159
rect 114381 69126 114382 69158
rect 22510 69094 22516 69126
rect 22440 68886 22516 69094
rect 22440 68822 22446 68886
rect 22510 68822 22516 68886
rect 22440 68816 22516 68822
rect 114376 69094 114382 69126
rect 114446 69126 114447 69158
rect 114789 69158 114855 69159
rect 114789 69126 114790 69158
rect 114446 69094 114452 69126
rect 114376 68886 114452 69094
rect 114376 68822 114382 68886
rect 114446 68822 114452 68886
rect 114376 68816 114452 68822
rect 114784 69094 114790 69126
rect 114854 69126 114855 69158
rect 115192 69158 115268 69164
rect 114854 69094 114860 69126
rect 114784 68886 114860 69094
rect 114784 68822 114790 68886
rect 114854 68822 114860 68886
rect 115192 69094 115198 69158
rect 115262 69094 115268 69158
rect 115192 68886 115268 69094
rect 115192 68854 115198 68886
rect 114784 68816 114860 68822
rect 115197 68822 115198 68854
rect 115262 68854 115268 68886
rect 116008 68886 116084 68892
rect 115262 68822 115263 68854
rect 115197 68821 115263 68822
rect 116008 68822 116014 68886
rect 116078 68822 116084 68886
rect 22037 68750 22103 68751
rect 22037 68718 22038 68750
rect 20808 68550 20814 68614
rect 20878 68550 20884 68614
rect 20808 68544 20884 68550
rect 22032 68686 22038 68718
rect 22102 68718 22103 68750
rect 22440 68750 22516 68756
rect 22102 68686 22108 68718
rect 22032 68478 22108 68686
rect 22032 68414 22038 68478
rect 22102 68414 22108 68478
rect 22440 68686 22446 68750
rect 22510 68686 22516 68750
rect 114381 68750 114447 68751
rect 114381 68718 114382 68750
rect 22440 68478 22516 68686
rect 22440 68446 22446 68478
rect 22032 68408 22108 68414
rect 22445 68414 22446 68446
rect 22510 68446 22516 68478
rect 114376 68686 114382 68718
rect 114446 68718 114447 68750
rect 114648 68750 114724 68756
rect 114446 68686 114452 68718
rect 114376 68478 114452 68686
rect 22510 68414 22511 68446
rect 22445 68413 22511 68414
rect 114376 68414 114382 68478
rect 114446 68414 114452 68478
rect 114648 68686 114654 68750
rect 114718 68686 114724 68750
rect 114648 68478 114724 68686
rect 116008 68614 116084 68822
rect 116008 68582 116014 68614
rect 116013 68550 116014 68582
rect 116078 68582 116084 68614
rect 116078 68550 116079 68582
rect 116013 68549 116079 68550
rect 114648 68446 114654 68478
rect 114376 68408 114452 68414
rect 114653 68414 114654 68446
rect 114718 68446 114724 68478
rect 114718 68414 114719 68446
rect 114653 68413 114719 68414
rect 21896 68342 21972 68348
rect 21896 68278 21902 68342
rect 21966 68278 21972 68342
rect 20813 68070 20879 68071
rect 20813 68038 20814 68070
rect 20808 68006 20814 68038
rect 20878 68038 20879 68070
rect 21896 68070 21972 68278
rect 115328 68342 115404 68348
rect 115328 68278 115334 68342
rect 115398 68278 115404 68342
rect 21896 68038 21902 68070
rect 20878 68006 20884 68038
rect 20808 67798 20884 68006
rect 21901 68006 21902 68038
rect 21966 68038 21972 68070
rect 27472 68206 27548 68212
rect 27472 68142 27478 68206
rect 27542 68142 27548 68206
rect 109485 68206 109551 68207
rect 109485 68174 109486 68206
rect 21966 68006 21967 68038
rect 21901 68005 21967 68006
rect 27341 67934 27407 67935
rect 27341 67902 27342 67934
rect 20808 67734 20814 67798
rect 20878 67734 20884 67798
rect 20808 67728 20884 67734
rect 27336 67870 27342 67902
rect 27406 67902 27407 67934
rect 27472 67934 27548 68142
rect 27472 67902 27478 67934
rect 27406 67870 27412 67902
rect 952 67462 1230 67526
rect 1294 67462 1300 67526
rect 952 66030 1300 67462
rect 20808 67662 20884 67668
rect 20808 67598 20814 67662
rect 20878 67598 20884 67662
rect 20808 67390 20884 67598
rect 20808 67358 20814 67390
rect 20813 67326 20814 67358
rect 20878 67358 20884 67390
rect 21216 67662 21292 67668
rect 21216 67598 21222 67662
rect 21286 67598 21292 67662
rect 21216 67390 21292 67598
rect 21216 67358 21222 67390
rect 20878 67326 20879 67358
rect 20813 67325 20879 67326
rect 21221 67326 21222 67358
rect 21286 67358 21292 67390
rect 21624 67662 21700 67668
rect 21624 67598 21630 67662
rect 21694 67598 21700 67662
rect 21624 67390 21700 67598
rect 27336 67662 27412 67870
rect 27477 67870 27478 67902
rect 27542 67902 27548 67934
rect 109480 68142 109486 68174
rect 109550 68174 109551 68206
rect 109550 68142 109556 68174
rect 109480 67934 109556 68142
rect 115328 68070 115404 68278
rect 115328 68038 115334 68070
rect 115333 68006 115334 68038
rect 115398 68038 115404 68070
rect 115877 68070 115943 68071
rect 115877 68038 115878 68070
rect 115398 68006 115399 68038
rect 115333 68005 115399 68006
rect 115872 68006 115878 68038
rect 115942 68038 115943 68070
rect 115942 68006 115948 68038
rect 27542 67870 27543 67902
rect 27477 67869 27543 67870
rect 109480 67870 109486 67934
rect 109550 67870 109556 67934
rect 109480 67864 109556 67870
rect 27336 67598 27342 67662
rect 27406 67598 27412 67662
rect 27336 67592 27412 67598
rect 109344 67798 109420 67804
rect 109344 67734 109350 67798
rect 109414 67734 109420 67798
rect 21624 67358 21630 67390
rect 21286 67326 21287 67358
rect 21221 67325 21287 67326
rect 21629 67326 21630 67358
rect 21694 67358 21700 67390
rect 109344 67390 109420 67734
rect 115872 67798 115948 68006
rect 115872 67734 115878 67798
rect 115942 67734 115948 67798
rect 115872 67728 115948 67734
rect 115600 67662 115676 67668
rect 115600 67598 115606 67662
rect 115670 67598 115676 67662
rect 109344 67358 109350 67390
rect 21694 67326 21695 67358
rect 21629 67325 21695 67326
rect 109349 67326 109350 67358
rect 109414 67358 109420 67390
rect 109480 67390 109556 67396
rect 109414 67326 109415 67358
rect 109349 67325 109415 67326
rect 109480 67326 109486 67390
rect 109550 67326 109556 67390
rect 115600 67390 115676 67598
rect 115600 67358 115606 67390
rect 20808 67254 20884 67260
rect 20808 67190 20814 67254
rect 20878 67190 20884 67254
rect 21493 67254 21559 67255
rect 21493 67222 21494 67254
rect 20808 66982 20884 67190
rect 20808 66950 20814 66982
rect 20813 66918 20814 66950
rect 20878 66950 20884 66982
rect 21488 67190 21494 67222
rect 21558 67222 21559 67254
rect 22032 67254 22108 67260
rect 21558 67190 21564 67222
rect 21488 66982 21564 67190
rect 20878 66918 20879 66950
rect 20813 66917 20879 66918
rect 21488 66918 21494 66982
rect 21558 66918 21564 66982
rect 22032 67190 22038 67254
rect 22102 67190 22108 67254
rect 22032 66982 22108 67190
rect 22032 66950 22038 66982
rect 21488 66912 21564 66918
rect 22037 66918 22038 66950
rect 22102 66950 22108 66982
rect 22440 67254 22516 67260
rect 22440 67190 22446 67254
rect 22510 67190 22516 67254
rect 22440 66982 22516 67190
rect 109480 67118 109556 67326
rect 115605 67326 115606 67358
rect 115670 67358 115676 67390
rect 116008 67662 116084 67668
rect 116008 67598 116014 67662
rect 116078 67598 116084 67662
rect 116008 67390 116084 67598
rect 116008 67358 116014 67390
rect 115670 67326 115671 67358
rect 115605 67325 115671 67326
rect 116013 67326 116014 67358
rect 116078 67358 116084 67390
rect 116078 67326 116079 67358
rect 116013 67325 116079 67326
rect 109480 67086 109486 67118
rect 109485 67054 109486 67086
rect 109550 67086 109556 67118
rect 114376 67254 114452 67260
rect 114376 67190 114382 67254
rect 114446 67190 114452 67254
rect 114653 67254 114719 67255
rect 114653 67222 114654 67254
rect 109550 67054 109551 67086
rect 109485 67053 109551 67054
rect 22440 66950 22446 66982
rect 22102 66918 22103 66950
rect 22037 66917 22103 66918
rect 22445 66918 22446 66950
rect 22510 66950 22516 66982
rect 114376 66982 114452 67190
rect 114376 66950 114382 66982
rect 22510 66918 22511 66950
rect 22445 66917 22511 66918
rect 114381 66918 114382 66950
rect 114446 66950 114452 66982
rect 114648 67190 114654 67222
rect 114718 67222 114719 67254
rect 115872 67254 115948 67260
rect 114718 67190 114724 67222
rect 114648 66982 114724 67190
rect 114446 66918 114447 66950
rect 114381 66917 114447 66918
rect 114648 66918 114654 66982
rect 114718 66918 114724 66982
rect 115872 67190 115878 67254
rect 115942 67190 115948 67254
rect 115872 66982 115948 67190
rect 133144 67118 133220 69774
rect 133144 67086 133150 67118
rect 133149 67054 133150 67086
rect 133214 67086 133220 67118
rect 133214 67054 133215 67086
rect 133149 67053 133215 67054
rect 115872 66950 115878 66982
rect 114648 66912 114724 66918
rect 115877 66918 115878 66950
rect 115942 66950 115948 66982
rect 132600 66982 132676 66988
rect 115942 66918 115943 66950
rect 115877 66917 115943 66918
rect 132600 66918 132606 66982
rect 132670 66918 132676 66982
rect 20813 66846 20879 66847
rect 20813 66814 20814 66846
rect 20808 66782 20814 66814
rect 20878 66814 20879 66846
rect 21629 66846 21695 66847
rect 21629 66814 21630 66846
rect 20878 66782 20884 66814
rect 20808 66574 20884 66782
rect 20808 66510 20814 66574
rect 20878 66510 20884 66574
rect 20808 66504 20884 66510
rect 21624 66782 21630 66814
rect 21694 66814 21695 66846
rect 22032 66846 22108 66852
rect 21694 66782 21700 66814
rect 21624 66574 21700 66782
rect 21624 66510 21630 66574
rect 21694 66510 21700 66574
rect 22032 66782 22038 66846
rect 22102 66782 22108 66846
rect 22445 66846 22511 66847
rect 22445 66814 22446 66846
rect 22032 66574 22108 66782
rect 22032 66542 22038 66574
rect 21624 66504 21700 66510
rect 22037 66510 22038 66542
rect 22102 66542 22108 66574
rect 22440 66782 22446 66814
rect 22510 66814 22511 66846
rect 114376 66846 114452 66852
rect 22510 66782 22516 66814
rect 22440 66574 22516 66782
rect 22102 66510 22103 66542
rect 22037 66509 22103 66510
rect 22440 66510 22446 66574
rect 22510 66510 22516 66574
rect 114376 66782 114382 66846
rect 114446 66782 114452 66846
rect 114376 66574 114452 66782
rect 114376 66542 114382 66574
rect 22440 66504 22516 66510
rect 114381 66510 114382 66542
rect 114446 66542 114452 66574
rect 114784 66846 114860 66852
rect 114784 66782 114790 66846
rect 114854 66782 114860 66846
rect 114784 66574 114860 66782
rect 114784 66542 114790 66574
rect 114446 66510 114447 66542
rect 114381 66509 114447 66510
rect 114789 66510 114790 66542
rect 114854 66542 114860 66574
rect 115600 66846 115676 66852
rect 115600 66782 115606 66846
rect 115670 66782 115676 66846
rect 115877 66846 115943 66847
rect 115877 66814 115878 66846
rect 115600 66574 115676 66782
rect 115600 66542 115606 66574
rect 114854 66510 114855 66542
rect 114789 66509 114855 66510
rect 115605 66510 115606 66542
rect 115670 66542 115676 66574
rect 115872 66782 115878 66814
rect 115942 66814 115943 66846
rect 115942 66782 115948 66814
rect 115872 66574 115948 66782
rect 115670 66510 115671 66542
rect 115605 66509 115671 66510
rect 115872 66510 115878 66574
rect 115942 66510 115948 66574
rect 115872 66504 115948 66510
rect 20944 66438 21020 66444
rect 20944 66374 20950 66438
rect 21014 66374 21020 66438
rect 21357 66438 21423 66439
rect 21357 66406 21358 66438
rect 20944 66166 21020 66374
rect 20944 66134 20950 66166
rect 20949 66102 20950 66134
rect 21014 66134 21020 66166
rect 21352 66374 21358 66406
rect 21422 66406 21423 66438
rect 21493 66438 21559 66439
rect 21493 66406 21494 66438
rect 21422 66374 21428 66406
rect 21352 66166 21428 66374
rect 21014 66102 21015 66134
rect 20949 66101 21015 66102
rect 21352 66102 21358 66166
rect 21422 66102 21428 66166
rect 21352 66096 21428 66102
rect 21488 66374 21494 66406
rect 21558 66406 21559 66438
rect 22173 66438 22239 66439
rect 22173 66406 22174 66438
rect 21558 66374 21564 66406
rect 21488 66166 21564 66374
rect 21488 66102 21494 66166
rect 21558 66102 21564 66166
rect 21488 66096 21564 66102
rect 22168 66374 22174 66406
rect 22238 66406 22239 66438
rect 22576 66438 22652 66444
rect 22238 66374 22244 66406
rect 22168 66166 22244 66374
rect 22168 66102 22174 66166
rect 22238 66102 22244 66166
rect 22576 66374 22582 66438
rect 22646 66374 22652 66438
rect 114245 66438 114311 66439
rect 114245 66406 114246 66438
rect 22576 66166 22652 66374
rect 22576 66134 22582 66166
rect 22168 66096 22244 66102
rect 22581 66102 22582 66134
rect 22646 66134 22652 66166
rect 114240 66374 114246 66406
rect 114310 66406 114311 66438
rect 114653 66438 114719 66439
rect 114653 66406 114654 66438
rect 114310 66374 114316 66406
rect 114240 66166 114316 66374
rect 22646 66102 22647 66134
rect 22581 66101 22647 66102
rect 114240 66102 114246 66166
rect 114310 66102 114316 66166
rect 114240 66096 114316 66102
rect 114648 66374 114654 66406
rect 114718 66406 114719 66438
rect 115061 66438 115127 66439
rect 115061 66406 115062 66438
rect 114718 66374 114724 66406
rect 114648 66166 114724 66374
rect 114648 66102 114654 66166
rect 114718 66102 114724 66166
rect 114648 66096 114724 66102
rect 115056 66374 115062 66406
rect 115126 66406 115127 66438
rect 115333 66438 115399 66439
rect 115333 66406 115334 66438
rect 115126 66374 115132 66406
rect 115056 66166 115132 66374
rect 115056 66102 115062 66166
rect 115126 66102 115132 66166
rect 115056 66096 115132 66102
rect 115328 66374 115334 66406
rect 115398 66406 115399 66438
rect 116013 66438 116079 66439
rect 116013 66406 116014 66438
rect 115398 66374 115404 66406
rect 115328 66166 115404 66374
rect 115328 66102 115334 66166
rect 115398 66102 115404 66166
rect 115328 66096 115404 66102
rect 116008 66374 116014 66406
rect 116078 66406 116079 66438
rect 116078 66374 116084 66406
rect 116008 66166 116084 66374
rect 116008 66102 116014 66166
rect 116078 66102 116084 66166
rect 116008 66096 116084 66102
rect 952 65966 1230 66030
rect 1294 65966 1300 66030
rect 952 64126 1300 65966
rect 20808 66030 20884 66036
rect 20808 65966 20814 66030
rect 20878 65966 20884 66030
rect 21765 66030 21831 66031
rect 21765 65998 21766 66030
rect 20808 65758 20884 65966
rect 20808 65726 20814 65758
rect 20813 65694 20814 65726
rect 20878 65726 20884 65758
rect 21760 65966 21766 65998
rect 21830 65998 21831 66030
rect 22032 66030 22108 66036
rect 21830 65966 21836 65998
rect 21760 65758 21836 65966
rect 20878 65694 20879 65726
rect 20813 65693 20879 65694
rect 21760 65694 21766 65758
rect 21830 65694 21836 65758
rect 22032 65966 22038 66030
rect 22102 65966 22108 66030
rect 22581 66030 22647 66031
rect 22581 65998 22582 66030
rect 22032 65758 22108 65966
rect 22032 65726 22038 65758
rect 21760 65688 21836 65694
rect 22037 65694 22038 65726
rect 22102 65726 22108 65758
rect 22576 65966 22582 65998
rect 22646 65998 22647 66030
rect 114376 66030 114452 66036
rect 22646 65966 22652 65998
rect 22576 65758 22652 65966
rect 22102 65694 22103 65726
rect 22037 65693 22103 65694
rect 22576 65694 22582 65758
rect 22646 65694 22652 65758
rect 114376 65966 114382 66030
rect 114446 65966 114452 66030
rect 114653 66030 114719 66031
rect 114653 65998 114654 66030
rect 114376 65758 114452 65966
rect 114376 65726 114382 65758
rect 22576 65688 22652 65694
rect 114381 65694 114382 65726
rect 114446 65726 114452 65758
rect 114648 65966 114654 65998
rect 114718 65998 114719 66030
rect 115605 66030 115671 66031
rect 115605 65998 115606 66030
rect 114718 65966 114724 65998
rect 114648 65758 114724 65966
rect 114446 65694 114447 65726
rect 114381 65693 114447 65694
rect 114648 65694 114654 65758
rect 114718 65694 114724 65758
rect 114648 65688 114724 65694
rect 115600 65966 115606 65998
rect 115670 65998 115671 66030
rect 116013 66030 116079 66031
rect 116013 65998 116014 66030
rect 115670 65966 115676 65998
rect 115600 65758 115676 65966
rect 115600 65694 115606 65758
rect 115670 65694 115676 65758
rect 115600 65688 115676 65694
rect 116008 65966 116014 65998
rect 116078 65998 116079 66030
rect 116078 65966 116084 65998
rect 116008 65758 116084 65966
rect 116008 65694 116014 65758
rect 116078 65694 116084 65758
rect 116008 65688 116084 65694
rect 20949 65622 21015 65623
rect 20949 65590 20950 65622
rect 20944 65558 20950 65590
rect 21014 65590 21015 65622
rect 21352 65622 21428 65628
rect 21014 65558 21020 65590
rect 20944 65350 21020 65558
rect 20944 65286 20950 65350
rect 21014 65286 21020 65350
rect 21352 65558 21358 65622
rect 21422 65558 21428 65622
rect 21352 65350 21428 65558
rect 21352 65318 21358 65350
rect 20944 65280 21020 65286
rect 21357 65286 21358 65318
rect 21422 65318 21428 65350
rect 21488 65622 21564 65628
rect 21488 65558 21494 65622
rect 21558 65558 21564 65622
rect 22037 65622 22103 65623
rect 22037 65590 22038 65622
rect 21488 65350 21564 65558
rect 21488 65318 21494 65350
rect 21422 65286 21423 65318
rect 21357 65285 21423 65286
rect 21493 65286 21494 65318
rect 21558 65318 21564 65350
rect 22032 65558 22038 65590
rect 22102 65590 22103 65622
rect 22440 65622 22516 65628
rect 22102 65558 22108 65590
rect 22032 65350 22108 65558
rect 21558 65286 21559 65318
rect 21493 65285 21559 65286
rect 22032 65286 22038 65350
rect 22102 65286 22108 65350
rect 22440 65558 22446 65622
rect 22510 65558 22516 65622
rect 114381 65622 114447 65623
rect 114381 65590 114382 65622
rect 22440 65350 22516 65558
rect 22440 65318 22446 65350
rect 22032 65280 22108 65286
rect 22445 65286 22446 65318
rect 22510 65318 22516 65350
rect 114376 65558 114382 65590
rect 114446 65590 114447 65622
rect 114648 65622 114724 65628
rect 114446 65558 114452 65590
rect 114376 65350 114452 65558
rect 22510 65286 22511 65318
rect 22445 65285 22511 65286
rect 114376 65286 114382 65350
rect 114446 65286 114452 65350
rect 114648 65558 114654 65622
rect 114718 65558 114724 65622
rect 115197 65622 115263 65623
rect 115197 65590 115198 65622
rect 114648 65350 114724 65558
rect 114648 65318 114654 65350
rect 114376 65280 114452 65286
rect 114653 65286 114654 65318
rect 114718 65318 114724 65350
rect 115192 65558 115198 65590
rect 115262 65590 115263 65622
rect 115333 65622 115399 65623
rect 115333 65590 115334 65622
rect 115262 65558 115268 65590
rect 115192 65350 115268 65558
rect 114718 65286 114719 65318
rect 114653 65285 114719 65286
rect 115192 65286 115198 65350
rect 115262 65286 115268 65350
rect 115192 65280 115268 65286
rect 115328 65558 115334 65590
rect 115398 65590 115399 65622
rect 115877 65622 115943 65623
rect 115877 65590 115878 65622
rect 115398 65558 115404 65590
rect 115328 65350 115404 65558
rect 115328 65286 115334 65350
rect 115398 65286 115404 65350
rect 115328 65280 115404 65286
rect 115872 65558 115878 65590
rect 115942 65590 115943 65622
rect 115942 65558 115948 65590
rect 115872 65350 115948 65558
rect 115872 65286 115878 65350
rect 115942 65286 115948 65350
rect 115872 65280 115948 65286
rect 21901 65214 21967 65215
rect 21901 65182 21902 65214
rect 21896 65150 21902 65182
rect 21966 65182 21967 65214
rect 22168 65214 22244 65220
rect 21966 65150 21972 65182
rect 21896 64942 21972 65150
rect 22168 65150 22174 65214
rect 22238 65150 22244 65214
rect 22445 65214 22511 65215
rect 22445 65182 22446 65214
rect 22037 65078 22103 65079
rect 22037 65046 22038 65078
rect 21896 64878 21902 64942
rect 21966 64878 21972 64942
rect 21896 64872 21972 64878
rect 22032 65014 22038 65046
rect 22102 65046 22103 65078
rect 22102 65014 22108 65046
rect 22032 64534 22108 65014
rect 22168 64942 22244 65150
rect 22168 64910 22174 64942
rect 22173 64878 22174 64910
rect 22238 64910 22244 64942
rect 22440 65150 22446 65182
rect 22510 65182 22511 65214
rect 114245 65214 114311 65215
rect 114245 65182 114246 65214
rect 22510 65150 22516 65182
rect 22440 64942 22516 65150
rect 114240 65150 114246 65182
rect 114310 65182 114311 65214
rect 114653 65214 114719 65215
rect 114653 65182 114654 65214
rect 114310 65150 114316 65182
rect 27613 65078 27679 65079
rect 27613 65046 27614 65078
rect 22238 64878 22239 64910
rect 22173 64877 22239 64878
rect 22440 64878 22446 64942
rect 22510 64878 22516 64942
rect 22440 64872 22516 64878
rect 27608 65014 27614 65046
rect 27678 65046 27679 65078
rect 27678 65014 27684 65046
rect 22173 64806 22239 64807
rect 22173 64774 22174 64806
rect 22032 64470 22038 64534
rect 22102 64470 22108 64534
rect 22032 64464 22108 64470
rect 22168 64742 22174 64774
rect 22238 64774 22239 64806
rect 22576 64806 22652 64812
rect 22238 64742 22244 64774
rect 22168 64534 22244 64742
rect 22168 64470 22174 64534
rect 22238 64470 22244 64534
rect 22576 64742 22582 64806
rect 22646 64742 22652 64806
rect 22576 64534 22652 64742
rect 27608 64806 27684 65014
rect 114240 64942 114316 65150
rect 114240 64878 114246 64942
rect 114310 64878 114316 64942
rect 114240 64872 114316 64878
rect 114648 65150 114654 65182
rect 114718 65182 114719 65214
rect 115056 65214 115132 65220
rect 114718 65150 114724 65182
rect 114648 64942 114724 65150
rect 114648 64878 114654 64942
rect 114718 64878 114724 64942
rect 115056 65150 115062 65214
rect 115126 65150 115132 65214
rect 115469 65214 115535 65215
rect 115469 65182 115470 65214
rect 115056 64942 115132 65150
rect 115056 64910 115062 64942
rect 114648 64872 114724 64878
rect 115061 64878 115062 64910
rect 115126 64910 115132 64942
rect 115464 65150 115470 65182
rect 115534 65182 115535 65214
rect 115534 65150 115540 65182
rect 115464 64942 115540 65150
rect 115126 64878 115127 64910
rect 115061 64877 115127 64878
rect 115464 64878 115470 64942
rect 115534 64878 115540 64942
rect 115464 64872 115540 64878
rect 27608 64742 27614 64806
rect 27678 64742 27684 64806
rect 109349 64806 109415 64807
rect 109349 64774 109350 64806
rect 27608 64736 27684 64742
rect 109344 64742 109350 64774
rect 109414 64774 109415 64806
rect 114376 64806 114452 64812
rect 109414 64742 109420 64774
rect 22576 64502 22582 64534
rect 22168 64464 22244 64470
rect 22581 64470 22582 64502
rect 22646 64502 22652 64534
rect 27336 64534 27412 64540
rect 22646 64470 22647 64502
rect 22581 64469 22647 64470
rect 27336 64470 27342 64534
rect 27406 64470 27412 64534
rect 21760 64398 21836 64404
rect 21760 64334 21766 64398
rect 21830 64334 21836 64398
rect 952 64062 1230 64126
rect 1294 64062 1300 64126
rect 20813 64126 20879 64127
rect 20813 64094 20814 64126
rect 952 62630 1300 64062
rect 20808 64062 20814 64094
rect 20878 64094 20879 64126
rect 21760 64126 21836 64334
rect 27336 64262 27412 64470
rect 109344 64398 109420 64742
rect 114376 64742 114382 64806
rect 114446 64742 114452 64806
rect 114653 64806 114719 64807
rect 114653 64774 114654 64806
rect 114376 64534 114452 64742
rect 114376 64502 114382 64534
rect 114381 64470 114382 64502
rect 114446 64502 114452 64534
rect 114648 64742 114654 64774
rect 114718 64774 114719 64806
rect 114718 64742 114724 64774
rect 114648 64534 114724 64742
rect 114446 64470 114447 64502
rect 114381 64469 114447 64470
rect 114648 64470 114654 64534
rect 114718 64470 114724 64534
rect 114648 64464 114724 64470
rect 109344 64334 109350 64398
rect 109414 64334 109420 64398
rect 115333 64398 115399 64399
rect 115333 64366 115334 64398
rect 109344 64328 109420 64334
rect 115328 64334 115334 64366
rect 115398 64366 115399 64398
rect 132600 64398 132676 66918
rect 132600 64366 132606 64398
rect 115398 64334 115404 64366
rect 27336 64230 27342 64262
rect 27341 64198 27342 64230
rect 27406 64230 27412 64262
rect 27613 64262 27679 64263
rect 27613 64230 27614 64262
rect 27406 64198 27407 64230
rect 27341 64197 27407 64198
rect 27608 64198 27614 64230
rect 27678 64230 27679 64262
rect 109485 64262 109551 64263
rect 109485 64230 109486 64262
rect 27678 64198 27684 64230
rect 21760 64094 21766 64126
rect 20878 64062 20884 64094
rect 20808 63854 20884 64062
rect 21765 64062 21766 64094
rect 21830 64094 21836 64126
rect 21830 64062 21831 64094
rect 21765 64061 21831 64062
rect 27608 63990 27684 64198
rect 109480 64198 109486 64230
rect 109550 64230 109551 64262
rect 109550 64198 109556 64230
rect 27608 63926 27614 63990
rect 27678 63926 27684 63990
rect 27608 63920 27684 63926
rect 109208 63990 109284 63996
rect 109208 63926 109214 63990
rect 109278 63926 109284 63990
rect 20808 63790 20814 63854
rect 20878 63790 20884 63854
rect 20808 63784 20884 63790
rect 27472 63854 27548 63860
rect 27472 63790 27478 63854
rect 27542 63790 27548 63854
rect 20813 63718 20879 63719
rect 20813 63686 20814 63718
rect 20808 63654 20814 63686
rect 20878 63686 20879 63718
rect 21901 63718 21967 63719
rect 21901 63686 21902 63718
rect 20878 63654 20884 63686
rect 20808 63446 20884 63654
rect 20808 63382 20814 63446
rect 20878 63382 20884 63446
rect 20808 63376 20884 63382
rect 21896 63654 21902 63686
rect 21966 63686 21967 63718
rect 21966 63654 21972 63686
rect 21896 63446 21972 63654
rect 27472 63582 27548 63790
rect 27472 63550 27478 63582
rect 27477 63518 27478 63550
rect 27542 63550 27548 63582
rect 109208 63582 109284 63926
rect 109480 63990 109556 64198
rect 115328 64126 115404 64334
rect 132605 64334 132606 64366
rect 132670 64366 132676 64398
rect 132670 64334 132671 64366
rect 132605 64333 132671 64334
rect 133421 64262 133487 64263
rect 133421 64230 133422 64262
rect 133416 64198 133422 64230
rect 133486 64230 133487 64262
rect 133486 64198 133492 64230
rect 115328 64062 115334 64126
rect 115398 64062 115404 64126
rect 116013 64126 116079 64127
rect 116013 64094 116014 64126
rect 115328 64056 115404 64062
rect 116008 64062 116014 64094
rect 116078 64094 116079 64126
rect 116078 64062 116084 64094
rect 109480 63926 109486 63990
rect 109550 63926 109556 63990
rect 109480 63920 109556 63926
rect 109208 63550 109214 63582
rect 27542 63518 27543 63550
rect 27477 63517 27543 63518
rect 109213 63518 109214 63550
rect 109278 63550 109284 63582
rect 109344 63854 109420 63860
rect 109344 63790 109350 63854
rect 109414 63790 109420 63854
rect 109344 63582 109420 63790
rect 116008 63854 116084 64062
rect 116008 63790 116014 63854
rect 116078 63790 116084 63854
rect 116008 63784 116084 63790
rect 109344 63550 109350 63582
rect 109278 63518 109279 63550
rect 109213 63517 109279 63518
rect 109349 63518 109350 63550
rect 109414 63550 109420 63582
rect 115464 63718 115540 63724
rect 115464 63654 115470 63718
rect 115534 63654 115540 63718
rect 109414 63518 109415 63550
rect 109349 63517 109415 63518
rect 21896 63382 21902 63446
rect 21966 63382 21972 63446
rect 115464 63446 115540 63654
rect 115464 63414 115470 63446
rect 21896 63376 21972 63382
rect 115469 63382 115470 63414
rect 115534 63414 115540 63446
rect 115872 63718 115948 63724
rect 115872 63654 115878 63718
rect 115942 63654 115948 63718
rect 115872 63446 115948 63654
rect 115872 63414 115878 63446
rect 115534 63382 115535 63414
rect 115469 63381 115535 63382
rect 115877 63382 115878 63414
rect 115942 63414 115948 63446
rect 115942 63382 115943 63414
rect 115877 63381 115943 63382
rect 20808 63310 20884 63316
rect 20808 63246 20814 63310
rect 20878 63246 20884 63310
rect 22037 63310 22103 63311
rect 22037 63278 22038 63310
rect 20808 63038 20884 63246
rect 20808 63006 20814 63038
rect 20813 62974 20814 63006
rect 20878 63006 20884 63038
rect 22032 63246 22038 63278
rect 22102 63278 22103 63310
rect 22581 63310 22647 63311
rect 22581 63278 22582 63310
rect 22102 63246 22108 63278
rect 22032 63038 22108 63246
rect 20878 62974 20879 63006
rect 20813 62973 20879 62974
rect 22032 62974 22038 63038
rect 22102 62974 22108 63038
rect 22032 62968 22108 62974
rect 22576 63246 22582 63278
rect 22646 63278 22647 63310
rect 114240 63310 114316 63316
rect 22646 63246 22652 63278
rect 22576 63038 22652 63246
rect 22576 62974 22582 63038
rect 22646 62974 22652 63038
rect 114240 63246 114246 63310
rect 114310 63246 114316 63310
rect 114789 63310 114855 63311
rect 114789 63278 114790 63310
rect 114240 63038 114316 63246
rect 114240 63006 114246 63038
rect 22576 62968 22652 62974
rect 114245 62974 114246 63006
rect 114310 63006 114316 63038
rect 114784 63246 114790 63278
rect 114854 63278 114855 63310
rect 116008 63310 116084 63316
rect 114854 63246 114860 63278
rect 114784 63038 114860 63246
rect 114310 62974 114311 63006
rect 114245 62973 114311 62974
rect 114784 62974 114790 63038
rect 114854 62974 114860 63038
rect 116008 63246 116014 63310
rect 116078 63246 116084 63310
rect 116008 63038 116084 63246
rect 116008 63006 116014 63038
rect 114784 62968 114860 62974
rect 116013 62974 116014 63006
rect 116078 63006 116084 63038
rect 116078 62974 116079 63006
rect 116013 62973 116079 62974
rect 20813 62902 20879 62903
rect 20813 62870 20814 62902
rect 952 62566 1230 62630
rect 1294 62566 1300 62630
rect 952 60998 1300 62566
rect 20808 62838 20814 62870
rect 20878 62870 20879 62902
rect 21765 62902 21831 62903
rect 21765 62870 21766 62902
rect 20878 62838 20884 62870
rect 20808 62630 20884 62838
rect 20808 62566 20814 62630
rect 20878 62566 20884 62630
rect 20808 62560 20884 62566
rect 21760 62838 21766 62870
rect 21830 62870 21831 62902
rect 22032 62902 22108 62908
rect 21830 62838 21836 62870
rect 21760 62630 21836 62838
rect 21760 62566 21766 62630
rect 21830 62566 21836 62630
rect 22032 62838 22038 62902
rect 22102 62838 22108 62902
rect 22032 62630 22108 62838
rect 22032 62598 22038 62630
rect 21760 62560 21836 62566
rect 22037 62566 22038 62598
rect 22102 62598 22108 62630
rect 22440 62902 22516 62908
rect 22440 62838 22446 62902
rect 22510 62838 22516 62902
rect 114245 62902 114311 62903
rect 114245 62870 114246 62902
rect 22440 62630 22516 62838
rect 114240 62838 114246 62870
rect 114310 62870 114311 62902
rect 114653 62902 114719 62903
rect 114653 62870 114654 62902
rect 114310 62838 114316 62870
rect 22440 62598 22446 62630
rect 22102 62566 22103 62598
rect 22037 62565 22103 62566
rect 22445 62566 22446 62598
rect 22510 62598 22516 62630
rect 109349 62630 109415 62631
rect 109349 62598 109350 62630
rect 22510 62566 22511 62598
rect 22445 62565 22511 62566
rect 109344 62566 109350 62598
rect 109414 62598 109415 62630
rect 114240 62630 114316 62838
rect 109414 62566 109420 62598
rect 20813 62494 20879 62495
rect 20813 62462 20814 62494
rect 20808 62430 20814 62462
rect 20878 62462 20879 62494
rect 21221 62494 21287 62495
rect 21221 62462 21222 62494
rect 20878 62430 20884 62462
rect 20808 62222 20884 62430
rect 20808 62158 20814 62222
rect 20878 62158 20884 62222
rect 20808 62152 20884 62158
rect 21216 62430 21222 62462
rect 21286 62462 21287 62494
rect 21624 62494 21700 62500
rect 21286 62430 21292 62462
rect 21216 62222 21292 62430
rect 21216 62158 21222 62222
rect 21286 62158 21292 62222
rect 21624 62430 21630 62494
rect 21694 62430 21700 62494
rect 22037 62494 22103 62495
rect 22037 62462 22038 62494
rect 21624 62222 21700 62430
rect 21624 62190 21630 62222
rect 21216 62152 21292 62158
rect 21629 62158 21630 62190
rect 21694 62190 21700 62222
rect 22032 62430 22038 62462
rect 22102 62462 22103 62494
rect 22576 62494 22652 62500
rect 22102 62430 22108 62462
rect 22032 62222 22108 62430
rect 21694 62158 21695 62190
rect 21629 62157 21695 62158
rect 22032 62158 22038 62222
rect 22102 62158 22108 62222
rect 22576 62430 22582 62494
rect 22646 62430 22652 62494
rect 22576 62222 22652 62430
rect 109344 62358 109420 62566
rect 114240 62566 114246 62630
rect 114310 62566 114316 62630
rect 114240 62560 114316 62566
rect 114648 62838 114654 62870
rect 114718 62870 114719 62902
rect 115061 62902 115127 62903
rect 115061 62870 115062 62902
rect 114718 62838 114724 62870
rect 114648 62630 114724 62838
rect 114648 62566 114654 62630
rect 114718 62566 114724 62630
rect 114648 62560 114724 62566
rect 115056 62838 115062 62870
rect 115126 62870 115127 62902
rect 115464 62902 115540 62908
rect 115126 62838 115132 62870
rect 115056 62630 115132 62838
rect 115056 62566 115062 62630
rect 115126 62566 115132 62630
rect 115464 62838 115470 62902
rect 115534 62838 115540 62902
rect 115464 62630 115540 62838
rect 115464 62598 115470 62630
rect 115056 62560 115132 62566
rect 115469 62566 115470 62598
rect 115534 62598 115540 62630
rect 115872 62902 115948 62908
rect 115872 62838 115878 62902
rect 115942 62838 115948 62902
rect 115872 62630 115948 62838
rect 115872 62598 115878 62630
rect 115534 62566 115535 62598
rect 115469 62565 115535 62566
rect 115877 62566 115878 62598
rect 115942 62598 115948 62630
rect 115942 62566 115943 62598
rect 115877 62565 115943 62566
rect 109344 62294 109350 62358
rect 109414 62294 109420 62358
rect 109344 62288 109420 62294
rect 114376 62494 114452 62500
rect 114376 62430 114382 62494
rect 114446 62430 114452 62494
rect 22576 62190 22582 62222
rect 22032 62152 22108 62158
rect 22581 62158 22582 62190
rect 22646 62190 22652 62222
rect 114376 62222 114452 62430
rect 114376 62190 114382 62222
rect 22646 62158 22647 62190
rect 22581 62157 22647 62158
rect 114381 62158 114382 62190
rect 114446 62190 114452 62222
rect 114784 62494 114860 62500
rect 114784 62430 114790 62494
rect 114854 62430 114860 62494
rect 114784 62222 114860 62430
rect 114784 62190 114790 62222
rect 114446 62158 114447 62190
rect 114381 62157 114447 62158
rect 114789 62158 114790 62190
rect 114854 62190 114860 62222
rect 115192 62494 115268 62500
rect 115192 62430 115198 62494
rect 115262 62430 115268 62494
rect 115877 62494 115943 62495
rect 115877 62462 115878 62494
rect 115192 62222 115268 62430
rect 115192 62190 115198 62222
rect 114854 62158 114855 62190
rect 114789 62157 114855 62158
rect 115197 62158 115198 62190
rect 115262 62190 115268 62222
rect 115872 62430 115878 62462
rect 115942 62462 115943 62494
rect 115942 62430 115948 62462
rect 115872 62222 115948 62430
rect 115262 62158 115263 62190
rect 115197 62157 115263 62158
rect 115872 62158 115878 62222
rect 115942 62158 115948 62222
rect 115872 62152 115948 62158
rect 20944 62086 21020 62092
rect 20944 62022 20950 62086
rect 21014 62022 21020 62086
rect 20944 61814 21020 62022
rect 20944 61782 20950 61814
rect 20949 61750 20950 61782
rect 21014 61782 21020 61814
rect 21352 62086 21428 62092
rect 21352 62022 21358 62086
rect 21422 62022 21428 62086
rect 22173 62086 22239 62087
rect 22173 62054 22174 62086
rect 21352 61814 21428 62022
rect 21352 61782 21358 61814
rect 21014 61750 21015 61782
rect 20949 61749 21015 61750
rect 21357 61750 21358 61782
rect 21422 61782 21428 61814
rect 22168 62022 22174 62054
rect 22238 62054 22239 62086
rect 22445 62086 22511 62087
rect 22445 62054 22446 62086
rect 22238 62022 22244 62054
rect 22168 61814 22244 62022
rect 21422 61750 21423 61782
rect 21357 61749 21423 61750
rect 22168 61750 22174 61814
rect 22238 61750 22244 61814
rect 22168 61744 22244 61750
rect 22440 62022 22446 62054
rect 22510 62054 22511 62086
rect 114245 62086 114311 62087
rect 114245 62054 114246 62086
rect 22510 62022 22516 62054
rect 22440 61814 22516 62022
rect 22440 61750 22446 61814
rect 22510 61750 22516 61814
rect 22440 61744 22516 61750
rect 114240 62022 114246 62054
rect 114310 62054 114311 62086
rect 114648 62086 114724 62092
rect 114310 62022 114316 62054
rect 114240 61814 114316 62022
rect 114240 61750 114246 61814
rect 114310 61750 114316 61814
rect 114648 62022 114654 62086
rect 114718 62022 114724 62086
rect 115469 62086 115535 62087
rect 115469 62054 115470 62086
rect 114648 61814 114724 62022
rect 114648 61782 114654 61814
rect 114240 61744 114316 61750
rect 114653 61750 114654 61782
rect 114718 61782 114724 61814
rect 115464 62022 115470 62054
rect 115534 62054 115535 62086
rect 116013 62086 116079 62087
rect 116013 62054 116014 62086
rect 115534 62022 115540 62054
rect 115464 61814 115540 62022
rect 114718 61750 114719 61782
rect 114653 61749 114719 61750
rect 115464 61750 115470 61814
rect 115534 61750 115540 61814
rect 115464 61744 115540 61750
rect 116008 62022 116014 62054
rect 116078 62054 116079 62086
rect 116078 62022 116084 62054
rect 116008 61814 116084 62022
rect 116008 61750 116014 61814
rect 116078 61750 116084 61814
rect 116008 61744 116084 61750
rect 20949 61678 21015 61679
rect 20949 61646 20950 61678
rect 20944 61614 20950 61646
rect 21014 61646 21015 61678
rect 21765 61678 21831 61679
rect 21765 61646 21766 61678
rect 21014 61614 21020 61646
rect 20944 61406 21020 61614
rect 20944 61342 20950 61406
rect 21014 61342 21020 61406
rect 20944 61336 21020 61342
rect 21760 61614 21766 61646
rect 21830 61646 21831 61678
rect 22032 61678 22108 61684
rect 21830 61614 21836 61646
rect 21760 61406 21836 61614
rect 21760 61342 21766 61406
rect 21830 61342 21836 61406
rect 22032 61614 22038 61678
rect 22102 61614 22108 61678
rect 22032 61406 22108 61614
rect 22032 61374 22038 61406
rect 21760 61336 21836 61342
rect 22037 61342 22038 61374
rect 22102 61374 22108 61406
rect 22440 61678 22516 61684
rect 22440 61614 22446 61678
rect 22510 61614 22516 61678
rect 114245 61678 114311 61679
rect 114245 61646 114246 61678
rect 22440 61406 22516 61614
rect 22440 61374 22446 61406
rect 22102 61342 22103 61374
rect 22037 61341 22103 61342
rect 22445 61342 22446 61374
rect 22510 61374 22516 61406
rect 114240 61614 114246 61646
rect 114310 61646 114311 61678
rect 114653 61678 114719 61679
rect 114653 61646 114654 61678
rect 114310 61614 114316 61646
rect 114240 61406 114316 61614
rect 22510 61342 22511 61374
rect 22445 61341 22511 61342
rect 114240 61342 114246 61406
rect 114310 61342 114316 61406
rect 114240 61336 114316 61342
rect 114648 61614 114654 61646
rect 114718 61646 114719 61678
rect 115061 61678 115127 61679
rect 115061 61646 115062 61678
rect 114718 61614 114724 61646
rect 114648 61406 114724 61614
rect 114648 61342 114654 61406
rect 114718 61342 114724 61406
rect 114648 61336 114724 61342
rect 115056 61614 115062 61646
rect 115126 61646 115127 61678
rect 115605 61678 115671 61679
rect 115605 61646 115606 61678
rect 115126 61614 115132 61646
rect 115056 61406 115132 61614
rect 115056 61342 115062 61406
rect 115126 61342 115132 61406
rect 115056 61336 115132 61342
rect 115600 61614 115606 61646
rect 115670 61646 115671 61678
rect 115872 61678 115948 61684
rect 115670 61614 115676 61646
rect 115600 61406 115676 61614
rect 115600 61342 115606 61406
rect 115670 61342 115676 61406
rect 115872 61614 115878 61678
rect 115942 61614 115948 61678
rect 115872 61406 115948 61614
rect 133416 61542 133492 64198
rect 134095 62124 134155 72293
rect 134781 71334 134847 71335
rect 134781 71302 134782 71334
rect 134776 71270 134782 71302
rect 134846 71302 134847 71334
rect 134846 71270 134852 71302
rect 134776 71062 134852 71270
rect 134776 70998 134782 71062
rect 134846 70998 134852 71062
rect 134776 70992 134852 70998
rect 135320 70926 135668 72494
rect 135320 70862 135326 70926
rect 135390 70862 135668 70926
rect 135320 69430 135668 70862
rect 135320 69366 135326 69430
rect 135390 69366 135668 69430
rect 134776 69158 134852 69164
rect 134776 69094 134782 69158
rect 134846 69094 134852 69158
rect 134776 68614 134852 69094
rect 134776 68582 134782 68614
rect 134781 68550 134782 68582
rect 134846 68582 134852 68614
rect 134846 68550 134847 68582
rect 134781 68549 134847 68550
rect 135320 67662 135668 69366
rect 135320 67598 135326 67662
rect 135390 67598 135668 67662
rect 135320 65894 135668 67598
rect 135320 65830 135326 65894
rect 135390 65830 135668 65894
rect 135320 64126 135668 65830
rect 135320 64062 135326 64126
rect 135390 64062 135668 64126
rect 135320 62494 135668 64062
rect 135320 62430 135326 62494
rect 135390 62430 135668 62494
rect 134092 62123 134158 62124
rect 134092 62059 134093 62123
rect 134157 62059 134158 62123
rect 134092 62058 134158 62059
rect 133416 61478 133422 61542
rect 133486 61478 133492 61542
rect 133416 61472 133492 61478
rect 115872 61374 115878 61406
rect 115600 61336 115676 61342
rect 115877 61342 115878 61374
rect 115942 61374 115948 61406
rect 115942 61342 115943 61374
rect 115877 61341 115943 61342
rect 952 60934 1230 60998
rect 1294 60934 1300 60998
rect 21352 61270 21428 61276
rect 21352 61206 21358 61270
rect 21422 61206 21428 61270
rect 21352 60998 21428 61206
rect 21352 60966 21358 60998
rect 952 59230 1300 60934
rect 21357 60934 21358 60966
rect 21422 60966 21428 60998
rect 22168 61270 22244 61276
rect 22168 61206 22174 61270
rect 22238 61206 22244 61270
rect 22445 61270 22511 61271
rect 22445 61238 22446 61270
rect 22168 60998 22244 61206
rect 22168 60966 22174 60998
rect 21422 60934 21423 60966
rect 21357 60933 21423 60934
rect 22173 60934 22174 60966
rect 22238 60966 22244 60998
rect 22440 61206 22446 61238
rect 22510 61238 22511 61270
rect 114240 61270 114316 61276
rect 22510 61206 22516 61238
rect 22440 60998 22516 61206
rect 114240 61206 114246 61270
rect 114310 61206 114316 61270
rect 22238 60934 22239 60966
rect 22173 60933 22239 60934
rect 22440 60934 22446 60998
rect 22510 60934 22516 60998
rect 22440 60928 22516 60934
rect 109480 61134 109556 61140
rect 109480 61070 109486 61134
rect 109550 61070 109556 61134
rect 22173 60862 22239 60863
rect 22173 60830 22174 60862
rect 22168 60798 22174 60830
rect 22238 60830 22239 60862
rect 22576 60862 22652 60868
rect 22238 60798 22244 60830
rect 22168 60590 22244 60798
rect 22168 60526 22174 60590
rect 22238 60526 22244 60590
rect 22576 60798 22582 60862
rect 22646 60798 22652 60862
rect 109480 60862 109556 61070
rect 114240 60998 114316 61206
rect 114240 60966 114246 60998
rect 114245 60934 114246 60966
rect 114310 60966 114316 60998
rect 114648 61270 114724 61276
rect 114648 61206 114654 61270
rect 114718 61206 114724 61270
rect 115333 61270 115399 61271
rect 115333 61238 115334 61270
rect 114648 60998 114724 61206
rect 114648 60966 114654 60998
rect 114310 60934 114311 60966
rect 114245 60933 114311 60934
rect 114653 60934 114654 60966
rect 114718 60966 114724 60998
rect 115328 61206 115334 61238
rect 115398 61238 115399 61270
rect 115398 61206 115404 61238
rect 115328 60998 115404 61206
rect 114718 60934 114719 60966
rect 114653 60933 114719 60934
rect 115328 60934 115334 60998
rect 115398 60934 115404 60998
rect 115328 60928 115404 60934
rect 109480 60830 109486 60862
rect 22576 60590 22652 60798
rect 109485 60798 109486 60830
rect 109550 60830 109556 60862
rect 114240 60862 114316 60868
rect 109550 60798 109551 60830
rect 109485 60797 109551 60798
rect 114240 60798 114246 60862
rect 114310 60798 114316 60862
rect 22576 60558 22582 60590
rect 22168 60520 22244 60526
rect 22581 60526 22582 60558
rect 22646 60558 22652 60590
rect 114240 60590 114316 60798
rect 114240 60558 114246 60590
rect 22646 60526 22647 60558
rect 22581 60525 22647 60526
rect 114245 60526 114246 60558
rect 114310 60558 114316 60590
rect 114648 60862 114724 60868
rect 114648 60798 114654 60862
rect 114718 60798 114724 60862
rect 114648 60590 114724 60798
rect 114648 60558 114654 60590
rect 114310 60526 114311 60558
rect 114245 60525 114311 60526
rect 114653 60526 114654 60558
rect 114718 60558 114724 60590
rect 135320 60862 135668 62430
rect 135320 60798 135326 60862
rect 135390 60798 135668 60862
rect 114718 60526 114719 60558
rect 114653 60525 114719 60526
rect 21901 60454 21967 60455
rect 21901 60422 21902 60454
rect 21896 60390 21902 60422
rect 21966 60422 21967 60454
rect 22037 60454 22103 60455
rect 22037 60422 22038 60454
rect 21966 60390 21972 60422
rect 20808 60182 20884 60188
rect 20808 60118 20814 60182
rect 20878 60118 20884 60182
rect 20808 59910 20884 60118
rect 21896 60182 21972 60390
rect 21896 60118 21902 60182
rect 21966 60118 21972 60182
rect 21896 60112 21972 60118
rect 22032 60390 22038 60422
rect 22102 60422 22103 60454
rect 22445 60454 22511 60455
rect 22445 60422 22446 60454
rect 22102 60390 22108 60422
rect 22032 60182 22108 60390
rect 22032 60118 22038 60182
rect 22102 60118 22108 60182
rect 22032 60112 22108 60118
rect 22440 60390 22446 60422
rect 22510 60422 22511 60454
rect 114376 60454 114452 60460
rect 22510 60390 22516 60422
rect 22440 60182 22516 60390
rect 22440 60118 22446 60182
rect 22510 60118 22516 60182
rect 114376 60390 114382 60454
rect 114446 60390 114452 60454
rect 114653 60454 114719 60455
rect 114653 60422 114654 60454
rect 114376 60182 114452 60390
rect 114376 60150 114382 60182
rect 22440 60112 22516 60118
rect 114381 60118 114382 60150
rect 114446 60150 114452 60182
rect 114648 60390 114654 60422
rect 114718 60422 114719 60454
rect 115192 60454 115268 60460
rect 114718 60390 114724 60422
rect 114648 60182 114724 60390
rect 114446 60118 114447 60150
rect 114381 60117 114447 60118
rect 114648 60118 114654 60182
rect 114718 60118 114724 60182
rect 115192 60390 115198 60454
rect 115262 60390 115268 60454
rect 115192 60182 115268 60390
rect 115192 60150 115198 60182
rect 114648 60112 114724 60118
rect 115197 60118 115198 60150
rect 115262 60150 115268 60182
rect 115328 60454 115404 60460
rect 115328 60390 115334 60454
rect 115398 60390 115404 60454
rect 115328 60182 115404 60390
rect 115328 60150 115334 60182
rect 115262 60118 115263 60150
rect 115197 60117 115263 60118
rect 115333 60118 115334 60150
rect 115398 60150 115404 60182
rect 116008 60182 116084 60188
rect 115398 60118 115399 60150
rect 115333 60117 115399 60118
rect 116008 60118 116014 60182
rect 116078 60118 116084 60182
rect 20808 59878 20814 59910
rect 20813 59846 20814 59878
rect 20878 59878 20884 59910
rect 27336 59910 27412 59916
rect 20878 59846 20879 59878
rect 20813 59845 20879 59846
rect 27336 59846 27342 59910
rect 27406 59846 27412 59910
rect 109485 59910 109551 59911
rect 109485 59878 109486 59910
rect 20813 59774 20879 59775
rect 20813 59742 20814 59774
rect 20808 59710 20814 59742
rect 20878 59742 20879 59774
rect 21765 59774 21831 59775
rect 21765 59742 21766 59774
rect 20878 59710 20884 59742
rect 20808 59502 20884 59710
rect 20808 59438 20814 59502
rect 20878 59438 20884 59502
rect 20808 59432 20884 59438
rect 21760 59710 21766 59742
rect 21830 59742 21831 59774
rect 21830 59710 21836 59742
rect 21760 59502 21836 59710
rect 27336 59638 27412 59846
rect 27336 59606 27342 59638
rect 27341 59574 27342 59606
rect 27406 59606 27412 59638
rect 109480 59846 109486 59878
rect 109550 59878 109551 59910
rect 116008 59910 116084 60118
rect 116008 59878 116014 59910
rect 109550 59846 109556 59878
rect 109480 59638 109556 59846
rect 116013 59846 116014 59878
rect 116078 59878 116084 59910
rect 116078 59846 116079 59878
rect 116013 59845 116079 59846
rect 115469 59774 115535 59775
rect 115469 59742 115470 59774
rect 27406 59574 27407 59606
rect 27341 59573 27407 59574
rect 109480 59574 109486 59638
rect 109550 59574 109556 59638
rect 109480 59568 109556 59574
rect 115464 59710 115470 59742
rect 115534 59742 115535 59774
rect 116013 59774 116079 59775
rect 116013 59742 116014 59774
rect 115534 59710 115540 59742
rect 21760 59438 21766 59502
rect 21830 59438 21836 59502
rect 21760 59432 21836 59438
rect 115464 59502 115540 59710
rect 115464 59438 115470 59502
rect 115534 59438 115540 59502
rect 115464 59432 115540 59438
rect 116008 59710 116014 59742
rect 116078 59742 116079 59774
rect 116078 59710 116084 59742
rect 116008 59502 116084 59710
rect 116008 59438 116014 59502
rect 116078 59438 116084 59502
rect 116008 59432 116084 59438
rect 20813 59366 20879 59367
rect 20813 59334 20814 59366
rect 952 59166 1230 59230
rect 1294 59166 1300 59230
rect 952 57598 1300 59166
rect 20808 59302 20814 59334
rect 20878 59334 20879 59366
rect 22037 59366 22103 59367
rect 22037 59334 22038 59366
rect 20878 59302 20884 59334
rect 20808 59094 20884 59302
rect 20808 59030 20814 59094
rect 20878 59030 20884 59094
rect 20808 59024 20884 59030
rect 22032 59302 22038 59334
rect 22102 59334 22103 59366
rect 22445 59366 22511 59367
rect 22445 59334 22446 59366
rect 22102 59302 22108 59334
rect 22032 59094 22108 59302
rect 22032 59030 22038 59094
rect 22102 59030 22108 59094
rect 22032 59024 22108 59030
rect 22440 59302 22446 59334
rect 22510 59334 22511 59366
rect 114376 59366 114452 59372
rect 22510 59302 22516 59334
rect 22440 59094 22516 59302
rect 22440 59030 22446 59094
rect 22510 59030 22516 59094
rect 114376 59302 114382 59366
rect 114446 59302 114452 59366
rect 114376 59094 114452 59302
rect 114376 59062 114382 59094
rect 22440 59024 22516 59030
rect 114381 59030 114382 59062
rect 114446 59062 114452 59094
rect 114784 59366 114860 59372
rect 114784 59302 114790 59366
rect 114854 59302 114860 59366
rect 114784 59094 114860 59302
rect 114784 59062 114790 59094
rect 114446 59030 114447 59062
rect 114381 59029 114447 59030
rect 114789 59030 114790 59062
rect 114854 59062 114860 59094
rect 115872 59366 115948 59372
rect 115872 59302 115878 59366
rect 115942 59302 115948 59366
rect 115872 59094 115948 59302
rect 115872 59062 115878 59094
rect 114854 59030 114855 59062
rect 114789 59029 114855 59030
rect 115877 59030 115878 59062
rect 115942 59062 115948 59094
rect 135320 59230 135668 60798
rect 135320 59166 135326 59230
rect 135390 59166 135668 59230
rect 115942 59030 115943 59062
rect 115877 59029 115943 59030
rect 20808 58958 20884 58964
rect 20808 58894 20814 58958
rect 20878 58894 20884 58958
rect 21221 58958 21287 58959
rect 21221 58926 21222 58958
rect 20808 58686 20884 58894
rect 20808 58654 20814 58686
rect 20813 58622 20814 58654
rect 20878 58654 20884 58686
rect 21216 58894 21222 58926
rect 21286 58926 21287 58958
rect 22168 58958 22244 58964
rect 21286 58894 21292 58926
rect 21216 58686 21292 58894
rect 20878 58622 20879 58654
rect 20813 58621 20879 58622
rect 21216 58622 21222 58686
rect 21286 58622 21292 58686
rect 22168 58894 22174 58958
rect 22238 58894 22244 58958
rect 22168 58686 22244 58894
rect 22168 58654 22174 58686
rect 21216 58616 21292 58622
rect 22173 58622 22174 58654
rect 22238 58654 22244 58686
rect 22440 58958 22516 58964
rect 22440 58894 22446 58958
rect 22510 58894 22516 58958
rect 114381 58958 114447 58959
rect 114381 58926 114382 58958
rect 22440 58686 22516 58894
rect 114376 58894 114382 58926
rect 114446 58926 114447 58958
rect 114789 58958 114855 58959
rect 114789 58926 114790 58958
rect 114446 58894 114452 58926
rect 22440 58654 22446 58686
rect 22238 58622 22239 58654
rect 22173 58621 22239 58622
rect 22445 58622 22446 58654
rect 22510 58654 22516 58686
rect 27613 58686 27679 58687
rect 27613 58654 27614 58686
rect 22510 58622 22511 58654
rect 22445 58621 22511 58622
rect 27608 58622 27614 58654
rect 27678 58654 27679 58686
rect 109485 58686 109551 58687
rect 109485 58654 109486 58686
rect 27678 58622 27684 58654
rect 20813 58550 20879 58551
rect 20813 58518 20814 58550
rect 20808 58486 20814 58518
rect 20878 58518 20879 58550
rect 21357 58550 21423 58551
rect 21357 58518 21358 58550
rect 20878 58486 20884 58518
rect 20808 58278 20884 58486
rect 20808 58214 20814 58278
rect 20878 58214 20884 58278
rect 20808 58208 20884 58214
rect 21352 58486 21358 58518
rect 21422 58518 21423 58550
rect 21765 58550 21831 58551
rect 21765 58518 21766 58550
rect 21422 58486 21428 58518
rect 21352 58278 21428 58486
rect 21352 58214 21358 58278
rect 21422 58214 21428 58278
rect 21352 58208 21428 58214
rect 21760 58486 21766 58518
rect 21830 58518 21831 58550
rect 22173 58550 22239 58551
rect 22173 58518 22174 58550
rect 21830 58486 21836 58518
rect 21760 58278 21836 58486
rect 21760 58214 21766 58278
rect 21830 58214 21836 58278
rect 21760 58208 21836 58214
rect 22168 58486 22174 58518
rect 22238 58518 22239 58550
rect 22445 58550 22511 58551
rect 22445 58518 22446 58550
rect 22238 58486 22244 58518
rect 22168 58278 22244 58486
rect 22168 58214 22174 58278
rect 22238 58214 22244 58278
rect 22168 58208 22244 58214
rect 22440 58486 22446 58518
rect 22510 58518 22511 58550
rect 22510 58486 22516 58518
rect 22440 58278 22516 58486
rect 27608 58414 27684 58622
rect 27608 58350 27614 58414
rect 27678 58350 27684 58414
rect 27608 58344 27684 58350
rect 109480 58622 109486 58654
rect 109550 58654 109551 58686
rect 114376 58686 114452 58894
rect 109550 58622 109556 58654
rect 109480 58414 109556 58622
rect 114376 58622 114382 58686
rect 114446 58622 114452 58686
rect 114376 58616 114452 58622
rect 114784 58894 114790 58926
rect 114854 58926 114855 58958
rect 115464 58958 115540 58964
rect 114854 58894 114860 58926
rect 114784 58686 114860 58894
rect 114784 58622 114790 58686
rect 114854 58622 114860 58686
rect 115464 58894 115470 58958
rect 115534 58894 115540 58958
rect 115877 58958 115943 58959
rect 115877 58926 115878 58958
rect 115464 58686 115540 58894
rect 115464 58654 115470 58686
rect 114784 58616 114860 58622
rect 115469 58622 115470 58654
rect 115534 58654 115540 58686
rect 115872 58894 115878 58926
rect 115942 58926 115943 58958
rect 115942 58894 115948 58926
rect 115872 58686 115948 58894
rect 115534 58622 115535 58654
rect 115469 58621 115535 58622
rect 115872 58622 115878 58686
rect 115942 58622 115948 58686
rect 115872 58616 115948 58622
rect 114245 58550 114311 58551
rect 114245 58518 114246 58550
rect 109480 58350 109486 58414
rect 109550 58350 109556 58414
rect 109480 58344 109556 58350
rect 114240 58486 114246 58518
rect 114310 58518 114311 58550
rect 114784 58550 114860 58556
rect 114310 58486 114316 58518
rect 22440 58214 22446 58278
rect 22510 58214 22516 58278
rect 22440 58208 22516 58214
rect 114240 58278 114316 58486
rect 114240 58214 114246 58278
rect 114310 58214 114316 58278
rect 114784 58486 114790 58550
rect 114854 58486 114860 58550
rect 115061 58550 115127 58551
rect 115061 58518 115062 58550
rect 114784 58278 114860 58486
rect 114784 58246 114790 58278
rect 114240 58208 114316 58214
rect 114789 58214 114790 58246
rect 114854 58246 114860 58278
rect 115056 58486 115062 58518
rect 115126 58518 115127 58550
rect 115328 58550 115404 58556
rect 115126 58486 115132 58518
rect 115056 58278 115132 58486
rect 114854 58214 114855 58246
rect 114789 58213 114855 58214
rect 115056 58214 115062 58278
rect 115126 58214 115132 58278
rect 115328 58486 115334 58550
rect 115398 58486 115404 58550
rect 116013 58550 116079 58551
rect 116013 58518 116014 58550
rect 115328 58278 115404 58486
rect 115328 58246 115334 58278
rect 115056 58208 115132 58214
rect 115333 58214 115334 58246
rect 115398 58246 115404 58278
rect 116008 58486 116014 58518
rect 116078 58518 116079 58550
rect 116078 58486 116084 58518
rect 116008 58278 116084 58486
rect 115398 58214 115399 58246
rect 115333 58213 115399 58214
rect 116008 58214 116014 58278
rect 116078 58214 116084 58278
rect 116008 58208 116084 58214
rect 20944 58142 21020 58148
rect 20944 58078 20950 58142
rect 21014 58078 21020 58142
rect 20944 57870 21020 58078
rect 20944 57838 20950 57870
rect 20949 57806 20950 57838
rect 21014 57838 21020 57870
rect 21488 58142 21564 58148
rect 21488 58078 21494 58142
rect 21558 58078 21564 58142
rect 22037 58142 22103 58143
rect 22037 58110 22038 58142
rect 21488 57870 21564 58078
rect 21488 57838 21494 57870
rect 21014 57806 21015 57838
rect 20949 57805 21015 57806
rect 21493 57806 21494 57838
rect 21558 57838 21564 57870
rect 22032 58078 22038 58110
rect 22102 58110 22103 58142
rect 22445 58142 22511 58143
rect 22445 58110 22446 58142
rect 22102 58078 22108 58110
rect 22032 57870 22108 58078
rect 21558 57806 21559 57838
rect 21493 57805 21559 57806
rect 22032 57806 22038 57870
rect 22102 57806 22108 57870
rect 22032 57800 22108 57806
rect 22440 58078 22446 58110
rect 22510 58110 22511 58142
rect 114376 58142 114452 58148
rect 22510 58078 22516 58110
rect 22440 57870 22516 58078
rect 22440 57806 22446 57870
rect 22510 57806 22516 57870
rect 114376 58078 114382 58142
rect 114446 58078 114452 58142
rect 114789 58142 114855 58143
rect 114789 58110 114790 58142
rect 114376 57870 114452 58078
rect 114376 57838 114382 57870
rect 22440 57800 22516 57806
rect 114381 57806 114382 57838
rect 114446 57838 114452 57870
rect 114784 58078 114790 58110
rect 114854 58110 114855 58142
rect 115192 58142 115268 58148
rect 114854 58078 114860 58110
rect 114784 57870 114860 58078
rect 114446 57806 114447 57838
rect 114381 57805 114447 57806
rect 114784 57806 114790 57870
rect 114854 57806 114860 57870
rect 115192 58078 115198 58142
rect 115262 58078 115268 58142
rect 115192 57870 115268 58078
rect 115192 57838 115198 57870
rect 114784 57800 114860 57806
rect 115197 57806 115198 57838
rect 115262 57838 115268 57870
rect 115328 58142 115404 58148
rect 115328 58078 115334 58142
rect 115398 58078 115404 58142
rect 115328 57870 115404 58078
rect 115328 57838 115334 57870
rect 115262 57806 115263 57838
rect 115197 57805 115263 57806
rect 115333 57806 115334 57838
rect 115398 57838 115404 57870
rect 115872 58142 115948 58148
rect 115872 58078 115878 58142
rect 115942 58078 115948 58142
rect 115872 57870 115948 58078
rect 115872 57838 115878 57870
rect 115398 57806 115399 57838
rect 115333 57805 115399 57806
rect 115877 57806 115878 57838
rect 115942 57838 115948 57870
rect 115942 57806 115943 57838
rect 115877 57805 115943 57806
rect 20813 57734 20879 57735
rect 20813 57702 20814 57734
rect 952 57534 1230 57598
rect 1294 57534 1300 57598
rect 952 55966 1300 57534
rect 20808 57670 20814 57702
rect 20878 57702 20879 57734
rect 22173 57734 22239 57735
rect 22173 57702 22174 57734
rect 20878 57670 20884 57702
rect 20808 57462 20884 57670
rect 20808 57398 20814 57462
rect 20878 57398 20884 57462
rect 20808 57392 20884 57398
rect 22168 57670 22174 57702
rect 22238 57702 22239 57734
rect 22576 57734 22652 57740
rect 22238 57670 22244 57702
rect 22168 57462 22244 57670
rect 22168 57398 22174 57462
rect 22238 57398 22244 57462
rect 22576 57670 22582 57734
rect 22646 57670 22652 57734
rect 22576 57462 22652 57670
rect 22576 57430 22582 57462
rect 22168 57392 22244 57398
rect 22581 57398 22582 57430
rect 22646 57430 22652 57462
rect 114240 57734 114316 57740
rect 114240 57670 114246 57734
rect 114310 57670 114316 57734
rect 114240 57462 114316 57670
rect 114240 57430 114246 57462
rect 22646 57398 22647 57430
rect 22581 57397 22647 57398
rect 114245 57398 114246 57430
rect 114310 57430 114316 57462
rect 114648 57734 114724 57740
rect 114648 57670 114654 57734
rect 114718 57670 114724 57734
rect 114648 57462 114724 57670
rect 114648 57430 114654 57462
rect 114310 57398 114311 57430
rect 114245 57397 114311 57398
rect 114653 57398 114654 57430
rect 114718 57430 114724 57462
rect 115600 57734 115676 57740
rect 115600 57670 115606 57734
rect 115670 57670 115676 57734
rect 116013 57734 116079 57735
rect 116013 57702 116014 57734
rect 115600 57462 115676 57670
rect 115600 57430 115606 57462
rect 114718 57398 114719 57430
rect 114653 57397 114719 57398
rect 115605 57398 115606 57430
rect 115670 57430 115676 57462
rect 116008 57670 116014 57702
rect 116078 57702 116079 57734
rect 116078 57670 116084 57702
rect 116008 57462 116084 57670
rect 115670 57398 115671 57430
rect 115605 57397 115671 57398
rect 116008 57398 116014 57462
rect 116078 57398 116084 57462
rect 116008 57392 116084 57398
rect 135320 57598 135668 59166
rect 135320 57534 135326 57598
rect 135390 57534 135668 57598
rect 21216 57326 21292 57332
rect 21216 57262 21222 57326
rect 21286 57262 21292 57326
rect 21765 57326 21831 57327
rect 21765 57294 21766 57326
rect 21216 57054 21292 57262
rect 21216 57022 21222 57054
rect 21221 56990 21222 57022
rect 21286 57022 21292 57054
rect 21760 57262 21766 57294
rect 21830 57294 21831 57326
rect 22032 57326 22108 57332
rect 21830 57262 21836 57294
rect 21760 57054 21836 57262
rect 21286 56990 21287 57022
rect 21221 56989 21287 56990
rect 21760 56990 21766 57054
rect 21830 56990 21836 57054
rect 22032 57262 22038 57326
rect 22102 57262 22108 57326
rect 22032 57054 22108 57262
rect 22032 57022 22038 57054
rect 21760 56984 21836 56990
rect 22037 56990 22038 57022
rect 22102 57022 22108 57054
rect 22440 57326 22516 57332
rect 22440 57262 22446 57326
rect 22510 57262 22516 57326
rect 114245 57326 114311 57327
rect 114245 57294 114246 57326
rect 22440 57054 22516 57262
rect 22440 57022 22446 57054
rect 22102 56990 22103 57022
rect 22037 56989 22103 56990
rect 22445 56990 22446 57022
rect 22510 57022 22516 57054
rect 114240 57262 114246 57294
rect 114310 57294 114311 57326
rect 114653 57326 114719 57327
rect 114653 57294 114654 57326
rect 114310 57262 114316 57294
rect 114240 57054 114316 57262
rect 22510 56990 22511 57022
rect 22445 56989 22511 56990
rect 114240 56990 114246 57054
rect 114310 56990 114316 57054
rect 114240 56984 114316 56990
rect 114648 57262 114654 57294
rect 114718 57294 114719 57326
rect 115192 57326 115268 57332
rect 114718 57262 114724 57294
rect 114648 57054 114724 57262
rect 114648 56990 114654 57054
rect 114718 56990 114724 57054
rect 115192 57262 115198 57326
rect 115262 57262 115268 57326
rect 115605 57326 115671 57327
rect 115605 57294 115606 57326
rect 115192 57054 115268 57262
rect 115192 57022 115198 57054
rect 114648 56984 114724 56990
rect 115197 56990 115198 57022
rect 115262 57022 115268 57054
rect 115600 57262 115606 57294
rect 115670 57294 115671 57326
rect 115670 57262 115676 57294
rect 115600 57054 115676 57262
rect 115262 56990 115263 57022
rect 115197 56989 115263 56990
rect 115600 56990 115606 57054
rect 115670 56990 115676 57054
rect 115600 56984 115676 56990
rect 22037 56918 22103 56919
rect 22037 56886 22038 56918
rect 22032 56854 22038 56886
rect 22102 56886 22103 56918
rect 22445 56918 22511 56919
rect 22445 56886 22446 56918
rect 22102 56854 22108 56886
rect 22032 56646 22108 56854
rect 22032 56582 22038 56646
rect 22102 56582 22108 56646
rect 22032 56576 22108 56582
rect 22440 56854 22446 56886
rect 22510 56886 22511 56918
rect 114240 56918 114316 56924
rect 22510 56854 22516 56886
rect 22440 56646 22516 56854
rect 22440 56582 22446 56646
rect 22510 56582 22516 56646
rect 114240 56854 114246 56918
rect 114310 56854 114316 56918
rect 114789 56918 114855 56919
rect 114789 56886 114790 56918
rect 114240 56646 114316 56854
rect 114240 56614 114246 56646
rect 22440 56576 22516 56582
rect 114245 56582 114246 56614
rect 114310 56614 114316 56646
rect 114784 56854 114790 56886
rect 114854 56886 114855 56918
rect 114854 56854 114860 56886
rect 114784 56646 114860 56854
rect 114310 56582 114311 56614
rect 114245 56581 114311 56582
rect 114784 56582 114790 56646
rect 114854 56582 114860 56646
rect 114784 56576 114860 56582
rect 21352 56510 21428 56516
rect 21352 56446 21358 56510
rect 21422 56446 21428 56510
rect 20949 56238 21015 56239
rect 20949 56206 20950 56238
rect 952 55902 1230 55966
rect 1294 55902 1300 55966
rect 952 54198 1300 55902
rect 20944 56174 20950 56206
rect 21014 56206 21015 56238
rect 21352 56238 21428 56446
rect 21352 56206 21358 56238
rect 21014 56174 21020 56206
rect 20944 55966 21020 56174
rect 21357 56174 21358 56206
rect 21422 56206 21428 56238
rect 21624 56510 21700 56516
rect 21624 56446 21630 56510
rect 21694 56446 21700 56510
rect 22173 56510 22239 56511
rect 22173 56478 22174 56510
rect 21624 56238 21700 56446
rect 21624 56206 21630 56238
rect 21422 56174 21423 56206
rect 21357 56173 21423 56174
rect 21629 56174 21630 56206
rect 21694 56206 21700 56238
rect 22168 56446 22174 56478
rect 22238 56478 22239 56510
rect 22445 56510 22511 56511
rect 22445 56478 22446 56510
rect 22238 56446 22244 56478
rect 22168 56238 22244 56446
rect 21694 56174 21695 56206
rect 21629 56173 21695 56174
rect 22168 56174 22174 56238
rect 22238 56174 22244 56238
rect 22168 56168 22244 56174
rect 22440 56446 22446 56478
rect 22510 56478 22511 56510
rect 114245 56510 114311 56511
rect 114245 56478 114246 56510
rect 22510 56446 22516 56478
rect 22440 56238 22516 56446
rect 22440 56174 22446 56238
rect 22510 56174 22516 56238
rect 22440 56168 22516 56174
rect 114240 56446 114246 56478
rect 114310 56478 114311 56510
rect 114648 56510 114724 56516
rect 114310 56446 114316 56478
rect 114240 56238 114316 56446
rect 114240 56174 114246 56238
rect 114310 56174 114316 56238
rect 114648 56446 114654 56510
rect 114718 56446 114724 56510
rect 114648 56238 114724 56446
rect 114648 56206 114654 56238
rect 114240 56168 114316 56174
rect 114653 56174 114654 56206
rect 114718 56206 114724 56238
rect 115056 56510 115132 56516
rect 115056 56446 115062 56510
rect 115126 56446 115132 56510
rect 115056 56238 115132 56446
rect 115056 56206 115062 56238
rect 114718 56174 114719 56206
rect 114653 56173 114719 56174
rect 115061 56174 115062 56206
rect 115126 56206 115132 56238
rect 116013 56238 116079 56239
rect 116013 56206 116014 56238
rect 115126 56174 115127 56206
rect 115061 56173 115127 56174
rect 116008 56174 116014 56206
rect 116078 56206 116079 56238
rect 116078 56174 116084 56206
rect 109349 56102 109415 56103
rect 109349 56070 109350 56102
rect 109344 56038 109350 56070
rect 109414 56070 109415 56102
rect 115192 56102 115404 56108
rect 109414 56038 109420 56070
rect 20944 55902 20950 55966
rect 21014 55902 21020 55966
rect 27477 55966 27543 55967
rect 27477 55934 27478 55966
rect 20944 55896 21020 55902
rect 27472 55902 27478 55934
rect 27542 55934 27543 55966
rect 27542 55902 27548 55934
rect 20808 55830 20884 55836
rect 20808 55766 20814 55830
rect 20878 55766 20884 55830
rect 20808 55558 20884 55766
rect 20808 55526 20814 55558
rect 20813 55494 20814 55526
rect 20878 55526 20884 55558
rect 21488 55830 21564 55836
rect 21488 55766 21494 55830
rect 21558 55766 21564 55830
rect 21488 55558 21564 55766
rect 21488 55526 21494 55558
rect 20878 55494 20879 55526
rect 20813 55493 20879 55494
rect 21493 55494 21494 55526
rect 21558 55526 21564 55558
rect 27472 55558 27548 55902
rect 109344 55694 109420 56038
rect 115192 56038 115334 56102
rect 115398 56038 115404 56102
rect 115192 56032 115404 56038
rect 109485 55966 109551 55967
rect 109485 55934 109486 55966
rect 109344 55630 109350 55694
rect 109414 55630 109420 55694
rect 109344 55624 109420 55630
rect 109480 55902 109486 55934
rect 109550 55934 109551 55966
rect 115192 55966 115268 56032
rect 115192 55934 115198 55966
rect 109550 55902 109556 55934
rect 109480 55694 109556 55902
rect 115197 55902 115198 55934
rect 115262 55934 115268 55966
rect 116008 55966 116084 56174
rect 115262 55902 115263 55934
rect 115197 55901 115263 55902
rect 116008 55902 116014 55966
rect 116078 55902 116084 55966
rect 116008 55896 116084 55902
rect 135320 55966 135668 57534
rect 135320 55902 135326 55966
rect 135390 55902 135668 55966
rect 115333 55830 115399 55831
rect 115333 55798 115334 55830
rect 109480 55630 109486 55694
rect 109550 55630 109556 55694
rect 109480 55624 109556 55630
rect 115328 55766 115334 55798
rect 115398 55798 115399 55830
rect 116008 55830 116084 55836
rect 115398 55766 115404 55798
rect 21558 55494 21559 55526
rect 21493 55493 21559 55494
rect 27472 55494 27478 55558
rect 27542 55494 27548 55558
rect 27613 55558 27679 55559
rect 27613 55526 27614 55558
rect 27472 55488 27548 55494
rect 27608 55494 27614 55526
rect 27678 55526 27679 55558
rect 109485 55558 109551 55559
rect 109485 55526 109486 55558
rect 27678 55494 27684 55526
rect 20944 55422 21020 55428
rect 20944 55358 20950 55422
rect 21014 55358 21020 55422
rect 20944 55150 21020 55358
rect 27608 55286 27684 55494
rect 27608 55222 27614 55286
rect 27678 55222 27684 55286
rect 27608 55216 27684 55222
rect 109480 55494 109486 55526
rect 109550 55526 109551 55558
rect 115328 55558 115404 55766
rect 109550 55494 109556 55526
rect 109480 55286 109556 55494
rect 115328 55494 115334 55558
rect 115398 55494 115404 55558
rect 116008 55766 116014 55830
rect 116078 55766 116084 55830
rect 116008 55558 116084 55766
rect 116008 55526 116014 55558
rect 115328 55488 115404 55494
rect 116013 55494 116014 55526
rect 116078 55526 116084 55558
rect 116078 55494 116079 55526
rect 116013 55493 116079 55494
rect 116013 55422 116079 55423
rect 116013 55390 116014 55422
rect 109480 55222 109486 55286
rect 109550 55222 109556 55286
rect 109480 55216 109556 55222
rect 116008 55358 116014 55390
rect 116078 55390 116079 55422
rect 116078 55358 116084 55390
rect 20944 55118 20950 55150
rect 20949 55086 20950 55118
rect 21014 55118 21020 55150
rect 116008 55150 116084 55358
rect 21014 55086 21015 55118
rect 20949 55085 21015 55086
rect 116008 55086 116014 55150
rect 116078 55086 116084 55150
rect 116008 55080 116084 55086
rect 20813 55014 20879 55015
rect 20813 54982 20814 55014
rect 20808 54950 20814 54982
rect 20878 54982 20879 55014
rect 21624 55014 21700 55020
rect 20878 54950 20884 54982
rect 20808 54742 20884 54950
rect 20808 54678 20814 54742
rect 20878 54678 20884 54742
rect 21624 54950 21630 55014
rect 21694 54950 21700 55014
rect 21624 54742 21700 54950
rect 21624 54710 21630 54742
rect 20808 54672 20884 54678
rect 21629 54678 21630 54710
rect 21694 54710 21700 54742
rect 22032 55014 22108 55020
rect 22032 54950 22038 55014
rect 22102 54950 22108 55014
rect 22445 55014 22511 55015
rect 22445 54982 22446 55014
rect 22032 54742 22108 54950
rect 22032 54710 22038 54742
rect 21694 54678 21695 54710
rect 21629 54677 21695 54678
rect 22037 54678 22038 54710
rect 22102 54710 22108 54742
rect 22440 54950 22446 54982
rect 22510 54982 22511 55014
rect 114376 55014 114452 55020
rect 22510 54950 22516 54982
rect 22440 54742 22516 54950
rect 22102 54678 22103 54710
rect 22037 54677 22103 54678
rect 22440 54678 22446 54742
rect 22510 54678 22516 54742
rect 114376 54950 114382 55014
rect 114446 54950 114452 55014
rect 114376 54742 114452 54950
rect 114376 54710 114382 54742
rect 22440 54672 22516 54678
rect 114381 54678 114382 54710
rect 114446 54710 114452 54742
rect 114784 55014 114860 55020
rect 114784 54950 114790 55014
rect 114854 54950 114860 55014
rect 115197 55014 115263 55015
rect 115197 54982 115198 55014
rect 114784 54742 114860 54950
rect 114784 54710 114790 54742
rect 114446 54678 114447 54710
rect 114381 54677 114447 54678
rect 114789 54678 114790 54710
rect 114854 54710 114860 54742
rect 115192 54950 115198 54982
rect 115262 54982 115263 55014
rect 115328 55014 115404 55020
rect 115262 54950 115268 54982
rect 115192 54742 115268 54950
rect 114854 54678 114855 54710
rect 114789 54677 114855 54678
rect 115192 54678 115198 54742
rect 115262 54678 115268 54742
rect 115328 54950 115334 55014
rect 115398 54950 115404 55014
rect 115877 55014 115943 55015
rect 115877 54982 115878 55014
rect 115328 54742 115404 54950
rect 115328 54710 115334 54742
rect 115192 54672 115268 54678
rect 115333 54678 115334 54710
rect 115398 54710 115404 54742
rect 115872 54950 115878 54982
rect 115942 54982 115943 55014
rect 115942 54950 115948 54982
rect 115872 54742 115948 54950
rect 115398 54678 115399 54710
rect 115333 54677 115399 54678
rect 115872 54678 115878 54742
rect 115942 54678 115948 54742
rect 115872 54672 115948 54678
rect 20944 54606 21020 54612
rect 20944 54542 20950 54606
rect 21014 54542 21020 54606
rect 20944 54334 21020 54542
rect 20944 54302 20950 54334
rect 20949 54270 20950 54302
rect 21014 54302 21020 54334
rect 21352 54606 21428 54612
rect 21352 54542 21358 54606
rect 21422 54542 21428 54606
rect 21352 54334 21428 54542
rect 21352 54302 21358 54334
rect 21014 54270 21015 54302
rect 20949 54269 21015 54270
rect 21357 54270 21358 54302
rect 21422 54302 21428 54334
rect 21488 54606 21564 54612
rect 21488 54542 21494 54606
rect 21558 54542 21564 54606
rect 21488 54334 21564 54542
rect 21488 54302 21494 54334
rect 21422 54270 21423 54302
rect 21357 54269 21423 54270
rect 21493 54270 21494 54302
rect 21558 54302 21564 54334
rect 22168 54606 22244 54612
rect 22168 54542 22174 54606
rect 22238 54542 22244 54606
rect 22581 54606 22647 54607
rect 22581 54574 22582 54606
rect 22168 54334 22244 54542
rect 22168 54302 22174 54334
rect 21558 54270 21559 54302
rect 21493 54269 21559 54270
rect 22173 54270 22174 54302
rect 22238 54302 22244 54334
rect 22576 54542 22582 54574
rect 22646 54574 22647 54606
rect 114240 54606 114316 54612
rect 22646 54542 22652 54574
rect 22576 54334 22652 54542
rect 22238 54270 22239 54302
rect 22173 54269 22239 54270
rect 22576 54270 22582 54334
rect 22646 54270 22652 54334
rect 114240 54542 114246 54606
rect 114310 54542 114316 54606
rect 114789 54606 114855 54607
rect 114789 54574 114790 54606
rect 114240 54334 114316 54542
rect 114240 54302 114246 54334
rect 22576 54264 22652 54270
rect 114245 54270 114246 54302
rect 114310 54302 114316 54334
rect 114784 54542 114790 54574
rect 114854 54574 114855 54606
rect 115464 54606 115540 54612
rect 114854 54542 114860 54574
rect 114784 54334 114860 54542
rect 114310 54270 114311 54302
rect 114245 54269 114311 54270
rect 114784 54270 114790 54334
rect 114854 54270 114860 54334
rect 115464 54542 115470 54606
rect 115534 54542 115540 54606
rect 115464 54334 115540 54542
rect 115464 54302 115470 54334
rect 114784 54264 114860 54270
rect 115469 54270 115470 54302
rect 115534 54302 115540 54334
rect 116008 54606 116084 54612
rect 116008 54542 116014 54606
rect 116078 54542 116084 54606
rect 116008 54334 116084 54542
rect 116008 54302 116014 54334
rect 115534 54270 115535 54302
rect 115469 54269 115535 54270
rect 116013 54270 116014 54302
rect 116078 54302 116084 54334
rect 116078 54270 116079 54302
rect 116013 54269 116079 54270
rect 952 54134 1230 54198
rect 1294 54134 1300 54198
rect 20813 54198 20879 54199
rect 20813 54166 20814 54198
rect 952 52566 1300 54134
rect 20808 54134 20814 54166
rect 20878 54166 20879 54198
rect 21765 54198 21831 54199
rect 21765 54166 21766 54198
rect 20878 54134 20884 54166
rect 20808 53926 20884 54134
rect 20808 53862 20814 53926
rect 20878 53862 20884 53926
rect 20808 53856 20884 53862
rect 21760 54134 21766 54166
rect 21830 54166 21831 54198
rect 22173 54198 22239 54199
rect 22173 54166 22174 54198
rect 21830 54134 21836 54166
rect 21760 53926 21836 54134
rect 21760 53862 21766 53926
rect 21830 53862 21836 53926
rect 21760 53856 21836 53862
rect 22168 54134 22174 54166
rect 22238 54166 22239 54198
rect 22440 54198 22516 54204
rect 22238 54134 22244 54166
rect 22168 53926 22244 54134
rect 22168 53862 22174 53926
rect 22238 53862 22244 53926
rect 22440 54134 22446 54198
rect 22510 54134 22516 54198
rect 22440 53926 22516 54134
rect 22440 53894 22446 53926
rect 22168 53856 22244 53862
rect 22445 53862 22446 53894
rect 22510 53894 22516 53926
rect 114376 54198 114452 54204
rect 114376 54134 114382 54198
rect 114446 54134 114452 54198
rect 114376 53926 114452 54134
rect 114376 53894 114382 53926
rect 22510 53862 22511 53894
rect 22445 53861 22511 53862
rect 114381 53862 114382 53894
rect 114446 53894 114452 53926
rect 114784 54198 114860 54204
rect 114784 54134 114790 54198
rect 114854 54134 114860 54198
rect 114784 53926 114860 54134
rect 114784 53894 114790 53926
rect 114446 53862 114447 53894
rect 114381 53861 114447 53862
rect 114789 53862 114790 53894
rect 114854 53894 114860 53926
rect 115192 54198 115268 54204
rect 115192 54134 115198 54198
rect 115262 54134 115268 54198
rect 115192 53926 115268 54134
rect 115192 53894 115198 53926
rect 114854 53862 114855 53894
rect 114789 53861 114855 53862
rect 115197 53862 115198 53894
rect 115262 53894 115268 53926
rect 115328 54198 115404 54204
rect 115328 54134 115334 54198
rect 115398 54134 115404 54198
rect 116013 54198 116079 54199
rect 116013 54166 116014 54198
rect 115328 53926 115404 54134
rect 115328 53894 115334 53926
rect 115262 53862 115263 53894
rect 115197 53861 115263 53862
rect 115333 53862 115334 53894
rect 115398 53894 115404 53926
rect 116008 54134 116014 54166
rect 116078 54166 116079 54198
rect 116078 54134 116084 54166
rect 116008 53926 116084 54134
rect 115398 53862 115399 53894
rect 115333 53861 115399 53862
rect 116008 53862 116014 53926
rect 116078 53862 116084 53926
rect 116008 53856 116084 53862
rect 135320 54062 135668 55902
rect 135320 53998 135326 54062
rect 135390 53998 135668 54062
rect 20813 53790 20879 53791
rect 20813 53758 20814 53790
rect 20808 53726 20814 53758
rect 20878 53758 20879 53790
rect 21624 53790 21700 53796
rect 20878 53726 20884 53758
rect 20808 53518 20884 53726
rect 20808 53454 20814 53518
rect 20878 53454 20884 53518
rect 21624 53726 21630 53790
rect 21694 53726 21700 53790
rect 22037 53790 22103 53791
rect 22037 53758 22038 53790
rect 21624 53518 21700 53726
rect 21624 53486 21630 53518
rect 20808 53448 20884 53454
rect 21629 53454 21630 53486
rect 21694 53486 21700 53518
rect 22032 53726 22038 53758
rect 22102 53758 22103 53790
rect 22445 53790 22511 53791
rect 22445 53758 22446 53790
rect 22102 53726 22108 53758
rect 22032 53518 22108 53726
rect 21694 53454 21695 53486
rect 21629 53453 21695 53454
rect 22032 53454 22038 53518
rect 22102 53454 22108 53518
rect 22032 53448 22108 53454
rect 22440 53726 22446 53758
rect 22510 53758 22511 53790
rect 114381 53790 114447 53791
rect 114381 53758 114382 53790
rect 22510 53726 22516 53758
rect 22440 53518 22516 53726
rect 22440 53454 22446 53518
rect 22510 53454 22516 53518
rect 22440 53448 22516 53454
rect 114376 53726 114382 53758
rect 114446 53758 114447 53790
rect 114789 53790 114855 53791
rect 114789 53758 114790 53790
rect 114446 53726 114452 53758
rect 114376 53518 114452 53726
rect 114376 53454 114382 53518
rect 114446 53454 114452 53518
rect 114376 53448 114452 53454
rect 114784 53726 114790 53758
rect 114854 53758 114855 53790
rect 115872 53790 115948 53796
rect 114854 53726 114860 53758
rect 114784 53518 114860 53726
rect 114784 53454 114790 53518
rect 114854 53454 114860 53518
rect 115872 53726 115878 53790
rect 115942 53726 115948 53790
rect 115872 53518 115948 53726
rect 115872 53486 115878 53518
rect 114784 53448 114860 53454
rect 115877 53454 115878 53486
rect 115942 53486 115948 53518
rect 115942 53454 115943 53486
rect 115877 53453 115943 53454
rect 21357 53382 21423 53383
rect 21357 53350 21358 53382
rect 21352 53318 21358 53350
rect 21422 53350 21423 53382
rect 21493 53382 21559 53383
rect 21493 53350 21494 53382
rect 21422 53318 21428 53350
rect 21352 53110 21428 53318
rect 21352 53046 21358 53110
rect 21422 53046 21428 53110
rect 21352 53040 21428 53046
rect 21488 53318 21494 53350
rect 21558 53350 21559 53382
rect 22168 53382 22244 53388
rect 21558 53318 21564 53350
rect 21488 53110 21564 53318
rect 21488 53046 21494 53110
rect 21558 53046 21564 53110
rect 22168 53318 22174 53382
rect 22238 53318 22244 53382
rect 22445 53382 22511 53383
rect 22445 53350 22446 53382
rect 22168 53110 22244 53318
rect 22168 53078 22174 53110
rect 21488 53040 21564 53046
rect 22173 53046 22174 53078
rect 22238 53078 22244 53110
rect 22440 53318 22446 53350
rect 22510 53350 22511 53382
rect 114240 53382 114316 53388
rect 22510 53318 22516 53350
rect 22440 53110 22516 53318
rect 22238 53046 22239 53078
rect 22173 53045 22239 53046
rect 22440 53046 22446 53110
rect 22510 53046 22516 53110
rect 114240 53318 114246 53382
rect 114310 53318 114316 53382
rect 114653 53382 114719 53383
rect 114653 53350 114654 53382
rect 114240 53110 114316 53318
rect 114240 53078 114246 53110
rect 22440 53040 22516 53046
rect 114245 53046 114246 53078
rect 114310 53078 114316 53110
rect 114648 53318 114654 53350
rect 114718 53350 114719 53382
rect 115469 53382 115535 53383
rect 115469 53350 115470 53382
rect 114718 53318 114724 53350
rect 114648 53110 114724 53318
rect 114310 53046 114311 53078
rect 114245 53045 114311 53046
rect 114648 53046 114654 53110
rect 114718 53046 114724 53110
rect 114648 53040 114724 53046
rect 115464 53318 115470 53350
rect 115534 53350 115535 53382
rect 115534 53318 115540 53350
rect 115464 53110 115540 53318
rect 115464 53046 115470 53110
rect 115534 53046 115540 53110
rect 115464 53040 115540 53046
rect 20949 52974 21015 52975
rect 20949 52942 20950 52974
rect 20944 52910 20950 52942
rect 21014 52942 21015 52974
rect 21216 52974 21292 52980
rect 21014 52910 21020 52942
rect 20944 52702 21020 52910
rect 20944 52638 20950 52702
rect 21014 52638 21020 52702
rect 21216 52910 21222 52974
rect 21286 52910 21292 52974
rect 21765 52974 21831 52975
rect 21765 52942 21766 52974
rect 21216 52702 21292 52910
rect 21216 52670 21222 52702
rect 20944 52632 21020 52638
rect 21221 52638 21222 52670
rect 21286 52670 21292 52702
rect 21760 52910 21766 52942
rect 21830 52942 21831 52974
rect 22173 52974 22239 52975
rect 22173 52942 22174 52974
rect 21830 52910 21836 52942
rect 21760 52702 21836 52910
rect 21286 52638 21287 52670
rect 21221 52637 21287 52638
rect 21760 52638 21766 52702
rect 21830 52638 21836 52702
rect 21760 52632 21836 52638
rect 22168 52910 22174 52942
rect 22238 52942 22239 52974
rect 22576 52974 22652 52980
rect 22238 52910 22244 52942
rect 22168 52702 22244 52910
rect 22168 52638 22174 52702
rect 22238 52638 22244 52702
rect 22576 52910 22582 52974
rect 22646 52910 22652 52974
rect 114245 52974 114311 52975
rect 114245 52942 114246 52974
rect 22576 52702 22652 52910
rect 22576 52670 22582 52702
rect 22168 52632 22244 52638
rect 22581 52638 22582 52670
rect 22646 52670 22652 52702
rect 114240 52910 114246 52942
rect 114310 52942 114311 52974
rect 114784 52974 114860 52980
rect 114310 52910 114316 52942
rect 114240 52702 114316 52910
rect 22646 52638 22647 52670
rect 22581 52637 22647 52638
rect 114240 52638 114246 52702
rect 114310 52638 114316 52702
rect 114784 52910 114790 52974
rect 114854 52910 114860 52974
rect 114784 52702 114860 52910
rect 114784 52670 114790 52702
rect 114240 52632 114316 52638
rect 114789 52638 114790 52670
rect 114854 52670 114860 52702
rect 115192 52974 115268 52980
rect 115192 52910 115198 52974
rect 115262 52910 115268 52974
rect 115192 52702 115268 52910
rect 115192 52670 115198 52702
rect 114854 52638 114855 52670
rect 114789 52637 114855 52638
rect 115197 52638 115198 52670
rect 115262 52670 115268 52702
rect 115600 52974 115676 52980
rect 115600 52910 115606 52974
rect 115670 52910 115676 52974
rect 115600 52702 115676 52910
rect 115600 52670 115606 52702
rect 115262 52638 115263 52670
rect 115197 52637 115263 52638
rect 115605 52638 115606 52670
rect 115670 52670 115676 52702
rect 115872 52974 115948 52980
rect 115872 52910 115878 52974
rect 115942 52910 115948 52974
rect 115872 52702 115948 52910
rect 115872 52670 115878 52702
rect 115670 52638 115671 52670
rect 115605 52637 115671 52638
rect 115877 52638 115878 52670
rect 115942 52670 115948 52702
rect 115942 52638 115943 52670
rect 115877 52637 115943 52638
rect 952 52502 1230 52566
rect 1294 52502 1300 52566
rect 952 50934 1300 52502
rect 22168 52566 22244 52572
rect 22168 52502 22174 52566
rect 22238 52502 22244 52566
rect 22445 52566 22511 52567
rect 22445 52534 22446 52566
rect 20813 52294 20879 52295
rect 20813 52262 20814 52294
rect 20808 52230 20814 52262
rect 20878 52262 20879 52294
rect 22168 52294 22244 52502
rect 22168 52262 22174 52294
rect 20878 52230 20884 52262
rect 20808 52022 20884 52230
rect 22173 52230 22174 52262
rect 22238 52262 22244 52294
rect 22440 52502 22446 52534
rect 22510 52534 22511 52566
rect 114381 52566 114447 52567
rect 114381 52534 114382 52566
rect 22510 52502 22516 52534
rect 22440 52294 22516 52502
rect 114376 52502 114382 52534
rect 114446 52534 114447 52566
rect 114789 52566 114855 52567
rect 114789 52534 114790 52566
rect 114446 52502 114452 52534
rect 27477 52430 27543 52431
rect 27477 52398 27478 52430
rect 22238 52230 22239 52262
rect 22173 52229 22239 52230
rect 22440 52230 22446 52294
rect 22510 52230 22516 52294
rect 22440 52224 22516 52230
rect 27472 52366 27478 52398
rect 27542 52398 27543 52430
rect 27542 52366 27548 52398
rect 22173 52158 22239 52159
rect 22173 52126 22174 52158
rect 20808 51958 20814 52022
rect 20878 51958 20884 52022
rect 20808 51952 20884 51958
rect 22168 52094 22174 52126
rect 22238 52126 22239 52158
rect 22576 52158 22652 52164
rect 22238 52094 22244 52126
rect 22168 51886 22244 52094
rect 22168 51822 22174 51886
rect 22238 51822 22244 51886
rect 22576 52094 22582 52158
rect 22646 52094 22652 52158
rect 22576 51886 22652 52094
rect 27472 52158 27548 52366
rect 114376 52294 114452 52502
rect 114376 52230 114382 52294
rect 114446 52230 114452 52294
rect 114376 52224 114452 52230
rect 114784 52502 114790 52534
rect 114854 52534 114855 52566
rect 115197 52566 115263 52567
rect 115197 52534 115198 52566
rect 114854 52502 114860 52534
rect 114784 52294 114860 52502
rect 114784 52230 114790 52294
rect 114854 52230 114860 52294
rect 114784 52224 114860 52230
rect 115192 52502 115198 52534
rect 115262 52534 115263 52566
rect 115262 52502 115268 52534
rect 115192 52294 115268 52502
rect 135320 52430 135668 53998
rect 135320 52366 135326 52430
rect 135390 52366 135668 52430
rect 115192 52230 115198 52294
rect 115262 52230 115268 52294
rect 116013 52294 116079 52295
rect 116013 52262 116014 52294
rect 115192 52224 115268 52230
rect 116008 52230 116014 52262
rect 116078 52262 116079 52294
rect 116078 52230 116084 52262
rect 27472 52094 27478 52158
rect 27542 52094 27548 52158
rect 27472 52088 27548 52094
rect 114240 52158 114316 52164
rect 114240 52094 114246 52158
rect 114310 52094 114316 52158
rect 22576 51854 22582 51886
rect 22168 51816 22244 51822
rect 22581 51822 22582 51854
rect 22646 51854 22652 51886
rect 114240 51886 114316 52094
rect 114240 51854 114246 51886
rect 22646 51822 22647 51854
rect 22581 51821 22647 51822
rect 114245 51822 114246 51854
rect 114310 51854 114316 51886
rect 114648 52158 114724 52164
rect 114648 52094 114654 52158
rect 114718 52094 114724 52158
rect 114648 51886 114724 52094
rect 116008 52022 116084 52230
rect 116008 51958 116014 52022
rect 116078 51958 116084 52022
rect 116008 51952 116084 51958
rect 114648 51854 114654 51886
rect 114310 51822 114311 51854
rect 114245 51821 114311 51822
rect 114653 51822 114654 51854
rect 114718 51854 114724 51886
rect 114718 51822 114719 51854
rect 114653 51821 114719 51822
rect 21760 51750 21836 51756
rect 21760 51686 21766 51750
rect 21830 51686 21836 51750
rect 20813 51478 20879 51479
rect 20813 51446 20814 51478
rect 20808 51414 20814 51446
rect 20878 51446 20879 51478
rect 21760 51478 21836 51686
rect 21760 51446 21766 51478
rect 20878 51414 20884 51446
rect 20808 51206 20884 51414
rect 21765 51414 21766 51446
rect 21830 51446 21836 51478
rect 115192 51750 115268 51756
rect 115192 51686 115198 51750
rect 115262 51686 115268 51750
rect 115192 51478 115268 51686
rect 115192 51446 115198 51478
rect 21830 51414 21831 51446
rect 21765 51413 21831 51414
rect 115197 51414 115198 51446
rect 115262 51446 115268 51478
rect 115877 51478 115943 51479
rect 115877 51446 115878 51478
rect 115262 51414 115263 51446
rect 115197 51413 115263 51414
rect 115872 51414 115878 51446
rect 115942 51446 115943 51478
rect 115942 51414 115948 51446
rect 27341 51342 27407 51343
rect 27341 51310 27342 51342
rect 20808 51142 20814 51206
rect 20878 51142 20884 51206
rect 20808 51136 20884 51142
rect 27336 51278 27342 51310
rect 27406 51310 27407 51342
rect 27406 51278 27412 51310
rect 20813 51070 20879 51071
rect 20813 51038 20814 51070
rect 952 50870 1230 50934
rect 1294 50870 1300 50934
rect 952 49030 1300 50870
rect 20808 51006 20814 51038
rect 20878 51038 20879 51070
rect 21357 51070 21423 51071
rect 21357 51038 21358 51070
rect 20878 51006 20884 51038
rect 20808 50798 20884 51006
rect 20808 50734 20814 50798
rect 20878 50734 20884 50798
rect 20808 50728 20884 50734
rect 21352 51006 21358 51038
rect 21422 51038 21423 51070
rect 21896 51070 21972 51076
rect 21422 51006 21428 51038
rect 21352 50798 21428 51006
rect 21352 50734 21358 50798
rect 21422 50734 21428 50798
rect 21896 51006 21902 51070
rect 21966 51006 21972 51070
rect 22173 51070 22239 51071
rect 22173 51038 22174 51070
rect 21896 50798 21972 51006
rect 21896 50766 21902 50798
rect 21352 50728 21428 50734
rect 21901 50734 21902 50766
rect 21966 50766 21972 50798
rect 22168 51006 22174 51038
rect 22238 51038 22239 51070
rect 22576 51070 22652 51076
rect 22238 51006 22244 51038
rect 22168 50798 22244 51006
rect 21966 50734 21967 50766
rect 21901 50733 21967 50734
rect 22168 50734 22174 50798
rect 22238 50734 22244 50798
rect 22576 51006 22582 51070
rect 22646 51006 22652 51070
rect 22576 50798 22652 51006
rect 27336 51070 27412 51278
rect 115872 51206 115948 51414
rect 115872 51142 115878 51206
rect 115942 51142 115948 51206
rect 115872 51136 115948 51142
rect 27336 51006 27342 51070
rect 27406 51006 27412 51070
rect 27336 51000 27412 51006
rect 114240 51070 114316 51076
rect 114240 51006 114246 51070
rect 114310 51006 114316 51070
rect 22576 50766 22582 50798
rect 22168 50728 22244 50734
rect 22581 50734 22582 50766
rect 22646 50766 22652 50798
rect 114240 50798 114316 51006
rect 114240 50766 114246 50798
rect 22646 50734 22647 50766
rect 22581 50733 22647 50734
rect 114245 50734 114246 50766
rect 114310 50766 114316 50798
rect 114648 51070 114724 51076
rect 114648 51006 114654 51070
rect 114718 51006 114724 51070
rect 114648 50798 114724 51006
rect 114648 50766 114654 50798
rect 114310 50734 114311 50766
rect 114245 50733 114311 50734
rect 114653 50734 114654 50766
rect 114718 50766 114724 50798
rect 115056 51070 115132 51076
rect 115056 51006 115062 51070
rect 115126 51006 115132 51070
rect 115469 51070 115535 51071
rect 115469 51038 115470 51070
rect 115056 50798 115132 51006
rect 115056 50766 115062 50798
rect 114718 50734 114719 50766
rect 114653 50733 114719 50734
rect 115061 50734 115062 50766
rect 115126 50766 115132 50798
rect 115464 51006 115470 51038
rect 115534 51038 115535 51070
rect 116013 51070 116079 51071
rect 116013 51038 116014 51070
rect 115534 51006 115540 51038
rect 115464 50798 115540 51006
rect 115126 50734 115127 50766
rect 115061 50733 115127 50734
rect 115464 50734 115470 50798
rect 115534 50734 115540 50798
rect 115464 50728 115540 50734
rect 116008 51006 116014 51038
rect 116078 51038 116079 51070
rect 116078 51006 116084 51038
rect 116008 50798 116084 51006
rect 116008 50734 116014 50798
rect 116078 50734 116084 50798
rect 116008 50728 116084 50734
rect 135320 50798 135668 52366
rect 135320 50734 135326 50798
rect 135390 50734 135668 50798
rect 20813 50662 20879 50663
rect 20813 50630 20814 50662
rect 20808 50598 20814 50630
rect 20878 50630 20879 50662
rect 21901 50662 21967 50663
rect 21901 50630 21902 50662
rect 20878 50598 20884 50630
rect 20808 50390 20884 50598
rect 20808 50326 20814 50390
rect 20878 50326 20884 50390
rect 20808 50320 20884 50326
rect 21896 50598 21902 50630
rect 21966 50630 21967 50662
rect 22032 50662 22108 50668
rect 21966 50598 21972 50630
rect 21896 50390 21972 50598
rect 21896 50326 21902 50390
rect 21966 50326 21972 50390
rect 22032 50598 22038 50662
rect 22102 50598 22108 50662
rect 22445 50662 22511 50663
rect 22445 50630 22446 50662
rect 22032 50390 22108 50598
rect 22032 50358 22038 50390
rect 21896 50320 21972 50326
rect 22037 50326 22038 50358
rect 22102 50358 22108 50390
rect 22440 50598 22446 50630
rect 22510 50630 22511 50662
rect 114381 50662 114447 50663
rect 114381 50630 114382 50662
rect 22510 50598 22516 50630
rect 22440 50390 22516 50598
rect 22102 50326 22103 50358
rect 22037 50325 22103 50326
rect 22440 50326 22446 50390
rect 22510 50326 22516 50390
rect 22440 50320 22516 50326
rect 114376 50598 114382 50630
rect 114446 50630 114447 50662
rect 114784 50662 114860 50668
rect 114446 50598 114452 50630
rect 114376 50390 114452 50598
rect 114376 50326 114382 50390
rect 114446 50326 114452 50390
rect 114784 50598 114790 50662
rect 114854 50598 114860 50662
rect 114784 50390 114860 50598
rect 114784 50358 114790 50390
rect 114376 50320 114452 50326
rect 114789 50326 114790 50358
rect 114854 50358 114860 50390
rect 115872 50662 115948 50668
rect 115872 50598 115878 50662
rect 115942 50598 115948 50662
rect 115872 50390 115948 50598
rect 115872 50358 115878 50390
rect 114854 50326 114855 50358
rect 114789 50325 114855 50326
rect 115877 50326 115878 50358
rect 115942 50358 115948 50390
rect 115942 50326 115943 50358
rect 115877 50325 115943 50326
rect 20949 50254 21015 50255
rect 20949 50222 20950 50254
rect 20944 50190 20950 50222
rect 21014 50222 21015 50254
rect 21221 50254 21287 50255
rect 21221 50222 21222 50254
rect 21014 50190 21020 50222
rect 20944 49982 21020 50190
rect 20944 49918 20950 49982
rect 21014 49918 21020 49982
rect 20944 49912 21020 49918
rect 21216 50190 21222 50222
rect 21286 50222 21287 50254
rect 21488 50254 21564 50260
rect 21286 50190 21292 50222
rect 21216 49982 21292 50190
rect 21216 49918 21222 49982
rect 21286 49918 21292 49982
rect 21488 50190 21494 50254
rect 21558 50190 21564 50254
rect 21488 49982 21564 50190
rect 21488 49950 21494 49982
rect 21216 49912 21292 49918
rect 21493 49918 21494 49950
rect 21558 49950 21564 49982
rect 22168 50254 22244 50260
rect 22168 50190 22174 50254
rect 22238 50190 22244 50254
rect 22581 50254 22647 50255
rect 22581 50222 22582 50254
rect 22168 49982 22244 50190
rect 22168 49950 22174 49982
rect 21558 49918 21559 49950
rect 21493 49917 21559 49918
rect 22173 49918 22174 49950
rect 22238 49950 22244 49982
rect 22576 50190 22582 50222
rect 22646 50222 22647 50254
rect 114240 50254 114316 50260
rect 22646 50190 22652 50222
rect 22576 49982 22652 50190
rect 22238 49918 22239 49950
rect 22173 49917 22239 49918
rect 22576 49918 22582 49982
rect 22646 49918 22652 49982
rect 114240 50190 114246 50254
rect 114310 50190 114316 50254
rect 114789 50254 114855 50255
rect 114789 50222 114790 50254
rect 114240 49982 114316 50190
rect 114240 49950 114246 49982
rect 22576 49912 22652 49918
rect 114245 49918 114246 49950
rect 114310 49950 114316 49982
rect 114784 50190 114790 50222
rect 114854 50222 114855 50254
rect 115605 50254 115671 50255
rect 115605 50222 115606 50254
rect 114854 50190 114860 50222
rect 114784 49982 114860 50190
rect 114310 49918 114311 49950
rect 114245 49917 114311 49918
rect 114784 49918 114790 49982
rect 114854 49918 114860 49982
rect 114784 49912 114860 49918
rect 115600 50190 115606 50222
rect 115670 50222 115671 50254
rect 115877 50254 115943 50255
rect 115877 50222 115878 50254
rect 115670 50190 115676 50222
rect 115600 49982 115676 50190
rect 115600 49918 115606 49982
rect 115670 49918 115676 49982
rect 115600 49912 115676 49918
rect 115872 50190 115878 50222
rect 115942 50222 115943 50254
rect 115942 50190 115948 50222
rect 115872 49982 115948 50190
rect 115872 49918 115878 49982
rect 115942 49918 115948 49982
rect 115872 49912 115948 49918
rect 20808 49846 20884 49852
rect 20808 49782 20814 49846
rect 20878 49782 20884 49846
rect 21765 49846 21831 49847
rect 21765 49814 21766 49846
rect 20808 49574 20884 49782
rect 20808 49542 20814 49574
rect 20813 49510 20814 49542
rect 20878 49542 20884 49574
rect 21760 49782 21766 49814
rect 21830 49814 21831 49846
rect 22173 49846 22239 49847
rect 22173 49814 22174 49846
rect 21830 49782 21836 49814
rect 21760 49574 21836 49782
rect 20878 49510 20879 49542
rect 20813 49509 20879 49510
rect 21760 49510 21766 49574
rect 21830 49510 21836 49574
rect 21760 49504 21836 49510
rect 22168 49782 22174 49814
rect 22238 49814 22239 49846
rect 22440 49846 22516 49852
rect 22238 49782 22244 49814
rect 22168 49574 22244 49782
rect 22168 49510 22174 49574
rect 22238 49510 22244 49574
rect 22440 49782 22446 49846
rect 22510 49782 22516 49846
rect 114245 49846 114311 49847
rect 114245 49814 114246 49846
rect 22440 49574 22516 49782
rect 22440 49542 22446 49574
rect 22168 49504 22244 49510
rect 22445 49510 22446 49542
rect 22510 49542 22516 49574
rect 114240 49782 114246 49814
rect 114310 49814 114311 49846
rect 114653 49846 114719 49847
rect 114653 49814 114654 49846
rect 114310 49782 114316 49814
rect 114240 49574 114316 49782
rect 22510 49510 22511 49542
rect 22445 49509 22511 49510
rect 114240 49510 114246 49574
rect 114310 49510 114316 49574
rect 114240 49504 114316 49510
rect 114648 49782 114654 49814
rect 114718 49814 114719 49846
rect 115192 49846 115268 49852
rect 114718 49782 114724 49814
rect 114648 49574 114724 49782
rect 114648 49510 114654 49574
rect 114718 49510 114724 49574
rect 115192 49782 115198 49846
rect 115262 49782 115268 49846
rect 115192 49574 115268 49782
rect 115192 49542 115198 49574
rect 114648 49504 114724 49510
rect 115197 49510 115198 49542
rect 115262 49542 115268 49574
rect 115328 49846 115404 49852
rect 115328 49782 115334 49846
rect 115398 49782 115404 49846
rect 115328 49574 115404 49782
rect 115328 49542 115334 49574
rect 115262 49510 115263 49542
rect 115197 49509 115263 49510
rect 115333 49510 115334 49542
rect 115398 49542 115404 49574
rect 115872 49846 115948 49852
rect 115872 49782 115878 49846
rect 115942 49782 115948 49846
rect 115872 49574 115948 49782
rect 115872 49542 115878 49574
rect 115398 49510 115399 49542
rect 115333 49509 115399 49510
rect 115877 49510 115878 49542
rect 115942 49542 115948 49574
rect 115942 49510 115943 49542
rect 115877 49509 115943 49510
rect 20944 49438 21020 49444
rect 20944 49374 20950 49438
rect 21014 49374 21020 49438
rect 21221 49438 21287 49439
rect 21221 49406 21222 49438
rect 20944 49166 21020 49374
rect 20944 49134 20950 49166
rect 20949 49102 20950 49134
rect 21014 49134 21020 49166
rect 21216 49374 21222 49406
rect 21286 49406 21287 49438
rect 21624 49438 21700 49444
rect 21286 49374 21292 49406
rect 21216 49166 21292 49374
rect 21014 49102 21015 49134
rect 20949 49101 21015 49102
rect 21216 49102 21222 49166
rect 21286 49102 21292 49166
rect 21624 49374 21630 49438
rect 21694 49374 21700 49438
rect 22037 49438 22103 49439
rect 22037 49406 22038 49438
rect 21624 49166 21700 49374
rect 21624 49134 21630 49166
rect 21216 49096 21292 49102
rect 21629 49102 21630 49134
rect 21694 49134 21700 49166
rect 22032 49374 22038 49406
rect 22102 49406 22103 49438
rect 22445 49438 22511 49439
rect 22445 49406 22446 49438
rect 22102 49374 22108 49406
rect 22032 49166 22108 49374
rect 21694 49102 21695 49134
rect 21629 49101 21695 49102
rect 22032 49102 22038 49166
rect 22102 49102 22108 49166
rect 22032 49096 22108 49102
rect 22440 49374 22446 49406
rect 22510 49406 22511 49438
rect 114376 49438 114452 49444
rect 22510 49374 22516 49406
rect 22440 49166 22516 49374
rect 22440 49102 22446 49166
rect 22510 49102 22516 49166
rect 114376 49374 114382 49438
rect 114446 49374 114452 49438
rect 114376 49166 114452 49374
rect 114376 49134 114382 49166
rect 22440 49096 22516 49102
rect 114381 49102 114382 49134
rect 114446 49134 114452 49166
rect 114648 49438 114724 49444
rect 114648 49374 114654 49438
rect 114718 49374 114724 49438
rect 115877 49438 115943 49439
rect 115877 49406 115878 49438
rect 114648 49166 114724 49374
rect 114648 49134 114654 49166
rect 114446 49102 114447 49134
rect 114381 49101 114447 49102
rect 114653 49102 114654 49134
rect 114718 49134 114724 49166
rect 115872 49374 115878 49406
rect 115942 49406 115943 49438
rect 115942 49374 115948 49406
rect 115872 49166 115948 49374
rect 114718 49102 114719 49134
rect 114653 49101 114719 49102
rect 115872 49102 115878 49166
rect 115942 49102 115948 49166
rect 115872 49096 115948 49102
rect 952 48966 1230 49030
rect 1294 48966 1300 49030
rect 20813 49030 20879 49031
rect 20813 48998 20814 49030
rect 952 47534 1300 48966
rect 20808 48966 20814 48998
rect 20878 48998 20879 49030
rect 21352 49030 21428 49036
rect 20878 48966 20884 48998
rect 20808 48758 20884 48966
rect 20808 48694 20814 48758
rect 20878 48694 20884 48758
rect 21352 48966 21358 49030
rect 21422 48966 21428 49030
rect 21352 48758 21428 48966
rect 21352 48726 21358 48758
rect 20808 48688 20884 48694
rect 21357 48694 21358 48726
rect 21422 48726 21428 48758
rect 21488 49030 21564 49036
rect 21488 48966 21494 49030
rect 21558 48966 21564 49030
rect 21488 48758 21564 48966
rect 21488 48726 21494 48758
rect 21422 48694 21423 48726
rect 21357 48693 21423 48694
rect 21493 48694 21494 48726
rect 21558 48726 21564 48758
rect 22168 49030 22244 49036
rect 22168 48966 22174 49030
rect 22238 48966 22244 49030
rect 22168 48758 22244 48966
rect 22168 48726 22174 48758
rect 21558 48694 21559 48726
rect 21493 48693 21559 48694
rect 22173 48694 22174 48726
rect 22238 48726 22244 48758
rect 22576 49030 22652 49036
rect 22576 48966 22582 49030
rect 22646 48966 22652 49030
rect 114245 49030 114311 49031
rect 114245 48998 114246 49030
rect 22576 48758 22652 48966
rect 22576 48726 22582 48758
rect 22238 48694 22239 48726
rect 22173 48693 22239 48694
rect 22581 48694 22582 48726
rect 22646 48726 22652 48758
rect 114240 48966 114246 48998
rect 114310 48998 114311 49030
rect 114648 49030 114724 49036
rect 114310 48966 114316 48998
rect 114240 48758 114316 48966
rect 22646 48694 22647 48726
rect 22581 48693 22647 48694
rect 114240 48694 114246 48758
rect 114310 48694 114316 48758
rect 114648 48966 114654 49030
rect 114718 48966 114724 49030
rect 114648 48758 114724 48966
rect 114648 48726 114654 48758
rect 114240 48688 114316 48694
rect 114653 48694 114654 48726
rect 114718 48726 114724 48758
rect 115600 49030 115676 49036
rect 115600 48966 115606 49030
rect 115670 48966 115676 49030
rect 116013 49030 116079 49031
rect 116013 48998 116014 49030
rect 115600 48758 115676 48966
rect 115600 48726 115606 48758
rect 114718 48694 114719 48726
rect 114653 48693 114719 48694
rect 115605 48694 115606 48726
rect 115670 48726 115676 48758
rect 116008 48966 116014 48998
rect 116078 48998 116079 49030
rect 135320 49030 135668 50734
rect 116078 48966 116084 48998
rect 116008 48758 116084 48966
rect 115670 48694 115671 48726
rect 115605 48693 115671 48694
rect 116008 48694 116014 48758
rect 116078 48694 116084 48758
rect 116008 48688 116084 48694
rect 135320 48966 135326 49030
rect 135390 48966 135668 49030
rect 21765 48622 21831 48623
rect 21765 48590 21766 48622
rect 21760 48558 21766 48590
rect 21830 48590 21831 48622
rect 22173 48622 22239 48623
rect 22173 48590 22174 48622
rect 21830 48558 21836 48590
rect 20813 48350 20879 48351
rect 20813 48318 20814 48350
rect 20808 48286 20814 48318
rect 20878 48318 20879 48350
rect 21760 48350 21836 48558
rect 20878 48286 20884 48318
rect 20808 48078 20884 48286
rect 21760 48286 21766 48350
rect 21830 48286 21836 48350
rect 21760 48280 21836 48286
rect 22168 48558 22174 48590
rect 22238 48590 22239 48622
rect 22440 48622 22516 48628
rect 22238 48558 22244 48590
rect 22168 48350 22244 48558
rect 22168 48286 22174 48350
rect 22238 48286 22244 48350
rect 22440 48558 22446 48622
rect 22510 48558 22516 48622
rect 22440 48350 22516 48558
rect 22440 48318 22446 48350
rect 22168 48280 22244 48286
rect 22445 48286 22446 48318
rect 22510 48318 22516 48350
rect 114376 48622 114452 48628
rect 114376 48558 114382 48622
rect 114446 48558 114452 48622
rect 114653 48622 114719 48623
rect 114653 48590 114654 48622
rect 114376 48350 114452 48558
rect 114376 48318 114382 48350
rect 22510 48286 22511 48318
rect 22445 48285 22511 48286
rect 114381 48286 114382 48318
rect 114446 48318 114452 48350
rect 114648 48558 114654 48590
rect 114718 48590 114719 48622
rect 115061 48622 115127 48623
rect 115061 48590 115062 48622
rect 114718 48558 114724 48590
rect 114648 48350 114724 48558
rect 114446 48286 114447 48318
rect 114381 48285 114447 48286
rect 114648 48286 114654 48350
rect 114718 48286 114724 48350
rect 114648 48280 114724 48286
rect 115056 48558 115062 48590
rect 115126 48590 115127 48622
rect 115464 48622 115540 48628
rect 115126 48558 115132 48590
rect 115056 48350 115132 48558
rect 115464 48558 115470 48622
rect 115534 48558 115540 48622
rect 115056 48286 115062 48350
rect 115126 48286 115132 48350
rect 115333 48350 115399 48351
rect 115333 48318 115334 48350
rect 115056 48280 115132 48286
rect 115328 48286 115334 48318
rect 115398 48318 115399 48350
rect 115464 48350 115540 48558
rect 115464 48318 115470 48350
rect 115398 48286 115404 48318
rect 20808 48014 20814 48078
rect 20878 48014 20884 48078
rect 20808 48008 20884 48014
rect 22168 48214 22244 48220
rect 22168 48150 22174 48214
rect 22238 48150 22244 48214
rect 22168 47942 22244 48150
rect 22168 47910 22174 47942
rect 22173 47878 22174 47910
rect 22238 47910 22244 47942
rect 22440 48214 22516 48220
rect 22440 48150 22446 48214
rect 22510 48150 22516 48214
rect 22440 47942 22516 48150
rect 22440 47910 22446 47942
rect 22238 47878 22239 47910
rect 22173 47877 22239 47878
rect 22445 47878 22446 47910
rect 22510 47910 22516 47942
rect 114240 48214 114316 48220
rect 114240 48150 114246 48214
rect 114310 48150 114316 48214
rect 114789 48214 114855 48215
rect 114789 48182 114790 48214
rect 114240 47942 114316 48150
rect 114240 47910 114246 47942
rect 22510 47878 22511 47910
rect 22445 47877 22511 47878
rect 114245 47878 114246 47910
rect 114310 47910 114316 47942
rect 114784 48150 114790 48182
rect 114854 48182 114855 48214
rect 114854 48150 114860 48182
rect 114784 47942 114860 48150
rect 115328 48078 115404 48286
rect 115469 48286 115470 48318
rect 115534 48318 115540 48350
rect 115877 48350 115943 48351
rect 115877 48318 115878 48350
rect 115534 48286 115535 48318
rect 115469 48285 115535 48286
rect 115872 48286 115878 48318
rect 115942 48318 115943 48350
rect 115942 48286 115948 48318
rect 115328 48014 115334 48078
rect 115398 48014 115404 48078
rect 115328 48008 115404 48014
rect 115872 48078 115948 48286
rect 115872 48014 115878 48078
rect 115942 48014 115948 48078
rect 115872 48008 115948 48014
rect 114310 47878 114311 47910
rect 114245 47877 114311 47878
rect 114784 47878 114790 47942
rect 114854 47878 114860 47942
rect 114784 47872 114860 47878
rect 21493 47806 21559 47807
rect 21493 47774 21494 47806
rect 21488 47742 21494 47774
rect 21558 47774 21559 47806
rect 115056 47806 115132 47812
rect 21558 47742 21564 47774
rect 952 47470 1230 47534
rect 1294 47470 1300 47534
rect 952 45630 1300 47470
rect 20808 47534 20884 47540
rect 20808 47470 20814 47534
rect 20878 47470 20884 47534
rect 20808 47262 20884 47470
rect 21488 47534 21564 47742
rect 21488 47470 21494 47534
rect 21558 47470 21564 47534
rect 115056 47742 115062 47806
rect 115126 47742 115132 47806
rect 115056 47534 115132 47742
rect 115056 47502 115062 47534
rect 21488 47464 21564 47470
rect 115061 47470 115062 47502
rect 115126 47502 115132 47534
rect 115872 47534 115948 47540
rect 115126 47470 115127 47502
rect 115061 47469 115127 47470
rect 115872 47470 115878 47534
rect 115942 47470 115948 47534
rect 20808 47230 20814 47262
rect 20813 47198 20814 47230
rect 20878 47230 20884 47262
rect 27336 47262 27412 47268
rect 20878 47198 20879 47230
rect 20813 47197 20879 47198
rect 27336 47198 27342 47262
rect 27406 47198 27412 47262
rect 109349 47262 109415 47263
rect 109349 47230 109350 47262
rect 20949 47126 21015 47127
rect 20949 47094 20950 47126
rect 20944 47062 20950 47094
rect 21014 47094 21015 47126
rect 21352 47126 21428 47132
rect 21014 47062 21020 47094
rect 20944 46854 21020 47062
rect 20944 46790 20950 46854
rect 21014 46790 21020 46854
rect 21352 47062 21358 47126
rect 21422 47062 21428 47126
rect 21765 47126 21831 47127
rect 21765 47094 21766 47126
rect 21352 46854 21428 47062
rect 21352 46822 21358 46854
rect 20944 46784 21020 46790
rect 21357 46790 21358 46822
rect 21422 46822 21428 46854
rect 21760 47062 21766 47094
rect 21830 47094 21831 47126
rect 21830 47062 21836 47094
rect 21760 46854 21836 47062
rect 27336 46990 27412 47198
rect 27336 46958 27342 46990
rect 27341 46926 27342 46958
rect 27406 46958 27412 46990
rect 109344 47198 109350 47230
rect 109414 47230 109415 47262
rect 115872 47262 115948 47470
rect 115872 47230 115878 47262
rect 109414 47198 109420 47230
rect 109344 46990 109420 47198
rect 115877 47198 115878 47230
rect 115942 47230 115948 47262
rect 135320 47534 135668 48966
rect 135320 47470 135326 47534
rect 135390 47470 135668 47534
rect 115942 47198 115943 47230
rect 115877 47197 115943 47198
rect 115333 47126 115399 47127
rect 115333 47094 115334 47126
rect 27406 46926 27407 46958
rect 27341 46925 27407 46926
rect 109344 46926 109350 46990
rect 109414 46926 109420 46990
rect 109344 46920 109420 46926
rect 115328 47062 115334 47094
rect 115398 47094 115399 47126
rect 115877 47126 115943 47127
rect 115877 47094 115878 47126
rect 115398 47062 115404 47094
rect 21422 46790 21423 46822
rect 21357 46789 21423 46790
rect 21760 46790 21766 46854
rect 21830 46790 21836 46854
rect 21760 46784 21836 46790
rect 27336 46854 27412 46860
rect 27336 46790 27342 46854
rect 27406 46790 27412 46854
rect 20813 46718 20879 46719
rect 20813 46686 20814 46718
rect 20808 46654 20814 46686
rect 20878 46686 20879 46718
rect 22173 46718 22239 46719
rect 22173 46686 22174 46718
rect 20878 46654 20884 46686
rect 20808 46446 20884 46654
rect 20808 46382 20814 46446
rect 20878 46382 20884 46446
rect 20808 46376 20884 46382
rect 22168 46654 22174 46686
rect 22238 46686 22239 46718
rect 22576 46718 22652 46724
rect 22238 46654 22244 46686
rect 22168 46446 22244 46654
rect 22168 46382 22174 46446
rect 22238 46382 22244 46446
rect 22576 46654 22582 46718
rect 22646 46654 22652 46718
rect 22576 46446 22652 46654
rect 27336 46582 27412 46790
rect 27336 46550 27342 46582
rect 27341 46518 27342 46550
rect 27406 46550 27412 46582
rect 109480 46854 109556 46860
rect 109480 46790 109486 46854
rect 109550 46790 109556 46854
rect 109480 46582 109556 46790
rect 115328 46854 115404 47062
rect 115328 46790 115334 46854
rect 115398 46790 115404 46854
rect 115328 46784 115404 46790
rect 115872 47062 115878 47094
rect 115942 47094 115943 47126
rect 115942 47062 115948 47094
rect 115872 46854 115948 47062
rect 115872 46790 115878 46854
rect 115942 46790 115948 46854
rect 115872 46784 115948 46790
rect 109480 46550 109486 46582
rect 27406 46518 27407 46550
rect 27341 46517 27407 46518
rect 109485 46518 109486 46550
rect 109550 46550 109556 46582
rect 114240 46718 114316 46724
rect 114240 46654 114246 46718
rect 114310 46654 114316 46718
rect 109550 46518 109551 46550
rect 109485 46517 109551 46518
rect 22576 46414 22582 46446
rect 22168 46376 22244 46382
rect 22581 46382 22582 46414
rect 22646 46414 22652 46446
rect 114240 46446 114316 46654
rect 114240 46414 114246 46446
rect 22646 46382 22647 46414
rect 22581 46381 22647 46382
rect 114245 46382 114246 46414
rect 114310 46414 114316 46446
rect 114648 46718 114724 46724
rect 114648 46654 114654 46718
rect 114718 46654 114724 46718
rect 114648 46446 114724 46654
rect 114648 46414 114654 46446
rect 114310 46382 114311 46414
rect 114245 46381 114311 46382
rect 114653 46382 114654 46414
rect 114718 46414 114724 46446
rect 116008 46718 116084 46724
rect 116008 46654 116014 46718
rect 116078 46654 116084 46718
rect 116008 46446 116084 46654
rect 116008 46414 116014 46446
rect 114718 46382 114719 46414
rect 114653 46381 114719 46382
rect 116013 46382 116014 46414
rect 116078 46414 116084 46446
rect 116078 46382 116079 46414
rect 116013 46381 116079 46382
rect 20944 46310 21020 46316
rect 20944 46246 20950 46310
rect 21014 46246 21020 46310
rect 21221 46310 21287 46311
rect 21221 46278 21222 46310
rect 20944 46038 21020 46246
rect 20944 46006 20950 46038
rect 20949 45974 20950 46006
rect 21014 46006 21020 46038
rect 21216 46246 21222 46278
rect 21286 46278 21287 46310
rect 22032 46310 22108 46316
rect 21286 46246 21292 46278
rect 21216 46038 21292 46246
rect 21014 45974 21015 46006
rect 20949 45973 21015 45974
rect 21216 45974 21222 46038
rect 21286 45974 21292 46038
rect 22032 46246 22038 46310
rect 22102 46246 22108 46310
rect 22032 46038 22108 46246
rect 22032 46006 22038 46038
rect 21216 45968 21292 45974
rect 22037 45974 22038 46006
rect 22102 46006 22108 46038
rect 22576 46310 22652 46316
rect 22576 46246 22582 46310
rect 22646 46246 22652 46310
rect 114381 46310 114447 46311
rect 114381 46278 114382 46310
rect 22576 46038 22652 46246
rect 22576 46006 22582 46038
rect 22102 45974 22103 46006
rect 22037 45973 22103 45974
rect 22581 45974 22582 46006
rect 22646 46006 22652 46038
rect 114376 46246 114382 46278
rect 114446 46278 114447 46310
rect 114789 46310 114855 46311
rect 114789 46278 114790 46310
rect 114446 46246 114452 46278
rect 114376 46038 114452 46246
rect 22646 45974 22647 46006
rect 22581 45973 22647 45974
rect 114376 45974 114382 46038
rect 114446 45974 114452 46038
rect 114376 45968 114452 45974
rect 114784 46246 114790 46278
rect 114854 46278 114855 46310
rect 115197 46310 115263 46311
rect 115197 46278 115198 46310
rect 114854 46246 114860 46278
rect 114784 46038 114860 46246
rect 114784 45974 114790 46038
rect 114854 45974 114860 46038
rect 114784 45968 114860 45974
rect 115192 46246 115198 46278
rect 115262 46278 115263 46310
rect 115328 46310 115404 46316
rect 115262 46246 115268 46278
rect 115192 46038 115268 46246
rect 115192 45974 115198 46038
rect 115262 45974 115268 46038
rect 115328 46246 115334 46310
rect 115398 46246 115404 46310
rect 115469 46310 115535 46311
rect 115469 46278 115470 46310
rect 115328 46038 115404 46246
rect 115328 46006 115334 46038
rect 115192 45968 115268 45974
rect 115333 45974 115334 46006
rect 115398 46006 115404 46038
rect 115464 46246 115470 46278
rect 115534 46278 115535 46310
rect 115877 46310 115943 46311
rect 115877 46278 115878 46310
rect 115534 46246 115540 46278
rect 115464 46038 115540 46246
rect 115398 45974 115399 46006
rect 115333 45973 115399 45974
rect 115464 45974 115470 46038
rect 115534 45974 115540 46038
rect 115464 45968 115540 45974
rect 115872 46246 115878 46278
rect 115942 46278 115943 46310
rect 115942 46246 115948 46278
rect 115872 46038 115948 46246
rect 115872 45974 115878 46038
rect 115942 45974 115948 46038
rect 115872 45968 115948 45974
rect 20949 45902 21015 45903
rect 20949 45870 20950 45902
rect 952 45566 1230 45630
rect 1294 45566 1300 45630
rect 952 44134 1300 45566
rect 20944 45838 20950 45870
rect 21014 45870 21015 45902
rect 21352 45902 21428 45908
rect 21014 45838 21020 45870
rect 20944 45630 21020 45838
rect 20944 45566 20950 45630
rect 21014 45566 21020 45630
rect 21352 45838 21358 45902
rect 21422 45838 21428 45902
rect 22037 45902 22103 45903
rect 22037 45870 22038 45902
rect 21352 45630 21428 45838
rect 21352 45598 21358 45630
rect 20944 45560 21020 45566
rect 21357 45566 21358 45598
rect 21422 45598 21428 45630
rect 22032 45838 22038 45870
rect 22102 45870 22103 45902
rect 22440 45902 22516 45908
rect 22102 45838 22108 45870
rect 22032 45630 22108 45838
rect 21422 45566 21423 45598
rect 21357 45565 21423 45566
rect 22032 45566 22038 45630
rect 22102 45566 22108 45630
rect 22440 45838 22446 45902
rect 22510 45838 22516 45902
rect 114381 45902 114447 45903
rect 114381 45870 114382 45902
rect 22440 45630 22516 45838
rect 22440 45598 22446 45630
rect 22032 45560 22108 45566
rect 22445 45566 22446 45598
rect 22510 45598 22516 45630
rect 114376 45838 114382 45870
rect 114446 45870 114447 45902
rect 114648 45902 114724 45908
rect 114446 45838 114452 45870
rect 114376 45630 114452 45838
rect 22510 45566 22511 45598
rect 22445 45565 22511 45566
rect 114376 45566 114382 45630
rect 114446 45566 114452 45630
rect 114648 45838 114654 45902
rect 114718 45838 114724 45902
rect 114648 45630 114724 45838
rect 114648 45598 114654 45630
rect 114376 45560 114452 45566
rect 114653 45566 114654 45598
rect 114718 45598 114724 45630
rect 115464 45902 115540 45908
rect 115464 45838 115470 45902
rect 115534 45838 115540 45902
rect 115464 45630 115540 45838
rect 115464 45598 115470 45630
rect 114718 45566 114719 45598
rect 114653 45565 114719 45566
rect 115469 45566 115470 45598
rect 115534 45598 115540 45630
rect 116008 45902 116084 45908
rect 116008 45838 116014 45902
rect 116078 45838 116084 45902
rect 116008 45630 116084 45838
rect 116008 45598 116014 45630
rect 115534 45566 115535 45598
rect 115469 45565 115535 45566
rect 116013 45566 116014 45598
rect 116078 45598 116084 45630
rect 135320 45766 135668 47470
rect 135320 45702 135326 45766
rect 135390 45702 135668 45766
rect 116078 45566 116079 45598
rect 116013 45565 116079 45566
rect 20813 45494 20879 45495
rect 20813 45462 20814 45494
rect 20808 45430 20814 45462
rect 20878 45462 20879 45494
rect 21760 45494 21836 45500
rect 20878 45430 20884 45462
rect 20808 45222 20884 45430
rect 20808 45158 20814 45222
rect 20878 45158 20884 45222
rect 21760 45430 21766 45494
rect 21830 45430 21836 45494
rect 21760 45222 21836 45430
rect 21760 45190 21766 45222
rect 20808 45152 20884 45158
rect 21765 45158 21766 45190
rect 21830 45190 21836 45222
rect 22032 45494 22108 45500
rect 22032 45430 22038 45494
rect 22102 45430 22108 45494
rect 22445 45494 22511 45495
rect 22445 45462 22446 45494
rect 22032 45222 22108 45430
rect 22032 45190 22038 45222
rect 21830 45158 21831 45190
rect 21765 45157 21831 45158
rect 22037 45158 22038 45190
rect 22102 45190 22108 45222
rect 22440 45430 22446 45462
rect 22510 45462 22511 45494
rect 25840 45494 25916 45500
rect 22510 45430 22516 45462
rect 22440 45222 22516 45430
rect 22102 45158 22103 45190
rect 22037 45157 22103 45158
rect 22440 45158 22446 45222
rect 22510 45158 22516 45222
rect 25840 45430 25846 45494
rect 25910 45430 25916 45494
rect 25840 45222 25916 45430
rect 25840 45190 25846 45222
rect 22440 45152 22516 45158
rect 25845 45158 25846 45190
rect 25910 45190 25916 45222
rect 113696 45494 113772 45500
rect 113696 45430 113702 45494
rect 113766 45430 113772 45494
rect 113696 45222 113772 45430
rect 113696 45190 113702 45222
rect 25910 45158 25911 45190
rect 25845 45157 25911 45158
rect 113701 45158 113702 45190
rect 113766 45190 113772 45222
rect 114376 45494 114452 45500
rect 114376 45430 114382 45494
rect 114446 45430 114452 45494
rect 114376 45222 114452 45430
rect 114376 45190 114382 45222
rect 113766 45158 113767 45190
rect 113701 45157 113767 45158
rect 114381 45158 114382 45190
rect 114446 45190 114452 45222
rect 114784 45494 114860 45500
rect 114784 45430 114790 45494
rect 114854 45430 114860 45494
rect 114784 45222 114860 45430
rect 114784 45190 114790 45222
rect 114446 45158 114447 45190
rect 114381 45157 114447 45158
rect 114789 45158 114790 45190
rect 114854 45190 114860 45222
rect 115192 45494 115268 45500
rect 115192 45430 115198 45494
rect 115262 45430 115268 45494
rect 115192 45222 115268 45430
rect 115192 45190 115198 45222
rect 114854 45158 114855 45190
rect 114789 45157 114855 45158
rect 115197 45158 115198 45190
rect 115262 45190 115268 45222
rect 115328 45494 115404 45500
rect 115328 45430 115334 45494
rect 115398 45430 115404 45494
rect 115328 45222 115404 45430
rect 115328 45190 115334 45222
rect 115262 45158 115263 45190
rect 115197 45157 115263 45158
rect 115333 45158 115334 45190
rect 115398 45190 115404 45222
rect 115872 45494 115948 45500
rect 115872 45430 115878 45494
rect 115942 45430 115948 45494
rect 115872 45222 115948 45430
rect 115872 45190 115878 45222
rect 115398 45158 115399 45190
rect 115333 45157 115399 45158
rect 115877 45158 115878 45190
rect 115942 45190 115948 45222
rect 115942 45158 115943 45190
rect 115877 45157 115943 45158
rect 20944 45086 21020 45092
rect 20944 45022 20950 45086
rect 21014 45022 21020 45086
rect 20944 44814 21020 45022
rect 20944 44782 20950 44814
rect 20949 44750 20950 44782
rect 21014 44782 21020 44814
rect 21216 45086 21292 45092
rect 21216 45022 21222 45086
rect 21286 45022 21292 45086
rect 21216 44814 21292 45022
rect 21216 44782 21222 44814
rect 21014 44750 21015 44782
rect 20949 44749 21015 44750
rect 21221 44750 21222 44782
rect 21286 44782 21292 44814
rect 21488 45086 21564 45092
rect 21488 45022 21494 45086
rect 21558 45022 21564 45086
rect 21488 44814 21564 45022
rect 21488 44782 21494 44814
rect 21286 44750 21287 44782
rect 21221 44749 21287 44750
rect 21493 44750 21494 44782
rect 21558 44782 21564 44814
rect 22032 45086 22108 45092
rect 22032 45022 22038 45086
rect 22102 45022 22108 45086
rect 22032 44814 22108 45022
rect 22032 44782 22038 44814
rect 21558 44750 21559 44782
rect 21493 44749 21559 44750
rect 22037 44750 22038 44782
rect 22102 44782 22108 44814
rect 22576 45086 22652 45092
rect 22576 45022 22582 45086
rect 22646 45022 22652 45086
rect 22576 44814 22652 45022
rect 22576 44782 22582 44814
rect 22102 44750 22103 44782
rect 22037 44749 22103 44750
rect 22581 44750 22582 44782
rect 22646 44782 22652 44814
rect 23256 45086 23332 45092
rect 23256 45022 23262 45086
rect 23326 45022 23332 45086
rect 23256 44814 23332 45022
rect 23256 44782 23262 44814
rect 22646 44750 22647 44782
rect 22581 44749 22647 44750
rect 23261 44750 23262 44782
rect 23326 44782 23332 44814
rect 112336 45086 112412 45092
rect 112336 45022 112342 45086
rect 112406 45022 112412 45086
rect 114381 45086 114447 45087
rect 114381 45054 114382 45086
rect 23326 44750 23327 44782
rect 23261 44749 23327 44750
rect 21357 44678 21423 44679
rect 21357 44646 21358 44678
rect 21352 44614 21358 44646
rect 21422 44646 21423 44678
rect 22168 44678 22244 44684
rect 21422 44614 21428 44646
rect 21352 44406 21428 44614
rect 21352 44342 21358 44406
rect 21422 44342 21428 44406
rect 22168 44614 22174 44678
rect 22238 44614 22244 44678
rect 22445 44678 22511 44679
rect 22445 44646 22446 44678
rect 22168 44406 22244 44614
rect 22168 44374 22174 44406
rect 21352 44336 21428 44342
rect 22173 44342 22174 44374
rect 22238 44374 22244 44406
rect 22440 44614 22446 44646
rect 22510 44646 22511 44678
rect 112336 44678 112412 45022
rect 114376 45022 114382 45054
rect 114446 45054 114447 45086
rect 114648 45086 114724 45092
rect 114446 45022 114452 45054
rect 114376 44814 114452 45022
rect 114376 44750 114382 44814
rect 114446 44750 114452 44814
rect 114648 45022 114654 45086
rect 114718 45022 114724 45086
rect 114648 44814 114724 45022
rect 114648 44782 114654 44814
rect 114376 44744 114452 44750
rect 114653 44750 114654 44782
rect 114718 44782 114724 44814
rect 115872 45086 115948 45092
rect 115872 45022 115878 45086
rect 115942 45022 115948 45086
rect 115872 44814 115948 45022
rect 115872 44782 115878 44814
rect 114718 44750 114719 44782
rect 114653 44749 114719 44750
rect 115877 44750 115878 44782
rect 115942 44782 115948 44814
rect 115942 44750 115943 44782
rect 115877 44749 115943 44750
rect 112336 44646 112342 44678
rect 22510 44614 22516 44646
rect 22440 44406 22516 44614
rect 112341 44614 112342 44646
rect 112406 44646 112412 44678
rect 114240 44678 114316 44684
rect 112406 44614 112407 44646
rect 112341 44613 112407 44614
rect 114240 44614 114246 44678
rect 114310 44614 114316 44678
rect 114653 44678 114719 44679
rect 114653 44646 114654 44678
rect 22238 44342 22239 44374
rect 22173 44341 22239 44342
rect 22440 44342 22446 44406
rect 22510 44342 22516 44406
rect 114240 44406 114316 44614
rect 114240 44374 114246 44406
rect 22440 44336 22516 44342
rect 114245 44342 114246 44374
rect 114310 44374 114316 44406
rect 114648 44614 114654 44646
rect 114718 44646 114719 44678
rect 115469 44678 115535 44679
rect 115469 44646 115470 44678
rect 114718 44614 114724 44646
rect 114648 44406 114724 44614
rect 114310 44342 114311 44374
rect 114245 44341 114311 44342
rect 114648 44342 114654 44406
rect 114718 44342 114724 44406
rect 114648 44336 114724 44342
rect 115464 44614 115470 44646
rect 115534 44646 115535 44678
rect 115534 44614 115540 44646
rect 115464 44406 115540 44614
rect 115464 44342 115470 44406
rect 115534 44342 115540 44406
rect 115464 44336 115540 44342
rect 22173 44270 22239 44271
rect 22173 44238 22174 44270
rect 952 44070 1230 44134
rect 1294 44070 1300 44134
rect 952 42502 1300 44070
rect 22168 44206 22174 44238
rect 22238 44238 22239 44270
rect 22581 44270 22647 44271
rect 22581 44238 22582 44270
rect 22238 44206 22244 44238
rect 22168 43998 22244 44206
rect 22168 43934 22174 43998
rect 22238 43934 22244 43998
rect 22168 43928 22244 43934
rect 22576 44206 22582 44238
rect 22646 44238 22647 44270
rect 114376 44270 114452 44276
rect 22646 44206 22652 44238
rect 22576 43998 22652 44206
rect 22576 43934 22582 43998
rect 22646 43934 22652 43998
rect 114376 44206 114382 44270
rect 114446 44206 114452 44270
rect 114376 43998 114452 44206
rect 114376 43966 114382 43998
rect 22576 43928 22652 43934
rect 114381 43934 114382 43966
rect 114446 43966 114452 43998
rect 114784 44270 114860 44276
rect 114784 44206 114790 44270
rect 114854 44206 114860 44270
rect 114784 43998 114860 44206
rect 114784 43966 114790 43998
rect 114446 43934 114447 43966
rect 114381 43933 114447 43934
rect 114789 43934 114790 43966
rect 114854 43966 114860 43998
rect 135320 43998 135668 45702
rect 114854 43934 114855 43966
rect 114789 43933 114855 43934
rect 135320 43934 135326 43998
rect 135390 43934 135668 43998
rect 21760 43862 21836 43868
rect 21760 43798 21766 43862
rect 21830 43798 21836 43862
rect 22037 43862 22103 43863
rect 22037 43830 22038 43862
rect 20813 43590 20879 43591
rect 20813 43558 20814 43590
rect 20808 43526 20814 43558
rect 20878 43558 20879 43590
rect 21760 43590 21836 43798
rect 21760 43558 21766 43590
rect 20878 43526 20884 43558
rect 20808 43318 20884 43526
rect 21765 43526 21766 43558
rect 21830 43558 21836 43590
rect 22032 43798 22038 43830
rect 22102 43830 22103 43862
rect 22445 43862 22511 43863
rect 22445 43830 22446 43862
rect 22102 43798 22108 43830
rect 22032 43590 22108 43798
rect 21830 43526 21831 43558
rect 21765 43525 21831 43526
rect 22032 43526 22038 43590
rect 22102 43526 22108 43590
rect 22032 43520 22108 43526
rect 22440 43798 22446 43830
rect 22510 43830 22511 43862
rect 114381 43862 114447 43863
rect 114381 43830 114382 43862
rect 22510 43798 22516 43830
rect 22440 43590 22516 43798
rect 114376 43798 114382 43830
rect 114446 43830 114447 43862
rect 114789 43862 114855 43863
rect 114789 43830 114790 43862
rect 114446 43798 114452 43830
rect 27477 43726 27543 43727
rect 27477 43694 27478 43726
rect 22440 43526 22446 43590
rect 22510 43526 22516 43590
rect 22440 43520 22516 43526
rect 27472 43662 27478 43694
rect 27542 43694 27543 43726
rect 109349 43726 109415 43727
rect 109349 43694 109350 43726
rect 27542 43662 27548 43694
rect 20808 43254 20814 43318
rect 20878 43254 20884 43318
rect 20808 43248 20884 43254
rect 21488 43454 21700 43460
rect 21488 43390 21630 43454
rect 21694 43390 21700 43454
rect 21488 43384 21700 43390
rect 27472 43454 27548 43662
rect 27472 43390 27478 43454
rect 27542 43390 27548 43454
rect 27472 43384 27548 43390
rect 109344 43662 109350 43694
rect 109414 43694 109415 43726
rect 109414 43662 109420 43694
rect 109344 43454 109420 43662
rect 114376 43590 114452 43798
rect 114376 43526 114382 43590
rect 114446 43526 114452 43590
rect 114376 43520 114452 43526
rect 114784 43798 114790 43830
rect 114854 43830 114855 43862
rect 115197 43862 115263 43863
rect 115197 43830 115198 43862
rect 114854 43798 114860 43830
rect 114784 43590 114860 43798
rect 114784 43526 114790 43590
rect 114854 43526 114860 43590
rect 114784 43520 114860 43526
rect 115192 43798 115198 43830
rect 115262 43830 115263 43862
rect 115262 43798 115268 43830
rect 115192 43590 115268 43798
rect 115192 43526 115198 43590
rect 115262 43526 115268 43590
rect 115192 43520 115268 43526
rect 116008 43590 116084 43596
rect 116008 43526 116014 43590
rect 116078 43526 116084 43590
rect 109344 43390 109350 43454
rect 109414 43390 109420 43454
rect 109344 43384 109420 43390
rect 20808 43182 20884 43188
rect 20808 43118 20814 43182
rect 20878 43118 20884 43182
rect 20808 42910 20884 43118
rect 20808 42878 20814 42910
rect 20813 42846 20814 42878
rect 20878 42878 20884 42910
rect 21216 43182 21292 43188
rect 21216 43118 21222 43182
rect 21286 43118 21292 43182
rect 21488 43182 21564 43384
rect 27613 43318 27679 43319
rect 27613 43286 27614 43318
rect 21488 43150 21494 43182
rect 21216 42910 21292 43118
rect 21493 43118 21494 43150
rect 21558 43150 21564 43182
rect 27608 43254 27614 43286
rect 27678 43286 27679 43318
rect 109344 43318 109420 43324
rect 27678 43254 27684 43286
rect 21558 43118 21559 43150
rect 21493 43117 21559 43118
rect 27608 43046 27684 43254
rect 27608 42982 27614 43046
rect 27678 42982 27684 43046
rect 109344 43254 109350 43318
rect 109414 43254 109420 43318
rect 116008 43318 116084 43526
rect 116008 43286 116014 43318
rect 109344 43046 109420 43254
rect 116013 43254 116014 43286
rect 116078 43286 116084 43318
rect 116078 43254 116079 43286
rect 116013 43253 116079 43254
rect 115061 43182 115127 43183
rect 115061 43150 115062 43182
rect 109344 43014 109350 43046
rect 27608 42976 27684 42982
rect 109349 42982 109350 43014
rect 109414 43014 109420 43046
rect 115056 43118 115062 43150
rect 115126 43150 115127 43182
rect 116013 43182 116079 43183
rect 116013 43150 116014 43182
rect 115126 43118 115132 43150
rect 109414 42982 109415 43014
rect 109349 42981 109415 42982
rect 21216 42878 21222 42910
rect 20878 42846 20879 42878
rect 20813 42845 20879 42846
rect 21221 42846 21222 42878
rect 21286 42878 21292 42910
rect 109349 42910 109415 42911
rect 109349 42878 109350 42910
rect 21286 42846 21287 42878
rect 21221 42845 21287 42846
rect 109344 42846 109350 42878
rect 109414 42878 109415 42910
rect 115056 42910 115132 43118
rect 109414 42846 109420 42878
rect 20813 42774 20879 42775
rect 20813 42742 20814 42774
rect 952 42438 1230 42502
rect 1294 42438 1300 42502
rect 952 40870 1300 42438
rect 20808 42710 20814 42742
rect 20878 42742 20879 42774
rect 22168 42774 22244 42780
rect 20878 42710 20884 42742
rect 20808 42502 20884 42710
rect 20808 42438 20814 42502
rect 20878 42438 20884 42502
rect 22168 42710 22174 42774
rect 22238 42710 22244 42774
rect 22168 42502 22244 42710
rect 22168 42470 22174 42502
rect 20808 42432 20884 42438
rect 22173 42438 22174 42470
rect 22238 42470 22244 42502
rect 22440 42774 22516 42780
rect 22440 42710 22446 42774
rect 22510 42710 22516 42774
rect 22440 42502 22516 42710
rect 109344 42638 109420 42846
rect 115056 42846 115062 42910
rect 115126 42846 115132 42910
rect 115056 42840 115132 42846
rect 116008 43118 116014 43150
rect 116078 43150 116079 43182
rect 116078 43118 116084 43150
rect 116008 42910 116084 43118
rect 116008 42846 116014 42910
rect 116078 42846 116084 42910
rect 116008 42840 116084 42846
rect 109344 42574 109350 42638
rect 109414 42574 109420 42638
rect 109344 42568 109420 42574
rect 114240 42774 114316 42780
rect 114240 42710 114246 42774
rect 114310 42710 114316 42774
rect 114789 42774 114855 42775
rect 114789 42742 114790 42774
rect 22440 42470 22446 42502
rect 22238 42438 22239 42470
rect 22173 42437 22239 42438
rect 22445 42438 22446 42470
rect 22510 42470 22516 42502
rect 114240 42502 114316 42710
rect 114240 42470 114246 42502
rect 22510 42438 22511 42470
rect 22445 42437 22511 42438
rect 114245 42438 114246 42470
rect 114310 42470 114316 42502
rect 114784 42710 114790 42742
rect 114854 42742 114855 42774
rect 115877 42774 115943 42775
rect 115877 42742 115878 42774
rect 114854 42710 114860 42742
rect 114784 42502 114860 42710
rect 114310 42438 114311 42470
rect 114245 42437 114311 42438
rect 114784 42438 114790 42502
rect 114854 42438 114860 42502
rect 114784 42432 114860 42438
rect 115872 42710 115878 42742
rect 115942 42742 115943 42774
rect 115942 42710 115948 42742
rect 115872 42502 115948 42710
rect 115872 42438 115878 42502
rect 115942 42438 115948 42502
rect 115872 42432 115948 42438
rect 20944 42366 21020 42372
rect 20944 42302 20950 42366
rect 21014 42302 21020 42366
rect 21765 42366 21831 42367
rect 21765 42334 21766 42366
rect 20944 42094 21020 42302
rect 20944 42062 20950 42094
rect 20949 42030 20950 42062
rect 21014 42062 21020 42094
rect 21760 42302 21766 42334
rect 21830 42334 21831 42366
rect 22173 42366 22239 42367
rect 22173 42334 22174 42366
rect 21830 42302 21836 42334
rect 21760 42094 21836 42302
rect 21014 42030 21015 42062
rect 20949 42029 21015 42030
rect 21760 42030 21766 42094
rect 21830 42030 21836 42094
rect 21760 42024 21836 42030
rect 22168 42302 22174 42334
rect 22238 42334 22239 42366
rect 22576 42366 22652 42372
rect 22238 42302 22244 42334
rect 22168 42094 22244 42302
rect 22168 42030 22174 42094
rect 22238 42030 22244 42094
rect 22576 42302 22582 42366
rect 22646 42302 22652 42366
rect 22576 42094 22652 42302
rect 22576 42062 22582 42094
rect 22168 42024 22244 42030
rect 22581 42030 22582 42062
rect 22646 42062 22652 42094
rect 114240 42366 114316 42372
rect 114240 42302 114246 42366
rect 114310 42302 114316 42366
rect 114240 42094 114316 42302
rect 114240 42062 114246 42094
rect 22646 42030 22647 42062
rect 22581 42029 22647 42030
rect 114245 42030 114246 42062
rect 114310 42062 114316 42094
rect 114648 42366 114724 42372
rect 114648 42302 114654 42366
rect 114718 42302 114724 42366
rect 114648 42094 114724 42302
rect 114648 42062 114654 42094
rect 114310 42030 114311 42062
rect 114245 42029 114311 42030
rect 114653 42030 114654 42062
rect 114718 42062 114724 42094
rect 115056 42366 115132 42372
rect 115056 42302 115062 42366
rect 115126 42302 115132 42366
rect 116013 42366 116079 42367
rect 116013 42334 116014 42366
rect 115056 42094 115132 42302
rect 115056 42062 115062 42094
rect 114718 42030 114719 42062
rect 114653 42029 114719 42030
rect 115061 42030 115062 42062
rect 115126 42062 115132 42094
rect 116008 42302 116014 42334
rect 116078 42334 116079 42366
rect 135320 42366 135668 43934
rect 116078 42302 116084 42334
rect 116008 42094 116084 42302
rect 115126 42030 115127 42062
rect 115061 42029 115127 42030
rect 116008 42030 116014 42094
rect 116078 42030 116084 42094
rect 116008 42024 116084 42030
rect 135320 42302 135326 42366
rect 135390 42302 135668 42366
rect 20813 41958 20879 41959
rect 20813 41926 20814 41958
rect 20808 41894 20814 41926
rect 20878 41926 20879 41958
rect 21221 41958 21287 41959
rect 21221 41926 21222 41958
rect 20878 41894 20884 41926
rect 20808 41686 20884 41894
rect 20808 41622 20814 41686
rect 20878 41622 20884 41686
rect 20808 41616 20884 41622
rect 21216 41894 21222 41926
rect 21286 41926 21287 41958
rect 21624 41958 21700 41964
rect 21286 41894 21292 41926
rect 21216 41686 21292 41894
rect 21216 41622 21222 41686
rect 21286 41622 21292 41686
rect 21624 41894 21630 41958
rect 21694 41894 21700 41958
rect 21624 41686 21700 41894
rect 21624 41654 21630 41686
rect 21216 41616 21292 41622
rect 21629 41622 21630 41654
rect 21694 41654 21700 41686
rect 22032 41958 22108 41964
rect 22032 41894 22038 41958
rect 22102 41894 22108 41958
rect 22445 41958 22511 41959
rect 22445 41926 22446 41958
rect 22032 41686 22108 41894
rect 22032 41654 22038 41686
rect 21694 41622 21695 41654
rect 21629 41621 21695 41622
rect 22037 41622 22038 41654
rect 22102 41654 22108 41686
rect 22440 41894 22446 41926
rect 22510 41926 22511 41958
rect 114381 41958 114447 41959
rect 114381 41926 114382 41958
rect 22510 41894 22516 41926
rect 22440 41686 22516 41894
rect 22102 41622 22103 41654
rect 22037 41621 22103 41622
rect 22440 41622 22446 41686
rect 22510 41622 22516 41686
rect 22440 41616 22516 41622
rect 114376 41894 114382 41926
rect 114446 41926 114447 41958
rect 114784 41958 114860 41964
rect 114446 41894 114452 41926
rect 114376 41686 114452 41894
rect 114376 41622 114382 41686
rect 114446 41622 114452 41686
rect 114784 41894 114790 41958
rect 114854 41894 114860 41958
rect 114784 41686 114860 41894
rect 114784 41654 114790 41686
rect 114376 41616 114452 41622
rect 114789 41622 114790 41654
rect 114854 41654 114860 41686
rect 115192 41958 115268 41964
rect 115192 41894 115198 41958
rect 115262 41894 115268 41958
rect 115192 41686 115268 41894
rect 115192 41654 115198 41686
rect 114854 41622 114855 41654
rect 114789 41621 114855 41622
rect 115197 41622 115198 41654
rect 115262 41654 115268 41686
rect 115328 41958 115404 41964
rect 115328 41894 115334 41958
rect 115398 41894 115404 41958
rect 115328 41686 115404 41894
rect 115328 41654 115334 41686
rect 115262 41622 115263 41654
rect 115197 41621 115263 41622
rect 115333 41622 115334 41654
rect 115398 41654 115404 41686
rect 115872 41958 115948 41964
rect 115872 41894 115878 41958
rect 115942 41894 115948 41958
rect 115872 41686 115948 41894
rect 115872 41654 115878 41686
rect 115398 41622 115399 41654
rect 115333 41621 115399 41622
rect 115877 41622 115878 41654
rect 115942 41654 115948 41686
rect 115942 41622 115943 41654
rect 115877 41621 115943 41622
rect 20808 41550 20884 41556
rect 20808 41486 20814 41550
rect 20878 41486 20884 41550
rect 20808 41278 20884 41486
rect 20808 41246 20814 41278
rect 20813 41214 20814 41246
rect 20878 41246 20884 41278
rect 21352 41550 21428 41556
rect 21352 41486 21358 41550
rect 21422 41486 21428 41550
rect 22037 41550 22103 41551
rect 22037 41518 22038 41550
rect 21352 41278 21428 41486
rect 21352 41246 21358 41278
rect 20878 41214 20879 41246
rect 20813 41213 20879 41214
rect 21357 41214 21358 41246
rect 21422 41246 21428 41278
rect 22032 41486 22038 41518
rect 22102 41518 22103 41550
rect 22581 41550 22647 41551
rect 22581 41518 22582 41550
rect 22102 41486 22108 41518
rect 22032 41278 22108 41486
rect 21422 41214 21423 41246
rect 21357 41213 21423 41214
rect 22032 41214 22038 41278
rect 22102 41214 22108 41278
rect 22032 41208 22108 41214
rect 22576 41486 22582 41518
rect 22646 41518 22647 41550
rect 114381 41550 114447 41551
rect 114381 41518 114382 41550
rect 22646 41486 22652 41518
rect 22576 41278 22652 41486
rect 22576 41214 22582 41278
rect 22646 41214 22652 41278
rect 22576 41208 22652 41214
rect 114376 41486 114382 41518
rect 114446 41518 114447 41550
rect 114789 41550 114855 41551
rect 114789 41518 114790 41550
rect 114446 41486 114452 41518
rect 114376 41278 114452 41486
rect 114376 41214 114382 41278
rect 114446 41214 114452 41278
rect 114376 41208 114452 41214
rect 114784 41486 114790 41518
rect 114854 41518 114855 41550
rect 115605 41550 115671 41551
rect 115605 41518 115606 41550
rect 114854 41486 114860 41518
rect 114784 41278 114860 41486
rect 114784 41214 114790 41278
rect 114854 41214 114860 41278
rect 114784 41208 114860 41214
rect 115600 41486 115606 41518
rect 115670 41518 115671 41550
rect 116008 41550 116084 41556
rect 115670 41486 115676 41518
rect 115600 41278 115676 41486
rect 115600 41214 115606 41278
rect 115670 41214 115676 41278
rect 116008 41486 116014 41550
rect 116078 41486 116084 41550
rect 116008 41278 116084 41486
rect 116008 41246 116014 41278
rect 115600 41208 115676 41214
rect 116013 41214 116014 41246
rect 116078 41246 116084 41278
rect 116078 41214 116079 41246
rect 116013 41213 116079 41214
rect 20813 41142 20879 41143
rect 20813 41110 20814 41142
rect 952 40806 1230 40870
rect 1294 40806 1300 40870
rect 952 39102 1300 40806
rect 20808 41078 20814 41110
rect 20878 41110 20879 41142
rect 21765 41142 21831 41143
rect 21765 41110 21766 41142
rect 20878 41078 20884 41110
rect 20808 40870 20884 41078
rect 20808 40806 20814 40870
rect 20878 40806 20884 40870
rect 20808 40800 20884 40806
rect 21760 41078 21766 41110
rect 21830 41110 21831 41142
rect 22032 41142 22108 41148
rect 21830 41078 21836 41110
rect 21760 40870 21836 41078
rect 21760 40806 21766 40870
rect 21830 40806 21836 40870
rect 22032 41078 22038 41142
rect 22102 41078 22108 41142
rect 22445 41142 22511 41143
rect 22445 41110 22446 41142
rect 22032 40870 22108 41078
rect 22032 40838 22038 40870
rect 21760 40800 21836 40806
rect 22037 40806 22038 40838
rect 22102 40838 22108 40870
rect 22440 41078 22446 41110
rect 22510 41110 22511 41142
rect 114376 41142 114452 41148
rect 22510 41078 22516 41110
rect 22440 40870 22516 41078
rect 22102 40806 22103 40838
rect 22037 40805 22103 40806
rect 22440 40806 22446 40870
rect 22510 40806 22516 40870
rect 114376 41078 114382 41142
rect 114446 41078 114452 41142
rect 114653 41142 114719 41143
rect 114653 41110 114654 41142
rect 114376 40870 114452 41078
rect 114376 40838 114382 40870
rect 22440 40800 22516 40806
rect 114381 40806 114382 40838
rect 114446 40838 114452 40870
rect 114648 41078 114654 41110
rect 114718 41110 114719 41142
rect 115192 41142 115268 41148
rect 114718 41078 114724 41110
rect 114648 40870 114724 41078
rect 114446 40806 114447 40838
rect 114381 40805 114447 40806
rect 114648 40806 114654 40870
rect 114718 40806 114724 40870
rect 115192 41078 115198 41142
rect 115262 41078 115268 41142
rect 115192 40870 115268 41078
rect 115192 40838 115198 40870
rect 114648 40800 114724 40806
rect 115197 40806 115198 40838
rect 115262 40838 115268 40870
rect 115328 41142 115404 41148
rect 115328 41078 115334 41142
rect 115398 41078 115404 41142
rect 115328 40870 115404 41078
rect 115328 40838 115334 40870
rect 115262 40806 115263 40838
rect 115197 40805 115263 40806
rect 115333 40806 115334 40838
rect 115398 40838 115404 40870
rect 115464 41142 115540 41148
rect 115464 41078 115470 41142
rect 115534 41078 115540 41142
rect 116013 41142 116079 41143
rect 116013 41110 116014 41142
rect 115464 40870 115540 41078
rect 115464 40838 115470 40870
rect 115398 40806 115399 40838
rect 115333 40805 115399 40806
rect 115469 40806 115470 40838
rect 115534 40838 115540 40870
rect 116008 41078 116014 41110
rect 116078 41110 116079 41142
rect 116078 41078 116084 41110
rect 116008 40870 116084 41078
rect 115534 40806 115535 40838
rect 115469 40805 115535 40806
rect 116008 40806 116014 40870
rect 116078 40806 116084 40870
rect 116008 40800 116084 40806
rect 135320 40870 135668 42302
rect 135320 40806 135326 40870
rect 135390 40806 135668 40870
rect 21221 40734 21287 40735
rect 21221 40702 21222 40734
rect 21216 40670 21222 40702
rect 21286 40702 21287 40734
rect 21624 40734 21700 40740
rect 21286 40670 21292 40702
rect 21216 40462 21292 40670
rect 21216 40398 21222 40462
rect 21286 40398 21292 40462
rect 21624 40670 21630 40734
rect 21694 40670 21700 40734
rect 22037 40734 22103 40735
rect 22037 40702 22038 40734
rect 21624 40462 21700 40670
rect 21624 40430 21630 40462
rect 21216 40392 21292 40398
rect 21629 40398 21630 40430
rect 21694 40430 21700 40462
rect 22032 40670 22038 40702
rect 22102 40702 22103 40734
rect 22576 40734 22652 40740
rect 22102 40670 22108 40702
rect 22032 40462 22108 40670
rect 21694 40398 21695 40430
rect 21629 40397 21695 40398
rect 22032 40398 22038 40462
rect 22102 40398 22108 40462
rect 22576 40670 22582 40734
rect 22646 40670 22652 40734
rect 114381 40734 114447 40735
rect 114381 40702 114382 40734
rect 22576 40462 22652 40670
rect 114376 40670 114382 40702
rect 114446 40702 114447 40734
rect 114648 40734 114724 40740
rect 114446 40670 114452 40702
rect 27477 40598 27543 40599
rect 27477 40566 27478 40598
rect 22576 40430 22582 40462
rect 22032 40392 22108 40398
rect 22581 40398 22582 40430
rect 22646 40430 22652 40462
rect 27472 40534 27478 40566
rect 27542 40566 27543 40598
rect 109480 40598 109556 40604
rect 27542 40534 27548 40566
rect 22646 40398 22647 40430
rect 22581 40397 22647 40398
rect 22173 40326 22239 40327
rect 22173 40294 22174 40326
rect 22168 40262 22174 40294
rect 22238 40294 22239 40326
rect 22445 40326 22511 40327
rect 22445 40294 22446 40326
rect 22238 40262 22244 40294
rect 22168 40054 22244 40262
rect 22168 39990 22174 40054
rect 22238 39990 22244 40054
rect 22168 39984 22244 39990
rect 22440 40262 22446 40294
rect 22510 40294 22511 40326
rect 27472 40326 27548 40534
rect 109480 40534 109486 40598
rect 109550 40534 109556 40598
rect 22510 40262 22516 40294
rect 22440 40054 22516 40262
rect 27472 40262 27478 40326
rect 27542 40262 27548 40326
rect 109349 40326 109415 40327
rect 109349 40294 109350 40326
rect 27472 40256 27548 40262
rect 109344 40262 109350 40294
rect 109414 40294 109415 40326
rect 109480 40326 109556 40534
rect 114376 40462 114452 40670
rect 114376 40398 114382 40462
rect 114446 40398 114452 40462
rect 114648 40670 114654 40734
rect 114718 40670 114724 40734
rect 114648 40462 114724 40670
rect 114648 40430 114654 40462
rect 114376 40392 114452 40398
rect 114653 40398 114654 40430
rect 114718 40430 114724 40462
rect 115328 40734 115404 40740
rect 115328 40670 115334 40734
rect 115398 40670 115404 40734
rect 115328 40462 115404 40670
rect 115328 40430 115334 40462
rect 114718 40398 114719 40430
rect 114653 40397 114719 40398
rect 115333 40398 115334 40430
rect 115398 40430 115404 40462
rect 115398 40398 115399 40430
rect 115333 40397 115399 40398
rect 109480 40294 109486 40326
rect 109414 40262 109420 40294
rect 22440 39990 22446 40054
rect 22510 39990 22516 40054
rect 22440 39984 22516 39990
rect 21765 39918 21831 39919
rect 21765 39886 21766 39918
rect 21760 39854 21766 39886
rect 21830 39886 21831 39918
rect 22032 39918 22108 39924
rect 21830 39854 21836 39886
rect 20813 39646 20879 39647
rect 20813 39614 20814 39646
rect 20808 39582 20814 39614
rect 20878 39614 20879 39646
rect 21760 39646 21836 39854
rect 20878 39582 20884 39614
rect 20808 39374 20884 39582
rect 21760 39582 21766 39646
rect 21830 39582 21836 39646
rect 22032 39854 22038 39918
rect 22102 39854 22108 39918
rect 22032 39646 22108 39854
rect 22032 39614 22038 39646
rect 21760 39576 21836 39582
rect 22037 39582 22038 39614
rect 22102 39614 22108 39646
rect 22576 39918 22652 39924
rect 22576 39854 22582 39918
rect 22646 39854 22652 39918
rect 22576 39646 22652 39854
rect 109344 39918 109420 40262
rect 109485 40262 109486 40294
rect 109550 40294 109556 40326
rect 114240 40326 114316 40332
rect 109550 40262 109551 40294
rect 109485 40261 109551 40262
rect 114240 40262 114246 40326
rect 114310 40262 114316 40326
rect 114240 40054 114316 40262
rect 114240 40022 114246 40054
rect 114245 39990 114246 40022
rect 114310 40022 114316 40054
rect 114648 40326 114724 40332
rect 114648 40262 114654 40326
rect 114718 40262 114724 40326
rect 115197 40326 115263 40327
rect 115197 40294 115198 40326
rect 114648 40054 114724 40262
rect 115192 40262 115198 40294
rect 115262 40294 115263 40326
rect 115262 40262 115268 40294
rect 115192 40196 115268 40262
rect 115192 40190 115404 40196
rect 115192 40126 115334 40190
rect 115398 40126 115404 40190
rect 115192 40120 115404 40126
rect 114648 40022 114654 40054
rect 114310 39990 114311 40022
rect 114245 39989 114311 39990
rect 114653 39990 114654 40022
rect 114718 40022 114724 40054
rect 114718 39990 114719 40022
rect 114653 39989 114719 39990
rect 109344 39854 109350 39918
rect 109414 39854 109420 39918
rect 114245 39918 114311 39919
rect 114245 39886 114246 39918
rect 109344 39848 109420 39854
rect 114240 39854 114246 39886
rect 114310 39886 114311 39918
rect 114653 39918 114719 39919
rect 114653 39886 114654 39918
rect 114310 39854 114316 39886
rect 22576 39614 22582 39646
rect 22102 39582 22103 39614
rect 22037 39581 22103 39582
rect 22581 39582 22582 39614
rect 22646 39614 22652 39646
rect 114240 39646 114316 39854
rect 22646 39582 22647 39614
rect 22581 39581 22647 39582
rect 114240 39582 114246 39646
rect 114310 39582 114316 39646
rect 114240 39576 114316 39582
rect 114648 39854 114654 39886
rect 114718 39886 114719 39918
rect 115192 39918 115268 39924
rect 114718 39854 114724 39886
rect 114648 39646 114724 39854
rect 114648 39582 114654 39646
rect 114718 39582 114724 39646
rect 115192 39854 115198 39918
rect 115262 39854 115268 39918
rect 115192 39646 115268 39854
rect 115192 39614 115198 39646
rect 114648 39576 114724 39582
rect 115197 39582 115198 39614
rect 115262 39614 115268 39646
rect 115872 39646 115948 39652
rect 115262 39582 115263 39614
rect 115197 39581 115263 39582
rect 115872 39582 115878 39646
rect 115942 39582 115948 39646
rect 20808 39310 20814 39374
rect 20878 39310 20884 39374
rect 20808 39304 20884 39310
rect 27472 39374 27548 39380
rect 27472 39310 27478 39374
rect 27542 39310 27548 39374
rect 20813 39238 20879 39239
rect 20813 39206 20814 39238
rect 952 39038 1230 39102
rect 1294 39038 1300 39102
rect 952 37334 1300 39038
rect 20808 39174 20814 39206
rect 20878 39206 20879 39238
rect 21488 39238 21564 39244
rect 20878 39174 20884 39206
rect 20808 38966 20884 39174
rect 20808 38902 20814 38966
rect 20878 38902 20884 38966
rect 21488 39174 21494 39238
rect 21558 39174 21564 39238
rect 21488 38966 21564 39174
rect 27472 39102 27548 39310
rect 27472 39070 27478 39102
rect 27477 39038 27478 39070
rect 27542 39070 27548 39102
rect 109480 39374 109556 39380
rect 109480 39310 109486 39374
rect 109550 39310 109556 39374
rect 115872 39374 115948 39582
rect 115872 39342 115878 39374
rect 109480 39102 109556 39310
rect 115877 39310 115878 39342
rect 115942 39342 115948 39374
rect 115942 39310 115943 39342
rect 115877 39309 115943 39310
rect 115469 39238 115535 39239
rect 115469 39206 115470 39238
rect 109480 39070 109486 39102
rect 27542 39038 27543 39070
rect 27477 39037 27543 39038
rect 109485 39038 109486 39070
rect 109550 39070 109556 39102
rect 115464 39174 115470 39206
rect 115534 39206 115535 39238
rect 116008 39238 116084 39244
rect 115534 39174 115540 39206
rect 109550 39038 109551 39070
rect 109485 39037 109551 39038
rect 21488 38934 21494 38966
rect 20808 38896 20884 38902
rect 21493 38902 21494 38934
rect 21558 38934 21564 38966
rect 115464 38966 115540 39174
rect 21558 38902 21559 38934
rect 21493 38901 21559 38902
rect 115464 38902 115470 38966
rect 115534 38902 115540 38966
rect 116008 39174 116014 39238
rect 116078 39174 116084 39238
rect 116008 38966 116084 39174
rect 116008 38934 116014 38966
rect 115464 38896 115540 38902
rect 116013 38902 116014 38934
rect 116078 38934 116084 38966
rect 135320 39102 135668 40806
rect 135320 39038 135326 39102
rect 135390 39038 135668 39102
rect 116078 38902 116079 38934
rect 116013 38901 116079 38902
rect 20808 38830 20884 38836
rect 20808 38766 20814 38830
rect 20878 38766 20884 38830
rect 116013 38830 116079 38831
rect 116013 38798 116014 38830
rect 20808 38558 20884 38766
rect 20808 38526 20814 38558
rect 20813 38494 20814 38526
rect 20878 38526 20884 38558
rect 116008 38766 116014 38798
rect 116078 38798 116079 38830
rect 116078 38766 116084 38798
rect 116008 38558 116084 38766
rect 20878 38494 20879 38526
rect 20813 38493 20879 38494
rect 116008 38494 116014 38558
rect 116078 38494 116084 38558
rect 116008 38488 116084 38494
rect 20813 38422 20879 38423
rect 20813 38390 20814 38422
rect 20808 38358 20814 38390
rect 20878 38390 20879 38422
rect 21352 38422 21428 38428
rect 20878 38358 20884 38390
rect 20808 38150 20884 38358
rect 20808 38086 20814 38150
rect 20878 38086 20884 38150
rect 21352 38358 21358 38422
rect 21422 38358 21428 38422
rect 22037 38422 22103 38423
rect 22037 38390 22038 38422
rect 21352 38150 21428 38358
rect 21352 38118 21358 38150
rect 20808 38080 20884 38086
rect 21357 38086 21358 38118
rect 21422 38118 21428 38150
rect 22032 38358 22038 38390
rect 22102 38390 22103 38422
rect 22440 38422 22516 38428
rect 22102 38358 22108 38390
rect 22032 38150 22108 38358
rect 21422 38086 21423 38118
rect 21357 38085 21423 38086
rect 22032 38086 22038 38150
rect 22102 38086 22108 38150
rect 22440 38358 22446 38422
rect 22510 38358 22516 38422
rect 114381 38422 114447 38423
rect 114381 38390 114382 38422
rect 22440 38150 22516 38358
rect 114376 38358 114382 38390
rect 114446 38390 114447 38422
rect 114648 38422 114724 38428
rect 114446 38358 114452 38390
rect 22440 38118 22446 38150
rect 22032 38080 22108 38086
rect 22445 38086 22446 38118
rect 22510 38118 22516 38150
rect 27336 38150 27412 38156
rect 22510 38086 22511 38118
rect 22445 38085 22511 38086
rect 27336 38086 27342 38150
rect 27406 38086 27412 38150
rect 109485 38150 109551 38151
rect 109485 38118 109486 38150
rect 20944 38014 21020 38020
rect 20944 37950 20950 38014
rect 21014 37950 21020 38014
rect 21765 38014 21831 38015
rect 21765 37982 21766 38014
rect 20944 37742 21020 37950
rect 20944 37710 20950 37742
rect 20949 37678 20950 37710
rect 21014 37710 21020 37742
rect 21760 37950 21766 37982
rect 21830 37982 21831 38014
rect 22168 38014 22244 38020
rect 21830 37950 21836 37982
rect 21760 37742 21836 37950
rect 21014 37678 21015 37710
rect 20949 37677 21015 37678
rect 21760 37678 21766 37742
rect 21830 37678 21836 37742
rect 22168 37950 22174 38014
rect 22238 37950 22244 38014
rect 22445 38014 22511 38015
rect 22445 37982 22446 38014
rect 22168 37742 22244 37950
rect 22168 37710 22174 37742
rect 21760 37672 21836 37678
rect 22173 37678 22174 37710
rect 22238 37710 22244 37742
rect 22440 37950 22446 37982
rect 22510 37982 22511 38014
rect 22510 37950 22516 37982
rect 22440 37742 22516 37950
rect 27336 37878 27412 38086
rect 27336 37846 27342 37878
rect 27341 37814 27342 37846
rect 27406 37846 27412 37878
rect 109480 38086 109486 38118
rect 109550 38118 109551 38150
rect 114376 38150 114452 38358
rect 109550 38086 109556 38118
rect 109480 37878 109556 38086
rect 114376 38086 114382 38150
rect 114446 38086 114452 38150
rect 114648 38358 114654 38422
rect 114718 38358 114724 38422
rect 115197 38422 115263 38423
rect 115197 38390 115198 38422
rect 114648 38150 114724 38358
rect 114648 38118 114654 38150
rect 114376 38080 114452 38086
rect 114653 38086 114654 38118
rect 114718 38118 114724 38150
rect 115192 38358 115198 38390
rect 115262 38390 115263 38422
rect 115333 38422 115399 38423
rect 115333 38390 115334 38422
rect 115262 38358 115268 38390
rect 115192 38150 115268 38358
rect 114718 38086 114719 38118
rect 114653 38085 114719 38086
rect 115192 38086 115198 38150
rect 115262 38086 115268 38150
rect 115192 38080 115268 38086
rect 115328 38358 115334 38390
rect 115398 38390 115399 38422
rect 115877 38422 115943 38423
rect 115877 38390 115878 38422
rect 115398 38358 115404 38390
rect 115328 38150 115404 38358
rect 115328 38086 115334 38150
rect 115398 38086 115404 38150
rect 115328 38080 115404 38086
rect 115872 38358 115878 38390
rect 115942 38390 115943 38422
rect 115942 38358 115948 38390
rect 115872 38150 115948 38358
rect 115872 38086 115878 38150
rect 115942 38086 115948 38150
rect 115872 38080 115948 38086
rect 27406 37814 27407 37846
rect 27341 37813 27407 37814
rect 109480 37814 109486 37878
rect 109550 37814 109556 37878
rect 109480 37808 109556 37814
rect 114240 38014 114316 38020
rect 114240 37950 114246 38014
rect 114310 37950 114316 38014
rect 114653 38014 114719 38015
rect 114653 37982 114654 38014
rect 22238 37678 22239 37710
rect 22173 37677 22239 37678
rect 22440 37678 22446 37742
rect 22510 37678 22516 37742
rect 114240 37742 114316 37950
rect 114240 37710 114246 37742
rect 22440 37672 22516 37678
rect 114245 37678 114246 37710
rect 114310 37710 114316 37742
rect 114648 37950 114654 37982
rect 114718 37982 114719 38014
rect 115056 38014 115132 38020
rect 114718 37950 114724 37982
rect 114648 37742 114724 37950
rect 114310 37678 114311 37710
rect 114245 37677 114311 37678
rect 114648 37678 114654 37742
rect 114718 37678 114724 37742
rect 115056 37950 115062 38014
rect 115126 37950 115132 38014
rect 115469 38014 115535 38015
rect 115469 37982 115470 38014
rect 115056 37742 115132 37950
rect 115056 37710 115062 37742
rect 114648 37672 114724 37678
rect 115061 37678 115062 37710
rect 115126 37710 115132 37742
rect 115464 37950 115470 37982
rect 115534 37982 115535 38014
rect 116013 38014 116079 38015
rect 116013 37982 116014 38014
rect 115534 37950 115540 37982
rect 115464 37742 115540 37950
rect 115126 37678 115127 37710
rect 115061 37677 115127 37678
rect 115464 37678 115470 37742
rect 115534 37678 115540 37742
rect 115464 37672 115540 37678
rect 116008 37950 116014 37982
rect 116078 37982 116079 38014
rect 116078 37950 116084 37982
rect 116008 37742 116084 37950
rect 116008 37678 116014 37742
rect 116078 37678 116084 37742
rect 116008 37672 116084 37678
rect 952 37270 1230 37334
rect 1294 37270 1300 37334
rect 952 35702 1300 37270
rect 952 35638 1230 35702
rect 1294 35638 1300 35702
rect 952 34070 1300 35638
rect 14144 37606 14220 37612
rect 14144 37542 14150 37606
rect 14214 37542 14220 37606
rect 20813 37606 20879 37607
rect 20813 37574 20814 37606
rect 14144 34886 14220 37542
rect 20808 37542 20814 37574
rect 20878 37574 20879 37606
rect 21221 37606 21287 37607
rect 21221 37574 21222 37606
rect 20878 37542 20884 37574
rect 20808 37334 20884 37542
rect 20808 37270 20814 37334
rect 20878 37270 20884 37334
rect 20808 37264 20884 37270
rect 21216 37542 21222 37574
rect 21286 37574 21287 37606
rect 21624 37606 21700 37612
rect 21286 37542 21292 37574
rect 21216 37334 21292 37542
rect 21216 37270 21222 37334
rect 21286 37270 21292 37334
rect 21624 37542 21630 37606
rect 21694 37542 21700 37606
rect 22037 37606 22103 37607
rect 22037 37574 22038 37606
rect 21624 37334 21700 37542
rect 21624 37302 21630 37334
rect 21216 37264 21292 37270
rect 21629 37270 21630 37302
rect 21694 37302 21700 37334
rect 22032 37542 22038 37574
rect 22102 37574 22103 37606
rect 22576 37606 22652 37612
rect 22102 37542 22108 37574
rect 22032 37334 22108 37542
rect 21694 37270 21695 37302
rect 21629 37269 21695 37270
rect 22032 37270 22038 37334
rect 22102 37270 22108 37334
rect 22576 37542 22582 37606
rect 22646 37542 22652 37606
rect 22576 37334 22652 37542
rect 22576 37302 22582 37334
rect 22032 37264 22108 37270
rect 22581 37270 22582 37302
rect 22646 37302 22652 37334
rect 114376 37606 114452 37612
rect 114376 37542 114382 37606
rect 114446 37542 114452 37606
rect 114376 37334 114452 37542
rect 114376 37302 114382 37334
rect 22646 37270 22647 37302
rect 22581 37269 22647 37270
rect 114381 37270 114382 37302
rect 114446 37302 114452 37334
rect 114784 37606 114860 37612
rect 114784 37542 114790 37606
rect 114854 37542 114860 37606
rect 114784 37334 114860 37542
rect 114784 37302 114790 37334
rect 114446 37270 114447 37302
rect 114381 37269 114447 37270
rect 114789 37270 114790 37302
rect 114854 37302 114860 37334
rect 115872 37606 115948 37612
rect 115872 37542 115878 37606
rect 115942 37542 115948 37606
rect 115872 37334 115948 37542
rect 115872 37302 115878 37334
rect 114854 37270 114855 37302
rect 114789 37269 114855 37270
rect 115877 37270 115878 37302
rect 115942 37302 115948 37334
rect 135320 37470 135668 39038
rect 135320 37406 135326 37470
rect 135390 37406 135668 37470
rect 115942 37270 115943 37302
rect 115877 37269 115943 37270
rect 20808 37198 20884 37204
rect 20808 37134 20814 37198
rect 20878 37134 20884 37198
rect 20808 36926 20884 37134
rect 20808 36894 20814 36926
rect 20813 36862 20814 36894
rect 20878 36894 20884 36926
rect 21352 37198 21428 37204
rect 21352 37134 21358 37198
rect 21422 37134 21428 37198
rect 21352 36926 21428 37134
rect 21352 36894 21358 36926
rect 20878 36862 20879 36894
rect 20813 36861 20879 36862
rect 21357 36862 21358 36894
rect 21422 36894 21428 36926
rect 21488 37198 21564 37204
rect 21488 37134 21494 37198
rect 21558 37134 21564 37198
rect 21488 36926 21564 37134
rect 21488 36894 21494 36926
rect 21422 36862 21423 36894
rect 21357 36861 21423 36862
rect 21493 36862 21494 36894
rect 21558 36894 21564 36926
rect 22168 37198 22244 37204
rect 22168 37134 22174 37198
rect 22238 37134 22244 37198
rect 22581 37198 22647 37199
rect 22581 37166 22582 37198
rect 22168 36926 22244 37134
rect 22168 36894 22174 36926
rect 21558 36862 21559 36894
rect 21493 36861 21559 36862
rect 22173 36862 22174 36894
rect 22238 36894 22244 36926
rect 22576 37134 22582 37166
rect 22646 37166 22647 37198
rect 114240 37198 114316 37204
rect 22646 37134 22652 37166
rect 22576 36926 22652 37134
rect 22238 36862 22239 36894
rect 22173 36861 22239 36862
rect 22576 36862 22582 36926
rect 22646 36862 22652 36926
rect 114240 37134 114246 37198
rect 114310 37134 114316 37198
rect 114789 37198 114855 37199
rect 114789 37166 114790 37198
rect 114240 36926 114316 37134
rect 114240 36894 114246 36926
rect 22576 36856 22652 36862
rect 114245 36862 114246 36894
rect 114310 36894 114316 36926
rect 114784 37134 114790 37166
rect 114854 37166 114855 37198
rect 115605 37198 115671 37199
rect 115605 37166 115606 37198
rect 114854 37134 114860 37166
rect 114784 36926 114860 37134
rect 114310 36862 114311 36894
rect 114245 36861 114311 36862
rect 114784 36862 114790 36926
rect 114854 36862 114860 36926
rect 114784 36856 114860 36862
rect 115600 37134 115606 37166
rect 115670 37166 115671 37198
rect 115877 37198 115943 37199
rect 115877 37166 115878 37198
rect 115670 37134 115676 37166
rect 115600 36926 115676 37134
rect 115600 36862 115606 36926
rect 115670 36862 115676 36926
rect 115600 36856 115676 36862
rect 115872 37134 115878 37166
rect 115942 37166 115943 37198
rect 115942 37134 115948 37166
rect 115872 36926 115948 37134
rect 115872 36862 115878 36926
rect 115942 36862 115948 36926
rect 115872 36856 115948 36862
rect 21765 36790 21831 36791
rect 21765 36758 21766 36790
rect 21760 36726 21766 36758
rect 21830 36758 21831 36790
rect 22032 36790 22108 36796
rect 21830 36726 21836 36758
rect 21760 36518 21836 36726
rect 21760 36454 21766 36518
rect 21830 36454 21836 36518
rect 22032 36726 22038 36790
rect 22102 36726 22108 36790
rect 22032 36518 22108 36726
rect 22032 36486 22038 36518
rect 21760 36448 21836 36454
rect 22037 36454 22038 36486
rect 22102 36486 22108 36518
rect 22440 36790 22516 36796
rect 22440 36726 22446 36790
rect 22510 36726 22516 36790
rect 114245 36790 114311 36791
rect 114245 36758 114246 36790
rect 22440 36518 22516 36726
rect 22440 36486 22446 36518
rect 22102 36454 22103 36486
rect 22037 36453 22103 36454
rect 22445 36454 22446 36486
rect 22510 36486 22516 36518
rect 114240 36726 114246 36758
rect 114310 36758 114311 36790
rect 114653 36790 114719 36791
rect 114653 36758 114654 36790
rect 114310 36726 114316 36758
rect 114240 36518 114316 36726
rect 22510 36454 22511 36486
rect 22445 36453 22511 36454
rect 114240 36454 114246 36518
rect 114310 36454 114316 36518
rect 114240 36448 114316 36454
rect 114648 36726 114654 36758
rect 114718 36758 114719 36790
rect 115192 36790 115268 36796
rect 114718 36726 114724 36758
rect 114648 36518 114724 36726
rect 114648 36454 114654 36518
rect 114718 36454 114724 36518
rect 115192 36726 115198 36790
rect 115262 36726 115268 36790
rect 115192 36518 115268 36726
rect 115192 36486 115198 36518
rect 114648 36448 114724 36454
rect 115197 36454 115198 36486
rect 115262 36486 115268 36518
rect 115464 36790 115540 36796
rect 115464 36726 115470 36790
rect 115534 36726 115540 36790
rect 115464 36518 115540 36726
rect 115464 36486 115470 36518
rect 115262 36454 115263 36486
rect 115197 36453 115263 36454
rect 115469 36454 115470 36486
rect 115534 36486 115540 36518
rect 115534 36454 115535 36486
rect 115469 36453 115535 36454
rect 20949 36382 21015 36383
rect 20949 36350 20950 36382
rect 20944 36318 20950 36350
rect 21014 36350 21015 36382
rect 21493 36382 21559 36383
rect 21493 36350 21494 36382
rect 21014 36318 21020 36350
rect 14144 34854 14150 34886
rect 14149 34822 14150 34854
rect 14214 34854 14220 34886
rect 14280 36246 14356 36252
rect 14280 36182 14286 36246
rect 14350 36182 14356 36246
rect 14214 34822 14215 34854
rect 14149 34821 14215 34822
rect 952 34006 1230 34070
rect 1294 34006 1300 34070
rect 952 32438 1300 34006
rect 952 32374 1230 32438
rect 1294 32374 1300 32438
rect 952 30534 1300 32374
rect 14008 34750 14084 34756
rect 14008 34686 14014 34750
rect 14078 34686 14084 34750
rect 14008 32166 14084 34686
rect 14280 33526 14356 36182
rect 20944 36110 21020 36318
rect 20944 36046 20950 36110
rect 21014 36046 21020 36110
rect 20944 36040 21020 36046
rect 21488 36318 21494 36350
rect 21558 36350 21559 36382
rect 21624 36382 21700 36388
rect 21558 36318 21564 36350
rect 21488 36110 21564 36318
rect 21488 36046 21494 36110
rect 21558 36046 21564 36110
rect 21624 36318 21630 36382
rect 21694 36318 21700 36382
rect 22037 36382 22103 36383
rect 22037 36350 22038 36382
rect 21624 36110 21700 36318
rect 21624 36078 21630 36110
rect 21488 36040 21564 36046
rect 21629 36046 21630 36078
rect 21694 36078 21700 36110
rect 22032 36318 22038 36350
rect 22102 36350 22103 36382
rect 22445 36382 22511 36383
rect 22445 36350 22446 36382
rect 22102 36318 22108 36350
rect 22032 36110 22108 36318
rect 21694 36046 21695 36078
rect 21629 36045 21695 36046
rect 22032 36046 22038 36110
rect 22102 36046 22108 36110
rect 22032 36040 22108 36046
rect 22440 36318 22446 36350
rect 22510 36350 22511 36382
rect 114376 36382 114452 36388
rect 22510 36318 22516 36350
rect 22440 36110 22516 36318
rect 22440 36046 22446 36110
rect 22510 36046 22516 36110
rect 114376 36318 114382 36382
rect 114446 36318 114452 36382
rect 114376 36110 114452 36318
rect 114376 36078 114382 36110
rect 22440 36040 22516 36046
rect 114381 36046 114382 36078
rect 114446 36078 114452 36110
rect 114784 36382 114860 36388
rect 114784 36318 114790 36382
rect 114854 36318 114860 36382
rect 114784 36110 114860 36318
rect 114784 36078 114790 36110
rect 114446 36046 114447 36078
rect 114381 36045 114447 36046
rect 114789 36046 114790 36078
rect 114854 36078 114860 36110
rect 115192 36382 115268 36388
rect 115192 36318 115198 36382
rect 115262 36318 115268 36382
rect 115192 36110 115268 36318
rect 115192 36078 115198 36110
rect 114854 36046 114855 36078
rect 114789 36045 114855 36046
rect 115197 36046 115198 36078
rect 115262 36078 115268 36110
rect 115328 36382 115404 36388
rect 115328 36318 115334 36382
rect 115398 36318 115404 36382
rect 116013 36382 116079 36383
rect 116013 36350 116014 36382
rect 115328 36110 115404 36318
rect 115328 36078 115334 36110
rect 115262 36046 115263 36078
rect 115197 36045 115263 36046
rect 115333 36046 115334 36078
rect 115398 36078 115404 36110
rect 116008 36318 116014 36350
rect 116078 36350 116079 36382
rect 116078 36318 116084 36350
rect 116008 36110 116084 36318
rect 115398 36046 115399 36078
rect 115333 36045 115399 36046
rect 116008 36046 116014 36110
rect 116078 36046 116084 36110
rect 116008 36040 116084 36046
rect 21493 35974 21559 35975
rect 21493 35942 21494 35974
rect 21488 35910 21494 35942
rect 21558 35942 21559 35974
rect 22168 35974 22244 35980
rect 21558 35910 21564 35942
rect 20808 35702 20884 35708
rect 20808 35638 20814 35702
rect 20878 35638 20884 35702
rect 20808 35430 20884 35638
rect 21488 35702 21564 35910
rect 21488 35638 21494 35702
rect 21558 35638 21564 35702
rect 22168 35910 22174 35974
rect 22238 35910 22244 35974
rect 22445 35974 22511 35975
rect 22445 35942 22446 35974
rect 22168 35702 22244 35910
rect 22168 35670 22174 35702
rect 21488 35632 21564 35638
rect 22173 35638 22174 35670
rect 22238 35670 22244 35702
rect 22440 35910 22446 35942
rect 22510 35942 22511 35974
rect 114245 35974 114311 35975
rect 114245 35942 114246 35974
rect 22510 35910 22516 35942
rect 22440 35702 22516 35910
rect 22238 35638 22239 35670
rect 22173 35637 22239 35638
rect 22440 35638 22446 35702
rect 22510 35638 22516 35702
rect 22440 35632 22516 35638
rect 114240 35910 114246 35942
rect 114310 35942 114311 35974
rect 114648 35974 114724 35980
rect 114310 35910 114316 35942
rect 114240 35702 114316 35910
rect 114240 35638 114246 35702
rect 114310 35638 114316 35702
rect 114648 35910 114654 35974
rect 114718 35910 114724 35974
rect 115469 35974 115535 35975
rect 115469 35942 115470 35974
rect 114648 35702 114724 35910
rect 114648 35670 114654 35702
rect 114240 35632 114316 35638
rect 114653 35638 114654 35670
rect 114718 35670 114724 35702
rect 115464 35910 115470 35942
rect 115534 35942 115535 35974
rect 115534 35910 115540 35942
rect 115464 35702 115540 35910
rect 114718 35638 114719 35670
rect 114653 35637 114719 35638
rect 115464 35638 115470 35702
rect 115534 35638 115540 35702
rect 115464 35632 115540 35638
rect 115872 35702 115948 35708
rect 115872 35638 115878 35702
rect 115942 35638 115948 35702
rect 21390 35567 21700 35572
rect 21357 35566 21700 35567
rect 21357 35502 21358 35566
rect 21422 35502 21630 35566
rect 21694 35502 21700 35566
rect 21357 35501 21700 35502
rect 21390 35496 21700 35501
rect 20808 35398 20814 35430
rect 20813 35366 20814 35398
rect 20878 35398 20884 35430
rect 115872 35430 115948 35638
rect 115872 35398 115878 35430
rect 20878 35366 20879 35398
rect 20813 35365 20879 35366
rect 115877 35366 115878 35398
rect 115942 35398 115948 35430
rect 135320 35566 135668 37406
rect 135320 35502 135326 35566
rect 135390 35502 135668 35566
rect 115942 35366 115943 35398
rect 115877 35365 115943 35366
rect 20944 35294 21020 35300
rect 20944 35230 20950 35294
rect 21014 35230 21020 35294
rect 21901 35294 21967 35295
rect 21901 35262 21902 35294
rect 20944 35022 21020 35230
rect 20944 34990 20950 35022
rect 20949 34958 20950 34990
rect 21014 34990 21020 35022
rect 21896 35230 21902 35262
rect 21966 35262 21967 35294
rect 27472 35294 27548 35300
rect 21966 35230 21972 35262
rect 21014 34958 21015 34990
rect 20949 34957 21015 34958
rect 20813 34886 20879 34887
rect 20813 34854 20814 34886
rect 20808 34822 20814 34854
rect 20878 34854 20879 34886
rect 21896 34886 21972 35230
rect 27472 35230 27478 35294
rect 27542 35230 27548 35294
rect 27472 35022 27548 35230
rect 115464 35294 115540 35300
rect 115464 35230 115470 35294
rect 115534 35230 115540 35294
rect 27472 34990 27478 35022
rect 27477 34958 27478 34990
rect 27542 34990 27548 35022
rect 109344 35022 109420 35028
rect 27542 34958 27543 34990
rect 27477 34957 27543 34958
rect 109344 34958 109350 35022
rect 109414 34958 109420 35022
rect 20878 34822 20884 34854
rect 20808 34614 20884 34822
rect 21896 34822 21902 34886
rect 21966 34822 21972 34886
rect 21896 34816 21972 34822
rect 109344 34750 109420 34958
rect 115464 34886 115540 35230
rect 115872 35294 115948 35300
rect 115872 35230 115878 35294
rect 115942 35230 115948 35294
rect 115872 35022 115948 35230
rect 115872 34990 115878 35022
rect 115877 34958 115878 34990
rect 115942 34990 115948 35022
rect 115942 34958 115943 34990
rect 115877 34957 115943 34958
rect 115464 34854 115470 34886
rect 115469 34822 115470 34854
rect 115534 34854 115540 34886
rect 116013 34886 116079 34887
rect 116013 34854 116014 34886
rect 115534 34822 115535 34854
rect 115469 34821 115535 34822
rect 116008 34822 116014 34854
rect 116078 34854 116079 34886
rect 116078 34822 116084 34854
rect 109344 34718 109350 34750
rect 109349 34686 109350 34718
rect 109414 34718 109420 34750
rect 109485 34750 109551 34751
rect 109485 34718 109486 34750
rect 109414 34686 109415 34718
rect 109349 34685 109415 34686
rect 109480 34686 109486 34718
rect 109550 34718 109551 34750
rect 109550 34686 109556 34718
rect 20808 34550 20814 34614
rect 20878 34550 20884 34614
rect 20808 34544 20884 34550
rect 20808 34478 20884 34484
rect 20808 34414 20814 34478
rect 20878 34414 20884 34478
rect 20808 34206 20884 34414
rect 20808 34174 20814 34206
rect 20813 34142 20814 34174
rect 20878 34174 20884 34206
rect 21216 34478 21292 34484
rect 21216 34414 21222 34478
rect 21286 34414 21292 34478
rect 21216 34206 21292 34414
rect 21216 34174 21222 34206
rect 20878 34142 20879 34174
rect 20813 34141 20879 34142
rect 21221 34142 21222 34174
rect 21286 34174 21292 34206
rect 22032 34478 22108 34484
rect 22032 34414 22038 34478
rect 22102 34414 22108 34478
rect 22032 34206 22108 34414
rect 22032 34174 22038 34206
rect 21286 34142 21287 34174
rect 21221 34141 21287 34142
rect 22037 34142 22038 34174
rect 22102 34174 22108 34206
rect 22440 34478 22516 34484
rect 22440 34414 22446 34478
rect 22510 34414 22516 34478
rect 22440 34206 22516 34414
rect 109480 34478 109556 34686
rect 116008 34614 116084 34822
rect 116008 34550 116014 34614
rect 116078 34550 116084 34614
rect 116008 34544 116084 34550
rect 109480 34414 109486 34478
rect 109550 34414 109556 34478
rect 114245 34478 114311 34479
rect 114245 34446 114246 34478
rect 109480 34408 109556 34414
rect 114240 34414 114246 34446
rect 114310 34446 114311 34478
rect 114653 34478 114719 34479
rect 114653 34446 114654 34478
rect 114310 34414 114316 34446
rect 22440 34174 22446 34206
rect 22102 34142 22103 34174
rect 22037 34141 22103 34142
rect 22445 34142 22446 34174
rect 22510 34174 22516 34206
rect 109485 34206 109551 34207
rect 109485 34174 109486 34206
rect 22510 34142 22511 34174
rect 22445 34141 22511 34142
rect 109480 34142 109486 34174
rect 109550 34174 109551 34206
rect 114240 34206 114316 34414
rect 109550 34142 109556 34174
rect 20813 34070 20879 34071
rect 20813 34038 20814 34070
rect 20808 34006 20814 34038
rect 20878 34038 20879 34070
rect 21352 34070 21428 34076
rect 20878 34006 20884 34038
rect 20808 33798 20884 34006
rect 20808 33734 20814 33798
rect 20878 33734 20884 33798
rect 21352 34006 21358 34070
rect 21422 34006 21428 34070
rect 22037 34070 22103 34071
rect 22037 34038 22038 34070
rect 21352 33798 21428 34006
rect 21352 33766 21358 33798
rect 20808 33728 20884 33734
rect 21357 33734 21358 33766
rect 21422 33766 21428 33798
rect 22032 34006 22038 34038
rect 22102 34038 22103 34070
rect 22440 34070 22516 34076
rect 22102 34006 22108 34038
rect 22032 33798 22108 34006
rect 21422 33734 21423 33766
rect 21357 33733 21423 33734
rect 22032 33734 22038 33798
rect 22102 33734 22108 33798
rect 22440 34006 22446 34070
rect 22510 34006 22516 34070
rect 22440 33798 22516 34006
rect 109480 33934 109556 34142
rect 114240 34142 114246 34206
rect 114310 34142 114316 34206
rect 114240 34136 114316 34142
rect 114648 34414 114654 34446
rect 114718 34446 114719 34478
rect 115192 34478 115268 34484
rect 114718 34414 114724 34446
rect 114648 34206 114724 34414
rect 114648 34142 114654 34206
rect 114718 34142 114724 34206
rect 115192 34414 115198 34478
rect 115262 34414 115268 34478
rect 115605 34478 115671 34479
rect 115605 34446 115606 34478
rect 115192 34206 115268 34414
rect 115192 34174 115198 34206
rect 114648 34136 114724 34142
rect 115197 34142 115198 34174
rect 115262 34174 115268 34206
rect 115600 34414 115606 34446
rect 115670 34446 115671 34478
rect 116013 34478 116079 34479
rect 116013 34446 116014 34478
rect 115670 34414 115676 34446
rect 115600 34206 115676 34414
rect 115262 34142 115263 34174
rect 115197 34141 115263 34142
rect 115600 34142 115606 34206
rect 115670 34142 115676 34206
rect 115600 34136 115676 34142
rect 116008 34414 116014 34446
rect 116078 34446 116079 34478
rect 116078 34414 116084 34446
rect 116008 34206 116084 34414
rect 116008 34142 116014 34206
rect 116078 34142 116084 34206
rect 116008 34136 116084 34142
rect 109480 33870 109486 33934
rect 109550 33870 109556 33934
rect 109480 33864 109556 33870
rect 114240 34070 114316 34076
rect 114240 34006 114246 34070
rect 114310 34006 114316 34070
rect 114789 34070 114855 34071
rect 114789 34038 114790 34070
rect 22440 33766 22446 33798
rect 22032 33728 22108 33734
rect 22445 33734 22446 33766
rect 22510 33766 22516 33798
rect 114240 33798 114316 34006
rect 114240 33766 114246 33798
rect 22510 33734 22511 33766
rect 22445 33733 22511 33734
rect 114245 33734 114246 33766
rect 114310 33766 114316 33798
rect 114784 34006 114790 34038
rect 114854 34038 114855 34070
rect 115333 34070 115399 34071
rect 115333 34038 115334 34070
rect 114854 34006 114860 34038
rect 114784 33798 114860 34006
rect 114310 33734 114311 33766
rect 114245 33733 114311 33734
rect 114784 33734 114790 33798
rect 114854 33734 114860 33798
rect 114784 33728 114860 33734
rect 115328 34006 115334 34038
rect 115398 34038 115399 34070
rect 115605 34070 115671 34071
rect 115605 34038 115606 34070
rect 115398 34006 115404 34038
rect 115328 33798 115404 34006
rect 115328 33734 115334 33798
rect 115398 33734 115404 33798
rect 115328 33728 115404 33734
rect 115600 34006 115606 34038
rect 115670 34038 115671 34070
rect 116008 34070 116084 34076
rect 115670 34006 115676 34038
rect 115600 33798 115676 34006
rect 115600 33734 115606 33798
rect 115670 33734 115676 33798
rect 116008 34006 116014 34070
rect 116078 34006 116084 34070
rect 116008 33798 116084 34006
rect 116008 33766 116014 33798
rect 115600 33728 115676 33734
rect 116013 33734 116014 33766
rect 116078 33766 116084 33798
rect 135320 33934 135668 35502
rect 135320 33870 135326 33934
rect 135390 33870 135668 33934
rect 116078 33734 116079 33766
rect 116013 33733 116079 33734
rect 20813 33662 20879 33663
rect 20813 33630 20814 33662
rect 14280 33494 14286 33526
rect 14285 33462 14286 33494
rect 14350 33494 14356 33526
rect 20808 33598 20814 33630
rect 20878 33630 20879 33662
rect 21357 33662 21423 33663
rect 21357 33630 21358 33662
rect 20878 33598 20884 33630
rect 14350 33462 14351 33494
rect 14285 33461 14351 33462
rect 14008 32134 14014 32166
rect 14013 32102 14014 32134
rect 14078 32134 14084 32166
rect 14144 33390 14220 33396
rect 14144 33326 14150 33390
rect 14214 33326 14220 33390
rect 14078 32102 14079 32134
rect 14013 32101 14079 32102
rect 14144 32036 14220 33326
rect 20808 33390 20884 33598
rect 20808 33326 20814 33390
rect 20878 33326 20884 33390
rect 20808 33320 20884 33326
rect 21352 33598 21358 33630
rect 21422 33630 21423 33662
rect 21765 33662 21831 33663
rect 21765 33630 21766 33662
rect 21422 33598 21428 33630
rect 21352 33390 21428 33598
rect 21352 33326 21358 33390
rect 21422 33326 21428 33390
rect 21352 33320 21428 33326
rect 21760 33598 21766 33630
rect 21830 33630 21831 33662
rect 22173 33662 22239 33663
rect 22173 33630 22174 33662
rect 21830 33598 21836 33630
rect 21760 33390 21836 33598
rect 21760 33326 21766 33390
rect 21830 33326 21836 33390
rect 21760 33320 21836 33326
rect 22168 33598 22174 33630
rect 22238 33630 22239 33662
rect 22445 33662 22511 33663
rect 22445 33630 22446 33662
rect 22238 33598 22244 33630
rect 22168 33390 22244 33598
rect 22168 33326 22174 33390
rect 22238 33326 22244 33390
rect 22168 33320 22244 33326
rect 22440 33598 22446 33630
rect 22510 33630 22511 33662
rect 114245 33662 114311 33663
rect 114245 33630 114246 33662
rect 22510 33598 22516 33630
rect 22440 33390 22516 33598
rect 22440 33326 22446 33390
rect 22510 33326 22516 33390
rect 22440 33320 22516 33326
rect 114240 33598 114246 33630
rect 114310 33630 114311 33662
rect 114648 33662 114724 33668
rect 114310 33598 114316 33630
rect 114240 33390 114316 33598
rect 114240 33326 114246 33390
rect 114310 33326 114316 33390
rect 114648 33598 114654 33662
rect 114718 33598 114724 33662
rect 115061 33662 115127 33663
rect 115061 33630 115062 33662
rect 114648 33390 114724 33598
rect 114648 33358 114654 33390
rect 114240 33320 114316 33326
rect 114653 33326 114654 33358
rect 114718 33358 114724 33390
rect 115056 33598 115062 33630
rect 115126 33630 115127 33662
rect 115600 33662 115676 33668
rect 115126 33598 115132 33630
rect 115056 33390 115132 33598
rect 114718 33326 114719 33358
rect 114653 33325 114719 33326
rect 115056 33326 115062 33390
rect 115126 33326 115132 33390
rect 115600 33598 115606 33662
rect 115670 33598 115676 33662
rect 116013 33662 116079 33663
rect 116013 33630 116014 33662
rect 115600 33390 115676 33598
rect 115600 33358 115606 33390
rect 115056 33320 115132 33326
rect 115605 33326 115606 33358
rect 115670 33358 115676 33390
rect 116008 33598 116014 33630
rect 116078 33630 116079 33662
rect 116078 33598 116084 33630
rect 116008 33390 116084 33598
rect 115670 33326 115671 33358
rect 115605 33325 115671 33326
rect 116008 33326 116014 33390
rect 116078 33326 116084 33390
rect 116008 33320 116084 33326
rect 20813 33254 20879 33255
rect 20813 33222 20814 33254
rect 20808 33190 20814 33222
rect 20878 33222 20879 33254
rect 21624 33254 21700 33260
rect 20878 33190 20884 33222
rect 20808 32982 20884 33190
rect 20808 32918 20814 32982
rect 20878 32918 20884 32982
rect 21624 33190 21630 33254
rect 21694 33190 21700 33254
rect 21624 32982 21700 33190
rect 21624 32950 21630 32982
rect 20808 32912 20884 32918
rect 21629 32918 21630 32950
rect 21694 32950 21700 32982
rect 22032 33254 22108 33260
rect 22032 33190 22038 33254
rect 22102 33190 22108 33254
rect 22445 33254 22511 33255
rect 22445 33222 22446 33254
rect 22032 32982 22108 33190
rect 22032 32950 22038 32982
rect 21694 32918 21695 32950
rect 21629 32917 21695 32918
rect 22037 32918 22038 32950
rect 22102 32950 22108 32982
rect 22440 33190 22446 33222
rect 22510 33222 22511 33254
rect 114376 33254 114452 33260
rect 22510 33190 22516 33222
rect 22440 32982 22516 33190
rect 22102 32918 22103 32950
rect 22037 32917 22103 32918
rect 22440 32918 22446 32982
rect 22510 32918 22516 32982
rect 114376 33190 114382 33254
rect 114446 33190 114452 33254
rect 114376 32982 114452 33190
rect 114376 32950 114382 32982
rect 22440 32912 22516 32918
rect 114381 32918 114382 32950
rect 114446 32950 114452 32982
rect 114784 33254 114860 33260
rect 114784 33190 114790 33254
rect 114854 33190 114860 33254
rect 114784 32982 114860 33190
rect 114784 32950 114790 32982
rect 114446 32918 114447 32950
rect 114381 32917 114447 32918
rect 114789 32918 114790 32950
rect 114854 32950 114860 32982
rect 115192 33254 115268 33260
rect 115192 33190 115198 33254
rect 115262 33190 115268 33254
rect 115192 32982 115268 33190
rect 115192 32950 115198 32982
rect 114854 32918 114855 32950
rect 114789 32917 114855 32918
rect 115197 32918 115198 32950
rect 115262 32950 115268 32982
rect 115872 33254 115948 33260
rect 115872 33190 115878 33254
rect 115942 33190 115948 33254
rect 115872 32982 115948 33190
rect 115872 32950 115878 32982
rect 115262 32918 115263 32950
rect 115197 32917 115263 32918
rect 115877 32918 115878 32950
rect 115942 32950 115948 32982
rect 115942 32918 115943 32950
rect 115877 32917 115943 32918
rect 20944 32846 21020 32852
rect 20944 32782 20950 32846
rect 21014 32782 21020 32846
rect 21221 32846 21287 32847
rect 21221 32814 21222 32846
rect 20944 32574 21020 32782
rect 20944 32542 20950 32574
rect 20949 32510 20950 32542
rect 21014 32542 21020 32574
rect 21216 32782 21222 32814
rect 21286 32814 21287 32846
rect 22037 32846 22103 32847
rect 22037 32814 22038 32846
rect 21286 32782 21292 32814
rect 21216 32574 21292 32782
rect 21014 32510 21015 32542
rect 20949 32509 21015 32510
rect 21216 32510 21222 32574
rect 21286 32510 21292 32574
rect 21216 32504 21292 32510
rect 22032 32782 22038 32814
rect 22102 32814 22103 32846
rect 22581 32846 22647 32847
rect 22581 32814 22582 32846
rect 22102 32782 22108 32814
rect 22032 32574 22108 32782
rect 22032 32510 22038 32574
rect 22102 32510 22108 32574
rect 22032 32504 22108 32510
rect 22576 32782 22582 32814
rect 22646 32814 22647 32846
rect 114381 32846 114447 32847
rect 114381 32814 114382 32846
rect 22646 32782 22652 32814
rect 22576 32574 22652 32782
rect 22576 32510 22582 32574
rect 22646 32510 22652 32574
rect 22576 32504 22652 32510
rect 114376 32782 114382 32814
rect 114446 32814 114447 32846
rect 114789 32846 114855 32847
rect 114789 32814 114790 32846
rect 114446 32782 114452 32814
rect 114376 32574 114452 32782
rect 114376 32510 114382 32574
rect 114446 32510 114452 32574
rect 114376 32504 114452 32510
rect 114784 32782 114790 32814
rect 114854 32814 114855 32846
rect 115605 32846 115671 32847
rect 115605 32814 115606 32846
rect 114854 32782 114860 32814
rect 114784 32574 114860 32782
rect 114784 32510 114790 32574
rect 114854 32510 114860 32574
rect 114784 32504 114860 32510
rect 115600 32782 115606 32814
rect 115670 32814 115671 32846
rect 115877 32846 115943 32847
rect 115877 32814 115878 32846
rect 115670 32782 115676 32814
rect 115600 32574 115676 32782
rect 115600 32510 115606 32574
rect 115670 32510 115676 32574
rect 115600 32504 115676 32510
rect 115872 32782 115878 32814
rect 115942 32814 115943 32846
rect 115942 32782 115948 32814
rect 115872 32574 115948 32782
rect 115872 32510 115878 32574
rect 115942 32510 115948 32574
rect 115872 32504 115948 32510
rect 20949 32438 21015 32439
rect 20949 32406 20950 32438
rect 20944 32374 20950 32406
rect 21014 32406 21015 32438
rect 21765 32438 21831 32439
rect 21765 32406 21766 32438
rect 21014 32374 21020 32406
rect 20944 32166 21020 32374
rect 20944 32102 20950 32166
rect 21014 32102 21020 32166
rect 20944 32096 21020 32102
rect 21760 32374 21766 32406
rect 21830 32406 21831 32438
rect 22032 32438 22108 32444
rect 21830 32374 21836 32406
rect 21760 32166 21836 32374
rect 21760 32102 21766 32166
rect 21830 32102 21836 32166
rect 22032 32374 22038 32438
rect 22102 32374 22108 32438
rect 22445 32438 22511 32439
rect 22445 32406 22446 32438
rect 22032 32166 22108 32374
rect 22032 32134 22038 32166
rect 21760 32096 21836 32102
rect 22037 32102 22038 32134
rect 22102 32134 22108 32166
rect 22440 32374 22446 32406
rect 22510 32406 22511 32438
rect 114245 32438 114311 32439
rect 114245 32406 114246 32438
rect 22510 32374 22516 32406
rect 22440 32166 22516 32374
rect 22102 32102 22103 32134
rect 22037 32101 22103 32102
rect 22440 32102 22446 32166
rect 22510 32102 22516 32166
rect 22440 32096 22516 32102
rect 114240 32374 114246 32406
rect 114310 32406 114311 32438
rect 114653 32438 114719 32439
rect 114653 32406 114654 32438
rect 114310 32374 114316 32406
rect 114240 32166 114316 32374
rect 114240 32102 114246 32166
rect 114310 32102 114316 32166
rect 114240 32096 114316 32102
rect 114648 32374 114654 32406
rect 114718 32406 114719 32438
rect 115192 32438 115268 32444
rect 114718 32374 114724 32406
rect 114648 32166 114724 32374
rect 114648 32102 114654 32166
rect 114718 32102 114724 32166
rect 115192 32374 115198 32438
rect 115262 32374 115268 32438
rect 115192 32166 115268 32374
rect 115192 32134 115198 32166
rect 114648 32096 114724 32102
rect 115197 32102 115198 32134
rect 115262 32134 115268 32166
rect 115328 32438 115404 32444
rect 115328 32374 115334 32438
rect 115398 32374 115404 32438
rect 115328 32166 115404 32374
rect 115328 32134 115334 32166
rect 115262 32102 115263 32134
rect 115197 32101 115263 32102
rect 115333 32102 115334 32134
rect 115398 32134 115404 32166
rect 115872 32438 115948 32444
rect 115872 32374 115878 32438
rect 115942 32374 115948 32438
rect 115872 32166 115948 32374
rect 115872 32134 115878 32166
rect 115398 32102 115399 32134
rect 115333 32101 115399 32102
rect 115877 32102 115878 32134
rect 115942 32134 115948 32166
rect 135320 32302 135668 33870
rect 135320 32238 135326 32302
rect 135390 32238 135668 32302
rect 115942 32102 115943 32134
rect 115877 32101 115943 32102
rect 14008 31960 14220 32036
rect 21221 32030 21287 32031
rect 21221 31998 21222 32030
rect 21216 31966 21222 31998
rect 21286 31998 21287 32030
rect 21629 32030 21695 32031
rect 21629 31998 21630 32030
rect 21286 31966 21292 31998
rect 14008 30670 14084 31960
rect 14149 31894 14215 31895
rect 14149 31862 14150 31894
rect 14008 30638 14014 30670
rect 14013 30606 14014 30638
rect 14078 30638 14084 30670
rect 14144 31830 14150 31862
rect 14214 31862 14215 31894
rect 14214 31830 14220 31862
rect 14078 30606 14079 30638
rect 14013 30605 14079 30606
rect 952 30470 1230 30534
rect 1294 30470 1300 30534
rect 952 29038 1300 30470
rect 952 28974 1230 29038
rect 1294 28974 1300 29038
rect 952 27270 1300 28974
rect 14008 30534 14084 30540
rect 14008 30470 14014 30534
rect 14078 30470 14084 30534
rect 14008 27814 14084 30470
rect 14144 29310 14220 31830
rect 20949 31758 21015 31759
rect 20949 31726 20950 31758
rect 20944 31694 20950 31726
rect 21014 31726 21015 31758
rect 21216 31758 21292 31966
rect 21014 31694 21020 31726
rect 20944 31486 21020 31694
rect 21216 31694 21222 31758
rect 21286 31694 21292 31758
rect 21216 31688 21292 31694
rect 21624 31966 21630 31998
rect 21694 31998 21695 32030
rect 22037 32030 22103 32031
rect 22037 31998 22038 32030
rect 21694 31966 21700 31998
rect 21624 31758 21700 31966
rect 21624 31694 21630 31758
rect 21694 31694 21700 31758
rect 21624 31688 21700 31694
rect 22032 31966 22038 31998
rect 22102 31998 22103 32030
rect 22576 32030 22652 32036
rect 22102 31966 22108 31998
rect 22032 31758 22108 31966
rect 22032 31694 22038 31758
rect 22102 31694 22108 31758
rect 22576 31966 22582 32030
rect 22646 31966 22652 32030
rect 22576 31758 22652 31966
rect 114376 32030 114452 32036
rect 114376 31966 114382 32030
rect 114446 31966 114452 32030
rect 22576 31726 22582 31758
rect 22032 31688 22108 31694
rect 22581 31694 22582 31726
rect 22646 31726 22652 31758
rect 109480 31894 109556 31900
rect 109480 31830 109486 31894
rect 109550 31830 109556 31894
rect 22646 31694 22647 31726
rect 22581 31693 22647 31694
rect 22173 31622 22239 31623
rect 22173 31590 22174 31622
rect 20944 31422 20950 31486
rect 21014 31422 21020 31486
rect 20944 31416 21020 31422
rect 22168 31558 22174 31590
rect 22238 31590 22239 31622
rect 22445 31622 22511 31623
rect 22445 31590 22446 31622
rect 22238 31558 22244 31590
rect 22168 31350 22244 31558
rect 22168 31286 22174 31350
rect 22238 31286 22244 31350
rect 22168 31280 22244 31286
rect 22440 31558 22446 31590
rect 22510 31590 22511 31622
rect 109349 31622 109415 31623
rect 109349 31590 109350 31622
rect 22510 31558 22516 31590
rect 22440 31350 22516 31558
rect 22440 31286 22446 31350
rect 22510 31286 22516 31350
rect 22440 31280 22516 31286
rect 109344 31558 109350 31590
rect 109414 31590 109415 31622
rect 109480 31622 109556 31830
rect 114376 31758 114452 31966
rect 114376 31726 114382 31758
rect 114381 31694 114382 31726
rect 114446 31726 114452 31758
rect 114784 32030 114860 32036
rect 114784 31966 114790 32030
rect 114854 31966 114860 32030
rect 114784 31758 114860 31966
rect 114784 31726 114790 31758
rect 114446 31694 114447 31726
rect 114381 31693 114447 31694
rect 114789 31694 114790 31726
rect 114854 31726 114860 31758
rect 115872 31758 115948 31764
rect 114854 31694 114855 31726
rect 114789 31693 114855 31694
rect 115872 31694 115878 31758
rect 115942 31694 115948 31758
rect 109480 31590 109486 31622
rect 109414 31558 109420 31590
rect 21765 31214 21831 31215
rect 21765 31182 21766 31214
rect 21760 31150 21766 31182
rect 21830 31182 21831 31214
rect 109344 31214 109420 31558
rect 109485 31558 109486 31590
rect 109550 31590 109556 31622
rect 114245 31622 114311 31623
rect 114245 31590 114246 31622
rect 109550 31558 109551 31590
rect 109485 31557 109551 31558
rect 114240 31558 114246 31590
rect 114310 31590 114311 31622
rect 114653 31622 114719 31623
rect 114653 31590 114654 31622
rect 114310 31558 114316 31590
rect 114240 31350 114316 31558
rect 114240 31286 114246 31350
rect 114310 31286 114316 31350
rect 114240 31280 114316 31286
rect 114648 31558 114654 31590
rect 114718 31590 114719 31622
rect 114718 31558 114724 31590
rect 114648 31350 114724 31558
rect 115872 31486 115948 31694
rect 115872 31454 115878 31486
rect 115877 31422 115878 31454
rect 115942 31454 115948 31486
rect 115942 31422 115943 31454
rect 115877 31421 115943 31422
rect 114648 31286 114654 31350
rect 114718 31286 114724 31350
rect 114648 31280 114724 31286
rect 21830 31150 21836 31182
rect 20813 30942 20879 30943
rect 20813 30910 20814 30942
rect 20808 30878 20814 30910
rect 20878 30910 20879 30942
rect 21760 30942 21836 31150
rect 109344 31150 109350 31214
rect 109414 31150 109420 31214
rect 109344 31144 109420 31150
rect 115464 31214 115540 31220
rect 115464 31150 115470 31214
rect 115534 31150 115540 31214
rect 27341 31078 27407 31079
rect 27341 31046 27342 31078
rect 20878 30878 20884 30910
rect 20808 30670 20884 30878
rect 21760 30878 21766 30942
rect 21830 30878 21836 30942
rect 21760 30872 21836 30878
rect 27336 31014 27342 31046
rect 27406 31046 27407 31078
rect 27406 31014 27412 31046
rect 27336 30806 27412 31014
rect 115464 30942 115540 31150
rect 115464 30910 115470 30942
rect 115469 30878 115470 30910
rect 115534 30910 115540 30942
rect 115872 30942 115948 30948
rect 115534 30878 115535 30910
rect 115469 30877 115535 30878
rect 115872 30878 115878 30942
rect 115942 30878 115948 30942
rect 27336 30742 27342 30806
rect 27406 30742 27412 30806
rect 27336 30736 27412 30742
rect 20808 30606 20814 30670
rect 20878 30606 20884 30670
rect 27477 30670 27543 30671
rect 27477 30638 27478 30670
rect 20808 30600 20884 30606
rect 27472 30606 27478 30638
rect 27542 30638 27543 30670
rect 109349 30670 109415 30671
rect 109349 30638 109350 30670
rect 27542 30606 27548 30638
rect 20813 30534 20879 30535
rect 20813 30502 20814 30534
rect 20808 30470 20814 30502
rect 20878 30502 20879 30534
rect 21352 30534 21428 30540
rect 20878 30470 20884 30502
rect 20808 30262 20884 30470
rect 20808 30198 20814 30262
rect 20878 30198 20884 30262
rect 21352 30470 21358 30534
rect 21422 30470 21428 30534
rect 21352 30262 21428 30470
rect 27472 30398 27548 30606
rect 27472 30334 27478 30398
rect 27542 30334 27548 30398
rect 27472 30328 27548 30334
rect 109344 30606 109350 30638
rect 109414 30638 109415 30670
rect 115872 30670 115948 30878
rect 115872 30638 115878 30670
rect 109414 30606 109420 30638
rect 109344 30398 109420 30606
rect 115877 30606 115878 30638
rect 115942 30638 115948 30670
rect 115942 30606 115943 30638
rect 115877 30605 115943 30606
rect 115469 30534 115535 30535
rect 115469 30502 115470 30534
rect 109344 30334 109350 30398
rect 109414 30334 109420 30398
rect 109344 30328 109420 30334
rect 115464 30470 115470 30502
rect 115534 30502 115535 30534
rect 116008 30534 116084 30540
rect 115534 30470 115540 30502
rect 21352 30230 21358 30262
rect 20808 30192 20884 30198
rect 21357 30198 21358 30230
rect 21422 30230 21428 30262
rect 109344 30262 109420 30268
rect 21422 30198 21423 30230
rect 21357 30197 21423 30198
rect 109344 30198 109350 30262
rect 109414 30198 109420 30262
rect 20949 30126 21015 30127
rect 20949 30094 20950 30126
rect 20944 30062 20950 30094
rect 21014 30094 21015 30126
rect 22173 30126 22239 30127
rect 22173 30094 22174 30126
rect 21014 30062 21020 30094
rect 20944 29854 21020 30062
rect 20944 29790 20950 29854
rect 21014 29790 21020 29854
rect 20944 29784 21020 29790
rect 22168 30062 22174 30094
rect 22238 30094 22239 30126
rect 22581 30126 22647 30127
rect 22581 30094 22582 30126
rect 22238 30062 22244 30094
rect 22168 29854 22244 30062
rect 22168 29790 22174 29854
rect 22238 29790 22244 29854
rect 22168 29784 22244 29790
rect 22576 30062 22582 30094
rect 22646 30094 22647 30126
rect 22646 30062 22652 30094
rect 22576 29854 22652 30062
rect 109344 29990 109420 30198
rect 115464 30262 115540 30470
rect 115464 30198 115470 30262
rect 115534 30198 115540 30262
rect 116008 30470 116014 30534
rect 116078 30470 116084 30534
rect 116008 30262 116084 30470
rect 116008 30230 116014 30262
rect 115464 30192 115540 30198
rect 116013 30198 116014 30230
rect 116078 30230 116084 30262
rect 135320 30534 135668 32238
rect 135320 30470 135326 30534
rect 135390 30470 135668 30534
rect 116078 30198 116079 30230
rect 116013 30197 116079 30198
rect 114245 30126 114311 30127
rect 114245 30094 114246 30126
rect 109344 29958 109350 29990
rect 109349 29926 109350 29958
rect 109414 29958 109420 29990
rect 114240 30062 114246 30094
rect 114310 30094 114311 30126
rect 114653 30126 114719 30127
rect 114653 30094 114654 30126
rect 114310 30062 114316 30094
rect 109414 29926 109415 29958
rect 109349 29925 109415 29926
rect 22576 29790 22582 29854
rect 22646 29790 22652 29854
rect 22576 29784 22652 29790
rect 114240 29854 114316 30062
rect 114240 29790 114246 29854
rect 114310 29790 114316 29854
rect 114240 29784 114316 29790
rect 114648 30062 114654 30094
rect 114718 30094 114719 30126
rect 115872 30126 115948 30132
rect 114718 30062 114724 30094
rect 114648 29854 114724 30062
rect 114648 29790 114654 29854
rect 114718 29790 114724 29854
rect 115872 30062 115878 30126
rect 115942 30062 115948 30126
rect 115872 29854 115948 30062
rect 115872 29822 115878 29854
rect 114648 29784 114724 29790
rect 115877 29790 115878 29822
rect 115942 29822 115948 29854
rect 115942 29790 115943 29822
rect 115877 29789 115943 29790
rect 20808 29718 20884 29724
rect 20808 29654 20814 29718
rect 20878 29654 20884 29718
rect 20808 29446 20884 29654
rect 20808 29414 20814 29446
rect 20813 29382 20814 29414
rect 20878 29414 20884 29446
rect 21488 29718 21564 29724
rect 21488 29654 21494 29718
rect 21558 29654 21564 29718
rect 21765 29718 21831 29719
rect 21765 29686 21766 29718
rect 21488 29446 21564 29654
rect 21488 29414 21494 29446
rect 20878 29382 20879 29414
rect 20813 29381 20879 29382
rect 21493 29382 21494 29414
rect 21558 29414 21564 29446
rect 21760 29654 21766 29686
rect 21830 29686 21831 29718
rect 22037 29718 22103 29719
rect 22037 29686 22038 29718
rect 21830 29654 21836 29686
rect 21760 29446 21836 29654
rect 21558 29382 21559 29414
rect 21493 29381 21559 29382
rect 21760 29382 21766 29446
rect 21830 29382 21836 29446
rect 21760 29376 21836 29382
rect 22032 29654 22038 29686
rect 22102 29686 22103 29718
rect 22440 29718 22516 29724
rect 22102 29654 22108 29686
rect 22032 29446 22108 29654
rect 22032 29382 22038 29446
rect 22102 29382 22108 29446
rect 22440 29654 22446 29718
rect 22510 29654 22516 29718
rect 22440 29446 22516 29654
rect 22440 29414 22446 29446
rect 22032 29376 22108 29382
rect 22445 29382 22446 29414
rect 22510 29414 22516 29446
rect 114240 29718 114316 29724
rect 114240 29654 114246 29718
rect 114310 29654 114316 29718
rect 114240 29446 114316 29654
rect 114240 29414 114246 29446
rect 22510 29382 22511 29414
rect 22445 29381 22511 29382
rect 114245 29382 114246 29414
rect 114310 29414 114316 29446
rect 114648 29718 114724 29724
rect 114648 29654 114654 29718
rect 114718 29654 114724 29718
rect 115333 29718 115399 29719
rect 115333 29686 115334 29718
rect 114648 29446 114724 29654
rect 114648 29414 114654 29446
rect 114310 29382 114311 29414
rect 114245 29381 114311 29382
rect 114653 29382 114654 29414
rect 114718 29414 114724 29446
rect 115328 29654 115334 29686
rect 115398 29686 115399 29718
rect 115464 29718 115540 29724
rect 115398 29654 115404 29686
rect 115328 29446 115404 29654
rect 114718 29382 114719 29414
rect 114653 29381 114719 29382
rect 115328 29382 115334 29446
rect 115398 29382 115404 29446
rect 115464 29654 115470 29718
rect 115534 29654 115540 29718
rect 115877 29718 115943 29719
rect 115877 29686 115878 29718
rect 115464 29446 115540 29654
rect 115464 29414 115470 29446
rect 115328 29376 115404 29382
rect 115469 29382 115470 29414
rect 115534 29414 115540 29446
rect 115872 29654 115878 29686
rect 115942 29686 115943 29718
rect 115942 29654 115948 29686
rect 115872 29446 115948 29654
rect 115534 29382 115535 29414
rect 115469 29381 115535 29382
rect 115872 29382 115878 29446
rect 115942 29382 115948 29446
rect 115872 29376 115948 29382
rect 14144 29246 14150 29310
rect 14214 29246 14220 29310
rect 20813 29310 20879 29311
rect 20813 29278 20814 29310
rect 14144 29240 14220 29246
rect 20808 29246 20814 29278
rect 20878 29278 20879 29310
rect 21765 29310 21831 29311
rect 21765 29278 21766 29310
rect 20878 29246 20884 29278
rect 17821 29174 17887 29175
rect 17821 29142 17822 29174
rect 14008 27782 14014 27814
rect 14013 27750 14014 27782
rect 14078 27782 14084 27814
rect 17816 29110 17822 29142
rect 17886 29142 17887 29174
rect 17886 29110 17892 29142
rect 14078 27750 14079 27782
rect 14013 27749 14079 27750
rect 15917 27678 15983 27679
rect 15917 27646 15918 27678
rect 952 27206 1230 27270
rect 1294 27206 1300 27270
rect 952 25638 1300 27206
rect 15912 27614 15918 27646
rect 15982 27646 15983 27678
rect 15982 27614 15988 27646
rect 952 25574 1230 25638
rect 1294 25574 1300 25638
rect 952 24006 1300 25574
rect 3808 25910 3884 25916
rect 3808 25846 3814 25910
rect 3878 25846 3884 25910
rect 2536 25365 2602 25366
rect 2536 25301 2537 25365
rect 2601 25301 2602 25365
rect 2536 25300 2602 25301
rect 952 23942 1230 24006
rect 1294 23942 1300 24006
rect 2312 24550 2388 24556
rect 2312 24486 2318 24550
rect 2382 24486 2388 24550
rect 2312 24006 2388 24486
rect 2312 23974 2318 24006
rect 952 22374 1300 23942
rect 2317 23942 2318 23974
rect 2382 23974 2388 24006
rect 2382 23942 2383 23974
rect 2317 23941 2383 23942
rect 952 22310 1230 22374
rect 1294 22310 1300 22374
rect 952 20606 1300 22310
rect 952 20542 1230 20606
rect 1294 20542 1300 20606
rect 952 18838 1300 20542
rect 952 18774 1230 18838
rect 1294 18774 1300 18838
rect 952 17070 1300 18774
rect 2539 17959 2599 25300
rect 3808 23326 3884 25846
rect 15912 25094 15988 27614
rect 17816 27542 17892 29110
rect 20808 29038 20884 29246
rect 20808 28974 20814 29038
rect 20878 28974 20884 29038
rect 20808 28968 20884 28974
rect 21760 29246 21766 29278
rect 21830 29278 21831 29310
rect 22168 29310 22244 29316
rect 21830 29246 21836 29278
rect 21760 29038 21836 29246
rect 21760 28974 21766 29038
rect 21830 28974 21836 29038
rect 22168 29246 22174 29310
rect 22238 29246 22244 29310
rect 22168 29038 22244 29246
rect 22168 29006 22174 29038
rect 21760 28968 21836 28974
rect 22173 28974 22174 29006
rect 22238 29006 22244 29038
rect 22576 29310 22652 29316
rect 22576 29246 22582 29310
rect 22646 29246 22652 29310
rect 114245 29310 114311 29311
rect 114245 29278 114246 29310
rect 22576 29038 22652 29246
rect 22576 29006 22582 29038
rect 22238 28974 22239 29006
rect 22173 28973 22239 28974
rect 22581 28974 22582 29006
rect 22646 29006 22652 29038
rect 114240 29246 114246 29278
rect 114310 29278 114311 29310
rect 114653 29310 114719 29311
rect 114653 29278 114654 29310
rect 114310 29246 114316 29278
rect 114240 29038 114316 29246
rect 22646 28974 22647 29006
rect 22581 28973 22647 28974
rect 114240 28974 114246 29038
rect 114310 28974 114316 29038
rect 114240 28968 114316 28974
rect 114648 29246 114654 29278
rect 114718 29278 114719 29310
rect 115061 29310 115127 29311
rect 115061 29278 115062 29310
rect 114718 29246 114724 29278
rect 114648 29038 114724 29246
rect 114648 28974 114654 29038
rect 114718 28974 114724 29038
rect 114648 28968 114724 28974
rect 115056 29246 115062 29278
rect 115126 29278 115127 29310
rect 115328 29310 115404 29316
rect 115126 29246 115132 29278
rect 115056 29038 115132 29246
rect 115056 28974 115062 29038
rect 115126 28974 115132 29038
rect 115328 29246 115334 29310
rect 115398 29246 115404 29310
rect 115328 29038 115404 29246
rect 115328 29006 115334 29038
rect 115056 28968 115132 28974
rect 115333 28974 115334 29006
rect 115398 29006 115404 29038
rect 116008 29310 116084 29316
rect 116008 29246 116014 29310
rect 116078 29246 116084 29310
rect 116008 29038 116084 29246
rect 116008 29006 116014 29038
rect 115398 28974 115399 29006
rect 115333 28973 115399 28974
rect 116013 28974 116014 29006
rect 116078 29006 116084 29038
rect 135320 29038 135668 30470
rect 116078 28974 116079 29006
rect 116013 28973 116079 28974
rect 135320 28974 135326 29038
rect 135390 28974 135668 29038
rect 20944 28902 21020 28908
rect 20944 28838 20950 28902
rect 21014 28838 21020 28902
rect 21221 28902 21287 28903
rect 21221 28870 21222 28902
rect 20944 28630 21020 28838
rect 20944 28598 20950 28630
rect 20949 28566 20950 28598
rect 21014 28598 21020 28630
rect 21216 28838 21222 28870
rect 21286 28870 21287 28902
rect 21624 28902 21700 28908
rect 21286 28838 21292 28870
rect 21216 28630 21292 28838
rect 21014 28566 21015 28598
rect 20949 28565 21015 28566
rect 21216 28566 21222 28630
rect 21286 28566 21292 28630
rect 21624 28838 21630 28902
rect 21694 28838 21700 28902
rect 22037 28902 22103 28903
rect 22037 28870 22038 28902
rect 21624 28630 21700 28838
rect 21624 28598 21630 28630
rect 21216 28560 21292 28566
rect 21629 28566 21630 28598
rect 21694 28598 21700 28630
rect 22032 28838 22038 28870
rect 22102 28870 22103 28902
rect 22576 28902 22652 28908
rect 22102 28838 22108 28870
rect 22032 28630 22108 28838
rect 21694 28566 21695 28598
rect 21629 28565 21695 28566
rect 22032 28566 22038 28630
rect 22102 28566 22108 28630
rect 22576 28838 22582 28902
rect 22646 28838 22652 28902
rect 22576 28630 22652 28838
rect 22576 28598 22582 28630
rect 22032 28560 22108 28566
rect 22581 28566 22582 28598
rect 22646 28598 22652 28630
rect 114376 28902 114452 28908
rect 114376 28838 114382 28902
rect 114446 28838 114452 28902
rect 114376 28630 114452 28838
rect 114376 28598 114382 28630
rect 22646 28566 22647 28598
rect 22581 28565 22647 28566
rect 114381 28566 114382 28598
rect 114446 28598 114452 28630
rect 114784 28902 114860 28908
rect 114784 28838 114790 28902
rect 114854 28838 114860 28902
rect 114784 28630 114860 28838
rect 114784 28598 114790 28630
rect 114446 28566 114447 28598
rect 114381 28565 114447 28566
rect 114789 28566 114790 28598
rect 114854 28598 114860 28630
rect 115192 28902 115268 28908
rect 115192 28838 115198 28902
rect 115262 28838 115268 28902
rect 115877 28902 115943 28903
rect 115877 28870 115878 28902
rect 115192 28630 115268 28838
rect 115192 28598 115198 28630
rect 114854 28566 114855 28598
rect 114789 28565 114855 28566
rect 115197 28566 115198 28598
rect 115262 28598 115268 28630
rect 115872 28838 115878 28870
rect 115942 28870 115943 28902
rect 115942 28838 115948 28870
rect 115872 28630 115948 28838
rect 115262 28566 115263 28598
rect 115197 28565 115263 28566
rect 115872 28566 115878 28630
rect 115942 28566 115948 28630
rect 115872 28560 115948 28566
rect 20949 28494 21015 28495
rect 20949 28462 20950 28494
rect 20944 28430 20950 28462
rect 21014 28462 21015 28494
rect 21352 28494 21428 28500
rect 21014 28430 21020 28462
rect 20944 28222 21020 28430
rect 20944 28158 20950 28222
rect 21014 28158 21020 28222
rect 21352 28430 21358 28494
rect 21422 28430 21428 28494
rect 21352 28222 21428 28430
rect 21352 28190 21358 28222
rect 20944 28152 21020 28158
rect 21357 28158 21358 28190
rect 21422 28190 21428 28222
rect 21488 28494 21564 28500
rect 21488 28430 21494 28494
rect 21558 28430 21564 28494
rect 21488 28222 21564 28430
rect 21488 28190 21494 28222
rect 21422 28158 21423 28190
rect 21357 28157 21423 28158
rect 21493 28158 21494 28190
rect 21558 28190 21564 28222
rect 22168 28494 22244 28500
rect 22168 28430 22174 28494
rect 22238 28430 22244 28494
rect 22168 28222 22244 28430
rect 22168 28190 22174 28222
rect 21558 28158 21559 28190
rect 21493 28157 21559 28158
rect 22173 28158 22174 28190
rect 22238 28190 22244 28222
rect 22440 28494 22516 28500
rect 22440 28430 22446 28494
rect 22510 28430 22516 28494
rect 114381 28494 114447 28495
rect 114381 28462 114382 28494
rect 22440 28222 22516 28430
rect 22440 28190 22446 28222
rect 22238 28158 22239 28190
rect 22173 28157 22239 28158
rect 22445 28158 22446 28190
rect 22510 28190 22516 28222
rect 114376 28430 114382 28462
rect 114446 28462 114447 28494
rect 114789 28494 114855 28495
rect 114789 28462 114790 28494
rect 114446 28430 114452 28462
rect 114376 28222 114452 28430
rect 22510 28158 22511 28190
rect 22445 28157 22511 28158
rect 114376 28158 114382 28222
rect 114446 28158 114452 28222
rect 114376 28152 114452 28158
rect 114784 28430 114790 28462
rect 114854 28462 114855 28494
rect 115605 28494 115671 28495
rect 115605 28462 115606 28494
rect 114854 28430 114860 28462
rect 114784 28222 114860 28430
rect 114784 28158 114790 28222
rect 114854 28158 114860 28222
rect 114784 28152 114860 28158
rect 115600 28430 115606 28462
rect 115670 28462 115671 28494
rect 115877 28494 115943 28495
rect 115877 28462 115878 28494
rect 115670 28430 115676 28462
rect 115600 28222 115676 28430
rect 115600 28158 115606 28222
rect 115670 28158 115676 28222
rect 115600 28152 115676 28158
rect 115872 28430 115878 28462
rect 115942 28462 115943 28494
rect 115942 28430 115948 28462
rect 115872 28222 115948 28430
rect 115872 28158 115878 28222
rect 115942 28158 115948 28222
rect 115872 28152 115948 28158
rect 17816 27478 17822 27542
rect 17886 27478 17892 27542
rect 17816 27472 17892 27478
rect 18904 28086 18980 28092
rect 18904 28022 18910 28086
rect 18974 28022 18980 28086
rect 18904 27406 18980 28022
rect 21760 28086 21836 28092
rect 21760 28022 21766 28086
rect 21830 28022 21836 28086
rect 21760 27814 21836 28022
rect 21760 27782 21766 27814
rect 21765 27750 21766 27782
rect 21830 27782 21836 27814
rect 22032 28086 22108 28092
rect 22032 28022 22038 28086
rect 22102 28022 22108 28086
rect 22445 28086 22511 28087
rect 22445 28054 22446 28086
rect 22032 27814 22108 28022
rect 22032 27782 22038 27814
rect 21830 27750 21831 27782
rect 21765 27749 21831 27750
rect 22037 27750 22038 27782
rect 22102 27782 22108 27814
rect 22440 28022 22446 28054
rect 22510 28054 22511 28086
rect 114376 28086 114452 28092
rect 22510 28022 22516 28054
rect 22440 27814 22516 28022
rect 22102 27750 22103 27782
rect 22037 27749 22103 27750
rect 22440 27750 22446 27814
rect 22510 27750 22516 27814
rect 114376 28022 114382 28086
rect 114446 28022 114452 28086
rect 114376 27814 114452 28022
rect 114376 27782 114382 27814
rect 22440 27744 22516 27750
rect 114381 27750 114382 27782
rect 114446 27782 114452 27814
rect 114784 28086 114860 28092
rect 114784 28022 114790 28086
rect 114854 28022 114860 28086
rect 114784 27814 114860 28022
rect 114784 27782 114790 27814
rect 114446 27750 114447 27782
rect 114381 27749 114447 27750
rect 114789 27750 114790 27782
rect 114854 27782 114860 27814
rect 115192 28086 115268 28092
rect 115192 28022 115198 28086
rect 115262 28022 115268 28086
rect 115192 27814 115268 28022
rect 115192 27782 115198 27814
rect 114854 27750 114855 27782
rect 114789 27749 114855 27750
rect 115197 27750 115198 27782
rect 115262 27782 115268 27814
rect 115262 27750 115263 27782
rect 115197 27749 115263 27750
rect 22037 27678 22103 27679
rect 22037 27646 22038 27678
rect 18904 27374 18910 27406
rect 18909 27342 18910 27374
rect 18974 27374 18980 27406
rect 22032 27614 22038 27646
rect 22102 27646 22103 27678
rect 22576 27678 22652 27684
rect 22102 27614 22108 27646
rect 22032 27406 22108 27614
rect 18974 27342 18975 27374
rect 18909 27341 18975 27342
rect 22032 27342 22038 27406
rect 22102 27342 22108 27406
rect 22576 27614 22582 27678
rect 22646 27614 22652 27678
rect 22576 27406 22652 27614
rect 22576 27374 22582 27406
rect 22032 27336 22108 27342
rect 22581 27342 22582 27374
rect 22646 27374 22652 27406
rect 114376 27678 114452 27684
rect 114376 27614 114382 27678
rect 114446 27614 114452 27678
rect 114376 27406 114452 27614
rect 114376 27374 114382 27406
rect 22646 27342 22647 27374
rect 22581 27341 22647 27342
rect 114381 27342 114382 27374
rect 114446 27374 114452 27406
rect 114784 27678 114860 27684
rect 114784 27614 114790 27678
rect 114854 27614 114860 27678
rect 114784 27406 114860 27614
rect 114784 27374 114790 27406
rect 114446 27342 114447 27374
rect 114381 27341 114447 27342
rect 114789 27342 114790 27374
rect 114854 27374 114860 27406
rect 114854 27342 114855 27374
rect 114789 27341 114855 27342
rect 17413 27270 17479 27271
rect 17413 27238 17414 27270
rect 17408 27206 17414 27238
rect 17478 27238 17479 27270
rect 18360 27270 18436 27276
rect 17478 27206 17484 27238
rect 17408 26726 17484 27206
rect 17408 26662 17414 26726
rect 17478 26662 17484 26726
rect 18360 27206 18366 27270
rect 18430 27206 18436 27270
rect 18360 26726 18436 27206
rect 18360 26694 18366 26726
rect 17408 26656 17484 26662
rect 18365 26662 18366 26694
rect 18430 26694 18436 26726
rect 18632 27270 18708 27276
rect 18632 27206 18638 27270
rect 18702 27206 18708 27270
rect 18632 26726 18708 27206
rect 18632 26694 18638 26726
rect 18430 26662 18431 26694
rect 18365 26661 18431 26662
rect 18637 26662 18638 26694
rect 18702 26694 18708 26726
rect 19040 27270 19116 27276
rect 19040 27206 19046 27270
rect 19110 27206 19116 27270
rect 20677 27270 20743 27271
rect 20677 27238 20678 27270
rect 19040 26726 19116 27206
rect 20672 27206 20678 27238
rect 20742 27238 20743 27270
rect 21352 27270 21428 27276
rect 20742 27206 20748 27238
rect 20672 26862 20748 27206
rect 21352 27206 21358 27270
rect 21422 27206 21428 27270
rect 20672 26798 20678 26862
rect 20742 26798 20748 26862
rect 20672 26792 20748 26798
rect 20808 26998 20884 27004
rect 20808 26934 20814 26998
rect 20878 26934 20884 26998
rect 21352 26998 21428 27206
rect 21352 26966 21358 26998
rect 19040 26694 19046 26726
rect 18702 26662 18703 26694
rect 18637 26661 18703 26662
rect 19045 26662 19046 26694
rect 19110 26694 19116 26726
rect 20808 26726 20884 26934
rect 21357 26934 21358 26966
rect 21422 26966 21428 26998
rect 21488 27270 21564 27276
rect 21488 27206 21494 27270
rect 21558 27206 21564 27270
rect 115605 27270 115671 27271
rect 115605 27238 115606 27270
rect 21488 26998 21564 27206
rect 21488 26966 21494 26998
rect 21422 26934 21423 26966
rect 21357 26933 21423 26934
rect 21493 26934 21494 26966
rect 21558 26966 21564 26998
rect 115600 27206 115606 27238
rect 115670 27238 115671 27270
rect 115741 27270 115807 27271
rect 115741 27238 115742 27270
rect 115670 27206 115676 27238
rect 115600 26998 115676 27206
rect 21558 26934 21559 26966
rect 21493 26933 21559 26934
rect 115600 26934 115606 26998
rect 115670 26934 115676 26998
rect 115600 26928 115676 26934
rect 115736 27206 115742 27238
rect 115806 27238 115807 27270
rect 117640 27270 117716 27276
rect 115806 27206 115812 27238
rect 115736 26862 115812 27206
rect 117640 27206 117646 27270
rect 117710 27206 117716 27270
rect 117781 27270 117847 27271
rect 117781 27238 117782 27270
rect 115736 26798 115742 26862
rect 115806 26798 115812 26862
rect 115736 26792 115812 26798
rect 115872 26998 115948 27004
rect 115872 26934 115878 26998
rect 115942 26934 115948 26998
rect 20808 26694 20814 26726
rect 19110 26662 19111 26694
rect 19045 26661 19111 26662
rect 20813 26662 20814 26694
rect 20878 26694 20884 26726
rect 27341 26726 27407 26727
rect 27341 26694 27342 26726
rect 20878 26662 20879 26694
rect 20813 26661 20879 26662
rect 27336 26662 27342 26694
rect 27406 26694 27407 26726
rect 109344 26726 109420 26732
rect 27406 26662 27412 26694
rect 17549 26590 17615 26591
rect 17549 26558 17550 26590
rect 17544 26526 17550 26558
rect 17614 26558 17615 26590
rect 17685 26590 17751 26591
rect 17685 26558 17686 26590
rect 17614 26526 17620 26558
rect 17544 25910 17620 26526
rect 17680 26526 17686 26558
rect 17750 26558 17751 26590
rect 20813 26590 20879 26591
rect 20813 26558 20814 26590
rect 17750 26526 17756 26558
rect 17680 26318 17756 26526
rect 20808 26526 20814 26558
rect 20878 26558 20879 26590
rect 21221 26590 21287 26591
rect 21221 26558 21222 26590
rect 20878 26526 20884 26558
rect 18229 26454 18295 26455
rect 18229 26422 18230 26454
rect 17680 26254 17686 26318
rect 17750 26254 17756 26318
rect 17680 26248 17756 26254
rect 18224 26390 18230 26422
rect 18294 26422 18295 26454
rect 18637 26454 18703 26455
rect 18637 26422 18638 26454
rect 18294 26390 18300 26422
rect 17544 25846 17550 25910
rect 17614 25846 17620 25910
rect 17544 25840 17620 25846
rect 18224 25910 18300 26390
rect 18224 25846 18230 25910
rect 18294 25846 18300 25910
rect 18224 25840 18300 25846
rect 18632 26390 18638 26422
rect 18702 26422 18703 26454
rect 18702 26390 18708 26422
rect 18632 25910 18708 26390
rect 20808 26318 20884 26526
rect 20808 26254 20814 26318
rect 20878 26254 20884 26318
rect 20808 26248 20884 26254
rect 21216 26526 21222 26558
rect 21286 26558 21287 26590
rect 21896 26590 21972 26596
rect 21286 26526 21292 26558
rect 21216 26318 21292 26526
rect 21216 26254 21222 26318
rect 21286 26254 21292 26318
rect 21896 26526 21902 26590
rect 21966 26526 21972 26590
rect 21896 26318 21972 26526
rect 27336 26454 27412 26662
rect 27336 26390 27342 26454
rect 27406 26390 27412 26454
rect 109344 26662 109350 26726
rect 109414 26662 109420 26726
rect 115872 26726 115948 26934
rect 117640 26862 117716 27206
rect 117640 26830 117646 26862
rect 117645 26798 117646 26830
rect 117710 26830 117716 26862
rect 117776 27206 117782 27238
rect 117846 27238 117847 27270
rect 118184 27270 118260 27276
rect 117846 27206 117852 27238
rect 117710 26798 117711 26830
rect 117645 26797 117711 26798
rect 115872 26694 115878 26726
rect 109344 26454 109420 26662
rect 115877 26662 115878 26694
rect 115942 26694 115948 26726
rect 117776 26726 117852 27206
rect 115942 26662 115943 26694
rect 115877 26661 115943 26662
rect 117776 26662 117782 26726
rect 117846 26662 117852 26726
rect 118184 27206 118190 27270
rect 118254 27206 118260 27270
rect 118184 26726 118260 27206
rect 118184 26694 118190 26726
rect 117776 26656 117852 26662
rect 118189 26662 118190 26694
rect 118254 26694 118260 26726
rect 118728 27270 118940 27276
rect 118728 27206 118870 27270
rect 118934 27206 118940 27270
rect 118728 27200 118940 27206
rect 119272 27270 119348 27276
rect 119272 27206 119278 27270
rect 119342 27206 119348 27270
rect 118728 26726 118804 27200
rect 118728 26694 118734 26726
rect 118254 26662 118255 26694
rect 118189 26661 118255 26662
rect 118733 26662 118734 26694
rect 118798 26694 118804 26726
rect 119272 26726 119348 27206
rect 119272 26694 119278 26726
rect 118798 26662 118799 26694
rect 118733 26661 118799 26662
rect 119277 26662 119278 26694
rect 119342 26694 119348 26726
rect 135320 27270 135668 28974
rect 135320 27206 135326 27270
rect 135390 27206 135668 27270
rect 119342 26662 119343 26694
rect 119277 26661 119343 26662
rect 115469 26590 115535 26591
rect 115469 26558 115470 26590
rect 109344 26422 109350 26454
rect 27336 26384 27412 26390
rect 109349 26390 109350 26422
rect 109414 26422 109420 26454
rect 115464 26526 115470 26558
rect 115534 26558 115535 26590
rect 115877 26590 115943 26591
rect 115877 26558 115878 26590
rect 115534 26526 115540 26558
rect 109414 26390 109415 26422
rect 109349 26389 109415 26390
rect 21896 26286 21902 26318
rect 21216 26248 21292 26254
rect 21901 26254 21902 26286
rect 21966 26286 21972 26318
rect 27477 26318 27543 26319
rect 27477 26286 27478 26318
rect 21966 26254 21967 26286
rect 21901 26253 21967 26254
rect 27472 26254 27478 26286
rect 27542 26286 27543 26318
rect 109349 26318 109415 26319
rect 109349 26286 109350 26318
rect 27542 26254 27548 26286
rect 20813 26182 20879 26183
rect 20813 26150 20814 26182
rect 18632 25846 18638 25910
rect 18702 25846 18708 25910
rect 18632 25840 18708 25846
rect 20808 26118 20814 26150
rect 20878 26150 20879 26182
rect 22168 26182 22244 26188
rect 20878 26118 20884 26150
rect 20808 25910 20884 26118
rect 20808 25846 20814 25910
rect 20878 25846 20884 25910
rect 22168 26118 22174 26182
rect 22238 26118 22244 26182
rect 22168 25910 22244 26118
rect 22168 25878 22174 25910
rect 20808 25840 20884 25846
rect 22173 25846 22174 25878
rect 22238 25878 22244 25910
rect 22576 26182 22652 26188
rect 22576 26118 22582 26182
rect 22646 26118 22652 26182
rect 22576 25910 22652 26118
rect 27472 26046 27548 26254
rect 27472 25982 27478 26046
rect 27542 25982 27548 26046
rect 27472 25976 27548 25982
rect 109344 26254 109350 26286
rect 109414 26286 109415 26318
rect 115464 26318 115540 26526
rect 109414 26254 109420 26286
rect 109344 26046 109420 26254
rect 115464 26254 115470 26318
rect 115534 26254 115540 26318
rect 115464 26248 115540 26254
rect 115872 26526 115878 26558
rect 115942 26558 115943 26590
rect 119000 26590 119076 26596
rect 115942 26526 115948 26558
rect 115872 26318 115948 26526
rect 119000 26526 119006 26590
rect 119070 26526 119076 26590
rect 119277 26590 119343 26591
rect 119277 26558 119278 26590
rect 117645 26454 117711 26455
rect 117645 26422 117646 26454
rect 115872 26254 115878 26318
rect 115942 26254 115948 26318
rect 115872 26248 115948 26254
rect 117640 26390 117646 26422
rect 117710 26422 117711 26454
rect 118189 26454 118255 26455
rect 118189 26422 118190 26454
rect 117710 26390 117716 26422
rect 109344 25982 109350 26046
rect 109414 25982 109420 26046
rect 109344 25976 109420 25982
rect 114240 26182 114316 26188
rect 114240 26118 114246 26182
rect 114310 26118 114316 26182
rect 22576 25878 22582 25910
rect 22238 25846 22239 25878
rect 22173 25845 22239 25846
rect 22581 25846 22582 25878
rect 22646 25878 22652 25910
rect 114240 25910 114316 26118
rect 114240 25878 114246 25910
rect 22646 25846 22647 25878
rect 22581 25845 22647 25846
rect 114245 25846 114246 25878
rect 114310 25878 114316 25910
rect 114648 26182 114724 26188
rect 114648 26118 114654 26182
rect 114718 26118 114724 26182
rect 114648 25910 114724 26118
rect 114648 25878 114654 25910
rect 114310 25846 114311 25878
rect 114245 25845 114311 25846
rect 114653 25846 114654 25878
rect 114718 25878 114724 25910
rect 116008 26182 116084 26188
rect 116008 26118 116014 26182
rect 116078 26118 116084 26182
rect 116008 25910 116084 26118
rect 116008 25878 116014 25910
rect 114718 25846 114719 25878
rect 114653 25845 114719 25846
rect 116013 25846 116014 25878
rect 116078 25878 116084 25910
rect 117640 25910 117716 26390
rect 116078 25846 116079 25878
rect 116013 25845 116079 25846
rect 117640 25846 117646 25910
rect 117710 25846 117716 25910
rect 117640 25840 117716 25846
rect 118184 26390 118190 26422
rect 118254 26422 118255 26454
rect 118254 26390 118260 26422
rect 118184 25910 118260 26390
rect 118184 25846 118190 25910
rect 118254 25846 118260 25910
rect 119000 25910 119076 26526
rect 119000 25878 119006 25910
rect 118184 25840 118260 25846
rect 119005 25846 119006 25878
rect 119070 25878 119076 25910
rect 119272 26526 119278 26558
rect 119342 26558 119343 26590
rect 119342 26526 119348 26558
rect 119272 25910 119348 26526
rect 119070 25846 119071 25878
rect 119005 25845 119071 25846
rect 119272 25846 119278 25910
rect 119342 25846 119348 25910
rect 119272 25840 119348 25846
rect 15912 25030 15918 25094
rect 15982 25030 15988 25094
rect 17408 25774 17484 25780
rect 17408 25710 17414 25774
rect 17478 25710 17484 25774
rect 18229 25774 18295 25775
rect 18229 25742 18230 25774
rect 17408 25094 17484 25710
rect 17408 25062 17414 25094
rect 15912 25024 15988 25030
rect 17413 25030 17414 25062
rect 17478 25062 17484 25094
rect 18224 25710 18230 25742
rect 18294 25742 18295 25774
rect 18773 25774 18839 25775
rect 18773 25742 18774 25774
rect 18294 25710 18300 25742
rect 18224 25094 18300 25710
rect 17478 25030 17479 25062
rect 17413 25029 17479 25030
rect 18224 25030 18230 25094
rect 18294 25030 18300 25094
rect 18224 25024 18300 25030
rect 18768 25710 18774 25742
rect 18838 25742 18839 25774
rect 19176 25774 19252 25780
rect 18838 25710 18844 25742
rect 18768 25094 18844 25710
rect 18768 25030 18774 25094
rect 18838 25030 18844 25094
rect 19176 25710 19182 25774
rect 19246 25710 19252 25774
rect 19176 25094 19252 25710
rect 20808 25774 20884 25780
rect 20808 25710 20814 25774
rect 20878 25710 20884 25774
rect 22173 25774 22239 25775
rect 22173 25742 22174 25774
rect 20808 25502 20884 25710
rect 20808 25470 20814 25502
rect 20813 25438 20814 25470
rect 20878 25470 20884 25502
rect 22168 25710 22174 25742
rect 22238 25742 22239 25774
rect 22576 25774 22652 25780
rect 22238 25710 22244 25742
rect 22168 25502 22244 25710
rect 20878 25438 20879 25470
rect 20813 25437 20879 25438
rect 22168 25438 22174 25502
rect 22238 25438 22244 25502
rect 22576 25710 22582 25774
rect 22646 25710 22652 25774
rect 114245 25774 114311 25775
rect 114245 25742 114246 25774
rect 22576 25502 22652 25710
rect 22576 25470 22582 25502
rect 22168 25432 22244 25438
rect 22581 25438 22582 25470
rect 22646 25470 22652 25502
rect 114240 25710 114246 25742
rect 114310 25742 114311 25774
rect 114784 25774 114860 25780
rect 114310 25710 114316 25742
rect 114240 25502 114316 25710
rect 22646 25438 22647 25470
rect 22581 25437 22647 25438
rect 114240 25438 114246 25502
rect 114310 25438 114316 25502
rect 114784 25710 114790 25774
rect 114854 25710 114860 25774
rect 115061 25774 115127 25775
rect 115061 25742 115062 25774
rect 114784 25502 114860 25710
rect 114784 25470 114790 25502
rect 114240 25432 114316 25438
rect 114789 25438 114790 25470
rect 114854 25470 114860 25502
rect 115056 25710 115062 25742
rect 115126 25742 115127 25774
rect 115605 25774 115671 25775
rect 115605 25742 115606 25774
rect 115126 25710 115132 25742
rect 115056 25502 115132 25710
rect 114854 25438 114855 25470
rect 114789 25437 114855 25438
rect 115056 25438 115062 25502
rect 115126 25438 115132 25502
rect 115056 25432 115132 25438
rect 115600 25710 115606 25742
rect 115670 25742 115671 25774
rect 116013 25774 116079 25775
rect 116013 25742 116014 25774
rect 115670 25710 115676 25742
rect 115600 25502 115676 25710
rect 115600 25438 115606 25502
rect 115670 25438 115676 25502
rect 115600 25432 115676 25438
rect 116008 25710 116014 25742
rect 116078 25742 116079 25774
rect 117640 25774 117716 25780
rect 116078 25710 116084 25742
rect 116008 25502 116084 25710
rect 116008 25438 116014 25502
rect 116078 25438 116084 25502
rect 116008 25432 116084 25438
rect 117640 25710 117646 25774
rect 117710 25710 117716 25774
rect 19176 25062 19182 25094
rect 18768 25024 18844 25030
rect 19181 25030 19182 25062
rect 19246 25062 19252 25094
rect 20808 25366 20884 25372
rect 20808 25302 20814 25366
rect 20878 25302 20884 25366
rect 20808 25094 20884 25302
rect 20808 25062 20814 25094
rect 19246 25030 19247 25062
rect 19181 25029 19247 25030
rect 20813 25030 20814 25062
rect 20878 25062 20884 25094
rect 21352 25366 21428 25372
rect 21352 25302 21358 25366
rect 21422 25302 21428 25366
rect 21352 25094 21428 25302
rect 21352 25062 21358 25094
rect 20878 25030 20879 25062
rect 20813 25029 20879 25030
rect 21357 25030 21358 25062
rect 21422 25062 21428 25094
rect 21488 25366 21564 25372
rect 21488 25302 21494 25366
rect 21558 25302 21564 25366
rect 21765 25366 21831 25367
rect 21765 25334 21766 25366
rect 21488 25094 21564 25302
rect 21488 25062 21494 25094
rect 21422 25030 21423 25062
rect 21357 25029 21423 25030
rect 21493 25030 21494 25062
rect 21558 25062 21564 25094
rect 21760 25302 21766 25334
rect 21830 25334 21831 25366
rect 22168 25366 22244 25372
rect 21830 25302 21836 25334
rect 21760 25094 21836 25302
rect 21558 25030 21559 25062
rect 21493 25029 21559 25030
rect 21760 25030 21766 25094
rect 21830 25030 21836 25094
rect 22168 25302 22174 25366
rect 22238 25302 22244 25366
rect 22445 25366 22511 25367
rect 22445 25334 22446 25366
rect 22168 25094 22244 25302
rect 22168 25062 22174 25094
rect 21760 25024 21836 25030
rect 22173 25030 22174 25062
rect 22238 25062 22244 25094
rect 22440 25302 22446 25334
rect 22510 25334 22511 25366
rect 114240 25366 114316 25372
rect 22510 25302 22516 25334
rect 22440 25094 22516 25302
rect 22238 25030 22239 25062
rect 22173 25029 22239 25030
rect 22440 25030 22446 25094
rect 22510 25030 22516 25094
rect 114240 25302 114246 25366
rect 114310 25302 114316 25366
rect 114240 25094 114316 25302
rect 114240 25062 114246 25094
rect 22440 25024 22516 25030
rect 114245 25030 114246 25062
rect 114310 25062 114316 25094
rect 114648 25366 114724 25372
rect 114648 25302 114654 25366
rect 114718 25302 114724 25366
rect 115197 25366 115263 25367
rect 115197 25334 115198 25366
rect 114648 25094 114724 25302
rect 114648 25062 114654 25094
rect 114310 25030 114311 25062
rect 114245 25029 114311 25030
rect 114653 25030 114654 25062
rect 114718 25062 114724 25094
rect 115192 25302 115198 25334
rect 115262 25334 115263 25366
rect 115464 25366 115540 25372
rect 115262 25302 115268 25334
rect 115192 25094 115268 25302
rect 114718 25030 114719 25062
rect 114653 25029 114719 25030
rect 115192 25030 115198 25094
rect 115262 25030 115268 25094
rect 115464 25302 115470 25366
rect 115534 25302 115540 25366
rect 115877 25366 115943 25367
rect 115877 25334 115878 25366
rect 115464 25094 115540 25302
rect 115464 25062 115470 25094
rect 115192 25024 115268 25030
rect 115469 25030 115470 25062
rect 115534 25062 115540 25094
rect 115872 25302 115878 25334
rect 115942 25334 115943 25366
rect 115942 25302 115948 25334
rect 115872 25094 115948 25302
rect 115534 25030 115535 25062
rect 115469 25029 115535 25030
rect 115872 25030 115878 25094
rect 115942 25030 115948 25094
rect 117640 25094 117716 25710
rect 117640 25062 117646 25094
rect 115872 25024 115948 25030
rect 117645 25030 117646 25062
rect 117710 25062 117716 25094
rect 118184 25774 118260 25780
rect 118184 25710 118190 25774
rect 118254 25710 118260 25774
rect 118184 25094 118260 25710
rect 118184 25062 118190 25094
rect 117710 25030 117711 25062
rect 117645 25029 117711 25030
rect 118189 25030 118190 25062
rect 118254 25062 118260 25094
rect 119000 25774 119076 25780
rect 119000 25710 119006 25774
rect 119070 25710 119076 25774
rect 119413 25774 119479 25775
rect 119413 25742 119414 25774
rect 119000 25094 119076 25710
rect 119000 25062 119006 25094
rect 118254 25030 118255 25062
rect 118189 25029 118255 25030
rect 119005 25030 119006 25062
rect 119070 25062 119076 25094
rect 119408 25710 119414 25742
rect 119478 25742 119479 25774
rect 120773 25774 120839 25775
rect 120773 25742 120774 25774
rect 119478 25710 119484 25742
rect 119408 25094 119484 25710
rect 119070 25030 119071 25062
rect 119005 25029 119071 25030
rect 119408 25030 119414 25094
rect 119478 25030 119484 25094
rect 119408 25024 119484 25030
rect 120768 25710 120774 25742
rect 120838 25742 120839 25774
rect 120838 25710 120844 25742
rect 120768 25094 120844 25710
rect 120768 25030 120774 25094
rect 120838 25030 120844 25094
rect 120768 25024 120844 25030
rect 135320 25502 135668 27206
rect 135320 25438 135326 25502
rect 135390 25438 135668 25502
rect 17685 24958 17751 24959
rect 17685 24926 17686 24958
rect 17680 24894 17686 24926
rect 17750 24926 17751 24958
rect 18229 24958 18295 24959
rect 18229 24926 18230 24958
rect 17750 24894 17756 24926
rect 17680 23462 17756 24894
rect 17680 23398 17686 23462
rect 17750 23398 17756 23462
rect 17680 23392 17756 23398
rect 18224 24894 18230 24926
rect 18294 24926 18295 24958
rect 20813 24958 20879 24959
rect 20813 24926 20814 24958
rect 18294 24894 18300 24926
rect 18224 23462 18300 24894
rect 20808 24894 20814 24926
rect 20878 24926 20879 24958
rect 21896 24958 21972 24964
rect 20878 24894 20884 24926
rect 20808 24686 20884 24894
rect 20808 24622 20814 24686
rect 20878 24622 20884 24686
rect 21896 24894 21902 24958
rect 21966 24894 21972 24958
rect 22173 24958 22239 24959
rect 22173 24926 22174 24958
rect 21896 24686 21972 24894
rect 21896 24654 21902 24686
rect 20808 24616 20884 24622
rect 21901 24622 21902 24654
rect 21966 24654 21972 24686
rect 22168 24894 22174 24926
rect 22238 24926 22239 24958
rect 22576 24958 22652 24964
rect 22238 24894 22244 24926
rect 22168 24686 22244 24894
rect 21966 24622 21967 24654
rect 21901 24621 21967 24622
rect 22168 24622 22174 24686
rect 22238 24622 22244 24686
rect 22576 24894 22582 24958
rect 22646 24894 22652 24958
rect 114245 24958 114311 24959
rect 114245 24926 114246 24958
rect 22576 24686 22652 24894
rect 22576 24654 22582 24686
rect 22168 24616 22244 24622
rect 22581 24622 22582 24654
rect 22646 24654 22652 24686
rect 114240 24894 114246 24926
rect 114310 24926 114311 24958
rect 114653 24958 114719 24959
rect 114653 24926 114654 24958
rect 114310 24894 114316 24926
rect 114240 24686 114316 24894
rect 22646 24622 22647 24654
rect 22581 24621 22647 24622
rect 114240 24622 114246 24686
rect 114310 24622 114316 24686
rect 114240 24616 114316 24622
rect 114648 24894 114654 24926
rect 114718 24926 114719 24958
rect 115056 24958 115132 24964
rect 114718 24894 114724 24926
rect 114648 24686 114724 24894
rect 114648 24622 114654 24686
rect 114718 24622 114724 24686
rect 115056 24894 115062 24958
rect 115126 24894 115132 24958
rect 115469 24958 115535 24959
rect 115469 24926 115470 24958
rect 115056 24686 115132 24894
rect 115056 24654 115062 24686
rect 114648 24616 114724 24622
rect 115061 24622 115062 24654
rect 115126 24654 115132 24686
rect 115464 24894 115470 24926
rect 115534 24926 115535 24958
rect 116008 24958 116084 24964
rect 115534 24894 115540 24926
rect 115464 24686 115540 24894
rect 115126 24622 115127 24654
rect 115061 24621 115127 24622
rect 115464 24622 115470 24686
rect 115534 24622 115540 24686
rect 116008 24894 116014 24958
rect 116078 24894 116084 24958
rect 116008 24686 116084 24894
rect 116008 24654 116014 24686
rect 115464 24616 115540 24622
rect 116013 24622 116014 24654
rect 116078 24654 116084 24686
rect 117640 24958 117716 24964
rect 117640 24894 117646 24958
rect 117710 24894 117716 24958
rect 118189 24958 118255 24959
rect 118189 24926 118190 24958
rect 116078 24622 116079 24654
rect 116013 24621 116079 24622
rect 20944 24550 21020 24556
rect 20944 24486 20950 24550
rect 21014 24486 21020 24550
rect 20944 24278 21020 24486
rect 20944 24246 20950 24278
rect 20949 24214 20950 24246
rect 21014 24246 21020 24278
rect 21624 24550 21700 24556
rect 21624 24486 21630 24550
rect 21694 24486 21700 24550
rect 21624 24278 21700 24486
rect 21624 24246 21630 24278
rect 21014 24214 21015 24246
rect 20949 24213 21015 24214
rect 21629 24214 21630 24246
rect 21694 24246 21700 24278
rect 22032 24550 22108 24556
rect 22032 24486 22038 24550
rect 22102 24486 22108 24550
rect 22445 24550 22511 24551
rect 22445 24518 22446 24550
rect 22032 24278 22108 24486
rect 22032 24246 22038 24278
rect 21694 24214 21695 24246
rect 21629 24213 21695 24214
rect 22037 24214 22038 24246
rect 22102 24246 22108 24278
rect 22440 24486 22446 24518
rect 22510 24518 22511 24550
rect 114381 24550 114447 24551
rect 114381 24518 114382 24550
rect 22510 24486 22516 24518
rect 22440 24278 22516 24486
rect 22102 24214 22103 24246
rect 22037 24213 22103 24214
rect 22440 24214 22446 24278
rect 22510 24214 22516 24278
rect 22440 24208 22516 24214
rect 114376 24486 114382 24518
rect 114446 24518 114447 24550
rect 114784 24550 114860 24556
rect 114446 24486 114452 24518
rect 114376 24278 114452 24486
rect 114376 24214 114382 24278
rect 114446 24214 114452 24278
rect 114784 24486 114790 24550
rect 114854 24486 114860 24550
rect 115877 24550 115943 24551
rect 115877 24518 115878 24550
rect 114784 24278 114860 24486
rect 114784 24246 114790 24278
rect 114376 24208 114452 24214
rect 114789 24214 114790 24246
rect 114854 24246 114860 24278
rect 115872 24486 115878 24518
rect 115942 24518 115943 24550
rect 115942 24486 115948 24518
rect 115872 24278 115948 24486
rect 114854 24214 114855 24246
rect 114789 24213 114855 24214
rect 115872 24214 115878 24278
rect 115942 24214 115948 24278
rect 115872 24208 115948 24214
rect 21221 24142 21287 24143
rect 21221 24110 21222 24142
rect 21216 24078 21222 24110
rect 21286 24110 21287 24142
rect 21488 24142 21564 24148
rect 21286 24078 21292 24110
rect 21216 23870 21292 24078
rect 21216 23806 21222 23870
rect 21286 23806 21292 23870
rect 21488 24078 21494 24142
rect 21558 24078 21564 24142
rect 22037 24142 22103 24143
rect 22037 24110 22038 24142
rect 21488 23870 21564 24078
rect 21488 23838 21494 23870
rect 21216 23800 21292 23806
rect 21493 23806 21494 23838
rect 21558 23838 21564 23870
rect 22032 24078 22038 24110
rect 22102 24110 22103 24142
rect 22440 24142 22516 24148
rect 22102 24078 22108 24110
rect 22032 23870 22108 24078
rect 21558 23806 21559 23838
rect 21493 23805 21559 23806
rect 22032 23806 22038 23870
rect 22102 23806 22108 23870
rect 22440 24078 22446 24142
rect 22510 24078 22516 24142
rect 22440 23870 22516 24078
rect 114240 24142 114316 24148
rect 114240 24078 114246 24142
rect 114310 24078 114316 24142
rect 114789 24142 114855 24143
rect 114789 24110 114790 24142
rect 22440 23838 22446 23870
rect 22032 23800 22108 23806
rect 22445 23806 22446 23838
rect 22510 23838 22516 23870
rect 27608 24006 27684 24012
rect 27608 23942 27614 24006
rect 27678 23942 27684 24006
rect 22510 23806 22511 23838
rect 22445 23805 22511 23806
rect 22173 23734 22239 23735
rect 22173 23702 22174 23734
rect 18224 23398 18230 23462
rect 18294 23398 18300 23462
rect 18224 23392 18300 23398
rect 22168 23670 22174 23702
rect 22238 23702 22239 23734
rect 22440 23734 22516 23740
rect 22238 23670 22244 23702
rect 22168 23462 22244 23670
rect 22168 23398 22174 23462
rect 22238 23398 22244 23462
rect 22440 23670 22446 23734
rect 22510 23670 22516 23734
rect 27477 23734 27543 23735
rect 27477 23702 27478 23734
rect 22440 23462 22516 23670
rect 22440 23430 22446 23462
rect 22168 23392 22244 23398
rect 22445 23398 22446 23430
rect 22510 23430 22516 23462
rect 27472 23670 27478 23702
rect 27542 23702 27543 23734
rect 27608 23734 27684 23942
rect 114240 23870 114316 24078
rect 114240 23838 114246 23870
rect 114245 23806 114246 23838
rect 114310 23838 114316 23870
rect 114784 24078 114790 24110
rect 114854 24110 114855 24142
rect 115197 24142 115263 24143
rect 115197 24110 115198 24142
rect 114854 24078 114860 24110
rect 114784 23870 114860 24078
rect 114310 23806 114311 23838
rect 114245 23805 114311 23806
rect 114784 23806 114790 23870
rect 114854 23806 114860 23870
rect 114784 23800 114860 23806
rect 115192 24078 115198 24110
rect 115262 24110 115263 24142
rect 115605 24142 115671 24143
rect 115605 24110 115606 24142
rect 115262 24078 115268 24110
rect 115192 23870 115268 24078
rect 115192 23806 115198 23870
rect 115262 23806 115268 23870
rect 115192 23800 115268 23806
rect 115600 24078 115606 24110
rect 115670 24110 115671 24142
rect 115670 24078 115676 24110
rect 115600 23870 115676 24078
rect 115600 23806 115606 23870
rect 115670 23806 115676 23870
rect 115600 23800 115676 23806
rect 27608 23702 27614 23734
rect 27542 23670 27548 23702
rect 22510 23398 22511 23430
rect 22445 23397 22511 23398
rect 3808 23294 3814 23326
rect 3813 23262 3814 23294
rect 3878 23294 3884 23326
rect 18224 23326 18300 23332
rect 3878 23262 3879 23294
rect 3813 23261 3879 23262
rect 18224 23262 18230 23326
rect 18294 23262 18300 23326
rect 3813 23190 3879 23191
rect 3813 23158 3814 23190
rect 3808 23126 3814 23158
rect 3878 23158 3879 23190
rect 3878 23126 3884 23158
rect 3133 22238 3199 22239
rect 3133 22206 3134 22238
rect 3128 22174 3134 22206
rect 3198 22206 3199 22238
rect 3198 22174 3204 22206
rect 3128 21830 3204 22174
rect 3128 21766 3134 21830
rect 3198 21766 3204 21830
rect 3128 21760 3204 21766
rect 3677 20470 3743 20471
rect 3677 20438 3678 20470
rect 3672 20406 3678 20438
rect 3742 20438 3743 20470
rect 3808 20470 3884 23126
rect 18224 22782 18300 23262
rect 18224 22750 18230 22782
rect 18229 22718 18230 22750
rect 18294 22750 18300 22782
rect 18632 23326 18708 23332
rect 18632 23262 18638 23326
rect 18702 23262 18708 23326
rect 19045 23326 19111 23327
rect 19045 23294 19046 23326
rect 18632 22782 18708 23262
rect 18632 22750 18638 22782
rect 18294 22718 18295 22750
rect 18229 22717 18295 22718
rect 18637 22718 18638 22750
rect 18702 22750 18708 22782
rect 19040 23262 19046 23294
rect 19110 23294 19111 23326
rect 21357 23326 21423 23327
rect 21357 23294 21358 23326
rect 19110 23262 19116 23294
rect 19040 22782 19116 23262
rect 21352 23262 21358 23294
rect 21422 23294 21423 23326
rect 21629 23326 21695 23327
rect 21629 23294 21630 23326
rect 21422 23262 21428 23294
rect 20949 23054 21015 23055
rect 20949 23022 20950 23054
rect 18702 22718 18703 22750
rect 18637 22717 18703 22718
rect 19040 22718 19046 22782
rect 19110 22718 19116 22782
rect 19040 22712 19116 22718
rect 20944 22990 20950 23022
rect 21014 23022 21015 23054
rect 21352 23054 21428 23262
rect 21624 23262 21630 23294
rect 21694 23294 21695 23326
rect 22032 23326 22108 23332
rect 21694 23262 21700 23294
rect 21014 22990 21020 23022
rect 20944 22782 21020 22990
rect 21352 22990 21358 23054
rect 21422 22990 21428 23054
rect 21493 23054 21559 23055
rect 21493 23022 21494 23054
rect 21352 22984 21428 22990
rect 21488 22990 21494 23022
rect 21558 23022 21559 23054
rect 21624 23054 21700 23262
rect 21558 22990 21564 23022
rect 20944 22718 20950 22782
rect 21014 22718 21020 22782
rect 20944 22712 21020 22718
rect 21488 22782 21564 22990
rect 21624 22990 21630 23054
rect 21694 22990 21700 23054
rect 22032 23262 22038 23326
rect 22102 23262 22108 23326
rect 22032 23054 22108 23262
rect 22032 23022 22038 23054
rect 21624 22984 21700 22990
rect 22037 22990 22038 23022
rect 22102 23022 22108 23054
rect 22576 23326 22652 23332
rect 22576 23262 22582 23326
rect 22646 23262 22652 23326
rect 22576 23054 22652 23262
rect 27472 23326 27548 23670
rect 27613 23670 27614 23702
rect 27678 23702 27684 23734
rect 114245 23734 114311 23735
rect 114245 23702 114246 23734
rect 27678 23670 27679 23702
rect 27613 23669 27679 23670
rect 114240 23670 114246 23702
rect 114310 23702 114311 23734
rect 114784 23734 114860 23740
rect 114310 23670 114316 23702
rect 114240 23462 114316 23670
rect 114240 23398 114246 23462
rect 114310 23398 114316 23462
rect 114784 23670 114790 23734
rect 114854 23670 114860 23734
rect 114784 23462 114860 23670
rect 114784 23430 114790 23462
rect 114240 23392 114316 23398
rect 114789 23398 114790 23430
rect 114854 23430 114860 23462
rect 117640 23462 117716 24894
rect 117640 23430 117646 23462
rect 114854 23398 114855 23430
rect 114789 23397 114855 23398
rect 117645 23398 117646 23430
rect 117710 23430 117716 23462
rect 118184 24894 118190 24926
rect 118254 24926 118255 24958
rect 118254 24894 118260 24926
rect 118184 23462 118260 24894
rect 117710 23398 117711 23430
rect 117645 23397 117711 23398
rect 118184 23398 118190 23462
rect 118254 23398 118260 23462
rect 118184 23392 118260 23398
rect 135320 23870 135668 25438
rect 135320 23806 135326 23870
rect 135390 23806 135668 23870
rect 27472 23262 27478 23326
rect 27542 23262 27548 23326
rect 114381 23326 114447 23327
rect 114381 23294 114382 23326
rect 27472 23256 27548 23262
rect 114376 23262 114382 23294
rect 114446 23294 114447 23326
rect 114789 23326 114855 23327
rect 114789 23294 114790 23326
rect 114446 23262 114452 23294
rect 22576 23022 22582 23054
rect 22102 22990 22103 23022
rect 22037 22989 22103 22990
rect 22581 22990 22582 23022
rect 22646 23022 22652 23054
rect 27336 23190 27412 23196
rect 27336 23126 27342 23190
rect 27406 23126 27412 23190
rect 109349 23190 109415 23191
rect 109349 23158 109350 23190
rect 22646 22990 22647 23022
rect 22581 22989 22647 22990
rect 27336 22918 27412 23126
rect 27336 22886 27342 22918
rect 27341 22854 27342 22886
rect 27406 22886 27412 22918
rect 109344 23126 109350 23158
rect 109414 23158 109415 23190
rect 109414 23126 109420 23158
rect 109344 22918 109420 23126
rect 114376 23054 114452 23262
rect 114376 22990 114382 23054
rect 114446 22990 114452 23054
rect 114376 22984 114452 22990
rect 114784 23262 114790 23294
rect 114854 23294 114855 23326
rect 117640 23326 117716 23332
rect 114854 23262 114860 23294
rect 114784 23054 114860 23262
rect 117640 23262 117646 23326
rect 117710 23262 117716 23326
rect 114784 22990 114790 23054
rect 114854 22990 114860 23054
rect 114784 22984 114860 22990
rect 116008 23054 116084 23060
rect 116008 22990 116014 23054
rect 116078 22990 116084 23054
rect 27406 22854 27407 22886
rect 27341 22853 27407 22854
rect 109344 22854 109350 22918
rect 109414 22854 109420 22918
rect 109344 22848 109420 22854
rect 21488 22718 21494 22782
rect 21558 22718 21564 22782
rect 21488 22712 21564 22718
rect 27472 22782 27548 22788
rect 27472 22718 27478 22782
rect 27542 22718 27548 22782
rect 20813 22646 20879 22647
rect 20813 22614 20814 22646
rect 20808 22582 20814 22614
rect 20878 22614 20879 22646
rect 21624 22646 21700 22652
rect 20878 22582 20884 22614
rect 18360 22510 18436 22516
rect 18360 22446 18366 22510
rect 18430 22446 18436 22510
rect 18360 21150 18436 22446
rect 18360 21118 18366 21150
rect 18365 21086 18366 21118
rect 18430 21118 18436 21150
rect 18632 22510 18708 22516
rect 18632 22446 18638 22510
rect 18702 22446 18708 22510
rect 18632 21150 18708 22446
rect 20808 22374 20884 22582
rect 20808 22310 20814 22374
rect 20878 22310 20884 22374
rect 21624 22582 21630 22646
rect 21694 22582 21700 22646
rect 21624 22374 21700 22582
rect 27472 22510 27548 22718
rect 27472 22478 27478 22510
rect 27477 22446 27478 22478
rect 27542 22478 27548 22510
rect 109480 22782 109556 22788
rect 109480 22718 109486 22782
rect 109550 22718 109556 22782
rect 116008 22782 116084 22990
rect 116008 22750 116014 22782
rect 109480 22510 109556 22718
rect 116013 22718 116014 22750
rect 116078 22750 116084 22782
rect 117640 22782 117716 23262
rect 117640 22750 117646 22782
rect 116078 22718 116079 22750
rect 116013 22717 116079 22718
rect 117645 22718 117646 22750
rect 117710 22750 117716 22782
rect 118048 23326 118124 23332
rect 118048 23262 118054 23326
rect 118118 23262 118124 23326
rect 118048 22782 118124 23262
rect 118592 23326 118668 23332
rect 118592 23262 118598 23326
rect 118662 23262 118668 23326
rect 119005 23326 119071 23327
rect 119005 23294 119006 23326
rect 118048 22750 118054 22782
rect 117710 22718 117711 22750
rect 117645 22717 117711 22718
rect 118053 22718 118054 22750
rect 118118 22750 118124 22782
rect 118320 23054 118396 23060
rect 118320 22990 118326 23054
rect 118390 22990 118396 23054
rect 118320 22782 118396 22990
rect 118320 22750 118326 22782
rect 118118 22718 118119 22750
rect 118053 22717 118119 22718
rect 118325 22718 118326 22750
rect 118390 22750 118396 22782
rect 118592 22782 118668 23262
rect 119000 23262 119006 23294
rect 119070 23294 119071 23326
rect 119070 23262 119076 23294
rect 118869 23054 118935 23055
rect 118869 23022 118870 23054
rect 118592 22750 118598 22782
rect 118390 22718 118391 22750
rect 118325 22717 118391 22718
rect 118597 22718 118598 22750
rect 118662 22750 118668 22782
rect 118864 22990 118870 23022
rect 118934 23022 118935 23054
rect 118934 22990 118940 23022
rect 118864 22782 118940 22990
rect 118662 22718 118663 22750
rect 118597 22717 118663 22718
rect 118864 22718 118870 22782
rect 118934 22718 118940 22782
rect 118864 22712 118940 22718
rect 119000 22782 119076 23262
rect 119000 22718 119006 22782
rect 119070 22718 119076 22782
rect 119000 22712 119076 22718
rect 115061 22646 115127 22647
rect 115061 22614 115062 22646
rect 109480 22478 109486 22510
rect 27542 22446 27543 22478
rect 27477 22445 27543 22446
rect 109485 22446 109486 22478
rect 109550 22478 109556 22510
rect 115056 22582 115062 22614
rect 115126 22614 115127 22646
rect 115872 22646 115948 22652
rect 115126 22582 115132 22614
rect 109550 22446 109551 22478
rect 109485 22445 109551 22446
rect 21624 22342 21630 22374
rect 20808 22304 20884 22310
rect 21629 22310 21630 22342
rect 21694 22342 21700 22374
rect 27341 22374 27407 22375
rect 27341 22342 27342 22374
rect 21694 22310 21695 22342
rect 21629 22309 21695 22310
rect 27336 22310 27342 22342
rect 27406 22342 27407 22374
rect 109344 22374 109420 22380
rect 27406 22310 27412 22342
rect 20944 22238 21020 22244
rect 20944 22174 20950 22238
rect 21014 22174 21020 22238
rect 20944 21966 21020 22174
rect 27336 22102 27412 22310
rect 27336 22038 27342 22102
rect 27406 22038 27412 22102
rect 109344 22310 109350 22374
rect 109414 22310 109420 22374
rect 109344 22102 109420 22310
rect 115056 22374 115132 22582
rect 115056 22310 115062 22374
rect 115126 22310 115132 22374
rect 115872 22582 115878 22646
rect 115942 22582 115948 22646
rect 115872 22374 115948 22582
rect 115872 22342 115878 22374
rect 115056 22304 115132 22310
rect 115877 22310 115878 22342
rect 115942 22342 115948 22374
rect 118456 22510 118532 22516
rect 118456 22446 118462 22510
rect 118526 22446 118532 22510
rect 115942 22310 115943 22342
rect 115877 22309 115943 22310
rect 115877 22238 115943 22239
rect 115877 22206 115878 22238
rect 109344 22070 109350 22102
rect 27336 22032 27412 22038
rect 109349 22038 109350 22070
rect 109414 22070 109420 22102
rect 115872 22174 115878 22206
rect 115942 22206 115943 22238
rect 118320 22238 118396 22244
rect 115942 22174 115948 22206
rect 109414 22038 109415 22070
rect 109349 22037 109415 22038
rect 20944 21934 20950 21966
rect 20949 21902 20950 21934
rect 21014 21934 21020 21966
rect 115872 21966 115948 22174
rect 21014 21902 21015 21934
rect 20949 21901 21015 21902
rect 115872 21902 115878 21966
rect 115942 21902 115948 21966
rect 115872 21896 115948 21902
rect 118320 22174 118326 22238
rect 118390 22174 118396 22238
rect 20944 21830 21020 21836
rect 20944 21766 20950 21830
rect 21014 21766 21020 21830
rect 20944 21558 21020 21766
rect 20944 21526 20950 21558
rect 20949 21494 20950 21526
rect 21014 21526 21020 21558
rect 21352 21830 21428 21836
rect 21352 21766 21358 21830
rect 21422 21766 21428 21830
rect 21352 21558 21428 21766
rect 21352 21526 21358 21558
rect 21014 21494 21015 21526
rect 20949 21493 21015 21494
rect 21357 21494 21358 21526
rect 21422 21526 21428 21558
rect 21488 21830 21564 21836
rect 21488 21766 21494 21830
rect 21558 21766 21564 21830
rect 21488 21558 21564 21766
rect 21488 21526 21494 21558
rect 21422 21494 21423 21526
rect 21357 21493 21423 21494
rect 21493 21494 21494 21526
rect 21558 21526 21564 21558
rect 21760 21830 21836 21836
rect 21760 21766 21766 21830
rect 21830 21766 21836 21830
rect 21760 21558 21836 21766
rect 21760 21526 21766 21558
rect 21558 21494 21559 21526
rect 21493 21493 21559 21494
rect 21765 21494 21766 21526
rect 21830 21526 21836 21558
rect 22168 21830 22244 21836
rect 22168 21766 22174 21830
rect 22238 21766 22244 21830
rect 22445 21830 22511 21831
rect 22445 21798 22446 21830
rect 22168 21558 22244 21766
rect 22168 21526 22174 21558
rect 21830 21494 21831 21526
rect 21765 21493 21831 21494
rect 22173 21494 22174 21526
rect 22238 21526 22244 21558
rect 22440 21766 22446 21798
rect 22510 21798 22511 21830
rect 114245 21830 114311 21831
rect 114245 21798 114246 21830
rect 22510 21766 22516 21798
rect 22440 21558 22516 21766
rect 114240 21766 114246 21798
rect 114310 21798 114311 21830
rect 114648 21830 114724 21836
rect 114310 21766 114316 21798
rect 22238 21494 22239 21526
rect 22173 21493 22239 21494
rect 22440 21494 22446 21558
rect 22510 21494 22516 21558
rect 22440 21488 22516 21494
rect 109344 21558 109420 21564
rect 109344 21494 109350 21558
rect 109414 21494 109420 21558
rect 20949 21422 21015 21423
rect 20949 21390 20950 21422
rect 18632 21118 18638 21150
rect 18430 21086 18431 21118
rect 18365 21085 18431 21086
rect 18637 21086 18638 21118
rect 18702 21118 18708 21150
rect 20944 21358 20950 21390
rect 21014 21390 21015 21422
rect 21629 21422 21695 21423
rect 21629 21390 21630 21422
rect 21014 21358 21020 21390
rect 20944 21150 21020 21358
rect 18702 21086 18703 21118
rect 18637 21085 18703 21086
rect 20944 21086 20950 21150
rect 21014 21086 21020 21150
rect 20944 21080 21020 21086
rect 21624 21358 21630 21390
rect 21694 21390 21695 21422
rect 22173 21422 22239 21423
rect 22173 21390 22174 21422
rect 21694 21358 21700 21390
rect 21624 21150 21700 21358
rect 21624 21086 21630 21150
rect 21694 21086 21700 21150
rect 21624 21080 21700 21086
rect 22168 21358 22174 21390
rect 22238 21390 22239 21422
rect 22440 21422 22516 21428
rect 22238 21358 22244 21390
rect 22168 21150 22244 21358
rect 22168 21086 22174 21150
rect 22238 21086 22244 21150
rect 22440 21358 22446 21422
rect 22510 21358 22516 21422
rect 22440 21150 22516 21358
rect 109344 21286 109420 21494
rect 114240 21558 114316 21766
rect 114240 21494 114246 21558
rect 114310 21494 114316 21558
rect 114648 21766 114654 21830
rect 114718 21766 114724 21830
rect 115061 21830 115127 21831
rect 115061 21798 115062 21830
rect 114648 21558 114724 21766
rect 114648 21526 114654 21558
rect 114240 21488 114316 21494
rect 114653 21494 114654 21526
rect 114718 21526 114724 21558
rect 115056 21766 115062 21798
rect 115126 21798 115127 21830
rect 115600 21830 115676 21836
rect 115126 21766 115132 21798
rect 115056 21558 115132 21766
rect 114718 21494 114719 21526
rect 114653 21493 114719 21494
rect 115056 21494 115062 21558
rect 115126 21494 115132 21558
rect 115600 21766 115606 21830
rect 115670 21766 115676 21830
rect 116013 21830 116079 21831
rect 116013 21798 116014 21830
rect 115600 21558 115676 21766
rect 115600 21526 115606 21558
rect 115056 21488 115132 21494
rect 115605 21494 115606 21526
rect 115670 21526 115676 21558
rect 116008 21766 116014 21798
rect 116078 21798 116079 21830
rect 116078 21766 116084 21798
rect 116008 21558 116084 21766
rect 115670 21494 115671 21526
rect 115605 21493 115671 21494
rect 116008 21494 116014 21558
rect 116078 21494 116084 21558
rect 116008 21488 116084 21494
rect 114245 21422 114311 21423
rect 114245 21390 114246 21422
rect 109344 21254 109350 21286
rect 109349 21222 109350 21254
rect 109414 21254 109420 21286
rect 114240 21358 114246 21390
rect 114310 21390 114311 21422
rect 114653 21422 114719 21423
rect 114653 21390 114654 21422
rect 114310 21358 114316 21390
rect 109414 21222 109415 21254
rect 109349 21221 109415 21222
rect 22440 21118 22446 21150
rect 22168 21080 22244 21086
rect 22445 21086 22446 21118
rect 22510 21118 22516 21150
rect 114240 21150 114316 21358
rect 22510 21086 22511 21118
rect 22445 21085 22511 21086
rect 114240 21086 114246 21150
rect 114310 21086 114316 21150
rect 114240 21080 114316 21086
rect 114648 21358 114654 21390
rect 114718 21390 114719 21422
rect 115605 21422 115671 21423
rect 115605 21390 115606 21422
rect 114718 21358 114724 21390
rect 114648 21150 114724 21358
rect 114648 21086 114654 21150
rect 114718 21086 114724 21150
rect 114648 21080 114724 21086
rect 115600 21358 115606 21390
rect 115670 21390 115671 21422
rect 115872 21422 115948 21428
rect 115670 21358 115676 21390
rect 115600 21150 115676 21358
rect 115600 21086 115606 21150
rect 115670 21086 115676 21150
rect 115872 21358 115878 21422
rect 115942 21358 115948 21422
rect 118053 21422 118119 21423
rect 118053 21390 118054 21422
rect 115872 21150 115948 21358
rect 115872 21118 115878 21150
rect 115600 21080 115676 21086
rect 115877 21086 115878 21118
rect 115942 21118 115948 21150
rect 118048 21358 118054 21390
rect 118118 21390 118119 21422
rect 118118 21358 118124 21390
rect 118048 21150 118124 21358
rect 115942 21086 115943 21118
rect 115877 21085 115943 21086
rect 118048 21086 118054 21150
rect 118118 21086 118124 21150
rect 118320 21150 118396 22174
rect 118456 21286 118532 22446
rect 118864 22510 118940 22516
rect 118864 22446 118870 22510
rect 118934 22446 118940 22510
rect 118864 22238 118940 22446
rect 118864 22206 118870 22238
rect 118869 22174 118870 22206
rect 118934 22206 118940 22238
rect 135320 22238 135668 23806
rect 118934 22174 118935 22206
rect 118869 22173 118935 22174
rect 135320 22174 135326 22238
rect 135390 22174 135668 22238
rect 118456 21254 118462 21286
rect 118461 21222 118462 21254
rect 118526 21254 118532 21286
rect 118526 21222 118527 21254
rect 118461 21221 118527 21222
rect 118320 21118 118326 21150
rect 118048 21080 118124 21086
rect 118325 21086 118326 21118
rect 118390 21118 118396 21150
rect 118390 21086 118391 21118
rect 118325 21085 118391 21086
rect 3742 20406 3748 20438
rect 2536 17958 2602 17959
rect 2536 17894 2537 17958
rect 2601 17894 2602 17958
rect 2536 17893 2602 17894
rect 3672 17614 3748 20406
rect 3808 20406 3814 20470
rect 3878 20406 3884 20470
rect 3808 20400 3884 20406
rect 17816 21014 17892 21020
rect 17816 20950 17822 21014
rect 17886 20950 17892 21014
rect 18365 21014 18431 21015
rect 18365 20982 18366 21014
rect 17816 20334 17892 20950
rect 17816 20302 17822 20334
rect 17821 20270 17822 20302
rect 17886 20302 17892 20334
rect 18360 20950 18366 20982
rect 18430 20982 18431 21014
rect 18637 21014 18703 21015
rect 18637 20982 18638 21014
rect 18430 20950 18436 20982
rect 18360 20334 18436 20950
rect 17886 20270 17887 20302
rect 17821 20269 17887 20270
rect 18360 20270 18366 20334
rect 18430 20270 18436 20334
rect 18360 20264 18436 20270
rect 18632 20950 18638 20982
rect 18702 20982 18703 21014
rect 19176 21014 19252 21020
rect 18702 20950 18708 20982
rect 18632 20334 18708 20950
rect 18632 20270 18638 20334
rect 18702 20270 18708 20334
rect 19176 20950 19182 21014
rect 19246 20950 19252 21014
rect 20813 21014 20879 21015
rect 20813 20982 20814 21014
rect 19176 20334 19252 20950
rect 20808 20950 20814 20982
rect 20878 20982 20879 21014
rect 21352 21014 21428 21020
rect 20878 20950 20884 20982
rect 20808 20742 20884 20950
rect 20808 20678 20814 20742
rect 20878 20678 20884 20742
rect 21352 20950 21358 21014
rect 21422 20950 21428 21014
rect 21765 21014 21831 21015
rect 21765 20982 21766 21014
rect 21352 20742 21428 20950
rect 21352 20710 21358 20742
rect 20808 20672 20884 20678
rect 21357 20678 21358 20710
rect 21422 20710 21428 20742
rect 21760 20950 21766 20982
rect 21830 20982 21831 21014
rect 22037 21014 22103 21015
rect 22037 20982 22038 21014
rect 21830 20950 21836 20982
rect 21760 20742 21836 20950
rect 21422 20678 21423 20710
rect 21357 20677 21423 20678
rect 21760 20678 21766 20742
rect 21830 20678 21836 20742
rect 21760 20672 21836 20678
rect 22032 20950 22038 20982
rect 22102 20982 22103 21014
rect 22445 21014 22511 21015
rect 22445 20982 22446 21014
rect 22102 20950 22108 20982
rect 22032 20742 22108 20950
rect 22032 20678 22038 20742
rect 22102 20678 22108 20742
rect 22032 20672 22108 20678
rect 22440 20950 22446 20982
rect 22510 20982 22511 21014
rect 114240 21014 114316 21020
rect 22510 20950 22516 20982
rect 22440 20742 22516 20950
rect 22440 20678 22446 20742
rect 22510 20678 22516 20742
rect 114240 20950 114246 21014
rect 114310 20950 114316 21014
rect 114240 20742 114316 20950
rect 114240 20710 114246 20742
rect 22440 20672 22516 20678
rect 114245 20678 114246 20710
rect 114310 20710 114316 20742
rect 114648 21014 114724 21020
rect 114648 20950 114654 21014
rect 114718 20950 114724 21014
rect 115197 21014 115263 21015
rect 115197 20982 115198 21014
rect 114648 20742 114724 20950
rect 114648 20710 114654 20742
rect 114310 20678 114311 20710
rect 114245 20677 114311 20678
rect 114653 20678 114654 20710
rect 114718 20710 114724 20742
rect 115192 20950 115198 20982
rect 115262 20982 115263 21014
rect 115333 21014 115399 21015
rect 115333 20982 115334 21014
rect 115262 20950 115268 20982
rect 115192 20742 115268 20950
rect 114718 20678 114719 20710
rect 114653 20677 114719 20678
rect 115192 20678 115198 20742
rect 115262 20678 115268 20742
rect 115192 20672 115268 20678
rect 115328 20950 115334 20982
rect 115398 20982 115399 21014
rect 116008 21014 116084 21020
rect 115398 20950 115404 20982
rect 115328 20742 115404 20950
rect 115328 20678 115334 20742
rect 115398 20678 115404 20742
rect 116008 20950 116014 21014
rect 116078 20950 116084 21014
rect 117645 21014 117711 21015
rect 117645 20982 117646 21014
rect 116008 20742 116084 20950
rect 116008 20710 116014 20742
rect 115328 20672 115404 20678
rect 116013 20678 116014 20710
rect 116078 20710 116084 20742
rect 117640 20950 117646 20982
rect 117710 20982 117711 21014
rect 118184 21014 118260 21020
rect 117710 20950 117716 20982
rect 116078 20678 116079 20710
rect 116013 20677 116079 20678
rect 19176 20302 19182 20334
rect 18632 20264 18708 20270
rect 19181 20270 19182 20302
rect 19246 20302 19252 20334
rect 20944 20606 21020 20612
rect 20944 20542 20950 20606
rect 21014 20542 21020 20606
rect 21357 20606 21423 20607
rect 21357 20574 21358 20606
rect 20944 20334 21020 20542
rect 20944 20302 20950 20334
rect 19246 20270 19247 20302
rect 19181 20269 19247 20270
rect 20949 20270 20950 20302
rect 21014 20302 21020 20334
rect 21352 20542 21358 20574
rect 21422 20574 21423 20606
rect 21765 20606 21831 20607
rect 21765 20574 21766 20606
rect 21422 20542 21428 20574
rect 21352 20334 21428 20542
rect 21014 20270 21015 20302
rect 20949 20269 21015 20270
rect 21352 20270 21358 20334
rect 21422 20270 21428 20334
rect 21352 20264 21428 20270
rect 21760 20542 21766 20574
rect 21830 20574 21831 20606
rect 22168 20606 22244 20612
rect 21830 20542 21836 20574
rect 21760 20334 21836 20542
rect 21760 20270 21766 20334
rect 21830 20270 21836 20334
rect 22168 20542 22174 20606
rect 22238 20542 22244 20606
rect 22445 20606 22511 20607
rect 22445 20574 22446 20606
rect 22168 20334 22244 20542
rect 22168 20302 22174 20334
rect 21760 20264 21836 20270
rect 22173 20270 22174 20302
rect 22238 20302 22244 20334
rect 22440 20542 22446 20574
rect 22510 20574 22511 20606
rect 114240 20606 114316 20612
rect 22510 20542 22516 20574
rect 22440 20334 22516 20542
rect 22238 20270 22239 20302
rect 22173 20269 22239 20270
rect 22440 20270 22446 20334
rect 22510 20270 22516 20334
rect 114240 20542 114246 20606
rect 114310 20542 114316 20606
rect 114240 20334 114316 20542
rect 114240 20302 114246 20334
rect 22440 20264 22516 20270
rect 114245 20270 114246 20302
rect 114310 20302 114316 20334
rect 114648 20606 114724 20612
rect 114648 20542 114654 20606
rect 114718 20542 114724 20606
rect 114648 20334 114724 20542
rect 114648 20302 114654 20334
rect 114310 20270 114311 20302
rect 114245 20269 114311 20270
rect 114653 20270 114654 20302
rect 114718 20302 114724 20334
rect 115056 20606 115132 20612
rect 115056 20542 115062 20606
rect 115126 20542 115132 20606
rect 115469 20606 115535 20607
rect 115469 20574 115470 20606
rect 115056 20334 115132 20542
rect 115056 20302 115062 20334
rect 114718 20270 114719 20302
rect 114653 20269 114719 20270
rect 115061 20270 115062 20302
rect 115126 20302 115132 20334
rect 115464 20542 115470 20574
rect 115534 20574 115535 20606
rect 116013 20606 116079 20607
rect 116013 20574 116014 20606
rect 115534 20542 115540 20574
rect 115464 20334 115540 20542
rect 115126 20270 115127 20302
rect 115061 20269 115127 20270
rect 115464 20270 115470 20334
rect 115534 20270 115540 20334
rect 115464 20264 115540 20270
rect 116008 20542 116014 20574
rect 116078 20574 116079 20606
rect 116078 20542 116084 20574
rect 116008 20334 116084 20542
rect 116008 20270 116014 20334
rect 116078 20270 116084 20334
rect 116008 20264 116084 20270
rect 117640 20334 117716 20950
rect 117640 20270 117646 20334
rect 117710 20270 117716 20334
rect 118184 20950 118190 21014
rect 118254 20950 118260 21014
rect 118184 20334 118260 20950
rect 118184 20302 118190 20334
rect 117640 20264 117716 20270
rect 118189 20270 118190 20302
rect 118254 20302 118260 20334
rect 118592 21014 118668 21020
rect 118592 20950 118598 21014
rect 118662 20950 118668 21014
rect 118592 20334 118668 20950
rect 118592 20302 118598 20334
rect 118254 20270 118255 20302
rect 118189 20269 118255 20270
rect 118597 20270 118598 20302
rect 118662 20302 118668 20334
rect 119000 21014 119076 21020
rect 119000 20950 119006 21014
rect 119070 20950 119076 21014
rect 119000 20334 119076 20950
rect 119000 20302 119006 20334
rect 118662 20270 118663 20302
rect 118597 20269 118663 20270
rect 119005 20270 119006 20302
rect 119070 20302 119076 20334
rect 135320 20606 135668 22174
rect 135320 20542 135326 20606
rect 135390 20542 135668 20606
rect 119070 20270 119071 20302
rect 119005 20269 119071 20270
rect 16592 20198 16668 20204
rect 16592 20134 16598 20198
rect 16662 20134 16668 20198
rect 16592 19110 16668 20134
rect 16592 19078 16598 19110
rect 16597 19046 16598 19078
rect 16662 19078 16668 19110
rect 17000 20198 17076 20204
rect 17000 20134 17006 20198
rect 17070 20134 17076 20198
rect 21085 20198 21151 20199
rect 21085 20166 21086 20198
rect 16662 19046 16663 19078
rect 16597 19045 16663 19046
rect 14693 18838 14759 18839
rect 14693 18806 14694 18838
rect 3672 17550 3678 17614
rect 3742 17550 3748 17614
rect 3672 17544 3748 17550
rect 14688 18774 14694 18806
rect 14758 18806 14759 18838
rect 14758 18774 14764 18806
rect 952 17006 1230 17070
rect 1294 17006 1300 17070
rect 952 15574 1300 17006
rect 14552 17478 14628 17484
rect 14552 17414 14558 17478
rect 14622 17414 14628 17478
rect 952 15510 1230 15574
rect 1294 15510 1300 15574
rect 3128 16118 3204 16124
rect 3128 16054 3134 16118
rect 3198 16054 3204 16118
rect 3128 15574 3204 16054
rect 3128 15542 3134 15574
rect 952 13942 1300 15510
rect 3133 15510 3134 15542
rect 3198 15542 3204 15574
rect 3198 15510 3199 15542
rect 3133 15509 3199 15510
rect 14552 14758 14628 17414
rect 14688 16254 14764 18774
rect 17000 17614 17076 20134
rect 17000 17582 17006 17614
rect 17005 17550 17006 17582
rect 17070 17582 17076 17614
rect 21080 20134 21086 20166
rect 21150 20166 21151 20198
rect 22445 20198 22511 20199
rect 22445 20166 22446 20198
rect 21150 20134 21156 20166
rect 17070 17550 17071 17582
rect 17005 17549 17071 17550
rect 21080 17348 21156 20134
rect 22440 20134 22446 20166
rect 22510 20166 22511 20198
rect 119957 20198 120023 20199
rect 119957 20166 119958 20198
rect 22510 20134 22516 20166
rect 22440 19790 22516 20134
rect 119952 20134 119958 20166
rect 120022 20166 120023 20198
rect 122813 20198 122879 20199
rect 122813 20166 122814 20198
rect 120022 20134 120028 20166
rect 109621 20062 109687 20063
rect 109621 20030 109622 20062
rect 109616 19998 109622 20030
rect 109686 20030 109687 20062
rect 109686 19998 109692 20030
rect 22440 19726 22446 19790
rect 22510 19726 22516 19790
rect 28973 19790 29039 19791
rect 28973 19758 28974 19790
rect 22440 19720 22516 19726
rect 28968 19726 28974 19758
rect 29038 19758 29039 19790
rect 109616 19790 109692 19998
rect 29038 19726 29044 19758
rect 22440 19654 22516 19660
rect 22440 19590 22446 19654
rect 22510 19590 22516 19654
rect 26933 19654 26999 19655
rect 26933 19622 26934 19654
rect 21080 17342 21292 17348
rect 21080 17278 21222 17342
rect 21286 17278 21292 17342
rect 21080 17272 21292 17278
rect 21357 17206 21423 17207
rect 21357 17174 21358 17206
rect 14688 16190 14694 16254
rect 14758 16190 14764 16254
rect 14688 16184 14764 16190
rect 21352 17142 21358 17174
rect 21422 17174 21423 17206
rect 21422 17142 21428 17174
rect 14552 14726 14558 14758
rect 14557 14694 14558 14726
rect 14622 14726 14628 14758
rect 14688 16118 14764 16124
rect 14688 16054 14694 16118
rect 14758 16054 14764 16118
rect 14622 14694 14623 14726
rect 14557 14693 14623 14694
rect 14557 14622 14623 14623
rect 14557 14590 14558 14622
rect 952 13878 1230 13942
rect 1294 13878 1300 13942
rect 952 12310 1300 13878
rect 14552 14558 14558 14590
rect 14622 14590 14623 14622
rect 14622 14558 14628 14590
rect 3133 13806 3199 13807
rect 3133 13774 3134 13806
rect 3128 13742 3134 13774
rect 3198 13774 3199 13806
rect 3198 13742 3204 13774
rect 3128 13398 3204 13742
rect 3128 13334 3134 13398
rect 3198 13334 3204 13398
rect 3128 13328 3204 13334
rect 952 12246 1230 12310
rect 1294 12246 1300 12310
rect 952 10542 1300 12246
rect 14552 12038 14628 14558
rect 14688 13398 14764 16054
rect 21221 15846 21287 15847
rect 21221 15814 21222 15846
rect 21216 15782 21222 15814
rect 21286 15814 21287 15846
rect 21286 15782 21292 15814
rect 14688 13366 14694 13398
rect 14693 13334 14694 13366
rect 14758 13366 14764 13398
rect 20264 14350 20340 14356
rect 20264 14286 20270 14350
rect 20334 14286 20340 14350
rect 14758 13334 14759 13366
rect 14693 13333 14759 13334
rect 14552 11974 14558 12038
rect 14622 11974 14628 12038
rect 14552 11968 14628 11974
rect 14688 13262 14764 13268
rect 14688 13198 14694 13262
rect 14758 13198 14764 13262
rect 952 10478 1230 10542
rect 1294 10478 1300 10542
rect 952 8774 1300 10478
rect 14552 11766 14628 11772
rect 14552 11702 14558 11766
rect 14622 11702 14628 11766
rect 14552 9182 14628 11702
rect 14688 10542 14764 13198
rect 20264 11766 20340 14286
rect 21216 13126 21292 15782
rect 21352 14622 21428 17142
rect 22440 15846 22516 19590
rect 26928 19590 26934 19622
rect 26998 19622 26999 19654
rect 26998 19590 27004 19622
rect 26928 19382 27004 19590
rect 26928 19318 26934 19382
rect 26998 19318 27004 19382
rect 26928 19312 27004 19318
rect 28293 19246 28359 19247
rect 28293 19214 28294 19246
rect 28288 19182 28294 19214
rect 28358 19214 28359 19246
rect 28565 19246 28631 19247
rect 28565 19214 28566 19246
rect 28358 19182 28364 19214
rect 28288 18838 28364 19182
rect 28288 18774 28294 18838
rect 28358 18774 28364 18838
rect 28288 18768 28364 18774
rect 28560 19182 28566 19214
rect 28630 19214 28631 19246
rect 28630 19182 28636 19214
rect 28560 18838 28636 19182
rect 28560 18774 28566 18838
rect 28630 18774 28636 18838
rect 28560 18768 28636 18774
rect 28968 17206 29044 19726
rect 109616 19726 109622 19790
rect 109686 19726 109692 19790
rect 109616 19720 109692 19726
rect 94520 19382 94596 19388
rect 94520 19318 94526 19382
rect 94590 19318 94596 19382
rect 29517 19246 29583 19247
rect 29517 19214 29518 19246
rect 29512 19182 29518 19214
rect 29582 19214 29583 19246
rect 30741 19246 30807 19247
rect 30741 19214 30742 19246
rect 29582 19182 29588 19214
rect 29512 18838 29588 19182
rect 29512 18774 29518 18838
rect 29582 18774 29588 18838
rect 29512 18768 29588 18774
rect 30736 19182 30742 19214
rect 30806 19214 30807 19246
rect 32504 19246 32580 19252
rect 30806 19182 30812 19214
rect 30736 18838 30812 19182
rect 30736 18774 30742 18838
rect 30806 18774 30812 18838
rect 32504 19182 32510 19246
rect 32574 19182 32580 19246
rect 33189 19246 33255 19247
rect 33189 19214 33190 19246
rect 32504 18838 32580 19182
rect 32504 18806 32510 18838
rect 30736 18768 30812 18774
rect 32509 18774 32510 18806
rect 32574 18806 32580 18838
rect 33184 19182 33190 19214
rect 33254 19214 33255 19246
rect 33728 19246 33804 19252
rect 33254 19182 33260 19214
rect 33184 18838 33260 19182
rect 32574 18774 32575 18806
rect 32509 18773 32575 18774
rect 33184 18774 33190 18838
rect 33254 18774 33260 18838
rect 33728 19182 33734 19246
rect 33798 19182 33804 19246
rect 34549 19246 34615 19247
rect 34549 19214 34550 19246
rect 33728 18838 33804 19182
rect 33728 18806 33734 18838
rect 33184 18768 33260 18774
rect 33733 18774 33734 18806
rect 33798 18806 33804 18838
rect 34544 19182 34550 19214
rect 34614 19214 34615 19246
rect 35637 19246 35703 19247
rect 35637 19214 35638 19246
rect 34614 19182 34620 19214
rect 34544 18838 34620 19182
rect 33798 18774 33799 18806
rect 33733 18773 33799 18774
rect 34544 18774 34550 18838
rect 34614 18774 34620 18838
rect 34544 18768 34620 18774
rect 35632 19182 35638 19214
rect 35702 19214 35703 19246
rect 37269 19246 37335 19247
rect 37269 19214 37270 19246
rect 35702 19182 35708 19214
rect 35632 18838 35708 19182
rect 35632 18774 35638 18838
rect 35702 18774 35708 18838
rect 35632 18768 35708 18774
rect 37264 19182 37270 19214
rect 37334 19214 37335 19246
rect 38221 19246 38287 19247
rect 38221 19214 38222 19246
rect 37334 19182 37340 19214
rect 37264 18838 37340 19182
rect 37264 18774 37270 18838
rect 37334 18774 37340 18838
rect 37264 18768 37340 18774
rect 38216 19182 38222 19214
rect 38286 19214 38287 19246
rect 38760 19246 38836 19252
rect 38286 19182 38292 19214
rect 38216 18838 38292 19182
rect 38216 18774 38222 18838
rect 38286 18774 38292 18838
rect 38760 19182 38766 19246
rect 38830 19182 38836 19246
rect 39445 19246 39511 19247
rect 39445 19214 39446 19246
rect 38760 18838 38836 19182
rect 38760 18806 38766 18838
rect 38216 18768 38292 18774
rect 38765 18774 38766 18806
rect 38830 18806 38836 18838
rect 39440 19182 39446 19214
rect 39510 19214 39511 19246
rect 39984 19246 40060 19252
rect 39510 19182 39516 19214
rect 39440 18838 39516 19182
rect 38830 18774 38831 18806
rect 38765 18773 38831 18774
rect 39440 18774 39446 18838
rect 39510 18774 39516 18838
rect 39984 19182 39990 19246
rect 40054 19182 40060 19246
rect 40669 19246 40735 19247
rect 40669 19214 40670 19246
rect 39984 18838 40060 19182
rect 39984 18806 39990 18838
rect 39440 18768 39516 18774
rect 39989 18774 39990 18806
rect 40054 18806 40060 18838
rect 40664 19182 40670 19214
rect 40734 19214 40735 19246
rect 41208 19246 41284 19252
rect 40734 19182 40740 19214
rect 40664 18838 40740 19182
rect 40054 18774 40055 18806
rect 39989 18773 40055 18774
rect 40664 18774 40670 18838
rect 40734 18774 40740 18838
rect 41208 19182 41214 19246
rect 41278 19182 41284 19246
rect 42029 19246 42095 19247
rect 42029 19214 42030 19246
rect 41208 18838 41284 19182
rect 41208 18806 41214 18838
rect 40664 18768 40740 18774
rect 41213 18774 41214 18806
rect 41278 18806 41284 18838
rect 42024 19182 42030 19214
rect 42094 19214 42095 19246
rect 42432 19246 42508 19252
rect 42094 19182 42100 19214
rect 42024 18838 42100 19182
rect 41278 18774 41279 18806
rect 41213 18773 41279 18774
rect 42024 18774 42030 18838
rect 42094 18774 42100 18838
rect 42432 19182 42438 19246
rect 42502 19182 42508 19246
rect 43253 19246 43319 19247
rect 43253 19214 43254 19246
rect 42432 18838 42508 19182
rect 42432 18806 42438 18838
rect 42024 18768 42100 18774
rect 42437 18774 42438 18806
rect 42502 18806 42508 18838
rect 43248 19182 43254 19214
rect 43318 19214 43319 19246
rect 43384 19246 43460 19252
rect 43318 19182 43324 19214
rect 43248 18838 43324 19182
rect 42502 18774 42503 18806
rect 42437 18773 42503 18774
rect 43248 18774 43254 18838
rect 43318 18774 43324 18838
rect 43384 19182 43390 19246
rect 43454 19182 43460 19246
rect 44477 19246 44543 19247
rect 44477 19214 44478 19246
rect 43384 18838 43460 19182
rect 43384 18806 43390 18838
rect 43248 18768 43324 18774
rect 43389 18774 43390 18806
rect 43454 18806 43460 18838
rect 44472 19182 44478 19214
rect 44542 19214 44543 19246
rect 45701 19246 45767 19247
rect 45701 19214 45702 19246
rect 44542 19182 44548 19214
rect 44472 18838 44548 19182
rect 43454 18774 43455 18806
rect 43389 18773 43455 18774
rect 44472 18774 44478 18838
rect 44542 18774 44548 18838
rect 44472 18768 44548 18774
rect 45696 19182 45702 19214
rect 45766 19214 45767 19246
rect 46925 19246 46991 19247
rect 46925 19214 46926 19246
rect 45766 19182 45772 19214
rect 45696 18838 45772 19182
rect 45696 18774 45702 18838
rect 45766 18774 45772 18838
rect 45696 18768 45772 18774
rect 46920 19182 46926 19214
rect 46990 19214 46991 19246
rect 47464 19246 47540 19252
rect 46990 19182 46996 19214
rect 46920 18838 46996 19182
rect 46920 18774 46926 18838
rect 46990 18774 46996 18838
rect 47464 19182 47470 19246
rect 47534 19182 47540 19246
rect 48149 19246 48215 19247
rect 48149 19214 48150 19246
rect 47464 18838 47540 19182
rect 47464 18806 47470 18838
rect 46920 18768 46996 18774
rect 47469 18774 47470 18806
rect 47534 18806 47540 18838
rect 48144 19182 48150 19214
rect 48214 19214 48215 19246
rect 49912 19246 49988 19252
rect 48214 19182 48220 19214
rect 48144 18838 48220 19182
rect 47534 18774 47535 18806
rect 47469 18773 47535 18774
rect 48144 18774 48150 18838
rect 48214 18774 48220 18838
rect 49912 19182 49918 19246
rect 49982 19182 49988 19246
rect 49912 18838 49988 19182
rect 49912 18806 49918 18838
rect 48144 18768 48220 18774
rect 49917 18774 49918 18806
rect 49982 18806 49988 18838
rect 51272 19246 51348 19252
rect 51272 19182 51278 19246
rect 51342 19182 51348 19246
rect 51957 19246 52023 19247
rect 51957 19214 51958 19246
rect 51272 18838 51348 19182
rect 51272 18806 51278 18838
rect 49982 18774 49983 18806
rect 49917 18773 49983 18774
rect 51277 18774 51278 18806
rect 51342 18806 51348 18838
rect 51952 19182 51958 19214
rect 52022 19214 52023 19246
rect 53181 19246 53247 19247
rect 53181 19214 53182 19246
rect 52022 19182 52028 19214
rect 51952 18838 52028 19182
rect 51342 18774 51343 18806
rect 51277 18773 51343 18774
rect 51952 18774 51958 18838
rect 52022 18774 52028 18838
rect 51952 18768 52028 18774
rect 53176 19182 53182 19214
rect 53246 19214 53247 19246
rect 53720 19246 53796 19252
rect 53246 19182 53252 19214
rect 53176 18838 53252 19182
rect 53176 18774 53182 18838
rect 53246 18774 53252 18838
rect 53720 19182 53726 19246
rect 53790 19182 53796 19246
rect 54405 19246 54471 19247
rect 54405 19214 54406 19246
rect 53720 18838 53796 19182
rect 53720 18806 53726 18838
rect 53176 18768 53252 18774
rect 53725 18774 53726 18806
rect 53790 18806 53796 18838
rect 54400 19182 54406 19214
rect 54470 19214 54471 19246
rect 54944 19246 55020 19252
rect 54470 19182 54476 19214
rect 54400 18838 54476 19182
rect 53790 18774 53791 18806
rect 53725 18773 53791 18774
rect 54400 18774 54406 18838
rect 54470 18774 54476 18838
rect 54944 19182 54950 19246
rect 55014 19182 55020 19246
rect 55629 19246 55695 19247
rect 55629 19214 55630 19246
rect 54944 18838 55020 19182
rect 54944 18806 54950 18838
rect 54400 18768 54476 18774
rect 54949 18774 54950 18806
rect 55014 18806 55020 18838
rect 55624 19182 55630 19214
rect 55694 19214 55695 19246
rect 56168 19246 56244 19252
rect 55694 19182 55700 19214
rect 55624 18838 55700 19182
rect 55014 18774 55015 18806
rect 54949 18773 55015 18774
rect 55624 18774 55630 18838
rect 55694 18774 55700 18838
rect 56168 19182 56174 19246
rect 56238 19182 56244 19246
rect 56168 18838 56244 19182
rect 56168 18806 56174 18838
rect 55624 18768 55700 18774
rect 56173 18774 56174 18806
rect 56238 18806 56244 18838
rect 57392 19246 57468 19252
rect 57392 19182 57398 19246
rect 57462 19182 57468 19246
rect 58213 19246 58279 19247
rect 58213 19214 58214 19246
rect 57392 18838 57468 19182
rect 57392 18806 57398 18838
rect 56238 18774 56239 18806
rect 56173 18773 56239 18774
rect 57397 18774 57398 18806
rect 57462 18806 57468 18838
rect 58208 19182 58214 19214
rect 58278 19214 58279 19246
rect 59437 19246 59503 19247
rect 59437 19214 59438 19246
rect 58278 19182 58284 19214
rect 58208 18838 58284 19182
rect 57462 18774 57463 18806
rect 57397 18773 57463 18774
rect 58208 18774 58214 18838
rect 58278 18774 58284 18838
rect 58208 18768 58284 18774
rect 59432 19182 59438 19214
rect 59502 19214 59503 19246
rect 59976 19246 60052 19252
rect 59502 19182 59508 19214
rect 59432 18838 59508 19182
rect 59432 18774 59438 18838
rect 59502 18774 59508 18838
rect 59976 19182 59982 19246
rect 60046 19182 60052 19246
rect 60661 19246 60727 19247
rect 60661 19214 60662 19246
rect 59976 18838 60052 19182
rect 59976 18806 59982 18838
rect 59432 18768 59508 18774
rect 59981 18774 59982 18806
rect 60046 18806 60052 18838
rect 60656 19182 60662 19214
rect 60726 19214 60727 19246
rect 60792 19246 60868 19252
rect 60726 19182 60732 19214
rect 60656 18838 60732 19182
rect 60046 18774 60047 18806
rect 59981 18773 60047 18774
rect 60656 18774 60662 18838
rect 60726 18774 60732 18838
rect 60792 19182 60798 19246
rect 60862 19182 60868 19246
rect 61885 19246 61951 19247
rect 61885 19214 61886 19246
rect 60792 18838 60868 19182
rect 60792 18806 60798 18838
rect 60656 18768 60732 18774
rect 60797 18774 60798 18806
rect 60862 18806 60868 18838
rect 61880 19182 61886 19214
rect 61950 19214 61951 19246
rect 62424 19246 62500 19252
rect 61950 19182 61956 19214
rect 61880 18838 61956 19182
rect 60862 18774 60863 18806
rect 60797 18773 60863 18774
rect 61880 18774 61886 18838
rect 61950 18774 61956 18838
rect 62424 19182 62430 19246
rect 62494 19182 62500 19246
rect 63109 19246 63175 19247
rect 63109 19214 63110 19246
rect 62424 18838 62500 19182
rect 62424 18806 62430 18838
rect 61880 18768 61956 18774
rect 62429 18774 62430 18806
rect 62494 18806 62500 18838
rect 63104 19182 63110 19214
rect 63174 19214 63175 19246
rect 64469 19246 64535 19247
rect 64469 19214 64470 19246
rect 63174 19182 63180 19214
rect 63104 18838 63180 19182
rect 62494 18774 62495 18806
rect 62429 18773 62495 18774
rect 63104 18774 63110 18838
rect 63174 18774 63180 18838
rect 63104 18768 63180 18774
rect 64464 19182 64470 19214
rect 64534 19214 64535 19246
rect 66232 19246 66308 19252
rect 64534 19182 64540 19214
rect 64464 18838 64540 19182
rect 64464 18774 64470 18838
rect 64534 18774 64540 18838
rect 66232 19182 66238 19246
rect 66302 19182 66308 19246
rect 66917 19246 66983 19247
rect 66917 19214 66918 19246
rect 66232 18838 66308 19182
rect 66232 18806 66238 18838
rect 64464 18768 64540 18774
rect 66237 18774 66238 18806
rect 66302 18806 66308 18838
rect 66912 19182 66918 19214
rect 66982 19214 66983 19246
rect 67456 19246 67532 19252
rect 66982 19182 66988 19214
rect 66912 18838 66988 19182
rect 66302 18774 66303 18806
rect 66237 18773 66303 18774
rect 66912 18774 66918 18838
rect 66982 18774 66988 18838
rect 67456 19182 67462 19246
rect 67526 19182 67532 19246
rect 67456 18838 67532 19182
rect 67456 18806 67462 18838
rect 66912 18768 66988 18774
rect 67461 18774 67462 18806
rect 67526 18806 67532 18838
rect 68680 19246 68756 19252
rect 68680 19182 68686 19246
rect 68750 19182 68756 19246
rect 69365 19246 69431 19247
rect 69365 19214 69366 19246
rect 68680 18838 68756 19182
rect 68680 18806 68686 18838
rect 67526 18774 67527 18806
rect 67461 18773 67527 18774
rect 68685 18774 68686 18806
rect 68750 18806 68756 18838
rect 69360 19182 69366 19214
rect 69430 19214 69431 19246
rect 70997 19246 71063 19247
rect 70997 19214 70998 19246
rect 69430 19182 69436 19214
rect 69360 18838 69436 19182
rect 68750 18774 68751 18806
rect 68685 18773 68751 18774
rect 69360 18774 69366 18838
rect 69430 18774 69436 18838
rect 69360 18768 69436 18774
rect 70992 19182 70998 19214
rect 71062 19214 71063 19246
rect 71949 19246 72015 19247
rect 71949 19214 71950 19246
rect 71062 19182 71068 19214
rect 70992 18838 71068 19182
rect 70992 18774 70998 18838
rect 71062 18774 71068 18838
rect 70992 18768 71068 18774
rect 71944 19182 71950 19214
rect 72014 19214 72015 19246
rect 72352 19246 72428 19252
rect 72014 19182 72020 19214
rect 71944 18838 72020 19182
rect 71944 18774 71950 18838
rect 72014 18774 72020 18838
rect 72352 19182 72358 19246
rect 72422 19182 72428 19246
rect 73173 19246 73239 19247
rect 73173 19214 73174 19246
rect 72352 18838 72428 19182
rect 72352 18806 72358 18838
rect 71944 18768 72020 18774
rect 72357 18774 72358 18806
rect 72422 18806 72428 18838
rect 73168 19182 73174 19214
rect 73238 19214 73239 19246
rect 74936 19246 75012 19252
rect 73238 19182 73244 19214
rect 73168 18838 73244 19182
rect 72422 18774 72423 18806
rect 72357 18773 72423 18774
rect 73168 18774 73174 18838
rect 73238 18774 73244 18838
rect 74936 19182 74942 19246
rect 75006 19182 75012 19246
rect 75621 19246 75687 19247
rect 75621 19214 75622 19246
rect 74936 18838 75012 19182
rect 74936 18806 74942 18838
rect 73168 18768 73244 18774
rect 74941 18774 74942 18806
rect 75006 18806 75012 18838
rect 75616 19182 75622 19214
rect 75686 19214 75687 19246
rect 76160 19246 76236 19252
rect 75686 19182 75692 19214
rect 75616 18838 75692 19182
rect 75006 18774 75007 18806
rect 74941 18773 75007 18774
rect 75616 18774 75622 18838
rect 75686 18774 75692 18838
rect 76160 19182 76166 19246
rect 76230 19182 76236 19246
rect 76160 18838 76236 19182
rect 76160 18806 76166 18838
rect 75616 18768 75692 18774
rect 76165 18774 76166 18806
rect 76230 18806 76236 18838
rect 77384 19246 77460 19252
rect 77384 19182 77390 19246
rect 77454 19182 77460 19246
rect 78069 19246 78135 19247
rect 78069 19214 78070 19246
rect 77384 18838 77460 19182
rect 77384 18806 77390 18838
rect 76230 18774 76231 18806
rect 76165 18773 76231 18774
rect 77389 18774 77390 18806
rect 77454 18806 77460 18838
rect 78064 19182 78070 19214
rect 78134 19214 78135 19246
rect 79701 19246 79767 19247
rect 79701 19214 79702 19246
rect 78134 19182 78140 19214
rect 78064 18838 78140 19182
rect 77454 18774 77455 18806
rect 77389 18773 77455 18774
rect 78064 18774 78070 18838
rect 78134 18774 78140 18838
rect 78064 18768 78140 18774
rect 79696 19182 79702 19214
rect 79766 19214 79767 19246
rect 80653 19246 80719 19247
rect 80653 19214 80654 19246
rect 79766 19182 79772 19214
rect 79696 18838 79772 19182
rect 79696 18774 79702 18838
rect 79766 18774 79772 18838
rect 79696 18768 79772 18774
rect 80648 19182 80654 19214
rect 80718 19214 80719 19246
rect 81192 19246 81268 19252
rect 80718 19182 80724 19214
rect 80648 18838 80724 19182
rect 80648 18774 80654 18838
rect 80718 18774 80724 18838
rect 81192 19182 81198 19246
rect 81262 19182 81268 19246
rect 81877 19246 81943 19247
rect 81877 19214 81878 19246
rect 81192 18838 81268 19182
rect 81192 18806 81198 18838
rect 80648 18768 80724 18774
rect 81197 18774 81198 18806
rect 81262 18806 81268 18838
rect 81872 19182 81878 19214
rect 81942 19214 81943 19246
rect 83640 19246 83716 19252
rect 81942 19182 81948 19214
rect 81872 18838 81948 19182
rect 81262 18774 81263 18806
rect 81197 18773 81263 18774
rect 81872 18774 81878 18838
rect 81942 18774 81948 18838
rect 83640 19182 83646 19246
rect 83710 19182 83716 19246
rect 84325 19246 84391 19247
rect 84325 19214 84326 19246
rect 83640 18838 83716 19182
rect 83640 18806 83646 18838
rect 81872 18768 81948 18774
rect 83645 18774 83646 18806
rect 83710 18806 83716 18838
rect 84320 19182 84326 19214
rect 84390 19214 84391 19246
rect 84864 19246 84940 19252
rect 84390 19182 84396 19214
rect 84320 18838 84396 19182
rect 83710 18774 83711 18806
rect 83645 18773 83711 18774
rect 84320 18774 84326 18838
rect 84390 18774 84396 18838
rect 84864 19182 84870 19246
rect 84934 19182 84940 19246
rect 84864 18838 84940 19182
rect 84864 18806 84870 18838
rect 84320 18768 84396 18774
rect 84869 18774 84870 18806
rect 84934 18806 84940 18838
rect 86088 19246 86164 19252
rect 86088 19182 86094 19246
rect 86158 19182 86164 19246
rect 86909 19246 86975 19247
rect 86909 19214 86910 19246
rect 86088 18838 86164 19182
rect 86088 18806 86094 18838
rect 84934 18774 84935 18806
rect 84869 18773 84935 18774
rect 86093 18774 86094 18806
rect 86158 18806 86164 18838
rect 86904 19182 86910 19214
rect 86974 19214 86975 19246
rect 87312 19246 87388 19252
rect 86974 19182 86980 19214
rect 86904 18838 86980 19182
rect 86158 18774 86159 18806
rect 86093 18773 86159 18774
rect 86904 18774 86910 18838
rect 86974 18774 86980 18838
rect 87312 19182 87318 19246
rect 87382 19182 87388 19246
rect 88133 19246 88199 19247
rect 88133 19214 88134 19246
rect 87312 18838 87388 19182
rect 87312 18806 87318 18838
rect 86904 18768 86980 18774
rect 87317 18774 87318 18806
rect 87382 18806 87388 18838
rect 88128 19182 88134 19214
rect 88198 19214 88199 19246
rect 88264 19246 88340 19252
rect 88198 19182 88204 19214
rect 88128 18838 88204 19182
rect 87382 18774 87383 18806
rect 87317 18773 87383 18774
rect 88128 18774 88134 18838
rect 88198 18774 88204 18838
rect 88264 19182 88270 19246
rect 88334 19182 88340 19246
rect 89357 19246 89423 19247
rect 89357 19214 89358 19246
rect 88264 18838 88340 19182
rect 88264 18806 88270 18838
rect 88128 18768 88204 18774
rect 88269 18774 88270 18806
rect 88334 18806 88340 18838
rect 89352 19182 89358 19214
rect 89422 19214 89423 19246
rect 89896 19246 89972 19252
rect 89422 19182 89428 19214
rect 89352 18838 89428 19182
rect 88334 18774 88335 18806
rect 88269 18773 88335 18774
rect 89352 18774 89358 18838
rect 89422 18774 89428 18838
rect 89896 19182 89902 19246
rect 89966 19182 89972 19246
rect 90717 19246 90783 19247
rect 90717 19214 90718 19246
rect 89896 18838 89972 19182
rect 89896 18806 89902 18838
rect 89352 18768 89428 18774
rect 89901 18774 89902 18806
rect 89966 18806 89972 18838
rect 90712 19182 90718 19214
rect 90782 19214 90783 19246
rect 91805 19246 91871 19247
rect 91805 19214 91806 19246
rect 90782 19182 90788 19214
rect 90712 18838 90788 19182
rect 89966 18774 89967 18806
rect 89901 18773 89967 18774
rect 90712 18774 90718 18838
rect 90782 18774 90788 18838
rect 90712 18768 90788 18774
rect 91800 19182 91806 19214
rect 91870 19214 91871 19246
rect 92344 19246 92420 19252
rect 91870 19182 91876 19214
rect 91800 18838 91876 19182
rect 91800 18774 91806 18838
rect 91870 18774 91876 18838
rect 92344 19182 92350 19246
rect 92414 19182 92420 19246
rect 93437 19246 93503 19247
rect 93437 19214 93438 19246
rect 92344 18838 92420 19182
rect 92344 18806 92350 18838
rect 91800 18768 91876 18774
rect 92349 18774 92350 18806
rect 92414 18806 92420 18838
rect 93432 19182 93438 19214
rect 93502 19214 93503 19246
rect 93502 19182 93508 19214
rect 93432 18838 93508 19182
rect 92414 18774 92415 18806
rect 92349 18773 92415 18774
rect 93432 18774 93438 18838
rect 93502 18774 93508 18838
rect 94520 18838 94596 19318
rect 95613 19246 95679 19247
rect 95613 19214 95614 19246
rect 94520 18806 94526 18838
rect 93432 18768 93508 18774
rect 94525 18774 94526 18806
rect 94590 18806 94596 18838
rect 95608 19182 95614 19214
rect 95678 19214 95679 19246
rect 96152 19246 96228 19252
rect 95678 19182 95684 19214
rect 95608 18838 95684 19182
rect 94590 18774 94591 18806
rect 94525 18773 94591 18774
rect 95608 18774 95614 18838
rect 95678 18774 95684 18838
rect 96152 19182 96158 19246
rect 96222 19182 96228 19246
rect 96837 19246 96903 19247
rect 96837 19214 96838 19246
rect 96152 18838 96228 19182
rect 96152 18806 96158 18838
rect 95608 18768 95684 18774
rect 96157 18774 96158 18806
rect 96222 18806 96228 18838
rect 96832 19182 96838 19214
rect 96902 19214 96903 19246
rect 98197 19246 98263 19247
rect 98197 19214 98198 19246
rect 96902 19182 96908 19214
rect 96832 18838 96908 19182
rect 96222 18774 96223 18806
rect 96157 18773 96223 18774
rect 96832 18774 96838 18838
rect 96902 18774 96908 18838
rect 96832 18768 96908 18774
rect 98192 19182 98198 19214
rect 98262 19214 98263 19246
rect 98600 19246 98676 19252
rect 98262 19182 98268 19214
rect 98192 18838 98268 19182
rect 98192 18774 98198 18838
rect 98262 18774 98268 18838
rect 98600 19182 98606 19246
rect 98670 19182 98676 19246
rect 98600 18838 98676 19182
rect 98600 18806 98606 18838
rect 98192 18768 98268 18774
rect 98605 18774 98606 18806
rect 98670 18806 98676 18838
rect 99824 19246 99900 19252
rect 99824 19182 99830 19246
rect 99894 19182 99900 19246
rect 99824 18838 99900 19182
rect 99824 18806 99830 18838
rect 98670 18774 98671 18806
rect 98605 18773 98671 18774
rect 99829 18774 99830 18806
rect 99894 18806 99900 18838
rect 101184 19246 101260 19252
rect 101184 19182 101190 19246
rect 101254 19182 101260 19246
rect 101869 19246 101935 19247
rect 101869 19214 101870 19246
rect 101184 18838 101260 19182
rect 101184 18806 101190 18838
rect 99894 18774 99895 18806
rect 99829 18773 99895 18774
rect 101189 18774 101190 18806
rect 101254 18806 101260 18838
rect 101864 19182 101870 19214
rect 101934 19214 101935 19246
rect 102408 19246 102484 19252
rect 101934 19182 101940 19214
rect 101864 18838 101940 19182
rect 101254 18774 101255 18806
rect 101189 18773 101255 18774
rect 101864 18774 101870 18838
rect 101934 18774 101940 18838
rect 102408 19182 102414 19246
rect 102478 19182 102484 19246
rect 103093 19246 103159 19247
rect 103093 19214 103094 19246
rect 102408 18838 102484 19182
rect 102408 18806 102414 18838
rect 101864 18768 101940 18774
rect 102413 18774 102414 18806
rect 102478 18806 102484 18838
rect 103088 19182 103094 19214
rect 103158 19214 103159 19246
rect 104317 19246 104383 19247
rect 104317 19214 104318 19246
rect 103158 19182 103164 19214
rect 103088 18838 103164 19182
rect 102478 18774 102479 18806
rect 102413 18773 102479 18774
rect 103088 18774 103094 18838
rect 103158 18774 103164 18838
rect 103088 18768 103164 18774
rect 104312 19182 104318 19214
rect 104382 19214 104383 19246
rect 104856 19246 104932 19252
rect 104382 19182 104388 19214
rect 104312 18838 104388 19182
rect 104312 18774 104318 18838
rect 104382 18774 104388 18838
rect 104856 19182 104862 19246
rect 104926 19182 104932 19246
rect 105541 19246 105607 19247
rect 105541 19214 105542 19246
rect 104856 18838 104932 19182
rect 104856 18806 104862 18838
rect 104312 18768 104388 18774
rect 104861 18774 104862 18806
rect 104926 18806 104932 18838
rect 105536 19182 105542 19214
rect 105606 19214 105607 19246
rect 105808 19246 105884 19252
rect 105606 19182 105612 19214
rect 105536 18838 105612 19182
rect 104926 18774 104927 18806
rect 104861 18773 104927 18774
rect 105536 18774 105542 18838
rect 105606 18774 105612 18838
rect 105808 19182 105814 19246
rect 105878 19182 105884 19246
rect 107173 19246 107239 19247
rect 107173 19214 107174 19246
rect 105808 18838 105884 19182
rect 105808 18806 105814 18838
rect 105536 18768 105612 18774
rect 105813 18774 105814 18806
rect 105878 18806 105884 18838
rect 107168 19182 107174 19214
rect 107238 19214 107239 19246
rect 107304 19246 107380 19252
rect 107238 19182 107244 19214
rect 107168 18838 107244 19182
rect 105878 18774 105879 18806
rect 105813 18773 105879 18774
rect 107168 18774 107174 18838
rect 107238 18774 107244 18838
rect 107304 19182 107310 19246
rect 107374 19182 107380 19246
rect 107304 18838 107380 19182
rect 107304 18806 107310 18838
rect 107168 18768 107244 18774
rect 107309 18774 107310 18806
rect 107374 18806 107380 18838
rect 108528 19246 108604 19252
rect 108528 19182 108534 19246
rect 108598 19182 108604 19246
rect 108528 18838 108604 19182
rect 108528 18806 108534 18838
rect 107374 18774 107375 18806
rect 107309 18773 107375 18774
rect 108533 18774 108534 18806
rect 108598 18806 108604 18838
rect 108598 18774 108599 18806
rect 108533 18773 108599 18774
rect 58349 18702 58415 18703
rect 58349 18670 58350 18702
rect 28968 17142 28974 17206
rect 29038 17142 29044 17206
rect 28968 17136 29044 17142
rect 58344 18638 58350 18670
rect 58414 18670 58415 18702
rect 58414 18638 58420 18670
rect 22440 15814 22446 15846
rect 22445 15782 22446 15814
rect 22510 15814 22516 15846
rect 28968 17070 29044 17076
rect 28968 17006 28974 17070
rect 29038 17006 29044 17070
rect 22510 15782 22511 15814
rect 22445 15781 22511 15782
rect 28968 15166 29044 17006
rect 31688 17070 31764 17076
rect 31688 17006 31694 17070
rect 31758 17006 31764 17070
rect 28968 15134 28974 15166
rect 28973 15102 28974 15134
rect 29038 15134 29044 15166
rect 29104 15166 29180 15172
rect 29038 15102 29039 15134
rect 28973 15101 29039 15102
rect 29104 15102 29110 15166
rect 29174 15102 29180 15166
rect 21352 14558 21358 14622
rect 21422 14558 21428 14622
rect 21352 14552 21428 14558
rect 28837 14350 28903 14351
rect 28837 14318 28838 14350
rect 28832 14286 28838 14318
rect 28902 14318 28903 14350
rect 28902 14286 28908 14318
rect 28832 13670 28908 14286
rect 28832 13606 28838 13670
rect 28902 13606 28908 13670
rect 28832 13600 28908 13606
rect 28968 13534 29044 13540
rect 28968 13470 28974 13534
rect 29038 13470 29044 13534
rect 21216 13062 21222 13126
rect 21286 13062 21292 13126
rect 28293 13126 28359 13127
rect 28293 13094 28294 13126
rect 21216 13056 21292 13062
rect 28288 13062 28294 13094
rect 28358 13094 28359 13126
rect 28358 13062 28364 13094
rect 20264 11734 20270 11766
rect 20269 11702 20270 11734
rect 20334 11734 20340 11766
rect 20334 11702 20335 11734
rect 20269 11701 20335 11702
rect 14688 10510 14694 10542
rect 14693 10478 14694 10510
rect 14758 10510 14764 10542
rect 28152 11358 28228 11364
rect 28152 11294 28158 11358
rect 28222 11294 28228 11358
rect 14758 10478 14759 10510
rect 14693 10477 14759 10478
rect 14552 9150 14558 9182
rect 14557 9118 14558 9150
rect 14622 9150 14628 9182
rect 14688 10406 14764 10412
rect 14688 10342 14694 10406
rect 14758 10342 14764 10406
rect 14622 9118 14623 9150
rect 14557 9117 14623 9118
rect 952 8710 1230 8774
rect 1294 8710 1300 8774
rect 952 7278 1300 8710
rect 14688 7686 14764 10342
rect 28152 9590 28228 11294
rect 28152 9558 28158 9590
rect 28157 9526 28158 9558
rect 28222 9558 28228 9590
rect 28222 9526 28223 9558
rect 28157 9525 28223 9526
rect 16325 9046 16391 9047
rect 16325 9014 16326 9046
rect 14688 7654 14694 7686
rect 14693 7622 14694 7654
rect 14758 7654 14764 7686
rect 16320 8982 16326 9014
rect 16390 9014 16391 9046
rect 16390 8982 16396 9014
rect 14758 7622 14759 7654
rect 14693 7621 14759 7622
rect 952 7214 1230 7278
rect 1294 7214 1300 7278
rect 952 5510 1300 7214
rect 952 5446 1230 5510
rect 1294 5446 1300 5510
rect 952 3878 1300 5446
rect 952 3814 1230 3878
rect 1294 3814 1300 3878
rect 952 1294 1300 3814
rect 16320 3878 16396 8982
rect 16320 3814 16326 3878
rect 16390 3814 16396 3878
rect 16320 3808 16396 3814
rect 20269 3742 20335 3743
rect 20269 3710 20270 3742
rect 20264 3678 20270 3710
rect 20334 3710 20335 3742
rect 20334 3678 20340 3710
rect 16053 2926 16119 2927
rect 16053 2894 16054 2926
rect 16048 2862 16054 2894
rect 16118 2894 16119 2926
rect 17141 2926 17207 2927
rect 17141 2894 17142 2926
rect 16118 2862 16124 2894
rect 2045 1702 2111 1703
rect 2045 1670 2046 1702
rect 952 1230 958 1294
rect 1022 1230 1094 1294
rect 1158 1230 1230 1294
rect 1294 1230 1300 1294
rect 952 1158 1300 1230
rect 2040 1638 2046 1670
rect 2110 1670 2111 1702
rect 3813 1702 3879 1703
rect 3813 1670 3814 1702
rect 2110 1638 2116 1670
rect 2040 1294 2116 1638
rect 2040 1230 2046 1294
rect 2110 1230 2116 1294
rect 2040 1224 2116 1230
rect 3808 1638 3814 1670
rect 3878 1670 3879 1702
rect 5581 1702 5647 1703
rect 5581 1670 5582 1702
rect 3878 1638 3884 1670
rect 3808 1294 3884 1638
rect 3808 1230 3814 1294
rect 3878 1230 3884 1294
rect 3808 1224 3884 1230
rect 5576 1638 5582 1670
rect 5646 1670 5647 1702
rect 7077 1702 7143 1703
rect 7077 1670 7078 1702
rect 5646 1638 5652 1670
rect 5576 1294 5652 1638
rect 5576 1230 5582 1294
rect 5646 1230 5652 1294
rect 5576 1224 5652 1230
rect 7072 1638 7078 1670
rect 7142 1670 7143 1702
rect 8709 1702 8775 1703
rect 8709 1670 8710 1702
rect 7142 1638 7148 1670
rect 7072 1294 7148 1638
rect 7072 1230 7078 1294
rect 7142 1230 7148 1294
rect 7072 1224 7148 1230
rect 8704 1638 8710 1670
rect 8774 1670 8775 1702
rect 10477 1702 10543 1703
rect 10477 1670 10478 1702
rect 8774 1638 8780 1670
rect 8704 1294 8780 1638
rect 8704 1230 8710 1294
rect 8774 1230 8780 1294
rect 8704 1224 8780 1230
rect 10472 1638 10478 1670
rect 10542 1670 10543 1702
rect 12109 1702 12175 1703
rect 12109 1670 12110 1702
rect 10542 1638 10548 1670
rect 10472 1294 10548 1638
rect 10472 1230 10478 1294
rect 10542 1230 10548 1294
rect 10472 1224 10548 1230
rect 12104 1638 12110 1670
rect 12174 1670 12175 1702
rect 14013 1702 14079 1703
rect 14013 1670 14014 1702
rect 12174 1638 12180 1670
rect 12104 1294 12180 1638
rect 12104 1230 12110 1294
rect 12174 1230 12180 1294
rect 12104 1224 12180 1230
rect 14008 1638 14014 1670
rect 14078 1670 14079 1702
rect 15509 1702 15575 1703
rect 15509 1670 15510 1702
rect 14078 1638 14084 1670
rect 14008 1294 14084 1638
rect 14008 1230 14014 1294
rect 14078 1230 14084 1294
rect 14008 1224 14084 1230
rect 15504 1638 15510 1670
rect 15574 1670 15575 1702
rect 15574 1638 15580 1670
rect 15504 1294 15580 1638
rect 15504 1230 15510 1294
rect 15574 1230 15580 1294
rect 15504 1224 15580 1230
rect 952 1094 958 1158
rect 1022 1094 1094 1158
rect 1158 1094 1230 1158
rect 1294 1094 1300 1158
rect 952 1022 1300 1094
rect 952 958 958 1022
rect 1022 958 1094 1022
rect 1158 958 1230 1022
rect 1294 958 1300 1022
rect 952 952 1300 958
rect 272 550 278 614
rect 342 550 414 614
rect 478 550 550 614
rect 614 550 620 614
rect 272 478 620 550
rect 272 414 278 478
rect 342 414 414 478
rect 478 414 550 478
rect 614 414 620 478
rect 272 342 620 414
rect 272 278 278 342
rect 342 278 414 342
rect 478 278 550 342
rect 614 278 620 342
rect 272 272 620 278
rect 16048 0 16124 2862
rect 17136 2862 17142 2894
rect 17206 2894 17207 2926
rect 18229 2926 18295 2927
rect 18229 2894 18230 2926
rect 17206 2862 17212 2894
rect 17136 0 17212 2862
rect 18224 2862 18230 2894
rect 18294 2894 18295 2926
rect 19589 2926 19655 2927
rect 19589 2894 19590 2926
rect 18294 2862 18300 2894
rect 17413 1702 17479 1703
rect 17413 1670 17414 1702
rect 17408 1638 17414 1670
rect 17478 1670 17479 1702
rect 17478 1638 17484 1670
rect 17408 1294 17484 1638
rect 17408 1230 17414 1294
rect 17478 1230 17484 1294
rect 17408 1224 17484 1230
rect 18224 0 18300 2862
rect 19584 2862 19590 2894
rect 19654 2894 19655 2926
rect 19654 2862 19660 2894
rect 19045 1702 19111 1703
rect 19045 1670 19046 1702
rect 19040 1638 19046 1670
rect 19110 1670 19111 1702
rect 19110 1638 19116 1670
rect 19040 1294 19116 1638
rect 19040 1230 19046 1294
rect 19110 1230 19116 1294
rect 19040 1224 19116 1230
rect 19584 0 19660 2862
rect 20264 1838 20340 3678
rect 20541 2926 20607 2927
rect 20541 2894 20542 2926
rect 20264 1774 20270 1838
rect 20334 1774 20340 1838
rect 20264 1768 20340 1774
rect 20536 2862 20542 2894
rect 20606 2894 20607 2926
rect 21765 2926 21831 2927
rect 21765 2894 21766 2926
rect 20606 2862 20612 2894
rect 20536 0 20612 2862
rect 21760 2862 21766 2894
rect 21830 2894 21831 2926
rect 23125 2926 23191 2927
rect 23125 2894 23126 2926
rect 21830 2862 21836 2894
rect 20813 1702 20879 1703
rect 20813 1670 20814 1702
rect 20808 1638 20814 1670
rect 20878 1670 20879 1702
rect 20878 1638 20884 1670
rect 20808 1294 20884 1638
rect 20808 1230 20814 1294
rect 20878 1230 20884 1294
rect 20808 1224 20884 1230
rect 21760 0 21836 2862
rect 23120 2862 23126 2894
rect 23190 2894 23191 2926
rect 24213 2926 24279 2927
rect 24213 2894 24214 2926
rect 23190 2862 23196 2894
rect 22173 1702 22239 1703
rect 22173 1670 22174 1702
rect 22168 1638 22174 1670
rect 22238 1670 22239 1702
rect 22238 1638 22244 1670
rect 22168 1294 22244 1638
rect 22168 1230 22174 1294
rect 22238 1230 22244 1294
rect 22168 1224 22244 1230
rect 23120 0 23196 2862
rect 24208 2862 24214 2894
rect 24278 2894 24279 2926
rect 25437 2926 25503 2927
rect 25437 2894 25438 2926
rect 24278 2862 24284 2894
rect 23941 1702 24007 1703
rect 23941 1670 23942 1702
rect 23936 1638 23942 1670
rect 24006 1670 24007 1702
rect 24006 1638 24012 1670
rect 23936 1294 24012 1638
rect 23936 1230 23942 1294
rect 24006 1230 24012 1294
rect 23936 1224 24012 1230
rect 24208 0 24284 2862
rect 25432 2862 25438 2894
rect 25502 2894 25503 2926
rect 26525 2926 26591 2927
rect 26525 2894 26526 2926
rect 25502 2862 25508 2894
rect 25432 0 25508 2862
rect 26520 2862 26526 2894
rect 26590 2894 26591 2926
rect 27613 2926 27679 2927
rect 27613 2894 27614 2926
rect 26590 2862 26596 2894
rect 25709 1702 25775 1703
rect 25709 1670 25710 1702
rect 25704 1638 25710 1670
rect 25774 1670 25775 1702
rect 25774 1638 25780 1670
rect 25704 1294 25780 1638
rect 25704 1230 25710 1294
rect 25774 1230 25780 1294
rect 25704 1224 25780 1230
rect 26520 0 26596 2862
rect 27608 2862 27614 2894
rect 27678 2894 27679 2926
rect 27678 2862 27684 2894
rect 27341 1702 27407 1703
rect 27341 1670 27342 1702
rect 27336 1638 27342 1670
rect 27406 1670 27407 1702
rect 27406 1638 27412 1670
rect 27336 1294 27412 1638
rect 27336 1230 27342 1294
rect 27406 1230 27412 1294
rect 27336 1224 27412 1230
rect 27608 0 27684 2862
rect 28288 0 28364 13062
rect 28837 12310 28903 12311
rect 28837 12278 28838 12310
rect 28832 12246 28838 12278
rect 28902 12278 28903 12310
rect 28902 12246 28908 12278
rect 28701 11902 28767 11903
rect 28701 11870 28702 11902
rect 28696 11838 28702 11870
rect 28766 11870 28767 11902
rect 28766 11838 28772 11870
rect 28560 11086 28636 11092
rect 28560 11022 28566 11086
rect 28630 11022 28636 11086
rect 28560 10678 28636 11022
rect 28696 11086 28772 11838
rect 28832 11766 28908 12246
rect 28968 12038 29044 13470
rect 29104 13262 29180 15102
rect 31552 15166 31628 15172
rect 31552 15102 31558 15166
rect 31622 15102 31628 15166
rect 31688 15166 31764 17006
rect 31688 15134 31694 15166
rect 31421 14350 31487 14351
rect 31421 14318 31422 14350
rect 31416 14286 31422 14318
rect 31486 14318 31487 14350
rect 31486 14286 31492 14318
rect 31416 13670 31492 14286
rect 31416 13606 31422 13670
rect 31486 13606 31492 13670
rect 31416 13600 31492 13606
rect 29104 13230 29110 13262
rect 29109 13198 29110 13230
rect 29174 13230 29180 13262
rect 31280 13534 31356 13540
rect 31280 13470 31286 13534
rect 31350 13470 31356 13534
rect 29174 13198 29175 13230
rect 29109 13197 29175 13198
rect 29104 13126 29180 13132
rect 29104 13062 29110 13126
rect 29174 13062 29180 13126
rect 30741 13126 30807 13127
rect 30741 13094 30742 13126
rect 29104 12582 29180 13062
rect 29104 12550 29110 12582
rect 29109 12518 29110 12550
rect 29174 12550 29180 12582
rect 30736 13062 30742 13094
rect 30806 13094 30807 13126
rect 30806 13062 30812 13094
rect 29174 12518 29175 12550
rect 29109 12517 29175 12518
rect 28968 12006 28974 12038
rect 28973 11974 28974 12006
rect 29038 12006 29044 12038
rect 29038 11974 29039 12006
rect 28973 11973 29039 11974
rect 28832 11702 28838 11766
rect 28902 11702 28908 11766
rect 28832 11696 28908 11702
rect 28696 11022 28702 11086
rect 28766 11022 28772 11086
rect 28696 11016 28772 11022
rect 28560 10646 28566 10678
rect 28565 10614 28566 10646
rect 28630 10646 28636 10678
rect 28630 10614 28631 10646
rect 28565 10613 28631 10614
rect 28701 2926 28767 2927
rect 28701 2894 28702 2926
rect 28696 2862 28702 2894
rect 28766 2894 28767 2926
rect 30061 2926 30127 2927
rect 30061 2894 30062 2926
rect 28766 2862 28772 2894
rect 28696 0 28772 2862
rect 30056 2862 30062 2894
rect 30126 2894 30127 2926
rect 30126 2862 30132 2894
rect 28973 1702 29039 1703
rect 28973 1670 28974 1702
rect 28968 1638 28974 1670
rect 29038 1670 29039 1702
rect 29038 1638 29044 1670
rect 28968 1294 29044 1638
rect 28968 1230 28974 1294
rect 29038 1230 29044 1294
rect 28968 1224 29044 1230
rect 30056 0 30132 2862
rect 30469 1702 30535 1703
rect 30469 1670 30470 1702
rect 30464 1638 30470 1670
rect 30534 1670 30535 1702
rect 30534 1638 30540 1670
rect 30464 1294 30540 1638
rect 30464 1230 30470 1294
rect 30534 1230 30540 1294
rect 30464 1224 30540 1230
rect 30736 0 30812 13062
rect 31280 12038 31356 13470
rect 31552 13262 31628 15102
rect 31693 15102 31694 15134
rect 31758 15134 31764 15166
rect 34000 17070 34076 17076
rect 34000 17006 34006 17070
rect 34070 17006 34076 17070
rect 34000 15166 34076 17006
rect 36448 17070 36524 17076
rect 36448 17006 36454 17070
rect 36518 17006 36524 17070
rect 34000 15134 34006 15166
rect 31758 15102 31759 15134
rect 31693 15101 31759 15102
rect 34005 15102 34006 15134
rect 34070 15134 34076 15166
rect 34136 15166 34212 15172
rect 34070 15102 34071 15134
rect 34005 15101 34071 15102
rect 34136 15102 34142 15166
rect 34206 15102 34212 15166
rect 36448 15166 36524 17006
rect 39168 17070 39244 17076
rect 39168 17006 39174 17070
rect 39238 17006 39244 17070
rect 36448 15134 36454 15166
rect 33592 14350 33668 14356
rect 33592 14286 33598 14350
rect 33662 14286 33668 14350
rect 33869 14350 33935 14351
rect 33869 14318 33870 14350
rect 33592 13670 33668 14286
rect 33592 13638 33598 13670
rect 33597 13606 33598 13638
rect 33662 13638 33668 13670
rect 33864 14286 33870 14318
rect 33934 14318 33935 14350
rect 33934 14286 33940 14318
rect 33864 13670 33940 14286
rect 33662 13606 33663 13638
rect 33597 13605 33663 13606
rect 33864 13606 33870 13670
rect 33934 13606 33940 13670
rect 33864 13600 33940 13606
rect 31552 13230 31558 13262
rect 31557 13198 31558 13230
rect 31622 13230 31628 13262
rect 34000 13534 34076 13540
rect 34000 13470 34006 13534
rect 34070 13470 34076 13534
rect 31622 13198 31623 13230
rect 31557 13197 31623 13198
rect 31416 13126 31492 13132
rect 31416 13062 31422 13126
rect 31486 13062 31492 13126
rect 33597 13126 33663 13127
rect 33597 13094 33598 13126
rect 31416 12582 31492 13062
rect 31416 12550 31422 12582
rect 31421 12518 31422 12550
rect 31486 12550 31492 12582
rect 33592 13062 33598 13094
rect 33662 13094 33663 13126
rect 33864 13126 33940 13132
rect 33662 13062 33668 13094
rect 31486 12518 31487 12550
rect 31421 12517 31487 12518
rect 31421 12310 31487 12311
rect 31421 12278 31422 12310
rect 31280 12006 31286 12038
rect 31285 11974 31286 12006
rect 31350 12006 31356 12038
rect 31416 12246 31422 12278
rect 31486 12278 31487 12310
rect 33461 12310 33527 12311
rect 33461 12278 33462 12310
rect 31486 12246 31492 12278
rect 31350 11974 31351 12006
rect 31285 11973 31351 11974
rect 31149 11902 31215 11903
rect 31149 11870 31150 11902
rect 31144 11838 31150 11870
rect 31214 11870 31215 11902
rect 31214 11838 31220 11870
rect 31144 11086 31220 11838
rect 31416 11766 31492 12246
rect 31416 11702 31422 11766
rect 31486 11702 31492 11766
rect 31416 11696 31492 11702
rect 33456 12246 33462 12278
rect 33526 12278 33527 12310
rect 33526 12246 33532 12278
rect 33456 11766 33532 12246
rect 33456 11702 33462 11766
rect 33526 11702 33532 11766
rect 33456 11696 33532 11702
rect 31144 11022 31150 11086
rect 31214 11022 31220 11086
rect 31144 11016 31220 11022
rect 31285 2926 31351 2927
rect 31285 2894 31286 2926
rect 31280 2862 31286 2894
rect 31350 2894 31351 2926
rect 32373 2926 32439 2927
rect 32373 2894 32374 2926
rect 31350 2862 31356 2894
rect 31280 0 31356 2862
rect 32368 2862 32374 2894
rect 32438 2894 32439 2926
rect 33461 2926 33527 2927
rect 33461 2894 33462 2926
rect 32438 2862 32444 2894
rect 32101 1702 32167 1703
rect 32101 1670 32102 1702
rect 32096 1638 32102 1670
rect 32166 1670 32167 1702
rect 32166 1638 32172 1670
rect 32096 1294 32172 1638
rect 32096 1230 32102 1294
rect 32166 1230 32172 1294
rect 32096 1224 32172 1230
rect 32368 0 32444 2862
rect 33456 2862 33462 2894
rect 33526 2894 33527 2926
rect 33526 2862 33532 2894
rect 33456 0 33532 2862
rect 33592 0 33668 13062
rect 33864 13062 33870 13126
rect 33934 13062 33940 13126
rect 33864 12582 33940 13062
rect 33864 12550 33870 12582
rect 33869 12518 33870 12550
rect 33934 12550 33940 12582
rect 33934 12518 33935 12550
rect 33869 12517 33935 12518
rect 34000 12038 34076 13470
rect 34136 13262 34212 15102
rect 36453 15102 36454 15134
rect 36518 15134 36524 15166
rect 36584 15166 36660 15172
rect 36518 15102 36519 15134
rect 36453 15101 36519 15102
rect 36584 15102 36590 15166
rect 36654 15102 36660 15166
rect 36453 14350 36519 14351
rect 36453 14318 36454 14350
rect 36448 14286 36454 14318
rect 36518 14318 36519 14350
rect 36518 14286 36524 14318
rect 36448 13670 36524 14286
rect 36448 13606 36454 13670
rect 36518 13606 36524 13670
rect 36448 13600 36524 13606
rect 34136 13230 34142 13262
rect 34141 13198 34142 13230
rect 34206 13230 34212 13262
rect 36448 13534 36524 13540
rect 36448 13470 36454 13534
rect 36518 13470 36524 13534
rect 34206 13198 34207 13230
rect 34141 13197 34207 13198
rect 36045 13126 36111 13127
rect 36045 13094 36046 13126
rect 34000 12006 34006 12038
rect 34005 11974 34006 12006
rect 34070 12006 34076 12038
rect 36040 13062 36046 13094
rect 36110 13094 36111 13126
rect 36110 13062 36116 13094
rect 34070 11974 34071 12006
rect 34005 11973 34071 11974
rect 33869 11902 33935 11903
rect 33869 11870 33870 11902
rect 33864 11838 33870 11870
rect 33934 11870 33935 11902
rect 33934 11838 33940 11870
rect 33864 11086 33940 11838
rect 33864 11022 33870 11086
rect 33934 11022 33940 11086
rect 33864 11016 33940 11022
rect 34549 2926 34615 2927
rect 34549 2894 34550 2926
rect 34544 2862 34550 2894
rect 34614 2894 34615 2926
rect 35909 2926 35975 2927
rect 35909 2894 35910 2926
rect 34614 2862 34620 2894
rect 34005 1702 34071 1703
rect 34005 1670 34006 1702
rect 34000 1638 34006 1670
rect 34070 1670 34071 1702
rect 34070 1638 34076 1670
rect 34000 1294 34076 1638
rect 34000 1230 34006 1294
rect 34070 1230 34076 1294
rect 34000 1224 34076 1230
rect 34544 0 34620 2862
rect 35904 2862 35910 2894
rect 35974 2894 35975 2926
rect 35974 2862 35980 2894
rect 35773 1702 35839 1703
rect 35773 1670 35774 1702
rect 35768 1638 35774 1670
rect 35838 1670 35839 1702
rect 35838 1638 35844 1670
rect 35768 1294 35844 1638
rect 35768 1230 35774 1294
rect 35838 1230 35844 1294
rect 35768 1224 35844 1230
rect 35904 0 35980 2862
rect 36040 0 36116 13062
rect 36181 12310 36247 12311
rect 36181 12278 36182 12310
rect 36176 12246 36182 12278
rect 36246 12278 36247 12310
rect 36246 12246 36252 12278
rect 36176 11766 36252 12246
rect 36448 12038 36524 13470
rect 36584 13262 36660 15102
rect 39032 15166 39108 15172
rect 39032 15102 39038 15166
rect 39102 15102 39108 15166
rect 39168 15166 39244 17006
rect 41616 17070 41692 17076
rect 41616 17006 41622 17070
rect 41686 17006 41692 17070
rect 39168 15134 39174 15166
rect 38901 14350 38967 14351
rect 38901 14318 38902 14350
rect 38896 14286 38902 14318
rect 38966 14318 38967 14350
rect 38966 14286 38972 14318
rect 38896 13670 38972 14286
rect 38896 13606 38902 13670
rect 38966 13606 38972 13670
rect 38896 13600 38972 13606
rect 36584 13230 36590 13262
rect 36589 13198 36590 13230
rect 36654 13230 36660 13262
rect 38896 13534 38972 13540
rect 38896 13470 38902 13534
rect 38966 13470 38972 13534
rect 36654 13198 36655 13230
rect 36589 13197 36655 13198
rect 36584 13126 36660 13132
rect 36584 13062 36590 13126
rect 36654 13062 36660 13126
rect 38493 13126 38559 13127
rect 38493 13094 38494 13126
rect 36584 12582 36660 13062
rect 36584 12550 36590 12582
rect 36589 12518 36590 12550
rect 36654 12550 36660 12582
rect 38488 13062 38494 13094
rect 38558 13094 38559 13126
rect 38558 13062 38564 13094
rect 36654 12518 36655 12550
rect 36589 12517 36655 12518
rect 36448 12006 36454 12038
rect 36453 11974 36454 12006
rect 36518 12006 36524 12038
rect 36518 11974 36519 12006
rect 36453 11973 36519 11974
rect 36317 11902 36383 11903
rect 36317 11870 36318 11902
rect 36176 11702 36182 11766
rect 36246 11702 36252 11766
rect 36176 11696 36252 11702
rect 36312 11838 36318 11870
rect 36382 11870 36383 11902
rect 36382 11838 36388 11870
rect 36312 11086 36388 11838
rect 36312 11022 36318 11086
rect 36382 11022 36388 11086
rect 36312 11016 36388 11022
rect 36997 2926 37063 2927
rect 36997 2894 36998 2926
rect 36992 2862 36998 2894
rect 37062 2894 37063 2926
rect 38085 2926 38151 2927
rect 38085 2894 38086 2926
rect 37062 2862 37068 2894
rect 36992 0 37068 2862
rect 38080 2862 38086 2894
rect 38150 2894 38151 2926
rect 38150 2862 38156 2894
rect 37405 1702 37471 1703
rect 37405 1670 37406 1702
rect 37400 1638 37406 1670
rect 37470 1670 37471 1702
rect 37470 1638 37476 1670
rect 37400 1294 37476 1638
rect 37400 1230 37406 1294
rect 37470 1230 37476 1294
rect 37400 1224 37476 1230
rect 38080 0 38156 2862
rect 38488 0 38564 13062
rect 38629 12310 38695 12311
rect 38629 12278 38630 12310
rect 38624 12246 38630 12278
rect 38694 12278 38695 12310
rect 38694 12246 38700 12278
rect 38624 11766 38700 12246
rect 38896 12038 38972 13470
rect 39032 13262 39108 15102
rect 39173 15102 39174 15134
rect 39238 15134 39244 15166
rect 41480 15166 41556 15172
rect 39238 15102 39239 15134
rect 39173 15101 39239 15102
rect 41480 15102 41486 15166
rect 41550 15102 41556 15166
rect 41616 15166 41692 17006
rect 41616 15134 41622 15166
rect 41077 14350 41143 14351
rect 41077 14318 41078 14350
rect 41072 14286 41078 14318
rect 41142 14318 41143 14350
rect 41213 14350 41279 14351
rect 41213 14318 41214 14350
rect 41142 14286 41148 14318
rect 41072 13670 41148 14286
rect 41072 13606 41078 13670
rect 41142 13606 41148 13670
rect 41072 13600 41148 13606
rect 41208 14286 41214 14318
rect 41278 14318 41279 14350
rect 41278 14286 41284 14318
rect 41208 13670 41284 14286
rect 41208 13606 41214 13670
rect 41278 13606 41284 13670
rect 41208 13600 41284 13606
rect 39032 13230 39038 13262
rect 39037 13198 39038 13230
rect 39102 13230 39108 13262
rect 41344 13534 41420 13540
rect 41344 13470 41350 13534
rect 41414 13470 41420 13534
rect 39102 13198 39103 13230
rect 39037 13197 39103 13198
rect 39032 13126 39108 13132
rect 39032 13062 39038 13126
rect 39102 13062 39108 13126
rect 41077 13126 41143 13127
rect 41077 13094 41078 13126
rect 39032 12582 39108 13062
rect 39032 12550 39038 12582
rect 39037 12518 39038 12550
rect 39102 12550 39108 12582
rect 41072 13062 41078 13094
rect 41142 13094 41143 13126
rect 41142 13062 41148 13094
rect 39102 12518 39103 12550
rect 39037 12517 39103 12518
rect 38896 12006 38902 12038
rect 38901 11974 38902 12006
rect 38966 12006 38972 12038
rect 38966 11974 38967 12006
rect 38901 11973 38967 11974
rect 38765 11902 38831 11903
rect 38765 11870 38766 11902
rect 38624 11702 38630 11766
rect 38694 11702 38700 11766
rect 38624 11696 38700 11702
rect 38760 11838 38766 11870
rect 38830 11870 38831 11902
rect 38830 11838 38836 11870
rect 38760 11086 38836 11838
rect 38760 11022 38766 11086
rect 38830 11022 38836 11086
rect 38760 11016 38836 11022
rect 39445 2926 39511 2927
rect 39445 2894 39446 2926
rect 39440 2862 39446 2894
rect 39510 2894 39511 2926
rect 40669 2926 40735 2927
rect 40669 2894 40670 2926
rect 39510 2862 39516 2894
rect 39173 1702 39239 1703
rect 39173 1670 39174 1702
rect 39168 1638 39174 1670
rect 39238 1670 39239 1702
rect 39238 1638 39244 1670
rect 39168 1294 39244 1638
rect 39168 1230 39174 1294
rect 39238 1230 39244 1294
rect 39168 1224 39244 1230
rect 39440 0 39516 2862
rect 40664 2862 40670 2894
rect 40734 2894 40735 2926
rect 40734 2862 40740 2894
rect 39717 2382 39783 2383
rect 39717 2350 39718 2382
rect 39712 2318 39718 2350
rect 39782 2350 39783 2382
rect 39782 2318 39788 2350
rect 39712 614 39788 2318
rect 39712 550 39718 614
rect 39782 550 39788 614
rect 39712 544 39788 550
rect 40664 0 40740 2862
rect 40805 1702 40871 1703
rect 40805 1670 40806 1702
rect 40800 1638 40806 1670
rect 40870 1670 40871 1702
rect 40870 1638 40876 1670
rect 40800 1294 40876 1638
rect 40800 1230 40806 1294
rect 40870 1230 40876 1294
rect 40800 1224 40876 1230
rect 41072 0 41148 13062
rect 41344 12038 41420 13470
rect 41480 13262 41556 15102
rect 41621 15102 41622 15134
rect 41686 15134 41692 15166
rect 43928 17070 44140 17076
rect 43928 17006 44070 17070
rect 44134 17006 44140 17070
rect 43928 17000 44140 17006
rect 46648 17070 46724 17076
rect 46648 17006 46654 17070
rect 46718 17006 46724 17070
rect 43928 15166 44004 17000
rect 43928 15134 43934 15166
rect 41686 15102 41687 15134
rect 41621 15101 41687 15102
rect 43933 15102 43934 15134
rect 43998 15134 44004 15166
rect 44064 15166 44140 15172
rect 43998 15102 43999 15134
rect 43933 15101 43999 15102
rect 44064 15102 44070 15166
rect 44134 15102 44140 15166
rect 43797 14350 43863 14351
rect 43797 14318 43798 14350
rect 43792 14286 43798 14318
rect 43862 14318 43863 14350
rect 43862 14286 43868 14318
rect 43792 13670 43868 14286
rect 43792 13606 43798 13670
rect 43862 13606 43868 13670
rect 43792 13600 43868 13606
rect 41480 13230 41486 13262
rect 41485 13198 41486 13230
rect 41550 13230 41556 13262
rect 43928 13534 44004 13540
rect 43928 13470 43934 13534
rect 43998 13470 44004 13534
rect 41550 13198 41551 13230
rect 41485 13197 41551 13198
rect 41480 13126 41556 13132
rect 41480 13062 41486 13126
rect 41550 13062 41556 13126
rect 43525 13126 43591 13127
rect 43525 13094 43526 13126
rect 41480 12582 41556 13062
rect 41480 12550 41486 12582
rect 41485 12518 41486 12550
rect 41550 12550 41556 12582
rect 43520 13062 43526 13094
rect 43590 13094 43591 13126
rect 43590 13062 43596 13094
rect 41550 12518 41551 12550
rect 41485 12517 41551 12518
rect 41485 12310 41551 12311
rect 41485 12278 41486 12310
rect 41344 12006 41350 12038
rect 41349 11974 41350 12006
rect 41414 12006 41420 12038
rect 41480 12246 41486 12278
rect 41550 12278 41551 12310
rect 43384 12310 43460 12316
rect 41550 12246 41556 12278
rect 41414 11974 41415 12006
rect 41349 11973 41415 11974
rect 41349 11902 41415 11903
rect 41349 11870 41350 11902
rect 41344 11838 41350 11870
rect 41414 11870 41415 11902
rect 41414 11838 41420 11870
rect 41344 11086 41420 11838
rect 41480 11766 41556 12246
rect 41480 11702 41486 11766
rect 41550 11702 41556 11766
rect 41480 11696 41556 11702
rect 43384 12246 43390 12310
rect 43454 12246 43460 12310
rect 43384 11494 43460 12246
rect 43384 11462 43390 11494
rect 43389 11430 43390 11462
rect 43454 11462 43460 11494
rect 43454 11430 43455 11462
rect 43389 11429 43455 11430
rect 41344 11022 41350 11086
rect 41414 11022 41420 11086
rect 41344 11016 41420 11022
rect 41757 2926 41823 2927
rect 41757 2894 41758 2926
rect 41752 2862 41758 2894
rect 41822 2894 41823 2926
rect 42845 2926 42911 2927
rect 42845 2894 42846 2926
rect 41822 2862 41828 2894
rect 41752 0 41828 2862
rect 42840 2862 42846 2894
rect 42910 2894 42911 2926
rect 42910 2862 42916 2894
rect 42437 1702 42503 1703
rect 42437 1670 42438 1702
rect 42432 1638 42438 1670
rect 42502 1670 42503 1702
rect 42502 1638 42508 1670
rect 42432 1294 42508 1638
rect 42432 1230 42438 1294
rect 42502 1230 42508 1294
rect 42432 1224 42508 1230
rect 42840 0 42916 2862
rect 43520 0 43596 13062
rect 43928 12038 44004 13470
rect 44064 13262 44140 15102
rect 46512 15166 46588 15172
rect 46512 15102 46518 15166
rect 46582 15102 46588 15166
rect 46648 15166 46724 17006
rect 46648 15134 46654 15166
rect 46245 14350 46311 14351
rect 46245 14318 46246 14350
rect 46240 14286 46246 14318
rect 46310 14318 46311 14350
rect 46310 14286 46316 14318
rect 46240 13670 46316 14286
rect 46240 13606 46246 13670
rect 46310 13606 46316 13670
rect 46240 13600 46316 13606
rect 44064 13230 44070 13262
rect 44069 13198 44070 13230
rect 44134 13230 44140 13262
rect 46376 13534 46452 13540
rect 46376 13470 46382 13534
rect 46446 13470 46452 13534
rect 44134 13198 44135 13230
rect 44069 13197 44135 13198
rect 44064 13126 44140 13132
rect 44064 13062 44070 13126
rect 44134 13062 44140 13126
rect 45973 13126 46039 13127
rect 45973 13094 45974 13126
rect 44064 12582 44140 13062
rect 44064 12550 44070 12582
rect 44069 12518 44070 12550
rect 44134 12550 44140 12582
rect 45968 13062 45974 13094
rect 46038 13094 46039 13126
rect 46038 13062 46044 13094
rect 44134 12518 44135 12550
rect 44069 12517 44135 12518
rect 43928 12006 43934 12038
rect 43933 11974 43934 12006
rect 43998 12006 44004 12038
rect 43998 11974 43999 12006
rect 43933 11973 43999 11974
rect 43797 11902 43863 11903
rect 43797 11870 43798 11902
rect 43792 11838 43798 11870
rect 43862 11870 43863 11902
rect 43862 11838 43868 11870
rect 43792 11086 43868 11838
rect 43792 11022 43798 11086
rect 43862 11022 43868 11086
rect 43792 11016 43868 11022
rect 43933 2926 43999 2927
rect 43933 2894 43934 2926
rect 43928 2862 43934 2894
rect 43998 2894 43999 2926
rect 45293 2926 45359 2927
rect 45293 2894 45294 2926
rect 43998 2862 44004 2894
rect 43928 0 44004 2862
rect 45288 2862 45294 2894
rect 45358 2894 45359 2926
rect 45358 2862 45364 2894
rect 44205 1702 44271 1703
rect 44205 1670 44206 1702
rect 44200 1638 44206 1670
rect 44270 1670 44271 1702
rect 44270 1638 44276 1670
rect 44200 1294 44276 1638
rect 44200 1230 44206 1294
rect 44270 1230 44276 1294
rect 44200 1224 44276 1230
rect 45288 0 45364 2862
rect 45701 1702 45767 1703
rect 45701 1670 45702 1702
rect 45696 1638 45702 1670
rect 45766 1670 45767 1702
rect 45766 1638 45772 1670
rect 45696 1294 45772 1638
rect 45696 1230 45702 1294
rect 45766 1230 45772 1294
rect 45696 1224 45772 1230
rect 45968 0 46044 13062
rect 46376 12038 46452 13470
rect 46512 13262 46588 15102
rect 46653 15102 46654 15134
rect 46718 15134 46724 15166
rect 48960 17070 49036 17076
rect 48960 17006 48966 17070
rect 49030 17006 49036 17070
rect 48960 15166 49036 17006
rect 51408 17070 51620 17076
rect 51408 17006 51550 17070
rect 51614 17006 51620 17070
rect 51408 17000 51620 17006
rect 54128 17070 54204 17076
rect 54128 17006 54134 17070
rect 54198 17006 54204 17070
rect 48960 15134 48966 15166
rect 46718 15102 46719 15134
rect 46653 15101 46719 15102
rect 48965 15102 48966 15134
rect 49030 15134 49036 15166
rect 49096 15166 49172 15172
rect 49030 15102 49031 15134
rect 48965 15101 49031 15102
rect 49096 15102 49102 15166
rect 49166 15102 49172 15166
rect 51408 15166 51484 17000
rect 51408 15134 51414 15166
rect 48829 14350 48895 14351
rect 48829 14318 48830 14350
rect 48824 14286 48830 14318
rect 48894 14318 48895 14350
rect 48894 14286 48900 14318
rect 48824 13670 48900 14286
rect 48824 13606 48830 13670
rect 48894 13606 48900 13670
rect 48824 13600 48900 13606
rect 46512 13230 46518 13262
rect 46517 13198 46518 13230
rect 46582 13230 46588 13262
rect 48960 13534 49036 13540
rect 48960 13470 48966 13534
rect 49030 13470 49036 13534
rect 46582 13198 46583 13230
rect 46517 13197 46583 13198
rect 46512 13126 46588 13132
rect 46512 13062 46518 13126
rect 46582 13062 46588 13126
rect 48285 13126 48351 13127
rect 48285 13094 48286 13126
rect 46512 12582 46588 13062
rect 46512 12550 46518 12582
rect 46517 12518 46518 12550
rect 46582 12550 46588 12582
rect 48280 13062 48286 13094
rect 48350 13094 48351 13126
rect 48824 13126 48900 13132
rect 48350 13062 48356 13094
rect 46582 12518 46583 12550
rect 46517 12517 46583 12518
rect 46517 12310 46583 12311
rect 46517 12278 46518 12310
rect 46376 12006 46382 12038
rect 46381 11974 46382 12006
rect 46446 12006 46452 12038
rect 46512 12246 46518 12278
rect 46582 12278 46583 12310
rect 46582 12246 46588 12278
rect 46446 11974 46447 12006
rect 46381 11973 46447 11974
rect 46245 11902 46311 11903
rect 46245 11870 46246 11902
rect 46240 11838 46246 11870
rect 46310 11870 46311 11902
rect 46310 11838 46316 11870
rect 46240 11086 46316 11838
rect 46512 11766 46588 12246
rect 46512 11702 46518 11766
rect 46582 11702 46588 11766
rect 46512 11696 46588 11702
rect 46240 11022 46246 11086
rect 46310 11022 46316 11086
rect 46240 11016 46316 11022
rect 46381 2926 46447 2927
rect 46381 2894 46382 2926
rect 46376 2862 46382 2894
rect 46446 2894 46447 2926
rect 47605 2926 47671 2927
rect 47605 2894 47606 2926
rect 46446 2862 46452 2894
rect 46376 0 46452 2862
rect 47600 2862 47606 2894
rect 47670 2894 47671 2926
rect 47670 2862 47676 2894
rect 47333 1702 47399 1703
rect 47333 1670 47334 1702
rect 47328 1638 47334 1670
rect 47398 1670 47399 1702
rect 47398 1638 47404 1670
rect 47328 1294 47404 1638
rect 47328 1230 47334 1294
rect 47398 1230 47404 1294
rect 47328 1224 47404 1230
rect 47600 0 47676 2862
rect 48280 0 48356 13062
rect 48824 13062 48830 13126
rect 48894 13062 48900 13126
rect 48824 12582 48900 13062
rect 48824 12550 48830 12582
rect 48829 12518 48830 12550
rect 48894 12550 48900 12582
rect 48894 12518 48895 12550
rect 48829 12517 48895 12518
rect 48829 12310 48895 12311
rect 48829 12278 48830 12310
rect 48824 12246 48830 12278
rect 48894 12278 48895 12310
rect 48894 12246 48900 12278
rect 48693 11902 48759 11903
rect 48693 11870 48694 11902
rect 48688 11838 48694 11870
rect 48758 11870 48759 11902
rect 48758 11838 48764 11870
rect 48688 11086 48764 11838
rect 48824 11766 48900 12246
rect 48960 12038 49036 13470
rect 49096 13262 49172 15102
rect 51413 15102 51414 15134
rect 51478 15134 51484 15166
rect 51544 15166 51620 15172
rect 51478 15102 51479 15134
rect 51413 15101 51479 15102
rect 51544 15102 51550 15166
rect 51614 15102 51620 15166
rect 51413 14350 51479 14351
rect 51413 14318 51414 14350
rect 51408 14286 51414 14318
rect 51478 14318 51479 14350
rect 51478 14286 51484 14318
rect 51408 13670 51484 14286
rect 51408 13606 51414 13670
rect 51478 13606 51484 13670
rect 51408 13600 51484 13606
rect 49096 13230 49102 13262
rect 49101 13198 49102 13230
rect 49166 13230 49172 13262
rect 51408 13534 51484 13540
rect 51408 13470 51414 13534
rect 51478 13470 51484 13534
rect 49166 13198 49167 13230
rect 49101 13197 49167 13198
rect 51005 13126 51071 13127
rect 51005 13094 51006 13126
rect 48960 12006 48966 12038
rect 48965 11974 48966 12006
rect 49030 12006 49036 12038
rect 51000 13062 51006 13094
rect 51070 13094 51071 13126
rect 51070 13062 51076 13094
rect 49030 11974 49031 12006
rect 48965 11973 49031 11974
rect 48824 11702 48830 11766
rect 48894 11702 48900 11766
rect 48824 11696 48900 11702
rect 48688 11022 48694 11086
rect 48758 11022 48764 11086
rect 48688 11016 48764 11022
rect 48693 2926 48759 2927
rect 48693 2894 48694 2926
rect 48688 2862 48694 2894
rect 48758 2894 48759 2926
rect 49781 2926 49847 2927
rect 49781 2894 49782 2926
rect 48758 2862 48764 2894
rect 48688 0 48764 2862
rect 49776 2862 49782 2894
rect 49846 2894 49847 2926
rect 49846 2862 49852 2894
rect 49101 1702 49167 1703
rect 49101 1670 49102 1702
rect 49096 1638 49102 1670
rect 49166 1670 49167 1702
rect 49166 1638 49172 1670
rect 49096 1294 49172 1638
rect 49096 1230 49102 1294
rect 49166 1230 49172 1294
rect 49096 1224 49172 1230
rect 49776 0 49852 2862
rect 50733 1702 50799 1703
rect 50733 1670 50734 1702
rect 50728 1638 50734 1670
rect 50798 1670 50799 1702
rect 50798 1638 50804 1670
rect 50728 1294 50804 1638
rect 50728 1230 50734 1294
rect 50798 1230 50804 1294
rect 50728 1224 50804 1230
rect 51000 0 51076 13062
rect 51277 12310 51343 12311
rect 51277 12278 51278 12310
rect 51272 12246 51278 12278
rect 51342 12278 51343 12310
rect 51342 12246 51348 12278
rect 51141 11902 51207 11903
rect 51141 11870 51142 11902
rect 51136 11838 51142 11870
rect 51206 11870 51207 11902
rect 51206 11838 51212 11870
rect 51136 11086 51212 11838
rect 51272 11766 51348 12246
rect 51408 12038 51484 13470
rect 51544 13262 51620 15102
rect 53992 15166 54068 15172
rect 53992 15102 53998 15166
rect 54062 15102 54068 15166
rect 54128 15166 54204 17006
rect 54128 15134 54134 15166
rect 53861 14350 53927 14351
rect 53861 14318 53862 14350
rect 53856 14286 53862 14318
rect 53926 14318 53927 14350
rect 53926 14286 53932 14318
rect 53856 13670 53932 14286
rect 53856 13606 53862 13670
rect 53926 13606 53932 13670
rect 53856 13600 53932 13606
rect 51544 13230 51550 13262
rect 51549 13198 51550 13230
rect 51614 13230 51620 13262
rect 53856 13534 53932 13540
rect 53856 13470 53862 13534
rect 53926 13470 53932 13534
rect 51614 13198 51615 13230
rect 51549 13197 51615 13198
rect 51544 13126 51620 13132
rect 51544 13062 51550 13126
rect 51614 13062 51620 13126
rect 53589 13126 53655 13127
rect 53589 13094 53590 13126
rect 51544 12582 51620 13062
rect 51544 12550 51550 12582
rect 51549 12518 51550 12550
rect 51614 12550 51620 12582
rect 53584 13062 53590 13094
rect 53654 13094 53655 13126
rect 53654 13062 53660 13094
rect 51614 12518 51615 12550
rect 51549 12517 51615 12518
rect 51408 12006 51414 12038
rect 51413 11974 51414 12006
rect 51478 12006 51484 12038
rect 51478 11974 51479 12006
rect 51413 11973 51479 11974
rect 51272 11702 51278 11766
rect 51342 11702 51348 11766
rect 51272 11696 51348 11702
rect 51136 11022 51142 11086
rect 51206 11022 51212 11086
rect 51136 11016 51212 11022
rect 51141 2926 51207 2927
rect 51141 2894 51142 2926
rect 51136 2862 51142 2894
rect 51206 2894 51207 2926
rect 52229 2926 52295 2927
rect 52229 2894 52230 2926
rect 51206 2862 51212 2894
rect 51136 0 51212 2862
rect 52224 2862 52230 2894
rect 52294 2894 52295 2926
rect 53317 2926 53383 2927
rect 53317 2894 53318 2926
rect 52294 2862 52300 2894
rect 52224 0 52300 2862
rect 53312 2862 53318 2894
rect 53382 2894 53383 2926
rect 53382 2862 53388 2894
rect 52501 1702 52567 1703
rect 52501 1670 52502 1702
rect 52496 1638 52502 1670
rect 52566 1670 52567 1702
rect 52566 1638 52572 1670
rect 52496 1294 52572 1638
rect 52496 1230 52502 1294
rect 52566 1230 52572 1294
rect 52496 1224 52572 1230
rect 53312 0 53388 2862
rect 53584 0 53660 13062
rect 53856 12038 53932 13470
rect 53992 13262 54068 15102
rect 54133 15102 54134 15134
rect 54198 15134 54204 15166
rect 56440 17070 56516 17076
rect 56440 17006 56446 17070
rect 56510 17006 56516 17070
rect 56440 15166 56516 17006
rect 56440 15134 56446 15166
rect 54198 15102 54199 15134
rect 54133 15101 54199 15102
rect 56445 15102 56446 15134
rect 56510 15134 56516 15166
rect 56576 15166 56652 15172
rect 56510 15102 56511 15134
rect 56445 15101 56511 15102
rect 56576 15102 56582 15166
rect 56646 15102 56652 15166
rect 56445 14350 56511 14351
rect 56445 14318 56446 14350
rect 56440 14286 56446 14318
rect 56510 14318 56511 14350
rect 56510 14286 56516 14318
rect 56440 13670 56516 14286
rect 56440 13606 56446 13670
rect 56510 13606 56516 13670
rect 56440 13600 56516 13606
rect 53992 13230 53998 13262
rect 53997 13198 53998 13230
rect 54062 13230 54068 13262
rect 56304 13534 56380 13540
rect 56304 13470 56310 13534
rect 56374 13470 56380 13534
rect 54062 13198 54063 13230
rect 53997 13197 54063 13198
rect 53992 13126 54068 13132
rect 53992 13062 53998 13126
rect 54062 13062 54068 13126
rect 56037 13126 56103 13127
rect 56037 13094 56038 13126
rect 53992 12582 54068 13062
rect 53992 12550 53998 12582
rect 53997 12518 53998 12550
rect 54062 12550 54068 12582
rect 56032 13062 56038 13094
rect 56102 13094 56103 13126
rect 56102 13062 56108 13094
rect 54062 12518 54063 12550
rect 53997 12517 54063 12518
rect 53997 12310 54063 12311
rect 53997 12278 53998 12310
rect 53856 12006 53862 12038
rect 53861 11974 53862 12006
rect 53926 12006 53932 12038
rect 53992 12246 53998 12278
rect 54062 12278 54063 12310
rect 54062 12246 54068 12278
rect 53926 11974 53927 12006
rect 53861 11973 53927 11974
rect 53861 11902 53927 11903
rect 53861 11870 53862 11902
rect 53856 11838 53862 11870
rect 53926 11870 53927 11902
rect 53926 11838 53932 11870
rect 53856 11086 53932 11838
rect 53992 11766 54068 12246
rect 53992 11702 53998 11766
rect 54062 11702 54068 11766
rect 53992 11696 54068 11702
rect 53856 11022 53862 11086
rect 53926 11022 53932 11086
rect 53856 11016 53932 11022
rect 54405 2926 54471 2927
rect 54405 2894 54406 2926
rect 54400 2862 54406 2894
rect 54470 2894 54471 2926
rect 55765 2926 55831 2927
rect 55765 2894 55766 2926
rect 54470 2862 54476 2894
rect 54133 1702 54199 1703
rect 54133 1670 54134 1702
rect 54128 1638 54134 1670
rect 54198 1670 54199 1702
rect 54198 1638 54204 1670
rect 54128 1294 54204 1638
rect 54128 1230 54134 1294
rect 54198 1230 54204 1294
rect 54128 1224 54204 1230
rect 54400 0 54476 2862
rect 55760 2862 55766 2894
rect 55830 2894 55831 2926
rect 55830 2862 55836 2894
rect 55493 1702 55559 1703
rect 55493 1670 55494 1702
rect 55488 1638 55494 1670
rect 55558 1670 55559 1702
rect 55558 1638 55564 1670
rect 55488 1294 55564 1638
rect 55488 1230 55494 1294
rect 55558 1230 55564 1294
rect 55488 1224 55564 1230
rect 55760 0 55836 2862
rect 56032 0 56108 13062
rect 56304 12038 56380 13470
rect 56576 13262 56652 15102
rect 58344 14486 58420 18638
rect 119952 18566 120028 20134
rect 122808 20134 122814 20166
rect 122878 20166 122879 20198
rect 122878 20134 122884 20166
rect 122808 19926 122884 20134
rect 122808 19862 122814 19926
rect 122878 19862 122884 19926
rect 122808 19856 122884 19862
rect 119952 18502 119958 18566
rect 120022 18502 120028 18566
rect 119952 18496 120028 18502
rect 122808 19790 122884 19796
rect 122808 19726 122814 19790
rect 122878 19726 122884 19790
rect 59160 17070 59236 17076
rect 59160 17006 59166 17070
rect 59230 17006 59236 17070
rect 58344 14422 58350 14486
rect 58414 14422 58420 14486
rect 58344 14416 58420 14422
rect 59024 15166 59100 15172
rect 59024 15102 59030 15166
rect 59094 15102 59100 15166
rect 59160 15166 59236 17006
rect 61608 17070 61684 17076
rect 61608 17006 61614 17070
rect 61678 17006 61684 17070
rect 59160 15134 59166 15166
rect 58616 14350 58692 14356
rect 58616 14286 58622 14350
rect 58686 14286 58692 14350
rect 58893 14350 58959 14351
rect 58893 14318 58894 14350
rect 58616 13670 58692 14286
rect 58616 13638 58622 13670
rect 58621 13606 58622 13638
rect 58686 13638 58692 13670
rect 58888 14286 58894 14318
rect 58958 14318 58959 14350
rect 58958 14286 58964 14318
rect 58888 13670 58964 14286
rect 58686 13606 58687 13638
rect 58621 13605 58687 13606
rect 58888 13606 58894 13670
rect 58958 13606 58964 13670
rect 58888 13600 58964 13606
rect 56576 13230 56582 13262
rect 56581 13198 56582 13230
rect 56646 13230 56652 13262
rect 58888 13534 58964 13540
rect 58888 13470 58894 13534
rect 58958 13470 58964 13534
rect 56646 13198 56647 13230
rect 56581 13197 56647 13198
rect 56440 13126 56516 13132
rect 56440 13062 56446 13126
rect 56510 13062 56516 13126
rect 58485 13126 58551 13127
rect 58485 13094 58486 13126
rect 56440 12582 56516 13062
rect 56440 12550 56446 12582
rect 56445 12518 56446 12550
rect 56510 12550 56516 12582
rect 58480 13062 58486 13094
rect 58550 13094 58551 13126
rect 58550 13062 58556 13094
rect 56510 12518 56511 12550
rect 56445 12517 56511 12518
rect 56445 12310 56511 12311
rect 56445 12278 56446 12310
rect 56304 12006 56310 12038
rect 56309 11974 56310 12006
rect 56374 12006 56380 12038
rect 56440 12246 56446 12278
rect 56510 12278 56511 12310
rect 56510 12246 56516 12278
rect 56374 11974 56375 12006
rect 56309 11973 56375 11974
rect 56309 11902 56375 11903
rect 56309 11870 56310 11902
rect 56304 11838 56310 11870
rect 56374 11870 56375 11902
rect 56374 11838 56380 11870
rect 56304 11086 56380 11838
rect 56440 11766 56516 12246
rect 56440 11702 56446 11766
rect 56510 11702 56516 11766
rect 56440 11696 56516 11702
rect 56304 11022 56310 11086
rect 56374 11022 56380 11086
rect 56304 11016 56380 11022
rect 56989 2926 57055 2927
rect 56989 2894 56990 2926
rect 56984 2862 56990 2894
rect 57054 2894 57055 2926
rect 58077 2926 58143 2927
rect 58077 2894 58078 2926
rect 57054 2862 57060 2894
rect 56984 0 57060 2862
rect 58072 2862 58078 2894
rect 58142 2894 58143 2926
rect 58142 2862 58148 2894
rect 57533 1702 57599 1703
rect 57533 1670 57534 1702
rect 57528 1638 57534 1670
rect 57598 1670 57599 1702
rect 57598 1638 57604 1670
rect 57528 1294 57604 1638
rect 57528 1230 57534 1294
rect 57598 1230 57604 1294
rect 57528 1224 57604 1230
rect 58072 0 58148 2862
rect 58480 0 58556 13062
rect 58888 12038 58964 13470
rect 59024 13262 59100 15102
rect 59165 15102 59166 15134
rect 59230 15134 59236 15166
rect 61472 15166 61548 15172
rect 59230 15102 59231 15134
rect 59165 15101 59231 15102
rect 61472 15102 61478 15166
rect 61542 15102 61548 15166
rect 61608 15166 61684 17006
rect 61608 15134 61614 15166
rect 61064 14350 61140 14356
rect 61064 14286 61070 14350
rect 61134 14286 61140 14350
rect 61341 14350 61407 14351
rect 61341 14318 61342 14350
rect 61064 13670 61140 14286
rect 61336 14286 61342 14318
rect 61406 14318 61407 14350
rect 61406 14286 61412 14318
rect 61064 13638 61070 13670
rect 61069 13606 61070 13638
rect 61134 13638 61140 13670
rect 61200 13670 61276 13676
rect 61134 13606 61135 13638
rect 61069 13605 61135 13606
rect 61200 13606 61206 13670
rect 61270 13606 61276 13670
rect 59024 13230 59030 13262
rect 59029 13198 59030 13230
rect 59094 13230 59100 13262
rect 59094 13198 59095 13230
rect 59029 13197 59095 13198
rect 59024 13126 59100 13132
rect 59024 13062 59030 13126
rect 59094 13062 59100 13126
rect 60933 13126 60999 13127
rect 60933 13094 60934 13126
rect 59024 12582 59100 13062
rect 59024 12550 59030 12582
rect 59029 12518 59030 12550
rect 59094 12550 59100 12582
rect 60928 13062 60934 13094
rect 60998 13094 60999 13126
rect 60998 13062 61004 13094
rect 59094 12518 59095 12550
rect 59029 12517 59095 12518
rect 59029 12310 59095 12311
rect 59029 12278 59030 12310
rect 58888 12006 58894 12038
rect 58893 11974 58894 12006
rect 58958 12006 58964 12038
rect 59024 12246 59030 12278
rect 59094 12278 59095 12310
rect 59094 12246 59100 12278
rect 58958 11974 58959 12006
rect 58893 11973 58959 11974
rect 58757 11902 58823 11903
rect 58757 11870 58758 11902
rect 58752 11838 58758 11870
rect 58822 11870 58823 11902
rect 58822 11838 58828 11870
rect 58752 11086 58828 11838
rect 59024 11766 59100 12246
rect 59024 11702 59030 11766
rect 59094 11702 59100 11766
rect 59024 11696 59100 11702
rect 58752 11022 58758 11086
rect 58822 11022 58828 11086
rect 58752 11016 58828 11022
rect 59165 2926 59231 2927
rect 59165 2894 59166 2926
rect 59160 2862 59166 2894
rect 59230 2894 59231 2926
rect 59230 2862 59236 2894
rect 59160 0 59236 2862
rect 59437 1702 59503 1703
rect 59437 1670 59438 1702
rect 59432 1638 59438 1670
rect 59502 1670 59503 1702
rect 60797 1702 60863 1703
rect 60797 1670 60798 1702
rect 59502 1638 59508 1670
rect 59432 1294 59508 1638
rect 59432 1230 59438 1294
rect 59502 1230 59508 1294
rect 59432 1224 59508 1230
rect 60792 1638 60798 1670
rect 60862 1670 60863 1702
rect 60862 1638 60868 1670
rect 60792 1294 60868 1638
rect 60792 1230 60798 1294
rect 60862 1230 60868 1294
rect 60792 1224 60868 1230
rect 60928 0 61004 13062
rect 61200 12038 61276 13606
rect 61336 13670 61412 14286
rect 61336 13606 61342 13670
rect 61406 13606 61412 13670
rect 61336 13600 61412 13606
rect 61336 13126 61412 13132
rect 61336 13062 61342 13126
rect 61406 13062 61412 13126
rect 61472 13126 61548 15102
rect 61613 15102 61614 15134
rect 61678 15134 61684 15166
rect 63920 17070 63996 17076
rect 63920 17006 63926 17070
rect 63990 17006 63996 17070
rect 63920 15166 63996 17006
rect 66640 17070 66716 17076
rect 66640 17006 66646 17070
rect 66710 17006 66716 17070
rect 63920 15134 63926 15166
rect 61678 15102 61679 15134
rect 61613 15101 61679 15102
rect 63925 15102 63926 15134
rect 63990 15134 63996 15166
rect 64056 15166 64132 15172
rect 63990 15102 63991 15134
rect 63925 15101 63991 15102
rect 64056 15102 64062 15166
rect 64126 15102 64132 15166
rect 63648 14350 63724 14356
rect 63648 14286 63654 14350
rect 63718 14286 63724 14350
rect 63789 14350 63855 14351
rect 63789 14318 63790 14350
rect 63648 13670 63724 14286
rect 63648 13638 63654 13670
rect 63653 13606 63654 13638
rect 63718 13638 63724 13670
rect 63784 14286 63790 14318
rect 63854 14318 63855 14350
rect 63854 14286 63860 14318
rect 63784 13670 63860 14286
rect 63718 13606 63719 13638
rect 63653 13605 63719 13606
rect 63784 13606 63790 13670
rect 63854 13606 63860 13670
rect 63784 13600 63860 13606
rect 63920 13534 63996 13540
rect 63920 13470 63926 13534
rect 63990 13470 63996 13534
rect 61472 13094 61478 13126
rect 61336 12582 61412 13062
rect 61477 13062 61478 13094
rect 61542 13094 61548 13126
rect 63517 13126 63583 13127
rect 63517 13094 63518 13126
rect 61542 13062 61543 13094
rect 61477 13061 61543 13062
rect 63512 13062 63518 13094
rect 63582 13094 63583 13126
rect 63582 13062 63588 13094
rect 61336 12550 61342 12582
rect 61341 12518 61342 12550
rect 61406 12550 61412 12582
rect 61406 12518 61407 12550
rect 61341 12517 61407 12518
rect 61341 12310 61407 12311
rect 61341 12278 61342 12310
rect 61200 12006 61206 12038
rect 61205 11974 61206 12006
rect 61270 12006 61276 12038
rect 61336 12246 61342 12278
rect 61406 12278 61407 12310
rect 61406 12246 61412 12278
rect 61270 11974 61271 12006
rect 61205 11973 61271 11974
rect 61205 11902 61271 11903
rect 61205 11870 61206 11902
rect 61200 11838 61206 11870
rect 61270 11870 61271 11902
rect 61270 11838 61276 11870
rect 61200 11086 61276 11838
rect 61336 11766 61412 12246
rect 61336 11702 61342 11766
rect 61406 11702 61412 11766
rect 61336 11696 61412 11702
rect 61200 11022 61206 11086
rect 61270 11022 61276 11086
rect 61200 11016 61276 11022
rect 62565 1702 62631 1703
rect 62565 1670 62566 1702
rect 62560 1638 62566 1670
rect 62630 1670 62631 1702
rect 62630 1638 62636 1670
rect 62560 1294 62636 1638
rect 62560 1230 62566 1294
rect 62630 1230 62636 1294
rect 62560 1224 62636 1230
rect 63512 0 63588 13062
rect 63653 12310 63719 12311
rect 63653 12278 63654 12310
rect 63648 12246 63654 12278
rect 63718 12278 63719 12310
rect 63718 12246 63724 12278
rect 63648 11766 63724 12246
rect 63920 12038 63996 13470
rect 64056 13262 64132 15102
rect 66504 15166 66580 15172
rect 66504 15102 66510 15166
rect 66574 15102 66580 15166
rect 66640 15166 66716 17006
rect 69088 17070 69164 17076
rect 69088 17006 69094 17070
rect 69158 17006 69164 17070
rect 66640 15134 66646 15166
rect 66237 14350 66303 14351
rect 66237 14318 66238 14350
rect 66232 14286 66238 14318
rect 66302 14318 66303 14350
rect 66302 14286 66308 14318
rect 66232 13670 66308 14286
rect 66232 13606 66238 13670
rect 66302 13606 66308 13670
rect 66232 13600 66308 13606
rect 64056 13230 64062 13262
rect 64061 13198 64062 13230
rect 64126 13230 64132 13262
rect 66368 13534 66444 13540
rect 66368 13470 66374 13534
rect 66438 13470 66444 13534
rect 64126 13198 64127 13230
rect 64061 13197 64127 13198
rect 64056 13126 64132 13132
rect 64056 13062 64062 13126
rect 64126 13062 64132 13126
rect 65965 13126 66031 13127
rect 65965 13094 65966 13126
rect 64056 12582 64132 13062
rect 64056 12550 64062 12582
rect 64061 12518 64062 12550
rect 64126 12550 64132 12582
rect 65960 13062 65966 13094
rect 66030 13094 66031 13126
rect 66030 13062 66036 13094
rect 64126 12518 64127 12550
rect 64061 12517 64127 12518
rect 63920 12006 63926 12038
rect 63925 11974 63926 12006
rect 63990 12006 63996 12038
rect 63990 11974 63991 12006
rect 63925 11973 63991 11974
rect 63789 11902 63855 11903
rect 63789 11870 63790 11902
rect 63648 11702 63654 11766
rect 63718 11702 63724 11766
rect 63648 11696 63724 11702
rect 63784 11838 63790 11870
rect 63854 11870 63855 11902
rect 63854 11838 63860 11870
rect 63784 11086 63860 11838
rect 63784 11022 63790 11086
rect 63854 11022 63860 11086
rect 63784 11016 63860 11022
rect 64333 1702 64399 1703
rect 64333 1670 64334 1702
rect 64328 1638 64334 1670
rect 64398 1670 64399 1702
rect 65829 1702 65895 1703
rect 65829 1670 65830 1702
rect 64398 1638 64404 1670
rect 64328 1294 64404 1638
rect 64328 1230 64334 1294
rect 64398 1230 64404 1294
rect 64328 1224 64404 1230
rect 65824 1638 65830 1670
rect 65894 1670 65895 1702
rect 65894 1638 65900 1670
rect 65824 1294 65900 1638
rect 65824 1230 65830 1294
rect 65894 1230 65900 1294
rect 65824 1224 65900 1230
rect 65960 0 66036 13062
rect 66237 12310 66303 12311
rect 66237 12278 66238 12310
rect 66232 12246 66238 12278
rect 66302 12278 66303 12310
rect 66302 12246 66308 12278
rect 66101 11902 66167 11903
rect 66101 11870 66102 11902
rect 66096 11838 66102 11870
rect 66166 11870 66167 11902
rect 66166 11838 66172 11870
rect 66096 11086 66172 11838
rect 66232 11766 66308 12246
rect 66368 12038 66444 13470
rect 66504 13262 66580 15102
rect 66645 15102 66646 15134
rect 66710 15134 66716 15166
rect 68952 15166 69028 15172
rect 66710 15102 66711 15134
rect 66645 15101 66711 15102
rect 68952 15102 68958 15166
rect 69022 15102 69028 15166
rect 69088 15166 69164 17006
rect 69088 15134 69094 15166
rect 68821 14350 68887 14351
rect 68821 14318 68822 14350
rect 68816 14286 68822 14318
rect 68886 14318 68887 14350
rect 68886 14286 68892 14318
rect 66504 13230 66510 13262
rect 66509 13198 66510 13230
rect 66574 13230 66580 13262
rect 68680 13670 68756 13676
rect 68680 13606 68686 13670
rect 68750 13606 68756 13670
rect 66574 13198 66575 13230
rect 66509 13197 66575 13198
rect 66504 13126 66580 13132
rect 66504 13062 66510 13126
rect 66574 13062 66580 13126
rect 68277 13126 68343 13127
rect 68277 13094 68278 13126
rect 66504 12582 66580 13062
rect 66504 12550 66510 12582
rect 66509 12518 66510 12550
rect 66574 12550 66580 12582
rect 68272 13062 68278 13094
rect 68342 13094 68343 13126
rect 68342 13062 68348 13094
rect 66574 12518 66575 12550
rect 66509 12517 66575 12518
rect 66368 12006 66374 12038
rect 66373 11974 66374 12006
rect 66438 12006 66444 12038
rect 66438 11974 66439 12006
rect 66373 11973 66439 11974
rect 66232 11702 66238 11766
rect 66302 11702 66308 11766
rect 66232 11696 66308 11702
rect 66096 11022 66102 11086
rect 66166 11022 66172 11086
rect 66096 11016 66172 11022
rect 67597 1702 67663 1703
rect 67597 1670 67598 1702
rect 67592 1638 67598 1670
rect 67662 1670 67663 1702
rect 67662 1638 67668 1670
rect 67592 1294 67668 1638
rect 67592 1230 67598 1294
rect 67662 1230 67668 1294
rect 67592 1224 67668 1230
rect 68272 0 68348 13062
rect 68549 12310 68615 12311
rect 68549 12278 68550 12310
rect 68544 12246 68550 12278
rect 68614 12278 68615 12310
rect 68614 12246 68620 12278
rect 68544 11766 68620 12246
rect 68680 12038 68756 13606
rect 68816 13670 68892 14286
rect 68816 13606 68822 13670
rect 68886 13606 68892 13670
rect 68816 13600 68892 13606
rect 68816 13126 68892 13132
rect 68816 13062 68822 13126
rect 68886 13062 68892 13126
rect 68952 13126 69028 15102
rect 69093 15102 69094 15134
rect 69158 15134 69164 15166
rect 71400 17070 71476 17076
rect 71400 17006 71406 17070
rect 71470 17006 71476 17070
rect 71400 15166 71476 17006
rect 74120 17070 74196 17076
rect 74120 17006 74126 17070
rect 74190 17006 74196 17070
rect 71400 15134 71406 15166
rect 69158 15102 69159 15134
rect 69093 15101 69159 15102
rect 71405 15102 71406 15134
rect 71470 15134 71476 15166
rect 71536 15166 71612 15172
rect 71470 15102 71471 15134
rect 71405 15101 71471 15102
rect 71536 15102 71542 15166
rect 71606 15102 71612 15166
rect 71269 14350 71335 14351
rect 71269 14318 71270 14350
rect 71264 14286 71270 14318
rect 71334 14318 71335 14350
rect 71334 14286 71340 14318
rect 71264 13670 71340 14286
rect 71264 13606 71270 13670
rect 71334 13606 71340 13670
rect 71264 13600 71340 13606
rect 71400 13534 71476 13540
rect 71400 13470 71406 13534
rect 71470 13470 71476 13534
rect 68952 13094 68958 13126
rect 68816 12582 68892 13062
rect 68957 13062 68958 13094
rect 69022 13094 69028 13126
rect 70997 13126 71063 13127
rect 70997 13094 70998 13126
rect 69022 13062 69023 13094
rect 68957 13061 69023 13062
rect 70992 13062 70998 13094
rect 71062 13094 71063 13126
rect 71062 13062 71068 13094
rect 68816 12550 68822 12582
rect 68821 12518 68822 12550
rect 68886 12550 68892 12582
rect 68886 12518 68887 12550
rect 68821 12517 68887 12518
rect 68680 12006 68686 12038
rect 68685 11974 68686 12006
rect 68750 12006 68756 12038
rect 68750 11974 68751 12006
rect 68685 11973 68751 11974
rect 68821 11902 68887 11903
rect 68821 11870 68822 11902
rect 68544 11702 68550 11766
rect 68614 11702 68620 11766
rect 68544 11696 68620 11702
rect 68816 11838 68822 11870
rect 68886 11870 68887 11902
rect 68886 11838 68892 11870
rect 68816 11086 68892 11838
rect 68816 11022 68822 11086
rect 68886 11022 68892 11086
rect 68816 11016 68892 11022
rect 69229 1702 69295 1703
rect 69229 1670 69230 1702
rect 69224 1638 69230 1670
rect 69294 1670 69295 1702
rect 70861 1702 70927 1703
rect 70861 1670 70862 1702
rect 69294 1638 69300 1670
rect 69224 1294 69300 1638
rect 69224 1230 69230 1294
rect 69294 1230 69300 1294
rect 69224 1224 69300 1230
rect 70856 1638 70862 1670
rect 70926 1670 70927 1702
rect 70926 1638 70932 1670
rect 70856 1294 70932 1638
rect 70856 1230 70862 1294
rect 70926 1230 70932 1294
rect 70856 1224 70932 1230
rect 70992 0 71068 13062
rect 71400 12038 71476 13470
rect 71536 13262 71612 15102
rect 73984 15166 74060 15172
rect 73984 15102 73990 15166
rect 74054 15102 74060 15166
rect 74120 15166 74196 17006
rect 74120 15134 74126 15166
rect 73853 14350 73919 14351
rect 73853 14318 73854 14350
rect 73848 14286 73854 14318
rect 73918 14318 73919 14350
rect 73918 14286 73924 14318
rect 73848 13670 73924 14286
rect 73848 13606 73854 13670
rect 73918 13606 73924 13670
rect 73848 13600 73924 13606
rect 71536 13230 71542 13262
rect 71541 13198 71542 13230
rect 71606 13230 71612 13262
rect 73848 13534 73924 13540
rect 73848 13470 73854 13534
rect 73918 13470 73924 13534
rect 71606 13198 71607 13230
rect 71541 13197 71607 13198
rect 71536 13126 71612 13132
rect 71536 13062 71542 13126
rect 71606 13062 71612 13126
rect 73445 13126 73511 13127
rect 73445 13094 73446 13126
rect 71536 12582 71612 13062
rect 71536 12550 71542 12582
rect 71541 12518 71542 12550
rect 71606 12550 71612 12582
rect 73440 13062 73446 13094
rect 73510 13094 73511 13126
rect 73510 13062 73516 13094
rect 71606 12518 71607 12550
rect 71541 12517 71607 12518
rect 71541 12310 71607 12311
rect 71541 12278 71542 12310
rect 71400 12006 71406 12038
rect 71405 11974 71406 12006
rect 71470 12006 71476 12038
rect 71536 12246 71542 12278
rect 71606 12278 71607 12310
rect 73304 12310 73380 12316
rect 71606 12246 71612 12278
rect 71470 11974 71471 12006
rect 71405 11973 71471 11974
rect 71269 11902 71335 11903
rect 71269 11870 71270 11902
rect 71264 11838 71270 11870
rect 71334 11870 71335 11902
rect 71334 11838 71340 11870
rect 71264 11086 71340 11838
rect 71536 11766 71612 12246
rect 71536 11702 71542 11766
rect 71606 11702 71612 11766
rect 71536 11696 71612 11702
rect 73304 12246 73310 12310
rect 73374 12246 73380 12310
rect 73304 11494 73380 12246
rect 73304 11462 73310 11494
rect 73309 11430 73310 11462
rect 73374 11462 73380 11494
rect 73374 11430 73375 11462
rect 73309 11429 73375 11430
rect 71264 11022 71270 11086
rect 71334 11022 71340 11086
rect 71264 11016 71340 11022
rect 72765 1702 72831 1703
rect 72765 1670 72766 1702
rect 72760 1638 72766 1670
rect 72830 1670 72831 1702
rect 72830 1638 72836 1670
rect 72760 1294 72836 1638
rect 72760 1230 72766 1294
rect 72830 1230 72836 1294
rect 72760 1224 72836 1230
rect 73440 0 73516 13062
rect 73848 12038 73924 13470
rect 73984 13262 74060 15102
rect 74125 15102 74126 15134
rect 74190 15134 74196 15166
rect 76432 17070 76508 17076
rect 76432 17006 76438 17070
rect 76502 17006 76508 17070
rect 76432 15166 76508 17006
rect 78880 17070 78956 17076
rect 78880 17006 78886 17070
rect 78950 17006 78956 17070
rect 76432 15134 76438 15166
rect 74190 15102 74191 15134
rect 74125 15101 74191 15102
rect 76437 15102 76438 15134
rect 76502 15134 76508 15166
rect 76568 15166 76644 15172
rect 76502 15102 76503 15134
rect 76437 15101 76503 15102
rect 76568 15102 76574 15166
rect 76638 15102 76644 15166
rect 78880 15166 78956 17006
rect 81600 17070 81676 17076
rect 81600 17006 81606 17070
rect 81670 17006 81676 17070
rect 78880 15134 78886 15166
rect 76024 14350 76100 14356
rect 76024 14286 76030 14350
rect 76094 14286 76100 14350
rect 76301 14350 76367 14351
rect 76301 14318 76302 14350
rect 76024 13670 76100 14286
rect 76024 13638 76030 13670
rect 76029 13606 76030 13638
rect 76094 13638 76100 13670
rect 76296 14286 76302 14318
rect 76366 14318 76367 14350
rect 76366 14286 76372 14318
rect 76296 13670 76372 14286
rect 76094 13606 76095 13638
rect 76029 13605 76095 13606
rect 76296 13606 76302 13670
rect 76366 13606 76372 13670
rect 76296 13600 76372 13606
rect 73984 13230 73990 13262
rect 73989 13198 73990 13230
rect 74054 13230 74060 13262
rect 76432 13534 76508 13540
rect 76432 13470 76438 13534
rect 76502 13470 76508 13534
rect 74054 13198 74055 13230
rect 73989 13197 74055 13198
rect 73984 13126 74060 13132
rect 73984 13062 73990 13126
rect 74054 13062 74060 13126
rect 75893 13126 75959 13127
rect 75893 13094 75894 13126
rect 73984 12582 74060 13062
rect 73984 12550 73990 12582
rect 73989 12518 73990 12550
rect 74054 12550 74060 12582
rect 75888 13062 75894 13094
rect 75958 13094 75959 13126
rect 76296 13126 76372 13132
rect 75958 13062 75964 13094
rect 74054 12518 74055 12550
rect 73989 12517 74055 12518
rect 73848 12006 73854 12038
rect 73853 11974 73854 12006
rect 73918 12006 73924 12038
rect 73918 11974 73919 12006
rect 73853 11973 73919 11974
rect 73717 11902 73783 11903
rect 73717 11870 73718 11902
rect 73712 11838 73718 11870
rect 73782 11870 73783 11902
rect 73782 11838 73788 11870
rect 73712 11086 73788 11838
rect 73712 11022 73718 11086
rect 73782 11022 73788 11086
rect 73712 11016 73788 11022
rect 74261 1702 74327 1703
rect 74261 1670 74262 1702
rect 74256 1638 74262 1670
rect 74326 1670 74327 1702
rect 74326 1638 74332 1670
rect 74256 1294 74332 1638
rect 74256 1230 74262 1294
rect 74326 1230 74332 1294
rect 74256 1224 74332 1230
rect 75888 0 75964 13062
rect 76296 13062 76302 13126
rect 76366 13062 76372 13126
rect 76296 12582 76372 13062
rect 76296 12550 76302 12582
rect 76301 12518 76302 12550
rect 76366 12550 76372 12582
rect 76366 12518 76367 12550
rect 76301 12517 76367 12518
rect 76165 12310 76231 12311
rect 76165 12278 76166 12310
rect 76160 12246 76166 12278
rect 76230 12278 76231 12310
rect 76230 12246 76236 12278
rect 76160 11766 76236 12246
rect 76432 12038 76508 13470
rect 76568 13262 76644 15102
rect 78885 15102 78886 15134
rect 78950 15134 78956 15166
rect 79016 15166 79092 15172
rect 78950 15102 78951 15134
rect 78885 15101 78951 15102
rect 79016 15102 79022 15166
rect 79086 15102 79092 15166
rect 78885 14350 78951 14351
rect 78885 14318 78886 14350
rect 78880 14286 78886 14318
rect 78950 14318 78951 14350
rect 78950 14286 78956 14318
rect 78880 13670 78956 14286
rect 78880 13606 78886 13670
rect 78950 13606 78956 13670
rect 78880 13600 78956 13606
rect 76568 13230 76574 13262
rect 76573 13198 76574 13230
rect 76638 13230 76644 13262
rect 78880 13534 78956 13540
rect 78880 13470 78886 13534
rect 78950 13470 78956 13534
rect 76638 13198 76639 13230
rect 76573 13197 76639 13198
rect 78477 13126 78543 13127
rect 78477 13094 78478 13126
rect 76432 12006 76438 12038
rect 76437 11974 76438 12006
rect 76502 12006 76508 12038
rect 78472 13062 78478 13094
rect 78542 13094 78543 13126
rect 78542 13062 78548 13094
rect 76502 11974 76503 12006
rect 76437 11973 76503 11974
rect 76301 11902 76367 11903
rect 76301 11870 76302 11902
rect 76160 11702 76166 11766
rect 76230 11702 76236 11766
rect 76160 11696 76236 11702
rect 76296 11838 76302 11870
rect 76366 11870 76367 11902
rect 76366 11838 76372 11870
rect 76296 11086 76372 11838
rect 76296 11022 76302 11086
rect 76366 11022 76372 11086
rect 76296 11016 76372 11022
rect 76165 1702 76231 1703
rect 76165 1670 76166 1702
rect 76160 1638 76166 1670
rect 76230 1670 76231 1702
rect 77661 1702 77727 1703
rect 77661 1670 77662 1702
rect 76230 1638 76236 1670
rect 76160 1294 76236 1638
rect 76160 1230 76166 1294
rect 76230 1230 76236 1294
rect 76160 1224 76236 1230
rect 77656 1638 77662 1670
rect 77726 1670 77727 1702
rect 77726 1638 77732 1670
rect 77656 1294 77732 1638
rect 77656 1230 77662 1294
rect 77726 1230 77732 1294
rect 77656 1224 77732 1230
rect 78472 0 78548 13062
rect 78613 12310 78679 12311
rect 78613 12278 78614 12310
rect 78608 12246 78614 12278
rect 78678 12278 78679 12310
rect 78678 12246 78684 12278
rect 78608 11766 78684 12246
rect 78880 12038 78956 13470
rect 79016 13262 79092 15102
rect 81464 15166 81540 15172
rect 81464 15102 81470 15166
rect 81534 15102 81540 15166
rect 81600 15166 81676 17006
rect 81600 15134 81606 15166
rect 81333 14350 81399 14351
rect 81333 14318 81334 14350
rect 81328 14286 81334 14318
rect 81398 14318 81399 14350
rect 81398 14286 81404 14318
rect 81328 13670 81404 14286
rect 81328 13606 81334 13670
rect 81398 13606 81404 13670
rect 81328 13600 81404 13606
rect 79016 13230 79022 13262
rect 79021 13198 79022 13230
rect 79086 13230 79092 13262
rect 81328 13534 81404 13540
rect 81328 13470 81334 13534
rect 81398 13470 81404 13534
rect 79086 13198 79087 13230
rect 79021 13197 79087 13198
rect 79016 13126 79092 13132
rect 79016 13062 79022 13126
rect 79086 13062 79092 13126
rect 80925 13126 80991 13127
rect 80925 13094 80926 13126
rect 79016 12582 79092 13062
rect 79016 12550 79022 12582
rect 79021 12518 79022 12550
rect 79086 12550 79092 12582
rect 80920 13062 80926 13094
rect 80990 13094 80991 13126
rect 80990 13062 80996 13094
rect 79086 12518 79087 12550
rect 79021 12517 79087 12518
rect 78880 12006 78886 12038
rect 78885 11974 78886 12006
rect 78950 12006 78956 12038
rect 78950 11974 78951 12006
rect 78885 11973 78951 11974
rect 78749 11902 78815 11903
rect 78749 11870 78750 11902
rect 78608 11702 78614 11766
rect 78678 11702 78684 11766
rect 78608 11696 78684 11702
rect 78744 11838 78750 11870
rect 78814 11870 78815 11902
rect 78814 11838 78820 11870
rect 78744 11086 78820 11838
rect 78744 11022 78750 11086
rect 78814 11022 78820 11086
rect 78744 11016 78820 11022
rect 79293 1702 79359 1703
rect 79293 1670 79294 1702
rect 79288 1638 79294 1670
rect 79358 1670 79359 1702
rect 79358 1638 79364 1670
rect 79288 1294 79364 1638
rect 79288 1230 79294 1294
rect 79358 1230 79364 1294
rect 79288 1224 79364 1230
rect 80920 0 80996 13062
rect 81061 12310 81127 12311
rect 81061 12278 81062 12310
rect 81056 12246 81062 12278
rect 81126 12278 81127 12310
rect 81126 12246 81132 12278
rect 81056 11766 81132 12246
rect 81328 12038 81404 13470
rect 81464 13262 81540 15102
rect 81605 15102 81606 15134
rect 81670 15134 81676 15166
rect 83912 17070 83988 17076
rect 83912 17006 83918 17070
rect 83982 17006 83988 17070
rect 83912 15166 83988 17006
rect 86360 17070 86436 17076
rect 86360 17006 86366 17070
rect 86430 17006 86436 17070
rect 83912 15134 83918 15166
rect 81670 15102 81671 15134
rect 81605 15101 81671 15102
rect 83917 15102 83918 15134
rect 83982 15134 83988 15166
rect 84048 15166 84124 15172
rect 83982 15102 83983 15134
rect 83917 15101 83983 15102
rect 84048 15102 84054 15166
rect 84118 15102 84124 15166
rect 86360 15166 86436 17006
rect 89080 17070 89156 17076
rect 89080 17006 89086 17070
rect 89150 17006 89156 17070
rect 86360 15134 86366 15166
rect 83645 14350 83711 14351
rect 83645 14318 83646 14350
rect 83640 14286 83646 14318
rect 83710 14318 83711 14350
rect 83710 14286 83716 14318
rect 83640 13670 83716 14286
rect 83640 13606 83646 13670
rect 83710 13606 83716 13670
rect 83640 13600 83716 13606
rect 81464 13230 81470 13262
rect 81469 13198 81470 13230
rect 81534 13230 81540 13262
rect 83912 13534 83988 13540
rect 83912 13470 83918 13534
rect 83982 13470 83988 13534
rect 81534 13198 81535 13230
rect 81469 13197 81535 13198
rect 81464 13126 81540 13132
rect 81464 13062 81470 13126
rect 81534 13062 81540 13126
rect 83509 13126 83575 13127
rect 83509 13094 83510 13126
rect 81464 12582 81540 13062
rect 81464 12550 81470 12582
rect 81469 12518 81470 12550
rect 81534 12550 81540 12582
rect 83504 13062 83510 13094
rect 83574 13094 83575 13126
rect 83776 13126 83852 13132
rect 83574 13062 83580 13094
rect 81534 12518 81535 12550
rect 81469 12517 81535 12518
rect 81328 12006 81334 12038
rect 81333 11974 81334 12006
rect 81398 12006 81404 12038
rect 81398 11974 81399 12006
rect 81333 11973 81399 11974
rect 81197 11902 81263 11903
rect 81197 11870 81198 11902
rect 81056 11702 81062 11766
rect 81126 11702 81132 11766
rect 81056 11696 81132 11702
rect 81192 11838 81198 11870
rect 81262 11870 81263 11902
rect 81262 11838 81268 11870
rect 81192 11086 81268 11838
rect 81192 11022 81198 11086
rect 81262 11022 81268 11086
rect 81192 11016 81268 11022
rect 81061 1702 81127 1703
rect 81061 1670 81062 1702
rect 81056 1638 81062 1670
rect 81126 1670 81127 1702
rect 82829 1702 82895 1703
rect 82829 1670 82830 1702
rect 81126 1638 81132 1670
rect 81056 1294 81132 1638
rect 81056 1230 81062 1294
rect 81126 1230 81132 1294
rect 81056 1224 81132 1230
rect 82824 1638 82830 1670
rect 82894 1670 82895 1702
rect 82894 1638 82900 1670
rect 82824 1294 82900 1638
rect 82824 1230 82830 1294
rect 82894 1230 82900 1294
rect 82824 1224 82900 1230
rect 83504 0 83580 13062
rect 83776 13062 83782 13126
rect 83846 13062 83852 13126
rect 83776 12582 83852 13062
rect 83776 12550 83782 12582
rect 83781 12518 83782 12550
rect 83846 12550 83852 12582
rect 83846 12518 83847 12550
rect 83781 12517 83847 12518
rect 83912 12038 83988 13470
rect 84048 13262 84124 15102
rect 86365 15102 86366 15134
rect 86430 15134 86436 15166
rect 86496 15166 86572 15172
rect 86430 15102 86431 15134
rect 86365 15101 86431 15102
rect 86496 15102 86502 15166
rect 86566 15102 86572 15166
rect 86088 14350 86164 14356
rect 86088 14286 86094 14350
rect 86158 14286 86164 14350
rect 86229 14350 86295 14351
rect 86229 14318 86230 14350
rect 86088 13670 86164 14286
rect 86088 13638 86094 13670
rect 86093 13606 86094 13638
rect 86158 13638 86164 13670
rect 86224 14286 86230 14318
rect 86294 14318 86295 14350
rect 86294 14286 86300 14318
rect 86224 13670 86300 14286
rect 86158 13606 86159 13638
rect 86093 13605 86159 13606
rect 86224 13606 86230 13670
rect 86294 13606 86300 13670
rect 86224 13600 86300 13606
rect 84048 13230 84054 13262
rect 84053 13198 84054 13230
rect 84118 13230 84124 13262
rect 86360 13534 86436 13540
rect 86360 13470 86366 13534
rect 86430 13470 86436 13534
rect 84118 13198 84119 13230
rect 84053 13197 84119 13198
rect 85957 13126 86023 13127
rect 85957 13094 85958 13126
rect 85952 13062 85958 13094
rect 86022 13094 86023 13126
rect 86022 13062 86028 13094
rect 84053 12310 84119 12311
rect 84053 12278 84054 12310
rect 83912 12006 83918 12038
rect 83917 11974 83918 12006
rect 83982 12006 83988 12038
rect 84048 12246 84054 12278
rect 84118 12278 84119 12310
rect 84118 12246 84124 12278
rect 83982 11974 83983 12006
rect 83917 11973 83983 11974
rect 83781 11902 83847 11903
rect 83781 11870 83782 11902
rect 83776 11838 83782 11870
rect 83846 11870 83847 11902
rect 83846 11838 83852 11870
rect 83776 11086 83852 11838
rect 84048 11766 84124 12246
rect 84048 11702 84054 11766
rect 84118 11702 84124 11766
rect 84048 11696 84124 11702
rect 83776 11022 83782 11086
rect 83846 11022 83852 11086
rect 83776 11016 83852 11022
rect 84325 1702 84391 1703
rect 84325 1670 84326 1702
rect 84320 1638 84326 1670
rect 84390 1670 84391 1702
rect 84390 1638 84396 1670
rect 84320 1294 84396 1638
rect 84320 1230 84326 1294
rect 84390 1230 84396 1294
rect 84320 1224 84396 1230
rect 85952 0 86028 13062
rect 86360 12038 86436 13470
rect 86496 13262 86572 15102
rect 88944 15166 89020 15172
rect 88944 15102 88950 15166
rect 89014 15102 89020 15166
rect 89080 15166 89156 17006
rect 89080 15134 89086 15166
rect 88677 14350 88743 14351
rect 88677 14318 88678 14350
rect 88672 14286 88678 14318
rect 88742 14318 88743 14350
rect 88742 14286 88748 14318
rect 88672 13670 88748 14286
rect 88672 13606 88678 13670
rect 88742 13606 88748 13670
rect 88672 13600 88748 13606
rect 86496 13230 86502 13262
rect 86501 13198 86502 13230
rect 86566 13230 86572 13262
rect 88808 13534 88884 13540
rect 88808 13470 88814 13534
rect 88878 13470 88884 13534
rect 86566 13198 86567 13230
rect 86501 13197 86567 13198
rect 86496 13126 86572 13132
rect 86496 13062 86502 13126
rect 86566 13062 86572 13126
rect 88541 13126 88607 13127
rect 88541 13094 88542 13126
rect 86496 12582 86572 13062
rect 86496 12550 86502 12582
rect 86501 12518 86502 12550
rect 86566 12550 86572 12582
rect 88536 13062 88542 13094
rect 88606 13094 88607 13126
rect 88606 13062 88612 13094
rect 86566 12518 86567 12550
rect 86501 12517 86567 12518
rect 86501 12310 86567 12311
rect 86501 12278 86502 12310
rect 86360 12006 86366 12038
rect 86365 11974 86366 12006
rect 86430 12006 86436 12038
rect 86496 12246 86502 12278
rect 86566 12278 86567 12310
rect 86566 12246 86572 12278
rect 86430 11974 86431 12006
rect 86365 11973 86431 11974
rect 86229 11902 86295 11903
rect 86229 11870 86230 11902
rect 86224 11838 86230 11870
rect 86294 11870 86295 11902
rect 86294 11838 86300 11870
rect 86224 11086 86300 11838
rect 86496 11766 86572 12246
rect 86496 11702 86502 11766
rect 86566 11702 86572 11766
rect 86496 11696 86572 11702
rect 86224 11022 86230 11086
rect 86294 11022 86300 11086
rect 86224 11016 86300 11022
rect 86229 1702 86295 1703
rect 86229 1670 86230 1702
rect 86224 1638 86230 1670
rect 86294 1670 86295 1702
rect 87725 1702 87791 1703
rect 87725 1670 87726 1702
rect 86294 1638 86300 1670
rect 86224 1294 86300 1638
rect 86224 1230 86230 1294
rect 86294 1230 86300 1294
rect 86224 1224 86300 1230
rect 87720 1638 87726 1670
rect 87790 1670 87791 1702
rect 87790 1638 87796 1670
rect 87720 1294 87796 1638
rect 87720 1230 87726 1294
rect 87790 1230 87796 1294
rect 87720 1224 87796 1230
rect 88536 0 88612 13062
rect 88808 12038 88884 13470
rect 88944 13262 89020 15102
rect 89085 15102 89086 15134
rect 89150 15134 89156 15166
rect 91392 17070 91468 17076
rect 91392 17006 91398 17070
rect 91462 17006 91468 17070
rect 91392 15166 91468 17006
rect 93840 17070 94052 17076
rect 93840 17006 93982 17070
rect 94046 17006 94052 17070
rect 93840 17000 94052 17006
rect 96560 17070 96636 17076
rect 96560 17006 96566 17070
rect 96630 17006 96636 17070
rect 91392 15134 91398 15166
rect 89150 15102 89151 15134
rect 89085 15101 89151 15102
rect 91397 15102 91398 15134
rect 91462 15134 91468 15166
rect 91528 15166 91604 15172
rect 91462 15102 91463 15134
rect 91397 15101 91463 15102
rect 91528 15102 91534 15166
rect 91598 15102 91604 15166
rect 93840 15166 93916 17000
rect 93840 15134 93846 15166
rect 91261 14350 91327 14351
rect 91261 14318 91262 14350
rect 91256 14286 91262 14318
rect 91326 14318 91327 14350
rect 91326 14286 91332 14318
rect 91256 13670 91332 14286
rect 91256 13606 91262 13670
rect 91326 13606 91332 13670
rect 91256 13600 91332 13606
rect 88944 13230 88950 13262
rect 88949 13198 88950 13230
rect 89014 13230 89020 13262
rect 91392 13534 91468 13540
rect 91392 13470 91398 13534
rect 91462 13470 91468 13534
rect 89014 13198 89015 13230
rect 88949 13197 89015 13198
rect 88944 13126 89020 13132
rect 88944 13062 88950 13126
rect 89014 13062 89020 13126
rect 90989 13126 91055 13127
rect 90989 13094 90990 13126
rect 88944 12582 89020 13062
rect 88944 12550 88950 12582
rect 88949 12518 88950 12550
rect 89014 12550 89020 12582
rect 90984 13062 90990 13094
rect 91054 13094 91055 13126
rect 91256 13126 91332 13132
rect 91054 13062 91060 13094
rect 89014 12518 89015 12550
rect 88949 12517 89015 12518
rect 88949 12310 89015 12311
rect 88949 12278 88950 12310
rect 88808 12006 88814 12038
rect 88813 11974 88814 12006
rect 88878 12006 88884 12038
rect 88944 12246 88950 12278
rect 89014 12278 89015 12310
rect 89014 12246 89020 12278
rect 88878 11974 88879 12006
rect 88813 11973 88879 11974
rect 88813 11902 88879 11903
rect 88813 11870 88814 11902
rect 88808 11838 88814 11870
rect 88878 11870 88879 11902
rect 88878 11838 88884 11870
rect 88808 11086 88884 11838
rect 88944 11766 89020 12246
rect 88944 11702 88950 11766
rect 89014 11702 89020 11766
rect 88944 11696 89020 11702
rect 88808 11022 88814 11086
rect 88878 11022 88884 11086
rect 88808 11016 88884 11022
rect 89357 1702 89423 1703
rect 89357 1670 89358 1702
rect 89352 1638 89358 1670
rect 89422 1670 89423 1702
rect 89422 1638 89428 1670
rect 89352 1294 89428 1638
rect 89352 1230 89358 1294
rect 89422 1230 89428 1294
rect 89352 1224 89428 1230
rect 90984 0 91060 13062
rect 91256 13062 91262 13126
rect 91326 13062 91332 13126
rect 91256 12582 91332 13062
rect 91256 12550 91262 12582
rect 91261 12518 91262 12550
rect 91326 12550 91332 12582
rect 91326 12518 91327 12550
rect 91261 12517 91327 12518
rect 91261 12310 91327 12311
rect 91261 12278 91262 12310
rect 91256 12246 91262 12278
rect 91326 12278 91327 12310
rect 91326 12246 91332 12278
rect 91125 11902 91191 11903
rect 91125 11870 91126 11902
rect 91120 11838 91126 11870
rect 91190 11870 91191 11902
rect 91190 11838 91196 11870
rect 91120 11086 91196 11838
rect 91256 11766 91332 12246
rect 91392 12038 91468 13470
rect 91528 13262 91604 15102
rect 93845 15102 93846 15134
rect 93910 15134 93916 15166
rect 93976 15166 94052 15172
rect 93910 15102 93911 15134
rect 93845 15101 93911 15102
rect 93976 15102 93982 15166
rect 94046 15102 94052 15166
rect 93845 14350 93911 14351
rect 93845 14318 93846 14350
rect 93840 14286 93846 14318
rect 93910 14318 93911 14350
rect 93910 14286 93916 14318
rect 93840 13670 93916 14286
rect 93840 13606 93846 13670
rect 93910 13606 93916 13670
rect 93840 13600 93916 13606
rect 91528 13230 91534 13262
rect 91533 13198 91534 13230
rect 91598 13230 91604 13262
rect 93840 13534 93916 13540
rect 93840 13470 93846 13534
rect 93910 13470 93916 13534
rect 91598 13198 91599 13230
rect 91533 13197 91599 13198
rect 93437 13126 93503 13127
rect 93437 13094 93438 13126
rect 91392 12006 91398 12038
rect 91397 11974 91398 12006
rect 91462 12006 91468 12038
rect 93432 13062 93438 13094
rect 93502 13094 93503 13126
rect 93502 13062 93508 13094
rect 91462 11974 91463 12006
rect 91397 11973 91463 11974
rect 91256 11702 91262 11766
rect 91326 11702 91332 11766
rect 91256 11696 91332 11702
rect 91120 11022 91126 11086
rect 91190 11022 91196 11086
rect 91120 11016 91196 11022
rect 91261 1702 91327 1703
rect 91261 1670 91262 1702
rect 91256 1638 91262 1670
rect 91326 1670 91327 1702
rect 92757 1702 92823 1703
rect 92757 1670 92758 1702
rect 91326 1638 91332 1670
rect 91256 1294 91332 1638
rect 91256 1230 91262 1294
rect 91326 1230 91332 1294
rect 91256 1224 91332 1230
rect 92752 1638 92758 1670
rect 92822 1670 92823 1702
rect 92822 1638 92828 1670
rect 92752 1294 92828 1638
rect 92752 1230 92758 1294
rect 92822 1230 92828 1294
rect 92752 1224 92828 1230
rect 93432 0 93508 13062
rect 93704 12310 93780 12316
rect 93704 12246 93710 12310
rect 93774 12246 93780 12310
rect 93573 11902 93639 11903
rect 93573 11870 93574 11902
rect 93568 11838 93574 11870
rect 93638 11870 93639 11902
rect 93638 11838 93644 11870
rect 93568 11086 93644 11838
rect 93704 11494 93780 12246
rect 93840 12038 93916 13470
rect 93976 13262 94052 15102
rect 96424 15166 96500 15172
rect 96424 15102 96430 15166
rect 96494 15102 96500 15166
rect 96560 15166 96636 17006
rect 96560 15134 96566 15166
rect 96293 14350 96359 14351
rect 96293 14318 96294 14350
rect 96288 14286 96294 14318
rect 96358 14318 96359 14350
rect 96358 14286 96364 14318
rect 96288 13670 96364 14286
rect 96288 13606 96294 13670
rect 96358 13606 96364 13670
rect 96288 13600 96364 13606
rect 93976 13230 93982 13262
rect 93981 13198 93982 13230
rect 94046 13230 94052 13262
rect 96288 13534 96364 13540
rect 96288 13470 96294 13534
rect 96358 13470 96364 13534
rect 94046 13198 94047 13230
rect 93981 13197 94047 13198
rect 93976 13126 94052 13132
rect 93976 13062 93982 13126
rect 94046 13062 94052 13126
rect 95885 13126 95951 13127
rect 95885 13094 95886 13126
rect 93976 12582 94052 13062
rect 93976 12550 93982 12582
rect 93981 12518 93982 12550
rect 94046 12550 94052 12582
rect 95880 13062 95886 13094
rect 95950 13094 95951 13126
rect 95950 13062 95956 13094
rect 94046 12518 94047 12550
rect 93981 12517 94047 12518
rect 93840 12006 93846 12038
rect 93845 11974 93846 12006
rect 93910 12006 93916 12038
rect 93910 11974 93911 12006
rect 93845 11973 93911 11974
rect 93704 11462 93710 11494
rect 93709 11430 93710 11462
rect 93774 11462 93780 11494
rect 93774 11430 93775 11462
rect 93709 11429 93775 11430
rect 93568 11022 93574 11086
rect 93638 11022 93644 11086
rect 93568 11016 93644 11022
rect 94389 1702 94455 1703
rect 94389 1670 94390 1702
rect 94384 1638 94390 1670
rect 94454 1670 94455 1702
rect 94454 1638 94460 1670
rect 94384 1294 94460 1638
rect 94384 1230 94390 1294
rect 94454 1230 94460 1294
rect 94384 1224 94460 1230
rect 95880 0 95956 13062
rect 96021 12310 96087 12311
rect 96021 12278 96022 12310
rect 96016 12246 96022 12278
rect 96086 12278 96087 12310
rect 96086 12246 96092 12278
rect 96016 11766 96092 12246
rect 96288 12038 96364 13470
rect 96424 13262 96500 15102
rect 96565 15102 96566 15134
rect 96630 15134 96636 15166
rect 98872 17070 98948 17076
rect 98872 17006 98878 17070
rect 98942 17006 98948 17070
rect 98872 15166 98948 17006
rect 101592 17070 101668 17076
rect 101592 17006 101598 17070
rect 101662 17006 101668 17070
rect 98872 15134 98878 15166
rect 96630 15102 96631 15134
rect 96565 15101 96631 15102
rect 98877 15102 98878 15134
rect 98942 15134 98948 15166
rect 99008 15166 99084 15172
rect 98942 15102 98943 15134
rect 98877 15101 98943 15102
rect 99008 15102 99014 15166
rect 99078 15102 99084 15166
rect 98877 14350 98943 14351
rect 98877 14318 98878 14350
rect 98872 14286 98878 14318
rect 98942 14318 98943 14350
rect 98942 14286 98948 14318
rect 98872 13670 98948 14286
rect 98872 13606 98878 13670
rect 98942 13606 98948 13670
rect 98872 13600 98948 13606
rect 96424 13230 96430 13262
rect 96429 13198 96430 13230
rect 96494 13230 96500 13262
rect 98872 13534 98948 13540
rect 98872 13470 98878 13534
rect 98942 13470 98948 13534
rect 96494 13198 96495 13230
rect 96429 13197 96495 13198
rect 96424 13126 96500 13132
rect 96424 13062 96430 13126
rect 96494 13062 96500 13126
rect 98469 13126 98535 13127
rect 98469 13094 98470 13126
rect 96424 12582 96500 13062
rect 96424 12550 96430 12582
rect 96429 12518 96430 12550
rect 96494 12550 96500 12582
rect 98464 13062 98470 13094
rect 98534 13094 98535 13126
rect 98534 13062 98540 13094
rect 96494 12518 96495 12550
rect 96429 12517 96495 12518
rect 96288 12006 96294 12038
rect 96293 11974 96294 12006
rect 96358 12006 96364 12038
rect 96358 11974 96359 12006
rect 96293 11973 96359 11974
rect 96157 11902 96223 11903
rect 96157 11870 96158 11902
rect 96016 11702 96022 11766
rect 96086 11702 96092 11766
rect 96016 11696 96092 11702
rect 96152 11838 96158 11870
rect 96222 11870 96223 11902
rect 96222 11838 96228 11870
rect 96152 11086 96228 11838
rect 96152 11022 96158 11086
rect 96222 11022 96228 11086
rect 96152 11016 96228 11022
rect 96157 1702 96223 1703
rect 96157 1670 96158 1702
rect 96152 1638 96158 1670
rect 96222 1670 96223 1702
rect 97789 1702 97855 1703
rect 97789 1670 97790 1702
rect 96222 1638 96228 1670
rect 96152 1294 96228 1638
rect 96152 1230 96158 1294
rect 96222 1230 96228 1294
rect 96152 1224 96228 1230
rect 97784 1638 97790 1670
rect 97854 1670 97855 1702
rect 97854 1638 97860 1670
rect 97784 1294 97860 1638
rect 97784 1230 97790 1294
rect 97854 1230 97860 1294
rect 97784 1224 97860 1230
rect 98464 0 98540 13062
rect 98872 12038 98948 13470
rect 99008 13262 99084 15102
rect 101456 15166 101532 15172
rect 101456 15102 101462 15166
rect 101526 15102 101532 15166
rect 101592 15166 101668 17006
rect 104040 17070 104116 17076
rect 104040 17006 104046 17070
rect 104110 17006 104116 17070
rect 101592 15134 101598 15166
rect 101325 14350 101391 14351
rect 101325 14318 101326 14350
rect 101320 14286 101326 14318
rect 101390 14318 101391 14350
rect 101390 14286 101396 14318
rect 101320 13670 101396 14286
rect 101320 13606 101326 13670
rect 101390 13606 101396 13670
rect 101320 13600 101396 13606
rect 99008 13230 99014 13262
rect 99013 13198 99014 13230
rect 99078 13230 99084 13262
rect 101320 13534 101396 13540
rect 101320 13470 101326 13534
rect 101390 13470 101396 13534
rect 99078 13198 99079 13230
rect 99013 13197 99079 13198
rect 99008 13126 99084 13132
rect 99008 13062 99014 13126
rect 99078 13062 99084 13126
rect 100917 13126 100983 13127
rect 100917 13094 100918 13126
rect 99008 12582 99084 13062
rect 99008 12550 99014 12582
rect 99013 12518 99014 12550
rect 99078 12550 99084 12582
rect 100912 13062 100918 13094
rect 100982 13094 100983 13126
rect 100982 13062 100988 13094
rect 99078 12518 99079 12550
rect 99013 12517 99079 12518
rect 99013 12310 99079 12311
rect 99013 12278 99014 12310
rect 98872 12006 98878 12038
rect 98877 11974 98878 12006
rect 98942 12006 98948 12038
rect 99008 12246 99014 12278
rect 99078 12278 99079 12310
rect 99078 12246 99084 12278
rect 98942 11974 98943 12006
rect 98877 11973 98943 11974
rect 98741 11902 98807 11903
rect 98741 11870 98742 11902
rect 98736 11838 98742 11870
rect 98806 11870 98807 11902
rect 98806 11838 98812 11870
rect 98736 11086 98812 11838
rect 99008 11766 99084 12246
rect 99008 11702 99014 11766
rect 99078 11702 99084 11766
rect 99008 11696 99084 11702
rect 98736 11022 98742 11086
rect 98806 11022 98812 11086
rect 98736 11016 98812 11022
rect 99557 1702 99623 1703
rect 99557 1670 99558 1702
rect 99552 1638 99558 1670
rect 99622 1670 99623 1702
rect 99622 1638 99628 1670
rect 99552 1294 99628 1638
rect 99552 1230 99558 1294
rect 99622 1230 99628 1294
rect 99552 1224 99628 1230
rect 100912 0 100988 13062
rect 101320 12038 101396 13470
rect 101456 13262 101532 15102
rect 101597 15102 101598 15134
rect 101662 15134 101668 15166
rect 103904 15166 103980 15172
rect 101662 15102 101663 15134
rect 101597 15101 101663 15102
rect 103904 15102 103910 15166
rect 103974 15102 103980 15166
rect 104040 15166 104116 17006
rect 104040 15134 104046 15166
rect 103496 14350 103572 14356
rect 103496 14286 103502 14350
rect 103566 14286 103572 14350
rect 103773 14350 103839 14351
rect 103773 14318 103774 14350
rect 103496 13670 103572 14286
rect 103768 14286 103774 14318
rect 103838 14318 103839 14350
rect 103838 14286 103844 14318
rect 103496 13638 103502 13670
rect 103501 13606 103502 13638
rect 103566 13638 103572 13670
rect 103632 13670 103708 13676
rect 103566 13606 103567 13638
rect 103501 13605 103567 13606
rect 103632 13606 103638 13670
rect 103702 13606 103708 13670
rect 101456 13230 101462 13262
rect 101461 13198 101462 13230
rect 101526 13230 101532 13262
rect 101526 13198 101527 13230
rect 101461 13197 101527 13198
rect 101456 13126 101532 13132
rect 101456 13062 101462 13126
rect 101526 13062 101532 13126
rect 103365 13126 103431 13127
rect 103365 13094 103366 13126
rect 101456 12582 101532 13062
rect 101456 12550 101462 12582
rect 101461 12518 101462 12550
rect 101526 12550 101532 12582
rect 103360 13062 103366 13094
rect 103430 13094 103431 13126
rect 103430 13062 103436 13094
rect 101526 12518 101527 12550
rect 101461 12517 101527 12518
rect 101461 12310 101527 12311
rect 101461 12278 101462 12310
rect 101320 12006 101326 12038
rect 101325 11974 101326 12006
rect 101390 12006 101396 12038
rect 101456 12246 101462 12278
rect 101526 12278 101527 12310
rect 101526 12246 101532 12278
rect 101390 11974 101391 12006
rect 101325 11973 101391 11974
rect 101189 11902 101255 11903
rect 101189 11870 101190 11902
rect 101184 11838 101190 11870
rect 101254 11870 101255 11902
rect 101254 11838 101260 11870
rect 101184 11086 101260 11838
rect 101456 11766 101532 12246
rect 101456 11702 101462 11766
rect 101526 11702 101532 11766
rect 101456 11696 101532 11702
rect 101184 11022 101190 11086
rect 101254 11022 101260 11086
rect 101184 11016 101260 11022
rect 101325 1702 101391 1703
rect 101325 1670 101326 1702
rect 101320 1638 101326 1670
rect 101390 1670 101391 1702
rect 102821 1702 102887 1703
rect 102821 1670 102822 1702
rect 101390 1638 101396 1670
rect 101320 1294 101396 1638
rect 101320 1230 101326 1294
rect 101390 1230 101396 1294
rect 101320 1224 101396 1230
rect 102816 1638 102822 1670
rect 102886 1670 102887 1702
rect 102886 1638 102892 1670
rect 102816 1294 102892 1638
rect 102816 1230 102822 1294
rect 102886 1230 102892 1294
rect 102816 1224 102892 1230
rect 103360 0 103436 13062
rect 103632 12038 103708 13606
rect 103768 13670 103844 14286
rect 103768 13606 103774 13670
rect 103838 13606 103844 13670
rect 103768 13600 103844 13606
rect 103768 13126 103844 13132
rect 103768 13062 103774 13126
rect 103838 13062 103844 13126
rect 103904 13126 103980 15102
rect 104045 15102 104046 15134
rect 104110 15134 104116 15166
rect 106352 17070 106428 17076
rect 106352 17006 106358 17070
rect 106422 17006 106428 17070
rect 122808 17070 122884 19726
rect 135320 18974 135668 20542
rect 135320 18910 135326 18974
rect 135390 18910 135668 18974
rect 122949 18430 123015 18431
rect 122949 18398 122950 18430
rect 122808 17038 122814 17070
rect 106352 15166 106428 17006
rect 122813 17006 122814 17038
rect 122878 17038 122884 17070
rect 122944 18366 122950 18398
rect 123014 18398 123015 18430
rect 123014 18366 123020 18398
rect 122878 17006 122879 17038
rect 122813 17005 122879 17006
rect 122813 16934 122879 16935
rect 122813 16902 122814 16934
rect 122808 16870 122814 16902
rect 122878 16902 122879 16934
rect 122878 16870 122884 16902
rect 106352 15134 106358 15166
rect 104110 15102 104111 15134
rect 104045 15101 104111 15102
rect 106357 15102 106358 15134
rect 106422 15134 106428 15166
rect 106488 15166 106564 15172
rect 106422 15102 106423 15134
rect 106357 15101 106423 15102
rect 106488 15102 106494 15166
rect 106558 15102 106564 15166
rect 106357 14350 106423 14351
rect 106357 14318 106358 14350
rect 106352 14286 106358 14318
rect 106422 14318 106423 14350
rect 106422 14286 106428 14318
rect 106352 13670 106428 14286
rect 106352 13606 106358 13670
rect 106422 13606 106428 13670
rect 106352 13600 106428 13606
rect 106352 13534 106428 13540
rect 106352 13470 106358 13534
rect 106422 13470 106428 13534
rect 103904 13094 103910 13126
rect 103768 12582 103844 13062
rect 103909 13062 103910 13094
rect 103974 13094 103980 13126
rect 105949 13126 106015 13127
rect 105949 13094 105950 13126
rect 103974 13062 103975 13094
rect 103909 13061 103975 13062
rect 105944 13062 105950 13094
rect 106014 13094 106015 13126
rect 106014 13062 106020 13094
rect 103768 12550 103774 12582
rect 103773 12518 103774 12550
rect 103838 12550 103844 12582
rect 103838 12518 103839 12550
rect 103773 12517 103839 12518
rect 103773 12310 103839 12311
rect 103773 12278 103774 12310
rect 103632 12006 103638 12038
rect 103637 11974 103638 12006
rect 103702 12006 103708 12038
rect 103768 12246 103774 12278
rect 103838 12278 103839 12310
rect 103838 12246 103844 12278
rect 103702 11974 103703 12006
rect 103637 11973 103703 11974
rect 103637 11902 103703 11903
rect 103637 11870 103638 11902
rect 103632 11838 103638 11870
rect 103702 11870 103703 11902
rect 103702 11838 103708 11870
rect 103632 11086 103708 11838
rect 103768 11766 103844 12246
rect 103768 11702 103774 11766
rect 103838 11702 103844 11766
rect 103768 11696 103844 11702
rect 103632 11022 103638 11086
rect 103702 11022 103708 11086
rect 103632 11016 103708 11022
rect 104589 1702 104655 1703
rect 104589 1670 104590 1702
rect 104584 1638 104590 1670
rect 104654 1670 104655 1702
rect 104654 1638 104660 1670
rect 104584 1294 104660 1638
rect 104584 1230 104590 1294
rect 104654 1230 104660 1294
rect 104584 1224 104660 1230
rect 105944 0 106020 13062
rect 106085 12310 106151 12311
rect 106085 12278 106086 12310
rect 106080 12246 106086 12278
rect 106150 12278 106151 12310
rect 106150 12246 106156 12278
rect 106080 11766 106156 12246
rect 106352 12038 106428 13470
rect 106488 13262 106564 15102
rect 122808 14350 122884 16870
rect 122944 15710 123020 18366
rect 122944 15646 122950 15710
rect 123014 15646 123020 15710
rect 122944 15640 123020 15646
rect 135320 17206 135668 18910
rect 135320 17142 135326 17206
rect 135390 17142 135668 17206
rect 122808 14286 122814 14350
rect 122878 14286 122884 14350
rect 122808 14280 122884 14286
rect 122944 15574 123020 15580
rect 122944 15510 122950 15574
rect 123014 15510 123020 15574
rect 106488 13230 106494 13262
rect 106493 13198 106494 13230
rect 106558 13230 106564 13262
rect 122808 14078 122884 14084
rect 122808 14014 122814 14078
rect 122878 14014 122884 14078
rect 106558 13198 106559 13230
rect 106493 13197 106559 13198
rect 106488 13126 106564 13132
rect 106488 13062 106494 13126
rect 106558 13062 106564 13126
rect 106488 12582 106564 13062
rect 106488 12550 106494 12582
rect 106493 12518 106494 12550
rect 106558 12550 106564 12582
rect 106558 12518 106559 12550
rect 106493 12517 106559 12518
rect 106352 12006 106358 12038
rect 106357 11974 106358 12006
rect 106422 12006 106428 12038
rect 106422 11974 106423 12006
rect 106357 11973 106423 11974
rect 106221 11902 106287 11903
rect 106221 11870 106222 11902
rect 106080 11702 106086 11766
rect 106150 11702 106156 11766
rect 106080 11696 106156 11702
rect 106216 11838 106222 11870
rect 106286 11870 106287 11902
rect 106286 11838 106292 11870
rect 106216 11086 106292 11838
rect 122808 11494 122884 14014
rect 122944 12854 123020 15510
rect 122944 12822 122950 12854
rect 122949 12790 122950 12822
rect 123014 12822 123020 12854
rect 135320 15438 135668 17142
rect 135320 15374 135326 15438
rect 135390 15374 135668 15438
rect 135320 13942 135668 15374
rect 135320 13878 135326 13942
rect 135390 13878 135668 13942
rect 123014 12790 123015 12822
rect 122949 12789 123015 12790
rect 122949 12718 123015 12719
rect 122949 12686 122950 12718
rect 122808 11462 122814 11494
rect 122813 11430 122814 11462
rect 122878 11462 122884 11494
rect 122944 12654 122950 12686
rect 123014 12686 123015 12718
rect 123014 12654 123020 12686
rect 122878 11430 122879 11462
rect 122813 11429 122879 11430
rect 108397 11358 108463 11359
rect 108397 11326 108398 11358
rect 108392 11294 108398 11326
rect 108462 11326 108463 11358
rect 108462 11294 108468 11326
rect 106216 11022 106222 11086
rect 106286 11022 106292 11086
rect 108261 11086 108327 11087
rect 108261 11054 108262 11086
rect 106216 11016 106292 11022
rect 108256 11022 108262 11054
rect 108326 11054 108327 11086
rect 108326 11022 108332 11054
rect 108256 10678 108332 11022
rect 108256 10614 108262 10678
rect 108326 10614 108332 10678
rect 108256 10608 108332 10614
rect 108392 9590 108468 11294
rect 122944 9998 123020 12654
rect 135320 12310 135668 13878
rect 135320 12246 135326 12310
rect 135390 12246 135668 12310
rect 123221 11902 123287 11903
rect 123221 11870 123222 11902
rect 122944 9934 122950 9998
rect 123014 9934 123020 9998
rect 122944 9928 123020 9934
rect 123216 11838 123222 11870
rect 123286 11870 123287 11902
rect 123286 11838 123292 11870
rect 108392 9526 108398 9590
rect 108462 9526 108468 9590
rect 108392 9520 108468 9526
rect 106221 1702 106287 1703
rect 106221 1670 106222 1702
rect 106216 1638 106222 1670
rect 106286 1670 106287 1702
rect 107853 1702 107919 1703
rect 107853 1670 107854 1702
rect 106286 1638 106292 1670
rect 106216 1294 106292 1638
rect 106216 1230 106222 1294
rect 106286 1230 106292 1294
rect 106216 1224 106292 1230
rect 107848 1638 107854 1670
rect 107918 1670 107919 1702
rect 109757 1702 109823 1703
rect 109757 1670 109758 1702
rect 107918 1638 107924 1670
rect 107848 1294 107924 1638
rect 107848 1230 107854 1294
rect 107918 1230 107924 1294
rect 107848 1224 107924 1230
rect 109752 1638 109758 1670
rect 109822 1670 109823 1702
rect 111253 1702 111319 1703
rect 111253 1670 111254 1702
rect 109822 1638 109828 1670
rect 109752 1294 109828 1638
rect 109752 1230 109758 1294
rect 109822 1230 109828 1294
rect 109752 1224 109828 1230
rect 111248 1638 111254 1670
rect 111318 1670 111319 1702
rect 113021 1702 113087 1703
rect 113021 1670 113022 1702
rect 111318 1638 111324 1670
rect 111248 1294 111324 1638
rect 111248 1230 111254 1294
rect 111318 1230 111324 1294
rect 111248 1224 111324 1230
rect 113016 1638 113022 1670
rect 113086 1670 113087 1702
rect 114789 1702 114855 1703
rect 114789 1670 114790 1702
rect 113086 1638 113092 1670
rect 113016 1294 113092 1638
rect 113016 1230 113022 1294
rect 113086 1230 113092 1294
rect 113016 1224 113092 1230
rect 114784 1638 114790 1670
rect 114854 1670 114855 1702
rect 116285 1702 116351 1703
rect 116285 1670 116286 1702
rect 114854 1638 114860 1670
rect 114784 1294 114860 1638
rect 114784 1230 114790 1294
rect 114854 1230 114860 1294
rect 114784 1224 114860 1230
rect 116280 1638 116286 1670
rect 116350 1670 116351 1702
rect 118053 1702 118119 1703
rect 118053 1670 118054 1702
rect 116350 1638 116356 1670
rect 116280 1294 116356 1638
rect 116280 1230 116286 1294
rect 116350 1230 116356 1294
rect 116280 1224 116356 1230
rect 118048 1638 118054 1670
rect 118118 1670 118119 1702
rect 119821 1702 119887 1703
rect 119821 1670 119822 1702
rect 118118 1638 118124 1670
rect 118048 1294 118124 1638
rect 118048 1230 118054 1294
rect 118118 1230 118124 1294
rect 118048 1224 118124 1230
rect 119816 1638 119822 1670
rect 119886 1670 119887 1702
rect 121317 1702 121383 1703
rect 121317 1670 121318 1702
rect 119886 1638 119892 1670
rect 119816 1294 119892 1638
rect 119816 1230 119822 1294
rect 119886 1230 119892 1294
rect 119816 1224 119892 1230
rect 121312 1638 121318 1670
rect 121382 1670 121383 1702
rect 123085 1702 123151 1703
rect 123085 1670 123086 1702
rect 121382 1638 121388 1670
rect 121312 1294 121388 1638
rect 121312 1230 121318 1294
rect 121382 1230 121388 1294
rect 121312 1224 121388 1230
rect 123080 1638 123086 1670
rect 123150 1670 123151 1702
rect 123150 1638 123156 1670
rect 123080 1294 123156 1638
rect 123080 1230 123086 1294
rect 123150 1230 123156 1294
rect 123080 1224 123156 1230
rect 123216 0 123292 11838
rect 123357 10814 123423 10815
rect 123357 10782 123358 10814
rect 123352 10750 123358 10782
rect 123422 10782 123423 10814
rect 123422 10750 123428 10782
rect 123352 0 123428 10750
rect 135320 10406 135668 12246
rect 135320 10342 135326 10406
rect 135390 10342 135668 10406
rect 135320 8774 135668 10342
rect 135320 8710 135326 8774
rect 135390 8710 135668 8774
rect 135320 7142 135668 8710
rect 135320 7078 135326 7142
rect 135390 7078 135668 7142
rect 135320 5374 135668 7078
rect 135320 5310 135326 5374
rect 135390 5310 135668 5374
rect 135320 3742 135668 5310
rect 135320 3678 135326 3742
rect 135390 3678 135668 3742
rect 135320 2110 135668 3678
rect 135320 2046 135326 2110
rect 135390 2046 135668 2110
rect 124717 1702 124783 1703
rect 124717 1670 124718 1702
rect 124712 1638 124718 1670
rect 124782 1670 124783 1702
rect 126349 1702 126415 1703
rect 126349 1670 126350 1702
rect 124782 1638 124788 1670
rect 124712 1294 124788 1638
rect 124712 1230 124718 1294
rect 124782 1230 124788 1294
rect 124712 1224 124788 1230
rect 126344 1638 126350 1670
rect 126414 1670 126415 1702
rect 127981 1702 128047 1703
rect 127981 1670 127982 1702
rect 126414 1638 126420 1670
rect 126344 1294 126420 1638
rect 126344 1230 126350 1294
rect 126414 1230 126420 1294
rect 126344 1224 126420 1230
rect 127976 1638 127982 1670
rect 128046 1670 128047 1702
rect 129749 1702 129815 1703
rect 129749 1670 129750 1702
rect 128046 1638 128052 1670
rect 127976 1294 128052 1638
rect 127976 1230 127982 1294
rect 128046 1230 128052 1294
rect 127976 1224 128052 1230
rect 129744 1638 129750 1670
rect 129814 1670 129815 1702
rect 131517 1702 131583 1703
rect 131517 1670 131518 1702
rect 129814 1638 129820 1670
rect 129744 1294 129820 1638
rect 129744 1230 129750 1294
rect 129814 1230 129820 1294
rect 129744 1224 129820 1230
rect 131512 1638 131518 1670
rect 131582 1670 131583 1702
rect 133149 1702 133215 1703
rect 133149 1670 133150 1702
rect 131582 1638 131588 1670
rect 131512 1294 131588 1638
rect 131512 1230 131518 1294
rect 131582 1230 131588 1294
rect 131512 1224 131588 1230
rect 133144 1638 133150 1670
rect 133214 1670 133215 1702
rect 133214 1638 133220 1670
rect 133144 1294 133220 1638
rect 133144 1230 133150 1294
rect 133214 1230 133220 1294
rect 133144 1224 133220 1230
rect 135320 1294 135668 2046
rect 135320 1230 135326 1294
rect 135390 1230 135462 1294
rect 135526 1230 135598 1294
rect 135662 1230 135668 1294
rect 135320 1158 135668 1230
rect 135320 1094 135326 1158
rect 135390 1094 135462 1158
rect 135526 1094 135598 1158
rect 135662 1094 135668 1158
rect 135320 1022 135668 1094
rect 135320 958 135326 1022
rect 135390 958 135462 1022
rect 135526 958 135598 1022
rect 135662 958 135668 1022
rect 135320 952 135668 958
rect 136000 79902 136348 82694
rect 136000 79838 136006 79902
rect 136070 79838 136348 79902
rect 136000 72830 136348 79838
rect 136000 72766 136006 72830
rect 136070 72766 136348 72830
rect 136000 64534 136348 72766
rect 136000 64470 136006 64534
rect 136070 64470 136348 64534
rect 136000 614 136348 64470
rect 136000 550 136006 614
rect 136070 550 136142 614
rect 136206 550 136278 614
rect 136342 550 136348 614
rect 136000 478 136348 550
rect 136000 414 136006 478
rect 136070 414 136142 478
rect 136206 414 136278 478
rect 136342 414 136348 478
rect 136000 342 136348 414
rect 136000 278 136006 342
rect 136070 278 136142 342
rect 136206 278 136278 342
rect 136342 278 136348 342
rect 136000 272 136348 278
use sky130_sram_2kbyte_1rw1r_32x512_8_bank  sky130_sram_2kbyte_1rw1r_32x512_8_bank_0
timestamp 1649977179
transform 1 0 14862 0 1 9422
box 0 0 107270 69282
use sky130_sram_2kbyte_1rw1r_32x512_8_col_addr_dff  sky130_sram_2kbyte_1rw1r_32x512_8_col_addr_dff_0
timestamp 1649977179
transform 1 0 15862 0 1 2396
box -36 -49 2372 1467
use sky130_sram_2kbyte_1rw1r_32x512_8_col_addr_dff  sky130_sram_2kbyte_1rw1r_32x512_8_col_addr_dff_1
timestamp 1649977179
transform -1 0 119964 0 -1 80801
box -36 -49 2372 1467
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_0
timestamp 1649977179
transform 1 0 134839 0 1 2023
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_1
timestamp 1649977179
transform 1 0 133165 0 1 1687
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_2
timestamp 1649977179
transform 1 0 131485 0 1 1687
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_3
timestamp 1649977179
transform 1 0 129805 0 1 1687
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_4
timestamp 1649977179
transform 1 0 128125 0 1 1687
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_5
timestamp 1649977179
transform 1 0 134839 0 1 3703
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_6
timestamp 1649977179
transform 1 0 124765 0 1 1687
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_7
timestamp 1649977179
transform 1 0 123085 0 1 1687
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_8
timestamp 1649977179
transform 1 0 121405 0 1 1687
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_9
timestamp 1649977179
transform 1 0 119725 0 1 1687
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_10
timestamp 1649977179
transform 1 0 126445 0 1 1687
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_11
timestamp 1649977179
transform 1 0 134839 0 1 10423
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_12
timestamp 1649977179
transform 1 0 134839 0 1 8743
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_13
timestamp 1649977179
transform 1 0 134839 0 1 7063
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_14
timestamp 1649977179
transform 1 0 134839 0 1 5383
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_15
timestamp 1649977179
transform 1 0 114685 0 1 1687
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_16
timestamp 1649977179
transform 1 0 111325 0 1 1687
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_17
timestamp 1649977179
transform 1 0 113005 0 1 1687
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_18
timestamp 1649977179
transform 1 0 118045 0 1 1687
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_19
timestamp 1649977179
transform 1 0 116365 0 1 1687
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_20
timestamp 1649977179
transform 1 0 102925 0 1 1687
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_21
timestamp 1649977179
transform 1 0 107965 0 1 1687
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_22
timestamp 1649977179
transform 1 0 104605 0 1 1687
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_23
timestamp 1649977179
transform 1 0 106285 0 1 1687
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_24
timestamp 1649977179
transform 1 0 109645 0 1 1687
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_25
timestamp 1649977179
transform 1 0 105989 0 1 13196
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_26
timestamp 1649977179
transform 1 0 103493 0 1 13196
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_27
timestamp 1649977179
transform 1 0 134839 0 1 13783
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_28
timestamp 1649977179
transform 1 0 134839 0 1 12103
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_29
timestamp 1649977179
transform 1 0 134839 0 1 15463
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_30
timestamp 1649977179
transform 1 0 122320 0 1 14788
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_31
timestamp 1649977179
transform 1 0 123265 0 1 10761
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_32
timestamp 1649977179
transform 1 0 123265 0 1 11889
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_33
timestamp 1649977179
transform 1 0 123265 0 1 13589
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_34
timestamp 1649977179
transform 1 0 123265 0 1 14717
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_35
timestamp 1649977179
transform 1 0 121662 0 1 13518
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_36
timestamp 1649977179
transform 1 0 122320 0 1 13518
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_37
timestamp 1649977179
transform 1 0 121742 0 1 14788
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_38
timestamp 1649977179
transform 1 0 121502 0 1 10690
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_39
timestamp 1649977179
transform 1 0 122320 0 1 10690
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_40
timestamp 1649977179
transform 1 0 121582 0 1 11960
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_41
timestamp 1649977179
transform 1 0 122320 0 1 11960
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_42
timestamp 1649977179
transform 1 0 121822 0 1 16346
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_43
timestamp 1649977179
transform 1 0 122320 0 1 16346
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_44
timestamp 1649977179
transform 1 0 121902 0 1 17616
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_45
timestamp 1649977179
transform 1 0 122320 0 1 17616
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_46
timestamp 1649977179
transform 1 0 121982 0 1 19174
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_47
timestamp 1649977179
transform 1 0 122320 0 1 19174
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_48
timestamp 1649977179
transform 1 0 123265 0 1 16417
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_49
timestamp 1649977179
transform 1 0 123265 0 1 17545
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_50
timestamp 1649977179
transform 1 0 123265 0 1 19245
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_51
timestamp 1649977179
transform 1 0 134839 0 1 20503
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_52
timestamp 1649977179
transform 1 0 134839 0 1 18823
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_53
timestamp 1649977179
transform 1 0 134839 0 1 17143
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_54
timestamp 1649977179
transform 1 0 94525 0 1 1687
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_55
timestamp 1649977179
transform 1 0 96205 0 1 1687
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_56
timestamp 1649977179
transform 1 0 101245 0 1 1687
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_57
timestamp 1649977179
transform 1 0 97885 0 1 1687
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_58
timestamp 1649977179
transform 1 0 99565 0 1 1687
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_59
timestamp 1649977179
transform 1 0 86125 0 1 1687
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_60
timestamp 1649977179
transform 1 0 89485 0 1 1687
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_61
timestamp 1649977179
transform 1 0 91165 0 1 1687
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_62
timestamp 1649977179
transform 1 0 87805 0 1 1687
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_63
timestamp 1649977179
transform 1 0 92845 0 1 1687
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_64
timestamp 1649977179
transform 1 0 77725 0 1 1687
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_65
timestamp 1649977179
transform 1 0 84445 0 1 1687
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_66
timestamp 1649977179
transform 1 0 81085 0 1 1687
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_67
timestamp 1649977179
transform 1 0 82765 0 1 1687
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_68
timestamp 1649977179
transform 1 0 79405 0 1 1687
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_69
timestamp 1649977179
transform 1 0 74365 0 1 1687
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_70
timestamp 1649977179
transform 1 0 76045 0 1 1687
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_71
timestamp 1649977179
transform 1 0 72685 0 1 1687
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_72
timestamp 1649977179
transform 1 0 71005 0 1 1687
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_73
timestamp 1649977179
transform 1 0 69325 0 1 1687
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_74
timestamp 1649977179
transform 1 0 83525 0 1 13196
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_75
timestamp 1649977179
transform 1 0 81029 0 1 13196
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_76
timestamp 1649977179
transform 1 0 78533 0 1 13196
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_77
timestamp 1649977179
transform 1 0 76037 0 1 13196
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_78
timestamp 1649977179
transform 1 0 73541 0 1 13196
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_79
timestamp 1649977179
transform 1 0 71045 0 1 13196
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_80
timestamp 1649977179
transform 1 0 68549 0 1 13196
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_81
timestamp 1649977179
transform 1 0 100997 0 1 13196
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_82
timestamp 1649977179
transform 1 0 98501 0 1 13196
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_83
timestamp 1649977179
transform 1 0 96005 0 1 13196
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_84
timestamp 1649977179
transform 1 0 93509 0 1 13196
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_85
timestamp 1649977179
transform 1 0 91013 0 1 13196
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_86
timestamp 1649977179
transform 1 0 88517 0 1 13196
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_87
timestamp 1649977179
transform 1 0 86021 0 1 13196
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_88
timestamp 1649977179
transform 1 0 134839 0 1 23863
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_89
timestamp 1649977179
transform 1 0 134839 0 1 22183
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_90
timestamp 1649977179
transform 1 0 134839 0 1 25543
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_91
timestamp 1649977179
transform 1 0 134839 0 1 27223
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_92
timestamp 1649977179
transform 1 0 134839 0 1 30583
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_93
timestamp 1649977179
transform 1 0 134839 0 1 28903
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_94
timestamp 1649977179
transform 1 0 134839 0 1 35623
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_95
timestamp 1649977179
transform 1 0 134839 0 1 33943
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_96
timestamp 1649977179
transform 1 0 134839 0 1 32263
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_97
timestamp 1649977179
transform 1 0 134839 0 1 40663
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_98
timestamp 1649977179
transform 1 0 134839 0 1 38983
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_99
timestamp 1649977179
transform 1 0 134839 0 1 37303
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_100
timestamp 1649977179
transform 1 0 65965 0 1 1687
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_101
timestamp 1649977179
transform 1 0 60925 0 1 1687
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_102
timestamp 1649977179
transform 1 0 64285 0 1 1687
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_103
timestamp 1649977179
transform 1 0 62605 0 1 1687
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_104
timestamp 1649977179
transform 1 0 67645 0 1 1687
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_105
timestamp 1649977179
transform 1 0 59245 0 1 1687
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_106
timestamp 1649977179
transform 1 0 55885 0 1 1687
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_107
timestamp 1649977179
transform 1 0 57565 0 1 1687
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_108
timestamp 1649977179
transform 1 0 52207 0 1 2923
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_109
timestamp 1649977179
transform 1 0 54205 0 1 1687
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_110
timestamp 1649977179
transform 1 0 52525 0 1 1687
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_111
timestamp 1649977179
transform 1 0 59215 0 1 2923
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_112
timestamp 1649977179
transform 1 0 58047 0 1 2923
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_113
timestamp 1649977179
transform 1 0 56879 0 1 2923
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_114
timestamp 1649977179
transform 1 0 55711 0 1 2923
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_115
timestamp 1649977179
transform 1 0 54543 0 1 2923
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_116
timestamp 1649977179
transform 1 0 53375 0 1 2923
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_117
timestamp 1649977179
transform 1 0 47485 0 1 1687
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_118
timestamp 1649977179
transform 1 0 49871 0 1 2923
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_119
timestamp 1649977179
transform 1 0 48703 0 1 2923
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_120
timestamp 1649977179
transform 1 0 45805 0 1 1687
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_121
timestamp 1649977179
transform 1 0 47535 0 1 2923
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_122
timestamp 1649977179
transform 1 0 46367 0 1 2923
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_123
timestamp 1649977179
transform 1 0 51039 0 1 2923
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_124
timestamp 1649977179
transform 1 0 50845 0 1 1687
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_125
timestamp 1649977179
transform 1 0 42863 0 1 2923
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_126
timestamp 1649977179
transform 1 0 45199 0 1 2923
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_127
timestamp 1649977179
transform 1 0 49165 0 1 1687
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_128
timestamp 1649977179
transform 1 0 44031 0 1 2923
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_129
timestamp 1649977179
transform 1 0 44125 0 1 1687
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_130
timestamp 1649977179
transform 1 0 39085 0 1 1687
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_131
timestamp 1649977179
transform 1 0 37405 0 1 1687
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_132
timestamp 1649977179
transform 1 0 35725 0 1 1687
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_133
timestamp 1649977179
transform 1 0 35855 0 1 2923
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_134
timestamp 1649977179
transform 1 0 41695 0 1 2923
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_135
timestamp 1649977179
transform 1 0 40527 0 1 2923
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_136
timestamp 1649977179
transform 1 0 39359 0 1 2923
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_137
timestamp 1649977179
transform 1 0 34687 0 1 2923
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_138
timestamp 1649977179
transform 1 0 38191 0 1 2923
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_139
timestamp 1649977179
transform 1 0 42445 0 1 1687
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_140
timestamp 1649977179
transform 1 0 40765 0 1 1687
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_141
timestamp 1649977179
transform 1 0 37023 0 1 2923
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_142
timestamp 1649977179
transform 1 0 51077 0 1 13196
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_143
timestamp 1649977179
transform 1 0 48581 0 1 13196
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_144
timestamp 1649977179
transform 1 0 46085 0 1 13196
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_145
timestamp 1649977179
transform 1 0 43589 0 1 13196
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_146
timestamp 1649977179
transform 1 0 41093 0 1 13196
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_147
timestamp 1649977179
transform 1 0 38597 0 1 13196
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_148
timestamp 1649977179
transform 1 0 36101 0 1 13196
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_149
timestamp 1649977179
transform 1 0 66053 0 1 13196
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_150
timestamp 1649977179
transform 1 0 63557 0 1 13196
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_151
timestamp 1649977179
transform 1 0 61061 0 1 13196
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_152
timestamp 1649977179
transform 1 0 58565 0 1 13196
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_153
timestamp 1649977179
transform 1 0 56069 0 1 13196
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_154
timestamp 1649977179
transform 1 0 53573 0 1 13196
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_155
timestamp 1649977179
transform 1 0 27325 0 1 1687
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_156
timestamp 1649977179
transform 1 0 32365 0 1 1687
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_157
timestamp 1649977179
transform 1 0 33519 0 1 2923
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_158
timestamp 1649977179
transform 1 0 32351 0 1 2923
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_159
timestamp 1649977179
transform 1 0 31183 0 1 2923
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_160
timestamp 1649977179
transform 1 0 30015 0 1 2923
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_161
timestamp 1649977179
transform 1 0 28847 0 1 2923
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_162
timestamp 1649977179
transform 1 0 27679 0 1 2923
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_163
timestamp 1649977179
transform 1 0 26511 0 1 2923
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_164
timestamp 1649977179
transform 1 0 30685 0 1 1687
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_165
timestamp 1649977179
transform 1 0 34045 0 1 1687
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_166
timestamp 1649977179
transform 1 0 29005 0 1 1687
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_167
timestamp 1649977179
transform 1 0 20605 0 1 1687
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_168
timestamp 1649977179
transform 1 0 25343 0 1 2923
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_169
timestamp 1649977179
transform 1 0 24175 0 1 2923
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_170
timestamp 1649977179
transform 1 0 23007 0 1 2923
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_171
timestamp 1649977179
transform 1 0 25645 0 1 1687
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_172
timestamp 1649977179
transform 1 0 23965 0 1 1687
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_173
timestamp 1649977179
transform 1 0 22285 0 1 1687
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_174
timestamp 1649977179
transform 1 0 18925 0 1 1687
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_175
timestamp 1649977179
transform 1 0 21839 0 1 2923
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_176
timestamp 1649977179
transform 1 0 20671 0 1 2923
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_177
timestamp 1649977179
transform 1 0 19503 0 1 2923
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_178
timestamp 1649977179
transform 1 0 18335 0 1 2923
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_179
timestamp 1649977179
transform 1 0 8845 0 1 1687
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_180
timestamp 1649977179
transform 1 0 12205 0 1 1687
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_181
timestamp 1649977179
transform 1 0 17167 0 1 2923
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_182
timestamp 1649977179
transform 1 0 15999 0 1 2923
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_183
timestamp 1649977179
transform 1 0 10525 0 1 1687
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_184
timestamp 1649977179
transform 1 0 15565 0 1 1687
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_185
timestamp 1649977179
transform 1 0 13885 0 1 1687
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_186
timestamp 1649977179
transform 1 0 5485 0 1 1687
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_187
timestamp 1649977179
transform 1 0 7165 0 1 1687
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_188
timestamp 1649977179
transform 1 0 3805 0 1 1687
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_189
timestamp 1649977179
transform 1 0 2125 0 1 1687
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_190
timestamp 1649977179
transform 1 0 1789 0 1 2023
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_191
timestamp 1649977179
transform 1 0 1789 0 1 3703
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_192
timestamp 1649977179
transform 1 0 1789 0 1 10423
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_193
timestamp 1649977179
transform 1 0 5970 0 1 8252
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_194
timestamp 1649977179
transform 1 0 2749 0 1 9847
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_195
timestamp 1649977179
transform 1 0 2749 0 1 8147
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_196
timestamp 1649977179
transform 1 0 1789 0 1 8743
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_197
timestamp 1649977179
transform 1 0 1789 0 1 7063
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_198
timestamp 1649977179
transform 1 0 1789 0 1 5383
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_199
timestamp 1649977179
transform 1 0 14661 0 1 15360
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_200
timestamp 1649977179
transform 1 0 14661 0 1 13946
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_201
timestamp 1649977179
transform 1 0 14661 0 1 12532
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_202
timestamp 1649977179
transform 1 0 1789 0 1 15463
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_203
timestamp 1649977179
transform 1 0 1789 0 1 12103
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_204
timestamp 1649977179
transform 1 0 1789 0 1 13783
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_205
timestamp 1649977179
transform 1 0 1789 0 1 20503
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_206
timestamp 1649977179
transform 1 0 1789 0 1 18823
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_207
timestamp 1649977179
transform 1 0 1789 0 1 17143
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_208
timestamp 1649977179
transform 1 0 14661 0 1 18188
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_209
timestamp 1649977179
transform 1 0 31109 0 1 13196
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_210
timestamp 1649977179
transform 1 0 28613 0 1 13196
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_211
timestamp 1649977179
transform 1 0 26754 0 1 13946
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_212
timestamp 1649977179
transform 1 0 26630 0 1 12532
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_213
timestamp 1649977179
transform 1 0 26506 0 1 15360
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_214
timestamp 1649977179
transform 1 0 33605 0 1 13196
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_215
timestamp 1649977179
transform 1 0 22803 0 1 18188
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_216
timestamp 1649977179
transform 1 0 17245 0 1 1687
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_217
timestamp 1649977179
transform 1 0 1789 0 1 22183
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_218
timestamp 1649977179
transform 1 0 2536 0 1 25296
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_219
timestamp 1649977179
transform 1 0 1789 0 1 25543
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_220
timestamp 1649977179
transform 1 0 1789 0 1 23863
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_221
timestamp 1649977179
transform 1 0 1789 0 1 28903
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_222
timestamp 1649977179
transform 1 0 1789 0 1 27223
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_223
timestamp 1649977179
transform 1 0 1789 0 1 30583
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_224
timestamp 1649977179
transform 1 0 13663 0 1 31101
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_225
timestamp 1649977179
transform 1 0 14608 0 1 29902
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_226
timestamp 1649977179
transform 1 0 14862 0 1 28344
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_227
timestamp 1649977179
transform 1 0 13663 0 1 29973
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_228
timestamp 1649977179
transform 1 0 13663 0 1 28273
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_229
timestamp 1649977179
transform 1 0 14608 0 1 28344
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_230
timestamp 1649977179
transform 1 0 15022 0 1 31172
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_231
timestamp 1649977179
transform 1 0 14608 0 1 31172
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_232
timestamp 1649977179
transform 1 0 14942 0 1 29902
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_233
timestamp 1649977179
transform 1 0 13663 0 1 35629
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_234
timestamp 1649977179
transform 1 0 14608 0 1 35558
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_235
timestamp 1649977179
transform 1 0 14608 0 1 32730
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_236
timestamp 1649977179
transform 1 0 15182 0 1 34000
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_237
timestamp 1649977179
transform 1 0 15262 0 1 35558
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_238
timestamp 1649977179
transform 1 0 14608 0 1 34000
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_239
timestamp 1649977179
transform 1 0 15102 0 1 32730
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_240
timestamp 1649977179
transform 1 0 13663 0 1 33929
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_241
timestamp 1649977179
transform 1 0 13663 0 1 32801
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_242
timestamp 1649977179
transform 1 0 1789 0 1 32263
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_243
timestamp 1649977179
transform 1 0 1789 0 1 35623
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_244
timestamp 1649977179
transform 1 0 1789 0 1 33943
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_245
timestamp 1649977179
transform 1 0 1789 0 1 40663
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_246
timestamp 1649977179
transform 1 0 1789 0 1 38983
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_247
timestamp 1649977179
transform 1 0 1789 0 1 37303
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_248
timestamp 1649977179
transform 1 0 15342 0 1 36828
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_249
timestamp 1649977179
transform 1 0 14608 0 1 36828
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_250
timestamp 1649977179
transform 1 0 13663 0 1 36757
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_251
timestamp 1649977179
transform 1 0 1789 0 1 45703
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_252
timestamp 1649977179
transform 1 0 1789 0 1 44023
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_253
timestamp 1649977179
transform 1 0 1789 0 1 42343
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_254
timestamp 1649977179
transform 1 0 1789 0 1 47383
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_255
timestamp 1649977179
transform 1 0 1789 0 1 49063
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_256
timestamp 1649977179
transform 1 0 1789 0 1 50743
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_257
timestamp 1649977179
transform 1 0 1789 0 1 52423
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_258
timestamp 1649977179
transform 1 0 1789 0 1 55783
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_259
timestamp 1649977179
transform 1 0 1789 0 1 54103
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_260
timestamp 1649977179
transform 1 0 1789 0 1 60823
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_261
timestamp 1649977179
transform 1 0 1789 0 1 59143
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_262
timestamp 1649977179
transform 1 0 1789 0 1 57463
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_263
timestamp 1649977179
transform 1 0 1789 0 1 62503
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_264
timestamp 1649977179
transform 1 0 1789 0 1 65863
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_265
timestamp 1649977179
transform 1 0 1789 0 1 64183
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_266
timestamp 1649977179
transform 1 0 1789 0 1 67543
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_267
timestamp 1649977179
transform 1 0 1789 0 1 69223
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_268
timestamp 1649977179
transform 1 0 1789 0 1 72583
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_269
timestamp 1649977179
transform 1 0 1789 0 1 70903
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_270
timestamp 1649977179
transform 1 0 1789 0 1 77623
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_271
timestamp 1649977179
transform 1 0 1789 0 1 75943
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_272
timestamp 1649977179
transform 1 0 1789 0 1 74263
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_273
timestamp 1649977179
transform 1 0 1789 0 1 79303
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_274
timestamp 1649977179
transform 1 0 2125 0 1 81436
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_275
timestamp 1649977179
transform 1 0 1789 0 1 80983
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_276
timestamp 1649977179
transform 1 0 3805 0 1 81436
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_277
timestamp 1649977179
transform 1 0 7165 0 1 81436
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_278
timestamp 1649977179
transform 1 0 5485 0 1 81436
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_279
timestamp 1649977179
transform 1 0 15565 0 1 81436
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_280
timestamp 1649977179
transform 1 0 13885 0 1 81436
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_281
timestamp 1649977179
transform 1 0 12205 0 1 81436
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_282
timestamp 1649977179
transform 1 0 10525 0 1 81436
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_283
timestamp 1649977179
transform 1 0 8845 0 1 81436
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_284
timestamp 1649977179
transform 1 0 31109 0 1 76982
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_285
timestamp 1649977179
transform 1 0 28613 0 1 76982
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_286
timestamp 1649977179
transform 1 0 33605 0 1 76982
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_287
timestamp 1649977179
transform 1 0 23965 0 1 81436
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_288
timestamp 1649977179
transform 1 0 22285 0 1 81436
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_289
timestamp 1649977179
transform 1 0 20605 0 1 81436
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_290
timestamp 1649977179
transform 1 0 18925 0 1 81436
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_291
timestamp 1649977179
transform 1 0 25645 0 1 81436
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_292
timestamp 1649977179
transform 1 0 34045 0 1 81436
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_293
timestamp 1649977179
transform 1 0 32365 0 1 81436
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_294
timestamp 1649977179
transform 1 0 30685 0 1 81436
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_295
timestamp 1649977179
transform 1 0 29005 0 1 81436
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_296
timestamp 1649977179
transform 1 0 27325 0 1 81436
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_297
timestamp 1649977179
transform 1 0 17245 0 1 81436
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_298
timestamp 1649977179
transform 1 0 51077 0 1 76982
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_299
timestamp 1649977179
transform 1 0 48581 0 1 76982
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_300
timestamp 1649977179
transform 1 0 46085 0 1 76982
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_301
timestamp 1649977179
transform 1 0 43589 0 1 76982
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_302
timestamp 1649977179
transform 1 0 41093 0 1 76982
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_303
timestamp 1649977179
transform 1 0 38597 0 1 76982
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_304
timestamp 1649977179
transform 1 0 36101 0 1 76982
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_305
timestamp 1649977179
transform 1 0 35725 0 1 81436
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_306
timestamp 1649977179
transform 1 0 42445 0 1 81436
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_307
timestamp 1649977179
transform 1 0 40765 0 1 81436
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_308
timestamp 1649977179
transform 1 0 39085 0 1 81436
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_309
timestamp 1649977179
transform 1 0 37405 0 1 81436
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_310
timestamp 1649977179
transform 1 0 45805 0 1 81436
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_311
timestamp 1649977179
transform 1 0 44125 0 1 81436
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_312
timestamp 1649977179
transform 1 0 50845 0 1 81436
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_313
timestamp 1649977179
transform 1 0 49165 0 1 81436
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_314
timestamp 1649977179
transform 1 0 47485 0 1 81436
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_315
timestamp 1649977179
transform 1 0 66053 0 1 76982
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_316
timestamp 1649977179
transform 1 0 63557 0 1 76982
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_317
timestamp 1649977179
transform 1 0 61061 0 1 76982
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_318
timestamp 1649977179
transform 1 0 58565 0 1 76982
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_319
timestamp 1649977179
transform 1 0 56069 0 1 76982
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_320
timestamp 1649977179
transform 1 0 53573 0 1 76982
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_321
timestamp 1649977179
transform 1 0 57565 0 1 81436
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_322
timestamp 1649977179
transform 1 0 55885 0 1 81436
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_323
timestamp 1649977179
transform 1 0 54205 0 1 81436
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_324
timestamp 1649977179
transform 1 0 52525 0 1 81436
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_325
timestamp 1649977179
transform 1 0 59245 0 1 81436
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_326
timestamp 1649977179
transform 1 0 67645 0 1 81436
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_327
timestamp 1649977179
transform 1 0 65965 0 1 81436
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_328
timestamp 1649977179
transform 1 0 64285 0 1 81436
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_329
timestamp 1649977179
transform 1 0 62605 0 1 81436
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_330
timestamp 1649977179
transform 1 0 60925 0 1 81436
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_331
timestamp 1649977179
transform 1 0 134839 0 1 42343
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_332
timestamp 1649977179
transform 1 0 134839 0 1 45703
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_333
timestamp 1649977179
transform 1 0 134839 0 1 44023
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_334
timestamp 1649977179
transform 1 0 134839 0 1 47383
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_335
timestamp 1649977179
transform 1 0 134839 0 1 49063
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_336
timestamp 1649977179
transform 1 0 134839 0 1 50743
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_337
timestamp 1649977179
transform 1 0 134839 0 1 55783
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_338
timestamp 1649977179
transform 1 0 134839 0 1 54103
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_339
timestamp 1649977179
transform 1 0 134839 0 1 52423
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_340
timestamp 1649977179
transform 1 0 134092 0 1 62054
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_341
timestamp 1649977179
transform 1 0 134839 0 1 60823
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_342
timestamp 1649977179
transform 1 0 134839 0 1 59143
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_343
timestamp 1649977179
transform 1 0 134839 0 1 57463
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_344
timestamp 1649977179
transform 1 0 78533 0 1 76982
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_345
timestamp 1649977179
transform 1 0 83525 0 1 76982
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_346
timestamp 1649977179
transform 1 0 81029 0 1 76982
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_347
timestamp 1649977179
transform 1 0 71045 0 1 76982
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_348
timestamp 1649977179
transform 1 0 68549 0 1 76982
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_349
timestamp 1649977179
transform 1 0 76037 0 1 76982
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_350
timestamp 1649977179
transform 1 0 73541 0 1 76982
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_351
timestamp 1649977179
transform 1 0 76045 0 1 81436
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_352
timestamp 1649977179
transform 1 0 74365 0 1 81436
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_353
timestamp 1649977179
transform 1 0 72685 0 1 81436
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_354
timestamp 1649977179
transform 1 0 71005 0 1 81436
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_355
timestamp 1649977179
transform 1 0 69325 0 1 81436
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_356
timestamp 1649977179
transform 1 0 84445 0 1 81436
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_357
timestamp 1649977179
transform 1 0 82765 0 1 81436
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_358
timestamp 1649977179
transform 1 0 81085 0 1 81436
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_359
timestamp 1649977179
transform 1 0 79405 0 1 81436
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_360
timestamp 1649977179
transform 1 0 77725 0 1 81436
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_361
timestamp 1649977179
transform 1 0 96005 0 1 76982
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_362
timestamp 1649977179
transform 1 0 100997 0 1 76982
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_363
timestamp 1649977179
transform 1 0 98501 0 1 76982
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_364
timestamp 1649977179
transform 1 0 93509 0 1 76982
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_365
timestamp 1649977179
transform 1 0 91013 0 1 76982
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_366
timestamp 1649977179
transform 1 0 88517 0 1 76982
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_367
timestamp 1649977179
transform 1 0 86021 0 1 76982
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_368
timestamp 1649977179
transform 1 0 86125 0 1 81436
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_369
timestamp 1649977179
transform 1 0 92845 0 1 81436
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_370
timestamp 1649977179
transform 1 0 91165 0 1 81436
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_371
timestamp 1649977179
transform 1 0 89485 0 1 81436
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_372
timestamp 1649977179
transform 1 0 87805 0 1 81436
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_373
timestamp 1649977179
transform 1 0 101245 0 1 81436
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_374
timestamp 1649977179
transform 1 0 99565 0 1 81436
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_375
timestamp 1649977179
transform 1 0 97885 0 1 81436
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_376
timestamp 1649977179
transform 1 0 96205 0 1 81436
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_377
timestamp 1649977179
transform 1 0 94525 0 1 81436
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_378
timestamp 1649977179
transform 1 0 134839 0 1 62503
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_379
timestamp 1649977179
transform 1 0 134839 0 1 65863
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_380
timestamp 1649977179
transform 1 0 134839 0 1 64183
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_381
timestamp 1649977179
transform 1 0 122267 0 1 71990
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_382
timestamp 1649977179
transform 1 0 134839 0 1 67543
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_383
timestamp 1649977179
transform 1 0 134839 0 1 72583
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_384
timestamp 1649977179
transform 1 0 134839 0 1 70903
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_385
timestamp 1649977179
transform 1 0 134839 0 1 69223
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_386
timestamp 1649977179
transform 1 0 114041 0 1 71990
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_387
timestamp 1649977179
transform 1 0 105989 0 1 76982
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_388
timestamp 1649977179
transform 1 0 103493 0 1 76982
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_389
timestamp 1649977179
transform 1 0 110056 0 1 74818
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_390
timestamp 1649977179
transform 1 0 110180 0 1 73404
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_391
timestamp 1649977179
transform 1 0 104605 0 1 81436
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_392
timestamp 1649977179
transform 1 0 102925 0 1 81436
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_393
timestamp 1649977179
transform 1 0 109645 0 1 81436
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_394
timestamp 1649977179
transform 1 0 107965 0 1 81436
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_395
timestamp 1649977179
transform 1 0 106285 0 1 81436
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_396
timestamp 1649977179
transform 1 0 118593 0 1 80200
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_397
timestamp 1649977179
transform 1 0 118045 0 1 81436
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_398
timestamp 1649977179
transform 1 0 116365 0 1 81436
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_399
timestamp 1649977179
transform 1 0 114685 0 1 81436
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_400
timestamp 1649977179
transform 1 0 113005 0 1 81436
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_401
timestamp 1649977179
transform 1 0 111325 0 1 81436
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_402
timestamp 1649977179
transform 1 0 134839 0 1 75943
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_403
timestamp 1649977179
transform 1 0 134839 0 1 74263
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_404
timestamp 1649977179
transform 1 0 134839 0 1 77623
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_405
timestamp 1649977179
transform 1 0 122267 0 1 74818
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_406
timestamp 1649977179
transform 1 0 122267 0 1 73404
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_407
timestamp 1649977179
transform 1 0 124765 0 1 81436
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_408
timestamp 1649977179
transform 1 0 123085 0 1 81436
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_409
timestamp 1649977179
transform 1 0 121405 0 1 81436
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_410
timestamp 1649977179
transform 1 0 119725 0 1 81436
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_411
timestamp 1649977179
transform 1 0 119761 0 1 80200
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_412
timestamp 1649977179
transform 1 0 126445 0 1 81436
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_413
timestamp 1649977179
transform 1 0 133879 0 1 79203
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_414
timestamp 1649977179
transform 1 0 134839 0 1 79303
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_415
timestamp 1649977179
transform 1 0 130742 0 1 79098
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_416
timestamp 1649977179
transform 1 0 128125 0 1 81436
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_417
timestamp 1649977179
transform 1 0 131485 0 1 81436
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_418
timestamp 1649977179
transform 1 0 129805 0 1 81436
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_419
timestamp 1649977179
transform 1 0 134839 0 1 80983
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_420
timestamp 1649977179
transform 1 0 133165 0 1 81436
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_0
timestamp 1649977179
transform 1 0 134847 0 1 2691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1
timestamp 1649977179
transform 1 0 132837 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_2
timestamp 1649977179
transform 1 0 134847 0 1 2355
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_3
timestamp 1649977179
transform 1 0 132501 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_4
timestamp 1649977179
transform 1 0 132165 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_5
timestamp 1649977179
transform 1 0 134181 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_6
timestamp 1649977179
transform 1 0 133845 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_7
timestamp 1649977179
transform 1 0 134847 0 1 2019
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_8
timestamp 1649977179
transform 1 0 133509 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_9
timestamp 1649977179
transform 1 0 133173 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_10
timestamp 1649977179
transform 1 0 128133 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_11
timestamp 1649977179
transform 1 0 131829 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_12
timestamp 1649977179
transform 1 0 131493 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_13
timestamp 1649977179
transform 1 0 131157 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_14
timestamp 1649977179
transform 1 0 130821 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_15
timestamp 1649977179
transform 1 0 130485 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_16
timestamp 1649977179
transform 1 0 130149 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_17
timestamp 1649977179
transform 1 0 129813 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_18
timestamp 1649977179
transform 1 0 129477 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_19
timestamp 1649977179
transform 1 0 129141 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_20
timestamp 1649977179
transform 1 0 128805 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_21
timestamp 1649977179
transform 1 0 128469 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_22
timestamp 1649977179
transform 1 0 134847 0 1 3027
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_23
timestamp 1649977179
transform 1 0 134847 0 1 3363
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_24
timestamp 1649977179
transform 1 0 134847 0 1 4371
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_25
timestamp 1649977179
transform 1 0 134847 0 1 3699
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_26
timestamp 1649977179
transform 1 0 134847 0 1 4035
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_27
timestamp 1649977179
transform 1 0 134847 0 1 5043
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_28
timestamp 1649977179
transform 1 0 134847 0 1 4707
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_29
timestamp 1649977179
transform 1 0 126453 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_30
timestamp 1649977179
transform 1 0 126117 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_31
timestamp 1649977179
transform 1 0 125781 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_32
timestamp 1649977179
transform 1 0 125445 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_33
timestamp 1649977179
transform 1 0 125109 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_34
timestamp 1649977179
transform 1 0 124773 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_35
timestamp 1649977179
transform 1 0 124437 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_36
timestamp 1649977179
transform 1 0 124101 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_37
timestamp 1649977179
transform 1 0 123765 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_38
timestamp 1649977179
transform 1 0 123429 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_39
timestamp 1649977179
transform 1 0 123093 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_40
timestamp 1649977179
transform 1 0 122757 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_41
timestamp 1649977179
transform 1 0 122421 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_42
timestamp 1649977179
transform 1 0 122085 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_43
timestamp 1649977179
transform 1 0 121749 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_44
timestamp 1649977179
transform 1 0 121413 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_45
timestamp 1649977179
transform 1 0 121077 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_46
timestamp 1649977179
transform 1 0 120741 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_47
timestamp 1649977179
transform 1 0 120405 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_48
timestamp 1649977179
transform 1 0 120069 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_49
timestamp 1649977179
transform 1 0 119733 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_50
timestamp 1649977179
transform 1 0 127461 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_51
timestamp 1649977179
transform 1 0 127125 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_52
timestamp 1649977179
transform 1 0 126789 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_53
timestamp 1649977179
transform 1 0 134847 0 1 10419
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_54
timestamp 1649977179
transform 1 0 134847 0 1 10083
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_55
timestamp 1649977179
transform 1 0 134847 0 1 9747
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_56
timestamp 1649977179
transform 1 0 134847 0 1 9411
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_57
timestamp 1649977179
transform 1 0 134847 0 1 9075
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_58
timestamp 1649977179
transform 1 0 134847 0 1 8739
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_59
timestamp 1649977179
transform 1 0 134847 0 1 8403
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_60
timestamp 1649977179
transform 1 0 134847 0 1 8067
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_61
timestamp 1649977179
transform 1 0 134847 0 1 7731
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_62
timestamp 1649977179
transform 1 0 134847 0 1 7395
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_63
timestamp 1649977179
transform 1 0 134847 0 1 7059
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_64
timestamp 1649977179
transform 1 0 134847 0 1 6723
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_65
timestamp 1649977179
transform 1 0 134847 0 1 6387
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_66
timestamp 1649977179
transform 1 0 134847 0 1 6051
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_67
timestamp 1649977179
transform 1 0 134847 0 1 5715
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_68
timestamp 1649977179
transform 1 0 134847 0 1 5379
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_69
timestamp 1649977179
transform 1 0 127797 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_70
timestamp 1649977179
transform 1 0 117717 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_71
timestamp 1649977179
transform 1 0 115029 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_72
timestamp 1649977179
transform 1 0 111669 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_73
timestamp 1649977179
transform 1 0 114693 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_74
timestamp 1649977179
transform 1 0 114357 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_75
timestamp 1649977179
transform 1 0 115365 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_76
timestamp 1649977179
transform 1 0 111333 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_77
timestamp 1649977179
transform 1 0 117381 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_78
timestamp 1649977179
transform 1 0 114021 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_79
timestamp 1649977179
transform 1 0 119061 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_80
timestamp 1649977179
transform 1 0 110997 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_81
timestamp 1649977179
transform 1 0 118725 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_82
timestamp 1649977179
transform 1 0 115701 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_83
timestamp 1649977179
transform 1 0 113685 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_84
timestamp 1649977179
transform 1 0 117045 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_85
timestamp 1649977179
transform 1 0 116373 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_86
timestamp 1649977179
transform 1 0 118389 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_87
timestamp 1649977179
transform 1 0 116709 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_88
timestamp 1649977179
transform 1 0 113349 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_89
timestamp 1649977179
transform 1 0 113013 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_90
timestamp 1649977179
transform 1 0 116037 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_91
timestamp 1649977179
transform 1 0 112677 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_92
timestamp 1649977179
transform 1 0 112341 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_93
timestamp 1649977179
transform 1 0 118053 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_94
timestamp 1649977179
transform 1 0 112005 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_95
timestamp 1649977179
transform 1 0 108981 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_96
timestamp 1649977179
transform 1 0 108645 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_97
timestamp 1649977179
transform 1 0 107637 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_98
timestamp 1649977179
transform 1 0 108309 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_99
timestamp 1649977179
transform 1 0 105957 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_100
timestamp 1649977179
transform 1 0 105621 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_101
timestamp 1649977179
transform 1 0 104277 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_102
timestamp 1649977179
transform 1 0 103941 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_103
timestamp 1649977179
transform 1 0 103605 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_104
timestamp 1649977179
transform 1 0 103269 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_105
timestamp 1649977179
transform 1 0 102933 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_106
timestamp 1649977179
transform 1 0 102597 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_107
timestamp 1649977179
transform 1 0 105285 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_108
timestamp 1649977179
transform 1 0 107301 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_109
timestamp 1649977179
transform 1 0 104949 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_110
timestamp 1649977179
transform 1 0 106965 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_111
timestamp 1649977179
transform 1 0 106629 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_112
timestamp 1649977179
transform 1 0 110661 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_113
timestamp 1649977179
transform 1 0 110325 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_114
timestamp 1649977179
transform 1 0 107973 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_115
timestamp 1649977179
transform 1 0 109989 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_116
timestamp 1649977179
transform 1 0 104613 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_117
timestamp 1649977179
transform 1 0 106293 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_118
timestamp 1649977179
transform 1 0 109653 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_119
timestamp 1649977179
transform 1 0 109317 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_120
timestamp 1649977179
transform 1 0 134847 0 1 15123
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_121
timestamp 1649977179
transform 1 0 134847 0 1 14787
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_122
timestamp 1649977179
transform 1 0 134847 0 1 14451
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_123
timestamp 1649977179
transform 1 0 134847 0 1 14115
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_124
timestamp 1649977179
transform 1 0 134847 0 1 13779
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_125
timestamp 1649977179
transform 1 0 134847 0 1 13443
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_126
timestamp 1649977179
transform 1 0 134847 0 1 13107
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_127
timestamp 1649977179
transform 1 0 134847 0 1 12771
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_128
timestamp 1649977179
transform 1 0 134847 0 1 12435
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_129
timestamp 1649977179
transform 1 0 134847 0 1 12099
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_130
timestamp 1649977179
transform 1 0 134847 0 1 11763
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_131
timestamp 1649977179
transform 1 0 134847 0 1 11427
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_132
timestamp 1649977179
transform 1 0 134847 0 1 11091
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_133
timestamp 1649977179
transform 1 0 134847 0 1 10755
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_134
timestamp 1649977179
transform 1 0 134847 0 1 15459
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_135
timestamp 1649977179
transform 1 0 134847 0 1 20835
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_136
timestamp 1649977179
transform 1 0 134847 0 1 20499
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_137
timestamp 1649977179
transform 1 0 134847 0 1 20163
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_138
timestamp 1649977179
transform 1 0 134847 0 1 19827
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_139
timestamp 1649977179
transform 1 0 134847 0 1 19491
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_140
timestamp 1649977179
transform 1 0 134847 0 1 19155
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_141
timestamp 1649977179
transform 1 0 134847 0 1 18819
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_142
timestamp 1649977179
transform 1 0 134847 0 1 18483
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_143
timestamp 1649977179
transform 1 0 134847 0 1 18147
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_144
timestamp 1649977179
transform 1 0 134847 0 1 17811
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_145
timestamp 1649977179
transform 1 0 134847 0 1 17475
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_146
timestamp 1649977179
transform 1 0 134847 0 1 17139
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_147
timestamp 1649977179
transform 1 0 134847 0 1 16803
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_148
timestamp 1649977179
transform 1 0 134847 0 1 16467
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_149
timestamp 1649977179
transform 1 0 134847 0 1 16131
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_150
timestamp 1649977179
transform 1 0 134847 0 1 15795
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_151
timestamp 1649977179
transform 1 0 119397 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_152
timestamp 1649977179
transform 1 0 97893 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_153
timestamp 1649977179
transform 1 0 97557 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_154
timestamp 1649977179
transform 1 0 97221 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_155
timestamp 1649977179
transform 1 0 94533 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_156
timestamp 1649977179
transform 1 0 101925 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_157
timestamp 1649977179
transform 1 0 96885 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_158
timestamp 1649977179
transform 1 0 96549 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_159
timestamp 1649977179
transform 1 0 101589 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_160
timestamp 1649977179
transform 1 0 94197 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_161
timestamp 1649977179
transform 1 0 101253 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_162
timestamp 1649977179
transform 1 0 100917 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_163
timestamp 1649977179
transform 1 0 99237 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_164
timestamp 1649977179
transform 1 0 100581 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_165
timestamp 1649977179
transform 1 0 96213 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_166
timestamp 1649977179
transform 1 0 100245 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_167
timestamp 1649977179
transform 1 0 95877 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_168
timestamp 1649977179
transform 1 0 95205 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_169
timestamp 1649977179
transform 1 0 95541 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_170
timestamp 1649977179
transform 1 0 98901 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_171
timestamp 1649977179
transform 1 0 98565 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_172
timestamp 1649977179
transform 1 0 98229 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_173
timestamp 1649977179
transform 1 0 94869 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_174
timestamp 1649977179
transform 1 0 99573 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_175
timestamp 1649977179
transform 1 0 99909 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_176
timestamp 1649977179
transform 1 0 92517 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_177
timestamp 1649977179
transform 1 0 86469 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_178
timestamp 1649977179
transform 1 0 86133 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_179
timestamp 1649977179
transform 1 0 85797 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_180
timestamp 1649977179
transform 1 0 85461 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_181
timestamp 1649977179
transform 1 0 92181 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_182
timestamp 1649977179
transform 1 0 92853 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_183
timestamp 1649977179
transform 1 0 93189 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_184
timestamp 1649977179
transform 1 0 89829 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_185
timestamp 1649977179
transform 1 0 91845 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_186
timestamp 1649977179
transform 1 0 89493 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_187
timestamp 1649977179
transform 1 0 89157 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_188
timestamp 1649977179
transform 1 0 88821 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_189
timestamp 1649977179
transform 1 0 91509 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_190
timestamp 1649977179
transform 1 0 88485 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_191
timestamp 1649977179
transform 1 0 91173 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_192
timestamp 1649977179
transform 1 0 88149 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_193
timestamp 1649977179
transform 1 0 93525 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_194
timestamp 1649977179
transform 1 0 90837 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_195
timestamp 1649977179
transform 1 0 90501 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_196
timestamp 1649977179
transform 1 0 90165 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_197
timestamp 1649977179
transform 1 0 87813 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_198
timestamp 1649977179
transform 1 0 87477 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_199
timestamp 1649977179
transform 1 0 87141 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_200
timestamp 1649977179
transform 1 0 86805 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_201
timestamp 1649977179
transform 1 0 93861 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_202
timestamp 1649977179
transform 1 0 80421 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_203
timestamp 1649977179
transform 1 0 79413 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_204
timestamp 1649977179
transform 1 0 80085 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_205
timestamp 1649977179
transform 1 0 85125 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_206
timestamp 1649977179
transform 1 0 79077 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_207
timestamp 1649977179
transform 1 0 78405 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_208
timestamp 1649977179
transform 1 0 82437 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_209
timestamp 1649977179
transform 1 0 84789 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_210
timestamp 1649977179
transform 1 0 83109 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_211
timestamp 1649977179
transform 1 0 83445 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_212
timestamp 1649977179
transform 1 0 82101 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_213
timestamp 1649977179
transform 1 0 77733 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_214
timestamp 1649977179
transform 1 0 84453 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_215
timestamp 1649977179
transform 1 0 77397 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_216
timestamp 1649977179
transform 1 0 81765 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_217
timestamp 1649977179
transform 1 0 84117 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_218
timestamp 1649977179
transform 1 0 81429 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_219
timestamp 1649977179
transform 1 0 78069 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_220
timestamp 1649977179
transform 1 0 81093 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_221
timestamp 1649977179
transform 1 0 82773 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_222
timestamp 1649977179
transform 1 0 80757 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_223
timestamp 1649977179
transform 1 0 79749 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_224
timestamp 1649977179
transform 1 0 77061 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_225
timestamp 1649977179
transform 1 0 83781 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_226
timestamp 1649977179
transform 1 0 78741 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_227
timestamp 1649977179
transform 1 0 75381 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_228
timestamp 1649977179
transform 1 0 75045 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_229
timestamp 1649977179
transform 1 0 74709 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_230
timestamp 1649977179
transform 1 0 74373 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_231
timestamp 1649977179
transform 1 0 76053 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_232
timestamp 1649977179
transform 1 0 74037 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_233
timestamp 1649977179
transform 1 0 73701 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_234
timestamp 1649977179
transform 1 0 73365 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_235
timestamp 1649977179
transform 1 0 73029 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_236
timestamp 1649977179
transform 1 0 72693 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_237
timestamp 1649977179
transform 1 0 72357 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_238
timestamp 1649977179
transform 1 0 72021 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_239
timestamp 1649977179
transform 1 0 71685 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_240
timestamp 1649977179
transform 1 0 71349 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_241
timestamp 1649977179
transform 1 0 71013 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_242
timestamp 1649977179
transform 1 0 70677 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_243
timestamp 1649977179
transform 1 0 70341 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_244
timestamp 1649977179
transform 1 0 70005 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_245
timestamp 1649977179
transform 1 0 69669 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_246
timestamp 1649977179
transform 1 0 69333 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_247
timestamp 1649977179
transform 1 0 68997 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_248
timestamp 1649977179
transform 1 0 68661 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_249
timestamp 1649977179
transform 1 0 75717 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_250
timestamp 1649977179
transform 1 0 76389 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_251
timestamp 1649977179
transform 1 0 76725 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_252
timestamp 1649977179
transform 1 0 134847 0 1 21171
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_253
timestamp 1649977179
transform 1 0 134847 0 1 22515
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_254
timestamp 1649977179
transform 1 0 134847 0 1 24867
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_255
timestamp 1649977179
transform 1 0 134847 0 1 24531
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_256
timestamp 1649977179
transform 1 0 134847 0 1 24195
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_257
timestamp 1649977179
transform 1 0 134847 0 1 23859
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_258
timestamp 1649977179
transform 1 0 134847 0 1 23523
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_259
timestamp 1649977179
transform 1 0 134847 0 1 25875
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_260
timestamp 1649977179
transform 1 0 134847 0 1 25539
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_261
timestamp 1649977179
transform 1 0 134847 0 1 25203
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_262
timestamp 1649977179
transform 1 0 134847 0 1 22179
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_263
timestamp 1649977179
transform 1 0 134847 0 1 23187
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_264
timestamp 1649977179
transform 1 0 134847 0 1 21843
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_265
timestamp 1649977179
transform 1 0 134847 0 1 22851
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_266
timestamp 1649977179
transform 1 0 134847 0 1 21507
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_267
timestamp 1649977179
transform 1 0 134847 0 1 27219
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_268
timestamp 1649977179
transform 1 0 134847 0 1 26883
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_269
timestamp 1649977179
transform 1 0 134847 0 1 26547
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_270
timestamp 1649977179
transform 1 0 134847 0 1 26211
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_271
timestamp 1649977179
transform 1 0 134847 0 1 30915
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_272
timestamp 1649977179
transform 1 0 134847 0 1 30579
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_273
timestamp 1649977179
transform 1 0 134847 0 1 30243
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_274
timestamp 1649977179
transform 1 0 134847 0 1 29907
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_275
timestamp 1649977179
transform 1 0 134847 0 1 29571
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_276
timestamp 1649977179
transform 1 0 134847 0 1 29235
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_277
timestamp 1649977179
transform 1 0 134847 0 1 28899
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_278
timestamp 1649977179
transform 1 0 134847 0 1 28563
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_279
timestamp 1649977179
transform 1 0 134847 0 1 28227
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_280
timestamp 1649977179
transform 1 0 134847 0 1 27891
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_281
timestamp 1649977179
transform 1 0 134847 0 1 27555
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_282
timestamp 1649977179
transform 1 0 134847 0 1 36291
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_283
timestamp 1649977179
transform 1 0 134847 0 1 35955
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_284
timestamp 1649977179
transform 1 0 134847 0 1 35619
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_285
timestamp 1649977179
transform 1 0 134847 0 1 35283
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_286
timestamp 1649977179
transform 1 0 134847 0 1 34947
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_287
timestamp 1649977179
transform 1 0 134847 0 1 34611
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_288
timestamp 1649977179
transform 1 0 134847 0 1 34275
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_289
timestamp 1649977179
transform 1 0 134847 0 1 31587
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_290
timestamp 1649977179
transform 1 0 134847 0 1 33939
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_291
timestamp 1649977179
transform 1 0 134847 0 1 33603
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_292
timestamp 1649977179
transform 1 0 134847 0 1 33267
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_293
timestamp 1649977179
transform 1 0 134847 0 1 32931
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_294
timestamp 1649977179
transform 1 0 134847 0 1 32595
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_295
timestamp 1649977179
transform 1 0 134847 0 1 32259
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_296
timestamp 1649977179
transform 1 0 134847 0 1 31923
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_297
timestamp 1649977179
transform 1 0 134847 0 1 41331
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_298
timestamp 1649977179
transform 1 0 134847 0 1 40995
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_299
timestamp 1649977179
transform 1 0 134847 0 1 40659
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_300
timestamp 1649977179
transform 1 0 134847 0 1 40323
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_301
timestamp 1649977179
transform 1 0 134847 0 1 39987
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_302
timestamp 1649977179
transform 1 0 134847 0 1 39651
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_303
timestamp 1649977179
transform 1 0 134847 0 1 39315
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_304
timestamp 1649977179
transform 1 0 134847 0 1 38979
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_305
timestamp 1649977179
transform 1 0 134847 0 1 38643
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_306
timestamp 1649977179
transform 1 0 134847 0 1 38307
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_307
timestamp 1649977179
transform 1 0 134847 0 1 37971
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_308
timestamp 1649977179
transform 1 0 134847 0 1 37635
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_309
timestamp 1649977179
transform 1 0 134847 0 1 37299
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_310
timestamp 1649977179
transform 1 0 134847 0 1 36963
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_311
timestamp 1649977179
transform 1 0 134847 0 1 36627
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_312
timestamp 1649977179
transform 1 0 134847 0 1 31251
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_313
timestamp 1649977179
transform 1 0 102261 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_314
timestamp 1649977179
transform 1 0 60261 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_315
timestamp 1649977179
transform 1 0 63285 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_316
timestamp 1649977179
transform 1 0 60933 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_317
timestamp 1649977179
transform 1 0 62949 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_318
timestamp 1649977179
transform 1 0 61269 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_319
timestamp 1649977179
transform 1 0 65301 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_320
timestamp 1649977179
transform 1 0 64629 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_321
timestamp 1649977179
transform 1 0 62277 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_322
timestamp 1649977179
transform 1 0 60597 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_323
timestamp 1649977179
transform 1 0 63957 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_324
timestamp 1649977179
transform 1 0 63621 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_325
timestamp 1649977179
transform 1 0 62613 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_326
timestamp 1649977179
transform 1 0 67653 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_327
timestamp 1649977179
transform 1 0 59925 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_328
timestamp 1649977179
transform 1 0 67317 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_329
timestamp 1649977179
transform 1 0 61941 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_330
timestamp 1649977179
transform 1 0 64293 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_331
timestamp 1649977179
transform 1 0 65973 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_332
timestamp 1649977179
transform 1 0 67989 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_333
timestamp 1649977179
transform 1 0 66981 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_334
timestamp 1649977179
transform 1 0 66645 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_335
timestamp 1649977179
transform 1 0 65637 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_336
timestamp 1649977179
transform 1 0 66309 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_337
timestamp 1649977179
transform 1 0 64965 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_338
timestamp 1649977179
transform 1 0 61605 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_339
timestamp 1649977179
transform 1 0 57237 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_340
timestamp 1649977179
transform 1 0 56901 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_341
timestamp 1649977179
transform 1 0 56565 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_342
timestamp 1649977179
transform 1 0 56229 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_343
timestamp 1649977179
transform 1 0 55893 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_344
timestamp 1649977179
transform 1 0 58917 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_345
timestamp 1649977179
transform 1 0 55557 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_346
timestamp 1649977179
transform 1 0 55221 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_347
timestamp 1649977179
transform 1 0 58245 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_348
timestamp 1649977179
transform 1 0 54885 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_349
timestamp 1649977179
transform 1 0 54549 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_350
timestamp 1649977179
transform 1 0 54213 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_351
timestamp 1649977179
transform 1 0 53877 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_352
timestamp 1649977179
transform 1 0 53541 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_353
timestamp 1649977179
transform 1 0 53205 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_354
timestamp 1649977179
transform 1 0 52869 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_355
timestamp 1649977179
transform 1 0 52533 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_356
timestamp 1649977179
transform 1 0 52197 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_357
timestamp 1649977179
transform 1 0 51861 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_358
timestamp 1649977179
transform 1 0 51525 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_359
timestamp 1649977179
transform 1 0 57573 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_360
timestamp 1649977179
transform 1 0 59589 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_361
timestamp 1649977179
transform 1 0 57909 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_362
timestamp 1649977179
transform 1 0 58581 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_363
timestamp 1649977179
transform 1 0 59253 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_364
timestamp 1649977179
transform 1 0 47829 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_365
timestamp 1649977179
transform 1 0 44133 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_366
timestamp 1649977179
transform 1 0 47493 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_367
timestamp 1649977179
transform 1 0 47157 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_368
timestamp 1649977179
transform 1 0 46821 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_369
timestamp 1649977179
transform 1 0 46485 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_370
timestamp 1649977179
transform 1 0 43797 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_371
timestamp 1649977179
transform 1 0 43461 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_372
timestamp 1649977179
transform 1 0 46149 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_373
timestamp 1649977179
transform 1 0 51189 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_374
timestamp 1649977179
transform 1 0 45813 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_375
timestamp 1649977179
transform 1 0 45477 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_376
timestamp 1649977179
transform 1 0 43125 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_377
timestamp 1649977179
transform 1 0 45141 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_378
timestamp 1649977179
transform 1 0 50853 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_379
timestamp 1649977179
transform 1 0 50517 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_380
timestamp 1649977179
transform 1 0 50181 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_381
timestamp 1649977179
transform 1 0 49845 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_382
timestamp 1649977179
transform 1 0 44805 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_383
timestamp 1649977179
transform 1 0 44469 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_384
timestamp 1649977179
transform 1 0 49509 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_385
timestamp 1649977179
transform 1 0 49173 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_386
timestamp 1649977179
transform 1 0 48837 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_387
timestamp 1649977179
transform 1 0 48501 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_388
timestamp 1649977179
transform 1 0 48165 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_389
timestamp 1649977179
transform 1 0 39429 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_390
timestamp 1649977179
transform 1 0 39093 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_391
timestamp 1649977179
transform 1 0 38757 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_392
timestamp 1649977179
transform 1 0 38421 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_393
timestamp 1649977179
transform 1 0 38085 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_394
timestamp 1649977179
transform 1 0 37749 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_395
timestamp 1649977179
transform 1 0 37413 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_396
timestamp 1649977179
transform 1 0 37077 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_397
timestamp 1649977179
transform 1 0 36741 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_398
timestamp 1649977179
transform 1 0 36405 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_399
timestamp 1649977179
transform 1 0 36069 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_400
timestamp 1649977179
transform 1 0 35733 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_401
timestamp 1649977179
transform 1 0 34389 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_402
timestamp 1649977179
transform 1 0 35397 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_403
timestamp 1649977179
transform 1 0 35061 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_404
timestamp 1649977179
transform 1 0 34725 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_405
timestamp 1649977179
transform 1 0 39765 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_406
timestamp 1649977179
transform 1 0 42453 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_407
timestamp 1649977179
transform 1 0 42117 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_408
timestamp 1649977179
transform 1 0 41781 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_409
timestamp 1649977179
transform 1 0 41445 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_410
timestamp 1649977179
transform 1 0 41109 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_411
timestamp 1649977179
transform 1 0 40773 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_412
timestamp 1649977179
transform 1 0 40437 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_413
timestamp 1649977179
transform 1 0 40101 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_414
timestamp 1649977179
transform 1 0 42789 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_415
timestamp 1649977179
transform 1 0 28005 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_416
timestamp 1649977179
transform 1 0 27669 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_417
timestamp 1649977179
transform 1 0 29013 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_418
timestamp 1649977179
transform 1 0 33045 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_419
timestamp 1649977179
transform 1 0 32709 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_420
timestamp 1649977179
transform 1 0 28677 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_421
timestamp 1649977179
transform 1 0 32373 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_422
timestamp 1649977179
transform 1 0 32037 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_423
timestamp 1649977179
transform 1 0 27333 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_424
timestamp 1649977179
transform 1 0 26997 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_425
timestamp 1649977179
transform 1 0 28341 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_426
timestamp 1649977179
transform 1 0 31701 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_427
timestamp 1649977179
transform 1 0 26661 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_428
timestamp 1649977179
transform 1 0 31365 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_429
timestamp 1649977179
transform 1 0 26325 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_430
timestamp 1649977179
transform 1 0 31029 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_431
timestamp 1649977179
transform 1 0 30693 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_432
timestamp 1649977179
transform 1 0 25989 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_433
timestamp 1649977179
transform 1 0 30357 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_434
timestamp 1649977179
transform 1 0 30021 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_435
timestamp 1649977179
transform 1 0 29685 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_436
timestamp 1649977179
transform 1 0 34053 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_437
timestamp 1649977179
transform 1 0 29349 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_438
timestamp 1649977179
transform 1 0 33717 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_439
timestamp 1649977179
transform 1 0 33381 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_440
timestamp 1649977179
transform 1 0 18597 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_441
timestamp 1649977179
transform 1 0 18261 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_442
timestamp 1649977179
transform 1 0 20613 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_443
timestamp 1649977179
transform 1 0 20277 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_444
timestamp 1649977179
transform 1 0 19941 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_445
timestamp 1649977179
transform 1 0 25653 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_446
timestamp 1649977179
transform 1 0 25317 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_447
timestamp 1649977179
transform 1 0 24981 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_448
timestamp 1649977179
transform 1 0 24645 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_449
timestamp 1649977179
transform 1 0 24309 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_450
timestamp 1649977179
transform 1 0 23973 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_451
timestamp 1649977179
transform 1 0 23637 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_452
timestamp 1649977179
transform 1 0 23301 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_453
timestamp 1649977179
transform 1 0 22965 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_454
timestamp 1649977179
transform 1 0 19605 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_455
timestamp 1649977179
transform 1 0 22629 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_456
timestamp 1649977179
transform 1 0 19269 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_457
timestamp 1649977179
transform 1 0 22293 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_458
timestamp 1649977179
transform 1 0 17925 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_459
timestamp 1649977179
transform 1 0 21957 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_460
timestamp 1649977179
transform 1 0 21621 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_461
timestamp 1649977179
transform 1 0 21285 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_462
timestamp 1649977179
transform 1 0 17589 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_463
timestamp 1649977179
transform 1 0 20949 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_464
timestamp 1649977179
transform 1 0 18933 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_465
timestamp 1649977179
transform 1 0 9189 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_466
timestamp 1649977179
transform 1 0 8853 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_467
timestamp 1649977179
transform 1 0 13557 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_468
timestamp 1649977179
transform 1 0 10197 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_469
timestamp 1649977179
transform 1 0 9525 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_470
timestamp 1649977179
transform 1 0 13221 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_471
timestamp 1649977179
transform 1 0 12885 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_472
timestamp 1649977179
transform 1 0 12549 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_473
timestamp 1649977179
transform 1 0 12213 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_474
timestamp 1649977179
transform 1 0 9861 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_475
timestamp 1649977179
transform 1 0 11877 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_476
timestamp 1649977179
transform 1 0 11541 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_477
timestamp 1649977179
transform 1 0 11205 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_478
timestamp 1649977179
transform 1 0 10869 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_479
timestamp 1649977179
transform 1 0 16917 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_480
timestamp 1649977179
transform 1 0 16581 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_481
timestamp 1649977179
transform 1 0 16245 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_482
timestamp 1649977179
transform 1 0 10533 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_483
timestamp 1649977179
transform 1 0 15909 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_484
timestamp 1649977179
transform 1 0 15573 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_485
timestamp 1649977179
transform 1 0 15237 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_486
timestamp 1649977179
transform 1 0 14901 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_487
timestamp 1649977179
transform 1 0 14565 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_488
timestamp 1649977179
transform 1 0 14229 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_489
timestamp 1649977179
transform 1 0 13893 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_490
timestamp 1649977179
transform 1 0 4821 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_491
timestamp 1649977179
transform 1 0 5829 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_492
timestamp 1649977179
transform 1 0 5157 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_493
timestamp 1649977179
transform 1 0 6165 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_494
timestamp 1649977179
transform 1 0 7173 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_495
timestamp 1649977179
transform 1 0 6837 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_496
timestamp 1649977179
transform 1 0 6501 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_497
timestamp 1649977179
transform 1 0 7845 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_498
timestamp 1649977179
transform 1 0 8517 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_499
timestamp 1649977179
transform 1 0 5493 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_500
timestamp 1649977179
transform 1 0 7509 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_501
timestamp 1649977179
transform 1 0 8181 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_502
timestamp 1649977179
transform 1 0 4149 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_503
timestamp 1649977179
transform 1 0 3813 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_504
timestamp 1649977179
transform 1 0 3477 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_505
timestamp 1649977179
transform 1 0 3141 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_506
timestamp 1649977179
transform 1 0 2805 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_507
timestamp 1649977179
transform 1 0 2469 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_508
timestamp 1649977179
transform 1 0 2133 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_509
timestamp 1649977179
transform 1 0 1797 0 1 2691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_510
timestamp 1649977179
transform 1 0 1797 0 1 2355
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_511
timestamp 1649977179
transform 1 0 1797 0 1 2019
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_512
timestamp 1649977179
transform 1 0 1797 0 1 4371
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_513
timestamp 1649977179
transform 1 0 1797 0 1 4035
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_514
timestamp 1649977179
transform 1 0 1797 0 1 3699
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_515
timestamp 1649977179
transform 1 0 1797 0 1 3363
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_516
timestamp 1649977179
transform 1 0 1797 0 1 3027
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_517
timestamp 1649977179
transform 1 0 1797 0 1 5043
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_518
timestamp 1649977179
transform 1 0 1797 0 1 4707
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_519
timestamp 1649977179
transform 1 0 4485 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_520
timestamp 1649977179
transform 1 0 1797 0 1 10419
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_521
timestamp 1649977179
transform 1 0 1797 0 1 10083
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_522
timestamp 1649977179
transform 1 0 1797 0 1 9747
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_523
timestamp 1649977179
transform 1 0 1797 0 1 9411
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_524
timestamp 1649977179
transform 1 0 1797 0 1 9075
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_525
timestamp 1649977179
transform 1 0 1797 0 1 8739
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_526
timestamp 1649977179
transform 1 0 1797 0 1 8403
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_527
timestamp 1649977179
transform 1 0 1797 0 1 8067
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_528
timestamp 1649977179
transform 1 0 1797 0 1 7731
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_529
timestamp 1649977179
transform 1 0 1797 0 1 7395
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_530
timestamp 1649977179
transform 1 0 1797 0 1 7059
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_531
timestamp 1649977179
transform 1 0 1797 0 1 6723
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_532
timestamp 1649977179
transform 1 0 1797 0 1 6387
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_533
timestamp 1649977179
transform 1 0 1797 0 1 6051
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_534
timestamp 1649977179
transform 1 0 1797 0 1 5715
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_535
timestamp 1649977179
transform 1 0 1797 0 1 5379
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_536
timestamp 1649977179
transform 1 0 1797 0 1 13443
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_537
timestamp 1649977179
transform 1 0 1797 0 1 15459
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_538
timestamp 1649977179
transform 1 0 1797 0 1 15123
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_539
timestamp 1649977179
transform 1 0 1797 0 1 11427
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_540
timestamp 1649977179
transform 1 0 1797 0 1 11091
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_541
timestamp 1649977179
transform 1 0 1797 0 1 14787
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_542
timestamp 1649977179
transform 1 0 1797 0 1 10755
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_543
timestamp 1649977179
transform 1 0 1797 0 1 13107
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_544
timestamp 1649977179
transform 1 0 1797 0 1 14451
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_545
timestamp 1649977179
transform 1 0 1797 0 1 12771
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_546
timestamp 1649977179
transform 1 0 1797 0 1 12435
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_547
timestamp 1649977179
transform 1 0 1797 0 1 14115
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_548
timestamp 1649977179
transform 1 0 1797 0 1 12099
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_549
timestamp 1649977179
transform 1 0 1797 0 1 11763
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_550
timestamp 1649977179
transform 1 0 1797 0 1 13779
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_551
timestamp 1649977179
transform 1 0 1797 0 1 16131
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_552
timestamp 1649977179
transform 1 0 1797 0 1 17139
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_553
timestamp 1649977179
transform 1 0 1797 0 1 16803
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_554
timestamp 1649977179
transform 1 0 1797 0 1 16467
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_555
timestamp 1649977179
transform 1 0 1797 0 1 20835
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_556
timestamp 1649977179
transform 1 0 1797 0 1 20499
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_557
timestamp 1649977179
transform 1 0 1797 0 1 20163
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_558
timestamp 1649977179
transform 1 0 1797 0 1 19827
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_559
timestamp 1649977179
transform 1 0 1797 0 1 19491
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_560
timestamp 1649977179
transform 1 0 1797 0 1 19155
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_561
timestamp 1649977179
transform 1 0 1797 0 1 18819
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_562
timestamp 1649977179
transform 1 0 1797 0 1 18483
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_563
timestamp 1649977179
transform 1 0 1797 0 1 18147
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_564
timestamp 1649977179
transform 1 0 1797 0 1 17811
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_565
timestamp 1649977179
transform 1 0 1797 0 1 17475
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_566
timestamp 1649977179
transform 1 0 1797 0 1 15795
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_567
timestamp 1649977179
transform 1 0 17253 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_568
timestamp 1649977179
transform 1 0 1797 0 1 24195
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_569
timestamp 1649977179
transform 1 0 1797 0 1 21507
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_570
timestamp 1649977179
transform 1 0 1797 0 1 21171
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_571
timestamp 1649977179
transform 1 0 1797 0 1 24867
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_572
timestamp 1649977179
transform 1 0 1797 0 1 25203
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_573
timestamp 1649977179
transform 1 0 1797 0 1 22515
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_574
timestamp 1649977179
transform 1 0 1797 0 1 24531
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_575
timestamp 1649977179
transform 1 0 1797 0 1 25875
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_576
timestamp 1649977179
transform 1 0 1797 0 1 25539
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_577
timestamp 1649977179
transform 1 0 1797 0 1 22179
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_578
timestamp 1649977179
transform 1 0 1797 0 1 23859
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_579
timestamp 1649977179
transform 1 0 1797 0 1 23523
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_580
timestamp 1649977179
transform 1 0 1797 0 1 21843
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_581
timestamp 1649977179
transform 1 0 1797 0 1 23187
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_582
timestamp 1649977179
transform 1 0 1797 0 1 22851
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_583
timestamp 1649977179
transform 1 0 1797 0 1 26211
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_584
timestamp 1649977179
transform 1 0 1797 0 1 29907
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_585
timestamp 1649977179
transform 1 0 1797 0 1 30579
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_586
timestamp 1649977179
transform 1 0 1797 0 1 29571
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_587
timestamp 1649977179
transform 1 0 1797 0 1 29235
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_588
timestamp 1649977179
transform 1 0 1797 0 1 28899
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_589
timestamp 1649977179
transform 1 0 1797 0 1 28563
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_590
timestamp 1649977179
transform 1 0 1797 0 1 30243
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_591
timestamp 1649977179
transform 1 0 1797 0 1 28227
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_592
timestamp 1649977179
transform 1 0 1797 0 1 27891
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_593
timestamp 1649977179
transform 1 0 1797 0 1 30915
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_594
timestamp 1649977179
transform 1 0 1797 0 1 27555
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_595
timestamp 1649977179
transform 1 0 1797 0 1 27219
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_596
timestamp 1649977179
transform 1 0 1797 0 1 26883
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_597
timestamp 1649977179
transform 1 0 1797 0 1 26547
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_598
timestamp 1649977179
transform 1 0 1797 0 1 31923
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_599
timestamp 1649977179
transform 1 0 1797 0 1 36291
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_600
timestamp 1649977179
transform 1 0 1797 0 1 35955
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_601
timestamp 1649977179
transform 1 0 1797 0 1 35619
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_602
timestamp 1649977179
transform 1 0 1797 0 1 35283
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_603
timestamp 1649977179
transform 1 0 1797 0 1 31587
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_604
timestamp 1649977179
transform 1 0 1797 0 1 34947
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_605
timestamp 1649977179
transform 1 0 1797 0 1 34611
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_606
timestamp 1649977179
transform 1 0 1797 0 1 34275
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_607
timestamp 1649977179
transform 1 0 1797 0 1 33939
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_608
timestamp 1649977179
transform 1 0 1797 0 1 33603
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_609
timestamp 1649977179
transform 1 0 1797 0 1 33267
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_610
timestamp 1649977179
transform 1 0 1797 0 1 32931
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_611
timestamp 1649977179
transform 1 0 1797 0 1 32595
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_612
timestamp 1649977179
transform 1 0 1797 0 1 32259
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_613
timestamp 1649977179
transform 1 0 1797 0 1 36963
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_614
timestamp 1649977179
transform 1 0 1797 0 1 36627
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_615
timestamp 1649977179
transform 1 0 1797 0 1 37299
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_616
timestamp 1649977179
transform 1 0 1797 0 1 41331
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_617
timestamp 1649977179
transform 1 0 1797 0 1 40995
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_618
timestamp 1649977179
transform 1 0 1797 0 1 40659
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_619
timestamp 1649977179
transform 1 0 1797 0 1 40323
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_620
timestamp 1649977179
transform 1 0 1797 0 1 39987
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_621
timestamp 1649977179
transform 1 0 1797 0 1 39651
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_622
timestamp 1649977179
transform 1 0 1797 0 1 39315
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_623
timestamp 1649977179
transform 1 0 1797 0 1 38979
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_624
timestamp 1649977179
transform 1 0 1797 0 1 38643
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_625
timestamp 1649977179
transform 1 0 1797 0 1 38307
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_626
timestamp 1649977179
transform 1 0 1797 0 1 37971
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_627
timestamp 1649977179
transform 1 0 1797 0 1 37635
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_628
timestamp 1649977179
transform 1 0 1797 0 1 31251
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_629
timestamp 1649977179
transform 1 0 1797 0 1 45699
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_630
timestamp 1649977179
transform 1 0 1797 0 1 45363
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_631
timestamp 1649977179
transform 1 0 1797 0 1 45027
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_632
timestamp 1649977179
transform 1 0 1797 0 1 44691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_633
timestamp 1649977179
transform 1 0 1797 0 1 44355
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_634
timestamp 1649977179
transform 1 0 1797 0 1 44019
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_635
timestamp 1649977179
transform 1 0 1797 0 1 43683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_636
timestamp 1649977179
transform 1 0 1797 0 1 43347
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_637
timestamp 1649977179
transform 1 0 1797 0 1 43011
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_638
timestamp 1649977179
transform 1 0 1797 0 1 42675
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_639
timestamp 1649977179
transform 1 0 1797 0 1 42339
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_640
timestamp 1649977179
transform 1 0 1797 0 1 46371
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_641
timestamp 1649977179
transform 1 0 1797 0 1 46035
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_642
timestamp 1649977179
transform 1 0 1797 0 1 42003
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_643
timestamp 1649977179
transform 1 0 1797 0 1 48723
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_644
timestamp 1649977179
transform 1 0 1797 0 1 48387
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_645
timestamp 1649977179
transform 1 0 1797 0 1 48051
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_646
timestamp 1649977179
transform 1 0 1797 0 1 49059
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_647
timestamp 1649977179
transform 1 0 1797 0 1 50403
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_648
timestamp 1649977179
transform 1 0 1797 0 1 49731
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_649
timestamp 1649977179
transform 1 0 1797 0 1 47715
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_650
timestamp 1649977179
transform 1 0 1797 0 1 49395
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_651
timestamp 1649977179
transform 1 0 1797 0 1 51747
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_652
timestamp 1649977179
transform 1 0 1797 0 1 51411
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_653
timestamp 1649977179
transform 1 0 1797 0 1 47379
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_654
timestamp 1649977179
transform 1 0 1797 0 1 47043
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_655
timestamp 1649977179
transform 1 0 1797 0 1 51075
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_656
timestamp 1649977179
transform 1 0 1797 0 1 50739
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_657
timestamp 1649977179
transform 1 0 1797 0 1 50067
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_658
timestamp 1649977179
transform 1 0 1797 0 1 46707
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_659
timestamp 1649977179
transform 1 0 1797 0 1 54099
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_660
timestamp 1649977179
transform 1 0 1797 0 1 53763
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_661
timestamp 1649977179
transform 1 0 1797 0 1 53427
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_662
timestamp 1649977179
transform 1 0 1797 0 1 53091
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_663
timestamp 1649977179
transform 1 0 1797 0 1 52755
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_664
timestamp 1649977179
transform 1 0 1797 0 1 52083
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_665
timestamp 1649977179
transform 1 0 1797 0 1 52419
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_666
timestamp 1649977179
transform 1 0 1797 0 1 56451
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_667
timestamp 1649977179
transform 1 0 1797 0 1 56115
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_668
timestamp 1649977179
transform 1 0 1797 0 1 55779
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_669
timestamp 1649977179
transform 1 0 1797 0 1 55443
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_670
timestamp 1649977179
transform 1 0 1797 0 1 55107
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_671
timestamp 1649977179
transform 1 0 1797 0 1 54771
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_672
timestamp 1649977179
transform 1 0 1797 0 1 54435
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_673
timestamp 1649977179
transform 1 0 1797 0 1 56787
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_674
timestamp 1649977179
transform 1 0 1797 0 1 62163
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_675
timestamp 1649977179
transform 1 0 1797 0 1 61827
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_676
timestamp 1649977179
transform 1 0 1797 0 1 61491
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_677
timestamp 1649977179
transform 1 0 1797 0 1 61155
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_678
timestamp 1649977179
transform 1 0 1797 0 1 60819
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_679
timestamp 1649977179
transform 1 0 1797 0 1 60483
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_680
timestamp 1649977179
transform 1 0 1797 0 1 60147
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_681
timestamp 1649977179
transform 1 0 1797 0 1 59811
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_682
timestamp 1649977179
transform 1 0 1797 0 1 59475
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_683
timestamp 1649977179
transform 1 0 1797 0 1 59139
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_684
timestamp 1649977179
transform 1 0 1797 0 1 58803
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_685
timestamp 1649977179
transform 1 0 1797 0 1 58467
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_686
timestamp 1649977179
transform 1 0 1797 0 1 58131
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_687
timestamp 1649977179
transform 1 0 1797 0 1 57795
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_688
timestamp 1649977179
transform 1 0 1797 0 1 57459
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_689
timestamp 1649977179
transform 1 0 1797 0 1 57123
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_690
timestamp 1649977179
transform 1 0 1797 0 1 63507
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_691
timestamp 1649977179
transform 1 0 1797 0 1 63171
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_692
timestamp 1649977179
transform 1 0 1797 0 1 62835
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_693
timestamp 1649977179
transform 1 0 1797 0 1 67203
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_694
timestamp 1649977179
transform 1 0 1797 0 1 66867
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_695
timestamp 1649977179
transform 1 0 1797 0 1 62499
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_696
timestamp 1649977179
transform 1 0 1797 0 1 66531
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_697
timestamp 1649977179
transform 1 0 1797 0 1 66195
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_698
timestamp 1649977179
transform 1 0 1797 0 1 65859
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_699
timestamp 1649977179
transform 1 0 1797 0 1 65523
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_700
timestamp 1649977179
transform 1 0 1797 0 1 65187
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_701
timestamp 1649977179
transform 1 0 1797 0 1 64851
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_702
timestamp 1649977179
transform 1 0 1797 0 1 64515
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_703
timestamp 1649977179
transform 1 0 1797 0 1 64179
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_704
timestamp 1649977179
transform 1 0 1797 0 1 63843
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_705
timestamp 1649977179
transform 1 0 1797 0 1 68211
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_706
timestamp 1649977179
transform 1 0 1797 0 1 67875
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_707
timestamp 1649977179
transform 1 0 1797 0 1 69219
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_708
timestamp 1649977179
transform 1 0 1797 0 1 68883
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_709
timestamp 1649977179
transform 1 0 1797 0 1 68547
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_710
timestamp 1649977179
transform 1 0 1797 0 1 72243
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_711
timestamp 1649977179
transform 1 0 1797 0 1 71907
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_712
timestamp 1649977179
transform 1 0 1797 0 1 71571
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_713
timestamp 1649977179
transform 1 0 1797 0 1 71235
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_714
timestamp 1649977179
transform 1 0 1797 0 1 70899
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_715
timestamp 1649977179
transform 1 0 1797 0 1 70563
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_716
timestamp 1649977179
transform 1 0 1797 0 1 70227
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_717
timestamp 1649977179
transform 1 0 1797 0 1 69891
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_718
timestamp 1649977179
transform 1 0 1797 0 1 69555
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_719
timestamp 1649977179
transform 1 0 1797 0 1 67539
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_720
timestamp 1649977179
transform 1 0 1797 0 1 77619
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_721
timestamp 1649977179
transform 1 0 1797 0 1 72915
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_722
timestamp 1649977179
transform 1 0 1797 0 1 76611
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_723
timestamp 1649977179
transform 1 0 1797 0 1 76275
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_724
timestamp 1649977179
transform 1 0 1797 0 1 77283
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_725
timestamp 1649977179
transform 1 0 1797 0 1 75939
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_726
timestamp 1649977179
transform 1 0 1797 0 1 75603
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_727
timestamp 1649977179
transform 1 0 1797 0 1 75267
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_728
timestamp 1649977179
transform 1 0 1797 0 1 74931
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_729
timestamp 1649977179
transform 1 0 1797 0 1 74595
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_730
timestamp 1649977179
transform 1 0 1797 0 1 74259
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_731
timestamp 1649977179
transform 1 0 1797 0 1 73923
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_732
timestamp 1649977179
transform 1 0 1797 0 1 76947
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_733
timestamp 1649977179
transform 1 0 1797 0 1 73587
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_734
timestamp 1649977179
transform 1 0 1797 0 1 73251
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_735
timestamp 1649977179
transform 1 0 1797 0 1 78627
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_736
timestamp 1649977179
transform 1 0 1797 0 1 78291
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_737
timestamp 1649977179
transform 1 0 1797 0 1 77955
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_738
timestamp 1649977179
transform 1 0 1797 0 1 80307
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_739
timestamp 1649977179
transform 1 0 1797 0 1 79971
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_740
timestamp 1649977179
transform 1 0 1797 0 1 79635
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_741
timestamp 1649977179
transform 1 0 1797 0 1 79299
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_742
timestamp 1649977179
transform 1 0 1797 0 1 78963
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_743
timestamp 1649977179
transform 1 0 3477 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_744
timestamp 1649977179
transform 1 0 3141 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_745
timestamp 1649977179
transform 1 0 2805 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_746
timestamp 1649977179
transform 1 0 2469 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_747
timestamp 1649977179
transform 1 0 2133 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_748
timestamp 1649977179
transform 1 0 1797 0 1 80979
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_749
timestamp 1649977179
transform 1 0 1797 0 1 80643
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_750
timestamp 1649977179
transform 1 0 4149 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_751
timestamp 1649977179
transform 1 0 3813 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_752
timestamp 1649977179
transform 1 0 8517 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_753
timestamp 1649977179
transform 1 0 8181 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_754
timestamp 1649977179
transform 1 0 7845 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_755
timestamp 1649977179
transform 1 0 7509 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_756
timestamp 1649977179
transform 1 0 7173 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_757
timestamp 1649977179
transform 1 0 6837 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_758
timestamp 1649977179
transform 1 0 6501 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_759
timestamp 1649977179
transform 1 0 6165 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_760
timestamp 1649977179
transform 1 0 5829 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_761
timestamp 1649977179
transform 1 0 5493 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_762
timestamp 1649977179
transform 1 0 5157 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_763
timestamp 1649977179
transform 1 0 4821 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_764
timestamp 1649977179
transform 1 0 4485 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_765
timestamp 1649977179
transform 1 0 8853 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_766
timestamp 1649977179
transform 1 0 16917 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_767
timestamp 1649977179
transform 1 0 16581 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_768
timestamp 1649977179
transform 1 0 16245 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_769
timestamp 1649977179
transform 1 0 15909 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_770
timestamp 1649977179
transform 1 0 15573 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_771
timestamp 1649977179
transform 1 0 15237 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_772
timestamp 1649977179
transform 1 0 14901 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_773
timestamp 1649977179
transform 1 0 14565 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_774
timestamp 1649977179
transform 1 0 14229 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_775
timestamp 1649977179
transform 1 0 13893 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_776
timestamp 1649977179
transform 1 0 13557 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_777
timestamp 1649977179
transform 1 0 13221 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_778
timestamp 1649977179
transform 1 0 12885 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_779
timestamp 1649977179
transform 1 0 12549 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_780
timestamp 1649977179
transform 1 0 12213 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_781
timestamp 1649977179
transform 1 0 11877 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_782
timestamp 1649977179
transform 1 0 11541 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_783
timestamp 1649977179
transform 1 0 11205 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_784
timestamp 1649977179
transform 1 0 10869 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_785
timestamp 1649977179
transform 1 0 10533 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_786
timestamp 1649977179
transform 1 0 10197 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_787
timestamp 1649977179
transform 1 0 9861 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_788
timestamp 1649977179
transform 1 0 9525 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_789
timestamp 1649977179
transform 1 0 9189 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_790
timestamp 1649977179
transform 1 0 24981 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_791
timestamp 1649977179
transform 1 0 24645 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_792
timestamp 1649977179
transform 1 0 24309 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_793
timestamp 1649977179
transform 1 0 23973 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_794
timestamp 1649977179
transform 1 0 23637 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_795
timestamp 1649977179
transform 1 0 23301 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_796
timestamp 1649977179
transform 1 0 22965 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_797
timestamp 1649977179
transform 1 0 22629 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_798
timestamp 1649977179
transform 1 0 22293 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_799
timestamp 1649977179
transform 1 0 21957 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_800
timestamp 1649977179
transform 1 0 21621 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_801
timestamp 1649977179
transform 1 0 21285 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_802
timestamp 1649977179
transform 1 0 20949 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_803
timestamp 1649977179
transform 1 0 20613 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_804
timestamp 1649977179
transform 1 0 20277 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_805
timestamp 1649977179
transform 1 0 19941 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_806
timestamp 1649977179
transform 1 0 19605 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_807
timestamp 1649977179
transform 1 0 19269 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_808
timestamp 1649977179
transform 1 0 18933 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_809
timestamp 1649977179
transform 1 0 18597 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_810
timestamp 1649977179
transform 1 0 18261 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_811
timestamp 1649977179
transform 1 0 17925 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_812
timestamp 1649977179
transform 1 0 17589 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_813
timestamp 1649977179
transform 1 0 25653 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_814
timestamp 1649977179
transform 1 0 25317 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_815
timestamp 1649977179
transform 1 0 34053 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_816
timestamp 1649977179
transform 1 0 33717 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_817
timestamp 1649977179
transform 1 0 33381 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_818
timestamp 1649977179
transform 1 0 33045 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_819
timestamp 1649977179
transform 1 0 32709 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_820
timestamp 1649977179
transform 1 0 32373 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_821
timestamp 1649977179
transform 1 0 32037 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_822
timestamp 1649977179
transform 1 0 31701 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_823
timestamp 1649977179
transform 1 0 31365 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_824
timestamp 1649977179
transform 1 0 31029 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_825
timestamp 1649977179
transform 1 0 30693 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_826
timestamp 1649977179
transform 1 0 30357 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_827
timestamp 1649977179
transform 1 0 30021 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_828
timestamp 1649977179
transform 1 0 29685 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_829
timestamp 1649977179
transform 1 0 29349 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_830
timestamp 1649977179
transform 1 0 29013 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_831
timestamp 1649977179
transform 1 0 28677 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_832
timestamp 1649977179
transform 1 0 28341 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_833
timestamp 1649977179
transform 1 0 28005 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_834
timestamp 1649977179
transform 1 0 27669 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_835
timestamp 1649977179
transform 1 0 27333 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_836
timestamp 1649977179
transform 1 0 26997 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_837
timestamp 1649977179
transform 1 0 26661 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_838
timestamp 1649977179
transform 1 0 26325 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_839
timestamp 1649977179
transform 1 0 25989 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_840
timestamp 1649977179
transform 1 0 17253 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_841
timestamp 1649977179
transform 1 0 1797 0 1 72579
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_842
timestamp 1649977179
transform 1 0 37413 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_843
timestamp 1649977179
transform 1 0 37077 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_844
timestamp 1649977179
transform 1 0 36741 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_845
timestamp 1649977179
transform 1 0 36405 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_846
timestamp 1649977179
transform 1 0 36069 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_847
timestamp 1649977179
transform 1 0 35733 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_848
timestamp 1649977179
transform 1 0 35397 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_849
timestamp 1649977179
transform 1 0 35061 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_850
timestamp 1649977179
transform 1 0 34725 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_851
timestamp 1649977179
transform 1 0 34389 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_852
timestamp 1649977179
transform 1 0 42453 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_853
timestamp 1649977179
transform 1 0 42117 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_854
timestamp 1649977179
transform 1 0 41781 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_855
timestamp 1649977179
transform 1 0 41445 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_856
timestamp 1649977179
transform 1 0 41109 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_857
timestamp 1649977179
transform 1 0 40773 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_858
timestamp 1649977179
transform 1 0 40437 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_859
timestamp 1649977179
transform 1 0 40101 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_860
timestamp 1649977179
transform 1 0 39765 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_861
timestamp 1649977179
transform 1 0 39429 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_862
timestamp 1649977179
transform 1 0 39093 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_863
timestamp 1649977179
transform 1 0 38757 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_864
timestamp 1649977179
transform 1 0 38421 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_865
timestamp 1649977179
transform 1 0 38085 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_866
timestamp 1649977179
transform 1 0 37749 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_867
timestamp 1649977179
transform 1 0 46485 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_868
timestamp 1649977179
transform 1 0 46149 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_869
timestamp 1649977179
transform 1 0 45813 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_870
timestamp 1649977179
transform 1 0 45477 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_871
timestamp 1649977179
transform 1 0 45141 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_872
timestamp 1649977179
transform 1 0 44805 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_873
timestamp 1649977179
transform 1 0 44469 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_874
timestamp 1649977179
transform 1 0 44133 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_875
timestamp 1649977179
transform 1 0 43797 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_876
timestamp 1649977179
transform 1 0 43461 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_877
timestamp 1649977179
transform 1 0 43125 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_878
timestamp 1649977179
transform 1 0 46821 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_879
timestamp 1649977179
transform 1 0 51189 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_880
timestamp 1649977179
transform 1 0 50853 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_881
timestamp 1649977179
transform 1 0 50517 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_882
timestamp 1649977179
transform 1 0 50181 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_883
timestamp 1649977179
transform 1 0 49845 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_884
timestamp 1649977179
transform 1 0 49509 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_885
timestamp 1649977179
transform 1 0 49173 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_886
timestamp 1649977179
transform 1 0 48837 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_887
timestamp 1649977179
transform 1 0 48501 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_888
timestamp 1649977179
transform 1 0 48165 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_889
timestamp 1649977179
transform 1 0 47829 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_890
timestamp 1649977179
transform 1 0 47493 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_891
timestamp 1649977179
transform 1 0 47157 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_892
timestamp 1649977179
transform 1 0 42789 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_893
timestamp 1649977179
transform 1 0 51525 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_894
timestamp 1649977179
transform 1 0 58581 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_895
timestamp 1649977179
transform 1 0 58245 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_896
timestamp 1649977179
transform 1 0 57909 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_897
timestamp 1649977179
transform 1 0 57573 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_898
timestamp 1649977179
transform 1 0 57237 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_899
timestamp 1649977179
transform 1 0 56901 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_900
timestamp 1649977179
transform 1 0 56565 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_901
timestamp 1649977179
transform 1 0 56229 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_902
timestamp 1649977179
transform 1 0 55893 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_903
timestamp 1649977179
transform 1 0 55557 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_904
timestamp 1649977179
transform 1 0 55221 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_905
timestamp 1649977179
transform 1 0 54885 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_906
timestamp 1649977179
transform 1 0 54549 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_907
timestamp 1649977179
transform 1 0 54213 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_908
timestamp 1649977179
transform 1 0 53877 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_909
timestamp 1649977179
transform 1 0 53541 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_910
timestamp 1649977179
transform 1 0 53205 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_911
timestamp 1649977179
transform 1 0 52869 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_912
timestamp 1649977179
transform 1 0 52533 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_913
timestamp 1649977179
transform 1 0 52197 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_914
timestamp 1649977179
transform 1 0 51861 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_915
timestamp 1649977179
transform 1 0 59589 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_916
timestamp 1649977179
transform 1 0 59253 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_917
timestamp 1649977179
transform 1 0 58917 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_918
timestamp 1649977179
transform 1 0 67989 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_919
timestamp 1649977179
transform 1 0 67653 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_920
timestamp 1649977179
transform 1 0 67317 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_921
timestamp 1649977179
transform 1 0 66981 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_922
timestamp 1649977179
transform 1 0 66645 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_923
timestamp 1649977179
transform 1 0 66309 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_924
timestamp 1649977179
transform 1 0 65973 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_925
timestamp 1649977179
transform 1 0 65637 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_926
timestamp 1649977179
transform 1 0 65301 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_927
timestamp 1649977179
transform 1 0 64965 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_928
timestamp 1649977179
transform 1 0 64629 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_929
timestamp 1649977179
transform 1 0 64293 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_930
timestamp 1649977179
transform 1 0 63957 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_931
timestamp 1649977179
transform 1 0 63621 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_932
timestamp 1649977179
transform 1 0 63285 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_933
timestamp 1649977179
transform 1 0 62949 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_934
timestamp 1649977179
transform 1 0 62613 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_935
timestamp 1649977179
transform 1 0 62277 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_936
timestamp 1649977179
transform 1 0 61941 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_937
timestamp 1649977179
transform 1 0 61605 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_938
timestamp 1649977179
transform 1 0 61269 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_939
timestamp 1649977179
transform 1 0 60933 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_940
timestamp 1649977179
transform 1 0 60597 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_941
timestamp 1649977179
transform 1 0 60261 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_942
timestamp 1649977179
transform 1 0 59925 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_943
timestamp 1649977179
transform 1 0 134847 0 1 44019
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_944
timestamp 1649977179
transform 1 0 134847 0 1 43683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_945
timestamp 1649977179
transform 1 0 134847 0 1 43347
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_946
timestamp 1649977179
transform 1 0 134847 0 1 43011
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_947
timestamp 1649977179
transform 1 0 134847 0 1 45027
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_948
timestamp 1649977179
transform 1 0 134847 0 1 46035
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_949
timestamp 1649977179
transform 1 0 134847 0 1 42675
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_950
timestamp 1649977179
transform 1 0 134847 0 1 42339
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_951
timestamp 1649977179
transform 1 0 134847 0 1 45363
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_952
timestamp 1649977179
transform 1 0 134847 0 1 42003
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_953
timestamp 1649977179
transform 1 0 134847 0 1 44691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_954
timestamp 1649977179
transform 1 0 134847 0 1 44355
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_955
timestamp 1649977179
transform 1 0 134847 0 1 46371
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_956
timestamp 1649977179
transform 1 0 134847 0 1 45699
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_957
timestamp 1649977179
transform 1 0 134847 0 1 47715
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_958
timestamp 1649977179
transform 1 0 134847 0 1 48723
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_959
timestamp 1649977179
transform 1 0 134847 0 1 47379
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_960
timestamp 1649977179
transform 1 0 134847 0 1 47043
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_961
timestamp 1649977179
transform 1 0 134847 0 1 48051
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_962
timestamp 1649977179
transform 1 0 134847 0 1 49731
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_963
timestamp 1649977179
transform 1 0 134847 0 1 49395
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_964
timestamp 1649977179
transform 1 0 134847 0 1 48387
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_965
timestamp 1649977179
transform 1 0 134847 0 1 51747
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_966
timestamp 1649977179
transform 1 0 134847 0 1 50403
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_967
timestamp 1649977179
transform 1 0 134847 0 1 51411
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_968
timestamp 1649977179
transform 1 0 134847 0 1 51075
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_969
timestamp 1649977179
transform 1 0 134847 0 1 50739
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_970
timestamp 1649977179
transform 1 0 134847 0 1 49059
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_971
timestamp 1649977179
transform 1 0 134847 0 1 50067
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_972
timestamp 1649977179
transform 1 0 134847 0 1 46707
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_973
timestamp 1649977179
transform 1 0 134847 0 1 52419
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_974
timestamp 1649977179
transform 1 0 134847 0 1 56787
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_975
timestamp 1649977179
transform 1 0 134847 0 1 52083
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_976
timestamp 1649977179
transform 1 0 134847 0 1 56451
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_977
timestamp 1649977179
transform 1 0 134847 0 1 56115
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_978
timestamp 1649977179
transform 1 0 134847 0 1 55779
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_979
timestamp 1649977179
transform 1 0 134847 0 1 55443
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_980
timestamp 1649977179
transform 1 0 134847 0 1 55107
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_981
timestamp 1649977179
transform 1 0 134847 0 1 54771
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_982
timestamp 1649977179
transform 1 0 134847 0 1 54435
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_983
timestamp 1649977179
transform 1 0 134847 0 1 54099
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_984
timestamp 1649977179
transform 1 0 134847 0 1 53763
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_985
timestamp 1649977179
transform 1 0 134847 0 1 53427
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_986
timestamp 1649977179
transform 1 0 134847 0 1 53091
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_987
timestamp 1649977179
transform 1 0 134847 0 1 52755
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_988
timestamp 1649977179
transform 1 0 134847 0 1 62163
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_989
timestamp 1649977179
transform 1 0 134847 0 1 61827
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_990
timestamp 1649977179
transform 1 0 134847 0 1 61491
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_991
timestamp 1649977179
transform 1 0 134847 0 1 61155
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_992
timestamp 1649977179
transform 1 0 134847 0 1 60819
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_993
timestamp 1649977179
transform 1 0 134847 0 1 60483
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_994
timestamp 1649977179
transform 1 0 134847 0 1 60147
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_995
timestamp 1649977179
transform 1 0 134847 0 1 59811
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_996
timestamp 1649977179
transform 1 0 134847 0 1 59475
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_997
timestamp 1649977179
transform 1 0 134847 0 1 59139
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_998
timestamp 1649977179
transform 1 0 134847 0 1 58803
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_999
timestamp 1649977179
transform 1 0 134847 0 1 58467
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1000
timestamp 1649977179
transform 1 0 134847 0 1 58131
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1001
timestamp 1649977179
transform 1 0 134847 0 1 57795
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1002
timestamp 1649977179
transform 1 0 134847 0 1 57459
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1003
timestamp 1649977179
transform 1 0 134847 0 1 57123
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1004
timestamp 1649977179
transform 1 0 76389 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1005
timestamp 1649977179
transform 1 0 76053 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1006
timestamp 1649977179
transform 1 0 75717 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1007
timestamp 1649977179
transform 1 0 75381 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1008
timestamp 1649977179
transform 1 0 75045 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1009
timestamp 1649977179
transform 1 0 74709 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1010
timestamp 1649977179
transform 1 0 74373 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1011
timestamp 1649977179
transform 1 0 74037 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1012
timestamp 1649977179
transform 1 0 73701 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1013
timestamp 1649977179
transform 1 0 68661 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1014
timestamp 1649977179
transform 1 0 73365 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1015
timestamp 1649977179
transform 1 0 73029 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1016
timestamp 1649977179
transform 1 0 72693 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1017
timestamp 1649977179
transform 1 0 72357 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1018
timestamp 1649977179
transform 1 0 72021 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1019
timestamp 1649977179
transform 1 0 71685 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1020
timestamp 1649977179
transform 1 0 71349 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1021
timestamp 1649977179
transform 1 0 71013 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1022
timestamp 1649977179
transform 1 0 70677 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1023
timestamp 1649977179
transform 1 0 70341 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1024
timestamp 1649977179
transform 1 0 70005 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1025
timestamp 1649977179
transform 1 0 69669 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1026
timestamp 1649977179
transform 1 0 69333 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1027
timestamp 1649977179
transform 1 0 68997 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1028
timestamp 1649977179
transform 1 0 85125 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1029
timestamp 1649977179
transform 1 0 84789 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1030
timestamp 1649977179
transform 1 0 84453 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1031
timestamp 1649977179
transform 1 0 84117 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1032
timestamp 1649977179
transform 1 0 83781 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1033
timestamp 1649977179
transform 1 0 83445 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1034
timestamp 1649977179
transform 1 0 83109 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1035
timestamp 1649977179
transform 1 0 82773 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1036
timestamp 1649977179
transform 1 0 82437 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1037
timestamp 1649977179
transform 1 0 82101 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1038
timestamp 1649977179
transform 1 0 81765 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1039
timestamp 1649977179
transform 1 0 81429 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1040
timestamp 1649977179
transform 1 0 81093 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1041
timestamp 1649977179
transform 1 0 80757 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1042
timestamp 1649977179
transform 1 0 80421 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1043
timestamp 1649977179
transform 1 0 80085 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1044
timestamp 1649977179
transform 1 0 79749 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1045
timestamp 1649977179
transform 1 0 79413 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1046
timestamp 1649977179
transform 1 0 79077 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1047
timestamp 1649977179
transform 1 0 78741 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1048
timestamp 1649977179
transform 1 0 78405 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1049
timestamp 1649977179
transform 1 0 78069 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1050
timestamp 1649977179
transform 1 0 77733 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1051
timestamp 1649977179
transform 1 0 77397 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1052
timestamp 1649977179
transform 1 0 77061 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1053
timestamp 1649977179
transform 1 0 76725 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1054
timestamp 1649977179
transform 1 0 86469 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1055
timestamp 1649977179
transform 1 0 86133 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1056
timestamp 1649977179
transform 1 0 85797 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1057
timestamp 1649977179
transform 1 0 85461 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1058
timestamp 1649977179
transform 1 0 93525 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1059
timestamp 1649977179
transform 1 0 93189 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1060
timestamp 1649977179
transform 1 0 92853 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1061
timestamp 1649977179
transform 1 0 92517 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1062
timestamp 1649977179
transform 1 0 92181 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1063
timestamp 1649977179
transform 1 0 91845 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1064
timestamp 1649977179
transform 1 0 91509 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1065
timestamp 1649977179
transform 1 0 91173 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1066
timestamp 1649977179
transform 1 0 90837 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1067
timestamp 1649977179
transform 1 0 90501 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1068
timestamp 1649977179
transform 1 0 90165 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1069
timestamp 1649977179
transform 1 0 89829 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1070
timestamp 1649977179
transform 1 0 89493 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1071
timestamp 1649977179
transform 1 0 89157 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1072
timestamp 1649977179
transform 1 0 88821 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1073
timestamp 1649977179
transform 1 0 88485 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1074
timestamp 1649977179
transform 1 0 88149 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1075
timestamp 1649977179
transform 1 0 87813 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1076
timestamp 1649977179
transform 1 0 87477 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1077
timestamp 1649977179
transform 1 0 87141 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1078
timestamp 1649977179
transform 1 0 86805 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1079
timestamp 1649977179
transform 1 0 101925 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1080
timestamp 1649977179
transform 1 0 101589 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1081
timestamp 1649977179
transform 1 0 101253 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1082
timestamp 1649977179
transform 1 0 100917 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1083
timestamp 1649977179
transform 1 0 100581 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1084
timestamp 1649977179
transform 1 0 100245 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1085
timestamp 1649977179
transform 1 0 99909 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1086
timestamp 1649977179
transform 1 0 99573 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1087
timestamp 1649977179
transform 1 0 99237 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1088
timestamp 1649977179
transform 1 0 98901 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1089
timestamp 1649977179
transform 1 0 98565 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1090
timestamp 1649977179
transform 1 0 98229 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1091
timestamp 1649977179
transform 1 0 97893 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1092
timestamp 1649977179
transform 1 0 97557 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1093
timestamp 1649977179
transform 1 0 97221 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1094
timestamp 1649977179
transform 1 0 96885 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1095
timestamp 1649977179
transform 1 0 96549 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1096
timestamp 1649977179
transform 1 0 96213 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1097
timestamp 1649977179
transform 1 0 95877 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1098
timestamp 1649977179
transform 1 0 95541 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1099
timestamp 1649977179
transform 1 0 95205 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1100
timestamp 1649977179
transform 1 0 94869 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1101
timestamp 1649977179
transform 1 0 94533 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1102
timestamp 1649977179
transform 1 0 94197 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1103
timestamp 1649977179
transform 1 0 93861 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1104
timestamp 1649977179
transform 1 0 134847 0 1 63507
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1105
timestamp 1649977179
transform 1 0 134847 0 1 62499
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1106
timestamp 1649977179
transform 1 0 134847 0 1 63171
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1107
timestamp 1649977179
transform 1 0 134847 0 1 62835
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1108
timestamp 1649977179
transform 1 0 134847 0 1 67203
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1109
timestamp 1649977179
transform 1 0 134847 0 1 66867
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1110
timestamp 1649977179
transform 1 0 134847 0 1 66531
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1111
timestamp 1649977179
transform 1 0 134847 0 1 66195
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1112
timestamp 1649977179
transform 1 0 134847 0 1 65859
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1113
timestamp 1649977179
transform 1 0 134847 0 1 65523
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1114
timestamp 1649977179
transform 1 0 134847 0 1 65187
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1115
timestamp 1649977179
transform 1 0 134847 0 1 64851
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1116
timestamp 1649977179
transform 1 0 134847 0 1 64515
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1117
timestamp 1649977179
transform 1 0 134847 0 1 64179
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1118
timestamp 1649977179
transform 1 0 134847 0 1 63843
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1119
timestamp 1649977179
transform 1 0 134847 0 1 67875
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1120
timestamp 1649977179
transform 1 0 134847 0 1 72243
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1121
timestamp 1649977179
transform 1 0 134847 0 1 71907
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1122
timestamp 1649977179
transform 1 0 134847 0 1 71571
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1123
timestamp 1649977179
transform 1 0 134847 0 1 71235
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1124
timestamp 1649977179
transform 1 0 134847 0 1 70899
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1125
timestamp 1649977179
transform 1 0 134847 0 1 70563
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1126
timestamp 1649977179
transform 1 0 134847 0 1 70227
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1127
timestamp 1649977179
transform 1 0 134847 0 1 69891
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1128
timestamp 1649977179
transform 1 0 134847 0 1 69555
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1129
timestamp 1649977179
transform 1 0 134847 0 1 69219
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1130
timestamp 1649977179
transform 1 0 134847 0 1 68883
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1131
timestamp 1649977179
transform 1 0 134847 0 1 68547
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1132
timestamp 1649977179
transform 1 0 134847 0 1 68211
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1133
timestamp 1649977179
transform 1 0 134847 0 1 67539
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1134
timestamp 1649977179
transform 1 0 102933 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1135
timestamp 1649977179
transform 1 0 102597 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1136
timestamp 1649977179
transform 1 0 106293 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1137
timestamp 1649977179
transform 1 0 105957 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1138
timestamp 1649977179
transform 1 0 105621 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1139
timestamp 1649977179
transform 1 0 105285 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1140
timestamp 1649977179
transform 1 0 104949 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1141
timestamp 1649977179
transform 1 0 104613 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1142
timestamp 1649977179
transform 1 0 104277 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1143
timestamp 1649977179
transform 1 0 103941 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1144
timestamp 1649977179
transform 1 0 103605 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1145
timestamp 1649977179
transform 1 0 103269 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1146
timestamp 1649977179
transform 1 0 110661 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1147
timestamp 1649977179
transform 1 0 110325 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1148
timestamp 1649977179
transform 1 0 109989 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1149
timestamp 1649977179
transform 1 0 109653 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1150
timestamp 1649977179
transform 1 0 109317 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1151
timestamp 1649977179
transform 1 0 108981 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1152
timestamp 1649977179
transform 1 0 108645 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1153
timestamp 1649977179
transform 1 0 108309 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1154
timestamp 1649977179
transform 1 0 107973 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1155
timestamp 1649977179
transform 1 0 107637 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1156
timestamp 1649977179
transform 1 0 107301 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1157
timestamp 1649977179
transform 1 0 106965 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1158
timestamp 1649977179
transform 1 0 106629 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1159
timestamp 1649977179
transform 1 0 119061 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1160
timestamp 1649977179
transform 1 0 118725 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1161
timestamp 1649977179
transform 1 0 110997 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1162
timestamp 1649977179
transform 1 0 118389 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1163
timestamp 1649977179
transform 1 0 118053 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1164
timestamp 1649977179
transform 1 0 117717 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1165
timestamp 1649977179
transform 1 0 117381 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1166
timestamp 1649977179
transform 1 0 117045 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1167
timestamp 1649977179
transform 1 0 116709 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1168
timestamp 1649977179
transform 1 0 116373 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1169
timestamp 1649977179
transform 1 0 116037 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1170
timestamp 1649977179
transform 1 0 115701 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1171
timestamp 1649977179
transform 1 0 115365 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1172
timestamp 1649977179
transform 1 0 115029 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1173
timestamp 1649977179
transform 1 0 114693 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1174
timestamp 1649977179
transform 1 0 114357 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1175
timestamp 1649977179
transform 1 0 114021 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1176
timestamp 1649977179
transform 1 0 113685 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1177
timestamp 1649977179
transform 1 0 113349 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1178
timestamp 1649977179
transform 1 0 113013 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1179
timestamp 1649977179
transform 1 0 112677 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1180
timestamp 1649977179
transform 1 0 112341 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1181
timestamp 1649977179
transform 1 0 112005 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1182
timestamp 1649977179
transform 1 0 111669 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1183
timestamp 1649977179
transform 1 0 111333 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1184
timestamp 1649977179
transform 1 0 134847 0 1 77283
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1185
timestamp 1649977179
transform 1 0 134847 0 1 76947
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1186
timestamp 1649977179
transform 1 0 134847 0 1 76611
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1187
timestamp 1649977179
transform 1 0 134847 0 1 76275
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1188
timestamp 1649977179
transform 1 0 134847 0 1 75939
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1189
timestamp 1649977179
transform 1 0 134847 0 1 75603
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1190
timestamp 1649977179
transform 1 0 134847 0 1 75267
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1191
timestamp 1649977179
transform 1 0 134847 0 1 74931
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1192
timestamp 1649977179
transform 1 0 134847 0 1 74595
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1193
timestamp 1649977179
transform 1 0 134847 0 1 74259
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1194
timestamp 1649977179
transform 1 0 134847 0 1 73923
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1195
timestamp 1649977179
transform 1 0 134847 0 1 73587
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1196
timestamp 1649977179
transform 1 0 134847 0 1 73251
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1197
timestamp 1649977179
transform 1 0 134847 0 1 72915
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1198
timestamp 1649977179
transform 1 0 134847 0 1 77619
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1199
timestamp 1649977179
transform 1 0 126453 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1200
timestamp 1649977179
transform 1 0 126117 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1201
timestamp 1649977179
transform 1 0 125781 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1202
timestamp 1649977179
transform 1 0 125445 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1203
timestamp 1649977179
transform 1 0 125109 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1204
timestamp 1649977179
transform 1 0 124773 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1205
timestamp 1649977179
transform 1 0 124437 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1206
timestamp 1649977179
transform 1 0 124101 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1207
timestamp 1649977179
transform 1 0 123765 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1208
timestamp 1649977179
transform 1 0 123429 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1209
timestamp 1649977179
transform 1 0 123093 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1210
timestamp 1649977179
transform 1 0 122757 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1211
timestamp 1649977179
transform 1 0 122421 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1212
timestamp 1649977179
transform 1 0 122085 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1213
timestamp 1649977179
transform 1 0 121749 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1214
timestamp 1649977179
transform 1 0 121413 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1215
timestamp 1649977179
transform 1 0 121077 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1216
timestamp 1649977179
transform 1 0 120741 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1217
timestamp 1649977179
transform 1 0 120405 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1218
timestamp 1649977179
transform 1 0 120069 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1219
timestamp 1649977179
transform 1 0 119733 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1220
timestamp 1649977179
transform 1 0 127461 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1221
timestamp 1649977179
transform 1 0 127125 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1222
timestamp 1649977179
transform 1 0 126789 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1223
timestamp 1649977179
transform 1 0 134847 0 1 78963
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1224
timestamp 1649977179
transform 1 0 134847 0 1 78627
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1225
timestamp 1649977179
transform 1 0 134847 0 1 78291
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1226
timestamp 1649977179
transform 1 0 134847 0 1 77955
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1227
timestamp 1649977179
transform 1 0 134847 0 1 80307
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1228
timestamp 1649977179
transform 1 0 134847 0 1 79971
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1229
timestamp 1649977179
transform 1 0 134847 0 1 79635
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1230
timestamp 1649977179
transform 1 0 134847 0 1 79299
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1231
timestamp 1649977179
transform 1 0 129813 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1232
timestamp 1649977179
transform 1 0 129477 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1233
timestamp 1649977179
transform 1 0 129141 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1234
timestamp 1649977179
transform 1 0 128805 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1235
timestamp 1649977179
transform 1 0 128469 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1236
timestamp 1649977179
transform 1 0 128133 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1237
timestamp 1649977179
transform 1 0 131829 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1238
timestamp 1649977179
transform 1 0 131493 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1239
timestamp 1649977179
transform 1 0 131157 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1240
timestamp 1649977179
transform 1 0 130821 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1241
timestamp 1649977179
transform 1 0 130485 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1242
timestamp 1649977179
transform 1 0 130149 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1243
timestamp 1649977179
transform 1 0 134847 0 1 80979
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1244
timestamp 1649977179
transform 1 0 134847 0 1 80643
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1245
timestamp 1649977179
transform 1 0 134181 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1246
timestamp 1649977179
transform 1 0 133845 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1247
timestamp 1649977179
transform 1 0 133509 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1248
timestamp 1649977179
transform 1 0 133173 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1249
timestamp 1649977179
transform 1 0 132837 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1250
timestamp 1649977179
transform 1 0 132501 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1251
timestamp 1649977179
transform 1 0 132165 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1252
timestamp 1649977179
transform 1 0 127797 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1253
timestamp 1649977179
transform 1 0 134847 0 1 72579
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1254
timestamp 1649977179
transform 1 0 119397 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1255
timestamp 1649977179
transform 1 0 102261 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1256
timestamp 1649977179
transform 1 0 134847 0 1 41667
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1257
timestamp 1649977179
transform 1 0 1797 0 1 41667
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1258
timestamp 1649977179
transform 1 0 68325 0 1 81432
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1259
timestamp 1649977179
transform 1 0 68325 0 1 1683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_0
timestamp 1649977179
transform 1 0 134843 0 1 2699
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1
timestamp 1649977179
transform 1 0 134843 0 1 2363
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_2
timestamp 1649977179
transform 1 0 132833 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_3
timestamp 1649977179
transform 1 0 132497 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_4
timestamp 1649977179
transform 1 0 132161 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_5
timestamp 1649977179
transform 1 0 134177 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_6
timestamp 1649977179
transform 1 0 133841 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_7
timestamp 1649977179
transform 1 0 134843 0 1 2027
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_8
timestamp 1649977179
transform 1 0 133505 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_9
timestamp 1649977179
transform 1 0 133169 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_10
timestamp 1649977179
transform 1 0 128129 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_11
timestamp 1649977179
transform 1 0 131825 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_12
timestamp 1649977179
transform 1 0 131489 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_13
timestamp 1649977179
transform 1 0 131153 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_14
timestamp 1649977179
transform 1 0 130817 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_15
timestamp 1649977179
transform 1 0 130481 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_16
timestamp 1649977179
transform 1 0 130145 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_17
timestamp 1649977179
transform 1 0 129809 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_18
timestamp 1649977179
transform 1 0 129473 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_19
timestamp 1649977179
transform 1 0 129137 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_20
timestamp 1649977179
transform 1 0 128801 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_21
timestamp 1649977179
transform 1 0 128465 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_22
timestamp 1649977179
transform 1 0 134843 0 1 3035
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_23
timestamp 1649977179
transform 1 0 134843 0 1 3707
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_24
timestamp 1649977179
transform 1 0 134843 0 1 4043
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_25
timestamp 1649977179
transform 1 0 134843 0 1 3371
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_26
timestamp 1649977179
transform 1 0 134843 0 1 5051
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_27
timestamp 1649977179
transform 1 0 134843 0 1 4715
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_28
timestamp 1649977179
transform 1 0 134843 0 1 4379
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_29
timestamp 1649977179
transform 1 0 126449 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_30
timestamp 1649977179
transform 1 0 126113 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_31
timestamp 1649977179
transform 1 0 125777 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_32
timestamp 1649977179
transform 1 0 125441 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_33
timestamp 1649977179
transform 1 0 125105 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_34
timestamp 1649977179
transform 1 0 124769 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_35
timestamp 1649977179
transform 1 0 124433 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_36
timestamp 1649977179
transform 1 0 124097 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_37
timestamp 1649977179
transform 1 0 123761 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_38
timestamp 1649977179
transform 1 0 123425 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_39
timestamp 1649977179
transform 1 0 123089 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_40
timestamp 1649977179
transform 1 0 122753 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_41
timestamp 1649977179
transform 1 0 122417 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_42
timestamp 1649977179
transform 1 0 122081 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_43
timestamp 1649977179
transform 1 0 121745 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_44
timestamp 1649977179
transform 1 0 121409 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_45
timestamp 1649977179
transform 1 0 121073 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_46
timestamp 1649977179
transform 1 0 120737 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_47
timestamp 1649977179
transform 1 0 120401 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_48
timestamp 1649977179
transform 1 0 120065 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_49
timestamp 1649977179
transform 1 0 119729 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_50
timestamp 1649977179
transform 1 0 119393 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_51
timestamp 1649977179
transform 1 0 127457 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_52
timestamp 1649977179
transform 1 0 127121 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_53
timestamp 1649977179
transform 1 0 126785 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_54
timestamp 1649977179
transform 1 0 134843 0 1 10427
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_55
timestamp 1649977179
transform 1 0 134843 0 1 10091
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_56
timestamp 1649977179
transform 1 0 134843 0 1 9755
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_57
timestamp 1649977179
transform 1 0 134843 0 1 9419
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_58
timestamp 1649977179
transform 1 0 134843 0 1 9083
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_59
timestamp 1649977179
transform 1 0 134843 0 1 8747
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_60
timestamp 1649977179
transform 1 0 134843 0 1 8411
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_61
timestamp 1649977179
transform 1 0 134843 0 1 8075
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_62
timestamp 1649977179
transform 1 0 134843 0 1 7739
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_63
timestamp 1649977179
transform 1 0 134843 0 1 7403
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_64
timestamp 1649977179
transform 1 0 134843 0 1 7067
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_65
timestamp 1649977179
transform 1 0 134843 0 1 6731
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_66
timestamp 1649977179
transform 1 0 134843 0 1 6395
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_67
timestamp 1649977179
transform 1 0 134843 0 1 6059
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_68
timestamp 1649977179
transform 1 0 134843 0 1 5723
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_69
timestamp 1649977179
transform 1 0 134843 0 1 5387
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_70
timestamp 1649977179
transform 1 0 127793 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_71
timestamp 1649977179
transform 1 0 115025 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_72
timestamp 1649977179
transform 1 0 111665 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_73
timestamp 1649977179
transform 1 0 114689 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_74
timestamp 1649977179
transform 1 0 114353 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_75
timestamp 1649977179
transform 1 0 117377 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_76
timestamp 1649977179
transform 1 0 111329 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_77
timestamp 1649977179
transform 1 0 115697 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_78
timestamp 1649977179
transform 1 0 114017 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_79
timestamp 1649977179
transform 1 0 110993 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_80
timestamp 1649977179
transform 1 0 119057 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_81
timestamp 1649977179
transform 1 0 118721 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_82
timestamp 1649977179
transform 1 0 113681 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_83
timestamp 1649977179
transform 1 0 117041 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_84
timestamp 1649977179
transform 1 0 116369 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_85
timestamp 1649977179
transform 1 0 116705 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_86
timestamp 1649977179
transform 1 0 118385 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_87
timestamp 1649977179
transform 1 0 113345 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_88
timestamp 1649977179
transform 1 0 116033 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_89
timestamp 1649977179
transform 1 0 113009 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_90
timestamp 1649977179
transform 1 0 112673 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_91
timestamp 1649977179
transform 1 0 112337 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_92
timestamp 1649977179
transform 1 0 118049 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_93
timestamp 1649977179
transform 1 0 112001 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_94
timestamp 1649977179
transform 1 0 115361 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_95
timestamp 1649977179
transform 1 0 117713 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_96
timestamp 1649977179
transform 1 0 104273 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_97
timestamp 1649977179
transform 1 0 108977 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_98
timestamp 1649977179
transform 1 0 105953 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_99
timestamp 1649977179
transform 1 0 108641 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_100
timestamp 1649977179
transform 1 0 107633 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_101
timestamp 1649977179
transform 1 0 108305 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_102
timestamp 1649977179
transform 1 0 105617 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_103
timestamp 1649977179
transform 1 0 107297 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_104
timestamp 1649977179
transform 1 0 103937 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_105
timestamp 1649977179
transform 1 0 103601 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_106
timestamp 1649977179
transform 1 0 104609 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_107
timestamp 1649977179
transform 1 0 103265 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_108
timestamp 1649977179
transform 1 0 102929 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_109
timestamp 1649977179
transform 1 0 102593 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_110
timestamp 1649977179
transform 1 0 105281 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_111
timestamp 1649977179
transform 1 0 104945 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_112
timestamp 1649977179
transform 1 0 106961 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_113
timestamp 1649977179
transform 1 0 106625 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_114
timestamp 1649977179
transform 1 0 110657 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_115
timestamp 1649977179
transform 1 0 110321 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_116
timestamp 1649977179
transform 1 0 107969 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_117
timestamp 1649977179
transform 1 0 109985 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_118
timestamp 1649977179
transform 1 0 106289 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_119
timestamp 1649977179
transform 1 0 109649 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_120
timestamp 1649977179
transform 1 0 109313 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_121
timestamp 1649977179
transform 1 0 134843 0 1 15131
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_122
timestamp 1649977179
transform 1 0 134843 0 1 14795
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_123
timestamp 1649977179
transform 1 0 134843 0 1 14459
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_124
timestamp 1649977179
transform 1 0 134843 0 1 14123
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_125
timestamp 1649977179
transform 1 0 134843 0 1 13787
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_126
timestamp 1649977179
transform 1 0 134843 0 1 13451
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_127
timestamp 1649977179
transform 1 0 134843 0 1 13115
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_128
timestamp 1649977179
transform 1 0 134843 0 1 12779
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_129
timestamp 1649977179
transform 1 0 134843 0 1 12443
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_130
timestamp 1649977179
transform 1 0 134843 0 1 12107
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_131
timestamp 1649977179
transform 1 0 134843 0 1 11771
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_132
timestamp 1649977179
transform 1 0 134843 0 1 11435
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_133
timestamp 1649977179
transform 1 0 134843 0 1 11099
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_134
timestamp 1649977179
transform 1 0 134843 0 1 10763
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_135
timestamp 1649977179
transform 1 0 134843 0 1 15467
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_136
timestamp 1649977179
transform 1 0 134843 0 1 20843
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_137
timestamp 1649977179
transform 1 0 134843 0 1 20507
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_138
timestamp 1649977179
transform 1 0 134843 0 1 20171
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_139
timestamp 1649977179
transform 1 0 134843 0 1 19835
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_140
timestamp 1649977179
transform 1 0 134843 0 1 19499
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_141
timestamp 1649977179
transform 1 0 134843 0 1 19163
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_142
timestamp 1649977179
transform 1 0 134843 0 1 18827
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_143
timestamp 1649977179
transform 1 0 134843 0 1 18491
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_144
timestamp 1649977179
transform 1 0 134843 0 1 18155
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_145
timestamp 1649977179
transform 1 0 134843 0 1 17819
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_146
timestamp 1649977179
transform 1 0 134843 0 1 17483
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_147
timestamp 1649977179
transform 1 0 134843 0 1 17147
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_148
timestamp 1649977179
transform 1 0 134843 0 1 16811
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_149
timestamp 1649977179
transform 1 0 134843 0 1 16475
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_150
timestamp 1649977179
transform 1 0 134843 0 1 16139
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_151
timestamp 1649977179
transform 1 0 134843 0 1 15803
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_152
timestamp 1649977179
transform 1 0 97889 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_153
timestamp 1649977179
transform 1 0 97553 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_154
timestamp 1649977179
transform 1 0 97217 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_155
timestamp 1649977179
transform 1 0 96881 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_156
timestamp 1649977179
transform 1 0 94529 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_157
timestamp 1649977179
transform 1 0 101921 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_158
timestamp 1649977179
transform 1 0 101585 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_159
timestamp 1649977179
transform 1 0 96545 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_160
timestamp 1649977179
transform 1 0 94193 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_161
timestamp 1649977179
transform 1 0 99233 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_162
timestamp 1649977179
transform 1 0 93857 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_163
timestamp 1649977179
transform 1 0 101249 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_164
timestamp 1649977179
transform 1 0 100913 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_165
timestamp 1649977179
transform 1 0 98897 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_166
timestamp 1649977179
transform 1 0 100577 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_167
timestamp 1649977179
transform 1 0 100241 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_168
timestamp 1649977179
transform 1 0 96209 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_169
timestamp 1649977179
transform 1 0 95873 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_170
timestamp 1649977179
transform 1 0 99905 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_171
timestamp 1649977179
transform 1 0 95537 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_172
timestamp 1649977179
transform 1 0 95201 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_173
timestamp 1649977179
transform 1 0 98561 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_174
timestamp 1649977179
transform 1 0 98225 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_175
timestamp 1649977179
transform 1 0 94865 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_176
timestamp 1649977179
transform 1 0 102257 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_177
timestamp 1649977179
transform 1 0 99569 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_178
timestamp 1649977179
transform 1 0 86129 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_179
timestamp 1649977179
transform 1 0 85793 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_180
timestamp 1649977179
transform 1 0 92177 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_181
timestamp 1649977179
transform 1 0 85457 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_182
timestamp 1649977179
transform 1 0 92849 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_183
timestamp 1649977179
transform 1 0 91841 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_184
timestamp 1649977179
transform 1 0 92513 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_185
timestamp 1649977179
transform 1 0 89825 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_186
timestamp 1649977179
transform 1 0 91505 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_187
timestamp 1649977179
transform 1 0 89489 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_188
timestamp 1649977179
transform 1 0 89153 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_189
timestamp 1649977179
transform 1 0 86465 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_190
timestamp 1649977179
transform 1 0 93521 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_191
timestamp 1649977179
transform 1 0 88817 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_192
timestamp 1649977179
transform 1 0 88481 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_193
timestamp 1649977179
transform 1 0 91169 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_194
timestamp 1649977179
transform 1 0 88145 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_195
timestamp 1649977179
transform 1 0 90833 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_196
timestamp 1649977179
transform 1 0 93185 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_197
timestamp 1649977179
transform 1 0 90497 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_198
timestamp 1649977179
transform 1 0 90161 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_199
timestamp 1649977179
transform 1 0 87809 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_200
timestamp 1649977179
transform 1 0 87473 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_201
timestamp 1649977179
transform 1 0 87137 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_202
timestamp 1649977179
transform 1 0 86801 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_203
timestamp 1649977179
transform 1 0 79409 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_204
timestamp 1649977179
transform 1 0 80081 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_205
timestamp 1649977179
transform 1 0 79073 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_206
timestamp 1649977179
transform 1 0 78401 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_207
timestamp 1649977179
transform 1 0 85121 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_208
timestamp 1649977179
transform 1 0 84785 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_209
timestamp 1649977179
transform 1 0 78737 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_210
timestamp 1649977179
transform 1 0 83441 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_211
timestamp 1649977179
transform 1 0 79745 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_212
timestamp 1649977179
transform 1 0 77729 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_213
timestamp 1649977179
transform 1 0 82097 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_214
timestamp 1649977179
transform 1 0 81761 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_215
timestamp 1649977179
transform 1 0 82769 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_216
timestamp 1649977179
transform 1 0 84449 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_217
timestamp 1649977179
transform 1 0 78065 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_218
timestamp 1649977179
transform 1 0 84113 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_219
timestamp 1649977179
transform 1 0 77057 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_220
timestamp 1649977179
transform 1 0 77393 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_221
timestamp 1649977179
transform 1 0 81425 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_222
timestamp 1649977179
transform 1 0 83777 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_223
timestamp 1649977179
transform 1 0 82433 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_224
timestamp 1649977179
transform 1 0 81089 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_225
timestamp 1649977179
transform 1 0 80753 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_226
timestamp 1649977179
transform 1 0 83105 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_227
timestamp 1649977179
transform 1 0 80417 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_228
timestamp 1649977179
transform 1 0 75041 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_229
timestamp 1649977179
transform 1 0 74705 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_230
timestamp 1649977179
transform 1 0 74369 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_231
timestamp 1649977179
transform 1 0 76049 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_232
timestamp 1649977179
transform 1 0 75713 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_233
timestamp 1649977179
transform 1 0 76721 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_234
timestamp 1649977179
transform 1 0 76385 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_235
timestamp 1649977179
transform 1 0 74033 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_236
timestamp 1649977179
transform 1 0 73697 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_237
timestamp 1649977179
transform 1 0 73361 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_238
timestamp 1649977179
transform 1 0 73025 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_239
timestamp 1649977179
transform 1 0 72689 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_240
timestamp 1649977179
transform 1 0 72353 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_241
timestamp 1649977179
transform 1 0 72017 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_242
timestamp 1649977179
transform 1 0 71681 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_243
timestamp 1649977179
transform 1 0 71345 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_244
timestamp 1649977179
transform 1 0 71009 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_245
timestamp 1649977179
transform 1 0 70673 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_246
timestamp 1649977179
transform 1 0 70337 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_247
timestamp 1649977179
transform 1 0 70001 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_248
timestamp 1649977179
transform 1 0 69665 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_249
timestamp 1649977179
transform 1 0 69329 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_250
timestamp 1649977179
transform 1 0 68993 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_251
timestamp 1649977179
transform 1 0 68657 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_252
timestamp 1649977179
transform 1 0 68321 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_253
timestamp 1649977179
transform 1 0 75377 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_254
timestamp 1649977179
transform 1 0 134843 0 1 21179
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_255
timestamp 1649977179
transform 1 0 134843 0 1 22523
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_256
timestamp 1649977179
transform 1 0 134843 0 1 24875
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_257
timestamp 1649977179
transform 1 0 134843 0 1 24539
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_258
timestamp 1649977179
transform 1 0 134843 0 1 24203
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_259
timestamp 1649977179
transform 1 0 134843 0 1 23867
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_260
timestamp 1649977179
transform 1 0 134843 0 1 23531
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_261
timestamp 1649977179
transform 1 0 134843 0 1 25883
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_262
timestamp 1649977179
transform 1 0 134843 0 1 25547
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_263
timestamp 1649977179
transform 1 0 134843 0 1 25211
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_264
timestamp 1649977179
transform 1 0 134843 0 1 23195
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_265
timestamp 1649977179
transform 1 0 134843 0 1 22187
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_266
timestamp 1649977179
transform 1 0 134843 0 1 21851
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_267
timestamp 1649977179
transform 1 0 134843 0 1 22859
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_268
timestamp 1649977179
transform 1 0 134843 0 1 21515
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_269
timestamp 1649977179
transform 1 0 134843 0 1 27227
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_270
timestamp 1649977179
transform 1 0 134843 0 1 26891
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_271
timestamp 1649977179
transform 1 0 134843 0 1 26555
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_272
timestamp 1649977179
transform 1 0 134843 0 1 26219
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_273
timestamp 1649977179
transform 1 0 134843 0 1 30923
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_274
timestamp 1649977179
transform 1 0 134843 0 1 30587
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_275
timestamp 1649977179
transform 1 0 134843 0 1 30251
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_276
timestamp 1649977179
transform 1 0 134843 0 1 29915
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_277
timestamp 1649977179
transform 1 0 134843 0 1 29579
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_278
timestamp 1649977179
transform 1 0 134843 0 1 29243
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_279
timestamp 1649977179
transform 1 0 134843 0 1 28907
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_280
timestamp 1649977179
transform 1 0 134843 0 1 28571
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_281
timestamp 1649977179
transform 1 0 134843 0 1 28235
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_282
timestamp 1649977179
transform 1 0 134843 0 1 27899
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_283
timestamp 1649977179
transform 1 0 134843 0 1 27563
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_284
timestamp 1649977179
transform 1 0 134843 0 1 31595
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_285
timestamp 1649977179
transform 1 0 134843 0 1 36299
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_286
timestamp 1649977179
transform 1 0 134843 0 1 35963
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_287
timestamp 1649977179
transform 1 0 134843 0 1 35627
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_288
timestamp 1649977179
transform 1 0 134843 0 1 35291
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_289
timestamp 1649977179
transform 1 0 134843 0 1 34955
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_290
timestamp 1649977179
transform 1 0 134843 0 1 34619
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_291
timestamp 1649977179
transform 1 0 134843 0 1 34283
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_292
timestamp 1649977179
transform 1 0 134843 0 1 33947
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_293
timestamp 1649977179
transform 1 0 134843 0 1 33611
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_294
timestamp 1649977179
transform 1 0 134843 0 1 33275
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_295
timestamp 1649977179
transform 1 0 134843 0 1 32939
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_296
timestamp 1649977179
transform 1 0 134843 0 1 32603
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_297
timestamp 1649977179
transform 1 0 134843 0 1 32267
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_298
timestamp 1649977179
transform 1 0 134843 0 1 31931
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_299
timestamp 1649977179
transform 1 0 134843 0 1 41339
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_300
timestamp 1649977179
transform 1 0 134843 0 1 41003
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_301
timestamp 1649977179
transform 1 0 134843 0 1 40667
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_302
timestamp 1649977179
transform 1 0 134843 0 1 40331
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_303
timestamp 1649977179
transform 1 0 134843 0 1 39995
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_304
timestamp 1649977179
transform 1 0 134843 0 1 39659
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_305
timestamp 1649977179
transform 1 0 134843 0 1 39323
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_306
timestamp 1649977179
transform 1 0 134843 0 1 38987
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_307
timestamp 1649977179
transform 1 0 134843 0 1 38651
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_308
timestamp 1649977179
transform 1 0 134843 0 1 38315
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_309
timestamp 1649977179
transform 1 0 134843 0 1 37979
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_310
timestamp 1649977179
transform 1 0 134843 0 1 37643
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_311
timestamp 1649977179
transform 1 0 134843 0 1 37307
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_312
timestamp 1649977179
transform 1 0 134843 0 1 36971
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_313
timestamp 1649977179
transform 1 0 134843 0 1 36635
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_314
timestamp 1649977179
transform 1 0 134843 0 1 31259
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_315
timestamp 1649977179
transform 1 0 63953 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_316
timestamp 1649977179
transform 1 0 64625 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_317
timestamp 1649977179
transform 1 0 65297 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_318
timestamp 1649977179
transform 1 0 62945 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_319
timestamp 1649977179
transform 1 0 60593 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_320
timestamp 1649977179
transform 1 0 61601 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_321
timestamp 1649977179
transform 1 0 61937 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_322
timestamp 1649977179
transform 1 0 62609 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_323
timestamp 1649977179
transform 1 0 63617 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_324
timestamp 1649977179
transform 1 0 59921 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_325
timestamp 1649977179
transform 1 0 67649 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_326
timestamp 1649977179
transform 1 0 61265 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_327
timestamp 1649977179
transform 1 0 60257 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_328
timestamp 1649977179
transform 1 0 64289 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_329
timestamp 1649977179
transform 1 0 67313 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_330
timestamp 1649977179
transform 1 0 67985 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_331
timestamp 1649977179
transform 1 0 64961 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_332
timestamp 1649977179
transform 1 0 65969 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_333
timestamp 1649977179
transform 1 0 66977 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_334
timestamp 1649977179
transform 1 0 66641 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_335
timestamp 1649977179
transform 1 0 65633 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_336
timestamp 1649977179
transform 1 0 66305 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_337
timestamp 1649977179
transform 1 0 62273 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_338
timestamp 1649977179
transform 1 0 60929 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_339
timestamp 1649977179
transform 1 0 63281 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_340
timestamp 1649977179
transform 1 0 57233 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_341
timestamp 1649977179
transform 1 0 58913 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_342
timestamp 1649977179
transform 1 0 56897 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_343
timestamp 1649977179
transform 1 0 56561 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_344
timestamp 1649977179
transform 1 0 56225 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_345
timestamp 1649977179
transform 1 0 55889 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_346
timestamp 1649977179
transform 1 0 55553 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_347
timestamp 1649977179
transform 1 0 59249 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_348
timestamp 1649977179
transform 1 0 55217 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_349
timestamp 1649977179
transform 1 0 57569 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_350
timestamp 1649977179
transform 1 0 59585 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_351
timestamp 1649977179
transform 1 0 54881 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_352
timestamp 1649977179
transform 1 0 54545 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_353
timestamp 1649977179
transform 1 0 54209 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_354
timestamp 1649977179
transform 1 0 53873 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_355
timestamp 1649977179
transform 1 0 53537 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_356
timestamp 1649977179
transform 1 0 53201 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_357
timestamp 1649977179
transform 1 0 52865 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_358
timestamp 1649977179
transform 1 0 52529 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_359
timestamp 1649977179
transform 1 0 52193 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_360
timestamp 1649977179
transform 1 0 51857 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_361
timestamp 1649977179
transform 1 0 51521 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_362
timestamp 1649977179
transform 1 0 57905 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_363
timestamp 1649977179
transform 1 0 58577 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_364
timestamp 1649977179
transform 1 0 58241 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_365
timestamp 1649977179
transform 1 0 47825 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_366
timestamp 1649977179
transform 1 0 44129 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_367
timestamp 1649977179
transform 1 0 43793 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_368
timestamp 1649977179
transform 1 0 47489 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_369
timestamp 1649977179
transform 1 0 47153 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_370
timestamp 1649977179
transform 1 0 46817 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_371
timestamp 1649977179
transform 1 0 46481 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_372
timestamp 1649977179
transform 1 0 43457 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_373
timestamp 1649977179
transform 1 0 43121 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_374
timestamp 1649977179
transform 1 0 46145 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_375
timestamp 1649977179
transform 1 0 51185 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_376
timestamp 1649977179
transform 1 0 45809 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_377
timestamp 1649977179
transform 1 0 45473 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_378
timestamp 1649977179
transform 1 0 45137 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_379
timestamp 1649977179
transform 1 0 50849 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_380
timestamp 1649977179
transform 1 0 50513 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_381
timestamp 1649977179
transform 1 0 50177 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_382
timestamp 1649977179
transform 1 0 49841 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_383
timestamp 1649977179
transform 1 0 44801 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_384
timestamp 1649977179
transform 1 0 44465 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_385
timestamp 1649977179
transform 1 0 49505 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_386
timestamp 1649977179
transform 1 0 49169 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_387
timestamp 1649977179
transform 1 0 48833 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_388
timestamp 1649977179
transform 1 0 48497 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_389
timestamp 1649977179
transform 1 0 48161 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_390
timestamp 1649977179
transform 1 0 39089 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_391
timestamp 1649977179
transform 1 0 38753 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_392
timestamp 1649977179
transform 1 0 38417 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_393
timestamp 1649977179
transform 1 0 38081 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_394
timestamp 1649977179
transform 1 0 37745 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_395
timestamp 1649977179
transform 1 0 37409 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_396
timestamp 1649977179
transform 1 0 37073 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_397
timestamp 1649977179
transform 1 0 36737 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_398
timestamp 1649977179
transform 1 0 36401 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_399
timestamp 1649977179
transform 1 0 36065 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_400
timestamp 1649977179
transform 1 0 35729 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_401
timestamp 1649977179
transform 1 0 35393 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_402
timestamp 1649977179
transform 1 0 35057 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_403
timestamp 1649977179
transform 1 0 34721 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_404
timestamp 1649977179
transform 1 0 34385 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_405
timestamp 1649977179
transform 1 0 39425 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_406
timestamp 1649977179
transform 1 0 42449 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_407
timestamp 1649977179
transform 1 0 42113 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_408
timestamp 1649977179
transform 1 0 41777 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_409
timestamp 1649977179
transform 1 0 41441 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_410
timestamp 1649977179
transform 1 0 41105 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_411
timestamp 1649977179
transform 1 0 40769 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_412
timestamp 1649977179
transform 1 0 40433 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_413
timestamp 1649977179
transform 1 0 40097 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_414
timestamp 1649977179
transform 1 0 39761 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_415
timestamp 1649977179
transform 1 0 42785 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_416
timestamp 1649977179
transform 1 0 28001 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_417
timestamp 1649977179
transform 1 0 27665 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_418
timestamp 1649977179
transform 1 0 28673 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_419
timestamp 1649977179
transform 1 0 32705 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_420
timestamp 1649977179
transform 1 0 32369 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_421
timestamp 1649977179
transform 1 0 28337 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_422
timestamp 1649977179
transform 1 0 32033 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_423
timestamp 1649977179
transform 1 0 27329 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_424
timestamp 1649977179
transform 1 0 26993 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_425
timestamp 1649977179
transform 1 0 31697 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_426
timestamp 1649977179
transform 1 0 31361 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_427
timestamp 1649977179
transform 1 0 26657 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_428
timestamp 1649977179
transform 1 0 31025 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_429
timestamp 1649977179
transform 1 0 26321 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_430
timestamp 1649977179
transform 1 0 30689 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_431
timestamp 1649977179
transform 1 0 30353 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_432
timestamp 1649977179
transform 1 0 25985 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_433
timestamp 1649977179
transform 1 0 30017 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_434
timestamp 1649977179
transform 1 0 29681 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_435
timestamp 1649977179
transform 1 0 29345 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_436
timestamp 1649977179
transform 1 0 34049 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_437
timestamp 1649977179
transform 1 0 33713 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_438
timestamp 1649977179
transform 1 0 33377 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_439
timestamp 1649977179
transform 1 0 29009 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_440
timestamp 1649977179
transform 1 0 33041 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_441
timestamp 1649977179
transform 1 0 18257 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_442
timestamp 1649977179
transform 1 0 18593 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_443
timestamp 1649977179
transform 1 0 17921 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_444
timestamp 1649977179
transform 1 0 20609 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_445
timestamp 1649977179
transform 1 0 20273 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_446
timestamp 1649977179
transform 1 0 19937 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_447
timestamp 1649977179
transform 1 0 25649 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_448
timestamp 1649977179
transform 1 0 25313 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_449
timestamp 1649977179
transform 1 0 24977 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_450
timestamp 1649977179
transform 1 0 24641 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_451
timestamp 1649977179
transform 1 0 24305 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_452
timestamp 1649977179
transform 1 0 23969 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_453
timestamp 1649977179
transform 1 0 23633 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_454
timestamp 1649977179
transform 1 0 23297 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_455
timestamp 1649977179
transform 1 0 22961 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_456
timestamp 1649977179
transform 1 0 19601 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_457
timestamp 1649977179
transform 1 0 22625 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_458
timestamp 1649977179
transform 1 0 19265 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_459
timestamp 1649977179
transform 1 0 22289 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_460
timestamp 1649977179
transform 1 0 17585 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_461
timestamp 1649977179
transform 1 0 21953 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_462
timestamp 1649977179
transform 1 0 21617 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_463
timestamp 1649977179
transform 1 0 21281 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_464
timestamp 1649977179
transform 1 0 18929 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_465
timestamp 1649977179
transform 1 0 20945 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_466
timestamp 1649977179
transform 1 0 9521 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_467
timestamp 1649977179
transform 1 0 8849 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_468
timestamp 1649977179
transform 1 0 13553 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_469
timestamp 1649977179
transform 1 0 10193 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_470
timestamp 1649977179
transform 1 0 13217 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_471
timestamp 1649977179
transform 1 0 12881 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_472
timestamp 1649977179
transform 1 0 12545 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_473
timestamp 1649977179
transform 1 0 12209 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_474
timestamp 1649977179
transform 1 0 11873 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_475
timestamp 1649977179
transform 1 0 9185 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_476
timestamp 1649977179
transform 1 0 9857 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_477
timestamp 1649977179
transform 1 0 11537 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_478
timestamp 1649977179
transform 1 0 11201 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_479
timestamp 1649977179
transform 1 0 10865 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_480
timestamp 1649977179
transform 1 0 10529 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_481
timestamp 1649977179
transform 1 0 16913 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_482
timestamp 1649977179
transform 1 0 16577 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_483
timestamp 1649977179
transform 1 0 16241 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_484
timestamp 1649977179
transform 1 0 15905 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_485
timestamp 1649977179
transform 1 0 15569 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_486
timestamp 1649977179
transform 1 0 15233 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_487
timestamp 1649977179
transform 1 0 14897 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_488
timestamp 1649977179
transform 1 0 14561 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_489
timestamp 1649977179
transform 1 0 14225 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_490
timestamp 1649977179
transform 1 0 13889 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_491
timestamp 1649977179
transform 1 0 5153 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_492
timestamp 1649977179
transform 1 0 7841 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_493
timestamp 1649977179
transform 1 0 4817 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_494
timestamp 1649977179
transform 1 0 7169 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_495
timestamp 1649977179
transform 1 0 8513 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_496
timestamp 1649977179
transform 1 0 5489 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_497
timestamp 1649977179
transform 1 0 6833 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_498
timestamp 1649977179
transform 1 0 6497 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_499
timestamp 1649977179
transform 1 0 6161 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_500
timestamp 1649977179
transform 1 0 5825 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_501
timestamp 1649977179
transform 1 0 8177 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_502
timestamp 1649977179
transform 1 0 7505 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_503
timestamp 1649977179
transform 1 0 4145 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_504
timestamp 1649977179
transform 1 0 3809 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_505
timestamp 1649977179
transform 1 0 3473 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_506
timestamp 1649977179
transform 1 0 3137 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_507
timestamp 1649977179
transform 1 0 2801 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_508
timestamp 1649977179
transform 1 0 2465 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_509
timestamp 1649977179
transform 1 0 2129 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_510
timestamp 1649977179
transform 1 0 1793 0 1 2699
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_511
timestamp 1649977179
transform 1 0 1793 0 1 2363
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_512
timestamp 1649977179
transform 1 0 1793 0 1 2027
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_513
timestamp 1649977179
transform 1 0 1793 0 1 4043
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_514
timestamp 1649977179
transform 1 0 1793 0 1 3707
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_515
timestamp 1649977179
transform 1 0 1793 0 1 3371
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_516
timestamp 1649977179
transform 1 0 1793 0 1 3035
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_517
timestamp 1649977179
transform 1 0 1793 0 1 5051
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_518
timestamp 1649977179
transform 1 0 1793 0 1 4715
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_519
timestamp 1649977179
transform 1 0 1793 0 1 4379
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_520
timestamp 1649977179
transform 1 0 4481 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_521
timestamp 1649977179
transform 1 0 1793 0 1 10427
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_522
timestamp 1649977179
transform 1 0 1793 0 1 10091
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_523
timestamp 1649977179
transform 1 0 1793 0 1 9755
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_524
timestamp 1649977179
transform 1 0 1793 0 1 9419
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_525
timestamp 1649977179
transform 1 0 1793 0 1 9083
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_526
timestamp 1649977179
transform 1 0 1793 0 1 8747
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_527
timestamp 1649977179
transform 1 0 1793 0 1 8411
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_528
timestamp 1649977179
transform 1 0 1793 0 1 8075
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_529
timestamp 1649977179
transform 1 0 1793 0 1 7739
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_530
timestamp 1649977179
transform 1 0 1793 0 1 7403
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_531
timestamp 1649977179
transform 1 0 1793 0 1 7067
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_532
timestamp 1649977179
transform 1 0 1793 0 1 6731
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_533
timestamp 1649977179
transform 1 0 1793 0 1 6395
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_534
timestamp 1649977179
transform 1 0 1793 0 1 6059
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_535
timestamp 1649977179
transform 1 0 1793 0 1 5723
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_536
timestamp 1649977179
transform 1 0 1793 0 1 5387
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_537
timestamp 1649977179
transform 1 0 1793 0 1 13451
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_538
timestamp 1649977179
transform 1 0 1793 0 1 15467
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_539
timestamp 1649977179
transform 1 0 1793 0 1 15131
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_540
timestamp 1649977179
transform 1 0 1793 0 1 11099
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_541
timestamp 1649977179
transform 1 0 1793 0 1 14795
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_542
timestamp 1649977179
transform 1 0 1793 0 1 10763
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_543
timestamp 1649977179
transform 1 0 1793 0 1 14459
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_544
timestamp 1649977179
transform 1 0 1793 0 1 13115
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_545
timestamp 1649977179
transform 1 0 1793 0 1 12779
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_546
timestamp 1649977179
transform 1 0 1793 0 1 12443
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_547
timestamp 1649977179
transform 1 0 1793 0 1 14123
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_548
timestamp 1649977179
transform 1 0 1793 0 1 12107
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_549
timestamp 1649977179
transform 1 0 1793 0 1 11435
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_550
timestamp 1649977179
transform 1 0 1793 0 1 11771
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_551
timestamp 1649977179
transform 1 0 1793 0 1 13787
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_552
timestamp 1649977179
transform 1 0 1793 0 1 15803
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_553
timestamp 1649977179
transform 1 0 1793 0 1 17147
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_554
timestamp 1649977179
transform 1 0 1793 0 1 16811
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_555
timestamp 1649977179
transform 1 0 1793 0 1 16475
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_556
timestamp 1649977179
transform 1 0 1793 0 1 16139
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_557
timestamp 1649977179
transform 1 0 1793 0 1 20843
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_558
timestamp 1649977179
transform 1 0 1793 0 1 20507
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_559
timestamp 1649977179
transform 1 0 1793 0 1 20171
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_560
timestamp 1649977179
transform 1 0 1793 0 1 19835
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_561
timestamp 1649977179
transform 1 0 1793 0 1 19499
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_562
timestamp 1649977179
transform 1 0 1793 0 1 19163
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_563
timestamp 1649977179
transform 1 0 1793 0 1 18827
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_564
timestamp 1649977179
transform 1 0 1793 0 1 18491
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_565
timestamp 1649977179
transform 1 0 1793 0 1 18155
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_566
timestamp 1649977179
transform 1 0 1793 0 1 17819
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_567
timestamp 1649977179
transform 1 0 1793 0 1 17483
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_568
timestamp 1649977179
transform 1 0 17249 0 1 1691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_569
timestamp 1649977179
transform 1 0 1793 0 1 21515
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_570
timestamp 1649977179
transform 1 0 1793 0 1 22523
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_571
timestamp 1649977179
transform 1 0 1793 0 1 24203
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_572
timestamp 1649977179
transform 1 0 1793 0 1 21179
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_573
timestamp 1649977179
transform 1 0 1793 0 1 24875
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_574
timestamp 1649977179
transform 1 0 1793 0 1 22187
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_575
timestamp 1649977179
transform 1 0 1793 0 1 24539
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_576
timestamp 1649977179
transform 1 0 1793 0 1 25883
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_577
timestamp 1649977179
transform 1 0 1793 0 1 25547
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_578
timestamp 1649977179
transform 1 0 1793 0 1 23867
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_579
timestamp 1649977179
transform 1 0 1793 0 1 23531
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_580
timestamp 1649977179
transform 1 0 1793 0 1 23195
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_581
timestamp 1649977179
transform 1 0 1793 0 1 25211
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_582
timestamp 1649977179
transform 1 0 1793 0 1 21851
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_583
timestamp 1649977179
transform 1 0 1793 0 1 22859
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_584
timestamp 1649977179
transform 1 0 1793 0 1 26219
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_585
timestamp 1649977179
transform 1 0 1793 0 1 29915
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_586
timestamp 1649977179
transform 1 0 1793 0 1 30923
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_587
timestamp 1649977179
transform 1 0 1793 0 1 30587
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_588
timestamp 1649977179
transform 1 0 1793 0 1 29579
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_589
timestamp 1649977179
transform 1 0 1793 0 1 29243
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_590
timestamp 1649977179
transform 1 0 1793 0 1 30251
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_591
timestamp 1649977179
transform 1 0 1793 0 1 28907
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_592
timestamp 1649977179
transform 1 0 1793 0 1 28571
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_593
timestamp 1649977179
transform 1 0 1793 0 1 28235
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_594
timestamp 1649977179
transform 1 0 1793 0 1 27899
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_595
timestamp 1649977179
transform 1 0 1793 0 1 27563
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_596
timestamp 1649977179
transform 1 0 1793 0 1 27227
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_597
timestamp 1649977179
transform 1 0 1793 0 1 26891
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_598
timestamp 1649977179
transform 1 0 1793 0 1 26555
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_599
timestamp 1649977179
transform 1 0 1793 0 1 31931
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_600
timestamp 1649977179
transform 1 0 1793 0 1 36299
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_601
timestamp 1649977179
transform 1 0 1793 0 1 35963
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_602
timestamp 1649977179
transform 1 0 1793 0 1 35627
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_603
timestamp 1649977179
transform 1 0 1793 0 1 35291
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_604
timestamp 1649977179
transform 1 0 1793 0 1 34955
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_605
timestamp 1649977179
transform 1 0 1793 0 1 31595
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_606
timestamp 1649977179
transform 1 0 1793 0 1 34619
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_607
timestamp 1649977179
transform 1 0 1793 0 1 34283
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_608
timestamp 1649977179
transform 1 0 1793 0 1 33947
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_609
timestamp 1649977179
transform 1 0 1793 0 1 33611
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_610
timestamp 1649977179
transform 1 0 1793 0 1 33275
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_611
timestamp 1649977179
transform 1 0 1793 0 1 32939
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_612
timestamp 1649977179
transform 1 0 1793 0 1 32603
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_613
timestamp 1649977179
transform 1 0 1793 0 1 32267
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_614
timestamp 1649977179
transform 1 0 1793 0 1 36635
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_615
timestamp 1649977179
transform 1 0 1793 0 1 37307
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_616
timestamp 1649977179
transform 1 0 1793 0 1 41339
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_617
timestamp 1649977179
transform 1 0 1793 0 1 41003
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_618
timestamp 1649977179
transform 1 0 1793 0 1 40667
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_619
timestamp 1649977179
transform 1 0 1793 0 1 40331
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_620
timestamp 1649977179
transform 1 0 1793 0 1 39995
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_621
timestamp 1649977179
transform 1 0 1793 0 1 39659
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_622
timestamp 1649977179
transform 1 0 1793 0 1 39323
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_623
timestamp 1649977179
transform 1 0 1793 0 1 38987
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_624
timestamp 1649977179
transform 1 0 1793 0 1 38651
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_625
timestamp 1649977179
transform 1 0 1793 0 1 38315
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_626
timestamp 1649977179
transform 1 0 1793 0 1 37979
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_627
timestamp 1649977179
transform 1 0 1793 0 1 37643
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_628
timestamp 1649977179
transform 1 0 1793 0 1 36971
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_629
timestamp 1649977179
transform 1 0 1793 0 1 31259
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_630
timestamp 1649977179
transform 1 0 1793 0 1 41675
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_631
timestamp 1649977179
transform 1 0 1793 0 1 45707
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_632
timestamp 1649977179
transform 1 0 1793 0 1 45371
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_633
timestamp 1649977179
transform 1 0 1793 0 1 45035
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_634
timestamp 1649977179
transform 1 0 1793 0 1 44699
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_635
timestamp 1649977179
transform 1 0 1793 0 1 44363
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_636
timestamp 1649977179
transform 1 0 1793 0 1 44027
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_637
timestamp 1649977179
transform 1 0 1793 0 1 43691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_638
timestamp 1649977179
transform 1 0 1793 0 1 43355
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_639
timestamp 1649977179
transform 1 0 1793 0 1 43019
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_640
timestamp 1649977179
transform 1 0 1793 0 1 42683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_641
timestamp 1649977179
transform 1 0 1793 0 1 42347
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_642
timestamp 1649977179
transform 1 0 1793 0 1 46715
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_643
timestamp 1649977179
transform 1 0 1793 0 1 46379
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_644
timestamp 1649977179
transform 1 0 1793 0 1 46043
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_645
timestamp 1649977179
transform 1 0 1793 0 1 42011
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_646
timestamp 1649977179
transform 1 0 1793 0 1 48395
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_647
timestamp 1649977179
transform 1 0 1793 0 1 48059
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_648
timestamp 1649977179
transform 1 0 1793 0 1 51755
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_649
timestamp 1649977179
transform 1 0 1793 0 1 49067
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_650
timestamp 1649977179
transform 1 0 1793 0 1 50411
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_651
timestamp 1649977179
transform 1 0 1793 0 1 47723
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_652
timestamp 1649977179
transform 1 0 1793 0 1 48731
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_653
timestamp 1649977179
transform 1 0 1793 0 1 49403
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_654
timestamp 1649977179
transform 1 0 1793 0 1 51419
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_655
timestamp 1649977179
transform 1 0 1793 0 1 47387
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_656
timestamp 1649977179
transform 1 0 1793 0 1 47051
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_657
timestamp 1649977179
transform 1 0 1793 0 1 51083
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_658
timestamp 1649977179
transform 1 0 1793 0 1 50747
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_659
timestamp 1649977179
transform 1 0 1793 0 1 50075
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_660
timestamp 1649977179
transform 1 0 1793 0 1 49739
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_661
timestamp 1649977179
transform 1 0 1793 0 1 53771
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_662
timestamp 1649977179
transform 1 0 1793 0 1 53435
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_663
timestamp 1649977179
transform 1 0 1793 0 1 53099
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_664
timestamp 1649977179
transform 1 0 1793 0 1 52091
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_665
timestamp 1649977179
transform 1 0 1793 0 1 52763
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_666
timestamp 1649977179
transform 1 0 1793 0 1 52427
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_667
timestamp 1649977179
transform 1 0 1793 0 1 56459
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_668
timestamp 1649977179
transform 1 0 1793 0 1 56123
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_669
timestamp 1649977179
transform 1 0 1793 0 1 55787
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_670
timestamp 1649977179
transform 1 0 1793 0 1 55451
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_671
timestamp 1649977179
transform 1 0 1793 0 1 55115
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_672
timestamp 1649977179
transform 1 0 1793 0 1 54779
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_673
timestamp 1649977179
transform 1 0 1793 0 1 54443
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_674
timestamp 1649977179
transform 1 0 1793 0 1 54107
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_675
timestamp 1649977179
transform 1 0 1793 0 1 56795
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_676
timestamp 1649977179
transform 1 0 1793 0 1 62171
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_677
timestamp 1649977179
transform 1 0 1793 0 1 61835
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_678
timestamp 1649977179
transform 1 0 1793 0 1 61499
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_679
timestamp 1649977179
transform 1 0 1793 0 1 61163
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_680
timestamp 1649977179
transform 1 0 1793 0 1 60827
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_681
timestamp 1649977179
transform 1 0 1793 0 1 60491
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_682
timestamp 1649977179
transform 1 0 1793 0 1 60155
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_683
timestamp 1649977179
transform 1 0 1793 0 1 59819
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_684
timestamp 1649977179
transform 1 0 1793 0 1 59483
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_685
timestamp 1649977179
transform 1 0 1793 0 1 59147
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_686
timestamp 1649977179
transform 1 0 1793 0 1 58811
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_687
timestamp 1649977179
transform 1 0 1793 0 1 58475
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_688
timestamp 1649977179
transform 1 0 1793 0 1 58139
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_689
timestamp 1649977179
transform 1 0 1793 0 1 57803
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_690
timestamp 1649977179
transform 1 0 1793 0 1 57467
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_691
timestamp 1649977179
transform 1 0 1793 0 1 57131
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_692
timestamp 1649977179
transform 1 0 1793 0 1 63179
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_693
timestamp 1649977179
transform 1 0 1793 0 1 62843
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_694
timestamp 1649977179
transform 1 0 1793 0 1 62507
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_695
timestamp 1649977179
transform 1 0 1793 0 1 67211
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_696
timestamp 1649977179
transform 1 0 1793 0 1 66875
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_697
timestamp 1649977179
transform 1 0 1793 0 1 66539
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_698
timestamp 1649977179
transform 1 0 1793 0 1 66203
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_699
timestamp 1649977179
transform 1 0 1793 0 1 65867
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_700
timestamp 1649977179
transform 1 0 1793 0 1 65531
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_701
timestamp 1649977179
transform 1 0 1793 0 1 65195
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_702
timestamp 1649977179
transform 1 0 1793 0 1 64859
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_703
timestamp 1649977179
transform 1 0 1793 0 1 64523
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_704
timestamp 1649977179
transform 1 0 1793 0 1 64187
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_705
timestamp 1649977179
transform 1 0 1793 0 1 63851
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_706
timestamp 1649977179
transform 1 0 1793 0 1 63515
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_707
timestamp 1649977179
transform 1 0 1793 0 1 68219
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_708
timestamp 1649977179
transform 1 0 1793 0 1 67883
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_709
timestamp 1649977179
transform 1 0 1793 0 1 67547
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_710
timestamp 1649977179
transform 1 0 1793 0 1 69227
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_711
timestamp 1649977179
transform 1 0 1793 0 1 68891
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_712
timestamp 1649977179
transform 1 0 1793 0 1 68555
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_713
timestamp 1649977179
transform 1 0 1793 0 1 72587
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_714
timestamp 1649977179
transform 1 0 1793 0 1 72251
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_715
timestamp 1649977179
transform 1 0 1793 0 1 71915
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_716
timestamp 1649977179
transform 1 0 1793 0 1 71579
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_717
timestamp 1649977179
transform 1 0 1793 0 1 71243
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_718
timestamp 1649977179
transform 1 0 1793 0 1 70907
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_719
timestamp 1649977179
transform 1 0 1793 0 1 70571
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_720
timestamp 1649977179
transform 1 0 1793 0 1 70235
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_721
timestamp 1649977179
transform 1 0 1793 0 1 69899
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_722
timestamp 1649977179
transform 1 0 1793 0 1 69563
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_723
timestamp 1649977179
transform 1 0 1793 0 1 72923
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_724
timestamp 1649977179
transform 1 0 1793 0 1 77291
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_725
timestamp 1649977179
transform 1 0 1793 0 1 77627
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_726
timestamp 1649977179
transform 1 0 1793 0 1 76619
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_727
timestamp 1649977179
transform 1 0 1793 0 1 76283
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_728
timestamp 1649977179
transform 1 0 1793 0 1 75947
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_729
timestamp 1649977179
transform 1 0 1793 0 1 76955
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_730
timestamp 1649977179
transform 1 0 1793 0 1 75611
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_731
timestamp 1649977179
transform 1 0 1793 0 1 75275
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_732
timestamp 1649977179
transform 1 0 1793 0 1 74939
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_733
timestamp 1649977179
transform 1 0 1793 0 1 74603
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_734
timestamp 1649977179
transform 1 0 1793 0 1 74267
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_735
timestamp 1649977179
transform 1 0 1793 0 1 73931
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_736
timestamp 1649977179
transform 1 0 1793 0 1 73595
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_737
timestamp 1649977179
transform 1 0 1793 0 1 73259
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_738
timestamp 1649977179
transform 1 0 1793 0 1 78635
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_739
timestamp 1649977179
transform 1 0 1793 0 1 78299
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_740
timestamp 1649977179
transform 1 0 1793 0 1 77963
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_741
timestamp 1649977179
transform 1 0 1793 0 1 80315
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_742
timestamp 1649977179
transform 1 0 1793 0 1 79979
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_743
timestamp 1649977179
transform 1 0 1793 0 1 79643
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_744
timestamp 1649977179
transform 1 0 1793 0 1 79307
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_745
timestamp 1649977179
transform 1 0 1793 0 1 78971
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_746
timestamp 1649977179
transform 1 0 3473 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_747
timestamp 1649977179
transform 1 0 3137 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_748
timestamp 1649977179
transform 1 0 2801 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_749
timestamp 1649977179
transform 1 0 2465 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_750
timestamp 1649977179
transform 1 0 2129 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_751
timestamp 1649977179
transform 1 0 1793 0 1 80987
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_752
timestamp 1649977179
transform 1 0 1793 0 1 80651
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_753
timestamp 1649977179
transform 1 0 4145 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_754
timestamp 1649977179
transform 1 0 3809 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_755
timestamp 1649977179
transform 1 0 8513 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_756
timestamp 1649977179
transform 1 0 8177 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_757
timestamp 1649977179
transform 1 0 7841 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_758
timestamp 1649977179
transform 1 0 7505 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_759
timestamp 1649977179
transform 1 0 7169 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_760
timestamp 1649977179
transform 1 0 6833 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_761
timestamp 1649977179
transform 1 0 6497 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_762
timestamp 1649977179
transform 1 0 6161 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_763
timestamp 1649977179
transform 1 0 5825 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_764
timestamp 1649977179
transform 1 0 5489 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_765
timestamp 1649977179
transform 1 0 5153 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_766
timestamp 1649977179
transform 1 0 4817 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_767
timestamp 1649977179
transform 1 0 4481 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_768
timestamp 1649977179
transform 1 0 8849 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_769
timestamp 1649977179
transform 1 0 16913 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_770
timestamp 1649977179
transform 1 0 16577 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_771
timestamp 1649977179
transform 1 0 16241 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_772
timestamp 1649977179
transform 1 0 15905 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_773
timestamp 1649977179
transform 1 0 15569 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_774
timestamp 1649977179
transform 1 0 15233 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_775
timestamp 1649977179
transform 1 0 14897 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_776
timestamp 1649977179
transform 1 0 14561 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_777
timestamp 1649977179
transform 1 0 14225 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_778
timestamp 1649977179
transform 1 0 13889 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_779
timestamp 1649977179
transform 1 0 13553 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_780
timestamp 1649977179
transform 1 0 13217 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_781
timestamp 1649977179
transform 1 0 12881 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_782
timestamp 1649977179
transform 1 0 12545 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_783
timestamp 1649977179
transform 1 0 12209 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_784
timestamp 1649977179
transform 1 0 11873 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_785
timestamp 1649977179
transform 1 0 11537 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_786
timestamp 1649977179
transform 1 0 11201 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_787
timestamp 1649977179
transform 1 0 10865 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_788
timestamp 1649977179
transform 1 0 10529 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_789
timestamp 1649977179
transform 1 0 10193 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_790
timestamp 1649977179
transform 1 0 9857 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_791
timestamp 1649977179
transform 1 0 9521 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_792
timestamp 1649977179
transform 1 0 9185 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_793
timestamp 1649977179
transform 1 0 24977 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_794
timestamp 1649977179
transform 1 0 24641 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_795
timestamp 1649977179
transform 1 0 24305 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_796
timestamp 1649977179
transform 1 0 23969 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_797
timestamp 1649977179
transform 1 0 23633 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_798
timestamp 1649977179
transform 1 0 23297 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_799
timestamp 1649977179
transform 1 0 22961 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_800
timestamp 1649977179
transform 1 0 22625 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_801
timestamp 1649977179
transform 1 0 22289 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_802
timestamp 1649977179
transform 1 0 21953 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_803
timestamp 1649977179
transform 1 0 21617 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_804
timestamp 1649977179
transform 1 0 21281 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_805
timestamp 1649977179
transform 1 0 20945 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_806
timestamp 1649977179
transform 1 0 20609 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_807
timestamp 1649977179
transform 1 0 20273 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_808
timestamp 1649977179
transform 1 0 19937 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_809
timestamp 1649977179
transform 1 0 19601 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_810
timestamp 1649977179
transform 1 0 19265 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_811
timestamp 1649977179
transform 1 0 18929 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_812
timestamp 1649977179
transform 1 0 18593 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_813
timestamp 1649977179
transform 1 0 18257 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_814
timestamp 1649977179
transform 1 0 17921 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_815
timestamp 1649977179
transform 1 0 17585 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_816
timestamp 1649977179
transform 1 0 25649 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_817
timestamp 1649977179
transform 1 0 25313 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_818
timestamp 1649977179
transform 1 0 34049 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_819
timestamp 1649977179
transform 1 0 33713 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_820
timestamp 1649977179
transform 1 0 33377 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_821
timestamp 1649977179
transform 1 0 33041 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_822
timestamp 1649977179
transform 1 0 32705 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_823
timestamp 1649977179
transform 1 0 32369 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_824
timestamp 1649977179
transform 1 0 32033 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_825
timestamp 1649977179
transform 1 0 31697 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_826
timestamp 1649977179
transform 1 0 31361 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_827
timestamp 1649977179
transform 1 0 31025 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_828
timestamp 1649977179
transform 1 0 30689 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_829
timestamp 1649977179
transform 1 0 30353 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_830
timestamp 1649977179
transform 1 0 30017 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_831
timestamp 1649977179
transform 1 0 29681 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_832
timestamp 1649977179
transform 1 0 29345 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_833
timestamp 1649977179
transform 1 0 29009 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_834
timestamp 1649977179
transform 1 0 28673 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_835
timestamp 1649977179
transform 1 0 28337 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_836
timestamp 1649977179
transform 1 0 28001 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_837
timestamp 1649977179
transform 1 0 27665 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_838
timestamp 1649977179
transform 1 0 27329 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_839
timestamp 1649977179
transform 1 0 26993 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_840
timestamp 1649977179
transform 1 0 26657 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_841
timestamp 1649977179
transform 1 0 26321 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_842
timestamp 1649977179
transform 1 0 25985 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_843
timestamp 1649977179
transform 1 0 17249 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_844
timestamp 1649977179
transform 1 0 37409 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_845
timestamp 1649977179
transform 1 0 37073 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_846
timestamp 1649977179
transform 1 0 36737 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_847
timestamp 1649977179
transform 1 0 36401 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_848
timestamp 1649977179
transform 1 0 36065 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_849
timestamp 1649977179
transform 1 0 35729 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_850
timestamp 1649977179
transform 1 0 35393 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_851
timestamp 1649977179
transform 1 0 35057 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_852
timestamp 1649977179
transform 1 0 34721 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_853
timestamp 1649977179
transform 1 0 34385 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_854
timestamp 1649977179
transform 1 0 42449 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_855
timestamp 1649977179
transform 1 0 42113 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_856
timestamp 1649977179
transform 1 0 41777 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_857
timestamp 1649977179
transform 1 0 41441 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_858
timestamp 1649977179
transform 1 0 41105 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_859
timestamp 1649977179
transform 1 0 40769 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_860
timestamp 1649977179
transform 1 0 40433 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_861
timestamp 1649977179
transform 1 0 40097 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_862
timestamp 1649977179
transform 1 0 39761 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_863
timestamp 1649977179
transform 1 0 39425 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_864
timestamp 1649977179
transform 1 0 39089 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_865
timestamp 1649977179
transform 1 0 38753 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_866
timestamp 1649977179
transform 1 0 38417 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_867
timestamp 1649977179
transform 1 0 38081 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_868
timestamp 1649977179
transform 1 0 37745 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_869
timestamp 1649977179
transform 1 0 46481 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_870
timestamp 1649977179
transform 1 0 46145 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_871
timestamp 1649977179
transform 1 0 45809 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_872
timestamp 1649977179
transform 1 0 45473 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_873
timestamp 1649977179
transform 1 0 45137 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_874
timestamp 1649977179
transform 1 0 44801 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_875
timestamp 1649977179
transform 1 0 44465 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_876
timestamp 1649977179
transform 1 0 44129 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_877
timestamp 1649977179
transform 1 0 43793 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_878
timestamp 1649977179
transform 1 0 43457 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_879
timestamp 1649977179
transform 1 0 43121 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_880
timestamp 1649977179
transform 1 0 51185 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_881
timestamp 1649977179
transform 1 0 50849 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_882
timestamp 1649977179
transform 1 0 50513 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_883
timestamp 1649977179
transform 1 0 50177 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_884
timestamp 1649977179
transform 1 0 49841 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_885
timestamp 1649977179
transform 1 0 49505 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_886
timestamp 1649977179
transform 1 0 49169 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_887
timestamp 1649977179
transform 1 0 48833 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_888
timestamp 1649977179
transform 1 0 48497 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_889
timestamp 1649977179
transform 1 0 48161 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_890
timestamp 1649977179
transform 1 0 47825 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_891
timestamp 1649977179
transform 1 0 47489 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_892
timestamp 1649977179
transform 1 0 47153 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_893
timestamp 1649977179
transform 1 0 46817 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_894
timestamp 1649977179
transform 1 0 42785 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_895
timestamp 1649977179
transform 1 0 58241 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_896
timestamp 1649977179
transform 1 0 57905 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_897
timestamp 1649977179
transform 1 0 57569 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_898
timestamp 1649977179
transform 1 0 57233 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_899
timestamp 1649977179
transform 1 0 56897 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_900
timestamp 1649977179
transform 1 0 56561 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_901
timestamp 1649977179
transform 1 0 56225 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_902
timestamp 1649977179
transform 1 0 55889 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_903
timestamp 1649977179
transform 1 0 55553 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_904
timestamp 1649977179
transform 1 0 55217 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_905
timestamp 1649977179
transform 1 0 54881 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_906
timestamp 1649977179
transform 1 0 54545 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_907
timestamp 1649977179
transform 1 0 54209 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_908
timestamp 1649977179
transform 1 0 53873 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_909
timestamp 1649977179
transform 1 0 53537 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_910
timestamp 1649977179
transform 1 0 53201 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_911
timestamp 1649977179
transform 1 0 52865 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_912
timestamp 1649977179
transform 1 0 52529 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_913
timestamp 1649977179
transform 1 0 52193 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_914
timestamp 1649977179
transform 1 0 51857 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_915
timestamp 1649977179
transform 1 0 51521 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_916
timestamp 1649977179
transform 1 0 59585 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_917
timestamp 1649977179
transform 1 0 59249 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_918
timestamp 1649977179
transform 1 0 58913 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_919
timestamp 1649977179
transform 1 0 58577 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_920
timestamp 1649977179
transform 1 0 67985 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_921
timestamp 1649977179
transform 1 0 67649 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_922
timestamp 1649977179
transform 1 0 67313 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_923
timestamp 1649977179
transform 1 0 66977 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_924
timestamp 1649977179
transform 1 0 66641 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_925
timestamp 1649977179
transform 1 0 66305 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_926
timestamp 1649977179
transform 1 0 65969 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_927
timestamp 1649977179
transform 1 0 65633 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_928
timestamp 1649977179
transform 1 0 65297 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_929
timestamp 1649977179
transform 1 0 64961 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_930
timestamp 1649977179
transform 1 0 64625 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_931
timestamp 1649977179
transform 1 0 64289 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_932
timestamp 1649977179
transform 1 0 63953 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_933
timestamp 1649977179
transform 1 0 63617 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_934
timestamp 1649977179
transform 1 0 63281 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_935
timestamp 1649977179
transform 1 0 62945 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_936
timestamp 1649977179
transform 1 0 62609 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_937
timestamp 1649977179
transform 1 0 62273 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_938
timestamp 1649977179
transform 1 0 61937 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_939
timestamp 1649977179
transform 1 0 61601 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_940
timestamp 1649977179
transform 1 0 61265 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_941
timestamp 1649977179
transform 1 0 60929 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_942
timestamp 1649977179
transform 1 0 60593 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_943
timestamp 1649977179
transform 1 0 60257 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_944
timestamp 1649977179
transform 1 0 59921 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_945
timestamp 1649977179
transform 1 0 134843 0 1 44027
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_946
timestamp 1649977179
transform 1 0 134843 0 1 46043
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_947
timestamp 1649977179
transform 1 0 134843 0 1 43691
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_948
timestamp 1649977179
transform 1 0 134843 0 1 43355
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_949
timestamp 1649977179
transform 1 0 134843 0 1 43019
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_950
timestamp 1649977179
transform 1 0 134843 0 1 44363
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_951
timestamp 1649977179
transform 1 0 134843 0 1 44699
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_952
timestamp 1649977179
transform 1 0 134843 0 1 46715
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_953
timestamp 1649977179
transform 1 0 134843 0 1 42683
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_954
timestamp 1649977179
transform 1 0 134843 0 1 42347
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_955
timestamp 1649977179
transform 1 0 134843 0 1 45371
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_956
timestamp 1649977179
transform 1 0 134843 0 1 45035
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_957
timestamp 1649977179
transform 1 0 134843 0 1 42011
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_958
timestamp 1649977179
transform 1 0 134843 0 1 41675
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_959
timestamp 1649977179
transform 1 0 134843 0 1 46379
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_960
timestamp 1649977179
transform 1 0 134843 0 1 45707
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_961
timestamp 1649977179
transform 1 0 134843 0 1 47051
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_962
timestamp 1649977179
transform 1 0 134843 0 1 49739
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_963
timestamp 1649977179
transform 1 0 134843 0 1 49403
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_964
timestamp 1649977179
transform 1 0 134843 0 1 48395
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_965
timestamp 1649977179
transform 1 0 134843 0 1 47723
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_966
timestamp 1649977179
transform 1 0 134843 0 1 47387
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_967
timestamp 1649977179
transform 1 0 134843 0 1 51755
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_968
timestamp 1649977179
transform 1 0 134843 0 1 48059
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_969
timestamp 1649977179
transform 1 0 134843 0 1 51419
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_970
timestamp 1649977179
transform 1 0 134843 0 1 51083
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_971
timestamp 1649977179
transform 1 0 134843 0 1 50747
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_972
timestamp 1649977179
transform 1 0 134843 0 1 50411
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_973
timestamp 1649977179
transform 1 0 134843 0 1 49067
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_974
timestamp 1649977179
transform 1 0 134843 0 1 50075
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_975
timestamp 1649977179
transform 1 0 134843 0 1 48731
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_976
timestamp 1649977179
transform 1 0 134843 0 1 52427
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_977
timestamp 1649977179
transform 1 0 134843 0 1 56795
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_978
timestamp 1649977179
transform 1 0 134843 0 1 52091
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_979
timestamp 1649977179
transform 1 0 134843 0 1 56459
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_980
timestamp 1649977179
transform 1 0 134843 0 1 56123
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_981
timestamp 1649977179
transform 1 0 134843 0 1 55787
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_982
timestamp 1649977179
transform 1 0 134843 0 1 55451
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_983
timestamp 1649977179
transform 1 0 134843 0 1 55115
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_984
timestamp 1649977179
transform 1 0 134843 0 1 54779
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_985
timestamp 1649977179
transform 1 0 134843 0 1 54443
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_986
timestamp 1649977179
transform 1 0 134843 0 1 54107
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_987
timestamp 1649977179
transform 1 0 134843 0 1 53771
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_988
timestamp 1649977179
transform 1 0 134843 0 1 53435
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_989
timestamp 1649977179
transform 1 0 134843 0 1 53099
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_990
timestamp 1649977179
transform 1 0 134843 0 1 52763
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_991
timestamp 1649977179
transform 1 0 134843 0 1 62171
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_992
timestamp 1649977179
transform 1 0 134843 0 1 61835
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_993
timestamp 1649977179
transform 1 0 134843 0 1 61499
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_994
timestamp 1649977179
transform 1 0 134843 0 1 61163
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_995
timestamp 1649977179
transform 1 0 134843 0 1 60827
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_996
timestamp 1649977179
transform 1 0 134843 0 1 60491
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_997
timestamp 1649977179
transform 1 0 134843 0 1 60155
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_998
timestamp 1649977179
transform 1 0 134843 0 1 59819
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_999
timestamp 1649977179
transform 1 0 134843 0 1 59483
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1000
timestamp 1649977179
transform 1 0 134843 0 1 59147
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1001
timestamp 1649977179
transform 1 0 134843 0 1 58811
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1002
timestamp 1649977179
transform 1 0 134843 0 1 58475
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1003
timestamp 1649977179
transform 1 0 134843 0 1 58139
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1004
timestamp 1649977179
transform 1 0 134843 0 1 57803
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1005
timestamp 1649977179
transform 1 0 134843 0 1 57467
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1006
timestamp 1649977179
transform 1 0 134843 0 1 57131
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1007
timestamp 1649977179
transform 1 0 76049 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1008
timestamp 1649977179
transform 1 0 75713 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1009
timestamp 1649977179
transform 1 0 75377 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1010
timestamp 1649977179
transform 1 0 75041 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1011
timestamp 1649977179
transform 1 0 74705 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1012
timestamp 1649977179
transform 1 0 74369 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1013
timestamp 1649977179
transform 1 0 74033 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1014
timestamp 1649977179
transform 1 0 73697 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1015
timestamp 1649977179
transform 1 0 73361 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1016
timestamp 1649977179
transform 1 0 68657 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1017
timestamp 1649977179
transform 1 0 68321 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1018
timestamp 1649977179
transform 1 0 73025 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1019
timestamp 1649977179
transform 1 0 72689 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1020
timestamp 1649977179
transform 1 0 72353 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1021
timestamp 1649977179
transform 1 0 72017 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1022
timestamp 1649977179
transform 1 0 71681 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1023
timestamp 1649977179
transform 1 0 71345 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1024
timestamp 1649977179
transform 1 0 71009 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1025
timestamp 1649977179
transform 1 0 70673 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1026
timestamp 1649977179
transform 1 0 70337 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1027
timestamp 1649977179
transform 1 0 70001 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1028
timestamp 1649977179
transform 1 0 69665 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1029
timestamp 1649977179
transform 1 0 69329 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1030
timestamp 1649977179
transform 1 0 68993 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1031
timestamp 1649977179
transform 1 0 76721 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1032
timestamp 1649977179
transform 1 0 76385 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1033
timestamp 1649977179
transform 1 0 85121 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1034
timestamp 1649977179
transform 1 0 84785 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1035
timestamp 1649977179
transform 1 0 84449 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1036
timestamp 1649977179
transform 1 0 84113 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1037
timestamp 1649977179
transform 1 0 83777 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1038
timestamp 1649977179
transform 1 0 83441 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1039
timestamp 1649977179
transform 1 0 83105 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1040
timestamp 1649977179
transform 1 0 82769 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1041
timestamp 1649977179
transform 1 0 82433 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1042
timestamp 1649977179
transform 1 0 82097 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1043
timestamp 1649977179
transform 1 0 81761 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1044
timestamp 1649977179
transform 1 0 81425 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1045
timestamp 1649977179
transform 1 0 81089 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1046
timestamp 1649977179
transform 1 0 80753 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1047
timestamp 1649977179
transform 1 0 80417 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1048
timestamp 1649977179
transform 1 0 80081 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1049
timestamp 1649977179
transform 1 0 79745 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1050
timestamp 1649977179
transform 1 0 79409 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1051
timestamp 1649977179
transform 1 0 79073 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1052
timestamp 1649977179
transform 1 0 78737 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1053
timestamp 1649977179
transform 1 0 78401 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1054
timestamp 1649977179
transform 1 0 78065 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1055
timestamp 1649977179
transform 1 0 77729 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1056
timestamp 1649977179
transform 1 0 77393 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1057
timestamp 1649977179
transform 1 0 77057 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1058
timestamp 1649977179
transform 1 0 86129 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1059
timestamp 1649977179
transform 1 0 85793 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1060
timestamp 1649977179
transform 1 0 85457 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1061
timestamp 1649977179
transform 1 0 93521 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1062
timestamp 1649977179
transform 1 0 93185 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1063
timestamp 1649977179
transform 1 0 92849 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1064
timestamp 1649977179
transform 1 0 92513 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1065
timestamp 1649977179
transform 1 0 92177 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1066
timestamp 1649977179
transform 1 0 91841 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1067
timestamp 1649977179
transform 1 0 91505 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1068
timestamp 1649977179
transform 1 0 91169 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1069
timestamp 1649977179
transform 1 0 90833 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1070
timestamp 1649977179
transform 1 0 90497 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1071
timestamp 1649977179
transform 1 0 90161 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1072
timestamp 1649977179
transform 1 0 89825 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1073
timestamp 1649977179
transform 1 0 89489 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1074
timestamp 1649977179
transform 1 0 89153 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1075
timestamp 1649977179
transform 1 0 88817 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1076
timestamp 1649977179
transform 1 0 88481 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1077
timestamp 1649977179
transform 1 0 88145 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1078
timestamp 1649977179
transform 1 0 87809 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1079
timestamp 1649977179
transform 1 0 87473 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1080
timestamp 1649977179
transform 1 0 87137 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1081
timestamp 1649977179
transform 1 0 86801 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1082
timestamp 1649977179
transform 1 0 86465 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1083
timestamp 1649977179
transform 1 0 102257 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1084
timestamp 1649977179
transform 1 0 101921 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1085
timestamp 1649977179
transform 1 0 101585 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1086
timestamp 1649977179
transform 1 0 101249 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1087
timestamp 1649977179
transform 1 0 100913 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1088
timestamp 1649977179
transform 1 0 100577 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1089
timestamp 1649977179
transform 1 0 100241 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1090
timestamp 1649977179
transform 1 0 99905 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1091
timestamp 1649977179
transform 1 0 99569 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1092
timestamp 1649977179
transform 1 0 99233 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1093
timestamp 1649977179
transform 1 0 98897 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1094
timestamp 1649977179
transform 1 0 98561 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1095
timestamp 1649977179
transform 1 0 98225 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1096
timestamp 1649977179
transform 1 0 97889 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1097
timestamp 1649977179
transform 1 0 97553 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1098
timestamp 1649977179
transform 1 0 97217 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1099
timestamp 1649977179
transform 1 0 96881 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1100
timestamp 1649977179
transform 1 0 96545 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1101
timestamp 1649977179
transform 1 0 96209 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1102
timestamp 1649977179
transform 1 0 95873 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1103
timestamp 1649977179
transform 1 0 95537 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1104
timestamp 1649977179
transform 1 0 95201 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1105
timestamp 1649977179
transform 1 0 94865 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1106
timestamp 1649977179
transform 1 0 94529 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1107
timestamp 1649977179
transform 1 0 94193 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1108
timestamp 1649977179
transform 1 0 93857 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1109
timestamp 1649977179
transform 1 0 134843 0 1 63515
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1110
timestamp 1649977179
transform 1 0 134843 0 1 63179
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1111
timestamp 1649977179
transform 1 0 134843 0 1 62843
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1112
timestamp 1649977179
transform 1 0 134843 0 1 62507
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1113
timestamp 1649977179
transform 1 0 134843 0 1 67211
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1114
timestamp 1649977179
transform 1 0 134843 0 1 66875
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1115
timestamp 1649977179
transform 1 0 134843 0 1 66539
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1116
timestamp 1649977179
transform 1 0 134843 0 1 66203
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1117
timestamp 1649977179
transform 1 0 134843 0 1 65867
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1118
timestamp 1649977179
transform 1 0 134843 0 1 65531
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1119
timestamp 1649977179
transform 1 0 134843 0 1 65195
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1120
timestamp 1649977179
transform 1 0 134843 0 1 64859
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1121
timestamp 1649977179
transform 1 0 134843 0 1 64523
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1122
timestamp 1649977179
transform 1 0 134843 0 1 64187
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1123
timestamp 1649977179
transform 1 0 134843 0 1 63851
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1124
timestamp 1649977179
transform 1 0 134843 0 1 67883
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1125
timestamp 1649977179
transform 1 0 134843 0 1 67547
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1126
timestamp 1649977179
transform 1 0 134843 0 1 72587
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1127
timestamp 1649977179
transform 1 0 134843 0 1 72251
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1128
timestamp 1649977179
transform 1 0 134843 0 1 71915
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1129
timestamp 1649977179
transform 1 0 134843 0 1 71579
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1130
timestamp 1649977179
transform 1 0 134843 0 1 71243
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1131
timestamp 1649977179
transform 1 0 134843 0 1 70907
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1132
timestamp 1649977179
transform 1 0 134843 0 1 70571
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1133
timestamp 1649977179
transform 1 0 134843 0 1 70235
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1134
timestamp 1649977179
transform 1 0 134843 0 1 69899
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1135
timestamp 1649977179
transform 1 0 134843 0 1 69563
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1136
timestamp 1649977179
transform 1 0 134843 0 1 69227
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1137
timestamp 1649977179
transform 1 0 134843 0 1 68891
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1138
timestamp 1649977179
transform 1 0 134843 0 1 68555
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1139
timestamp 1649977179
transform 1 0 134843 0 1 68219
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1140
timestamp 1649977179
transform 1 0 102929 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1141
timestamp 1649977179
transform 1 0 102593 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1142
timestamp 1649977179
transform 1 0 106289 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1143
timestamp 1649977179
transform 1 0 105953 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1144
timestamp 1649977179
transform 1 0 105617 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1145
timestamp 1649977179
transform 1 0 105281 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1146
timestamp 1649977179
transform 1 0 104945 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1147
timestamp 1649977179
transform 1 0 104609 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1148
timestamp 1649977179
transform 1 0 104273 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1149
timestamp 1649977179
transform 1 0 103937 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1150
timestamp 1649977179
transform 1 0 103601 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1151
timestamp 1649977179
transform 1 0 103265 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1152
timestamp 1649977179
transform 1 0 110657 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1153
timestamp 1649977179
transform 1 0 110321 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1154
timestamp 1649977179
transform 1 0 109985 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1155
timestamp 1649977179
transform 1 0 109649 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1156
timestamp 1649977179
transform 1 0 109313 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1157
timestamp 1649977179
transform 1 0 108977 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1158
timestamp 1649977179
transform 1 0 108641 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1159
timestamp 1649977179
transform 1 0 108305 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1160
timestamp 1649977179
transform 1 0 107969 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1161
timestamp 1649977179
transform 1 0 107633 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1162
timestamp 1649977179
transform 1 0 107297 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1163
timestamp 1649977179
transform 1 0 106961 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1164
timestamp 1649977179
transform 1 0 106625 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1165
timestamp 1649977179
transform 1 0 119057 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1166
timestamp 1649977179
transform 1 0 118721 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1167
timestamp 1649977179
transform 1 0 118385 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1168
timestamp 1649977179
transform 1 0 118049 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1169
timestamp 1649977179
transform 1 0 117713 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1170
timestamp 1649977179
transform 1 0 117377 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1171
timestamp 1649977179
transform 1 0 117041 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1172
timestamp 1649977179
transform 1 0 116705 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1173
timestamp 1649977179
transform 1 0 116369 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1174
timestamp 1649977179
transform 1 0 116033 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1175
timestamp 1649977179
transform 1 0 115697 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1176
timestamp 1649977179
transform 1 0 115361 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1177
timestamp 1649977179
transform 1 0 115025 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1178
timestamp 1649977179
transform 1 0 114689 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1179
timestamp 1649977179
transform 1 0 114353 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1180
timestamp 1649977179
transform 1 0 114017 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1181
timestamp 1649977179
transform 1 0 113681 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1182
timestamp 1649977179
transform 1 0 113345 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1183
timestamp 1649977179
transform 1 0 113009 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1184
timestamp 1649977179
transform 1 0 112673 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1185
timestamp 1649977179
transform 1 0 112337 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1186
timestamp 1649977179
transform 1 0 112001 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1187
timestamp 1649977179
transform 1 0 111665 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1188
timestamp 1649977179
transform 1 0 111329 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1189
timestamp 1649977179
transform 1 0 110993 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1190
timestamp 1649977179
transform 1 0 134843 0 1 77291
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1191
timestamp 1649977179
transform 1 0 134843 0 1 76955
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1192
timestamp 1649977179
transform 1 0 134843 0 1 76619
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1193
timestamp 1649977179
transform 1 0 134843 0 1 76283
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1194
timestamp 1649977179
transform 1 0 134843 0 1 75947
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1195
timestamp 1649977179
transform 1 0 134843 0 1 75611
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1196
timestamp 1649977179
transform 1 0 134843 0 1 75275
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1197
timestamp 1649977179
transform 1 0 134843 0 1 74939
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1198
timestamp 1649977179
transform 1 0 134843 0 1 74603
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1199
timestamp 1649977179
transform 1 0 134843 0 1 74267
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1200
timestamp 1649977179
transform 1 0 134843 0 1 73931
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1201
timestamp 1649977179
transform 1 0 134843 0 1 73595
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1202
timestamp 1649977179
transform 1 0 134843 0 1 73259
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1203
timestamp 1649977179
transform 1 0 134843 0 1 72923
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1204
timestamp 1649977179
transform 1 0 134843 0 1 77627
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1205
timestamp 1649977179
transform 1 0 126449 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1206
timestamp 1649977179
transform 1 0 126113 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1207
timestamp 1649977179
transform 1 0 125777 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1208
timestamp 1649977179
transform 1 0 125441 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1209
timestamp 1649977179
transform 1 0 125105 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1210
timestamp 1649977179
transform 1 0 124769 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1211
timestamp 1649977179
transform 1 0 124433 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1212
timestamp 1649977179
transform 1 0 124097 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1213
timestamp 1649977179
transform 1 0 123761 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1214
timestamp 1649977179
transform 1 0 123425 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1215
timestamp 1649977179
transform 1 0 123089 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1216
timestamp 1649977179
transform 1 0 122753 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1217
timestamp 1649977179
transform 1 0 122417 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1218
timestamp 1649977179
transform 1 0 122081 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1219
timestamp 1649977179
transform 1 0 121745 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1220
timestamp 1649977179
transform 1 0 121409 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1221
timestamp 1649977179
transform 1 0 121073 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1222
timestamp 1649977179
transform 1 0 120737 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1223
timestamp 1649977179
transform 1 0 120401 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1224
timestamp 1649977179
transform 1 0 120065 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1225
timestamp 1649977179
transform 1 0 119729 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1226
timestamp 1649977179
transform 1 0 119393 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1227
timestamp 1649977179
transform 1 0 127457 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1228
timestamp 1649977179
transform 1 0 127121 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1229
timestamp 1649977179
transform 1 0 126785 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1230
timestamp 1649977179
transform 1 0 134843 0 1 78971
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1231
timestamp 1649977179
transform 1 0 134843 0 1 78635
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1232
timestamp 1649977179
transform 1 0 134843 0 1 78299
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1233
timestamp 1649977179
transform 1 0 134843 0 1 77963
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1234
timestamp 1649977179
transform 1 0 134843 0 1 80315
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1235
timestamp 1649977179
transform 1 0 134843 0 1 79979
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1236
timestamp 1649977179
transform 1 0 134843 0 1 79643
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1237
timestamp 1649977179
transform 1 0 134843 0 1 79307
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1238
timestamp 1649977179
transform 1 0 129809 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1239
timestamp 1649977179
transform 1 0 129473 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1240
timestamp 1649977179
transform 1 0 129137 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1241
timestamp 1649977179
transform 1 0 128801 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1242
timestamp 1649977179
transform 1 0 128465 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1243
timestamp 1649977179
transform 1 0 128129 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1244
timestamp 1649977179
transform 1 0 131825 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1245
timestamp 1649977179
transform 1 0 131489 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1246
timestamp 1649977179
transform 1 0 131153 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1247
timestamp 1649977179
transform 1 0 130817 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1248
timestamp 1649977179
transform 1 0 130481 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1249
timestamp 1649977179
transform 1 0 130145 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1250
timestamp 1649977179
transform 1 0 134843 0 1 80987
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1251
timestamp 1649977179
transform 1 0 134843 0 1 80651
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1252
timestamp 1649977179
transform 1 0 134177 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1253
timestamp 1649977179
transform 1 0 133841 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1254
timestamp 1649977179
transform 1 0 133505 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1255
timestamp 1649977179
transform 1 0 133169 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1256
timestamp 1649977179
transform 1 0 132833 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1257
timestamp 1649977179
transform 1 0 132497 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1258
timestamp 1649977179
transform 1 0 132161 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1259
timestamp 1649977179
transform 1 0 127793 0 1 81440
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_0
timestamp 1649977179
transform 1 0 134840 0 1 2700
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_1
timestamp 1649977179
transform 1 0 134840 0 1 2364
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_2
timestamp 1649977179
transform 1 0 134840 0 1 2028
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_3
timestamp 1649977179
transform 1 0 133166 0 1 1692
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_4
timestamp 1649977179
transform 1 0 131486 0 1 1692
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_5
timestamp 1649977179
transform 1 0 129806 0 1 1692
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_6
timestamp 1649977179
transform 1 0 128126 0 1 1692
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_7
timestamp 1649977179
transform 1 0 134840 0 1 3036
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_8
timestamp 1649977179
transform 1 0 134840 0 1 4044
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_9
timestamp 1649977179
transform 1 0 134840 0 1 3372
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_10
timestamp 1649977179
transform 1 0 134840 0 1 3708
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_11
timestamp 1649977179
transform 1 0 134840 0 1 5052
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_12
timestamp 1649977179
transform 1 0 134840 0 1 4716
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_13
timestamp 1649977179
transform 1 0 134840 0 1 4380
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_14
timestamp 1649977179
transform 1 0 126446 0 1 1692
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_15
timestamp 1649977179
transform 1 0 124766 0 1 1692
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_16
timestamp 1649977179
transform 1 0 123086 0 1 1692
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_17
timestamp 1649977179
transform 1 0 121406 0 1 1692
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_18
timestamp 1649977179
transform 1 0 119726 0 1 1692
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_19
timestamp 1649977179
transform 1 0 134840 0 1 10428
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_20
timestamp 1649977179
transform 1 0 134840 0 1 10092
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_21
timestamp 1649977179
transform 1 0 134840 0 1 9756
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_22
timestamp 1649977179
transform 1 0 134840 0 1 9420
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_23
timestamp 1649977179
transform 1 0 134840 0 1 9084
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_24
timestamp 1649977179
transform 1 0 134840 0 1 8748
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_25
timestamp 1649977179
transform 1 0 134840 0 1 8412
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_26
timestamp 1649977179
transform 1 0 134840 0 1 8076
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_27
timestamp 1649977179
transform 1 0 134840 0 1 7740
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_28
timestamp 1649977179
transform 1 0 134840 0 1 7404
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_29
timestamp 1649977179
transform 1 0 134840 0 1 7068
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_30
timestamp 1649977179
transform 1 0 134840 0 1 6732
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_31
timestamp 1649977179
transform 1 0 134840 0 1 6396
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_32
timestamp 1649977179
transform 1 0 134840 0 1 6060
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_33
timestamp 1649977179
transform 1 0 134840 0 1 5724
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_34
timestamp 1649977179
transform 1 0 134840 0 1 5388
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_35
timestamp 1649977179
transform 1 0 114686 0 1 1692
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_36
timestamp 1649977179
transform 1 0 111326 0 1 1692
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_37
timestamp 1649977179
transform 1 0 113006 0 1 1692
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_38
timestamp 1649977179
transform 1 0 118046 0 1 1692
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_39
timestamp 1649977179
transform 1 0 116366 0 1 1692
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_40
timestamp 1649977179
transform 1 0 102926 0 1 1692
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_41
timestamp 1649977179
transform 1 0 107966 0 1 1692
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_42
timestamp 1649977179
transform 1 0 104606 0 1 1692
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_43
timestamp 1649977179
transform 1 0 106286 0 1 1692
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_44
timestamp 1649977179
transform 1 0 109646 0 1 1692
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_45
timestamp 1649977179
transform 1 0 105990 0 1 13201
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_46
timestamp 1649977179
transform 1 0 103494 0 1 13201
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_47
timestamp 1649977179
transform 1 0 134840 0 1 14796
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_48
timestamp 1649977179
transform 1 0 134840 0 1 14460
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_49
timestamp 1649977179
transform 1 0 134840 0 1 14124
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_50
timestamp 1649977179
transform 1 0 134840 0 1 13788
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_51
timestamp 1649977179
transform 1 0 134840 0 1 13452
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_52
timestamp 1649977179
transform 1 0 134840 0 1 13116
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_53
timestamp 1649977179
transform 1 0 134840 0 1 12780
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_54
timestamp 1649977179
transform 1 0 134840 0 1 12444
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_55
timestamp 1649977179
transform 1 0 134840 0 1 12108
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_56
timestamp 1649977179
transform 1 0 134840 0 1 11772
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_57
timestamp 1649977179
transform 1 0 134840 0 1 11436
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_58
timestamp 1649977179
transform 1 0 134840 0 1 11100
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_59
timestamp 1649977179
transform 1 0 134840 0 1 10764
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_60
timestamp 1649977179
transform 1 0 134840 0 1 15468
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_61
timestamp 1649977179
transform 1 0 134840 0 1 15132
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_62
timestamp 1649977179
transform 1 0 121743 0 1 14793
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_63
timestamp 1649977179
transform 1 0 121663 0 1 13523
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_64
timestamp 1649977179
transform 1 0 121503 0 1 10695
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_65
timestamp 1649977179
transform 1 0 121583 0 1 11965
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_66
timestamp 1649977179
transform 1 0 121823 0 1 16351
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_67
timestamp 1649977179
transform 1 0 121903 0 1 17621
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_68
timestamp 1649977179
transform 1 0 121983 0 1 19179
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_69
timestamp 1649977179
transform 1 0 134840 0 1 20844
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_70
timestamp 1649977179
transform 1 0 134840 0 1 20508
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_71
timestamp 1649977179
transform 1 0 134840 0 1 20172
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_72
timestamp 1649977179
transform 1 0 134840 0 1 19836
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_73
timestamp 1649977179
transform 1 0 134840 0 1 19500
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_74
timestamp 1649977179
transform 1 0 134840 0 1 19164
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_75
timestamp 1649977179
transform 1 0 134840 0 1 18828
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_76
timestamp 1649977179
transform 1 0 134840 0 1 18492
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_77
timestamp 1649977179
transform 1 0 134840 0 1 18156
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_78
timestamp 1649977179
transform 1 0 134840 0 1 17820
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_79
timestamp 1649977179
transform 1 0 134840 0 1 17484
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_80
timestamp 1649977179
transform 1 0 134840 0 1 17148
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_81
timestamp 1649977179
transform 1 0 134840 0 1 16812
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_82
timestamp 1649977179
transform 1 0 134840 0 1 16476
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_83
timestamp 1649977179
transform 1 0 134840 0 1 16140
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_84
timestamp 1649977179
transform 1 0 134840 0 1 15804
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_85
timestamp 1649977179
transform 1 0 94526 0 1 1692
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_86
timestamp 1649977179
transform 1 0 101246 0 1 1692
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_87
timestamp 1649977179
transform 1 0 96206 0 1 1692
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_88
timestamp 1649977179
transform 1 0 97886 0 1 1692
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_89
timestamp 1649977179
transform 1 0 99566 0 1 1692
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_90
timestamp 1649977179
transform 1 0 86126 0 1 1692
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_91
timestamp 1649977179
transform 1 0 92846 0 1 1692
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_92
timestamp 1649977179
transform 1 0 89486 0 1 1692
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_93
timestamp 1649977179
transform 1 0 91166 0 1 1692
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_94
timestamp 1649977179
transform 1 0 87806 0 1 1692
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_95
timestamp 1649977179
transform 1 0 79406 0 1 1692
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_96
timestamp 1649977179
transform 1 0 77726 0 1 1692
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_97
timestamp 1649977179
transform 1 0 84446 0 1 1692
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_98
timestamp 1649977179
transform 1 0 81086 0 1 1692
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_99
timestamp 1649977179
transform 1 0 82766 0 1 1692
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_100
timestamp 1649977179
transform 1 0 74366 0 1 1692
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_101
timestamp 1649977179
transform 1 0 76046 0 1 1692
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_102
timestamp 1649977179
transform 1 0 72686 0 1 1692
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_103
timestamp 1649977179
transform 1 0 71006 0 1 1692
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_104
timestamp 1649977179
transform 1 0 69326 0 1 1692
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_105
timestamp 1649977179
transform 1 0 83526 0 1 13201
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_106
timestamp 1649977179
transform 1 0 81030 0 1 13201
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_107
timestamp 1649977179
transform 1 0 78534 0 1 13201
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_108
timestamp 1649977179
transform 1 0 76038 0 1 13201
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_109
timestamp 1649977179
transform 1 0 73542 0 1 13201
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_110
timestamp 1649977179
transform 1 0 71046 0 1 13201
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_111
timestamp 1649977179
transform 1 0 68550 0 1 13201
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_112
timestamp 1649977179
transform 1 0 100998 0 1 13201
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_113
timestamp 1649977179
transform 1 0 98502 0 1 13201
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_114
timestamp 1649977179
transform 1 0 96006 0 1 13201
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_115
timestamp 1649977179
transform 1 0 93510 0 1 13201
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_116
timestamp 1649977179
transform 1 0 91014 0 1 13201
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_117
timestamp 1649977179
transform 1 0 88518 0 1 13201
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_118
timestamp 1649977179
transform 1 0 86022 0 1 13201
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_119
timestamp 1649977179
transform 1 0 134840 0 1 21180
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_120
timestamp 1649977179
transform 1 0 134840 0 1 22524
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_121
timestamp 1649977179
transform 1 0 134840 0 1 24876
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_122
timestamp 1649977179
transform 1 0 134840 0 1 24540
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_123
timestamp 1649977179
transform 1 0 134840 0 1 24204
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_124
timestamp 1649977179
transform 1 0 134840 0 1 23868
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_125
timestamp 1649977179
transform 1 0 134840 0 1 23532
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_126
timestamp 1649977179
transform 1 0 134840 0 1 25884
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_127
timestamp 1649977179
transform 1 0 134840 0 1 25548
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_128
timestamp 1649977179
transform 1 0 134840 0 1 25212
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_129
timestamp 1649977179
transform 1 0 134840 0 1 23196
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_130
timestamp 1649977179
transform 1 0 134840 0 1 22188
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_131
timestamp 1649977179
transform 1 0 134840 0 1 22860
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_132
timestamp 1649977179
transform 1 0 134840 0 1 21852
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_133
timestamp 1649977179
transform 1 0 134840 0 1 21516
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_134
timestamp 1649977179
transform 1 0 134840 0 1 27228
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_135
timestamp 1649977179
transform 1 0 134840 0 1 26892
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_136
timestamp 1649977179
transform 1 0 134840 0 1 26556
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_137
timestamp 1649977179
transform 1 0 134840 0 1 26220
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_138
timestamp 1649977179
transform 1 0 134840 0 1 30924
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_139
timestamp 1649977179
transform 1 0 134840 0 1 30588
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_140
timestamp 1649977179
transform 1 0 134840 0 1 30252
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_141
timestamp 1649977179
transform 1 0 134840 0 1 29916
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_142
timestamp 1649977179
transform 1 0 134840 0 1 29580
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_143
timestamp 1649977179
transform 1 0 134840 0 1 29244
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_144
timestamp 1649977179
transform 1 0 134840 0 1 28908
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_145
timestamp 1649977179
transform 1 0 134840 0 1 28572
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_146
timestamp 1649977179
transform 1 0 134840 0 1 28236
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_147
timestamp 1649977179
transform 1 0 134840 0 1 27900
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_148
timestamp 1649977179
transform 1 0 134840 0 1 27564
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_149
timestamp 1649977179
transform 1 0 134840 0 1 31596
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_150
timestamp 1649977179
transform 1 0 134840 0 1 36300
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_151
timestamp 1649977179
transform 1 0 134840 0 1 35964
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_152
timestamp 1649977179
transform 1 0 134840 0 1 35628
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_153
timestamp 1649977179
transform 1 0 134840 0 1 35292
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_154
timestamp 1649977179
transform 1 0 134840 0 1 34956
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_155
timestamp 1649977179
transform 1 0 134840 0 1 34620
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_156
timestamp 1649977179
transform 1 0 134840 0 1 34284
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_157
timestamp 1649977179
transform 1 0 134840 0 1 33948
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_158
timestamp 1649977179
transform 1 0 134840 0 1 33612
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_159
timestamp 1649977179
transform 1 0 134840 0 1 33276
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_160
timestamp 1649977179
transform 1 0 134840 0 1 32940
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_161
timestamp 1649977179
transform 1 0 134840 0 1 32604
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_162
timestamp 1649977179
transform 1 0 134840 0 1 32268
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_163
timestamp 1649977179
transform 1 0 134840 0 1 31932
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_164
timestamp 1649977179
transform 1 0 134840 0 1 41340
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_165
timestamp 1649977179
transform 1 0 134840 0 1 41004
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_166
timestamp 1649977179
transform 1 0 134840 0 1 40668
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_167
timestamp 1649977179
transform 1 0 134840 0 1 40332
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_168
timestamp 1649977179
transform 1 0 134840 0 1 39996
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_169
timestamp 1649977179
transform 1 0 134840 0 1 39660
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_170
timestamp 1649977179
transform 1 0 134840 0 1 39324
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_171
timestamp 1649977179
transform 1 0 134840 0 1 38988
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_172
timestamp 1649977179
transform 1 0 134840 0 1 38652
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_173
timestamp 1649977179
transform 1 0 134840 0 1 38316
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_174
timestamp 1649977179
transform 1 0 134840 0 1 37980
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_175
timestamp 1649977179
transform 1 0 134840 0 1 37644
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_176
timestamp 1649977179
transform 1 0 134840 0 1 37308
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_177
timestamp 1649977179
transform 1 0 134840 0 1 36972
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_178
timestamp 1649977179
transform 1 0 134840 0 1 36636
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_179
timestamp 1649977179
transform 1 0 134840 0 1 31260
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_180
timestamp 1649977179
transform 1 0 65966 0 1 1692
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_181
timestamp 1649977179
transform 1 0 67646 0 1 1692
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_182
timestamp 1649977179
transform 1 0 64286 0 1 1692
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_183
timestamp 1649977179
transform 1 0 62606 0 1 1692
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_184
timestamp 1649977179
transform 1 0 60926 0 1 1692
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_185
timestamp 1649977179
transform 1 0 55886 0 1 1692
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_186
timestamp 1649977179
transform 1 0 57566 0 1 1692
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_187
timestamp 1649977179
transform 1 0 54206 0 1 1692
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_188
timestamp 1649977179
transform 1 0 59246 0 1 1692
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_189
timestamp 1649977179
transform 1 0 52526 0 1 1692
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_190
timestamp 1649977179
transform 1 0 44126 0 1 1692
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_191
timestamp 1649977179
transform 1 0 47486 0 1 1692
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_192
timestamp 1649977179
transform 1 0 45806 0 1 1692
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_193
timestamp 1649977179
transform 1 0 50846 0 1 1692
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_194
timestamp 1649977179
transform 1 0 49166 0 1 1692
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_195
timestamp 1649977179
transform 1 0 39086 0 1 1692
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_196
timestamp 1649977179
transform 1 0 37406 0 1 1692
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_197
timestamp 1649977179
transform 1 0 35726 0 1 1692
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_198
timestamp 1649977179
transform 1 0 42446 0 1 1692
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_199
timestamp 1649977179
transform 1 0 40766 0 1 1692
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_200
timestamp 1649977179
transform 1 0 51078 0 1 13201
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_201
timestamp 1649977179
transform 1 0 48582 0 1 13201
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_202
timestamp 1649977179
transform 1 0 46086 0 1 13201
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_203
timestamp 1649977179
transform 1 0 43590 0 1 13201
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_204
timestamp 1649977179
transform 1 0 41094 0 1 13201
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_205
timestamp 1649977179
transform 1 0 38598 0 1 13201
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_206
timestamp 1649977179
transform 1 0 36102 0 1 13201
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_207
timestamp 1649977179
transform 1 0 66054 0 1 13201
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_208
timestamp 1649977179
transform 1 0 63558 0 1 13201
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_209
timestamp 1649977179
transform 1 0 61062 0 1 13201
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_210
timestamp 1649977179
transform 1 0 58566 0 1 13201
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_211
timestamp 1649977179
transform 1 0 56070 0 1 13201
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_212
timestamp 1649977179
transform 1 0 53574 0 1 13201
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_213
timestamp 1649977179
transform 1 0 32366 0 1 1692
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_214
timestamp 1649977179
transform 1 0 27326 0 1 1692
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_215
timestamp 1649977179
transform 1 0 30686 0 1 1692
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_216
timestamp 1649977179
transform 1 0 34046 0 1 1692
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_217
timestamp 1649977179
transform 1 0 29006 0 1 1692
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_218
timestamp 1649977179
transform 1 0 20606 0 1 1692
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_219
timestamp 1649977179
transform 1 0 25646 0 1 1692
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_220
timestamp 1649977179
transform 1 0 23966 0 1 1692
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_221
timestamp 1649977179
transform 1 0 22286 0 1 1692
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_222
timestamp 1649977179
transform 1 0 18926 0 1 1692
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_223
timestamp 1649977179
transform 1 0 8846 0 1 1692
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_224
timestamp 1649977179
transform 1 0 12206 0 1 1692
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_225
timestamp 1649977179
transform 1 0 10526 0 1 1692
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_226
timestamp 1649977179
transform 1 0 15566 0 1 1692
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_227
timestamp 1649977179
transform 1 0 13886 0 1 1692
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_228
timestamp 1649977179
transform 1 0 5486 0 1 1692
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_229
timestamp 1649977179
transform 1 0 7166 0 1 1692
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_230
timestamp 1649977179
transform 1 0 3806 0 1 1692
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_231
timestamp 1649977179
transform 1 0 2126 0 1 1692
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_232
timestamp 1649977179
transform 1 0 1790 0 1 2700
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_233
timestamp 1649977179
transform 1 0 1790 0 1 2364
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_234
timestamp 1649977179
transform 1 0 1790 0 1 2028
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_235
timestamp 1649977179
transform 1 0 1790 0 1 4044
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_236
timestamp 1649977179
transform 1 0 1790 0 1 3708
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_237
timestamp 1649977179
transform 1 0 1790 0 1 3372
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_238
timestamp 1649977179
transform 1 0 1790 0 1 3036
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_239
timestamp 1649977179
transform 1 0 1790 0 1 5052
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_240
timestamp 1649977179
transform 1 0 1790 0 1 4716
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_241
timestamp 1649977179
transform 1 0 1790 0 1 4380
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_242
timestamp 1649977179
transform 1 0 1790 0 1 10428
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_243
timestamp 1649977179
transform 1 0 1790 0 1 10092
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_244
timestamp 1649977179
transform 1 0 1790 0 1 9756
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_245
timestamp 1649977179
transform 1 0 1790 0 1 9420
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_246
timestamp 1649977179
transform 1 0 1790 0 1 9084
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_247
timestamp 1649977179
transform 1 0 1790 0 1 8748
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_248
timestamp 1649977179
transform 1 0 1790 0 1 8412
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_249
timestamp 1649977179
transform 1 0 1790 0 1 8076
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_250
timestamp 1649977179
transform 1 0 1790 0 1 7740
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_251
timestamp 1649977179
transform 1 0 1790 0 1 7404
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_252
timestamp 1649977179
transform 1 0 1790 0 1 7068
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_253
timestamp 1649977179
transform 1 0 1790 0 1 6732
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_254
timestamp 1649977179
transform 1 0 1790 0 1 6396
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_255
timestamp 1649977179
transform 1 0 1790 0 1 6060
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_256
timestamp 1649977179
transform 1 0 1790 0 1 5724
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_257
timestamp 1649977179
transform 1 0 1790 0 1 5388
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_258
timestamp 1649977179
transform 1 0 1790 0 1 13452
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_259
timestamp 1649977179
transform 1 0 1790 0 1 13116
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_260
timestamp 1649977179
transform 1 0 1790 0 1 15468
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_261
timestamp 1649977179
transform 1 0 1790 0 1 15132
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_262
timestamp 1649977179
transform 1 0 1790 0 1 14796
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_263
timestamp 1649977179
transform 1 0 1790 0 1 11100
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_264
timestamp 1649977179
transform 1 0 1790 0 1 10764
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_265
timestamp 1649977179
transform 1 0 1790 0 1 14460
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_266
timestamp 1649977179
transform 1 0 1790 0 1 14124
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_267
timestamp 1649977179
transform 1 0 1790 0 1 12780
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_268
timestamp 1649977179
transform 1 0 1790 0 1 12444
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_269
timestamp 1649977179
transform 1 0 1790 0 1 12108
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_270
timestamp 1649977179
transform 1 0 1790 0 1 13788
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_271
timestamp 1649977179
transform 1 0 1790 0 1 11772
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_272
timestamp 1649977179
transform 1 0 1790 0 1 11436
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_273
timestamp 1649977179
transform 1 0 1790 0 1 15804
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_274
timestamp 1649977179
transform 1 0 1790 0 1 16812
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_275
timestamp 1649977179
transform 1 0 1790 0 1 16476
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_276
timestamp 1649977179
transform 1 0 1790 0 1 16140
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_277
timestamp 1649977179
transform 1 0 1790 0 1 20844
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_278
timestamp 1649977179
transform 1 0 1790 0 1 20508
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_279
timestamp 1649977179
transform 1 0 1790 0 1 20172
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_280
timestamp 1649977179
transform 1 0 1790 0 1 19836
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_281
timestamp 1649977179
transform 1 0 1790 0 1 19500
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_282
timestamp 1649977179
transform 1 0 1790 0 1 19164
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_283
timestamp 1649977179
transform 1 0 1790 0 1 18828
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_284
timestamp 1649977179
transform 1 0 1790 0 1 18492
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_285
timestamp 1649977179
transform 1 0 1790 0 1 18156
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_286
timestamp 1649977179
transform 1 0 1790 0 1 17820
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_287
timestamp 1649977179
transform 1 0 1790 0 1 17484
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_288
timestamp 1649977179
transform 1 0 1790 0 1 17148
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_289
timestamp 1649977179
transform 1 0 33606 0 1 13201
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_290
timestamp 1649977179
transform 1 0 31110 0 1 13201
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_291
timestamp 1649977179
transform 1 0 28614 0 1 13201
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_292
timestamp 1649977179
transform 1 0 17246 0 1 1692
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_293
timestamp 1649977179
transform 1 0 1790 0 1 22524
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_294
timestamp 1649977179
transform 1 0 1790 0 1 24204
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_295
timestamp 1649977179
transform 1 0 1790 0 1 21180
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_296
timestamp 1649977179
transform 1 0 1790 0 1 24876
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_297
timestamp 1649977179
transform 1 0 1790 0 1 24540
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_298
timestamp 1649977179
transform 1 0 1790 0 1 22188
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_299
timestamp 1649977179
transform 1 0 1790 0 1 25884
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_300
timestamp 1649977179
transform 1 0 1790 0 1 25548
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_301
timestamp 1649977179
transform 1 0 1790 0 1 25212
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_302
timestamp 1649977179
transform 1 0 1790 0 1 23868
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_303
timestamp 1649977179
transform 1 0 1790 0 1 23532
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_304
timestamp 1649977179
transform 1 0 1790 0 1 23196
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_305
timestamp 1649977179
transform 1 0 1790 0 1 21852
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_306
timestamp 1649977179
transform 1 0 1790 0 1 22860
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_307
timestamp 1649977179
transform 1 0 1790 0 1 21516
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_308
timestamp 1649977179
transform 1 0 1790 0 1 29916
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_309
timestamp 1649977179
transform 1 0 1790 0 1 29580
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_310
timestamp 1649977179
transform 1 0 1790 0 1 30924
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_311
timestamp 1649977179
transform 1 0 1790 0 1 30588
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_312
timestamp 1649977179
transform 1 0 1790 0 1 29244
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_313
timestamp 1649977179
transform 1 0 1790 0 1 30252
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_314
timestamp 1649977179
transform 1 0 1790 0 1 28908
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_315
timestamp 1649977179
transform 1 0 1790 0 1 28572
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_316
timestamp 1649977179
transform 1 0 1790 0 1 28236
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_317
timestamp 1649977179
transform 1 0 1790 0 1 27900
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_318
timestamp 1649977179
transform 1 0 1790 0 1 27564
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_319
timestamp 1649977179
transform 1 0 1790 0 1 27228
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_320
timestamp 1649977179
transform 1 0 1790 0 1 26892
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_321
timestamp 1649977179
transform 1 0 1790 0 1 26556
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_322
timestamp 1649977179
transform 1 0 1790 0 1 26220
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_323
timestamp 1649977179
transform 1 0 14943 0 1 29907
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_324
timestamp 1649977179
transform 1 0 14863 0 1 28349
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_325
timestamp 1649977179
transform 1 0 15023 0 1 31177
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_326
timestamp 1649977179
transform 1 0 15103 0 1 32735
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_327
timestamp 1649977179
transform 1 0 15263 0 1 35563
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_328
timestamp 1649977179
transform 1 0 15183 0 1 34005
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_329
timestamp 1649977179
transform 1 0 1790 0 1 32268
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_330
timestamp 1649977179
transform 1 0 1790 0 1 36300
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_331
timestamp 1649977179
transform 1 0 1790 0 1 35964
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_332
timestamp 1649977179
transform 1 0 1790 0 1 35628
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_333
timestamp 1649977179
transform 1 0 1790 0 1 35292
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_334
timestamp 1649977179
transform 1 0 1790 0 1 34956
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_335
timestamp 1649977179
transform 1 0 1790 0 1 31596
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_336
timestamp 1649977179
transform 1 0 1790 0 1 31932
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_337
timestamp 1649977179
transform 1 0 1790 0 1 34620
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_338
timestamp 1649977179
transform 1 0 1790 0 1 34284
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_339
timestamp 1649977179
transform 1 0 1790 0 1 33948
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_340
timestamp 1649977179
transform 1 0 1790 0 1 33612
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_341
timestamp 1649977179
transform 1 0 1790 0 1 33276
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_342
timestamp 1649977179
transform 1 0 1790 0 1 32940
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_343
timestamp 1649977179
transform 1 0 1790 0 1 32604
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_344
timestamp 1649977179
transform 1 0 1790 0 1 36636
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_345
timestamp 1649977179
transform 1 0 1790 0 1 36972
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_346
timestamp 1649977179
transform 1 0 1790 0 1 41340
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_347
timestamp 1649977179
transform 1 0 1790 0 1 41004
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_348
timestamp 1649977179
transform 1 0 1790 0 1 40668
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_349
timestamp 1649977179
transform 1 0 1790 0 1 40332
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_350
timestamp 1649977179
transform 1 0 1790 0 1 39996
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_351
timestamp 1649977179
transform 1 0 1790 0 1 39660
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_352
timestamp 1649977179
transform 1 0 1790 0 1 39324
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_353
timestamp 1649977179
transform 1 0 1790 0 1 38988
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_354
timestamp 1649977179
transform 1 0 1790 0 1 38652
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_355
timestamp 1649977179
transform 1 0 1790 0 1 38316
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_356
timestamp 1649977179
transform 1 0 1790 0 1 37980
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_357
timestamp 1649977179
transform 1 0 1790 0 1 37644
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_358
timestamp 1649977179
transform 1 0 1790 0 1 37308
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_359
timestamp 1649977179
transform 1 0 15343 0 1 36833
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_360
timestamp 1649977179
transform 1 0 1790 0 1 31260
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_361
timestamp 1649977179
transform 1 0 1790 0 1 45708
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_362
timestamp 1649977179
transform 1 0 1790 0 1 45372
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_363
timestamp 1649977179
transform 1 0 1790 0 1 45036
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_364
timestamp 1649977179
transform 1 0 1790 0 1 44700
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_365
timestamp 1649977179
transform 1 0 1790 0 1 44364
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_366
timestamp 1649977179
transform 1 0 1790 0 1 44028
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_367
timestamp 1649977179
transform 1 0 1790 0 1 43692
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_368
timestamp 1649977179
transform 1 0 1790 0 1 43356
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_369
timestamp 1649977179
transform 1 0 1790 0 1 43020
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_370
timestamp 1649977179
transform 1 0 1790 0 1 42684
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_371
timestamp 1649977179
transform 1 0 1790 0 1 42348
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_372
timestamp 1649977179
transform 1 0 1790 0 1 46716
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_373
timestamp 1649977179
transform 1 0 1790 0 1 42012
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_374
timestamp 1649977179
transform 1 0 1790 0 1 46380
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_375
timestamp 1649977179
transform 1 0 1790 0 1 46044
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_376
timestamp 1649977179
transform 1 0 1790 0 1 41676
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_377
timestamp 1649977179
transform 1 0 1790 0 1 48396
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_378
timestamp 1649977179
transform 1 0 1790 0 1 48060
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_379
timestamp 1649977179
transform 1 0 1790 0 1 47724
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_380
timestamp 1649977179
transform 1 0 1790 0 1 50412
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_381
timestamp 1649977179
transform 1 0 1790 0 1 50076
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_382
timestamp 1649977179
transform 1 0 1790 0 1 48732
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_383
timestamp 1649977179
transform 1 0 1790 0 1 49404
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_384
timestamp 1649977179
transform 1 0 1790 0 1 51420
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_385
timestamp 1649977179
transform 1 0 1790 0 1 47388
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_386
timestamp 1649977179
transform 1 0 1790 0 1 47052
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_387
timestamp 1649977179
transform 1 0 1790 0 1 51756
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_388
timestamp 1649977179
transform 1 0 1790 0 1 51084
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_389
timestamp 1649977179
transform 1 0 1790 0 1 49068
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_390
timestamp 1649977179
transform 1 0 1790 0 1 50748
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_391
timestamp 1649977179
transform 1 0 1790 0 1 49740
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_392
timestamp 1649977179
transform 1 0 1790 0 1 53772
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_393
timestamp 1649977179
transform 1 0 1790 0 1 53436
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_394
timestamp 1649977179
transform 1 0 1790 0 1 53100
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_395
timestamp 1649977179
transform 1 0 1790 0 1 52092
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_396
timestamp 1649977179
transform 1 0 1790 0 1 52428
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_397
timestamp 1649977179
transform 1 0 1790 0 1 52764
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_398
timestamp 1649977179
transform 1 0 1790 0 1 56460
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_399
timestamp 1649977179
transform 1 0 1790 0 1 56124
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_400
timestamp 1649977179
transform 1 0 1790 0 1 55788
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_401
timestamp 1649977179
transform 1 0 1790 0 1 55452
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_402
timestamp 1649977179
transform 1 0 1790 0 1 55116
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_403
timestamp 1649977179
transform 1 0 1790 0 1 54780
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_404
timestamp 1649977179
transform 1 0 1790 0 1 54444
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_405
timestamp 1649977179
transform 1 0 1790 0 1 54108
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_406
timestamp 1649977179
transform 1 0 1790 0 1 56796
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_407
timestamp 1649977179
transform 1 0 1790 0 1 62172
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_408
timestamp 1649977179
transform 1 0 1790 0 1 61836
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_409
timestamp 1649977179
transform 1 0 1790 0 1 61500
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_410
timestamp 1649977179
transform 1 0 1790 0 1 61164
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_411
timestamp 1649977179
transform 1 0 1790 0 1 60828
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_412
timestamp 1649977179
transform 1 0 1790 0 1 60492
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_413
timestamp 1649977179
transform 1 0 1790 0 1 60156
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_414
timestamp 1649977179
transform 1 0 1790 0 1 59820
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_415
timestamp 1649977179
transform 1 0 1790 0 1 59484
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_416
timestamp 1649977179
transform 1 0 1790 0 1 59148
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_417
timestamp 1649977179
transform 1 0 1790 0 1 58812
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_418
timestamp 1649977179
transform 1 0 1790 0 1 58476
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_419
timestamp 1649977179
transform 1 0 1790 0 1 58140
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_420
timestamp 1649977179
transform 1 0 1790 0 1 57804
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_421
timestamp 1649977179
transform 1 0 1790 0 1 57468
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_422
timestamp 1649977179
transform 1 0 1790 0 1 57132
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_423
timestamp 1649977179
transform 1 0 1790 0 1 63180
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_424
timestamp 1649977179
transform 1 0 1790 0 1 62844
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_425
timestamp 1649977179
transform 1 0 1790 0 1 62508
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_426
timestamp 1649977179
transform 1 0 1790 0 1 67212
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_427
timestamp 1649977179
transform 1 0 1790 0 1 66876
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_428
timestamp 1649977179
transform 1 0 1790 0 1 66540
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_429
timestamp 1649977179
transform 1 0 1790 0 1 66204
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_430
timestamp 1649977179
transform 1 0 1790 0 1 65868
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_431
timestamp 1649977179
transform 1 0 1790 0 1 65532
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_432
timestamp 1649977179
transform 1 0 1790 0 1 65196
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_433
timestamp 1649977179
transform 1 0 1790 0 1 64860
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_434
timestamp 1649977179
transform 1 0 1790 0 1 64524
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_435
timestamp 1649977179
transform 1 0 1790 0 1 64188
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_436
timestamp 1649977179
transform 1 0 1790 0 1 63852
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_437
timestamp 1649977179
transform 1 0 1790 0 1 63516
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_438
timestamp 1649977179
transform 1 0 1790 0 1 68220
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_439
timestamp 1649977179
transform 1 0 1790 0 1 67884
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_440
timestamp 1649977179
transform 1 0 1790 0 1 67548
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_441
timestamp 1649977179
transform 1 0 1790 0 1 68892
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_442
timestamp 1649977179
transform 1 0 1790 0 1 68556
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_443
timestamp 1649977179
transform 1 0 1790 0 1 72588
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_444
timestamp 1649977179
transform 1 0 1790 0 1 72252
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_445
timestamp 1649977179
transform 1 0 1790 0 1 71916
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_446
timestamp 1649977179
transform 1 0 1790 0 1 71580
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_447
timestamp 1649977179
transform 1 0 1790 0 1 71244
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_448
timestamp 1649977179
transform 1 0 1790 0 1 70908
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_449
timestamp 1649977179
transform 1 0 1790 0 1 70572
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_450
timestamp 1649977179
transform 1 0 1790 0 1 70236
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_451
timestamp 1649977179
transform 1 0 1790 0 1 69228
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_452
timestamp 1649977179
transform 1 0 1790 0 1 69900
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_453
timestamp 1649977179
transform 1 0 1790 0 1 69564
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_454
timestamp 1649977179
transform 1 0 1790 0 1 72924
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_455
timestamp 1649977179
transform 1 0 1790 0 1 77292
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_456
timestamp 1649977179
transform 1 0 1790 0 1 77628
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_457
timestamp 1649977179
transform 1 0 1790 0 1 76620
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_458
timestamp 1649977179
transform 1 0 1790 0 1 76284
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_459
timestamp 1649977179
transform 1 0 1790 0 1 75948
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_460
timestamp 1649977179
transform 1 0 1790 0 1 76956
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_461
timestamp 1649977179
transform 1 0 1790 0 1 75612
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_462
timestamp 1649977179
transform 1 0 1790 0 1 75276
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_463
timestamp 1649977179
transform 1 0 1790 0 1 74940
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_464
timestamp 1649977179
transform 1 0 1790 0 1 74604
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_465
timestamp 1649977179
transform 1 0 1790 0 1 74268
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_466
timestamp 1649977179
transform 1 0 1790 0 1 73932
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_467
timestamp 1649977179
transform 1 0 1790 0 1 73596
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_468
timestamp 1649977179
transform 1 0 1790 0 1 73260
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_469
timestamp 1649977179
transform 1 0 1790 0 1 78636
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_470
timestamp 1649977179
transform 1 0 1790 0 1 78300
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_471
timestamp 1649977179
transform 1 0 1790 0 1 77964
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_472
timestamp 1649977179
transform 1 0 1790 0 1 80316
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_473
timestamp 1649977179
transform 1 0 1790 0 1 79980
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_474
timestamp 1649977179
transform 1 0 1790 0 1 79644
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_475
timestamp 1649977179
transform 1 0 1790 0 1 79308
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_476
timestamp 1649977179
transform 1 0 1790 0 1 78972
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_477
timestamp 1649977179
transform 1 0 2126 0 1 81441
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_478
timestamp 1649977179
transform 1 0 1790 0 1 80988
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_479
timestamp 1649977179
transform 1 0 1790 0 1 80652
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_480
timestamp 1649977179
transform 1 0 3806 0 1 81441
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_481
timestamp 1649977179
transform 1 0 7166 0 1 81441
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_482
timestamp 1649977179
transform 1 0 5486 0 1 81441
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_483
timestamp 1649977179
transform 1 0 15566 0 1 81441
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_484
timestamp 1649977179
transform 1 0 13886 0 1 81441
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_485
timestamp 1649977179
transform 1 0 12206 0 1 81441
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_486
timestamp 1649977179
transform 1 0 10526 0 1 81441
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_487
timestamp 1649977179
transform 1 0 8846 0 1 81441
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_488
timestamp 1649977179
transform 1 0 31110 0 1 76987
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_489
timestamp 1649977179
transform 1 0 28614 0 1 76987
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_490
timestamp 1649977179
transform 1 0 33606 0 1 76987
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_491
timestamp 1649977179
transform 1 0 23966 0 1 81441
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_492
timestamp 1649977179
transform 1 0 22286 0 1 81441
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_493
timestamp 1649977179
transform 1 0 20606 0 1 81441
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_494
timestamp 1649977179
transform 1 0 18926 0 1 81441
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_495
timestamp 1649977179
transform 1 0 25646 0 1 81441
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_496
timestamp 1649977179
transform 1 0 34046 0 1 81441
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_497
timestamp 1649977179
transform 1 0 32366 0 1 81441
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_498
timestamp 1649977179
transform 1 0 30686 0 1 81441
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_499
timestamp 1649977179
transform 1 0 29006 0 1 81441
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_500
timestamp 1649977179
transform 1 0 27326 0 1 81441
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_501
timestamp 1649977179
transform 1 0 17246 0 1 81441
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_502
timestamp 1649977179
transform 1 0 51078 0 1 76987
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_503
timestamp 1649977179
transform 1 0 48582 0 1 76987
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_504
timestamp 1649977179
transform 1 0 46086 0 1 76987
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_505
timestamp 1649977179
transform 1 0 43590 0 1 76987
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_506
timestamp 1649977179
transform 1 0 36102 0 1 76987
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_507
timestamp 1649977179
transform 1 0 41094 0 1 76987
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_508
timestamp 1649977179
transform 1 0 38598 0 1 76987
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_509
timestamp 1649977179
transform 1 0 35726 0 1 81441
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_510
timestamp 1649977179
transform 1 0 42446 0 1 81441
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_511
timestamp 1649977179
transform 1 0 40766 0 1 81441
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_512
timestamp 1649977179
transform 1 0 39086 0 1 81441
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_513
timestamp 1649977179
transform 1 0 37406 0 1 81441
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_514
timestamp 1649977179
transform 1 0 45806 0 1 81441
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_515
timestamp 1649977179
transform 1 0 44126 0 1 81441
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_516
timestamp 1649977179
transform 1 0 50846 0 1 81441
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_517
timestamp 1649977179
transform 1 0 49166 0 1 81441
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_518
timestamp 1649977179
transform 1 0 47486 0 1 81441
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_519
timestamp 1649977179
transform 1 0 66054 0 1 76987
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_520
timestamp 1649977179
transform 1 0 63558 0 1 76987
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_521
timestamp 1649977179
transform 1 0 61062 0 1 76987
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_522
timestamp 1649977179
transform 1 0 58566 0 1 76987
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_523
timestamp 1649977179
transform 1 0 56070 0 1 76987
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_524
timestamp 1649977179
transform 1 0 53574 0 1 76987
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_525
timestamp 1649977179
transform 1 0 57566 0 1 81441
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_526
timestamp 1649977179
transform 1 0 55886 0 1 81441
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_527
timestamp 1649977179
transform 1 0 54206 0 1 81441
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_528
timestamp 1649977179
transform 1 0 52526 0 1 81441
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_529
timestamp 1649977179
transform 1 0 59246 0 1 81441
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_530
timestamp 1649977179
transform 1 0 67646 0 1 81441
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_531
timestamp 1649977179
transform 1 0 65966 0 1 81441
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_532
timestamp 1649977179
transform 1 0 64286 0 1 81441
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_533
timestamp 1649977179
transform 1 0 62606 0 1 81441
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_534
timestamp 1649977179
transform 1 0 60926 0 1 81441
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_535
timestamp 1649977179
transform 1 0 134840 0 1 44700
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_536
timestamp 1649977179
transform 1 0 134840 0 1 44364
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_537
timestamp 1649977179
transform 1 0 134840 0 1 43692
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_538
timestamp 1649977179
transform 1 0 134840 0 1 43356
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_539
timestamp 1649977179
transform 1 0 134840 0 1 43020
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_540
timestamp 1649977179
transform 1 0 134840 0 1 46716
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_541
timestamp 1649977179
transform 1 0 134840 0 1 42684
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_542
timestamp 1649977179
transform 1 0 134840 0 1 42348
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_543
timestamp 1649977179
transform 1 0 134840 0 1 42012
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_544
timestamp 1649977179
transform 1 0 134840 0 1 45036
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_545
timestamp 1649977179
transform 1 0 134840 0 1 41676
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_546
timestamp 1649977179
transform 1 0 134840 0 1 45708
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_547
timestamp 1649977179
transform 1 0 134840 0 1 46380
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_548
timestamp 1649977179
transform 1 0 134840 0 1 46044
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_549
timestamp 1649977179
transform 1 0 134840 0 1 45372
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_550
timestamp 1649977179
transform 1 0 134840 0 1 44028
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_551
timestamp 1649977179
transform 1 0 134840 0 1 47724
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_552
timestamp 1649977179
transform 1 0 134840 0 1 47052
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_553
timestamp 1649977179
transform 1 0 134840 0 1 48396
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_554
timestamp 1649977179
transform 1 0 134840 0 1 49740
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_555
timestamp 1649977179
transform 1 0 134840 0 1 49404
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_556
timestamp 1649977179
transform 1 0 134840 0 1 47388
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_557
timestamp 1649977179
transform 1 0 134840 0 1 51756
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_558
timestamp 1649977179
transform 1 0 134840 0 1 48060
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_559
timestamp 1649977179
transform 1 0 134840 0 1 51420
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_560
timestamp 1649977179
transform 1 0 134840 0 1 51084
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_561
timestamp 1649977179
transform 1 0 134840 0 1 50076
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_562
timestamp 1649977179
transform 1 0 134840 0 1 49068
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_563
timestamp 1649977179
transform 1 0 134840 0 1 50748
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_564
timestamp 1649977179
transform 1 0 134840 0 1 50412
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_565
timestamp 1649977179
transform 1 0 134840 0 1 48732
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_566
timestamp 1649977179
transform 1 0 134840 0 1 52092
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_567
timestamp 1649977179
transform 1 0 134840 0 1 56796
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_568
timestamp 1649977179
transform 1 0 134840 0 1 56460
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_569
timestamp 1649977179
transform 1 0 134840 0 1 56124
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_570
timestamp 1649977179
transform 1 0 134840 0 1 55788
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_571
timestamp 1649977179
transform 1 0 134840 0 1 55452
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_572
timestamp 1649977179
transform 1 0 134840 0 1 55116
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_573
timestamp 1649977179
transform 1 0 134840 0 1 54780
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_574
timestamp 1649977179
transform 1 0 134840 0 1 54444
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_575
timestamp 1649977179
transform 1 0 134840 0 1 54108
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_576
timestamp 1649977179
transform 1 0 134840 0 1 53772
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_577
timestamp 1649977179
transform 1 0 134840 0 1 53436
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_578
timestamp 1649977179
transform 1 0 134840 0 1 53100
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_579
timestamp 1649977179
transform 1 0 134840 0 1 52764
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_580
timestamp 1649977179
transform 1 0 134840 0 1 52428
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_581
timestamp 1649977179
transform 1 0 134840 0 1 62172
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_582
timestamp 1649977179
transform 1 0 134840 0 1 61836
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_583
timestamp 1649977179
transform 1 0 134840 0 1 61500
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_584
timestamp 1649977179
transform 1 0 134840 0 1 61164
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_585
timestamp 1649977179
transform 1 0 134840 0 1 60828
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_586
timestamp 1649977179
transform 1 0 134840 0 1 60492
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_587
timestamp 1649977179
transform 1 0 134840 0 1 60156
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_588
timestamp 1649977179
transform 1 0 134840 0 1 59820
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_589
timestamp 1649977179
transform 1 0 134840 0 1 59484
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_590
timestamp 1649977179
transform 1 0 134840 0 1 59148
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_591
timestamp 1649977179
transform 1 0 134840 0 1 58812
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_592
timestamp 1649977179
transform 1 0 134840 0 1 58476
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_593
timestamp 1649977179
transform 1 0 134840 0 1 58140
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_594
timestamp 1649977179
transform 1 0 134840 0 1 57804
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_595
timestamp 1649977179
transform 1 0 134840 0 1 57468
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_596
timestamp 1649977179
transform 1 0 134840 0 1 57132
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_597
timestamp 1649977179
transform 1 0 81030 0 1 76987
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_598
timestamp 1649977179
transform 1 0 78534 0 1 76987
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_599
timestamp 1649977179
transform 1 0 83526 0 1 76987
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_600
timestamp 1649977179
transform 1 0 71046 0 1 76987
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_601
timestamp 1649977179
transform 1 0 68550 0 1 76987
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_602
timestamp 1649977179
transform 1 0 76038 0 1 76987
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_603
timestamp 1649977179
transform 1 0 73542 0 1 76987
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_604
timestamp 1649977179
transform 1 0 76046 0 1 81441
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_605
timestamp 1649977179
transform 1 0 74366 0 1 81441
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_606
timestamp 1649977179
transform 1 0 72686 0 1 81441
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_607
timestamp 1649977179
transform 1 0 71006 0 1 81441
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_608
timestamp 1649977179
transform 1 0 69326 0 1 81441
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_609
timestamp 1649977179
transform 1 0 84446 0 1 81441
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_610
timestamp 1649977179
transform 1 0 82766 0 1 81441
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_611
timestamp 1649977179
transform 1 0 81086 0 1 81441
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_612
timestamp 1649977179
transform 1 0 79406 0 1 81441
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_613
timestamp 1649977179
transform 1 0 77726 0 1 81441
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_614
timestamp 1649977179
transform 1 0 96006 0 1 76987
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_615
timestamp 1649977179
transform 1 0 100998 0 1 76987
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_616
timestamp 1649977179
transform 1 0 98502 0 1 76987
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_617
timestamp 1649977179
transform 1 0 93510 0 1 76987
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_618
timestamp 1649977179
transform 1 0 91014 0 1 76987
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_619
timestamp 1649977179
transform 1 0 88518 0 1 76987
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_620
timestamp 1649977179
transform 1 0 86022 0 1 76987
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_621
timestamp 1649977179
transform 1 0 86126 0 1 81441
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_622
timestamp 1649977179
transform 1 0 92846 0 1 81441
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_623
timestamp 1649977179
transform 1 0 91166 0 1 81441
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_624
timestamp 1649977179
transform 1 0 89486 0 1 81441
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_625
timestamp 1649977179
transform 1 0 87806 0 1 81441
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_626
timestamp 1649977179
transform 1 0 101246 0 1 81441
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_627
timestamp 1649977179
transform 1 0 99566 0 1 81441
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_628
timestamp 1649977179
transform 1 0 97886 0 1 81441
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_629
timestamp 1649977179
transform 1 0 96206 0 1 81441
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_630
timestamp 1649977179
transform 1 0 94526 0 1 81441
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_631
timestamp 1649977179
transform 1 0 134840 0 1 63516
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_632
timestamp 1649977179
transform 1 0 134840 0 1 63180
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_633
timestamp 1649977179
transform 1 0 134840 0 1 62844
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_634
timestamp 1649977179
transform 1 0 134840 0 1 62508
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_635
timestamp 1649977179
transform 1 0 134840 0 1 67212
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_636
timestamp 1649977179
transform 1 0 134840 0 1 66876
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_637
timestamp 1649977179
transform 1 0 134840 0 1 66540
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_638
timestamp 1649977179
transform 1 0 134840 0 1 66204
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_639
timestamp 1649977179
transform 1 0 134840 0 1 65868
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_640
timestamp 1649977179
transform 1 0 134840 0 1 65532
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_641
timestamp 1649977179
transform 1 0 134840 0 1 65196
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_642
timestamp 1649977179
transform 1 0 134840 0 1 64860
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_643
timestamp 1649977179
transform 1 0 134840 0 1 64524
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_644
timestamp 1649977179
transform 1 0 134840 0 1 64188
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_645
timestamp 1649977179
transform 1 0 134840 0 1 63852
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_646
timestamp 1649977179
transform 1 0 134840 0 1 67884
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_647
timestamp 1649977179
transform 1 0 134840 0 1 67548
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_648
timestamp 1649977179
transform 1 0 134840 0 1 72588
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_649
timestamp 1649977179
transform 1 0 134840 0 1 72252
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_650
timestamp 1649977179
transform 1 0 134840 0 1 71916
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_651
timestamp 1649977179
transform 1 0 134840 0 1 71580
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_652
timestamp 1649977179
transform 1 0 134840 0 1 71244
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_653
timestamp 1649977179
transform 1 0 134840 0 1 70908
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_654
timestamp 1649977179
transform 1 0 134840 0 1 70572
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_655
timestamp 1649977179
transform 1 0 134840 0 1 70236
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_656
timestamp 1649977179
transform 1 0 134840 0 1 69900
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_657
timestamp 1649977179
transform 1 0 134840 0 1 69564
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_658
timestamp 1649977179
transform 1 0 134840 0 1 69228
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_659
timestamp 1649977179
transform 1 0 134840 0 1 68892
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_660
timestamp 1649977179
transform 1 0 134840 0 1 68556
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_661
timestamp 1649977179
transform 1 0 134840 0 1 68220
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_662
timestamp 1649977179
transform 1 0 103494 0 1 76987
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_663
timestamp 1649977179
transform 1 0 105990 0 1 76987
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_664
timestamp 1649977179
transform 1 0 106286 0 1 81441
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_665
timestamp 1649977179
transform 1 0 104606 0 1 81441
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_666
timestamp 1649977179
transform 1 0 102926 0 1 81441
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_667
timestamp 1649977179
transform 1 0 109646 0 1 81441
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_668
timestamp 1649977179
transform 1 0 107966 0 1 81441
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_669
timestamp 1649977179
transform 1 0 118046 0 1 81441
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_670
timestamp 1649977179
transform 1 0 116366 0 1 81441
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_671
timestamp 1649977179
transform 1 0 114686 0 1 81441
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_672
timestamp 1649977179
transform 1 0 113006 0 1 81441
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_673
timestamp 1649977179
transform 1 0 111326 0 1 81441
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_674
timestamp 1649977179
transform 1 0 134840 0 1 76956
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_675
timestamp 1649977179
transform 1 0 134840 0 1 76620
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_676
timestamp 1649977179
transform 1 0 134840 0 1 76284
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_677
timestamp 1649977179
transform 1 0 134840 0 1 75948
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_678
timestamp 1649977179
transform 1 0 134840 0 1 75612
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_679
timestamp 1649977179
transform 1 0 134840 0 1 75276
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_680
timestamp 1649977179
transform 1 0 134840 0 1 74940
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_681
timestamp 1649977179
transform 1 0 134840 0 1 74604
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_682
timestamp 1649977179
transform 1 0 134840 0 1 74268
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_683
timestamp 1649977179
transform 1 0 134840 0 1 73932
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_684
timestamp 1649977179
transform 1 0 134840 0 1 73596
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_685
timestamp 1649977179
transform 1 0 134840 0 1 73260
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_686
timestamp 1649977179
transform 1 0 134840 0 1 72924
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_687
timestamp 1649977179
transform 1 0 134840 0 1 77628
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_688
timestamp 1649977179
transform 1 0 134840 0 1 77292
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_689
timestamp 1649977179
transform 1 0 126446 0 1 81441
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_690
timestamp 1649977179
transform 1 0 124766 0 1 81441
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_691
timestamp 1649977179
transform 1 0 123086 0 1 81441
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_692
timestamp 1649977179
transform 1 0 121406 0 1 81441
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_693
timestamp 1649977179
transform 1 0 119726 0 1 81441
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_694
timestamp 1649977179
transform 1 0 134840 0 1 78972
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_695
timestamp 1649977179
transform 1 0 134840 0 1 78636
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_696
timestamp 1649977179
transform 1 0 134840 0 1 78300
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_697
timestamp 1649977179
transform 1 0 134840 0 1 77964
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_698
timestamp 1649977179
transform 1 0 134840 0 1 80316
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_699
timestamp 1649977179
transform 1 0 134840 0 1 79980
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_700
timestamp 1649977179
transform 1 0 134840 0 1 79644
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_701
timestamp 1649977179
transform 1 0 134840 0 1 79308
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_702
timestamp 1649977179
transform 1 0 129806 0 1 81441
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_703
timestamp 1649977179
transform 1 0 128126 0 1 81441
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_704
timestamp 1649977179
transform 1 0 131486 0 1 81441
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_705
timestamp 1649977179
transform 1 0 134840 0 1 80988
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_706
timestamp 1649977179
transform 1 0 134840 0 1 80652
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_707
timestamp 1649977179
transform 1 0 133166 0 1 81441
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_32  sky130_sram_2kbyte_1rw1r_32x512_8_contact_32_0
timestamp 1649977179
transform 1 0 122183 0 1 19501
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_32  sky130_sram_2kbyte_1rw1r_32x512_8_contact_32_1
timestamp 1649977179
transform 1 0 14745 0 1 2667
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_32  sky130_sram_2kbyte_1rw1r_32x512_8_contact_32_2
timestamp 1649977179
transform 1 0 14745 0 1 28017
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_32  sky130_sram_2kbyte_1rw1r_32x512_8_contact_32_3
timestamp 1649977179
transform 1 0 122183 0 1 80456
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_0
timestamp 1649977179
transform 1 0 133144 0 1 1229
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1
timestamp 1649977179
transform 1 0 133144 0 1 1637
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2
timestamp 1649977179
transform 1 0 135320 0 1 2045
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3
timestamp 1649977179
transform 1 0 131512 0 1 1229
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_4
timestamp 1649977179
transform 1 0 131512 0 1 1637
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_5
timestamp 1649977179
transform 1 0 129744 0 1 1229
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_6
timestamp 1649977179
transform 1 0 129744 0 1 1637
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_7
timestamp 1649977179
transform 1 0 127976 0 1 1229
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_8
timestamp 1649977179
transform 1 0 127976 0 1 1637
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_9
timestamp 1649977179
transform 1 0 135320 0 1 3677
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_10
timestamp 1649977179
transform 1 0 135320 0 1 5309
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_11
timestamp 1649977179
transform 1 0 119816 0 1 1637
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_12
timestamp 1649977179
transform 1 0 126344 0 1 1229
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_13
timestamp 1649977179
transform 1 0 126344 0 1 1637
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_14
timestamp 1649977179
transform 1 0 124712 0 1 1229
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_15
timestamp 1649977179
transform 1 0 124712 0 1 1637
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_16
timestamp 1649977179
transform 1 0 123080 0 1 1229
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_17
timestamp 1649977179
transform 1 0 123080 0 1 1637
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_18
timestamp 1649977179
transform 1 0 121312 0 1 1229
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_19
timestamp 1649977179
transform 1 0 121312 0 1 1637
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_20
timestamp 1649977179
transform 1 0 119816 0 1 1229
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_21
timestamp 1649977179
transform 1 0 122944 0 1 9933
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_22
timestamp 1649977179
transform 1 0 135320 0 1 7077
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_23
timestamp 1649977179
transform 1 0 135320 0 1 8709
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_24
timestamp 1649977179
transform 1 0 135320 0 1 10341
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_25
timestamp 1649977179
transform 1 0 111248 0 1 1229
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_26
timestamp 1649977179
transform 1 0 111248 0 1 1637
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_27
timestamp 1649977179
transform 1 0 116280 0 1 1229
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_28
timestamp 1649977179
transform 1 0 116280 0 1 1637
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_29
timestamp 1649977179
transform 1 0 118048 0 1 1229
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_30
timestamp 1649977179
transform 1 0 118048 0 1 1637
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_31
timestamp 1649977179
transform 1 0 114784 0 1 1229
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_32
timestamp 1649977179
transform 1 0 114784 0 1 1637
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_33
timestamp 1649977179
transform 1 0 113016 0 1 1229
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_34
timestamp 1649977179
transform 1 0 113016 0 1 1637
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_35
timestamp 1649977179
transform 1 0 102816 0 1 1637
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_36
timestamp 1649977179
transform 1 0 106216 0 1 1229
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_37
timestamp 1649977179
transform 1 0 106216 0 1 1637
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_38
timestamp 1649977179
transform 1 0 109752 0 1 1229
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_39
timestamp 1649977179
transform 1 0 109752 0 1 1637
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_40
timestamp 1649977179
transform 1 0 107848 0 1 1229
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_41
timestamp 1649977179
transform 1 0 107848 0 1 1637
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_42
timestamp 1649977179
transform 1 0 102816 0 1 1229
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_43
timestamp 1649977179
transform 1 0 104584 0 1 1229
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_44
timestamp 1649977179
transform 1 0 104584 0 1 1637
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_45
timestamp 1649977179
transform 1 0 108392 0 1 9525
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_46
timestamp 1649977179
transform 1 0 103768 0 1 12517
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_47
timestamp 1649977179
transform 1 0 103768 0 1 11701
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_48
timestamp 1649977179
transform 1 0 103768 0 1 12245
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_49
timestamp 1649977179
transform 1 0 116008 0 1 20269
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_50
timestamp 1649977179
transform 1 0 116008 0 1 20541
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_51
timestamp 1649977179
transform 1 0 116008 0 1 20677
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_52
timestamp 1649977179
transform 1 0 107168 0 1 19181
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_53
timestamp 1649977179
transform 1 0 118592 0 1 20269
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_54
timestamp 1649977179
transform 1 0 114648 0 1 20541
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_55
timestamp 1649977179
transform 1 0 114648 0 1 20269
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_56
timestamp 1649977179
transform 1 0 115192 0 1 20677
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_57
timestamp 1649977179
transform 1 0 106352 0 1 13605
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_58
timestamp 1649977179
transform 1 0 106352 0 1 14285
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_59
timestamp 1649977179
transform 1 0 102408 0 1 19181
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_60
timestamp 1649977179
transform 1 0 108256 0 1 11021
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_61
timestamp 1649977179
transform 1 0 106352 0 1 13469
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_62
timestamp 1649977179
transform 1 0 106352 0 1 11973
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_63
timestamp 1649977179
transform 1 0 106216 0 1 11021
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_64
timestamp 1649977179
transform 1 0 106216 0 1 11837
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_65
timestamp 1649977179
transform 1 0 102408 0 1 18773
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_66
timestamp 1649977179
transform 1 0 119000 0 1 20269
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_67
timestamp 1649977179
transform 1 0 105944 0 1 13061
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_68
timestamp 1649977179
transform 1 0 103360 0 1 13061
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_69
timestamp 1649977179
transform 1 0 118184 0 1 20269
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_70
timestamp 1649977179
transform 1 0 115328 0 1 20677
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_71
timestamp 1649977179
transform 1 0 115464 0 1 20269
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_72
timestamp 1649977179
transform 1 0 109616 0 1 19725
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_73
timestamp 1649977179
transform 1 0 105808 0 1 19181
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_74
timestamp 1649977179
transform 1 0 105808 0 1 18773
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_75
timestamp 1649977179
transform 1 0 105536 0 1 18773
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_76
timestamp 1649977179
transform 1 0 105536 0 1 19181
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_77
timestamp 1649977179
transform 1 0 109616 0 1 19997
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_78
timestamp 1649977179
transform 1 0 103496 0 1 14285
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_79
timestamp 1649977179
transform 1 0 104856 0 1 19181
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_80
timestamp 1649977179
transform 1 0 104856 0 1 18773
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_81
timestamp 1649977179
transform 1 0 103496 0 1 13605
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_82
timestamp 1649977179
transform 1 0 106352 0 1 17005
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_83
timestamp 1649977179
transform 1 0 114648 0 1 20677
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_84
timestamp 1649977179
transform 1 0 104312 0 1 18773
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_85
timestamp 1649977179
transform 1 0 104312 0 1 19181
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_86
timestamp 1649977179
transform 1 0 115464 0 1 20541
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_87
timestamp 1649977179
transform 1 0 106352 0 1 15101
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_88
timestamp 1649977179
transform 1 0 103768 0 1 13605
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_89
timestamp 1649977179
transform 1 0 103768 0 1 14285
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_90
timestamp 1649977179
transform 1 0 103632 0 1 13605
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_91
timestamp 1649977179
transform 1 0 103632 0 1 11973
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_92
timestamp 1649977179
transform 1 0 103632 0 1 11021
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_93
timestamp 1649977179
transform 1 0 103632 0 1 11837
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_94
timestamp 1649977179
transform 1 0 115056 0 1 20541
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_95
timestamp 1649977179
transform 1 0 117640 0 1 20269
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_96
timestamp 1649977179
transform 1 0 115056 0 1 20269
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_97
timestamp 1649977179
transform 1 0 103088 0 1 18773
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_98
timestamp 1649977179
transform 1 0 114240 0 1 20677
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_99
timestamp 1649977179
transform 1 0 106488 0 1 15101
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_100
timestamp 1649977179
transform 1 0 106488 0 1 13197
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_101
timestamp 1649977179
transform 1 0 106488 0 1 13061
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_102
timestamp 1649977179
transform 1 0 106488 0 1 12517
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_103
timestamp 1649977179
transform 1 0 106080 0 1 11701
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_104
timestamp 1649977179
transform 1 0 106080 0 1 12245
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_105
timestamp 1649977179
transform 1 0 108528 0 1 19181
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_106
timestamp 1649977179
transform 1 0 108528 0 1 18773
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_107
timestamp 1649977179
transform 1 0 103088 0 1 19181
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_108
timestamp 1649977179
transform 1 0 114240 0 1 20541
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_109
timestamp 1649977179
transform 1 0 108392 0 1 11293
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_110
timestamp 1649977179
transform 1 0 104040 0 1 17005
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_111
timestamp 1649977179
transform 1 0 114240 0 1 20269
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_112
timestamp 1649977179
transform 1 0 104040 0 1 15101
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_113
timestamp 1649977179
transform 1 0 107304 0 1 19181
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_114
timestamp 1649977179
transform 1 0 103904 0 1 15101
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_115
timestamp 1649977179
transform 1 0 103904 0 1 13061
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_116
timestamp 1649977179
transform 1 0 107304 0 1 18773
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_117
timestamp 1649977179
transform 1 0 107168 0 1 18773
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_118
timestamp 1649977179
transform 1 0 103768 0 1 13061
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_119
timestamp 1649977179
transform 1 0 135320 0 1 13877
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_120
timestamp 1649977179
transform 1 0 135320 0 1 15373
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_121
timestamp 1649977179
transform 1 0 135320 0 1 12245
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_122
timestamp 1649977179
transform 1 0 122808 0 1 14013
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_123
timestamp 1649977179
transform 1 0 122808 0 1 11429
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_124
timestamp 1649977179
transform 1 0 122808 0 1 14285
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_125
timestamp 1649977179
transform 1 0 122944 0 1 15509
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_126
timestamp 1649977179
transform 1 0 122944 0 1 12789
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_127
timestamp 1649977179
transform 1 0 122944 0 1 15645
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_128
timestamp 1649977179
transform 1 0 123216 0 1 11837
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_129
timestamp 1649977179
transform 1 0 123352 0 1 10749
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_130
timestamp 1649977179
transform 1 0 122944 0 1 12653
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_131
timestamp 1649977179
transform 1 0 122808 0 1 19725
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_132
timestamp 1649977179
transform 1 0 122808 0 1 17005
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_133
timestamp 1649977179
transform 1 0 122808 0 1 16869
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_134
timestamp 1649977179
transform 1 0 122808 0 1 19861
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_135
timestamp 1649977179
transform 1 0 122808 0 1 20133
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_136
timestamp 1649977179
transform 1 0 122944 0 1 18365
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_137
timestamp 1649977179
transform 1 0 119952 0 1 18501
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_138
timestamp 1649977179
transform 1 0 119952 0 1 20133
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_139
timestamp 1649977179
transform 1 0 135320 0 1 18909
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_140
timestamp 1649977179
transform 1 0 135320 0 1 20541
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_141
timestamp 1649977179
transform 1 0 135320 0 1 17141
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_142
timestamp 1649977179
transform 1 0 108256 0 1 10613
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_143
timestamp 1649977179
transform 1 0 97784 0 1 1637
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_144
timestamp 1649977179
transform 1 0 97784 0 1 1229
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_145
timestamp 1649977179
transform 1 0 101320 0 1 1229
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_146
timestamp 1649977179
transform 1 0 101320 0 1 1637
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_147
timestamp 1649977179
transform 1 0 99552 0 1 1229
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_148
timestamp 1649977179
transform 1 0 99552 0 1 1637
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_149
timestamp 1649977179
transform 1 0 96152 0 1 1637
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_150
timestamp 1649977179
transform 1 0 94384 0 1 1229
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_151
timestamp 1649977179
transform 1 0 96152 0 1 1229
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_152
timestamp 1649977179
transform 1 0 94384 0 1 1637
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_153
timestamp 1649977179
transform 1 0 92752 0 1 1229
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_154
timestamp 1649977179
transform 1 0 92752 0 1 1637
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_155
timestamp 1649977179
transform 1 0 91256 0 1 1229
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_156
timestamp 1649977179
transform 1 0 91256 0 1 1637
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_157
timestamp 1649977179
transform 1 0 89352 0 1 1229
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_158
timestamp 1649977179
transform 1 0 89352 0 1 1637
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_159
timestamp 1649977179
transform 1 0 87720 0 1 1229
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_160
timestamp 1649977179
transform 1 0 87720 0 1 1637
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_161
timestamp 1649977179
transform 1 0 86224 0 1 1229
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_162
timestamp 1649977179
transform 1 0 86224 0 1 1637
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_163
timestamp 1649977179
transform 1 0 81056 0 1 1229
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_164
timestamp 1649977179
transform 1 0 81056 0 1 1637
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_165
timestamp 1649977179
transform 1 0 82824 0 1 1229
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_166
timestamp 1649977179
transform 1 0 82824 0 1 1637
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_167
timestamp 1649977179
transform 1 0 79288 0 1 1229
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_168
timestamp 1649977179
transform 1 0 79288 0 1 1637
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_169
timestamp 1649977179
transform 1 0 84320 0 1 1229
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_170
timestamp 1649977179
transform 1 0 84320 0 1 1637
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_171
timestamp 1649977179
transform 1 0 77656 0 1 1229
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_172
timestamp 1649977179
transform 1 0 77656 0 1 1637
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_173
timestamp 1649977179
transform 1 0 76160 0 1 1229
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_174
timestamp 1649977179
transform 1 0 76160 0 1 1637
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_175
timestamp 1649977179
transform 1 0 74256 0 1 1229
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_176
timestamp 1649977179
transform 1 0 74256 0 1 1637
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_177
timestamp 1649977179
transform 1 0 72760 0 1 1229
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_178
timestamp 1649977179
transform 1 0 72760 0 1 1637
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_179
timestamp 1649977179
transform 1 0 70856 0 1 1229
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_180
timestamp 1649977179
transform 1 0 70856 0 1 1637
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_181
timestamp 1649977179
transform 1 0 69224 0 1 1229
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_182
timestamp 1649977179
transform 1 0 69224 0 1 1637
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_183
timestamp 1649977179
transform 1 0 78608 0 1 11701
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_184
timestamp 1649977179
transform 1 0 78608 0 1 12245
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_185
timestamp 1649977179
transform 1 0 81464 0 1 13197
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_186
timestamp 1649977179
transform 1 0 83504 0 1 13061
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_187
timestamp 1649977179
transform 1 0 83912 0 1 15101
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_188
timestamp 1649977179
transform 1 0 80920 0 1 13061
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_189
timestamp 1649977179
transform 1 0 84048 0 1 15101
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_190
timestamp 1649977179
transform 1 0 84048 0 1 13197
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_191
timestamp 1649977179
transform 1 0 78880 0 1 13605
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_192
timestamp 1649977179
transform 1 0 78880 0 1 14285
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_193
timestamp 1649977179
transform 1 0 78880 0 1 13469
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_194
timestamp 1649977179
transform 1 0 78880 0 1 11973
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_195
timestamp 1649977179
transform 1 0 78744 0 1 11021
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_196
timestamp 1649977179
transform 1 0 78744 0 1 11837
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_197
timestamp 1649977179
transform 1 0 83776 0 1 13061
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_198
timestamp 1649977179
transform 1 0 83776 0 1 12517
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_199
timestamp 1649977179
transform 1 0 84048 0 1 11701
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_200
timestamp 1649977179
transform 1 0 83640 0 1 13605
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_201
timestamp 1649977179
transform 1 0 83640 0 1 14285
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_202
timestamp 1649977179
transform 1 0 83912 0 1 13469
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_203
timestamp 1649977179
transform 1 0 83912 0 1 11973
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_204
timestamp 1649977179
transform 1 0 83776 0 1 11021
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_205
timestamp 1649977179
transform 1 0 81464 0 1 13061
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_206
timestamp 1649977179
transform 1 0 81464 0 1 12517
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_207
timestamp 1649977179
transform 1 0 81056 0 1 11701
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_208
timestamp 1649977179
transform 1 0 81056 0 1 12245
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_209
timestamp 1649977179
transform 1 0 83776 0 1 11837
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_210
timestamp 1649977179
transform 1 0 84048 0 1 12245
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_211
timestamp 1649977179
transform 1 0 78880 0 1 15101
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_212
timestamp 1649977179
transform 1 0 79016 0 1 15101
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_213
timestamp 1649977179
transform 1 0 79016 0 1 13197
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_214
timestamp 1649977179
transform 1 0 78472 0 1 13061
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_215
timestamp 1649977179
transform 1 0 81600 0 1 15101
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_216
timestamp 1649977179
transform 1 0 81464 0 1 15101
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_217
timestamp 1649977179
transform 1 0 81328 0 1 13605
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_218
timestamp 1649977179
transform 1 0 81328 0 1 14285
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_219
timestamp 1649977179
transform 1 0 81328 0 1 13469
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_220
timestamp 1649977179
transform 1 0 81328 0 1 11973
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_221
timestamp 1649977179
transform 1 0 81192 0 1 11021
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_222
timestamp 1649977179
transform 1 0 81192 0 1 11837
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_223
timestamp 1649977179
transform 1 0 79016 0 1 13061
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_224
timestamp 1649977179
transform 1 0 79016 0 1 12517
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_225
timestamp 1649977179
transform 1 0 73984 0 1 12517
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_226
timestamp 1649977179
transform 1 0 73304 0 1 12245
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_227
timestamp 1649977179
transform 1 0 73304 0 1 11429
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_228
timestamp 1649977179
transform 1 0 75888 0 1 13061
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_229
timestamp 1649977179
transform 1 0 76432 0 1 11973
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_230
timestamp 1649977179
transform 1 0 71400 0 1 15101
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_231
timestamp 1649977179
transform 1 0 71536 0 1 15101
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_232
timestamp 1649977179
transform 1 0 71536 0 1 13197
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_233
timestamp 1649977179
transform 1 0 73440 0 1 13061
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_234
timestamp 1649977179
transform 1 0 71536 0 1 13061
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_235
timestamp 1649977179
transform 1 0 71536 0 1 12517
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_236
timestamp 1649977179
transform 1 0 71536 0 1 11701
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_237
timestamp 1649977179
transform 1 0 71536 0 1 12245
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_238
timestamp 1649977179
transform 1 0 76296 0 1 11021
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_239
timestamp 1649977179
transform 1 0 69088 0 1 15101
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_240
timestamp 1649977179
transform 1 0 68952 0 1 15101
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_241
timestamp 1649977179
transform 1 0 68952 0 1 13061
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_242
timestamp 1649977179
transform 1 0 68816 0 1 13061
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_243
timestamp 1649977179
transform 1 0 68816 0 1 12517
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_244
timestamp 1649977179
transform 1 0 68544 0 1 11701
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_245
timestamp 1649977179
transform 1 0 68544 0 1 12245
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_246
timestamp 1649977179
transform 1 0 70992 0 1 13061
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_247
timestamp 1649977179
transform 1 0 73984 0 1 13197
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_248
timestamp 1649977179
transform 1 0 76296 0 1 11837
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_249
timestamp 1649977179
transform 1 0 73984 0 1 13061
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_250
timestamp 1649977179
transform 1 0 71264 0 1 14285
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_251
timestamp 1649977179
transform 1 0 76432 0 1 15101
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_252
timestamp 1649977179
transform 1 0 71400 0 1 13469
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_253
timestamp 1649977179
transform 1 0 74120 0 1 15101
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_254
timestamp 1649977179
transform 1 0 73984 0 1 15101
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_255
timestamp 1649977179
transform 1 0 76568 0 1 15101
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_256
timestamp 1649977179
transform 1 0 76568 0 1 13197
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_257
timestamp 1649977179
transform 1 0 76296 0 1 13061
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_258
timestamp 1649977179
transform 1 0 76296 0 1 12517
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_259
timestamp 1649977179
transform 1 0 71400 0 1 11973
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_260
timestamp 1649977179
transform 1 0 71264 0 1 11021
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_261
timestamp 1649977179
transform 1 0 71264 0 1 11837
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_262
timestamp 1649977179
transform 1 0 68680 0 1 11973
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_263
timestamp 1649977179
transform 1 0 76160 0 1 11701
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_264
timestamp 1649977179
transform 1 0 76024 0 1 14285
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_265
timestamp 1649977179
transform 1 0 76024 0 1 13605
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_266
timestamp 1649977179
transform 1 0 73848 0 1 13605
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_267
timestamp 1649977179
transform 1 0 73848 0 1 14285
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_268
timestamp 1649977179
transform 1 0 73848 0 1 13469
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_269
timestamp 1649977179
transform 1 0 73848 0 1 11973
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_270
timestamp 1649977179
transform 1 0 73712 0 1 11021
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_271
timestamp 1649977179
transform 1 0 73712 0 1 11837
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_272
timestamp 1649977179
transform 1 0 68816 0 1 11021
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_273
timestamp 1649977179
transform 1 0 68816 0 1 11837
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_274
timestamp 1649977179
transform 1 0 76160 0 1 12245
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_275
timestamp 1649977179
transform 1 0 68816 0 1 13605
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_276
timestamp 1649977179
transform 1 0 68816 0 1 14285
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_277
timestamp 1649977179
transform 1 0 68680 0 1 13605
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_278
timestamp 1649977179
transform 1 0 71264 0 1 13605
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_279
timestamp 1649977179
transform 1 0 76296 0 1 13605
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_280
timestamp 1649977179
transform 1 0 76296 0 1 14285
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_281
timestamp 1649977179
transform 1 0 76432 0 1 13469
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_282
timestamp 1649977179
transform 1 0 71400 0 1 17005
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_283
timestamp 1649977179
transform 1 0 69088 0 1 17005
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_284
timestamp 1649977179
transform 1 0 68680 0 1 19181
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_285
timestamp 1649977179
transform 1 0 76432 0 1 17005
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_286
timestamp 1649977179
transform 1 0 74120 0 1 17005
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_287
timestamp 1649977179
transform 1 0 68680 0 1 18773
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_288
timestamp 1649977179
transform 1 0 76160 0 1 19181
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_289
timestamp 1649977179
transform 1 0 76160 0 1 18773
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_290
timestamp 1649977179
transform 1 0 75616 0 1 18773
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_291
timestamp 1649977179
transform 1 0 75616 0 1 19181
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_292
timestamp 1649977179
transform 1 0 74936 0 1 19181
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_293
timestamp 1649977179
transform 1 0 74936 0 1 18773
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_294
timestamp 1649977179
transform 1 0 73168 0 1 18773
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_295
timestamp 1649977179
transform 1 0 73168 0 1 19181
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_296
timestamp 1649977179
transform 1 0 72352 0 1 19181
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_297
timestamp 1649977179
transform 1 0 72352 0 1 18773
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_298
timestamp 1649977179
transform 1 0 71944 0 1 18773
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_299
timestamp 1649977179
transform 1 0 71944 0 1 19181
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_300
timestamp 1649977179
transform 1 0 70992 0 1 18773
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_301
timestamp 1649977179
transform 1 0 70992 0 1 19181
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_302
timestamp 1649977179
transform 1 0 69360 0 1 18773
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_303
timestamp 1649977179
transform 1 0 69360 0 1 19181
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_304
timestamp 1649977179
transform 1 0 78880 0 1 17005
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_305
timestamp 1649977179
transform 1 0 84864 0 1 19181
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_306
timestamp 1649977179
transform 1 0 84864 0 1 18773
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_307
timestamp 1649977179
transform 1 0 84320 0 1 18773
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_308
timestamp 1649977179
transform 1 0 84320 0 1 19181
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_309
timestamp 1649977179
transform 1 0 83912 0 1 17005
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_310
timestamp 1649977179
transform 1 0 83640 0 1 19181
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_311
timestamp 1649977179
transform 1 0 83640 0 1 18773
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_312
timestamp 1649977179
transform 1 0 81872 0 1 18773
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_313
timestamp 1649977179
transform 1 0 81872 0 1 19181
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_314
timestamp 1649977179
transform 1 0 81192 0 1 19181
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_315
timestamp 1649977179
transform 1 0 81192 0 1 18773
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_316
timestamp 1649977179
transform 1 0 80648 0 1 18773
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_317
timestamp 1649977179
transform 1 0 80648 0 1 19181
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_318
timestamp 1649977179
transform 1 0 79696 0 1 18773
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_319
timestamp 1649977179
transform 1 0 79696 0 1 19181
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_320
timestamp 1649977179
transform 1 0 78064 0 1 18773
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_321
timestamp 1649977179
transform 1 0 78064 0 1 19181
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_322
timestamp 1649977179
transform 1 0 77384 0 1 19181
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_323
timestamp 1649977179
transform 1 0 77384 0 1 18773
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_324
timestamp 1649977179
transform 1 0 81600 0 1 17005
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_325
timestamp 1649977179
transform 1 0 96424 0 1 13197
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_326
timestamp 1649977179
transform 1 0 96152 0 1 11837
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_327
timestamp 1649977179
transform 1 0 96424 0 1 13061
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_328
timestamp 1649977179
transform 1 0 96424 0 1 12517
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_329
timestamp 1649977179
transform 1 0 96016 0 1 11701
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_330
timestamp 1649977179
transform 1 0 96016 0 1 12245
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_331
timestamp 1649977179
transform 1 0 96288 0 1 11973
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_332
timestamp 1649977179
transform 1 0 93840 0 1 15101
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_333
timestamp 1649977179
transform 1 0 101320 0 1 13605
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_334
timestamp 1649977179
transform 1 0 101320 0 1 14285
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_335
timestamp 1649977179
transform 1 0 101320 0 1 13469
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_336
timestamp 1649977179
transform 1 0 101320 0 1 11973
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_337
timestamp 1649977179
transform 1 0 101184 0 1 11021
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_338
timestamp 1649977179
transform 1 0 101184 0 1 11837
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_339
timestamp 1649977179
transform 1 0 93976 0 1 15101
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_340
timestamp 1649977179
transform 1 0 93976 0 1 13197
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_341
timestamp 1649977179
transform 1 0 96288 0 1 13605
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_342
timestamp 1649977179
transform 1 0 93976 0 1 13061
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_343
timestamp 1649977179
transform 1 0 98872 0 1 13605
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_344
timestamp 1649977179
transform 1 0 98872 0 1 14285
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_345
timestamp 1649977179
transform 1 0 98872 0 1 13469
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_346
timestamp 1649977179
transform 1 0 98872 0 1 11973
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_347
timestamp 1649977179
transform 1 0 98736 0 1 11021
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_348
timestamp 1649977179
transform 1 0 98736 0 1 11837
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_349
timestamp 1649977179
transform 1 0 93976 0 1 12517
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_350
timestamp 1649977179
transform 1 0 96152 0 1 11021
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_351
timestamp 1649977179
transform 1 0 93840 0 1 13469
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_352
timestamp 1649977179
transform 1 0 96288 0 1 14285
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_353
timestamp 1649977179
transform 1 0 93840 0 1 11973
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_354
timestamp 1649977179
transform 1 0 101592 0 1 15101
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_355
timestamp 1649977179
transform 1 0 101456 0 1 15101
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_356
timestamp 1649977179
transform 1 0 101456 0 1 13197
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_357
timestamp 1649977179
transform 1 0 101456 0 1 13061
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_358
timestamp 1649977179
transform 1 0 101456 0 1 12517
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_359
timestamp 1649977179
transform 1 0 101456 0 1 11701
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_360
timestamp 1649977179
transform 1 0 101456 0 1 12245
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_361
timestamp 1649977179
transform 1 0 93840 0 1 13605
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_362
timestamp 1649977179
transform 1 0 98872 0 1 15101
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_363
timestamp 1649977179
transform 1 0 99008 0 1 15101
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_364
timestamp 1649977179
transform 1 0 99008 0 1 13197
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_365
timestamp 1649977179
transform 1 0 99008 0 1 13061
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_366
timestamp 1649977179
transform 1 0 99008 0 1 12517
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_367
timestamp 1649977179
transform 1 0 100912 0 1 13061
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_368
timestamp 1649977179
transform 1 0 98464 0 1 13061
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_369
timestamp 1649977179
transform 1 0 95880 0 1 13061
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_370
timestamp 1649977179
transform 1 0 99008 0 1 11701
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_371
timestamp 1649977179
transform 1 0 99008 0 1 12245
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_372
timestamp 1649977179
transform 1 0 96288 0 1 13469
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_373
timestamp 1649977179
transform 1 0 93840 0 1 14285
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_374
timestamp 1649977179
transform 1 0 96560 0 1 15101
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_375
timestamp 1649977179
transform 1 0 96424 0 1 15101
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_376
timestamp 1649977179
transform 1 0 88944 0 1 15101
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_377
timestamp 1649977179
transform 1 0 88944 0 1 13197
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_378
timestamp 1649977179
transform 1 0 88944 0 1 13061
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_379
timestamp 1649977179
transform 1 0 88944 0 1 12517
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_380
timestamp 1649977179
transform 1 0 88944 0 1 11701
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_381
timestamp 1649977179
transform 1 0 88944 0 1 12245
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_382
timestamp 1649977179
transform 1 0 91256 0 1 13605
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_383
timestamp 1649977179
transform 1 0 91256 0 1 14285
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_384
timestamp 1649977179
transform 1 0 91392 0 1 13469
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_385
timestamp 1649977179
transform 1 0 91392 0 1 11973
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_386
timestamp 1649977179
transform 1 0 91120 0 1 11021
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_387
timestamp 1649977179
transform 1 0 91120 0 1 11837
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_388
timestamp 1649977179
transform 1 0 86496 0 1 12245
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_389
timestamp 1649977179
transform 1 0 93568 0 1 11021
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_390
timestamp 1649977179
transform 1 0 86360 0 1 15101
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_391
timestamp 1649977179
transform 1 0 93568 0 1 11837
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_392
timestamp 1649977179
transform 1 0 86496 0 1 15101
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_393
timestamp 1649977179
transform 1 0 86496 0 1 13197
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_394
timestamp 1649977179
transform 1 0 88672 0 1 13605
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_395
timestamp 1649977179
transform 1 0 88672 0 1 14285
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_396
timestamp 1649977179
transform 1 0 88808 0 1 13469
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_397
timestamp 1649977179
transform 1 0 88808 0 1 11973
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_398
timestamp 1649977179
transform 1 0 88808 0 1 11021
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_399
timestamp 1649977179
transform 1 0 88808 0 1 11837
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_400
timestamp 1649977179
transform 1 0 86496 0 1 13061
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_401
timestamp 1649977179
transform 1 0 93704 0 1 12245
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_402
timestamp 1649977179
transform 1 0 93704 0 1 11429
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_403
timestamp 1649977179
transform 1 0 86496 0 1 12517
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_404
timestamp 1649977179
transform 1 0 91392 0 1 15101
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_405
timestamp 1649977179
transform 1 0 91528 0 1 15101
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_406
timestamp 1649977179
transform 1 0 91528 0 1 13197
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_407
timestamp 1649977179
transform 1 0 91256 0 1 13061
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_408
timestamp 1649977179
transform 1 0 86224 0 1 13605
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_409
timestamp 1649977179
transform 1 0 86224 0 1 14285
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_410
timestamp 1649977179
transform 1 0 86360 0 1 13469
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_411
timestamp 1649977179
transform 1 0 86360 0 1 11973
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_412
timestamp 1649977179
transform 1 0 86224 0 1 11021
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_413
timestamp 1649977179
transform 1 0 86224 0 1 11837
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_414
timestamp 1649977179
transform 1 0 91256 0 1 12517
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_415
timestamp 1649977179
transform 1 0 91256 0 1 11701
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_416
timestamp 1649977179
transform 1 0 86088 0 1 14285
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_417
timestamp 1649977179
transform 1 0 86088 0 1 13605
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_418
timestamp 1649977179
transform 1 0 93432 0 1 13061
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_419
timestamp 1649977179
transform 1 0 90984 0 1 13061
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_420
timestamp 1649977179
transform 1 0 88536 0 1 13061
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_421
timestamp 1649977179
transform 1 0 85952 0 1 13061
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_422
timestamp 1649977179
transform 1 0 91256 0 1 12245
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_423
timestamp 1649977179
transform 1 0 86496 0 1 11701
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_424
timestamp 1649977179
transform 1 0 89080 0 1 15101
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_425
timestamp 1649977179
transform 1 0 93432 0 1 18773
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_426
timestamp 1649977179
transform 1 0 93432 0 1 19181
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_427
timestamp 1649977179
transform 1 0 92344 0 1 19181
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_428
timestamp 1649977179
transform 1 0 92344 0 1 18773
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_429
timestamp 1649977179
transform 1 0 91800 0 1 18773
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_430
timestamp 1649977179
transform 1 0 91800 0 1 19181
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_431
timestamp 1649977179
transform 1 0 90712 0 1 18773
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_432
timestamp 1649977179
transform 1 0 90712 0 1 19181
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_433
timestamp 1649977179
transform 1 0 89896 0 1 19181
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_434
timestamp 1649977179
transform 1 0 89896 0 1 18773
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_435
timestamp 1649977179
transform 1 0 89352 0 1 18773
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_436
timestamp 1649977179
transform 1 0 89352 0 1 19181
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_437
timestamp 1649977179
transform 1 0 88264 0 1 19181
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_438
timestamp 1649977179
transform 1 0 88264 0 1 18773
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_439
timestamp 1649977179
transform 1 0 88128 0 1 18773
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_440
timestamp 1649977179
transform 1 0 88128 0 1 19181
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_441
timestamp 1649977179
transform 1 0 87312 0 1 19181
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_442
timestamp 1649977179
transform 1 0 87312 0 1 18773
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_443
timestamp 1649977179
transform 1 0 86904 0 1 18773
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_444
timestamp 1649977179
transform 1 0 86904 0 1 19181
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_445
timestamp 1649977179
transform 1 0 86088 0 1 19181
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_446
timestamp 1649977179
transform 1 0 86088 0 1 18773
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_447
timestamp 1649977179
transform 1 0 86360 0 1 17005
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_448
timestamp 1649977179
transform 1 0 91392 0 1 17005
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_449
timestamp 1649977179
transform 1 0 89080 0 1 17005
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_450
timestamp 1649977179
transform 1 0 101864 0 1 18773
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_451
timestamp 1649977179
transform 1 0 101864 0 1 19181
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_452
timestamp 1649977179
transform 1 0 101184 0 1 19181
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_453
timestamp 1649977179
transform 1 0 101184 0 1 18773
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_454
timestamp 1649977179
transform 1 0 99824 0 1 19181
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_455
timestamp 1649977179
transform 1 0 99824 0 1 18773
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_456
timestamp 1649977179
transform 1 0 98600 0 1 19181
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_457
timestamp 1649977179
transform 1 0 98600 0 1 18773
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_458
timestamp 1649977179
transform 1 0 98192 0 1 18773
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_459
timestamp 1649977179
transform 1 0 98192 0 1 19181
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_460
timestamp 1649977179
transform 1 0 101592 0 1 17005
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_461
timestamp 1649977179
transform 1 0 98872 0 1 17005
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_462
timestamp 1649977179
transform 1 0 96832 0 1 18773
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_463
timestamp 1649977179
transform 1 0 96560 0 1 17005
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_464
timestamp 1649977179
transform 1 0 96832 0 1 19181
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_465
timestamp 1649977179
transform 1 0 93976 0 1 17005
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_466
timestamp 1649977179
transform 1 0 96152 0 1 19181
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_467
timestamp 1649977179
transform 1 0 96152 0 1 18773
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_468
timestamp 1649977179
transform 1 0 95608 0 1 18773
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_469
timestamp 1649977179
transform 1 0 95608 0 1 19181
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_470
timestamp 1649977179
transform 1 0 94520 0 1 19317
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_471
timestamp 1649977179
transform 1 0 94520 0 1 18773
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_472
timestamp 1649977179
transform 1 0 135320 0 1 25437
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_473
timestamp 1649977179
transform 1 0 135320 0 1 23805
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_474
timestamp 1649977179
transform 1 0 135320 0 1 22173
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_475
timestamp 1649977179
transform 1 0 119408 0 1 25029
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_476
timestamp 1649977179
transform 1 0 119408 0 1 25709
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_477
timestamp 1649977179
transform 1 0 120768 0 1 25029
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_478
timestamp 1649977179
transform 1 0 120768 0 1 25709
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_479
timestamp 1649977179
transform 1 0 135320 0 1 27205
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_480
timestamp 1649977179
transform 1 0 135320 0 1 28973
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_481
timestamp 1649977179
transform 1 0 135320 0 1 30469
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_482
timestamp 1649977179
transform 1 0 117640 0 1 22717
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_483
timestamp 1649977179
transform 1 0 117640 0 1 23397
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_484
timestamp 1649977179
transform 1 0 115600 0 1 21765
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_485
timestamp 1649977179
transform 1 0 115600 0 1 21085
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_486
timestamp 1649977179
transform 1 0 118048 0 1 21085
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_487
timestamp 1649977179
transform 1 0 118048 0 1 21357
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_488
timestamp 1649977179
transform 1 0 115872 0 1 21901
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_489
timestamp 1649977179
transform 1 0 115872 0 1 22173
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_490
timestamp 1649977179
transform 1 0 115872 0 1 22581
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_491
timestamp 1649977179
transform 1 0 115872 0 1 22309
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_492
timestamp 1649977179
transform 1 0 116008 0 1 21493
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_493
timestamp 1649977179
transform 1 0 116008 0 1 21765
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_494
timestamp 1649977179
transform 1 0 119000 0 1 22717
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_495
timestamp 1649977179
transform 1 0 119000 0 1 23261
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_496
timestamp 1649977179
transform 1 0 115600 0 1 21357
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_497
timestamp 1649977179
transform 1 0 115600 0 1 21493
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_498
timestamp 1649977179
transform 1 0 116008 0 1 22989
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_499
timestamp 1649977179
transform 1 0 118864 0 1 22445
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_500
timestamp 1649977179
transform 1 0 118864 0 1 22173
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_501
timestamp 1649977179
transform 1 0 118320 0 1 22173
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_502
timestamp 1649977179
transform 1 0 118320 0 1 21085
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_503
timestamp 1649977179
transform 1 0 118184 0 1 23397
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_504
timestamp 1649977179
transform 1 0 116008 0 1 22717
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_505
timestamp 1649977179
transform 1 0 117640 0 1 23261
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_506
timestamp 1649977179
transform 1 0 118456 0 1 22445
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_507
timestamp 1649977179
transform 1 0 118864 0 1 22717
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_508
timestamp 1649977179
transform 1 0 118864 0 1 22989
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_509
timestamp 1649977179
transform 1 0 118320 0 1 22989
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_510
timestamp 1649977179
transform 1 0 118320 0 1 22717
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_511
timestamp 1649977179
transform 1 0 118048 0 1 23261
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_512
timestamp 1649977179
transform 1 0 118048 0 1 22717
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_513
timestamp 1649977179
transform 1 0 115872 0 1 21357
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_514
timestamp 1649977179
transform 1 0 118592 0 1 22717
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_515
timestamp 1649977179
transform 1 0 115872 0 1 21085
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_516
timestamp 1649977179
transform 1 0 118456 0 1 21221
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_517
timestamp 1649977179
transform 1 0 118592 0 1 23261
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_518
timestamp 1649977179
transform 1 0 114240 0 1 21085
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_519
timestamp 1649977179
transform 1 0 114648 0 1 21765
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_520
timestamp 1649977179
transform 1 0 114784 0 1 22989
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_521
timestamp 1649977179
transform 1 0 114784 0 1 23261
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_522
timestamp 1649977179
transform 1 0 114240 0 1 21357
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_523
timestamp 1649977179
transform 1 0 114376 0 1 23261
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_524
timestamp 1649977179
transform 1 0 114376 0 1 22989
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_525
timestamp 1649977179
transform 1 0 114240 0 1 23397
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_526
timestamp 1649977179
transform 1 0 114240 0 1 21493
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_527
timestamp 1649977179
transform 1 0 114240 0 1 21765
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_528
timestamp 1649977179
transform 1 0 114784 0 1 23397
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_529
timestamp 1649977179
transform 1 0 114648 0 1 21493
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_530
timestamp 1649977179
transform 1 0 114648 0 1 21085
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_531
timestamp 1649977179
transform 1 0 114648 0 1 21357
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_532
timestamp 1649977179
transform 1 0 114240 0 1 24893
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_533
timestamp 1649977179
transform 1 0 114240 0 1 25301
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_534
timestamp 1649977179
transform 1 0 114376 0 1 24213
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_535
timestamp 1649977179
transform 1 0 114376 0 1 24485
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_536
timestamp 1649977179
transform 1 0 114240 0 1 25437
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_537
timestamp 1649977179
transform 1 0 114240 0 1 25709
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_538
timestamp 1649977179
transform 1 0 114240 0 1 25029
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_539
timestamp 1649977179
transform 1 0 114784 0 1 24077
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_540
timestamp 1649977179
transform 1 0 114240 0 1 25845
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_541
timestamp 1649977179
transform 1 0 114648 0 1 25845
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_542
timestamp 1649977179
transform 1 0 114784 0 1 24485
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_543
timestamp 1649977179
transform 1 0 114784 0 1 23805
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_544
timestamp 1649977179
transform 1 0 114784 0 1 23669
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_545
timestamp 1649977179
transform 1 0 114784 0 1 24213
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_546
timestamp 1649977179
transform 1 0 114240 0 1 24621
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_547
timestamp 1649977179
transform 1 0 114648 0 1 24621
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_548
timestamp 1649977179
transform 1 0 114784 0 1 25709
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_549
timestamp 1649977179
transform 1 0 114648 0 1 24893
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_550
timestamp 1649977179
transform 1 0 114648 0 1 25301
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_551
timestamp 1649977179
transform 1 0 114784 0 1 25437
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_552
timestamp 1649977179
transform 1 0 114240 0 1 24077
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_553
timestamp 1649977179
transform 1 0 114240 0 1 23805
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_554
timestamp 1649977179
transform 1 0 114648 0 1 25029
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_555
timestamp 1649977179
transform 1 0 114240 0 1 23669
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_556
timestamp 1649977179
transform 1 0 119000 0 1 25709
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_557
timestamp 1649977179
transform 1 0 119000 0 1 25029
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_558
timestamp 1649977179
transform 1 0 115192 0 1 23805
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_559
timestamp 1649977179
transform 1 0 115192 0 1 24077
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_560
timestamp 1649977179
transform 1 0 116008 0 1 25845
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_561
timestamp 1649977179
transform 1 0 118184 0 1 24893
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_562
timestamp 1649977179
transform 1 0 118184 0 1 25709
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_563
timestamp 1649977179
transform 1 0 118184 0 1 25029
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_564
timestamp 1649977179
transform 1 0 115464 0 1 24621
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_565
timestamp 1649977179
transform 1 0 115872 0 1 24213
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_566
timestamp 1649977179
transform 1 0 115872 0 1 24485
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_567
timestamp 1649977179
transform 1 0 118184 0 1 25845
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_568
timestamp 1649977179
transform 1 0 115464 0 1 24893
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_569
timestamp 1649977179
transform 1 0 115464 0 1 25301
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_570
timestamp 1649977179
transform 1 0 115464 0 1 25029
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_571
timestamp 1649977179
transform 1 0 116008 0 1 25437
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_572
timestamp 1649977179
transform 1 0 115192 0 1 25029
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_573
timestamp 1649977179
transform 1 0 115192 0 1 25301
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_574
timestamp 1649977179
transform 1 0 117640 0 1 25845
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_575
timestamp 1649977179
transform 1 0 115872 0 1 25029
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_576
timestamp 1649977179
transform 1 0 115872 0 1 25301
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_577
timestamp 1649977179
transform 1 0 115600 0 1 23805
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_578
timestamp 1649977179
transform 1 0 116008 0 1 25709
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_579
timestamp 1649977179
transform 1 0 115600 0 1 25437
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_580
timestamp 1649977179
transform 1 0 115600 0 1 25709
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_581
timestamp 1649977179
transform 1 0 117640 0 1 25709
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_582
timestamp 1649977179
transform 1 0 117640 0 1 25029
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_583
timestamp 1649977179
transform 1 0 117640 0 1 24893
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_584
timestamp 1649977179
transform 1 0 116008 0 1 24893
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_585
timestamp 1649977179
transform 1 0 116008 0 1 24621
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_586
timestamp 1649977179
transform 1 0 119000 0 1 25845
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_587
timestamp 1649977179
transform 1 0 115600 0 1 24077
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_588
timestamp 1649977179
transform 1 0 115056 0 1 24621
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_589
timestamp 1649977179
transform 1 0 115056 0 1 21493
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_590
timestamp 1649977179
transform 1 0 115056 0 1 21765
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_591
timestamp 1649977179
transform 1 0 115056 0 1 22309
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_592
timestamp 1649977179
transform 1 0 115056 0 1 22581
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_593
timestamp 1649977179
transform 1 0 115056 0 1 24893
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_594
timestamp 1649977179
transform 1 0 115056 0 1 25437
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_595
timestamp 1649977179
transform 1 0 115056 0 1 25709
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_596
timestamp 1649977179
transform 1 0 109344 0 1 22853
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_597
timestamp 1649977179
transform 1 0 109344 0 1 22309
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_598
timestamp 1649977179
transform 1 0 109480 0 1 22717
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_599
timestamp 1649977179
transform 1 0 109344 0 1 23125
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_600
timestamp 1649977179
transform 1 0 109344 0 1 22037
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_601
timestamp 1649977179
transform 1 0 109344 0 1 21493
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_602
timestamp 1649977179
transform 1 0 109344 0 1 21221
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_603
timestamp 1649977179
transform 1 0 109480 0 1 22445
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_604
timestamp 1649977179
transform 1 0 109344 0 1 25981
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_605
timestamp 1649977179
transform 1 0 109344 0 1 26661
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_606
timestamp 1649977179
transform 1 0 109344 0 1 30333
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_607
timestamp 1649977179
transform 1 0 109344 0 1 30605
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_608
timestamp 1649977179
transform 1 0 109344 0 1 26389
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_609
timestamp 1649977179
transform 1 0 109344 0 1 26253
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_610
timestamp 1649977179
transform 1 0 109344 0 1 30197
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_611
timestamp 1649977179
transform 1 0 109344 0 1 29925
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_612
timestamp 1649977179
transform 1 0 109344 0 1 31149
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_613
timestamp 1649977179
transform 1 0 114240 0 1 29789
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_614
timestamp 1649977179
transform 1 0 114240 0 1 30061
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_615
timestamp 1649977179
transform 1 0 118184 0 1 27205
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_616
timestamp 1649977179
transform 1 0 118184 0 1 26661
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_617
timestamp 1649977179
transform 1 0 118184 0 1 26389
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_618
timestamp 1649977179
transform 1 0 114240 0 1 28973
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_619
timestamp 1649977179
transform 1 0 115600 0 1 28157
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_620
timestamp 1649977179
transform 1 0 114240 0 1 29245
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_621
timestamp 1649977179
transform 1 0 114240 0 1 29653
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_622
timestamp 1649977179
transform 1 0 114240 0 1 29381
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_623
timestamp 1649977179
transform 1 0 114784 0 1 28565
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_624
timestamp 1649977179
transform 1 0 115872 0 1 30877
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_625
timestamp 1649977179
transform 1 0 115872 0 1 30605
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_626
timestamp 1649977179
transform 1 0 114376 0 1 28021
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_627
timestamp 1649977179
transform 1 0 115600 0 1 28429
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_628
timestamp 1649977179
transform 1 0 115192 0 1 28021
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_629
timestamp 1649977179
transform 1 0 115192 0 1 27749
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_630
timestamp 1649977179
transform 1 0 114376 0 1 27749
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_631
timestamp 1649977179
transform 1 0 115056 0 1 28973
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_632
timestamp 1649977179
transform 1 0 115056 0 1 29245
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_633
timestamp 1649977179
transform 1 0 115464 0 1 29653
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_634
timestamp 1649977179
transform 1 0 115464 0 1 29381
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_635
timestamp 1649977179
transform 1 0 115192 0 1 28837
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_636
timestamp 1649977179
transform 1 0 115192 0 1 28565
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_637
timestamp 1649977179
transform 1 0 117640 0 1 27205
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_638
timestamp 1649977179
transform 1 0 117640 0 1 26797
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_639
timestamp 1649977179
transform 1 0 115736 0 1 26797
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_640
timestamp 1649977179
transform 1 0 114784 0 1 28021
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_641
timestamp 1649977179
transform 1 0 114784 0 1 27749
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_642
timestamp 1649977179
transform 1 0 115736 0 1 27205
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_643
timestamp 1649977179
transform 1 0 114784 0 1 28157
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_644
timestamp 1649977179
transform 1 0 115872 0 1 28157
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_645
timestamp 1649977179
transform 1 0 115872 0 1 28429
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_646
timestamp 1649977179
transform 1 0 114648 0 1 28973
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_647
timestamp 1649977179
transform 1 0 114648 0 1 29245
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_648
timestamp 1649977179
transform 1 0 114648 0 1 29653
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_649
timestamp 1649977179
transform 1 0 114648 0 1 29381
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_650
timestamp 1649977179
transform 1 0 119000 0 1 26525
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_651
timestamp 1649977179
transform 1 0 118864 0 1 27205
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_652
timestamp 1649977179
transform 1 0 118728 0 1 26661
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_653
timestamp 1649977179
transform 1 0 114376 0 1 28837
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_654
timestamp 1649977179
transform 1 0 114376 0 1 28565
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_655
timestamp 1649977179
transform 1 0 114376 0 1 28157
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_656
timestamp 1649977179
transform 1 0 114376 0 1 28429
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_657
timestamp 1649977179
transform 1 0 114648 0 1 29789
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_658
timestamp 1649977179
transform 1 0 114648 0 1 30061
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_659
timestamp 1649977179
transform 1 0 114784 0 1 28429
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_660
timestamp 1649977179
transform 1 0 115600 0 1 26933
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_661
timestamp 1649977179
transform 1 0 116008 0 1 30469
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_662
timestamp 1649977179
transform 1 0 116008 0 1 30197
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_663
timestamp 1649977179
transform 1 0 117640 0 1 26389
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_664
timestamp 1649977179
transform 1 0 115600 0 1 27205
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_665
timestamp 1649977179
transform 1 0 117776 0 1 26661
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_666
timestamp 1649977179
transform 1 0 117776 0 1 27205
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_667
timestamp 1649977179
transform 1 0 116008 0 1 29245
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_668
timestamp 1649977179
transform 1 0 116008 0 1 28973
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_669
timestamp 1649977179
transform 1 0 115872 0 1 28565
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_670
timestamp 1649977179
transform 1 0 115872 0 1 28837
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_671
timestamp 1649977179
transform 1 0 115328 0 1 29245
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_672
timestamp 1649977179
transform 1 0 115328 0 1 28973
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_673
timestamp 1649977179
transform 1 0 115464 0 1 31149
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_674
timestamp 1649977179
transform 1 0 115464 0 1 30877
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_675
timestamp 1649977179
transform 1 0 115464 0 1 26253
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_676
timestamp 1649977179
transform 1 0 115464 0 1 26525
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_677
timestamp 1649977179
transform 1 0 115872 0 1 26253
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_678
timestamp 1649977179
transform 1 0 115872 0 1 26525
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_679
timestamp 1649977179
transform 1 0 115872 0 1 26933
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_680
timestamp 1649977179
transform 1 0 115872 0 1 26661
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_681
timestamp 1649977179
transform 1 0 115464 0 1 30197
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_682
timestamp 1649977179
transform 1 0 115464 0 1 30469
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_683
timestamp 1649977179
transform 1 0 114784 0 1 27613
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_684
timestamp 1649977179
transform 1 0 114784 0 1 27341
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_685
timestamp 1649977179
transform 1 0 114376 0 1 27613
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_686
timestamp 1649977179
transform 1 0 114376 0 1 27341
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_687
timestamp 1649977179
transform 1 0 115872 0 1 29381
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_688
timestamp 1649977179
transform 1 0 115872 0 1 29653
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_689
timestamp 1649977179
transform 1 0 115872 0 1 30061
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_690
timestamp 1649977179
transform 1 0 115872 0 1 29789
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_691
timestamp 1649977179
transform 1 0 115328 0 1 29381
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_692
timestamp 1649977179
transform 1 0 115328 0 1 29653
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_693
timestamp 1649977179
transform 1 0 114784 0 1 28837
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_694
timestamp 1649977179
transform 1 0 114648 0 1 26117
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_695
timestamp 1649977179
transform 1 0 116008 0 1 26117
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_696
timestamp 1649977179
transform 1 0 114240 0 1 26117
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_697
timestamp 1649977179
transform 1 0 115328 0 1 34005
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_698
timestamp 1649977179
transform 1 0 114648 0 1 33597
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_699
timestamp 1649977179
transform 1 0 115328 0 1 36317
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_700
timestamp 1649977179
transform 1 0 114648 0 1 34141
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_701
timestamp 1649977179
transform 1 0 114648 0 1 34413
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_702
timestamp 1649977179
transform 1 0 114648 0 1 33325
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_703
timestamp 1649977179
transform 1 0 114376 0 1 31965
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_704
timestamp 1649977179
transform 1 0 114376 0 1 31693
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_705
timestamp 1649977179
transform 1 0 115192 0 1 32373
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_706
timestamp 1649977179
transform 1 0 114784 0 1 31965
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_707
timestamp 1649977179
transform 1 0 114240 0 1 31557
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_708
timestamp 1649977179
transform 1 0 115192 0 1 32101
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_709
timestamp 1649977179
transform 1 0 114240 0 1 35637
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_710
timestamp 1649977179
transform 1 0 114376 0 1 33189
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_711
timestamp 1649977179
transform 1 0 114376 0 1 32917
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_712
timestamp 1649977179
transform 1 0 114376 0 1 32509
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_713
timestamp 1649977179
transform 1 0 114376 0 1 32781
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_714
timestamp 1649977179
transform 1 0 115872 0 1 33189
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_715
timestamp 1649977179
transform 1 0 115872 0 1 32917
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_716
timestamp 1649977179
transform 1 0 115872 0 1 32509
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_717
timestamp 1649977179
transform 1 0 115872 0 1 32781
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_718
timestamp 1649977179
transform 1 0 115328 0 1 36045
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_719
timestamp 1649977179
transform 1 0 115192 0 1 36317
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_720
timestamp 1649977179
transform 1 0 115192 0 1 36045
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_721
timestamp 1649977179
transform 1 0 114240 0 1 35909
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_722
timestamp 1649977179
transform 1 0 116008 0 1 36045
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_723
timestamp 1649977179
transform 1 0 116008 0 1 36317
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_724
timestamp 1649977179
transform 1 0 115872 0 1 32373
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_725
timestamp 1649977179
transform 1 0 115872 0 1 32101
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_726
timestamp 1649977179
transform 1 0 114376 0 1 36317
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_727
timestamp 1649977179
transform 1 0 114376 0 1 36045
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_728
timestamp 1649977179
transform 1 0 114784 0 1 33733
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_729
timestamp 1649977179
transform 1 0 114784 0 1 33189
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_730
timestamp 1649977179
transform 1 0 114784 0 1 32917
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_731
timestamp 1649977179
transform 1 0 114784 0 1 32509
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_732
timestamp 1649977179
transform 1 0 114784 0 1 32781
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_733
timestamp 1649977179
transform 1 0 114648 0 1 35909
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_734
timestamp 1649977179
transform 1 0 114648 0 1 35637
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_735
timestamp 1649977179
transform 1 0 115056 0 1 33325
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_736
timestamp 1649977179
transform 1 0 115056 0 1 33597
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_737
timestamp 1649977179
transform 1 0 114784 0 1 34005
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_738
timestamp 1649977179
transform 1 0 114240 0 1 34141
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_739
timestamp 1649977179
transform 1 0 114784 0 1 31693
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_740
timestamp 1649977179
transform 1 0 115192 0 1 32917
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_741
timestamp 1649977179
transform 1 0 115872 0 1 31693
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_742
timestamp 1649977179
transform 1 0 115872 0 1 31421
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_743
timestamp 1649977179
transform 1 0 115600 0 1 34141
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_744
timestamp 1649977179
transform 1 0 115600 0 1 34413
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_745
timestamp 1649977179
transform 1 0 114240 0 1 34413
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_746
timestamp 1649977179
transform 1 0 114648 0 1 31557
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_747
timestamp 1649977179
transform 1 0 115328 0 1 32373
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_748
timestamp 1649977179
transform 1 0 115328 0 1 32101
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_749
timestamp 1649977179
transform 1 0 114240 0 1 32101
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_750
timestamp 1649977179
transform 1 0 115872 0 1 35229
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_751
timestamp 1649977179
transform 1 0 115872 0 1 34957
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_752
timestamp 1649977179
transform 1 0 116008 0 1 34549
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_753
timestamp 1649977179
transform 1 0 116008 0 1 34821
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_754
timestamp 1649977179
transform 1 0 114240 0 1 32373
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_755
timestamp 1649977179
transform 1 0 114648 0 1 32101
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_756
timestamp 1649977179
transform 1 0 115600 0 1 33597
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_757
timestamp 1649977179
transform 1 0 115600 0 1 33733
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_758
timestamp 1649977179
transform 1 0 115600 0 1 34005
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_759
timestamp 1649977179
transform 1 0 115600 0 1 33325
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_760
timestamp 1649977179
transform 1 0 115600 0 1 32509
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_761
timestamp 1649977179
transform 1 0 115600 0 1 32781
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_762
timestamp 1649977179
transform 1 0 114648 0 1 32373
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_763
timestamp 1649977179
transform 1 0 115872 0 1 35637
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_764
timestamp 1649977179
transform 1 0 115872 0 1 35365
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_765
timestamp 1649977179
transform 1 0 115464 0 1 35229
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_766
timestamp 1649977179
transform 1 0 115464 0 1 34821
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_767
timestamp 1649977179
transform 1 0 115464 0 1 35637
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_768
timestamp 1649977179
transform 1 0 115464 0 1 35909
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_769
timestamp 1649977179
transform 1 0 116008 0 1 33325
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_770
timestamp 1649977179
transform 1 0 116008 0 1 33597
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_771
timestamp 1649977179
transform 1 0 116008 0 1 34005
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_772
timestamp 1649977179
transform 1 0 116008 0 1 33733
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_773
timestamp 1649977179
transform 1 0 115192 0 1 34141
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_774
timestamp 1649977179
transform 1 0 115192 0 1 34413
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_775
timestamp 1649977179
transform 1 0 115192 0 1 33189
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_776
timestamp 1649977179
transform 1 0 115328 0 1 33733
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_777
timestamp 1649977179
transform 1 0 116008 0 1 34141
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_778
timestamp 1649977179
transform 1 0 116008 0 1 34413
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_779
timestamp 1649977179
transform 1 0 114784 0 1 36317
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_780
timestamp 1649977179
transform 1 0 114240 0 1 34005
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_781
timestamp 1649977179
transform 1 0 114240 0 1 33733
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_782
timestamp 1649977179
transform 1 0 114240 0 1 33325
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_783
timestamp 1649977179
transform 1 0 114240 0 1 33597
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_784
timestamp 1649977179
transform 1 0 114784 0 1 36045
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_785
timestamp 1649977179
transform 1 0 109480 0 1 33869
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_786
timestamp 1649977179
transform 1 0 109480 0 1 34141
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_787
timestamp 1649977179
transform 1 0 109344 0 1 34957
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_788
timestamp 1649977179
transform 1 0 109344 0 1 34685
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_789
timestamp 1649977179
transform 1 0 109480 0 1 31829
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_790
timestamp 1649977179
transform 1 0 109480 0 1 31557
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_791
timestamp 1649977179
transform 1 0 109344 0 1 31557
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_792
timestamp 1649977179
transform 1 0 109480 0 1 34413
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_793
timestamp 1649977179
transform 1 0 109480 0 1 34685
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_794
timestamp 1649977179
transform 1 0 109480 0 1 39309
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_795
timestamp 1649977179
transform 1 0 109480 0 1 39037
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_796
timestamp 1649977179
transform 1 0 109480 0 1 40533
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_797
timestamp 1649977179
transform 1 0 109480 0 1 40261
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_798
timestamp 1649977179
transform 1 0 109480 0 1 37813
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_799
timestamp 1649977179
transform 1 0 109480 0 1 38085
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_800
timestamp 1649977179
transform 1 0 109344 0 1 39853
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_801
timestamp 1649977179
transform 1 0 109344 0 1 40261
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_802
timestamp 1649977179
transform 1 0 114240 0 1 37949
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_803
timestamp 1649977179
transform 1 0 114240 0 1 37677
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_804
timestamp 1649977179
transform 1 0 114784 0 1 37541
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_805
timestamp 1649977179
transform 1 0 114784 0 1 37269
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_806
timestamp 1649977179
transform 1 0 114376 0 1 41213
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_807
timestamp 1649977179
transform 1 0 114376 0 1 41485
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_808
timestamp 1649977179
transform 1 0 114784 0 1 36861
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_809
timestamp 1649977179
transform 1 0 114784 0 1 37133
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_810
timestamp 1649977179
transform 1 0 115328 0 1 38085
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_811
timestamp 1649977179
transform 1 0 116008 0 1 37677
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_812
timestamp 1649977179
transform 1 0 116008 0 1 37949
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_813
timestamp 1649977179
transform 1 0 115328 0 1 38357
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_814
timestamp 1649977179
transform 1 0 115872 0 1 37541
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_815
timestamp 1649977179
transform 1 0 115872 0 1 37269
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_816
timestamp 1649977179
transform 1 0 115872 0 1 36861
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_817
timestamp 1649977179
transform 1 0 115872 0 1 37133
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_818
timestamp 1649977179
transform 1 0 115192 0 1 38085
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_819
timestamp 1649977179
transform 1 0 115192 0 1 38357
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_820
timestamp 1649977179
transform 1 0 115192 0 1 39853
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_821
timestamp 1649977179
transform 1 0 115192 0 1 39581
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_822
timestamp 1649977179
transform 1 0 114784 0 1 41213
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_823
timestamp 1649977179
transform 1 0 114376 0 1 40397
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_824
timestamp 1649977179
transform 1 0 115872 0 1 39581
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_825
timestamp 1649977179
transform 1 0 115872 0 1 39309
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_826
timestamp 1649977179
transform 1 0 114376 0 1 40669
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_827
timestamp 1649977179
transform 1 0 114376 0 1 41077
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_828
timestamp 1649977179
transform 1 0 114376 0 1 40805
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_829
timestamp 1649977179
transform 1 0 114376 0 1 37541
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_830
timestamp 1649977179
transform 1 0 114376 0 1 37269
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_831
timestamp 1649977179
transform 1 0 114784 0 1 41485
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_832
timestamp 1649977179
transform 1 0 114648 0 1 37677
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_833
timestamp 1649977179
transform 1 0 114648 0 1 37949
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_834
timestamp 1649977179
transform 1 0 114648 0 1 38357
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_835
timestamp 1649977179
transform 1 0 114648 0 1 38085
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_836
timestamp 1649977179
transform 1 0 115872 0 1 38085
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_837
timestamp 1649977179
transform 1 0 115872 0 1 38357
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_838
timestamp 1649977179
transform 1 0 114376 0 1 38085
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_839
timestamp 1649977179
transform 1 0 116008 0 1 39173
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_840
timestamp 1649977179
transform 1 0 116008 0 1 38901
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_841
timestamp 1649977179
transform 1 0 116008 0 1 38493
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_842
timestamp 1649977179
transform 1 0 116008 0 1 38765
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_843
timestamp 1649977179
transform 1 0 114376 0 1 38357
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_844
timestamp 1649977179
transform 1 0 115600 0 1 36861
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_845
timestamp 1649977179
transform 1 0 115600 0 1 37133
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_846
timestamp 1649977179
transform 1 0 116008 0 1 41485
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_847
timestamp 1649977179
transform 1 0 116008 0 1 41213
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_848
timestamp 1649977179
transform 1 0 116008 0 1 40805
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_849
timestamp 1649977179
transform 1 0 116008 0 1 41077
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_850
timestamp 1649977179
transform 1 0 115464 0 1 36725
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_851
timestamp 1649977179
transform 1 0 114648 0 1 39853
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_852
timestamp 1649977179
transform 1 0 115464 0 1 41077
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_853
timestamp 1649977179
transform 1 0 115464 0 1 40805
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_854
timestamp 1649977179
transform 1 0 115600 0 1 41213
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_855
timestamp 1649977179
transform 1 0 114648 0 1 40261
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_856
timestamp 1649977179
transform 1 0 114240 0 1 36725
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_857
timestamp 1649977179
transform 1 0 114240 0 1 37133
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_858
timestamp 1649977179
transform 1 0 114240 0 1 36861
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_859
timestamp 1649977179
transform 1 0 115600 0 1 41485
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_860
timestamp 1649977179
transform 1 0 115464 0 1 38901
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_861
timestamp 1649977179
transform 1 0 115464 0 1 39173
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_862
timestamp 1649977179
transform 1 0 115464 0 1 37677
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_863
timestamp 1649977179
transform 1 0 115464 0 1 37949
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_864
timestamp 1649977179
transform 1 0 115328 0 1 40125
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_865
timestamp 1649977179
transform 1 0 114240 0 1 40261
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_866
timestamp 1649977179
transform 1 0 114240 0 1 39989
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_867
timestamp 1649977179
transform 1 0 114240 0 1 39581
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_868
timestamp 1649977179
transform 1 0 115192 0 1 40261
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_869
timestamp 1649977179
transform 1 0 114240 0 1 39853
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_870
timestamp 1649977179
transform 1 0 115328 0 1 40669
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_871
timestamp 1649977179
transform 1 0 115328 0 1 40397
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_872
timestamp 1649977179
transform 1 0 115328 0 1 41077
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_873
timestamp 1649977179
transform 1 0 114648 0 1 40669
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_874
timestamp 1649977179
transform 1 0 114648 0 1 40397
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_875
timestamp 1649977179
transform 1 0 115328 0 1 40805
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_876
timestamp 1649977179
transform 1 0 115192 0 1 41077
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_877
timestamp 1649977179
transform 1 0 115192 0 1 40805
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_878
timestamp 1649977179
transform 1 0 115192 0 1 36725
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_879
timestamp 1649977179
transform 1 0 114648 0 1 39989
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_880
timestamp 1649977179
transform 1 0 115056 0 1 37677
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_881
timestamp 1649977179
transform 1 0 114648 0 1 36725
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_882
timestamp 1649977179
transform 1 0 114648 0 1 40805
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_883
timestamp 1649977179
transform 1 0 114648 0 1 41077
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_884
timestamp 1649977179
transform 1 0 115056 0 1 37949
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_885
timestamp 1649977179
transform 1 0 114648 0 1 39581
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_886
timestamp 1649977179
transform 1 0 115464 0 1 36453
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_887
timestamp 1649977179
transform 1 0 114240 0 1 36453
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_888
timestamp 1649977179
transform 1 0 115192 0 1 36453
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_889
timestamp 1649977179
transform 1 0 114648 0 1 36453
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_890
timestamp 1649977179
transform 1 0 135320 0 1 35501
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_891
timestamp 1649977179
transform 1 0 135320 0 1 33869
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_892
timestamp 1649977179
transform 1 0 135320 0 1 32237
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_893
timestamp 1649977179
transform 1 0 135320 0 1 39037
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_894
timestamp 1649977179
transform 1 0 135320 0 1 40805
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_895
timestamp 1649977179
transform 1 0 135320 0 1 37405
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_896
timestamp 1649977179
transform 1 0 119272 0 1 27205
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_897
timestamp 1649977179
transform 1 0 119272 0 1 26661
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_898
timestamp 1649977179
transform 1 0 119272 0 1 25845
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_899
timestamp 1649977179
transform 1 0 119272 0 1 26525
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_900
timestamp 1649977179
transform 1 0 114240 0 1 31285
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_901
timestamp 1649977179
transform 1 0 114648 0 1 31285
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_902
timestamp 1649977179
transform 1 0 119000 0 1 20949
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_903
timestamp 1649977179
transform 1 0 118184 0 1 20949
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_904
timestamp 1649977179
transform 1 0 114240 0 1 20949
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_905
timestamp 1649977179
transform 1 0 116008 0 1 20949
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_906
timestamp 1649977179
transform 1 0 114648 0 1 20949
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_907
timestamp 1649977179
transform 1 0 118592 0 1 20949
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_908
timestamp 1649977179
transform 1 0 117640 0 1 20949
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_909
timestamp 1649977179
transform 1 0 115328 0 1 20949
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_910
timestamp 1649977179
transform 1 0 115192 0 1 20949
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_911
timestamp 1649977179
transform 1 0 62560 0 1 1229
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_912
timestamp 1649977179
transform 1 0 62560 0 1 1637
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_913
timestamp 1649977179
transform 1 0 60792 0 1 1229
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_914
timestamp 1649977179
transform 1 0 67592 0 1 1229
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_915
timestamp 1649977179
transform 1 0 67592 0 1 1637
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_916
timestamp 1649977179
transform 1 0 60792 0 1 1637
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_917
timestamp 1649977179
transform 1 0 65824 0 1 1229
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_918
timestamp 1649977179
transform 1 0 65824 0 1 1637
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_919
timestamp 1649977179
transform 1 0 64328 0 1 1229
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_920
timestamp 1649977179
transform 1 0 64328 0 1 1637
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_921
timestamp 1649977179
transform 1 0 54128 0 1 1229
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_922
timestamp 1649977179
transform 1 0 54128 0 1 1637
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_923
timestamp 1649977179
transform 1 0 52496 0 1 1229
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_924
timestamp 1649977179
transform 1 0 52496 0 1 1637
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_925
timestamp 1649977179
transform 1 0 55488 0 1 1229
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_926
timestamp 1649977179
transform 1 0 55488 0 1 1637
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_927
timestamp 1649977179
transform 1 0 57528 0 1 1229
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_928
timestamp 1649977179
transform 1 0 57528 0 1 1637
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_929
timestamp 1649977179
transform 1 0 59160 0 1 2861
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_930
timestamp 1649977179
transform 1 0 58072 0 1 2861
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_931
timestamp 1649977179
transform 1 0 56984 0 1 2861
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_932
timestamp 1649977179
transform 1 0 55760 0 1 2861
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_933
timestamp 1649977179
transform 1 0 54400 0 1 2861
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_934
timestamp 1649977179
transform 1 0 53312 0 1 2861
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_935
timestamp 1649977179
transform 1 0 52224 0 1 2861
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_936
timestamp 1649977179
transform 1 0 59432 0 1 1229
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_937
timestamp 1649977179
transform 1 0 59432 0 1 1637
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_938
timestamp 1649977179
transform 1 0 51136 0 1 2861
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_939
timestamp 1649977179
transform 1 0 49776 0 1 2861
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_940
timestamp 1649977179
transform 1 0 48688 0 1 2861
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_941
timestamp 1649977179
transform 1 0 47600 0 1 2861
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_942
timestamp 1649977179
transform 1 0 46376 0 1 2861
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_943
timestamp 1649977179
transform 1 0 45288 0 1 2861
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_944
timestamp 1649977179
transform 1 0 43928 0 1 2861
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_945
timestamp 1649977179
transform 1 0 42840 0 1 2861
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_946
timestamp 1649977179
transform 1 0 50728 0 1 1229
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_947
timestamp 1649977179
transform 1 0 50728 0 1 1637
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_948
timestamp 1649977179
transform 1 0 47328 0 1 1229
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_949
timestamp 1649977179
transform 1 0 47328 0 1 1637
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_950
timestamp 1649977179
transform 1 0 45696 0 1 1229
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_951
timestamp 1649977179
transform 1 0 45696 0 1 1637
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_952
timestamp 1649977179
transform 1 0 44200 0 1 1229
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_953
timestamp 1649977179
transform 1 0 44200 0 1 1637
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_954
timestamp 1649977179
transform 1 0 49096 0 1 1229
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_955
timestamp 1649977179
transform 1 0 49096 0 1 1637
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_956
timestamp 1649977179
transform 1 0 41752 0 1 2861
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_957
timestamp 1649977179
transform 1 0 40664 0 1 2861
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_958
timestamp 1649977179
transform 1 0 39440 0 1 2861
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_959
timestamp 1649977179
transform 1 0 38080 0 1 2861
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_960
timestamp 1649977179
transform 1 0 36992 0 1 2861
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_961
timestamp 1649977179
transform 1 0 35904 0 1 2861
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_962
timestamp 1649977179
transform 1 0 34544 0 1 2861
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_963
timestamp 1649977179
transform 1 0 37400 0 1 1229
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_964
timestamp 1649977179
transform 1 0 37400 0 1 1637
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_965
timestamp 1649977179
transform 1 0 42432 0 1 1229
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_966
timestamp 1649977179
transform 1 0 42432 0 1 1637
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_967
timestamp 1649977179
transform 1 0 35768 0 1 1229
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_968
timestamp 1649977179
transform 1 0 35768 0 1 1637
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_969
timestamp 1649977179
transform 1 0 39168 0 1 1229
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_970
timestamp 1649977179
transform 1 0 39712 0 1 549
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_971
timestamp 1649977179
transform 1 0 39712 0 1 2317
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_972
timestamp 1649977179
transform 1 0 39168 0 1 1637
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_973
timestamp 1649977179
transform 1 0 40800 0 1 1229
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_974
timestamp 1649977179
transform 1 0 40800 0 1 1637
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_975
timestamp 1649977179
transform 1 0 43792 0 1 14285
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_976
timestamp 1649977179
transform 1 0 43928 0 1 13469
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_977
timestamp 1649977179
transform 1 0 43928 0 1 11973
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_978
timestamp 1649977179
transform 1 0 48824 0 1 13605
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_979
timestamp 1649977179
transform 1 0 48824 0 1 14285
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_980
timestamp 1649977179
transform 1 0 43792 0 1 11021
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_981
timestamp 1649977179
transform 1 0 43792 0 1 11837
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_982
timestamp 1649977179
transform 1 0 48960 0 1 13469
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_983
timestamp 1649977179
transform 1 0 48960 0 1 11973
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_984
timestamp 1649977179
transform 1 0 48688 0 1 11021
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_985
timestamp 1649977179
transform 1 0 48688 0 1 11837
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_986
timestamp 1649977179
transform 1 0 46512 0 1 12517
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_987
timestamp 1649977179
transform 1 0 46512 0 1 11701
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_988
timestamp 1649977179
transform 1 0 46512 0 1 12245
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_989
timestamp 1649977179
transform 1 0 44064 0 1 12517
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_990
timestamp 1649977179
transform 1 0 43384 0 1 12245
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_991
timestamp 1649977179
transform 1 0 43384 0 1 11429
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_992
timestamp 1649977179
transform 1 0 44064 0 1 13061
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_993
timestamp 1649977179
transform 1 0 43928 0 1 15101
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_994
timestamp 1649977179
transform 1 0 44064 0 1 15101
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_995
timestamp 1649977179
transform 1 0 46240 0 1 13605
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_996
timestamp 1649977179
transform 1 0 46240 0 1 14285
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_997
timestamp 1649977179
transform 1 0 46376 0 1 13469
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_998
timestamp 1649977179
transform 1 0 46376 0 1 11973
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_999
timestamp 1649977179
transform 1 0 46240 0 1 11021
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1000
timestamp 1649977179
transform 1 0 46240 0 1 11837
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1001
timestamp 1649977179
transform 1 0 44064 0 1 13197
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1002
timestamp 1649977179
transform 1 0 51136 0 1 11021
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1003
timestamp 1649977179
transform 1 0 51136 0 1 11837
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1004
timestamp 1649977179
transform 1 0 48960 0 1 15101
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1005
timestamp 1649977179
transform 1 0 49096 0 1 15101
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1006
timestamp 1649977179
transform 1 0 49096 0 1 13197
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1007
timestamp 1649977179
transform 1 0 46512 0 1 15101
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1008
timestamp 1649977179
transform 1 0 46512 0 1 13197
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1009
timestamp 1649977179
transform 1 0 48824 0 1 13061
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1010
timestamp 1649977179
transform 1 0 48824 0 1 12517
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1011
timestamp 1649977179
transform 1 0 48824 0 1 11701
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1012
timestamp 1649977179
transform 1 0 48824 0 1 12245
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1013
timestamp 1649977179
transform 1 0 46512 0 1 13061
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1014
timestamp 1649977179
transform 1 0 46648 0 1 15101
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1015
timestamp 1649977179
transform 1 0 51000 0 1 13061
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1016
timestamp 1649977179
transform 1 0 48280 0 1 13061
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1017
timestamp 1649977179
transform 1 0 45968 0 1 13061
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1018
timestamp 1649977179
transform 1 0 43520 0 1 13061
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1019
timestamp 1649977179
transform 1 0 43792 0 1 13605
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1020
timestamp 1649977179
transform 1 0 39168 0 1 15101
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1021
timestamp 1649977179
transform 1 0 41480 0 1 13197
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1022
timestamp 1649977179
transform 1 0 41480 0 1 12245
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1023
timestamp 1649977179
transform 1 0 38896 0 1 11973
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1024
timestamp 1649977179
transform 1 0 36448 0 1 13469
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1025
timestamp 1649977179
transform 1 0 39032 0 1 15101
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1026
timestamp 1649977179
transform 1 0 39032 0 1 13197
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1027
timestamp 1649977179
transform 1 0 39032 0 1 13061
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1028
timestamp 1649977179
transform 1 0 39032 0 1 12517
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1029
timestamp 1649977179
transform 1 0 38624 0 1 11701
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1030
timestamp 1649977179
transform 1 0 38624 0 1 12245
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1031
timestamp 1649977179
transform 1 0 36312 0 1 11837
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1032
timestamp 1649977179
transform 1 0 36448 0 1 15101
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1033
timestamp 1649977179
transform 1 0 38896 0 1 14285
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1034
timestamp 1649977179
transform 1 0 38896 0 1 13469
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1035
timestamp 1649977179
transform 1 0 36448 0 1 11973
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1036
timestamp 1649977179
transform 1 0 36312 0 1 11021
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1037
timestamp 1649977179
transform 1 0 36584 0 1 15101
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1038
timestamp 1649977179
transform 1 0 36584 0 1 13197
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1039
timestamp 1649977179
transform 1 0 36584 0 1 13061
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1040
timestamp 1649977179
transform 1 0 36584 0 1 12517
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1041
timestamp 1649977179
transform 1 0 36176 0 1 11701
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1042
timestamp 1649977179
transform 1 0 36176 0 1 12245
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1043
timestamp 1649977179
transform 1 0 41480 0 1 13061
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1044
timestamp 1649977179
transform 1 0 36448 0 1 13605
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1045
timestamp 1649977179
transform 1 0 36448 0 1 14285
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1046
timestamp 1649977179
transform 1 0 41480 0 1 12517
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1047
timestamp 1649977179
transform 1 0 41208 0 1 13605
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1048
timestamp 1649977179
transform 1 0 41208 0 1 14285
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1049
timestamp 1649977179
transform 1 0 41344 0 1 13469
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1050
timestamp 1649977179
transform 1 0 41072 0 1 13061
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1051
timestamp 1649977179
transform 1 0 38488 0 1 13061
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1052
timestamp 1649977179
transform 1 0 36040 0 1 13061
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1053
timestamp 1649977179
transform 1 0 41344 0 1 11973
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1054
timestamp 1649977179
transform 1 0 41344 0 1 11021
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1055
timestamp 1649977179
transform 1 0 41344 0 1 11837
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1056
timestamp 1649977179
transform 1 0 41072 0 1 13605
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1057
timestamp 1649977179
transform 1 0 41072 0 1 14285
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1058
timestamp 1649977179
transform 1 0 38896 0 1 13605
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1059
timestamp 1649977179
transform 1 0 41480 0 1 11701
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1060
timestamp 1649977179
transform 1 0 41616 0 1 15101
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1061
timestamp 1649977179
transform 1 0 38760 0 1 11021
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1062
timestamp 1649977179
transform 1 0 38760 0 1 11837
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1063
timestamp 1649977179
transform 1 0 41480 0 1 15101
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1064
timestamp 1649977179
transform 1 0 37264 0 1 19181
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1065
timestamp 1649977179
transform 1 0 38216 0 1 19181
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1066
timestamp 1649977179
transform 1 0 36448 0 1 17005
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1067
timestamp 1649977179
transform 1 0 35632 0 1 18773
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1068
timestamp 1649977179
transform 1 0 34544 0 1 19181
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1069
timestamp 1649977179
transform 1 0 35632 0 1 19181
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1070
timestamp 1649977179
transform 1 0 42432 0 1 18773
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1071
timestamp 1649977179
transform 1 0 42024 0 1 18773
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1072
timestamp 1649977179
transform 1 0 42024 0 1 19181
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1073
timestamp 1649977179
transform 1 0 41208 0 1 19181
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1074
timestamp 1649977179
transform 1 0 41208 0 1 18773
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1075
timestamp 1649977179
transform 1 0 40664 0 1 18773
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1076
timestamp 1649977179
transform 1 0 40664 0 1 19181
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1077
timestamp 1649977179
transform 1 0 39984 0 1 19181
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1078
timestamp 1649977179
transform 1 0 39984 0 1 18773
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1079
timestamp 1649977179
transform 1 0 39440 0 1 18773
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1080
timestamp 1649977179
transform 1 0 39440 0 1 19181
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1081
timestamp 1649977179
transform 1 0 38760 0 1 19181
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1082
timestamp 1649977179
transform 1 0 37264 0 1 18773
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1083
timestamp 1649977179
transform 1 0 39168 0 1 17005
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1084
timestamp 1649977179
transform 1 0 34544 0 1 18773
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1085
timestamp 1649977179
transform 1 0 38760 0 1 18773
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1086
timestamp 1649977179
transform 1 0 41616 0 1 17005
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1087
timestamp 1649977179
transform 1 0 38216 0 1 18773
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1088
timestamp 1649977179
transform 1 0 42432 0 1 19181
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1089
timestamp 1649977179
transform 1 0 48960 0 1 17005
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1090
timestamp 1649977179
transform 1 0 49912 0 1 19181
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1091
timestamp 1649977179
transform 1 0 49912 0 1 18773
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1092
timestamp 1649977179
transform 1 0 46648 0 1 17005
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1093
timestamp 1649977179
transform 1 0 48144 0 1 18773
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1094
timestamp 1649977179
transform 1 0 48144 0 1 19181
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1095
timestamp 1649977179
transform 1 0 47464 0 1 19181
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1096
timestamp 1649977179
transform 1 0 47464 0 1 18773
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1097
timestamp 1649977179
transform 1 0 46920 0 1 18773
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1098
timestamp 1649977179
transform 1 0 46920 0 1 19181
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1099
timestamp 1649977179
transform 1 0 45696 0 1 18773
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1100
timestamp 1649977179
transform 1 0 45696 0 1 19181
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1101
timestamp 1649977179
transform 1 0 44472 0 1 18773
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1102
timestamp 1649977179
transform 1 0 44472 0 1 19181
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1103
timestamp 1649977179
transform 1 0 43384 0 1 19181
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1104
timestamp 1649977179
transform 1 0 43384 0 1 18773
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1105
timestamp 1649977179
transform 1 0 43248 0 1 18773
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1106
timestamp 1649977179
transform 1 0 43248 0 1 19181
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1107
timestamp 1649977179
transform 1 0 44064 0 1 17005
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1108
timestamp 1649977179
transform 1 0 63648 0 1 13605
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1109
timestamp 1649977179
transform 1 0 61608 0 1 15101
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1110
timestamp 1649977179
transform 1 0 61472 0 1 15101
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1111
timestamp 1649977179
transform 1 0 61472 0 1 13061
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1112
timestamp 1649977179
transform 1 0 61336 0 1 13061
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1113
timestamp 1649977179
transform 1 0 61336 0 1 12517
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1114
timestamp 1649977179
transform 1 0 61336 0 1 11701
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1115
timestamp 1649977179
transform 1 0 61336 0 1 12245
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1116
timestamp 1649977179
transform 1 0 61336 0 1 13605
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1117
timestamp 1649977179
transform 1 0 61336 0 1 14285
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1118
timestamp 1649977179
transform 1 0 63784 0 1 13605
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1119
timestamp 1649977179
transform 1 0 63784 0 1 14285
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1120
timestamp 1649977179
transform 1 0 63920 0 1 13469
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1121
timestamp 1649977179
transform 1 0 63920 0 1 11973
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1122
timestamp 1649977179
transform 1 0 63784 0 1 11021
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1123
timestamp 1649977179
transform 1 0 63784 0 1 11837
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1124
timestamp 1649977179
transform 1 0 61200 0 1 13605
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1125
timestamp 1649977179
transform 1 0 61200 0 1 11973
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1126
timestamp 1649977179
transform 1 0 61200 0 1 11021
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1127
timestamp 1649977179
transform 1 0 61200 0 1 11837
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1128
timestamp 1649977179
transform 1 0 61064 0 1 14285
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1129
timestamp 1649977179
transform 1 0 61064 0 1 13605
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1130
timestamp 1649977179
transform 1 0 66232 0 1 13605
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1131
timestamp 1649977179
transform 1 0 66232 0 1 14285
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1132
timestamp 1649977179
transform 1 0 65960 0 1 13061
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1133
timestamp 1649977179
transform 1 0 63512 0 1 13061
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1134
timestamp 1649977179
transform 1 0 60928 0 1 13061
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1135
timestamp 1649977179
transform 1 0 66368 0 1 13469
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1136
timestamp 1649977179
transform 1 0 66368 0 1 11973
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1137
timestamp 1649977179
transform 1 0 66096 0 1 11021
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1138
timestamp 1649977179
transform 1 0 66096 0 1 11837
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1139
timestamp 1649977179
transform 1 0 66640 0 1 15101
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1140
timestamp 1649977179
transform 1 0 66504 0 1 15101
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1141
timestamp 1649977179
transform 1 0 66504 0 1 13197
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1142
timestamp 1649977179
transform 1 0 66504 0 1 13061
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1143
timestamp 1649977179
transform 1 0 66504 0 1 12517
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1144
timestamp 1649977179
transform 1 0 66232 0 1 11701
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1145
timestamp 1649977179
transform 1 0 66232 0 1 12245
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1146
timestamp 1649977179
transform 1 0 63648 0 1 14285
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1147
timestamp 1649977179
transform 1 0 63920 0 1 15101
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1148
timestamp 1649977179
transform 1 0 64056 0 1 15101
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1149
timestamp 1649977179
transform 1 0 64056 0 1 13197
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1150
timestamp 1649977179
transform 1 0 64056 0 1 13061
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1151
timestamp 1649977179
transform 1 0 64056 0 1 12517
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1152
timestamp 1649977179
transform 1 0 63648 0 1 11701
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1153
timestamp 1649977179
transform 1 0 63648 0 1 12245
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1154
timestamp 1649977179
transform 1 0 53856 0 1 13605
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1155
timestamp 1649977179
transform 1 0 53856 0 1 14285
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1156
timestamp 1649977179
transform 1 0 53856 0 1 13469
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1157
timestamp 1649977179
transform 1 0 53856 0 1 11973
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1158
timestamp 1649977179
transform 1 0 53856 0 1 11021
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1159
timestamp 1649977179
transform 1 0 53856 0 1 11837
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1160
timestamp 1649977179
transform 1 0 58344 0 1 14421
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1161
timestamp 1649977179
transform 1 0 56440 0 1 14285
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1162
timestamp 1649977179
transform 1 0 56304 0 1 13469
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1163
timestamp 1649977179
transform 1 0 56304 0 1 11973
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1164
timestamp 1649977179
transform 1 0 56304 0 1 11021
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1165
timestamp 1649977179
transform 1 0 56304 0 1 11837
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1166
timestamp 1649977179
transform 1 0 51408 0 1 13605
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1167
timestamp 1649977179
transform 1 0 51408 0 1 14285
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1168
timestamp 1649977179
transform 1 0 51408 0 1 13469
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1169
timestamp 1649977179
transform 1 0 51408 0 1 11973
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1170
timestamp 1649977179
transform 1 0 58616 0 1 14285
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1171
timestamp 1649977179
transform 1 0 58616 0 1 13605
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1172
timestamp 1649977179
transform 1 0 58480 0 1 13061
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1173
timestamp 1649977179
transform 1 0 56032 0 1 13061
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1174
timestamp 1649977179
transform 1 0 53584 0 1 13061
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1175
timestamp 1649977179
transform 1 0 56440 0 1 13605
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1176
timestamp 1649977179
transform 1 0 58888 0 1 13605
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1177
timestamp 1649977179
transform 1 0 58888 0 1 14285
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1178
timestamp 1649977179
transform 1 0 58888 0 1 13469
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1179
timestamp 1649977179
transform 1 0 59160 0 1 15101
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1180
timestamp 1649977179
transform 1 0 59024 0 1 15101
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1181
timestamp 1649977179
transform 1 0 59024 0 1 13197
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1182
timestamp 1649977179
transform 1 0 59024 0 1 13061
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1183
timestamp 1649977179
transform 1 0 59024 0 1 12517
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1184
timestamp 1649977179
transform 1 0 59024 0 1 11701
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1185
timestamp 1649977179
transform 1 0 59024 0 1 12245
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1186
timestamp 1649977179
transform 1 0 58888 0 1 11973
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1187
timestamp 1649977179
transform 1 0 56440 0 1 15101
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1188
timestamp 1649977179
transform 1 0 56576 0 1 15101
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1189
timestamp 1649977179
transform 1 0 56576 0 1 13197
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1190
timestamp 1649977179
transform 1 0 56440 0 1 13061
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1191
timestamp 1649977179
transform 1 0 56440 0 1 12517
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1192
timestamp 1649977179
transform 1 0 56440 0 1 11701
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1193
timestamp 1649977179
transform 1 0 56440 0 1 12245
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1194
timestamp 1649977179
transform 1 0 58752 0 1 11021
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1195
timestamp 1649977179
transform 1 0 54128 0 1 15101
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1196
timestamp 1649977179
transform 1 0 53992 0 1 15101
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1197
timestamp 1649977179
transform 1 0 53992 0 1 13197
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1198
timestamp 1649977179
transform 1 0 53992 0 1 13061
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1199
timestamp 1649977179
transform 1 0 53992 0 1 12517
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1200
timestamp 1649977179
transform 1 0 53992 0 1 11701
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1201
timestamp 1649977179
transform 1 0 53992 0 1 12245
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1202
timestamp 1649977179
transform 1 0 58752 0 1 11837
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1203
timestamp 1649977179
transform 1 0 51408 0 1 15101
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1204
timestamp 1649977179
transform 1 0 51544 0 1 15101
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1205
timestamp 1649977179
transform 1 0 51544 0 1 13197
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1206
timestamp 1649977179
transform 1 0 51544 0 1 13061
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1207
timestamp 1649977179
transform 1 0 51544 0 1 12517
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1208
timestamp 1649977179
transform 1 0 53720 0 1 19181
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1209
timestamp 1649977179
transform 1 0 53720 0 1 18773
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1210
timestamp 1649977179
transform 1 0 53176 0 1 18773
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1211
timestamp 1649977179
transform 1 0 53176 0 1 19181
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1212
timestamp 1649977179
transform 1 0 51952 0 1 18773
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1213
timestamp 1649977179
transform 1 0 51952 0 1 19181
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1214
timestamp 1649977179
transform 1 0 54944 0 1 19181
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1215
timestamp 1649977179
transform 1 0 54944 0 1 18773
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1216
timestamp 1649977179
transform 1 0 55624 0 1 19181
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1217
timestamp 1649977179
transform 1 0 59432 0 1 18773
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1218
timestamp 1649977179
transform 1 0 59432 0 1 19181
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1219
timestamp 1649977179
transform 1 0 59160 0 1 17005
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1220
timestamp 1649977179
transform 1 0 56440 0 1 17005
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1221
timestamp 1649977179
transform 1 0 54128 0 1 17005
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1222
timestamp 1649977179
transform 1 0 51544 0 1 17005
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1223
timestamp 1649977179
transform 1 0 54400 0 1 18773
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1224
timestamp 1649977179
transform 1 0 54400 0 1 19181
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1225
timestamp 1649977179
transform 1 0 58344 0 1 18637
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1226
timestamp 1649977179
transform 1 0 58208 0 1 18773
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1227
timestamp 1649977179
transform 1 0 58208 0 1 19181
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1228
timestamp 1649977179
transform 1 0 57392 0 1 19181
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1229
timestamp 1649977179
transform 1 0 57392 0 1 18773
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1230
timestamp 1649977179
transform 1 0 56168 0 1 19181
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1231
timestamp 1649977179
transform 1 0 56168 0 1 18773
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1232
timestamp 1649977179
transform 1 0 55624 0 1 18773
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1233
timestamp 1649977179
transform 1 0 66640 0 1 17005
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1234
timestamp 1649977179
transform 1 0 63920 0 1 17005
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1235
timestamp 1649977179
transform 1 0 61608 0 1 17005
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1236
timestamp 1649977179
transform 1 0 67456 0 1 19181
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1237
timestamp 1649977179
transform 1 0 67456 0 1 18773
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1238
timestamp 1649977179
transform 1 0 66912 0 1 18773
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1239
timestamp 1649977179
transform 1 0 66912 0 1 19181
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1240
timestamp 1649977179
transform 1 0 66232 0 1 19181
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1241
timestamp 1649977179
transform 1 0 66232 0 1 18773
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1242
timestamp 1649977179
transform 1 0 64464 0 1 18773
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1243
timestamp 1649977179
transform 1 0 64464 0 1 19181
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1244
timestamp 1649977179
transform 1 0 63104 0 1 18773
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1245
timestamp 1649977179
transform 1 0 63104 0 1 19181
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1246
timestamp 1649977179
transform 1 0 62424 0 1 19181
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1247
timestamp 1649977179
transform 1 0 62424 0 1 18773
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1248
timestamp 1649977179
transform 1 0 61880 0 1 18773
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1249
timestamp 1649977179
transform 1 0 61880 0 1 19181
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1250
timestamp 1649977179
transform 1 0 60792 0 1 19181
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1251
timestamp 1649977179
transform 1 0 60792 0 1 18773
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1252
timestamp 1649977179
transform 1 0 60656 0 1 18773
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1253
timestamp 1649977179
transform 1 0 60656 0 1 19181
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1254
timestamp 1649977179
transform 1 0 59976 0 1 19181
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1255
timestamp 1649977179
transform 1 0 59976 0 1 18773
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1256
timestamp 1649977179
transform 1 0 51272 0 1 19181
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1257
timestamp 1649977179
transform 1 0 51272 0 1 18773
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1258
timestamp 1649977179
transform 1 0 51272 0 1 11701
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1259
timestamp 1649977179
transform 1 0 51272 0 1 12245
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1260
timestamp 1649977179
transform 1 0 27336 0 1 1229
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1261
timestamp 1649977179
transform 1 0 27336 0 1 1637
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1262
timestamp 1649977179
transform 1 0 33456 0 1 2861
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1263
timestamp 1649977179
transform 1 0 32368 0 1 2861
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1264
timestamp 1649977179
transform 1 0 31280 0 1 2861
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1265
timestamp 1649977179
transform 1 0 30056 0 1 2861
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1266
timestamp 1649977179
transform 1 0 28696 0 1 2861
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1267
timestamp 1649977179
transform 1 0 27608 0 1 2861
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1268
timestamp 1649977179
transform 1 0 26520 0 1 2861
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1269
timestamp 1649977179
transform 1 0 34000 0 1 1229
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1270
timestamp 1649977179
transform 1 0 34000 0 1 1637
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1271
timestamp 1649977179
transform 1 0 28968 0 1 1229
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1272
timestamp 1649977179
transform 1 0 28968 0 1 1637
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1273
timestamp 1649977179
transform 1 0 32096 0 1 1229
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1274
timestamp 1649977179
transform 1 0 32096 0 1 1637
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1275
timestamp 1649977179
transform 1 0 30464 0 1 1229
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1276
timestamp 1649977179
transform 1 0 30464 0 1 1637
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1277
timestamp 1649977179
transform 1 0 25704 0 1 1229
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1278
timestamp 1649977179
transform 1 0 25704 0 1 1637
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1279
timestamp 1649977179
transform 1 0 23936 0 1 1229
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1280
timestamp 1649977179
transform 1 0 23936 0 1 1637
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1281
timestamp 1649977179
transform 1 0 21760 0 1 2861
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1282
timestamp 1649977179
transform 1 0 20536 0 1 2861
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1283
timestamp 1649977179
transform 1 0 19584 0 1 2861
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1284
timestamp 1649977179
transform 1 0 18224 0 1 2861
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1285
timestamp 1649977179
transform 1 0 17408 0 1 1229
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1286
timestamp 1649977179
transform 1 0 25432 0 1 2861
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1287
timestamp 1649977179
transform 1 0 24208 0 1 2861
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1288
timestamp 1649977179
transform 1 0 23120 0 1 2861
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1289
timestamp 1649977179
transform 1 0 17408 0 1 1637
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1290
timestamp 1649977179
transform 1 0 22168 0 1 1229
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1291
timestamp 1649977179
transform 1 0 22168 0 1 1637
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1292
timestamp 1649977179
transform 1 0 20808 0 1 1229
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1293
timestamp 1649977179
transform 1 0 20808 0 1 1637
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1294
timestamp 1649977179
transform 1 0 20264 0 1 1773
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1295
timestamp 1649977179
transform 1 0 20264 0 1 3677
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1296
timestamp 1649977179
transform 1 0 19040 0 1 1229
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1297
timestamp 1649977179
transform 1 0 19040 0 1 1637
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1298
timestamp 1649977179
transform 1 0 28152 0 1 9525
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1299
timestamp 1649977179
transform 1 0 15504 0 1 1229
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1300
timestamp 1649977179
transform 1 0 15504 0 1 1637
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1301
timestamp 1649977179
transform 1 0 17136 0 1 2861
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1302
timestamp 1649977179
transform 1 0 16048 0 1 2861
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1303
timestamp 1649977179
transform 1 0 16320 0 1 3813
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1304
timestamp 1649977179
transform 1 0 14008 0 1 1229
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1305
timestamp 1649977179
transform 1 0 14008 0 1 1637
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1306
timestamp 1649977179
transform 1 0 12104 0 1 1229
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1307
timestamp 1649977179
transform 1 0 12104 0 1 1637
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1308
timestamp 1649977179
transform 1 0 10472 0 1 1229
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1309
timestamp 1649977179
transform 1 0 10472 0 1 1637
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1310
timestamp 1649977179
transform 1 0 7072 0 1 1229
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1311
timestamp 1649977179
transform 1 0 7072 0 1 1637
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1312
timestamp 1649977179
transform 1 0 5576 0 1 1229
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1313
timestamp 1649977179
transform 1 0 5576 0 1 1637
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1314
timestamp 1649977179
transform 1 0 3808 0 1 1229
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1315
timestamp 1649977179
transform 1 0 3808 0 1 1637
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1316
timestamp 1649977179
transform 1 0 2040 0 1 1229
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1317
timestamp 1649977179
transform 1 0 2040 0 1 1637
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1318
timestamp 1649977179
transform 1 0 1224 0 1 3813
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1319
timestamp 1649977179
transform 1 0 1224 0 1 10477
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1320
timestamp 1649977179
transform 1 0 1224 0 1 7213
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1321
timestamp 1649977179
transform 1 0 1224 0 1 8709
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1322
timestamp 1649977179
transform 1 0 544 0 1 10205
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1323
timestamp 1649977179
transform 1 0 544 0 1 7621
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1324
timestamp 1649977179
transform 1 0 14688 0 1 10477
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1325
timestamp 1649977179
transform 1 0 14688 0 1 10341
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1326
timestamp 1649977179
transform 1 0 14688 0 1 7621
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1327
timestamp 1649977179
transform 1 0 16320 0 1 8981
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1328
timestamp 1649977179
transform 1 0 14552 0 1 9117
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1329
timestamp 1649977179
transform 1 0 8704 0 1 1229
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1330
timestamp 1649977179
transform 1 0 8704 0 1 1637
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1331
timestamp 1649977179
transform 1 0 1224 0 1 5445
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1332
timestamp 1649977179
transform 1 0 14552 0 1 11701
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1333
timestamp 1649977179
transform 1 0 14552 0 1 14557
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1334
timestamp 1649977179
transform 1 0 14552 0 1 14693
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1335
timestamp 1649977179
transform 1 0 14688 0 1 13333
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1336
timestamp 1649977179
transform 1 0 14688 0 1 13197
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1337
timestamp 1649977179
transform 1 0 14552 0 1 11973
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1338
timestamp 1649977179
transform 1 0 3128 0 1 13333
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1339
timestamp 1649977179
transform 1 0 3128 0 1 13741
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1340
timestamp 1649977179
transform 1 0 1224 0 1 15509
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1341
timestamp 1649977179
transform 1 0 3128 0 1 15509
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1342
timestamp 1649977179
transform 1 0 1224 0 1 12245
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1343
timestamp 1649977179
transform 1 0 1224 0 1 13877
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1344
timestamp 1649977179
transform 1 0 544 0 1 14693
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1345
timestamp 1649977179
transform 1 0 1224 0 1 17005
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1346
timestamp 1649977179
transform 1 0 1224 0 1 18773
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1347
timestamp 1649977179
transform 1 0 3128 0 1 16053
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1348
timestamp 1649977179
transform 1 0 1224 0 1 20541
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1349
timestamp 1649977179
transform 1 0 2531 0 1 17893
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1350
timestamp 1649977179
transform 1 0 3672 0 1 17549
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1351
timestamp 1649977179
transform 1 0 3672 0 1 20405
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1352
timestamp 1649977179
transform 1 0 3808 0 1 20405
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1353
timestamp 1649977179
transform 1 0 14552 0 1 17413
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1354
timestamp 1649977179
transform 1 0 16592 0 1 20133
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1355
timestamp 1649977179
transform 1 0 16592 0 1 19045
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1356
timestamp 1649977179
transform 1 0 14688 0 1 16189
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1357
timestamp 1649977179
transform 1 0 14688 0 1 18773
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1358
timestamp 1649977179
transform 1 0 14688 0 1 16053
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1359
timestamp 1649977179
transform 1 0 17000 0 1 20133
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1360
timestamp 1649977179
transform 1 0 17000 0 1 17549
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1361
timestamp 1649977179
transform 1 0 28560 0 1 11021
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1362
timestamp 1649977179
transform 1 0 33864 0 1 13605
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1363
timestamp 1649977179
transform 1 0 33864 0 1 14285
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1364
timestamp 1649977179
transform 1 0 34000 0 1 13469
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1365
timestamp 1649977179
transform 1 0 34000 0 1 11973
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1366
timestamp 1649977179
transform 1 0 33864 0 1 11021
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1367
timestamp 1649977179
transform 1 0 29104 0 1 15101
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1368
timestamp 1649977179
transform 1 0 33864 0 1 11837
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1369
timestamp 1649977179
transform 1 0 29104 0 1 13197
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1370
timestamp 1649977179
transform 1 0 29104 0 1 13061
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1371
timestamp 1649977179
transform 1 0 29104 0 1 12517
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1372
timestamp 1649977179
transform 1 0 28832 0 1 11701
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1373
timestamp 1649977179
transform 1 0 34000 0 1 15101
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1374
timestamp 1649977179
transform 1 0 34136 0 1 15101
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1375
timestamp 1649977179
transform 1 0 34136 0 1 13197
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1376
timestamp 1649977179
transform 1 0 33592 0 1 14285
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1377
timestamp 1649977179
transform 1 0 33864 0 1 13061
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1378
timestamp 1649977179
transform 1 0 33592 0 1 13605
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1379
timestamp 1649977179
transform 1 0 31416 0 1 13605
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1380
timestamp 1649977179
transform 1 0 33864 0 1 12517
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1381
timestamp 1649977179
transform 1 0 31416 0 1 14285
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1382
timestamp 1649977179
transform 1 0 31280 0 1 13469
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1383
timestamp 1649977179
transform 1 0 31280 0 1 11973
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1384
timestamp 1649977179
transform 1 0 31144 0 1 11021
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1385
timestamp 1649977179
transform 1 0 31144 0 1 11837
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1386
timestamp 1649977179
transform 1 0 33456 0 1 11701
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1387
timestamp 1649977179
transform 1 0 33456 0 1 12245
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1388
timestamp 1649977179
transform 1 0 28832 0 1 12245
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1389
timestamp 1649977179
transform 1 0 31688 0 1 15101
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1390
timestamp 1649977179
transform 1 0 31552 0 1 15101
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1391
timestamp 1649977179
transform 1 0 31552 0 1 13197
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1392
timestamp 1649977179
transform 1 0 31416 0 1 13061
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1393
timestamp 1649977179
transform 1 0 28832 0 1 13605
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1394
timestamp 1649977179
transform 1 0 28832 0 1 14285
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1395
timestamp 1649977179
transform 1 0 31416 0 1 12517
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1396
timestamp 1649977179
transform 1 0 31416 0 1 11701
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1397
timestamp 1649977179
transform 1 0 28968 0 1 13469
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1398
timestamp 1649977179
transform 1 0 28968 0 1 11973
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1399
timestamp 1649977179
transform 1 0 28696 0 1 11021
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1400
timestamp 1649977179
transform 1 0 28696 0 1 11837
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1401
timestamp 1649977179
transform 1 0 31416 0 1 12245
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1402
timestamp 1649977179
transform 1 0 28152 0 1 11293
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1403
timestamp 1649977179
transform 1 0 33592 0 1 13061
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1404
timestamp 1649977179
transform 1 0 30736 0 1 13061
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1405
timestamp 1649977179
transform 1 0 28288 0 1 13061
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1406
timestamp 1649977179
transform 1 0 28968 0 1 15101
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1407
timestamp 1649977179
transform 1 0 20264 0 1 14285
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1408
timestamp 1649977179
transform 1 0 20264 0 1 11701
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1409
timestamp 1649977179
transform 1 0 21216 0 1 13061
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1410
timestamp 1649977179
transform 1 0 21352 0 1 14557
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1411
timestamp 1649977179
transform 1 0 20944 0 1 20541
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1412
timestamp 1649977179
transform 1 0 21352 0 1 20677
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1413
timestamp 1649977179
transform 1 0 21352 0 1 20269
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1414
timestamp 1649977179
transform 1 0 22440 0 1 19725
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1415
timestamp 1649977179
transform 1 0 22440 0 1 20133
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1416
timestamp 1649977179
transform 1 0 22440 0 1 20269
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1417
timestamp 1649977179
transform 1 0 22440 0 1 20541
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1418
timestamp 1649977179
transform 1 0 20944 0 1 20269
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1419
timestamp 1649977179
transform 1 0 21352 0 1 20541
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1420
timestamp 1649977179
transform 1 0 22440 0 1 19589
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1421
timestamp 1649977179
transform 1 0 19176 0 1 20269
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1422
timestamp 1649977179
transform 1 0 22168 0 1 20541
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1423
timestamp 1649977179
transform 1 0 22168 0 1 20269
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1424
timestamp 1649977179
transform 1 0 18632 0 1 20269
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1425
timestamp 1649977179
transform 1 0 18360 0 1 20269
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1426
timestamp 1649977179
transform 1 0 22440 0 1 20677
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1427
timestamp 1649977179
transform 1 0 17816 0 1 20269
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1428
timestamp 1649977179
transform 1 0 21352 0 1 17141
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1429
timestamp 1649977179
transform 1 0 21216 0 1 17277
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1430
timestamp 1649977179
transform 1 0 21760 0 1 20269
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1431
timestamp 1649977179
transform 1 0 21760 0 1 20541
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1432
timestamp 1649977179
transform 1 0 21760 0 1 20677
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1433
timestamp 1649977179
transform 1 0 21080 0 1 20133
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1434
timestamp 1649977179
transform 1 0 22032 0 1 20677
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1435
timestamp 1649977179
transform 1 0 20808 0 1 20677
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1436
timestamp 1649977179
transform 1 0 28288 0 1 19181
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1437
timestamp 1649977179
transform 1 0 26928 0 1 19317
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1438
timestamp 1649977179
transform 1 0 26928 0 1 19589
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1439
timestamp 1649977179
transform 1 0 33728 0 1 19181
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1440
timestamp 1649977179
transform 1 0 33728 0 1 18773
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1441
timestamp 1649977179
transform 1 0 33184 0 1 18773
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1442
timestamp 1649977179
transform 1 0 33184 0 1 19181
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1443
timestamp 1649977179
transform 1 0 32504 0 1 19181
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1444
timestamp 1649977179
transform 1 0 32504 0 1 18773
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1445
timestamp 1649977179
transform 1 0 30736 0 1 18773
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1446
timestamp 1649977179
transform 1 0 30736 0 1 19181
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1447
timestamp 1649977179
transform 1 0 29512 0 1 18773
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1448
timestamp 1649977179
transform 1 0 29512 0 1 19181
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1449
timestamp 1649977179
transform 1 0 28560 0 1 18773
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1450
timestamp 1649977179
transform 1 0 28560 0 1 19181
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1451
timestamp 1649977179
transform 1 0 28288 0 1 18773
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1452
timestamp 1649977179
transform 1 0 28968 0 1 17141
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1453
timestamp 1649977179
transform 1 0 28968 0 1 19725
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1454
timestamp 1649977179
transform 1 0 34000 0 1 17005
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1455
timestamp 1649977179
transform 1 0 31688 0 1 17005
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1456
timestamp 1649977179
transform 1 0 28968 0 1 17005
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1457
timestamp 1649977179
transform 1 0 22440 0 1 15781
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1458
timestamp 1649977179
transform 1 0 21216 0 1 15781
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1459
timestamp 1649977179
transform 1 0 28560 0 1 10613
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1460
timestamp 1649977179
transform 1 0 27472 0 1 22445
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1461
timestamp 1649977179
transform 1 0 27608 0 1 23941
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1462
timestamp 1649977179
transform 1 0 27608 0 1 23669
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1463
timestamp 1649977179
transform 1 0 27472 0 1 23261
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1464
timestamp 1649977179
transform 1 0 27472 0 1 23669
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1465
timestamp 1649977179
transform 1 0 27336 0 1 22037
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1466
timestamp 1649977179
transform 1 0 27336 0 1 22853
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1467
timestamp 1649977179
transform 1 0 27336 0 1 22309
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1468
timestamp 1649977179
transform 1 0 27336 0 1 23125
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1469
timestamp 1649977179
transform 1 0 27472 0 1 25981
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1470
timestamp 1649977179
transform 1 0 27472 0 1 22717
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1471
timestamp 1649977179
transform 1 0 21760 0 1 21765
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1472
timestamp 1649977179
transform 1 0 21760 0 1 21493
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1473
timestamp 1649977179
transform 1 0 21624 0 1 21085
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1474
timestamp 1649977179
transform 1 0 21624 0 1 21357
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1475
timestamp 1649977179
transform 1 0 22168 0 1 21493
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1476
timestamp 1649977179
transform 1 0 22168 0 1 21085
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1477
timestamp 1649977179
transform 1 0 22168 0 1 21357
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1478
timestamp 1649977179
transform 1 0 22440 0 1 21493
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1479
timestamp 1649977179
transform 1 0 22440 0 1 21357
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1480
timestamp 1649977179
transform 1 0 22440 0 1 21085
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1481
timestamp 1649977179
transform 1 0 22440 0 1 21765
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1482
timestamp 1649977179
transform 1 0 22168 0 1 21765
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1483
timestamp 1649977179
transform 1 0 21624 0 1 22989
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1484
timestamp 1649977179
transform 1 0 22440 0 1 23397
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1485
timestamp 1649977179
transform 1 0 21624 0 1 23261
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1486
timestamp 1649977179
transform 1 0 21624 0 1 22581
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1487
timestamp 1649977179
transform 1 0 22168 0 1 23397
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1488
timestamp 1649977179
transform 1 0 22576 0 1 23261
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1489
timestamp 1649977179
transform 1 0 22576 0 1 22989
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1490
timestamp 1649977179
transform 1 0 22032 0 1 23261
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1491
timestamp 1649977179
transform 1 0 22032 0 1 22989
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1492
timestamp 1649977179
transform 1 0 21624 0 1 22309
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1493
timestamp 1649977179
transform 1 0 20944 0 1 21357
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1494
timestamp 1649977179
transform 1 0 21352 0 1 21493
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1495
timestamp 1649977179
transform 1 0 19040 0 1 23261
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1496
timestamp 1649977179
transform 1 0 21352 0 1 22989
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1497
timestamp 1649977179
transform 1 0 18360 0 1 21085
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1498
timestamp 1649977179
transform 1 0 18224 0 1 23397
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1499
timestamp 1649977179
transform 1 0 21352 0 1 23261
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1500
timestamp 1649977179
transform 1 0 18360 0 1 22445
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1501
timestamp 1649977179
transform 1 0 18632 0 1 23261
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1502
timestamp 1649977179
transform 1 0 21352 0 1 21765
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1503
timestamp 1649977179
transform 1 0 18632 0 1 22717
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1504
timestamp 1649977179
transform 1 0 20944 0 1 22717
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1505
timestamp 1649977179
transform 1 0 17680 0 1 23397
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1506
timestamp 1649977179
transform 1 0 20944 0 1 22989
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1507
timestamp 1649977179
transform 1 0 20808 0 1 22309
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1508
timestamp 1649977179
transform 1 0 18224 0 1 23261
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1509
timestamp 1649977179
transform 1 0 18632 0 1 22445
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1510
timestamp 1649977179
transform 1 0 18632 0 1 21085
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1511
timestamp 1649977179
transform 1 0 20808 0 1 22581
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1512
timestamp 1649977179
transform 1 0 18224 0 1 22717
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1513
timestamp 1649977179
transform 1 0 20944 0 1 22173
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1514
timestamp 1649977179
transform 1 0 20944 0 1 21901
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1515
timestamp 1649977179
transform 1 0 19040 0 1 22717
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1516
timestamp 1649977179
transform 1 0 20944 0 1 21765
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1517
timestamp 1649977179
transform 1 0 20944 0 1 21493
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1518
timestamp 1649977179
transform 1 0 20944 0 1 21085
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1519
timestamp 1649977179
transform 1 0 20808 0 1 24621
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1520
timestamp 1649977179
transform 1 0 20808 0 1 24893
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1521
timestamp 1649977179
transform 1 0 18224 0 1 25845
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1522
timestamp 1649977179
transform 1 0 20808 0 1 25301
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1523
timestamp 1649977179
transform 1 0 20808 0 1 25029
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1524
timestamp 1649977179
transform 1 0 18768 0 1 25029
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1525
timestamp 1649977179
transform 1 0 18768 0 1 25709
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1526
timestamp 1649977179
transform 1 0 17408 0 1 25029
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1527
timestamp 1649977179
transform 1 0 20808 0 1 25845
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1528
timestamp 1649977179
transform 1 0 21352 0 1 25301
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1529
timestamp 1649977179
transform 1 0 21216 0 1 23805
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1530
timestamp 1649977179
transform 1 0 21216 0 1 24077
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1531
timestamp 1649977179
transform 1 0 20808 0 1 25709
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1532
timestamp 1649977179
transform 1 0 17544 0 1 25845
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1533
timestamp 1649977179
transform 1 0 20944 0 1 24485
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1534
timestamp 1649977179
transform 1 0 17408 0 1 25709
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1535
timestamp 1649977179
transform 1 0 18632 0 1 25845
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1536
timestamp 1649977179
transform 1 0 21352 0 1 25029
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1537
timestamp 1649977179
transform 1 0 20944 0 1 24213
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1538
timestamp 1649977179
transform 1 0 20808 0 1 25437
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1539
timestamp 1649977179
transform 1 0 18224 0 1 24893
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1540
timestamp 1649977179
transform 1 0 18224 0 1 25029
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1541
timestamp 1649977179
transform 1 0 18224 0 1 25709
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1542
timestamp 1649977179
transform 1 0 19176 0 1 25709
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1543
timestamp 1649977179
transform 1 0 19176 0 1 25029
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1544
timestamp 1649977179
transform 1 0 17680 0 1 24893
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1545
timestamp 1649977179
transform 1 0 22168 0 1 25709
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1546
timestamp 1649977179
transform 1 0 22440 0 1 24077
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1547
timestamp 1649977179
transform 1 0 22440 0 1 23805
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1548
timestamp 1649977179
transform 1 0 22032 0 1 23805
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1549
timestamp 1649977179
transform 1 0 22032 0 1 24077
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1550
timestamp 1649977179
transform 1 0 22168 0 1 25301
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1551
timestamp 1649977179
transform 1 0 22576 0 1 25845
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1552
timestamp 1649977179
transform 1 0 22440 0 1 23669
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1553
timestamp 1649977179
transform 1 0 22168 0 1 25029
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1554
timestamp 1649977179
transform 1 0 22168 0 1 24621
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1555
timestamp 1649977179
transform 1 0 22168 0 1 23669
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1556
timestamp 1649977179
transform 1 0 22168 0 1 24893
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1557
timestamp 1649977179
transform 1 0 22440 0 1 24213
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1558
timestamp 1649977179
transform 1 0 22440 0 1 24485
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1559
timestamp 1649977179
transform 1 0 22576 0 1 24893
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1560
timestamp 1649977179
transform 1 0 22576 0 1 24621
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1561
timestamp 1649977179
transform 1 0 22032 0 1 24485
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1562
timestamp 1649977179
transform 1 0 22440 0 1 25029
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1563
timestamp 1649977179
transform 1 0 22440 0 1 25301
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1564
timestamp 1649977179
transform 1 0 22576 0 1 25709
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1565
timestamp 1649977179
transform 1 0 22576 0 1 25437
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1566
timestamp 1649977179
transform 1 0 22032 0 1 24213
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1567
timestamp 1649977179
transform 1 0 21896 0 1 24893
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1568
timestamp 1649977179
transform 1 0 21896 0 1 24621
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1569
timestamp 1649977179
transform 1 0 21760 0 1 25029
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1570
timestamp 1649977179
transform 1 0 21760 0 1 25301
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1571
timestamp 1649977179
transform 1 0 21624 0 1 24485
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1572
timestamp 1649977179
transform 1 0 21624 0 1 24213
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1573
timestamp 1649977179
transform 1 0 22168 0 1 25437
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1574
timestamp 1649977179
transform 1 0 22168 0 1 25845
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1575
timestamp 1649977179
transform 1 0 21488 0 1 25301
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1576
timestamp 1649977179
transform 1 0 21488 0 1 24077
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1577
timestamp 1649977179
transform 1 0 21488 0 1 23805
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1578
timestamp 1649977179
transform 1 0 21488 0 1 25029
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1579
timestamp 1649977179
transform 1 0 21488 0 1 22717
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1580
timestamp 1649977179
transform 1 0 21488 0 1 22989
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1581
timestamp 1649977179
transform 1 0 21488 0 1 21765
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1582
timestamp 1649977179
transform 1 0 21488 0 1 21493
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1583
timestamp 1649977179
transform 1 0 22168 0 1 29789
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1584
timestamp 1649977179
transform 1 0 22440 0 1 29653
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1585
timestamp 1649977179
transform 1 0 22440 0 1 29381
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1586
timestamp 1649977179
transform 1 0 22168 0 1 30061
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1587
timestamp 1649977179
transform 1 0 17680 0 1 26253
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1588
timestamp 1649977179
transform 1 0 18360 0 1 27205
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1589
timestamp 1649977179
transform 1 0 17680 0 1 26525
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1590
timestamp 1649977179
transform 1 0 18360 0 1 26661
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1591
timestamp 1649977179
transform 1 0 21352 0 1 28429
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1592
timestamp 1649977179
transform 1 0 22576 0 1 29245
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1593
timestamp 1649977179
transform 1 0 22576 0 1 28973
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1594
timestamp 1649977179
transform 1 0 22576 0 1 29789
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1595
timestamp 1649977179
transform 1 0 22576 0 1 30061
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1596
timestamp 1649977179
transform 1 0 22576 0 1 27613
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1597
timestamp 1649977179
transform 1 0 22576 0 1 27341
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1598
timestamp 1649977179
transform 1 0 20944 0 1 28837
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1599
timestamp 1649977179
transform 1 0 20944 0 1 28565
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1600
timestamp 1649977179
transform 1 0 22576 0 1 28837
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1601
timestamp 1649977179
transform 1 0 22576 0 1 28565
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1602
timestamp 1649977179
transform 1 0 20944 0 1 28157
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1603
timestamp 1649977179
transform 1 0 20944 0 1 28429
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1604
timestamp 1649977179
transform 1 0 17544 0 1 26525
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1605
timestamp 1649977179
transform 1 0 18224 0 1 26389
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1606
timestamp 1649977179
transform 1 0 17408 0 1 26661
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1607
timestamp 1649977179
transform 1 0 20808 0 1 28973
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1608
timestamp 1649977179
transform 1 0 20808 0 1 29245
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1609
timestamp 1649977179
transform 1 0 20808 0 1 29653
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1610
timestamp 1649977179
transform 1 0 22440 0 1 27749
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1611
timestamp 1649977179
transform 1 0 22440 0 1 28021
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1612
timestamp 1649977179
transform 1 0 22440 0 1 28429
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1613
timestamp 1649977179
transform 1 0 22440 0 1 28157
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1614
timestamp 1649977179
transform 1 0 20808 0 1 29381
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1615
timestamp 1649977179
transform 1 0 17408 0 1 27205
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1616
timestamp 1649977179
transform 1 0 22168 0 1 29245
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1617
timestamp 1649977179
transform 1 0 22168 0 1 28973
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1618
timestamp 1649977179
transform 1 0 21216 0 1 26253
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1619
timestamp 1649977179
transform 1 0 21216 0 1 26525
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1620
timestamp 1649977179
transform 1 0 21488 0 1 28429
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1621
timestamp 1649977179
transform 1 0 21488 0 1 28157
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1622
timestamp 1649977179
transform 1 0 22032 0 1 28565
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1623
timestamp 1649977179
transform 1 0 21624 0 1 28837
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1624
timestamp 1649977179
transform 1 0 21624 0 1 28565
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1625
timestamp 1649977179
transform 1 0 22032 0 1 28837
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1626
timestamp 1649977179
transform 1 0 21760 0 1 30877
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1627
timestamp 1649977179
transform 1 0 21760 0 1 31149
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1628
timestamp 1649977179
transform 1 0 21760 0 1 28973
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1629
timestamp 1649977179
transform 1 0 21760 0 1 29245
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1630
timestamp 1649977179
transform 1 0 20944 0 1 29789
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1631
timestamp 1649977179
transform 1 0 20944 0 1 30061
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1632
timestamp 1649977179
transform 1 0 17816 0 1 27477
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1633
timestamp 1649977179
transform 1 0 21760 0 1 28021
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1634
timestamp 1649977179
transform 1 0 21760 0 1 27749
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1635
timestamp 1649977179
transform 1 0 17816 0 1 29109
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1636
timestamp 1649977179
transform 1 0 21896 0 1 26525
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1637
timestamp 1649977179
transform 1 0 21896 0 1 26253
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1638
timestamp 1649977179
transform 1 0 20808 0 1 26253
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1639
timestamp 1649977179
transform 1 0 20808 0 1 26525
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1640
timestamp 1649977179
transform 1 0 20808 0 1 26933
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1641
timestamp 1649977179
transform 1 0 21352 0 1 30469
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1642
timestamp 1649977179
transform 1 0 21352 0 1 30197
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1643
timestamp 1649977179
transform 1 0 20808 0 1 26661
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1644
timestamp 1649977179
transform 1 0 21760 0 1 29381
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1645
timestamp 1649977179
transform 1 0 21760 0 1 29653
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1646
timestamp 1649977179
transform 1 0 21352 0 1 28157
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1647
timestamp 1649977179
transform 1 0 18904 0 1 28021
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1648
timestamp 1649977179
transform 1 0 18904 0 1 27341
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1649
timestamp 1649977179
transform 1 0 20808 0 1 30605
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1650
timestamp 1649977179
transform 1 0 20808 0 1 30877
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1651
timestamp 1649977179
transform 1 0 21488 0 1 29653
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1652
timestamp 1649977179
transform 1 0 21488 0 1 29381
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1653
timestamp 1649977179
transform 1 0 22032 0 1 29381
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1654
timestamp 1649977179
transform 1 0 22032 0 1 29653
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1655
timestamp 1649977179
transform 1 0 18632 0 1 26389
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1656
timestamp 1649977179
transform 1 0 20808 0 1 30197
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1657
timestamp 1649977179
transform 1 0 20672 0 1 26797
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1658
timestamp 1649977179
transform 1 0 20672 0 1 27205
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1659
timestamp 1649977179
transform 1 0 20808 0 1 30469
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1660
timestamp 1649977179
transform 1 0 18632 0 1 27205
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1661
timestamp 1649977179
transform 1 0 18632 0 1 26661
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1662
timestamp 1649977179
transform 1 0 19040 0 1 27205
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1663
timestamp 1649977179
transform 1 0 19040 0 1 26661
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1664
timestamp 1649977179
transform 1 0 22168 0 1 28429
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1665
timestamp 1649977179
transform 1 0 21488 0 1 27205
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1666
timestamp 1649977179
transform 1 0 21488 0 1 26933
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1667
timestamp 1649977179
transform 1 0 21352 0 1 27205
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1668
timestamp 1649977179
transform 1 0 21352 0 1 26933
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1669
timestamp 1649977179
transform 1 0 22168 0 1 28157
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1670
timestamp 1649977179
transform 1 0 21216 0 1 28565
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1671
timestamp 1649977179
transform 1 0 21216 0 1 28837
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1672
timestamp 1649977179
transform 1 0 22032 0 1 27341
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1673
timestamp 1649977179
transform 1 0 22032 0 1 27613
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1674
timestamp 1649977179
transform 1 0 22032 0 1 28021
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1675
timestamp 1649977179
transform 1 0 22032 0 1 27749
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1676
timestamp 1649977179
transform 1 0 27472 0 1 30333
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1677
timestamp 1649977179
transform 1 0 27472 0 1 30605
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1678
timestamp 1649977179
transform 1 0 27472 0 1 26253
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1679
timestamp 1649977179
transform 1 0 27336 0 1 30741
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1680
timestamp 1649977179
transform 1 0 27336 0 1 31013
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1681
timestamp 1649977179
transform 1 0 27336 0 1 26389
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1682
timestamp 1649977179
transform 1 0 27336 0 1 26661
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1683
timestamp 1649977179
transform 1 0 22576 0 1 26117
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1684
timestamp 1649977179
transform 1 0 20808 0 1 26117
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1685
timestamp 1649977179
transform 1 0 22168 0 1 26117
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1686
timestamp 1649977179
transform 1 0 15912 0 1 25029
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1687
timestamp 1649977179
transform 1 0 2531 0 1 25300
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1688
timestamp 1649977179
transform 1 0 1224 0 1 23941
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1689
timestamp 1649977179
transform 1 0 2312 0 1 24485
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1690
timestamp 1649977179
transform 1 0 2312 0 1 23941
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1691
timestamp 1649977179
transform 1 0 544 0 1 23125
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1692
timestamp 1649977179
transform 1 0 3808 0 1 25845
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1693
timestamp 1649977179
transform 1 0 3808 0 1 23261
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1694
timestamp 1649977179
transform 1 0 3808 0 1 23125
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1695
timestamp 1649977179
transform 1 0 1224 0 1 25573
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1696
timestamp 1649977179
transform 1 0 1224 0 1 22309
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1697
timestamp 1649977179
transform 1 0 3128 0 1 21765
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1698
timestamp 1649977179
transform 1 0 3128 0 1 22173
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1699
timestamp 1649977179
transform 1 0 1224 0 1 27205
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1700
timestamp 1649977179
transform 1 0 1224 0 1 28973
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1701
timestamp 1649977179
transform 1 0 1224 0 1 30469
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1702
timestamp 1649977179
transform 1 0 14008 0 1 30605
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1703
timestamp 1649977179
transform 1 0 15912 0 1 27613
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1704
timestamp 1649977179
transform 1 0 14008 0 1 30469
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1705
timestamp 1649977179
transform 1 0 14008 0 1 27749
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1706
timestamp 1649977179
transform 1 0 14144 0 1 29245
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1707
timestamp 1649977179
transform 1 0 14280 0 1 36181
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1708
timestamp 1649977179
transform 1 0 14280 0 1 33461
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1709
timestamp 1649977179
transform 1 0 14144 0 1 33325
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1710
timestamp 1649977179
transform 1 0 14144 0 1 34821
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1711
timestamp 1649977179
transform 1 0 14008 0 1 32101
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1712
timestamp 1649977179
transform 1 0 14144 0 1 31829
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1713
timestamp 1649977179
transform 1 0 14008 0 1 34685
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1714
timestamp 1649977179
transform 1 0 1224 0 1 35637
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1715
timestamp 1649977179
transform 1 0 1224 0 1 32373
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1716
timestamp 1649977179
transform 1 0 1224 0 1 34005
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1717
timestamp 1649977179
transform 1 0 1224 0 1 37269
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1718
timestamp 1649977179
transform 1 0 1224 0 1 40805
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1719
timestamp 1649977179
transform 1 0 1224 0 1 39037
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1720
timestamp 1649977179
transform 1 0 14144 0 1 37541
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1721
timestamp 1649977179
transform 1 0 27472 0 1 35229
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1722
timestamp 1649977179
transform 1 0 27472 0 1 34957
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1723
timestamp 1649977179
transform 1 0 22032 0 1 36317
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1724
timestamp 1649977179
transform 1 0 22168 0 1 35909
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1725
timestamp 1649977179
transform 1 0 22440 0 1 32101
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1726
timestamp 1649977179
transform 1 0 22440 0 1 32373
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1727
timestamp 1649977179
transform 1 0 22440 0 1 35637
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1728
timestamp 1649977179
transform 1 0 22440 0 1 35909
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1729
timestamp 1649977179
transform 1 0 22576 0 1 32509
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1730
timestamp 1649977179
transform 1 0 22576 0 1 32781
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1731
timestamp 1649977179
transform 1 0 22168 0 1 35637
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1732
timestamp 1649977179
transform 1 0 20944 0 1 36317
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1733
timestamp 1649977179
transform 1 0 20808 0 1 32917
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1734
timestamp 1649977179
transform 1 0 20808 0 1 33189
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1735
timestamp 1649977179
transform 1 0 20808 0 1 34549
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1736
timestamp 1649977179
transform 1 0 20808 0 1 34821
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1737
timestamp 1649977179
transform 1 0 20944 0 1 35229
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1738
timestamp 1649977179
transform 1 0 20944 0 1 34957
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1739
timestamp 1649977179
transform 1 0 22576 0 1 31965
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1740
timestamp 1649977179
transform 1 0 22576 0 1 31693
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1741
timestamp 1649977179
transform 1 0 20944 0 1 31693
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1742
timestamp 1649977179
transform 1 0 22440 0 1 31557
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1743
timestamp 1649977179
transform 1 0 22440 0 1 32917
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1744
timestamp 1649977179
transform 1 0 22440 0 1 33189
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1745
timestamp 1649977179
transform 1 0 21216 0 1 32509
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1746
timestamp 1649977179
transform 1 0 21216 0 1 32781
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1747
timestamp 1649977179
transform 1 0 20808 0 1 33597
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1748
timestamp 1649977179
transform 1 0 20944 0 1 31421
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1749
timestamp 1649977179
transform 1 0 22440 0 1 36045
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1750
timestamp 1649977179
transform 1 0 22440 0 1 36317
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1751
timestamp 1649977179
transform 1 0 22032 0 1 33189
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1752
timestamp 1649977179
transform 1 0 22032 0 1 32917
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1753
timestamp 1649977179
transform 1 0 22440 0 1 34413
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1754
timestamp 1649977179
transform 1 0 22440 0 1 34141
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1755
timestamp 1649977179
transform 1 0 22032 0 1 32509
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1756
timestamp 1649977179
transform 1 0 22032 0 1 32781
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1757
timestamp 1649977179
transform 1 0 22168 0 1 33325
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1758
timestamp 1649977179
transform 1 0 22168 0 1 33597
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1759
timestamp 1649977179
transform 1 0 22440 0 1 33325
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1760
timestamp 1649977179
transform 1 0 22440 0 1 33597
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1761
timestamp 1649977179
transform 1 0 22440 0 1 34005
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1762
timestamp 1649977179
transform 1 0 22440 0 1 33733
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1763
timestamp 1649977179
transform 1 0 21624 0 1 33189
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1764
timestamp 1649977179
transform 1 0 21624 0 1 32917
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1765
timestamp 1649977179
transform 1 0 20808 0 1 33325
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1766
timestamp 1649977179
transform 1 0 20808 0 1 35637
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1767
timestamp 1649977179
transform 1 0 21896 0 1 34821
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1768
timestamp 1649977179
transform 1 0 21896 0 1 35229
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1769
timestamp 1649977179
transform 1 0 20808 0 1 34413
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1770
timestamp 1649977179
transform 1 0 22168 0 1 31557
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1771
timestamp 1649977179
transform 1 0 20808 0 1 35365
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1772
timestamp 1649977179
transform 1 0 20944 0 1 32781
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1773
timestamp 1649977179
transform 1 0 20808 0 1 34141
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1774
timestamp 1649977179
transform 1 0 20944 0 1 32509
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1775
timestamp 1649977179
transform 1 0 21624 0 1 31693
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1776
timestamp 1649977179
transform 1 0 21624 0 1 31965
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1777
timestamp 1649977179
transform 1 0 21760 0 1 33325
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1778
timestamp 1649977179
transform 1 0 21760 0 1 33597
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1779
timestamp 1649977179
transform 1 0 21624 0 1 36317
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1780
timestamp 1649977179
transform 1 0 21624 0 1 36045
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1781
timestamp 1649977179
transform 1 0 21760 0 1 32101
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1782
timestamp 1649977179
transform 1 0 21760 0 1 32373
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1783
timestamp 1649977179
transform 1 0 20944 0 1 32101
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1784
timestamp 1649977179
transform 1 0 22032 0 1 33733
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1785
timestamp 1649977179
transform 1 0 22032 0 1 34005
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1786
timestamp 1649977179
transform 1 0 22032 0 1 34413
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1787
timestamp 1649977179
transform 1 0 21488 0 1 36045
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1788
timestamp 1649977179
transform 1 0 21488 0 1 36317
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1789
timestamp 1649977179
transform 1 0 22032 0 1 34141
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1790
timestamp 1649977179
transform 1 0 22032 0 1 32373
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1791
timestamp 1649977179
transform 1 0 21216 0 1 31693
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1792
timestamp 1649977179
transform 1 0 21216 0 1 31965
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1793
timestamp 1649977179
transform 1 0 21624 0 1 35501
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1794
timestamp 1649977179
transform 1 0 21352 0 1 35501
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1795
timestamp 1649977179
transform 1 0 22032 0 1 32101
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1796
timestamp 1649977179
transform 1 0 22032 0 1 31693
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1797
timestamp 1649977179
transform 1 0 21488 0 1 35637
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1798
timestamp 1649977179
transform 1 0 21488 0 1 35909
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1799
timestamp 1649977179
transform 1 0 21216 0 1 34413
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1800
timestamp 1649977179
transform 1 0 21216 0 1 34141
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1801
timestamp 1649977179
transform 1 0 21352 0 1 33325
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1802
timestamp 1649977179
transform 1 0 21352 0 1 33597
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1803
timestamp 1649977179
transform 1 0 21352 0 1 34005
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1804
timestamp 1649977179
transform 1 0 21352 0 1 33733
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1805
timestamp 1649977179
transform 1 0 22032 0 1 31965
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1806
timestamp 1649977179
transform 1 0 20808 0 1 33733
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1807
timestamp 1649977179
transform 1 0 20808 0 1 34005
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1808
timestamp 1649977179
transform 1 0 20944 0 1 32373
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1809
timestamp 1649977179
transform 1 0 20944 0 1 36045
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1810
timestamp 1649977179
transform 1 0 22032 0 1 36045
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1811
timestamp 1649977179
transform 1 0 22576 0 1 39853
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1812
timestamp 1649977179
transform 1 0 22576 0 1 39581
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1813
timestamp 1649977179
transform 1 0 22440 0 1 40805
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1814
timestamp 1649977179
transform 1 0 22440 0 1 41077
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1815
timestamp 1649977179
transform 1 0 22576 0 1 36861
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1816
timestamp 1649977179
transform 1 0 22576 0 1 37133
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1817
timestamp 1649977179
transform 1 0 22576 0 1 37541
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1818
timestamp 1649977179
transform 1 0 22576 0 1 37269
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1819
timestamp 1649977179
transform 1 0 22576 0 1 41213
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1820
timestamp 1649977179
transform 1 0 22576 0 1 41485
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1821
timestamp 1649977179
transform 1 0 22440 0 1 38357
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1822
timestamp 1649977179
transform 1 0 22440 0 1 38085
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1823
timestamp 1649977179
transform 1 0 22440 0 1 37677
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1824
timestamp 1649977179
transform 1 0 22440 0 1 37949
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1825
timestamp 1649977179
transform 1 0 22440 0 1 36725
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1826
timestamp 1649977179
transform 1 0 20808 0 1 39581
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1827
timestamp 1649977179
transform 1 0 22440 0 1 39989
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1828
timestamp 1649977179
transform 1 0 22440 0 1 40261
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1829
timestamp 1649977179
transform 1 0 22576 0 1 40669
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1830
timestamp 1649977179
transform 1 0 22576 0 1 40397
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1831
timestamp 1649977179
transform 1 0 21760 0 1 37677
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1832
timestamp 1649977179
transform 1 0 21760 0 1 37949
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1833
timestamp 1649977179
transform 1 0 20808 0 1 38085
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1834
timestamp 1649977179
transform 1 0 21760 0 1 36725
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1835
timestamp 1649977179
transform 1 0 21624 0 1 37541
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1836
timestamp 1649977179
transform 1 0 21624 0 1 37269
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1837
timestamp 1649977179
transform 1 0 21624 0 1 40669
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1838
timestamp 1649977179
transform 1 0 21624 0 1 40397
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1839
timestamp 1649977179
transform 1 0 21760 0 1 39581
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1840
timestamp 1649977179
transform 1 0 21760 0 1 39853
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1841
timestamp 1649977179
transform 1 0 21760 0 1 40805
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1842
timestamp 1649977179
transform 1 0 21760 0 1 41077
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1843
timestamp 1649977179
transform 1 0 21216 0 1 40397
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1844
timestamp 1649977179
transform 1 0 21216 0 1 40669
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1845
timestamp 1649977179
transform 1 0 21352 0 1 41485
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1846
timestamp 1649977179
transform 1 0 21352 0 1 41213
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1847
timestamp 1649977179
transform 1 0 21352 0 1 38357
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1848
timestamp 1649977179
transform 1 0 21352 0 1 38085
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1849
timestamp 1649977179
transform 1 0 20808 0 1 38357
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1850
timestamp 1649977179
transform 1 0 20808 0 1 38765
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1851
timestamp 1649977179
transform 1 0 20808 0 1 38493
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1852
timestamp 1649977179
transform 1 0 20808 0 1 40805
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1853
timestamp 1649977179
transform 1 0 20808 0 1 41077
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1854
timestamp 1649977179
transform 1 0 20808 0 1 41485
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1855
timestamp 1649977179
transform 1 0 21216 0 1 37269
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1856
timestamp 1649977179
transform 1 0 21216 0 1 37541
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1857
timestamp 1649977179
transform 1 0 21488 0 1 39173
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1858
timestamp 1649977179
transform 1 0 21488 0 1 38901
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1859
timestamp 1649977179
transform 1 0 21488 0 1 37133
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1860
timestamp 1649977179
transform 1 0 21488 0 1 36861
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1861
timestamp 1649977179
transform 1 0 21352 0 1 37133
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1862
timestamp 1649977179
transform 1 0 21352 0 1 36861
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1863
timestamp 1649977179
transform 1 0 22032 0 1 41213
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1864
timestamp 1649977179
transform 1 0 22032 0 1 41485
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1865
timestamp 1649977179
transform 1 0 22168 0 1 37133
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1866
timestamp 1649977179
transform 1 0 22168 0 1 36861
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1867
timestamp 1649977179
transform 1 0 22168 0 1 39989
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1868
timestamp 1649977179
transform 1 0 22168 0 1 40261
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1869
timestamp 1649977179
transform 1 0 22032 0 1 39853
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1870
timestamp 1649977179
transform 1 0 22032 0 1 39581
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1871
timestamp 1649977179
transform 1 0 22032 0 1 36725
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1872
timestamp 1649977179
transform 1 0 20808 0 1 41213
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1873
timestamp 1649977179
transform 1 0 22032 0 1 38085
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1874
timestamp 1649977179
transform 1 0 22032 0 1 38357
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1875
timestamp 1649977179
transform 1 0 22168 0 1 37949
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1876
timestamp 1649977179
transform 1 0 22168 0 1 37677
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1877
timestamp 1649977179
transform 1 0 22032 0 1 37269
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1878
timestamp 1649977179
transform 1 0 22032 0 1 37541
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1879
timestamp 1649977179
transform 1 0 22032 0 1 41077
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1880
timestamp 1649977179
transform 1 0 22032 0 1 40805
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1881
timestamp 1649977179
transform 1 0 22032 0 1 40397
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1882
timestamp 1649977179
transform 1 0 22032 0 1 40669
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1883
timestamp 1649977179
transform 1 0 20944 0 1 37949
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1884
timestamp 1649977179
transform 1 0 20944 0 1 37677
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1885
timestamp 1649977179
transform 1 0 20808 0 1 37269
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1886
timestamp 1649977179
transform 1 0 20808 0 1 37541
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1887
timestamp 1649977179
transform 1 0 20808 0 1 38901
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1888
timestamp 1649977179
transform 1 0 20808 0 1 39173
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1889
timestamp 1649977179
transform 1 0 20808 0 1 37133
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1890
timestamp 1649977179
transform 1 0 20808 0 1 36861
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1891
timestamp 1649977179
transform 1 0 20808 0 1 39309
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1892
timestamp 1649977179
transform 1 0 27336 0 1 38085
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1893
timestamp 1649977179
transform 1 0 27336 0 1 37813
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1894
timestamp 1649977179
transform 1 0 27472 0 1 39309
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1895
timestamp 1649977179
transform 1 0 27472 0 1 39037
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1896
timestamp 1649977179
transform 1 0 27472 0 1 40261
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1897
timestamp 1649977179
transform 1 0 27472 0 1 40533
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1898
timestamp 1649977179
transform 1 0 22440 0 1 36453
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1899
timestamp 1649977179
transform 1 0 21760 0 1 36453
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1900
timestamp 1649977179
transform 1 0 22032 0 1 36453
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1901
timestamp 1649977179
transform 1 0 22440 0 1 31285
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1902
timestamp 1649977179
transform 1 0 22168 0 1 31285
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1903
timestamp 1649977179
transform 1 0 22440 0 1 20949
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1904
timestamp 1649977179
transform 1 0 21760 0 1 20949
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1905
timestamp 1649977179
transform 1 0 22032 0 1 20949
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1906
timestamp 1649977179
transform 1 0 21352 0 1 20949
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1907
timestamp 1649977179
transform 1 0 19176 0 1 20949
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1908
timestamp 1649977179
transform 1 0 18360 0 1 20949
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1909
timestamp 1649977179
transform 1 0 20808 0 1 20949
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1910
timestamp 1649977179
transform 1 0 18632 0 1 20949
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1911
timestamp 1649977179
transform 1 0 17816 0 1 20949
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1912
timestamp 1649977179
transform 1 0 27608 0 1 43253
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1913
timestamp 1649977179
transform 1 0 27472 0 1 43661
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1914
timestamp 1649977179
transform 1 0 25840 0 1 45429
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1915
timestamp 1649977179
transform 1 0 25840 0 1 45157
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1916
timestamp 1649977179
transform 1 0 27336 0 1 46517
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1917
timestamp 1649977179
transform 1 0 27472 0 1 43389
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1918
timestamp 1649977179
transform 1 0 27608 0 1 42981
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1919
timestamp 1649977179
transform 1 0 22032 0 1 45429
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1920
timestamp 1649977179
transform 1 0 22168 0 1 42437
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1921
timestamp 1649977179
transform 1 0 22032 0 1 45157
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1922
timestamp 1649977179
transform 1 0 22168 0 1 44613
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1923
timestamp 1649977179
transform 1 0 21352 0 1 44613
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1924
timestamp 1649977179
transform 1 0 21216 0 1 41893
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1925
timestamp 1649977179
transform 1 0 21760 0 1 45429
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1926
timestamp 1649977179
transform 1 0 21760 0 1 45157
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1927
timestamp 1649977179
transform 1 0 20944 0 1 45021
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1928
timestamp 1649977179
transform 1 0 20944 0 1 44749
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1929
timestamp 1649977179
transform 1 0 21624 0 1 41893
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1930
timestamp 1649977179
transform 1 0 22168 0 1 42029
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1931
timestamp 1649977179
transform 1 0 21760 0 1 43797
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1932
timestamp 1649977179
transform 1 0 21760 0 1 43525
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1933
timestamp 1649977179
transform 1 0 22576 0 1 46653
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1934
timestamp 1649977179
transform 1 0 22576 0 1 46381
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1935
timestamp 1649977179
transform 1 0 22440 0 1 43525
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1936
timestamp 1649977179
transform 1 0 22440 0 1 43797
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1937
timestamp 1649977179
transform 1 0 21216 0 1 43117
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1938
timestamp 1649977179
transform 1 0 22032 0 1 43525
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1939
timestamp 1649977179
transform 1 0 22032 0 1 43797
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1940
timestamp 1649977179
transform 1 0 21216 0 1 45973
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1941
timestamp 1649977179
transform 1 0 20808 0 1 46381
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1942
timestamp 1649977179
transform 1 0 20808 0 1 46653
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1943
timestamp 1649977179
transform 1 0 21216 0 1 46245
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1944
timestamp 1649977179
transform 1 0 22440 0 1 45157
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1945
timestamp 1649977179
transform 1 0 22440 0 1 45429
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1946
timestamp 1649977179
transform 1 0 22440 0 1 45837
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1947
timestamp 1649977179
transform 1 0 22440 0 1 45565
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1948
timestamp 1649977179
transform 1 0 21216 0 1 42845
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1949
timestamp 1649977179
transform 1 0 22576 0 1 43933
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1950
timestamp 1649977179
transform 1 0 22576 0 1 44205
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1951
timestamp 1649977179
transform 1 0 21624 0 1 43389
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1952
timestamp 1649977179
transform 1 0 21488 0 1 43117
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1953
timestamp 1649977179
transform 1 0 22576 0 1 42301
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1954
timestamp 1649977179
transform 1 0 22576 0 1 42029
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1955
timestamp 1649977179
transform 1 0 22576 0 1 46245
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1956
timestamp 1649977179
transform 1 0 22440 0 1 41893
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1957
timestamp 1649977179
transform 1 0 22576 0 1 45973
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1958
timestamp 1649977179
transform 1 0 20808 0 1 43253
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1959
timestamp 1649977179
transform 1 0 20808 0 1 43525
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1960
timestamp 1649977179
transform 1 0 22168 0 1 46381
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1961
timestamp 1649977179
transform 1 0 21488 0 1 45021
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1962
timestamp 1649977179
transform 1 0 21216 0 1 45021
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1963
timestamp 1649977179
transform 1 0 21216 0 1 44749
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1964
timestamp 1649977179
transform 1 0 22168 0 1 42301
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1965
timestamp 1649977179
transform 1 0 21488 0 1 44749
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1966
timestamp 1649977179
transform 1 0 23256 0 1 45021
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1967
timestamp 1649977179
transform 1 0 23256 0 1 44749
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1968
timestamp 1649977179
transform 1 0 22440 0 1 42709
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1969
timestamp 1649977179
transform 1 0 22440 0 1 42437
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1970
timestamp 1649977179
transform 1 0 22576 0 1 45021
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1971
timestamp 1649977179
transform 1 0 22576 0 1 44749
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1972
timestamp 1649977179
transform 1 0 22440 0 1 44341
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1973
timestamp 1649977179
transform 1 0 21760 0 1 42029
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1974
timestamp 1649977179
transform 1 0 22168 0 1 46653
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1975
timestamp 1649977179
transform 1 0 22032 0 1 45021
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1976
timestamp 1649977179
transform 1 0 22440 0 1 44613
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1977
timestamp 1649977179
transform 1 0 21352 0 1 45837
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1978
timestamp 1649977179
transform 1 0 20808 0 1 45157
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1979
timestamp 1649977179
transform 1 0 20808 0 1 45429
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1980
timestamp 1649977179
transform 1 0 22032 0 1 44749
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1981
timestamp 1649977179
transform 1 0 21760 0 1 42301
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1982
timestamp 1649977179
transform 1 0 21352 0 1 45565
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1983
timestamp 1649977179
transform 1 0 22032 0 1 46245
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1984
timestamp 1649977179
transform 1 0 22168 0 1 44341
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1985
timestamp 1649977179
transform 1 0 22168 0 1 42709
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1986
timestamp 1649977179
transform 1 0 21352 0 1 44341
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1987
timestamp 1649977179
transform 1 0 22168 0 1 43933
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1988
timestamp 1649977179
transform 1 0 22168 0 1 44205
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1989
timestamp 1649977179
transform 1 0 22032 0 1 41893
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1990
timestamp 1649977179
transform 1 0 22032 0 1 45973
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1991
timestamp 1649977179
transform 1 0 22032 0 1 45565
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1992
timestamp 1649977179
transform 1 0 20944 0 1 46245
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1993
timestamp 1649977179
transform 1 0 20944 0 1 45973
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1994
timestamp 1649977179
transform 1 0 20944 0 1 45565
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1995
timestamp 1649977179
transform 1 0 20944 0 1 45837
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1996
timestamp 1649977179
transform 1 0 20808 0 1 43117
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1997
timestamp 1649977179
transform 1 0 20808 0 1 42845
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1998
timestamp 1649977179
transform 1 0 20808 0 1 42437
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1999
timestamp 1649977179
transform 1 0 20808 0 1 42709
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2000
timestamp 1649977179
transform 1 0 20944 0 1 42301
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2001
timestamp 1649977179
transform 1 0 20944 0 1 42029
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2002
timestamp 1649977179
transform 1 0 22032 0 1 45837
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2003
timestamp 1649977179
transform 1 0 20808 0 1 41893
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2004
timestamp 1649977179
transform 1 0 22168 0 1 51005
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2005
timestamp 1649977179
transform 1 0 21896 0 1 51005
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2006
timestamp 1649977179
transform 1 0 21896 0 1 50733
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2007
timestamp 1649977179
transform 1 0 21896 0 1 50325
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2008
timestamp 1649977179
transform 1 0 21896 0 1 50597
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2009
timestamp 1649977179
transform 1 0 20808 0 1 50325
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2010
timestamp 1649977179
transform 1 0 20808 0 1 50597
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2011
timestamp 1649977179
transform 1 0 20808 0 1 49781
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2012
timestamp 1649977179
transform 1 0 20808 0 1 49509
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2013
timestamp 1649977179
transform 1 0 20808 0 1 50733
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2014
timestamp 1649977179
transform 1 0 20808 0 1 51005
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2015
timestamp 1649977179
transform 1 0 21488 0 1 48965
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2016
timestamp 1649977179
transform 1 0 21488 0 1 48693
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2017
timestamp 1649977179
transform 1 0 21488 0 1 47469
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2018
timestamp 1649977179
transform 1 0 21488 0 1 47741
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2019
timestamp 1649977179
transform 1 0 21352 0 1 48965
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2020
timestamp 1649977179
transform 1 0 21352 0 1 48693
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2021
timestamp 1649977179
transform 1 0 20808 0 1 48693
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2022
timestamp 1649977179
transform 1 0 20808 0 1 48965
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2023
timestamp 1649977179
transform 1 0 20944 0 1 49373
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2024
timestamp 1649977179
transform 1 0 20944 0 1 49101
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2025
timestamp 1649977179
transform 1 0 20808 0 1 51141
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2026
timestamp 1649977179
transform 1 0 20808 0 1 51413
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2027
timestamp 1649977179
transform 1 0 21352 0 1 50733
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2028
timestamp 1649977179
transform 1 0 21352 0 1 51005
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2029
timestamp 1649977179
transform 1 0 21760 0 1 51413
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2030
timestamp 1649977179
transform 1 0 21488 0 1 50189
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2031
timestamp 1649977179
transform 1 0 21488 0 1 49917
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2032
timestamp 1649977179
transform 1 0 22168 0 1 49509
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2033
timestamp 1649977179
transform 1 0 22576 0 1 51821
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2034
timestamp 1649977179
transform 1 0 22576 0 1 48965
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2035
timestamp 1649977179
transform 1 0 22576 0 1 48693
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2036
timestamp 1649977179
transform 1 0 20808 0 1 48013
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2037
timestamp 1649977179
transform 1 0 20808 0 1 48285
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2038
timestamp 1649977179
transform 1 0 20808 0 1 47469
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2039
timestamp 1649977179
transform 1 0 20808 0 1 47197
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2040
timestamp 1649977179
transform 1 0 21216 0 1 49917
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2041
timestamp 1649977179
transform 1 0 20944 0 1 47061
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2042
timestamp 1649977179
transform 1 0 22576 0 1 49917
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2043
timestamp 1649977179
transform 1 0 22576 0 1 50189
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2044
timestamp 1649977179
transform 1 0 22168 0 1 49781
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2045
timestamp 1649977179
transform 1 0 20944 0 1 49917
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2046
timestamp 1649977179
transform 1 0 21216 0 1 50189
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2047
timestamp 1649977179
transform 1 0 21760 0 1 49509
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2048
timestamp 1649977179
transform 1 0 20944 0 1 50189
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2049
timestamp 1649977179
transform 1 0 22168 0 1 50189
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2050
timestamp 1649977179
transform 1 0 22168 0 1 48965
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2051
timestamp 1649977179
transform 1 0 22168 0 1 48693
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2052
timestamp 1649977179
transform 1 0 22168 0 1 48285
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2053
timestamp 1649977179
transform 1 0 22440 0 1 49101
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2054
timestamp 1649977179
transform 1 0 22440 0 1 49373
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2055
timestamp 1649977179
transform 1 0 22440 0 1 49781
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2056
timestamp 1649977179
transform 1 0 22440 0 1 49509
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2057
timestamp 1649977179
transform 1 0 22168 0 1 48557
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2058
timestamp 1649977179
transform 1 0 22168 0 1 49917
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2059
timestamp 1649977179
transform 1 0 22032 0 1 50597
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2060
timestamp 1649977179
transform 1 0 22032 0 1 50325
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2061
timestamp 1649977179
transform 1 0 22168 0 1 51821
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2062
timestamp 1649977179
transform 1 0 22168 0 1 48149
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2063
timestamp 1649977179
transform 1 0 22168 0 1 47877
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2064
timestamp 1649977179
transform 1 0 22032 0 1 49101
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2065
timestamp 1649977179
transform 1 0 22032 0 1 49373
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2066
timestamp 1649977179
transform 1 0 21760 0 1 49781
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2067
timestamp 1649977179
transform 1 0 21624 0 1 49373
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2068
timestamp 1649977179
transform 1 0 22440 0 1 48557
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2069
timestamp 1649977179
transform 1 0 21216 0 1 49101
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2070
timestamp 1649977179
transform 1 0 22440 0 1 48285
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2071
timestamp 1649977179
transform 1 0 21352 0 1 47061
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2072
timestamp 1649977179
transform 1 0 21216 0 1 49373
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2073
timestamp 1649977179
transform 1 0 21624 0 1 49101
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2074
timestamp 1649977179
transform 1 0 21760 0 1 48285
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2075
timestamp 1649977179
transform 1 0 21760 0 1 48557
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2076
timestamp 1649977179
transform 1 0 22576 0 1 51005
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2077
timestamp 1649977179
transform 1 0 22576 0 1 50733
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2078
timestamp 1649977179
transform 1 0 22440 0 1 50325
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2079
timestamp 1649977179
transform 1 0 22440 0 1 50597
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2080
timestamp 1649977179
transform 1 0 22168 0 1 50733
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2081
timestamp 1649977179
transform 1 0 21760 0 1 47061
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2082
timestamp 1649977179
transform 1 0 22440 0 1 48149
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2083
timestamp 1649977179
transform 1 0 22440 0 1 47877
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2084
timestamp 1649977179
transform 1 0 21760 0 1 51685
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2085
timestamp 1649977179
transform 1 0 27336 0 1 47197
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2086
timestamp 1649977179
transform 1 0 27336 0 1 46925
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2087
timestamp 1649977179
transform 1 0 27336 0 1 51005
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2088
timestamp 1649977179
transform 1 0 27336 0 1 51277
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2089
timestamp 1649977179
transform 1 0 27336 0 1 46789
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2090
timestamp 1649977179
transform 1 0 20944 0 1 46789
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2091
timestamp 1649977179
transform 1 0 21352 0 1 46789
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2092
timestamp 1649977179
transform 1 0 21760 0 1 46789
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2093
timestamp 1649977179
transform 1 0 1224 0 1 42437
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2094
timestamp 1649977179
transform 1 0 1224 0 1 44069
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2095
timestamp 1649977179
transform 1 0 1224 0 1 45565
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2096
timestamp 1649977179
transform 1 0 1224 0 1 50869
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2097
timestamp 1649977179
transform 1 0 1224 0 1 47469
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2098
timestamp 1649977179
transform 1 0 1224 0 1 48965
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2099
timestamp 1649977179
transform 1 0 1224 0 1 54133
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2100
timestamp 1649977179
transform 1 0 1224 0 1 55901
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2101
timestamp 1649977179
transform 1 0 1224 0 1 52501
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2102
timestamp 1649977179
transform 1 0 1224 0 1 59165
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2103
timestamp 1649977179
transform 1 0 1224 0 1 60933
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2104
timestamp 1649977179
transform 1 0 1224 0 1 57533
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2105
timestamp 1649977179
transform 1 0 27472 0 1 55901
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2106
timestamp 1649977179
transform 1 0 27608 0 1 55221
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2107
timestamp 1649977179
transform 1 0 27608 0 1 55493
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2108
timestamp 1649977179
transform 1 0 27472 0 1 52093
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2109
timestamp 1649977179
transform 1 0 27472 0 1 52365
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2110
timestamp 1649977179
transform 1 0 27472 0 1 55493
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2111
timestamp 1649977179
transform 1 0 21216 0 1 52637
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2112
timestamp 1649977179
transform 1 0 21488 0 1 54541
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2113
timestamp 1649977179
transform 1 0 21488 0 1 54269
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2114
timestamp 1649977179
transform 1 0 21352 0 1 54541
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2115
timestamp 1649977179
transform 1 0 22168 0 1 54133
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2116
timestamp 1649977179
transform 1 0 20808 0 1 55493
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2117
timestamp 1649977179
transform 1 0 20808 0 1 53453
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2118
timestamp 1649977179
transform 1 0 20808 0 1 53725
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2119
timestamp 1649977179
transform 1 0 22032 0 1 53453
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2120
timestamp 1649977179
transform 1 0 22032 0 1 53725
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2121
timestamp 1649977179
transform 1 0 22440 0 1 53453
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2122
timestamp 1649977179
transform 1 0 20944 0 1 52637
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2123
timestamp 1649977179
transform 1 0 20944 0 1 52909
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2124
timestamp 1649977179
transform 1 0 22440 0 1 53725
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2125
timestamp 1649977179
transform 1 0 22440 0 1 54133
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2126
timestamp 1649977179
transform 1 0 22440 0 1 53861
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2127
timestamp 1649977179
transform 1 0 22032 0 1 56581
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2128
timestamp 1649977179
transform 1 0 22032 0 1 56853
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2129
timestamp 1649977179
transform 1 0 22440 0 1 56581
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2130
timestamp 1649977179
transform 1 0 22440 0 1 56853
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2131
timestamp 1649977179
transform 1 0 22168 0 1 53317
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2132
timestamp 1649977179
transform 1 0 20944 0 1 54541
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2133
timestamp 1649977179
transform 1 0 20944 0 1 54269
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2134
timestamp 1649977179
transform 1 0 20808 0 1 53861
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2135
timestamp 1649977179
transform 1 0 20808 0 1 54133
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2136
timestamp 1649977179
transform 1 0 20808 0 1 54677
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2137
timestamp 1649977179
transform 1 0 20808 0 1 54949
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2138
timestamp 1649977179
transform 1 0 20944 0 1 55357
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2139
timestamp 1649977179
transform 1 0 20944 0 1 55085
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2140
timestamp 1649977179
transform 1 0 21624 0 1 53725
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2141
timestamp 1649977179
transform 1 0 21624 0 1 53453
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2142
timestamp 1649977179
transform 1 0 22440 0 1 56989
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2143
timestamp 1649977179
transform 1 0 21352 0 1 54269
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2144
timestamp 1649977179
transform 1 0 22032 0 1 56989
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2145
timestamp 1649977179
transform 1 0 21760 0 1 52637
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2146
timestamp 1649977179
transform 1 0 21760 0 1 52909
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2147
timestamp 1649977179
transform 1 0 21760 0 1 53861
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2148
timestamp 1649977179
transform 1 0 21760 0 1 54133
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2149
timestamp 1649977179
transform 1 0 21488 0 1 53045
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2150
timestamp 1649977179
transform 1 0 21760 0 1 56989
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2151
timestamp 1649977179
transform 1 0 22168 0 1 53045
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2152
timestamp 1649977179
transform 1 0 21488 0 1 53317
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2153
timestamp 1649977179
transform 1 0 21352 0 1 53045
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2154
timestamp 1649977179
transform 1 0 22168 0 1 52637
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2155
timestamp 1649977179
transform 1 0 22168 0 1 52909
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2156
timestamp 1649977179
transform 1 0 21352 0 1 53317
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2157
timestamp 1649977179
transform 1 0 21624 0 1 54949
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2158
timestamp 1649977179
transform 1 0 21624 0 1 54677
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2159
timestamp 1649977179
transform 1 0 20808 0 1 52229
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2160
timestamp 1649977179
transform 1 0 22168 0 1 52501
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2161
timestamp 1649977179
transform 1 0 22168 0 1 52229
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2162
timestamp 1649977179
transform 1 0 22168 0 1 52093
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2163
timestamp 1649977179
transform 1 0 20808 0 1 55765
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2164
timestamp 1649977179
transform 1 0 22440 0 1 52229
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2165
timestamp 1649977179
transform 1 0 21624 0 1 56445
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2166
timestamp 1649977179
transform 1 0 21624 0 1 56173
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2167
timestamp 1649977179
transform 1 0 21488 0 1 55765
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2168
timestamp 1649977179
transform 1 0 21488 0 1 55493
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2169
timestamp 1649977179
transform 1 0 22440 0 1 52501
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2170
timestamp 1649977179
transform 1 0 22576 0 1 52909
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2171
timestamp 1649977179
transform 1 0 22576 0 1 52637
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2172
timestamp 1649977179
transform 1 0 22440 0 1 54677
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2173
timestamp 1649977179
transform 1 0 22440 0 1 54949
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2174
timestamp 1649977179
transform 1 0 20944 0 1 55901
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2175
timestamp 1649977179
transform 1 0 21216 0 1 56989
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2176
timestamp 1649977179
transform 1 0 21352 0 1 56445
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2177
timestamp 1649977179
transform 1 0 22576 0 1 52093
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2178
timestamp 1649977179
transform 1 0 22440 0 1 53045
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2179
timestamp 1649977179
transform 1 0 22440 0 1 53317
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2180
timestamp 1649977179
transform 1 0 21352 0 1 56173
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2181
timestamp 1649977179
transform 1 0 22440 0 1 56173
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2182
timestamp 1649977179
transform 1 0 22440 0 1 56445
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2183
timestamp 1649977179
transform 1 0 20944 0 1 56173
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2184
timestamp 1649977179
transform 1 0 22168 0 1 54541
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2185
timestamp 1649977179
transform 1 0 22168 0 1 54269
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2186
timestamp 1649977179
transform 1 0 22168 0 1 53861
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2187
timestamp 1649977179
transform 1 0 22576 0 1 54269
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2188
timestamp 1649977179
transform 1 0 22576 0 1 54541
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2189
timestamp 1649977179
transform 1 0 22032 0 1 54949
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2190
timestamp 1649977179
transform 1 0 22032 0 1 54677
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2191
timestamp 1649977179
transform 1 0 22168 0 1 56173
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2192
timestamp 1649977179
transform 1 0 22168 0 1 56445
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2193
timestamp 1649977179
transform 1 0 21216 0 1 52909
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2194
timestamp 1649977179
transform 1 0 20808 0 1 58893
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2195
timestamp 1649977179
transform 1 0 20808 0 1 58621
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2196
timestamp 1649977179
transform 1 0 20944 0 1 61341
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2197
timestamp 1649977179
transform 1 0 20944 0 1 61613
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2198
timestamp 1649977179
transform 1 0 20944 0 1 62021
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2199
timestamp 1649977179
transform 1 0 20944 0 1 61749
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2200
timestamp 1649977179
transform 1 0 20808 0 1 62157
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2201
timestamp 1649977179
transform 1 0 20808 0 1 59029
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2202
timestamp 1649977179
transform 1 0 20808 0 1 59301
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2203
timestamp 1649977179
transform 1 0 20944 0 1 58077
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2204
timestamp 1649977179
transform 1 0 20944 0 1 57805
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2205
timestamp 1649977179
transform 1 0 20808 0 1 57397
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2206
timestamp 1649977179
transform 1 0 20808 0 1 57669
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2207
timestamp 1649977179
transform 1 0 20808 0 1 60117
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2208
timestamp 1649977179
transform 1 0 20808 0 1 59845
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2209
timestamp 1649977179
transform 1 0 20808 0 1 59437
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2210
timestamp 1649977179
transform 1 0 20808 0 1 59709
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2211
timestamp 1649977179
transform 1 0 21216 0 1 58621
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2212
timestamp 1649977179
transform 1 0 21624 0 1 62157
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2213
timestamp 1649977179
transform 1 0 21216 0 1 58893
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2214
timestamp 1649977179
transform 1 0 21760 0 1 57261
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2215
timestamp 1649977179
transform 1 0 21896 0 1 60117
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2216
timestamp 1649977179
transform 1 0 21896 0 1 60389
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2217
timestamp 1649977179
transform 1 0 21760 0 1 59437
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2218
timestamp 1649977179
transform 1 0 21760 0 1 59709
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2219
timestamp 1649977179
transform 1 0 21760 0 1 58213
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2220
timestamp 1649977179
transform 1 0 21760 0 1 58485
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2221
timestamp 1649977179
transform 1 0 21760 0 1 61341
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2222
timestamp 1649977179
transform 1 0 21760 0 1 61613
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2223
timestamp 1649977179
transform 1 0 21352 0 1 62021
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2224
timestamp 1649977179
transform 1 0 21352 0 1 61749
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2225
timestamp 1649977179
transform 1 0 21352 0 1 58213
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2226
timestamp 1649977179
transform 1 0 21352 0 1 58485
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2227
timestamp 1649977179
transform 1 0 21352 0 1 61205
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2228
timestamp 1649977179
transform 1 0 21352 0 1 60933
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2229
timestamp 1649977179
transform 1 0 21216 0 1 62157
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2230
timestamp 1649977179
transform 1 0 22440 0 1 60117
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2231
timestamp 1649977179
transform 1 0 22440 0 1 60389
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2232
timestamp 1649977179
transform 1 0 22576 0 1 60797
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2233
timestamp 1649977179
transform 1 0 22576 0 1 60525
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2234
timestamp 1649977179
transform 1 0 22440 0 1 57805
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2235
timestamp 1649977179
transform 1 0 22440 0 1 58077
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2236
timestamp 1649977179
transform 1 0 21488 0 1 58077
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2237
timestamp 1649977179
transform 1 0 21488 0 1 57805
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2238
timestamp 1649977179
transform 1 0 22440 0 1 58893
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2239
timestamp 1649977179
transform 1 0 22440 0 1 58621
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2240
timestamp 1649977179
transform 1 0 22440 0 1 58213
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2241
timestamp 1649977179
transform 1 0 22440 0 1 58485
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2242
timestamp 1649977179
transform 1 0 22576 0 1 57669
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2243
timestamp 1649977179
transform 1 0 22576 0 1 57397
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2244
timestamp 1649977179
transform 1 0 22440 0 1 57261
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2245
timestamp 1649977179
transform 1 0 22576 0 1 62157
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2246
timestamp 1649977179
transform 1 0 22440 0 1 61749
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2247
timestamp 1649977179
transform 1 0 22440 0 1 62021
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2248
timestamp 1649977179
transform 1 0 22440 0 1 59029
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2249
timestamp 1649977179
transform 1 0 22440 0 1 59301
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2250
timestamp 1649977179
transform 1 0 22440 0 1 60933
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2251
timestamp 1649977179
transform 1 0 22440 0 1 61205
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2252
timestamp 1649977179
transform 1 0 22440 0 1 61613
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2253
timestamp 1649977179
transform 1 0 22440 0 1 61341
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2254
timestamp 1649977179
transform 1 0 21216 0 1 57261
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2255
timestamp 1649977179
transform 1 0 22032 0 1 59029
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2256
timestamp 1649977179
transform 1 0 22032 0 1 59301
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2257
timestamp 1649977179
transform 1 0 20808 0 1 58485
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2258
timestamp 1649977179
transform 1 0 20808 0 1 58213
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2259
timestamp 1649977179
transform 1 0 22032 0 1 61613
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2260
timestamp 1649977179
transform 1 0 22032 0 1 61341
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2261
timestamp 1649977179
transform 1 0 22032 0 1 57261
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2262
timestamp 1649977179
transform 1 0 22168 0 1 61749
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2263
timestamp 1649977179
transform 1 0 22168 0 1 62021
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2264
timestamp 1649977179
transform 1 0 22168 0 1 57397
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2265
timestamp 1649977179
transform 1 0 22168 0 1 57669
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2266
timestamp 1649977179
transform 1 0 22032 0 1 62157
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2267
timestamp 1649977179
transform 1 0 22032 0 1 57805
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2268
timestamp 1649977179
transform 1 0 22032 0 1 58077
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2269
timestamp 1649977179
transform 1 0 22032 0 1 60117
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2270
timestamp 1649977179
transform 1 0 22032 0 1 60389
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2271
timestamp 1649977179
transform 1 0 22168 0 1 58893
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2272
timestamp 1649977179
transform 1 0 22168 0 1 58621
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2273
timestamp 1649977179
transform 1 0 22168 0 1 58213
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2274
timestamp 1649977179
transform 1 0 22168 0 1 58485
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2275
timestamp 1649977179
transform 1 0 22168 0 1 61205
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2276
timestamp 1649977179
transform 1 0 22168 0 1 60933
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2277
timestamp 1649977179
transform 1 0 22168 0 1 60525
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2278
timestamp 1649977179
transform 1 0 22168 0 1 60797
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2279
timestamp 1649977179
transform 1 0 27608 0 1 58349
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2280
timestamp 1649977179
transform 1 0 27608 0 1 58621
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2281
timestamp 1649977179
transform 1 0 27336 0 1 59845
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2282
timestamp 1649977179
transform 1 0 27336 0 1 59573
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2283
timestamp 1649977179
transform 1 0 20808 0 1 51957
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2284
timestamp 1649977179
transform 1 0 27608 0 1 65013
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2285
timestamp 1649977179
transform 1 0 27608 0 1 63925
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2286
timestamp 1649977179
transform 1 0 27608 0 1 64197
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2287
timestamp 1649977179
transform 1 0 27336 0 1 64469
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2288
timestamp 1649977179
transform 1 0 27336 0 1 64197
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2289
timestamp 1649977179
transform 1 0 27472 0 1 63789
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2290
timestamp 1649977179
transform 1 0 27472 0 1 63517
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2291
timestamp 1649977179
transform 1 0 27608 0 1 64741
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2292
timestamp 1649977179
transform 1 0 21488 0 1 65557
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2293
timestamp 1649977179
transform 1 0 21488 0 1 65285
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2294
timestamp 1649977179
transform 1 0 21352 0 1 65557
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2295
timestamp 1649977179
transform 1 0 21352 0 1 65285
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2296
timestamp 1649977179
transform 1 0 20808 0 1 62837
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2297
timestamp 1649977179
transform 1 0 22440 0 1 64877
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2298
timestamp 1649977179
transform 1 0 22440 0 1 65149
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2299
timestamp 1649977179
transform 1 0 22440 0 1 65557
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2300
timestamp 1649977179
transform 1 0 22440 0 1 65285
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2301
timestamp 1649977179
transform 1 0 22032 0 1 67189
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2302
timestamp 1649977179
transform 1 0 22032 0 1 66917
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2303
timestamp 1649977179
transform 1 0 20808 0 1 65965
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2304
timestamp 1649977179
transform 1 0 20808 0 1 65693
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2305
timestamp 1649977179
transform 1 0 20944 0 1 65285
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2306
timestamp 1649977179
transform 1 0 20944 0 1 65557
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2307
timestamp 1649977179
transform 1 0 22168 0 1 64469
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2308
timestamp 1649977179
transform 1 0 22168 0 1 64741
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2309
timestamp 1649977179
transform 1 0 22440 0 1 66509
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2310
timestamp 1649977179
transform 1 0 22440 0 1 66781
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2311
timestamp 1649977179
transform 1 0 22168 0 1 65149
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2312
timestamp 1649977179
transform 1 0 22168 0 1 64877
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2313
timestamp 1649977179
transform 1 0 22168 0 1 66101
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2314
timestamp 1649977179
transform 1 0 22168 0 1 66373
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2315
timestamp 1649977179
transform 1 0 22440 0 1 67189
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2316
timestamp 1649977179
transform 1 0 22440 0 1 66917
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2317
timestamp 1649977179
transform 1 0 22032 0 1 66781
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2318
timestamp 1649977179
transform 1 0 22032 0 1 66509
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2319
timestamp 1649977179
transform 1 0 21624 0 1 62429
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2320
timestamp 1649977179
transform 1 0 22576 0 1 62973
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2321
timestamp 1649977179
transform 1 0 22576 0 1 63245
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2322
timestamp 1649977179
transform 1 0 22032 0 1 62973
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2323
timestamp 1649977179
transform 1 0 22032 0 1 63245
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2324
timestamp 1649977179
transform 1 0 22576 0 1 64741
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2325
timestamp 1649977179
transform 1 0 22576 0 1 64469
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2326
timestamp 1649977179
transform 1 0 22440 0 1 62837
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2327
timestamp 1649977179
transform 1 0 22440 0 1 62565
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2328
timestamp 1649977179
transform 1 0 22576 0 1 66373
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2329
timestamp 1649977179
transform 1 0 22576 0 1 66101
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2330
timestamp 1649977179
transform 1 0 22576 0 1 65693
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2331
timestamp 1649977179
transform 1 0 22032 0 1 64469
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2332
timestamp 1649977179
transform 1 0 22032 0 1 65013
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2333
timestamp 1649977179
transform 1 0 20808 0 1 63789
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2334
timestamp 1649977179
transform 1 0 20808 0 1 67325
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2335
timestamp 1649977179
transform 1 0 22576 0 1 65965
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2336
timestamp 1649977179
transform 1 0 20808 0 1 64061
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2337
timestamp 1649977179
transform 1 0 22576 0 1 62429
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2338
timestamp 1649977179
transform 1 0 20944 0 1 66373
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2339
timestamp 1649977179
transform 1 0 21760 0 1 62565
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2340
timestamp 1649977179
transform 1 0 22032 0 1 65965
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2341
timestamp 1649977179
transform 1 0 22032 0 1 65693
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2342
timestamp 1649977179
transform 1 0 22032 0 1 65285
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2343
timestamp 1649977179
transform 1 0 22032 0 1 65557
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2344
timestamp 1649977179
transform 1 0 22032 0 1 62837
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2345
timestamp 1649977179
transform 1 0 22032 0 1 62565
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2346
timestamp 1649977179
transform 1 0 21760 0 1 62837
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2347
timestamp 1649977179
transform 1 0 21896 0 1 64877
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2348
timestamp 1649977179
transform 1 0 21896 0 1 65149
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2349
timestamp 1649977179
transform 1 0 21624 0 1 66509
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2350
timestamp 1649977179
transform 1 0 21624 0 1 66781
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2351
timestamp 1649977179
transform 1 0 20944 0 1 66101
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2352
timestamp 1649977179
transform 1 0 20808 0 1 66509
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2353
timestamp 1649977179
transform 1 0 20808 0 1 66781
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2354
timestamp 1649977179
transform 1 0 20808 0 1 67189
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2355
timestamp 1649977179
transform 1 0 20808 0 1 66917
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2356
timestamp 1649977179
transform 1 0 21624 0 1 67325
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2357
timestamp 1649977179
transform 1 0 21760 0 1 64333
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2358
timestamp 1649977179
transform 1 0 21760 0 1 64061
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2359
timestamp 1649977179
transform 1 0 21896 0 1 63381
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2360
timestamp 1649977179
transform 1 0 21896 0 1 63653
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2361
timestamp 1649977179
transform 1 0 21760 0 1 65693
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2362
timestamp 1649977179
transform 1 0 21760 0 1 65965
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2363
timestamp 1649977179
transform 1 0 22032 0 1 62429
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2364
timestamp 1649977179
transform 1 0 20808 0 1 62429
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2365
timestamp 1649977179
transform 1 0 20808 0 1 63381
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2366
timestamp 1649977179
transform 1 0 20808 0 1 63653
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2367
timestamp 1649977179
transform 1 0 20808 0 1 63245
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2368
timestamp 1649977179
transform 1 0 21216 0 1 62429
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2369
timestamp 1649977179
transform 1 0 21488 0 1 66917
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2370
timestamp 1649977179
transform 1 0 21488 0 1 67189
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2371
timestamp 1649977179
transform 1 0 20808 0 1 62973
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2372
timestamp 1649977179
transform 1 0 21216 0 1 67325
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2373
timestamp 1649977179
transform 1 0 21488 0 1 66101
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2374
timestamp 1649977179
transform 1 0 21488 0 1 66373
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2375
timestamp 1649977179
transform 1 0 21352 0 1 66101
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2376
timestamp 1649977179
transform 1 0 21352 0 1 66373
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2377
timestamp 1649977179
transform 1 0 20808 0 1 62565
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2378
timestamp 1649977179
transform 1 0 21896 0 1 68277
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2379
timestamp 1649977179
transform 1 0 22440 0 1 68821
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2380
timestamp 1649977179
transform 1 0 22440 0 1 69093
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2381
timestamp 1649977179
transform 1 0 21896 0 1 68005
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2382
timestamp 1649977179
transform 1 0 21352 0 1 69229
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2383
timestamp 1649977179
transform 1 0 21352 0 1 69501
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2384
timestamp 1649977179
transform 1 0 21216 0 1 67597
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2385
timestamp 1649977179
transform 1 0 22032 0 1 68413
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2386
timestamp 1649977179
transform 1 0 22032 0 1 68685
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2387
timestamp 1649977179
transform 1 0 22440 0 1 69229
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2388
timestamp 1649977179
transform 1 0 22440 0 1 69501
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2389
timestamp 1649977179
transform 1 0 22440 0 1 69909
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2390
timestamp 1649977179
transform 1 0 22440 0 1 69637
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2391
timestamp 1649977179
transform 1 0 22168 0 1 69501
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2392
timestamp 1649977179
transform 1 0 22168 0 1 69229
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2393
timestamp 1649977179
transform 1 0 22032 0 1 68821
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2394
timestamp 1649977179
transform 1 0 22032 0 1 69093
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2395
timestamp 1649977179
transform 1 0 20808 0 1 67733
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2396
timestamp 1649977179
transform 1 0 20808 0 1 68005
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2397
timestamp 1649977179
transform 1 0 22440 0 1 68685
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2398
timestamp 1649977179
transform 1 0 22440 0 1 68413
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2399
timestamp 1649977179
transform 1 0 20808 0 1 67597
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2400
timestamp 1649977179
transform 1 0 20808 0 1 68549
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2401
timestamp 1649977179
transform 1 0 20808 0 1 68821
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2402
timestamp 1649977179
transform 1 0 20808 0 1 69229
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2403
timestamp 1649977179
transform 1 0 20808 0 1 69501
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2404
timestamp 1649977179
transform 1 0 22168 0 1 69909
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2405
timestamp 1649977179
transform 1 0 22168 0 1 69637
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2406
timestamp 1649977179
transform 1 0 21624 0 1 69501
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2407
timestamp 1649977179
transform 1 0 21624 0 1 69229
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2408
timestamp 1649977179
transform 1 0 21760 0 1 69093
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2409
timestamp 1649977179
transform 1 0 21760 0 1 68821
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2410
timestamp 1649977179
transform 1 0 21624 0 1 67597
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2411
timestamp 1649977179
transform 1 0 31280 0 1 71405
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2412
timestamp 1649977179
transform 1 0 29784 0 1 71405
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2413
timestamp 1649977179
transform 1 0 29784 0 1 70997
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2414
timestamp 1649977179
transform 1 0 28696 0 1 70997
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2415
timestamp 1649977179
transform 1 0 28696 0 1 71405
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2416
timestamp 1649977179
transform 1 0 28560 0 1 71405
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2417
timestamp 1649977179
transform 1 0 28560 0 1 70997
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2418
timestamp 1649977179
transform 1 0 33728 0 1 70997
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2419
timestamp 1649977179
transform 1 0 33728 0 1 71405
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2420
timestamp 1649977179
transform 1 0 32504 0 1 70997
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2421
timestamp 1649977179
transform 1 0 32504 0 1 71405
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2422
timestamp 1649977179
transform 1 0 31960 0 1 71405
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2423
timestamp 1649977179
transform 1 0 31960 0 1 70997
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2424
timestamp 1649977179
transform 1 0 27336 0 1 67597
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2425
timestamp 1649977179
transform 1 0 27336 0 1 67869
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2426
timestamp 1649977179
transform 1 0 27472 0 1 68141
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2427
timestamp 1649977179
transform 1 0 27472 0 1 67869
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2428
timestamp 1649977179
transform 1 0 28968 0 1 70725
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2429
timestamp 1649977179
transform 1 0 31280 0 1 70997
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2430
timestamp 1649977179
transform 1 0 1224 0 1 64061
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2431
timestamp 1649977179
transform 1 0 1224 0 1 62565
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2432
timestamp 1649977179
transform 1 0 1224 0 1 65965
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2433
timestamp 1649977179
transform 1 0 1224 0 1 70997
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2434
timestamp 1649977179
transform 1 0 1224 0 1 69229
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2435
timestamp 1649977179
transform 1 0 1224 0 1 67461
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2436
timestamp 1649977179
transform 1 0 1224 0 1 74125
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2437
timestamp 1649977179
transform 1 0 1224 0 1 76029
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2438
timestamp 1649977179
transform 1 0 1224 0 1 77525
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2439
timestamp 1649977179
transform 1 0 1224 0 1 79429
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2440
timestamp 1649977179
transform 1 0 3944 0 1 82013
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2441
timestamp 1649977179
transform 1 0 3944 0 1 81469
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2442
timestamp 1649977179
transform 1 0 2176 0 1 82013
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2443
timestamp 1649977179
transform 1 0 2176 0 1 81469
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2444
timestamp 1649977179
transform 1 0 2040 0 1 81333
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2445
timestamp 1649977179
transform 1 0 2040 0 1 81061
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2446
timestamp 1649977179
transform 1 0 7208 0 1 82013
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2447
timestamp 1649977179
transform 1 0 7208 0 1 81469
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2448
timestamp 1649977179
transform 1 0 5440 0 1 82013
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2449
timestamp 1649977179
transform 1 0 5440 0 1 81469
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2450
timestamp 1649977179
transform 1 0 17136 0 1 82013
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2451
timestamp 1649977179
transform 1 0 17136 0 1 81469
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2452
timestamp 1649977179
transform 1 0 15640 0 1 82013
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2453
timestamp 1649977179
transform 1 0 15640 0 1 81469
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2454
timestamp 1649977179
transform 1 0 14008 0 1 82013
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2455
timestamp 1649977179
transform 1 0 14008 0 1 81469
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2456
timestamp 1649977179
transform 1 0 12104 0 1 82013
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2457
timestamp 1649977179
transform 1 0 12104 0 1 81469
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2458
timestamp 1649977179
transform 1 0 10472 0 1 82013
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2459
timestamp 1649977179
transform 1 0 10472 0 1 81469
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2460
timestamp 1649977179
transform 1 0 8704 0 1 82013
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2461
timestamp 1649977179
transform 1 0 8704 0 1 81469
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2462
timestamp 1649977179
transform 1 0 33456 0 1 77117
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2463
timestamp 1649977179
transform 1 0 31008 0 1 77117
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2464
timestamp 1649977179
transform 1 0 28696 0 1 77117
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2465
timestamp 1649977179
transform 1 0 28968 0 1 76981
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2466
timestamp 1649977179
transform 1 0 28968 0 1 73037
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2467
timestamp 1649977179
transform 1 0 31280 0 1 76573
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2468
timestamp 1649977179
transform 1 0 31280 0 1 75893
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2469
timestamp 1649977179
transform 1 0 33728 0 1 76573
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2470
timestamp 1649977179
transform 1 0 33728 0 1 75893
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2471
timestamp 1649977179
transform 1 0 28968 0 1 76573
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2472
timestamp 1649977179
transform 1 0 28968 0 1 75893
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2473
timestamp 1649977179
transform 1 0 34000 0 1 73173
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2474
timestamp 1649977179
transform 1 0 34000 0 1 75077
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2475
timestamp 1649977179
transform 1 0 34000 0 1 75213
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2476
timestamp 1649977179
transform 1 0 34000 0 1 76981
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2477
timestamp 1649977179
transform 1 0 31552 0 1 73173
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2478
timestamp 1649977179
transform 1 0 31552 0 1 75077
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2479
timestamp 1649977179
transform 1 0 31416 0 1 75213
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2480
timestamp 1649977179
transform 1 0 31416 0 1 76981
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2481
timestamp 1649977179
transform 1 0 28968 0 1 73173
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2482
timestamp 1649977179
transform 1 0 28968 0 1 75077
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2483
timestamp 1649977179
transform 1 0 28832 0 1 75213
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2484
timestamp 1649977179
transform 1 0 20672 0 1 82013
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2485
timestamp 1649977179
transform 1 0 20672 0 1 81469
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2486
timestamp 1649977179
transform 1 0 18904 0 1 82013
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2487
timestamp 1649977179
transform 1 0 18904 0 1 81469
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2488
timestamp 1649977179
transform 1 0 23936 0 1 81469
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2489
timestamp 1649977179
transform 1 0 22168 0 1 82013
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2490
timestamp 1649977179
transform 1 0 22168 0 1 81469
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2491
timestamp 1649977179
transform 1 0 23936 0 1 82013
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2492
timestamp 1649977179
transform 1 0 25704 0 1 82013
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2493
timestamp 1649977179
transform 1 0 25704 0 1 81469
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2494
timestamp 1649977179
transform 1 0 34136 0 1 82013
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2495
timestamp 1649977179
transform 1 0 34136 0 1 81469
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2496
timestamp 1649977179
transform 1 0 32368 0 1 82013
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2497
timestamp 1649977179
transform 1 0 32368 0 1 81469
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2498
timestamp 1649977179
transform 1 0 30600 0 1 82013
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2499
timestamp 1649977179
transform 1 0 30600 0 1 81469
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2500
timestamp 1649977179
transform 1 0 28968 0 1 82013
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2501
timestamp 1649977179
transform 1 0 28968 0 1 81469
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2502
timestamp 1649977179
transform 1 0 27200 0 1 82013
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2503
timestamp 1649977179
transform 1 0 27200 0 1 81469
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2504
timestamp 1649977179
transform 1 0 1224 0 1 72629
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2505
timestamp 1649977179
transform 1 0 53176 0 1 70997
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2506
timestamp 1649977179
transform 1 0 52496 0 1 70997
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2507
timestamp 1649977179
transform 1 0 61200 0 1 70997
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2508
timestamp 1649977179
transform 1 0 61200 0 1 71405
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2509
timestamp 1649977179
transform 1 0 52496 0 1 71405
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2510
timestamp 1649977179
transform 1 0 56032 0 1 71405
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2511
timestamp 1649977179
transform 1 0 59976 0 1 70997
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2512
timestamp 1649977179
transform 1 0 59976 0 1 71405
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2513
timestamp 1649977179
transform 1 0 59432 0 1 71405
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2514
timestamp 1649977179
transform 1 0 59432 0 1 70997
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2515
timestamp 1649977179
transform 1 0 56032 0 1 70997
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2516
timestamp 1649977179
transform 1 0 68136 0 1 71405
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2517
timestamp 1649977179
transform 1 0 68136 0 1 70997
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2518
timestamp 1649977179
transform 1 0 54944 0 1 70997
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2519
timestamp 1649977179
transform 1 0 59432 0 1 71541
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2520
timestamp 1649977179
transform 1 0 67456 0 1 70997
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2521
timestamp 1649977179
transform 1 0 67456 0 1 71405
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2522
timestamp 1649977179
transform 1 0 66912 0 1 71405
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2523
timestamp 1649977179
transform 1 0 66912 0 1 70997
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2524
timestamp 1649977179
transform 1 0 54944 0 1 71405
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2525
timestamp 1649977179
transform 1 0 54400 0 1 71405
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2526
timestamp 1649977179
transform 1 0 66096 0 1 70997
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2527
timestamp 1649977179
transform 1 0 66096 0 1 71405
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2528
timestamp 1649977179
transform 1 0 54400 0 1 70997
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2529
timestamp 1649977179
transform 1 0 58616 0 1 70997
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2530
timestamp 1649977179
transform 1 0 65008 0 1 70997
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2531
timestamp 1649977179
transform 1 0 65008 0 1 71405
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2532
timestamp 1649977179
transform 1 0 58616 0 1 71405
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2533
timestamp 1649977179
transform 1 0 53312 0 1 70997
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2534
timestamp 1649977179
transform 1 0 53312 0 1 71405
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2535
timestamp 1649977179
transform 1 0 57392 0 1 70997
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2536
timestamp 1649977179
transform 1 0 63648 0 1 70997
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2537
timestamp 1649977179
transform 1 0 63648 0 1 71405
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2538
timestamp 1649977179
transform 1 0 63104 0 1 71405
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2539
timestamp 1649977179
transform 1 0 63104 0 1 70997
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2540
timestamp 1649977179
transform 1 0 57392 0 1 71405
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2541
timestamp 1649977179
transform 1 0 53176 0 1 71405
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2542
timestamp 1649977179
transform 1 0 62424 0 1 70997
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2543
timestamp 1649977179
transform 1 0 62424 0 1 71405
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2544
timestamp 1649977179
transform 1 0 61880 0 1 71405
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2545
timestamp 1649977179
transform 1 0 61880 0 1 70997
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2546
timestamp 1649977179
transform 1 0 45696 0 1 70997
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2547
timestamp 1649977179
transform 1 0 44608 0 1 70861
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2548
timestamp 1649977179
transform 1 0 44608 0 1 71405
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2549
timestamp 1649977179
transform 1 0 36176 0 1 70997
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2550
timestamp 1649977179
transform 1 0 36176 0 1 71405
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2551
timestamp 1649977179
transform 1 0 38216 0 1 71405
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2552
timestamp 1649977179
transform 1 0 38216 0 1 70997
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2553
timestamp 1649977179
transform 1 0 43248 0 1 71405
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2554
timestamp 1649977179
transform 1 0 43248 0 1 70997
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2555
timestamp 1649977179
transform 1 0 37536 0 1 70997
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2556
timestamp 1649977179
transform 1 0 37536 0 1 71405
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2557
timestamp 1649977179
transform 1 0 42432 0 1 70997
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2558
timestamp 1649977179
transform 1 0 42432 0 1 71405
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2559
timestamp 1649977179
transform 1 0 41888 0 1 71405
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2560
timestamp 1649977179
transform 1 0 41888 0 1 70997
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2561
timestamp 1649977179
transform 1 0 34408 0 1 71405
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2562
timestamp 1649977179
transform 1 0 34408 0 1 70997
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2563
timestamp 1649977179
transform 1 0 36992 0 1 71405
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2564
timestamp 1649977179
transform 1 0 36992 0 1 70997
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2565
timestamp 1649977179
transform 1 0 50728 0 1 71405
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2566
timestamp 1649977179
transform 1 0 50728 0 1 70997
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2567
timestamp 1649977179
transform 1 0 49912 0 1 70997
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2568
timestamp 1649977179
transform 1 0 49912 0 1 71405
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2569
timestamp 1649977179
transform 1 0 41208 0 1 70997
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2570
timestamp 1649977179
transform 1 0 41208 0 1 71405
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2571
timestamp 1649977179
transform 1 0 35768 0 1 71405
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2572
timestamp 1649977179
transform 1 0 35768 0 1 70997
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2573
timestamp 1649977179
transform 1 0 48688 0 1 70997
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2574
timestamp 1649977179
transform 1 0 48688 0 1 71405
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2575
timestamp 1649977179
transform 1 0 40664 0 1 71405
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2576
timestamp 1649977179
transform 1 0 40664 0 1 70997
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2577
timestamp 1649977179
transform 1 0 46920 0 1 71405
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2578
timestamp 1649977179
transform 1 0 46920 0 1 70997
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2579
timestamp 1649977179
transform 1 0 39984 0 1 70997
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2580
timestamp 1649977179
transform 1 0 39984 0 1 71405
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2581
timestamp 1649977179
transform 1 0 46240 0 1 70997
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2582
timestamp 1649977179
transform 1 0 46240 0 1 71405
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2583
timestamp 1649977179
transform 1 0 34952 0 1 70997
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2584
timestamp 1649977179
transform 1 0 34952 0 1 71405
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2585
timestamp 1649977179
transform 1 0 45696 0 1 71405
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2586
timestamp 1649977179
transform 1 0 48688 0 1 75893
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2587
timestamp 1649977179
transform 1 0 48960 0 1 73173
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2588
timestamp 1649977179
transform 1 0 48960 0 1 75077
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2589
timestamp 1649977179
transform 1 0 48960 0 1 75213
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2590
timestamp 1649977179
transform 1 0 46376 0 1 76573
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2591
timestamp 1649977179
transform 1 0 46376 0 1 75893
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2592
timestamp 1649977179
transform 1 0 48960 0 1 76981
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2593
timestamp 1649977179
transform 1 0 46512 0 1 73173
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2594
timestamp 1649977179
transform 1 0 51136 0 1 77117
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2595
timestamp 1649977179
transform 1 0 48552 0 1 77117
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2596
timestamp 1649977179
transform 1 0 46104 0 1 77117
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2597
timestamp 1649977179
transform 1 0 43520 0 1 77117
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2598
timestamp 1649977179
transform 1 0 46512 0 1 75077
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2599
timestamp 1649977179
transform 1 0 46512 0 1 75213
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2600
timestamp 1649977179
transform 1 0 46512 0 1 76981
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2601
timestamp 1649977179
transform 1 0 44064 0 1 73173
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2602
timestamp 1649977179
transform 1 0 44064 0 1 75077
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2603
timestamp 1649977179
transform 1 0 43792 0 1 75213
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2604
timestamp 1649977179
transform 1 0 43928 0 1 76981
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2605
timestamp 1649977179
transform 1 0 43928 0 1 76573
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2606
timestamp 1649977179
transform 1 0 43928 0 1 75893
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2607
timestamp 1649977179
transform 1 0 43656 0 1 75893
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2608
timestamp 1649977179
transform 1 0 43656 0 1 76573
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2609
timestamp 1649977179
transform 1 0 48688 0 1 76573
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2610
timestamp 1649977179
transform 1 0 39032 0 1 75077
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2611
timestamp 1649977179
transform 1 0 39032 0 1 75213
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2612
timestamp 1649977179
transform 1 0 38624 0 1 75893
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2613
timestamp 1649977179
transform 1 0 38624 0 1 76573
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2614
timestamp 1649977179
transform 1 0 36312 0 1 76573
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2615
timestamp 1649977179
transform 1 0 36312 0 1 75893
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2616
timestamp 1649977179
transform 1 0 39032 0 1 76981
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2617
timestamp 1649977179
transform 1 0 41072 0 1 77117
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2618
timestamp 1649977179
transform 1 0 38488 0 1 77117
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2619
timestamp 1649977179
transform 1 0 36176 0 1 77117
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2620
timestamp 1649977179
transform 1 0 36448 0 1 73173
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2621
timestamp 1649977179
transform 1 0 36448 0 1 75077
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2622
timestamp 1649977179
transform 1 0 36448 0 1 75213
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2623
timestamp 1649977179
transform 1 0 36448 0 1 76981
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2624
timestamp 1649977179
transform 1 0 41480 0 1 73173
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2625
timestamp 1649977179
transform 1 0 41344 0 1 76573
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2626
timestamp 1649977179
transform 1 0 41344 0 1 75893
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2627
timestamp 1649977179
transform 1 0 41480 0 1 75077
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2628
timestamp 1649977179
transform 1 0 41480 0 1 75213
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2629
timestamp 1649977179
transform 1 0 41480 0 1 76981
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2630
timestamp 1649977179
transform 1 0 39032 0 1 73173
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2631
timestamp 1649977179
transform 1 0 38896 0 1 76573
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2632
timestamp 1649977179
transform 1 0 38896 0 1 75893
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2633
timestamp 1649977179
transform 1 0 35632 0 1 82013
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2634
timestamp 1649977179
transform 1 0 35632 0 1 81469
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2635
timestamp 1649977179
transform 1 0 42432 0 1 82013
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2636
timestamp 1649977179
transform 1 0 42432 0 1 81469
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2637
timestamp 1649977179
transform 1 0 40664 0 1 82013
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2638
timestamp 1649977179
transform 1 0 40664 0 1 81469
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2639
timestamp 1649977179
transform 1 0 39168 0 1 82013
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2640
timestamp 1649977179
transform 1 0 39168 0 1 81469
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2641
timestamp 1649977179
transform 1 0 37536 0 1 82013
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2642
timestamp 1649977179
transform 1 0 37536 0 1 81469
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2643
timestamp 1649977179
transform 1 0 47464 0 1 82013
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2644
timestamp 1649977179
transform 1 0 47464 0 1 81469
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2645
timestamp 1649977179
transform 1 0 45696 0 1 82013
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2646
timestamp 1649977179
transform 1 0 45696 0 1 81469
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2647
timestamp 1649977179
transform 1 0 49232 0 1 82013
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2648
timestamp 1649977179
transform 1 0 49232 0 1 81469
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2649
timestamp 1649977179
transform 1 0 44200 0 1 82013
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2650
timestamp 1649977179
transform 1 0 44200 0 1 81469
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2651
timestamp 1649977179
transform 1 0 50728 0 1 82013
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2652
timestamp 1649977179
transform 1 0 50728 0 1 81469
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2653
timestamp 1649977179
transform 1 0 66096 0 1 77117
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2654
timestamp 1649977179
transform 1 0 63648 0 1 77117
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2655
timestamp 1649977179
transform 1 0 60928 0 1 77117
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2656
timestamp 1649977179
transform 1 0 66368 0 1 76573
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2657
timestamp 1649977179
transform 1 0 66368 0 1 75893
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2658
timestamp 1649977179
transform 1 0 63784 0 1 76573
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2659
timestamp 1649977179
transform 1 0 66504 0 1 73173
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2660
timestamp 1649977179
transform 1 0 66504 0 1 75077
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2661
timestamp 1649977179
transform 1 0 66504 0 1 75213
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2662
timestamp 1649977179
transform 1 0 66504 0 1 76981
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2663
timestamp 1649977179
transform 1 0 63920 0 1 73173
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2664
timestamp 1649977179
transform 1 0 63920 0 1 75077
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2665
timestamp 1649977179
transform 1 0 63920 0 1 75213
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2666
timestamp 1649977179
transform 1 0 63920 0 1 76981
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2667
timestamp 1649977179
transform 1 0 61472 0 1 73173
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2668
timestamp 1649977179
transform 1 0 61472 0 1 75077
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2669
timestamp 1649977179
transform 1 0 61472 0 1 75213
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2670
timestamp 1649977179
transform 1 0 61472 0 1 77117
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2671
timestamp 1649977179
transform 1 0 63784 0 1 75893
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2672
timestamp 1649977179
transform 1 0 61336 0 1 76573
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2673
timestamp 1649977179
transform 1 0 61336 0 1 75893
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2674
timestamp 1649977179
transform 1 0 58480 0 1 77117
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2675
timestamp 1649977179
transform 1 0 56168 0 1 77117
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2676
timestamp 1649977179
transform 1 0 53584 0 1 77117
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2677
timestamp 1649977179
transform 1 0 59024 0 1 73173
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2678
timestamp 1649977179
transform 1 0 59024 0 1 75077
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2679
timestamp 1649977179
transform 1 0 58888 0 1 75213
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2680
timestamp 1649977179
transform 1 0 58888 0 1 76981
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2681
timestamp 1649977179
transform 1 0 56440 0 1 75213
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2682
timestamp 1649977179
transform 1 0 56440 0 1 76981
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2683
timestamp 1649977179
transform 1 0 56304 0 1 75077
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2684
timestamp 1649977179
transform 1 0 56304 0 1 73173
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2685
timestamp 1649977179
transform 1 0 53992 0 1 73173
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2686
timestamp 1649977179
transform 1 0 53992 0 1 75077
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2687
timestamp 1649977179
transform 1 0 53856 0 1 75213
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2688
timestamp 1649977179
transform 1 0 53856 0 1 76981
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2689
timestamp 1649977179
transform 1 0 51544 0 1 73173
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2690
timestamp 1649977179
transform 1 0 51544 0 1 75077
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2691
timestamp 1649977179
transform 1 0 59432 0 1 75757
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2692
timestamp 1649977179
transform 1 0 51408 0 1 76981
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2693
timestamp 1649977179
transform 1 0 58752 0 1 76573
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2694
timestamp 1649977179
transform 1 0 58752 0 1 75893
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2695
timestamp 1649977179
transform 1 0 56168 0 1 75893
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2696
timestamp 1649977179
transform 1 0 56168 0 1 76573
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2697
timestamp 1649977179
transform 1 0 56304 0 1 76573
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2698
timestamp 1649977179
transform 1 0 56304 0 1 75893
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2699
timestamp 1649977179
transform 1 0 53720 0 1 76573
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2700
timestamp 1649977179
transform 1 0 53720 0 1 75893
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2701
timestamp 1649977179
transform 1 0 51408 0 1 76573
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2702
timestamp 1649977179
transform 1 0 51408 0 1 75893
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2703
timestamp 1649977179
transform 1 0 59160 0 1 82013
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2704
timestamp 1649977179
transform 1 0 59160 0 1 81469
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2705
timestamp 1649977179
transform 1 0 57664 0 1 82013
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2706
timestamp 1649977179
transform 1 0 57664 0 1 81469
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2707
timestamp 1649977179
transform 1 0 55896 0 1 82013
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2708
timestamp 1649977179
transform 1 0 55896 0 1 81469
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2709
timestamp 1649977179
transform 1 0 54128 0 1 82013
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2710
timestamp 1649977179
transform 1 0 54128 0 1 81469
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2711
timestamp 1649977179
transform 1 0 52632 0 1 82013
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2712
timestamp 1649977179
transform 1 0 52632 0 1 81469
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2713
timestamp 1649977179
transform 1 0 67592 0 1 82013
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2714
timestamp 1649977179
transform 1 0 67592 0 1 81469
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2715
timestamp 1649977179
transform 1 0 65824 0 1 82013
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2716
timestamp 1649977179
transform 1 0 65824 0 1 81469
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2717
timestamp 1649977179
transform 1 0 64192 0 1 82013
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2718
timestamp 1649977179
transform 1 0 64192 0 1 81469
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2719
timestamp 1649977179
transform 1 0 62696 0 1 82013
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2720
timestamp 1649977179
transform 1 0 62696 0 1 81469
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2721
timestamp 1649977179
transform 1 0 60792 0 1 82013
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2722
timestamp 1649977179
transform 1 0 60792 0 1 81469
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2723
timestamp 1649977179
transform 1 0 51272 0 1 75213
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2724
timestamp 1649977179
transform 1 0 51272 0 1 70997
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2725
timestamp 1649977179
transform 1 0 51272 0 1 71405
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2726
timestamp 1649977179
transform 1 0 135320 0 1 43933
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2727
timestamp 1649977179
transform 1 0 135320 0 1 45701
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2728
timestamp 1649977179
transform 1 0 135320 0 1 42301
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2729
timestamp 1649977179
transform 1 0 135320 0 1 50733
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2730
timestamp 1649977179
transform 1 0 135320 0 1 47469
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2731
timestamp 1649977179
transform 1 0 135320 0 1 48965
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2732
timestamp 1649977179
transform 1 0 114784 0 1 43525
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2733
timestamp 1649977179
transform 1 0 114784 0 1 43797
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2734
timestamp 1649977179
transform 1 0 115872 0 1 45973
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2735
timestamp 1649977179
transform 1 0 115464 0 1 45837
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2736
timestamp 1649977179
transform 1 0 115872 0 1 46245
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2737
timestamp 1649977179
transform 1 0 115464 0 1 45565
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2738
timestamp 1649977179
transform 1 0 115056 0 1 42301
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2739
timestamp 1649977179
transform 1 0 115056 0 1 42029
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2740
timestamp 1649977179
transform 1 0 116008 0 1 46653
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2741
timestamp 1649977179
transform 1 0 114376 0 1 45565
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2742
timestamp 1649977179
transform 1 0 114376 0 1 45837
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2743
timestamp 1649977179
transform 1 0 116008 0 1 46381
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2744
timestamp 1649977179
transform 1 0 115328 0 1 45429
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2745
timestamp 1649977179
transform 1 0 115464 0 1 44613
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2746
timestamp 1649977179
transform 1 0 114648 0 1 42301
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2747
timestamp 1649977179
transform 1 0 114648 0 1 42029
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2748
timestamp 1649977179
transform 1 0 115192 0 1 45429
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2749
timestamp 1649977179
transform 1 0 114376 0 1 45973
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2750
timestamp 1649977179
transform 1 0 114784 0 1 45973
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2751
timestamp 1649977179
transform 1 0 114784 0 1 46245
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2752
timestamp 1649977179
transform 1 0 114648 0 1 46653
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2753
timestamp 1649977179
transform 1 0 114648 0 1 46381
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2754
timestamp 1649977179
transform 1 0 116008 0 1 42029
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2755
timestamp 1649977179
transform 1 0 116008 0 1 42301
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2756
timestamp 1649977179
transform 1 0 115192 0 1 45157
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2757
timestamp 1649977179
transform 1 0 114648 0 1 44341
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2758
timestamp 1649977179
transform 1 0 114648 0 1 44613
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2759
timestamp 1649977179
transform 1 0 114648 0 1 45021
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2760
timestamp 1649977179
transform 1 0 116008 0 1 45837
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2761
timestamp 1649977179
transform 1 0 116008 0 1 45565
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2762
timestamp 1649977179
transform 1 0 115056 0 1 42845
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2763
timestamp 1649977179
transform 1 0 114648 0 1 44749
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2764
timestamp 1649977179
transform 1 0 115056 0 1 43117
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2765
timestamp 1649977179
transform 1 0 114376 0 1 46245
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2766
timestamp 1649977179
transform 1 0 115872 0 1 42437
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2767
timestamp 1649977179
transform 1 0 115872 0 1 42709
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2768
timestamp 1649977179
transform 1 0 114240 0 1 42301
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2769
timestamp 1649977179
transform 1 0 114240 0 1 42029
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2770
timestamp 1649977179
transform 1 0 114376 0 1 43525
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2771
timestamp 1649977179
transform 1 0 115328 0 1 46245
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2772
timestamp 1649977179
transform 1 0 115872 0 1 45429
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2773
timestamp 1649977179
transform 1 0 115872 0 1 45157
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2774
timestamp 1649977179
transform 1 0 114376 0 1 41893
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2775
timestamp 1649977179
transform 1 0 115328 0 1 45973
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2776
timestamp 1649977179
transform 1 0 114376 0 1 43797
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2777
timestamp 1649977179
transform 1 0 114376 0 1 44205
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2778
timestamp 1649977179
transform 1 0 114376 0 1 43933
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2779
timestamp 1649977179
transform 1 0 115872 0 1 45021
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2780
timestamp 1649977179
transform 1 0 115872 0 1 44749
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2781
timestamp 1649977179
transform 1 0 114784 0 1 42709
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2782
timestamp 1649977179
transform 1 0 114376 0 1 45021
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2783
timestamp 1649977179
transform 1 0 114240 0 1 42709
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2784
timestamp 1649977179
transform 1 0 114240 0 1 42437
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2785
timestamp 1649977179
transform 1 0 115192 0 1 45973
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2786
timestamp 1649977179
transform 1 0 115192 0 1 46245
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2787
timestamp 1649977179
transform 1 0 115192 0 1 41893
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2788
timestamp 1649977179
transform 1 0 115464 0 1 45973
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2789
timestamp 1649977179
transform 1 0 115328 0 1 41893
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2790
timestamp 1649977179
transform 1 0 114648 0 1 45837
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2791
timestamp 1649977179
transform 1 0 114648 0 1 45565
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2792
timestamp 1649977179
transform 1 0 114784 0 1 45429
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2793
timestamp 1649977179
transform 1 0 115872 0 1 41893
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2794
timestamp 1649977179
transform 1 0 114240 0 1 44613
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2795
timestamp 1649977179
transform 1 0 114784 0 1 45157
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2796
timestamp 1649977179
transform 1 0 114376 0 1 45429
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2797
timestamp 1649977179
transform 1 0 114376 0 1 45157
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2798
timestamp 1649977179
transform 1 0 115464 0 1 46245
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2799
timestamp 1649977179
transform 1 0 114784 0 1 44205
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2800
timestamp 1649977179
transform 1 0 113696 0 1 45429
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2801
timestamp 1649977179
transform 1 0 113696 0 1 45157
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2802
timestamp 1649977179
transform 1 0 114784 0 1 43933
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2803
timestamp 1649977179
transform 1 0 114376 0 1 44749
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2804
timestamp 1649977179
transform 1 0 115192 0 1 43525
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2805
timestamp 1649977179
transform 1 0 116008 0 1 42845
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2806
timestamp 1649977179
transform 1 0 116008 0 1 43117
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2807
timestamp 1649977179
transform 1 0 116008 0 1 43525
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2808
timestamp 1649977179
transform 1 0 116008 0 1 43253
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2809
timestamp 1649977179
transform 1 0 114784 0 1 41893
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2810
timestamp 1649977179
transform 1 0 112336 0 1 45021
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2811
timestamp 1649977179
transform 1 0 112336 0 1 44613
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2812
timestamp 1649977179
transform 1 0 115192 0 1 43797
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2813
timestamp 1649977179
transform 1 0 114240 0 1 46653
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2814
timestamp 1649977179
transform 1 0 114240 0 1 46381
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2815
timestamp 1649977179
transform 1 0 114240 0 1 44341
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2816
timestamp 1649977179
transform 1 0 114784 0 1 42437
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2817
timestamp 1649977179
transform 1 0 115328 0 1 45157
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2818
timestamp 1649977179
transform 1 0 115464 0 1 44341
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2819
timestamp 1649977179
transform 1 0 109344 0 1 43389
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2820
timestamp 1649977179
transform 1 0 109344 0 1 43661
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2821
timestamp 1649977179
transform 1 0 109344 0 1 42845
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2822
timestamp 1649977179
transform 1 0 109344 0 1 43253
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2823
timestamp 1649977179
transform 1 0 109480 0 1 46517
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2824
timestamp 1649977179
transform 1 0 109344 0 1 42981
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2825
timestamp 1649977179
transform 1 0 109344 0 1 42573
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2826
timestamp 1649977179
transform 1 0 109344 0 1 46925
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2827
timestamp 1649977179
transform 1 0 109344 0 1 47197
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2828
timestamp 1649977179
transform 1 0 114376 0 1 48557
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2829
timestamp 1649977179
transform 1 0 114376 0 1 48285
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2830
timestamp 1649977179
transform 1 0 115328 0 1 48013
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2831
timestamp 1649977179
transform 1 0 115328 0 1 48285
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2832
timestamp 1649977179
transform 1 0 115056 0 1 47741
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2833
timestamp 1649977179
transform 1 0 115056 0 1 47469
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2834
timestamp 1649977179
transform 1 0 115600 0 1 49917
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2835
timestamp 1649977179
transform 1 0 115600 0 1 50189
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2836
timestamp 1649977179
transform 1 0 114240 0 1 48149
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2837
timestamp 1649977179
transform 1 0 114240 0 1 47877
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2838
timestamp 1649977179
transform 1 0 116008 0 1 48693
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2839
timestamp 1649977179
transform 1 0 116008 0 1 48965
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2840
timestamp 1649977179
transform 1 0 114240 0 1 51821
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2841
timestamp 1649977179
transform 1 0 115056 0 1 51005
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2842
timestamp 1649977179
transform 1 0 115056 0 1 50733
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2843
timestamp 1649977179
transform 1 0 115600 0 1 48965
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2844
timestamp 1649977179
transform 1 0 115600 0 1 48693
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2845
timestamp 1649977179
transform 1 0 115464 0 1 48557
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2846
timestamp 1649977179
transform 1 0 115464 0 1 48285
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2847
timestamp 1649977179
transform 1 0 115192 0 1 51685
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2848
timestamp 1649977179
transform 1 0 114240 0 1 48693
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2849
timestamp 1649977179
transform 1 0 114240 0 1 48965
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2850
timestamp 1649977179
transform 1 0 114376 0 1 49373
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2851
timestamp 1649977179
transform 1 0 115192 0 1 51413
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2852
timestamp 1649977179
transform 1 0 114376 0 1 49101
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2853
timestamp 1649977179
transform 1 0 115872 0 1 49917
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2854
timestamp 1649977179
transform 1 0 115872 0 1 50189
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2855
timestamp 1649977179
transform 1 0 115872 0 1 50597
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2856
timestamp 1649977179
transform 1 0 115872 0 1 50325
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2857
timestamp 1649977179
transform 1 0 116008 0 1 50733
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2858
timestamp 1649977179
transform 1 0 116008 0 1 51005
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2859
timestamp 1649977179
transform 1 0 115872 0 1 49781
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2860
timestamp 1649977179
transform 1 0 115872 0 1 49509
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2861
timestamp 1649977179
transform 1 0 115872 0 1 49101
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2862
timestamp 1649977179
transform 1 0 115872 0 1 49373
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2863
timestamp 1649977179
transform 1 0 114240 0 1 50189
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2864
timestamp 1649977179
transform 1 0 114784 0 1 50325
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2865
timestamp 1649977179
transform 1 0 115328 0 1 47061
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2866
timestamp 1649977179
transform 1 0 115056 0 1 48285
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2867
timestamp 1649977179
transform 1 0 115056 0 1 48557
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2868
timestamp 1649977179
transform 1 0 114376 0 1 50325
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2869
timestamp 1649977179
transform 1 0 115872 0 1 51141
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2870
timestamp 1649977179
transform 1 0 115872 0 1 51413
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2871
timestamp 1649977179
transform 1 0 115328 0 1 49781
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2872
timestamp 1649977179
transform 1 0 114376 0 1 50597
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2873
timestamp 1649977179
transform 1 0 114240 0 1 51005
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2874
timestamp 1649977179
transform 1 0 114240 0 1 50733
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2875
timestamp 1649977179
transform 1 0 115872 0 1 48013
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2876
timestamp 1649977179
transform 1 0 115872 0 1 48285
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2877
timestamp 1649977179
transform 1 0 115328 0 1 49509
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2878
timestamp 1649977179
transform 1 0 115192 0 1 49781
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2879
timestamp 1649977179
transform 1 0 115192 0 1 49509
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2880
timestamp 1649977179
transform 1 0 114240 0 1 49917
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2881
timestamp 1649977179
transform 1 0 114784 0 1 49917
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2882
timestamp 1649977179
transform 1 0 115872 0 1 47061
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2883
timestamp 1649977179
transform 1 0 115872 0 1 47469
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2884
timestamp 1649977179
transform 1 0 115872 0 1 47197
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2885
timestamp 1649977179
transform 1 0 114240 0 1 49509
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2886
timestamp 1649977179
transform 1 0 114648 0 1 51005
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2887
timestamp 1649977179
transform 1 0 114648 0 1 50733
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2888
timestamp 1649977179
transform 1 0 114784 0 1 50189
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2889
timestamp 1649977179
transform 1 0 114648 0 1 49373
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2890
timestamp 1649977179
transform 1 0 114648 0 1 49101
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2891
timestamp 1649977179
transform 1 0 114784 0 1 47877
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2892
timestamp 1649977179
transform 1 0 114784 0 1 48149
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2893
timestamp 1649977179
transform 1 0 114240 0 1 49781
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2894
timestamp 1649977179
transform 1 0 114648 0 1 48965
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2895
timestamp 1649977179
transform 1 0 114648 0 1 48693
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2896
timestamp 1649977179
transform 1 0 114648 0 1 48285
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2897
timestamp 1649977179
transform 1 0 114648 0 1 48557
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2898
timestamp 1649977179
transform 1 0 114648 0 1 49509
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2899
timestamp 1649977179
transform 1 0 114648 0 1 49781
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2900
timestamp 1649977179
transform 1 0 115464 0 1 50733
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2901
timestamp 1649977179
transform 1 0 115464 0 1 51005
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2902
timestamp 1649977179
transform 1 0 114648 0 1 51821
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2903
timestamp 1649977179
transform 1 0 114784 0 1 50597
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2904
timestamp 1649977179
transform 1 0 115328 0 1 46789
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2905
timestamp 1649977179
transform 1 0 115872 0 1 46789
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2906
timestamp 1649977179
transform 1 0 109480 0 1 46789
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2907
timestamp 1649977179
transform 1 0 115464 0 1 54269
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2908
timestamp 1649977179
transform 1 0 115600 0 1 56989
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2909
timestamp 1649977179
transform 1 0 115464 0 1 53317
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2910
timestamp 1649977179
transform 1 0 114240 0 1 52637
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2911
timestamp 1649977179
transform 1 0 114240 0 1 52909
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2912
timestamp 1649977179
transform 1 0 114240 0 1 53317
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2913
timestamp 1649977179
transform 1 0 114240 0 1 53045
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2914
timestamp 1649977179
transform 1 0 115192 0 1 52501
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2915
timestamp 1649977179
transform 1 0 114376 0 1 53725
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2916
timestamp 1649977179
transform 1 0 114376 0 1 54133
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2917
timestamp 1649977179
transform 1 0 114376 0 1 53861
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2918
timestamp 1649977179
transform 1 0 114376 0 1 54949
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2919
timestamp 1649977179
transform 1 0 114376 0 1 54677
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2920
timestamp 1649977179
transform 1 0 114240 0 1 56853
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2921
timestamp 1649977179
transform 1 0 114240 0 1 56581
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2922
timestamp 1649977179
transform 1 0 114240 0 1 56173
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2923
timestamp 1649977179
transform 1 0 114648 0 1 56989
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2924
timestamp 1649977179
transform 1 0 115192 0 1 52909
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2925
timestamp 1649977179
transform 1 0 114240 0 1 52093
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2926
timestamp 1649977179
transform 1 0 115872 0 1 53725
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2927
timestamp 1649977179
transform 1 0 115872 0 1 53453
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2928
timestamp 1649977179
transform 1 0 115872 0 1 54677
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2929
timestamp 1649977179
transform 1 0 115872 0 1 54949
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2930
timestamp 1649977179
transform 1 0 116008 0 1 53861
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2931
timestamp 1649977179
transform 1 0 116008 0 1 54133
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2932
timestamp 1649977179
transform 1 0 116008 0 1 54541
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2933
timestamp 1649977179
transform 1 0 116008 0 1 54269
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2934
timestamp 1649977179
transform 1 0 115192 0 1 52637
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2935
timestamp 1649977179
transform 1 0 115328 0 1 54949
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2936
timestamp 1649977179
transform 1 0 114240 0 1 56445
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2937
timestamp 1649977179
transform 1 0 115328 0 1 54677
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2938
timestamp 1649977179
transform 1 0 114376 0 1 52229
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2939
timestamp 1649977179
transform 1 0 115192 0 1 56989
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2940
timestamp 1649977179
transform 1 0 115192 0 1 52229
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2941
timestamp 1649977179
transform 1 0 116008 0 1 52229
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2942
timestamp 1649977179
transform 1 0 114376 0 1 52501
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2943
timestamp 1649977179
transform 1 0 115328 0 1 56037
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2944
timestamp 1649977179
transform 1 0 115192 0 1 55901
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2945
timestamp 1649977179
transform 1 0 115056 0 1 56445
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2946
timestamp 1649977179
transform 1 0 116008 0 1 55901
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2947
timestamp 1649977179
transform 1 0 116008 0 1 56173
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2948
timestamp 1649977179
transform 1 0 115056 0 1 56173
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2949
timestamp 1649977179
transform 1 0 114240 0 1 56989
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2950
timestamp 1649977179
transform 1 0 115872 0 1 52909
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2951
timestamp 1649977179
transform 1 0 115872 0 1 52637
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2952
timestamp 1649977179
transform 1 0 115192 0 1 54677
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2953
timestamp 1649977179
transform 1 0 116008 0 1 55765
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2954
timestamp 1649977179
transform 1 0 116008 0 1 55493
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2955
timestamp 1649977179
transform 1 0 116008 0 1 55085
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2956
timestamp 1649977179
transform 1 0 116008 0 1 55357
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2957
timestamp 1649977179
transform 1 0 115192 0 1 54949
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2958
timestamp 1649977179
transform 1 0 115328 0 1 55493
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2959
timestamp 1649977179
transform 1 0 115328 0 1 55765
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2960
timestamp 1649977179
transform 1 0 115328 0 1 54133
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2961
timestamp 1649977179
transform 1 0 114784 0 1 56581
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2962
timestamp 1649977179
transform 1 0 114784 0 1 56853
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2963
timestamp 1649977179
transform 1 0 114648 0 1 56445
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2964
timestamp 1649977179
transform 1 0 114648 0 1 56173
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2965
timestamp 1649977179
transform 1 0 115328 0 1 53861
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2966
timestamp 1649977179
transform 1 0 115192 0 1 54133
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2967
timestamp 1649977179
transform 1 0 114648 0 1 53045
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2968
timestamp 1649977179
transform 1 0 114648 0 1 53317
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2969
timestamp 1649977179
transform 1 0 114784 0 1 52229
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2970
timestamp 1649977179
transform 1 0 114784 0 1 52501
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2971
timestamp 1649977179
transform 1 0 114784 0 1 52909
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2972
timestamp 1649977179
transform 1 0 114784 0 1 52637
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2973
timestamp 1649977179
transform 1 0 115192 0 1 53861
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2974
timestamp 1649977179
transform 1 0 114240 0 1 54541
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2975
timestamp 1649977179
transform 1 0 114240 0 1 54269
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2976
timestamp 1649977179
transform 1 0 114784 0 1 54949
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2977
timestamp 1649977179
transform 1 0 114784 0 1 54677
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2978
timestamp 1649977179
transform 1 0 114784 0 1 54269
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2979
timestamp 1649977179
transform 1 0 114784 0 1 54541
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2980
timestamp 1649977179
transform 1 0 114784 0 1 53453
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2981
timestamp 1649977179
transform 1 0 114784 0 1 53725
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2982
timestamp 1649977179
transform 1 0 114784 0 1 54133
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2983
timestamp 1649977179
transform 1 0 114784 0 1 53861
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2984
timestamp 1649977179
transform 1 0 114648 0 1 52093
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2985
timestamp 1649977179
transform 1 0 114376 0 1 53453
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2986
timestamp 1649977179
transform 1 0 115600 0 1 52909
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2987
timestamp 1649977179
transform 1 0 115600 0 1 52637
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2988
timestamp 1649977179
transform 1 0 115464 0 1 53045
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2989
timestamp 1649977179
transform 1 0 115464 0 1 54541
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2990
timestamp 1649977179
transform 1 0 109480 0 1 55493
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2991
timestamp 1649977179
transform 1 0 109480 0 1 55629
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2992
timestamp 1649977179
transform 1 0 109480 0 1 55901
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2993
timestamp 1649977179
transform 1 0 109344 0 1 55629
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2994
timestamp 1649977179
transform 1 0 109344 0 1 56037
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2995
timestamp 1649977179
transform 1 0 109480 0 1 55221
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2996
timestamp 1649977179
transform 1 0 109480 0 1 59845
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2997
timestamp 1649977179
transform 1 0 109480 0 1 58349
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2998
timestamp 1649977179
transform 1 0 109480 0 1 58621
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2999
timestamp 1649977179
transform 1 0 109480 0 1 61069
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3000
timestamp 1649977179
transform 1 0 109480 0 1 60797
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3001
timestamp 1649977179
transform 1 0 109480 0 1 59573
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3002
timestamp 1649977179
transform 1 0 114240 0 1 60797
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3003
timestamp 1649977179
transform 1 0 114240 0 1 60525
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3004
timestamp 1649977179
transform 1 0 115056 0 1 58485
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3005
timestamp 1649977179
transform 1 0 114376 0 1 60389
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3006
timestamp 1649977179
transform 1 0 114376 0 1 60117
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3007
timestamp 1649977179
transform 1 0 114240 0 1 61341
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3008
timestamp 1649977179
transform 1 0 114240 0 1 61613
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3009
timestamp 1649977179
transform 1 0 116008 0 1 61749
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3010
timestamp 1649977179
transform 1 0 116008 0 1 62021
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3011
timestamp 1649977179
transform 1 0 114376 0 1 62157
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3012
timestamp 1649977179
transform 1 0 114240 0 1 61749
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3013
timestamp 1649977179
transform 1 0 114240 0 1 62021
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3014
timestamp 1649977179
transform 1 0 116008 0 1 57397
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3015
timestamp 1649977179
transform 1 0 116008 0 1 57669
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3016
timestamp 1649977179
transform 1 0 115872 0 1 58077
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3017
timestamp 1649977179
transform 1 0 115872 0 1 57805
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3018
timestamp 1649977179
transform 1 0 115872 0 1 61613
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3019
timestamp 1649977179
transform 1 0 115872 0 1 61341
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3020
timestamp 1649977179
transform 1 0 116008 0 1 59437
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3021
timestamp 1649977179
transform 1 0 116008 0 1 59709
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3022
timestamp 1649977179
transform 1 0 116008 0 1 60117
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3023
timestamp 1649977179
transform 1 0 116008 0 1 59845
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3024
timestamp 1649977179
transform 1 0 116008 0 1 58213
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3025
timestamp 1649977179
transform 1 0 116008 0 1 58485
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3026
timestamp 1649977179
transform 1 0 115872 0 1 62157
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3027
timestamp 1649977179
transform 1 0 115872 0 1 59301
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3028
timestamp 1649977179
transform 1 0 115872 0 1 59029
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3029
timestamp 1649977179
transform 1 0 115872 0 1 58621
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3030
timestamp 1649977179
transform 1 0 115872 0 1 58893
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3031
timestamp 1649977179
transform 1 0 114648 0 1 61205
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3032
timestamp 1649977179
transform 1 0 114648 0 1 60933
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3033
timestamp 1649977179
transform 1 0 114784 0 1 62157
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3034
timestamp 1649977179
transform 1 0 114648 0 1 60797
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3035
timestamp 1649977179
transform 1 0 114648 0 1 60525
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3036
timestamp 1649977179
transform 1 0 114648 0 1 60117
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3037
timestamp 1649977179
transform 1 0 114648 0 1 60389
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3038
timestamp 1649977179
transform 1 0 114784 0 1 58485
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3039
timestamp 1649977179
transform 1 0 114784 0 1 58213
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3040
timestamp 1649977179
transform 1 0 114784 0 1 57805
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3041
timestamp 1649977179
transform 1 0 114784 0 1 58077
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3042
timestamp 1649977179
transform 1 0 114648 0 1 57261
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3043
timestamp 1649977179
transform 1 0 114648 0 1 57669
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3044
timestamp 1649977179
transform 1 0 114648 0 1 57397
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3045
timestamp 1649977179
transform 1 0 114648 0 1 61341
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3046
timestamp 1649977179
transform 1 0 114648 0 1 61613
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3047
timestamp 1649977179
transform 1 0 114648 0 1 62021
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3048
timestamp 1649977179
transform 1 0 114648 0 1 61749
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3049
timestamp 1649977179
transform 1 0 114784 0 1 58621
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3050
timestamp 1649977179
transform 1 0 114784 0 1 58893
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3051
timestamp 1649977179
transform 1 0 114784 0 1 59301
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3052
timestamp 1649977179
transform 1 0 114784 0 1 59029
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3053
timestamp 1649977179
transform 1 0 114376 0 1 58621
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3054
timestamp 1649977179
transform 1 0 114376 0 1 58893
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3055
timestamp 1649977179
transform 1 0 114376 0 1 59301
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3056
timestamp 1649977179
transform 1 0 114376 0 1 59029
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3057
timestamp 1649977179
transform 1 0 115192 0 1 57261
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3058
timestamp 1649977179
transform 1 0 115328 0 1 60933
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3059
timestamp 1649977179
transform 1 0 115328 0 1 61205
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3060
timestamp 1649977179
transform 1 0 115328 0 1 60389
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3061
timestamp 1649977179
transform 1 0 115328 0 1 60117
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3062
timestamp 1649977179
transform 1 0 115192 0 1 60389
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3063
timestamp 1649977179
transform 1 0 115192 0 1 60117
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3064
timestamp 1649977179
transform 1 0 115056 0 1 61341
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3065
timestamp 1649977179
transform 1 0 115056 0 1 61613
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3066
timestamp 1649977179
transform 1 0 114240 0 1 58213
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3067
timestamp 1649977179
transform 1 0 114240 0 1 58485
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3068
timestamp 1649977179
transform 1 0 115192 0 1 62157
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3069
timestamp 1649977179
transform 1 0 115328 0 1 58077
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3070
timestamp 1649977179
transform 1 0 115328 0 1 57805
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3071
timestamp 1649977179
transform 1 0 115192 0 1 58077
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3072
timestamp 1649977179
transform 1 0 115192 0 1 57805
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3073
timestamp 1649977179
transform 1 0 114376 0 1 58077
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3074
timestamp 1649977179
transform 1 0 114376 0 1 57805
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3075
timestamp 1649977179
transform 1 0 114240 0 1 61205
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3076
timestamp 1649977179
transform 1 0 114240 0 1 60933
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3077
timestamp 1649977179
transform 1 0 114240 0 1 57261
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3078
timestamp 1649977179
transform 1 0 114240 0 1 57669
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3079
timestamp 1649977179
transform 1 0 114240 0 1 57397
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3080
timestamp 1649977179
transform 1 0 115464 0 1 58893
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3081
timestamp 1649977179
transform 1 0 115464 0 1 58621
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3082
timestamp 1649977179
transform 1 0 115600 0 1 57261
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3083
timestamp 1649977179
transform 1 0 115600 0 1 57669
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3084
timestamp 1649977179
transform 1 0 115600 0 1 57397
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3085
timestamp 1649977179
transform 1 0 115464 0 1 59437
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3086
timestamp 1649977179
transform 1 0 115464 0 1 59709
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3087
timestamp 1649977179
transform 1 0 115600 0 1 61341
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3088
timestamp 1649977179
transform 1 0 115600 0 1 61613
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3089
timestamp 1649977179
transform 1 0 115464 0 1 61749
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3090
timestamp 1649977179
transform 1 0 115464 0 1 62021
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3091
timestamp 1649977179
transform 1 0 115328 0 1 58485
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3092
timestamp 1649977179
transform 1 0 115328 0 1 58213
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3093
timestamp 1649977179
transform 1 0 115056 0 1 58213
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3094
timestamp 1649977179
transform 1 0 135320 0 1 53997
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3095
timestamp 1649977179
transform 1 0 135320 0 1 55901
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3096
timestamp 1649977179
transform 1 0 135320 0 1 52365
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3097
timestamp 1649977179
transform 1 0 133416 0 1 61477
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3098
timestamp 1649977179
transform 1 0 135320 0 1 59165
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3099
timestamp 1649977179
transform 1 0 135320 0 1 57533
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3100
timestamp 1649977179
transform 1 0 135320 0 1 60797
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3101
timestamp 1649977179
transform 1 0 134087 0 1 62058
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3102
timestamp 1649977179
transform 1 0 116008 0 1 51957
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3103
timestamp 1649977179
transform 1 0 94928 0 1 71405
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3104
timestamp 1649977179
transform 1 0 89896 0 1 70997
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3105
timestamp 1649977179
transform 1 0 89896 0 1 71405
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3106
timestamp 1649977179
transform 1 0 86088 0 1 70997
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3107
timestamp 1649977179
transform 1 0 86088 0 1 71405
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3108
timestamp 1649977179
transform 1 0 101864 0 1 71405
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3109
timestamp 1649977179
transform 1 0 101864 0 1 70997
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3110
timestamp 1649977179
transform 1 0 93296 0 1 70861
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3111
timestamp 1649977179
transform 1 0 93296 0 1 71405
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3112
timestamp 1649977179
transform 1 0 89352 0 1 71405
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3113
timestamp 1649977179
transform 1 0 89352 0 1 70997
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3114
timestamp 1649977179
transform 1 0 100912 0 1 71405
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3115
timestamp 1649977179
transform 1 0 100912 0 1 70997
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3116
timestamp 1649977179
transform 1 0 99824 0 1 70997
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3117
timestamp 1649977179
transform 1 0 99824 0 1 71405
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3118
timestamp 1649977179
transform 1 0 92344 0 1 70997
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3119
timestamp 1649977179
transform 1 0 92344 0 1 71405
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3120
timestamp 1649977179
transform 1 0 86904 0 1 71405
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3121
timestamp 1649977179
transform 1 0 86904 0 1 70997
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3122
timestamp 1649977179
transform 1 0 98600 0 1 70997
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3123
timestamp 1649977179
transform 1 0 98600 0 1 71269
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3124
timestamp 1649977179
transform 1 0 88672 0 1 70997
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3125
timestamp 1649977179
transform 1 0 88672 0 1 71405
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3126
timestamp 1649977179
transform 1 0 97376 0 1 70997
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3127
timestamp 1649977179
transform 1 0 97376 0 1 71405
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3128
timestamp 1649977179
transform 1 0 96832 0 1 71405
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3129
timestamp 1649977179
transform 1 0 96832 0 1 70997
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3130
timestamp 1649977179
transform 1 0 88128 0 1 71405
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3131
timestamp 1649977179
transform 1 0 88128 0 1 70997
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3132
timestamp 1649977179
transform 1 0 91120 0 1 70997
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3133
timestamp 1649977179
transform 1 0 91120 0 1 71405
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3134
timestamp 1649977179
transform 1 0 90712 0 1 71405
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3135
timestamp 1649977179
transform 1 0 90712 0 1 70997
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3136
timestamp 1649977179
transform 1 0 95608 0 1 71405
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3137
timestamp 1649977179
transform 1 0 95608 0 1 70997
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3138
timestamp 1649977179
transform 1 0 94928 0 1 70997
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3139
timestamp 1649977179
transform 1 0 79424 0 1 70997
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3140
timestamp 1649977179
transform 1 0 68680 0 1 70997
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3141
timestamp 1649977179
transform 1 0 68680 0 1 71405
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3142
timestamp 1649977179
transform 1 0 78472 0 1 71405
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3143
timestamp 1649977179
transform 1 0 78472 0 1 70997
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3144
timestamp 1649977179
transform 1 0 78200 0 1 71405
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3145
timestamp 1649977179
transform 1 0 78200 0 1 70997
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3146
timestamp 1649977179
transform 1 0 73712 0 1 70997
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3147
timestamp 1649977179
transform 1 0 73712 0 1 71405
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3148
timestamp 1649977179
transform 1 0 77384 0 1 70997
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3149
timestamp 1649977179
transform 1 0 77384 0 1 71405
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3150
timestamp 1649977179
transform 1 0 76840 0 1 71405
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3151
timestamp 1649977179
transform 1 0 76840 0 1 70997
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3152
timestamp 1649977179
transform 1 0 70584 0 1 71405
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3153
timestamp 1649977179
transform 1 0 70584 0 1 70997
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3154
timestamp 1649977179
transform 1 0 72080 0 1 70861
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3155
timestamp 1649977179
transform 1 0 72080 0 1 71405
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3156
timestamp 1649977179
transform 1 0 84592 0 1 70997
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3157
timestamp 1649977179
transform 1 0 84592 0 1 71405
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3158
timestamp 1649977179
transform 1 0 76160 0 1 70997
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3159
timestamp 1649977179
transform 1 0 76160 0 1 71405
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3160
timestamp 1649977179
transform 1 0 72216 0 1 71405
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3161
timestamp 1649977179
transform 1 0 72216 0 1 70997
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3162
timestamp 1649977179
transform 1 0 83640 0 1 70997
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3163
timestamp 1649977179
transform 1 0 83640 0 1 71405
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3164
timestamp 1649977179
transform 1 0 83096 0 1 71405
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3165
timestamp 1649977179
transform 1 0 83096 0 1 70997
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3166
timestamp 1649977179
transform 1 0 75616 0 1 71405
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3167
timestamp 1649977179
transform 1 0 75616 0 1 70997
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3168
timestamp 1649977179
transform 1 0 82416 0 1 70997
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3169
timestamp 1649977179
transform 1 0 82416 0 1 71405
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3170
timestamp 1649977179
transform 1 0 81872 0 1 71405
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3171
timestamp 1649977179
transform 1 0 81872 0 1 70997
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3172
timestamp 1649977179
transform 1 0 74936 0 1 70997
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3173
timestamp 1649977179
transform 1 0 74936 0 1 71405
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3174
timestamp 1649977179
transform 1 0 69904 0 1 70997
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3175
timestamp 1649977179
transform 1 0 69904 0 1 71405
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3176
timestamp 1649977179
transform 1 0 80648 0 1 71405
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3177
timestamp 1649977179
transform 1 0 80648 0 1 70997
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3178
timestamp 1649977179
transform 1 0 79968 0 1 70997
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3179
timestamp 1649977179
transform 1 0 79968 0 1 71405
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3180
timestamp 1649977179
transform 1 0 74392 0 1 71405
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3181
timestamp 1649977179
transform 1 0 74392 0 1 70997
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3182
timestamp 1649977179
transform 1 0 79424 0 1 71405
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3183
timestamp 1649977179
transform 1 0 81464 0 1 73173
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3184
timestamp 1649977179
transform 1 0 78744 0 1 76573
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3185
timestamp 1649977179
transform 1 0 83776 0 1 76573
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3186
timestamp 1649977179
transform 1 0 83776 0 1 75893
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3187
timestamp 1649977179
transform 1 0 78744 0 1 75893
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3188
timestamp 1649977179
transform 1 0 81464 0 1 75077
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3189
timestamp 1649977179
transform 1 0 81464 0 1 75213
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3190
timestamp 1649977179
transform 1 0 78608 0 1 75893
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3191
timestamp 1649977179
transform 1 0 78608 0 1 76573
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3192
timestamp 1649977179
transform 1 0 81464 0 1 76981
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3193
timestamp 1649977179
transform 1 0 81328 0 1 76573
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3194
timestamp 1649977179
transform 1 0 81328 0 1 75893
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3195
timestamp 1649977179
transform 1 0 78880 0 1 73173
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3196
timestamp 1649977179
transform 1 0 78880 0 1 75077
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3197
timestamp 1649977179
transform 1 0 78880 0 1 75213
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3198
timestamp 1649977179
transform 1 0 83504 0 1 77117
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3199
timestamp 1649977179
transform 1 0 81056 0 1 77117
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3200
timestamp 1649977179
transform 1 0 78608 0 1 77117
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3201
timestamp 1649977179
transform 1 0 78880 0 1 76981
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3202
timestamp 1649977179
transform 1 0 83912 0 1 73173
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3203
timestamp 1649977179
transform 1 0 83912 0 1 75077
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3204
timestamp 1649977179
transform 1 0 83912 0 1 75213
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3205
timestamp 1649977179
transform 1 0 83912 0 1 76981
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3206
timestamp 1649977179
transform 1 0 71128 0 1 75893
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3207
timestamp 1649977179
transform 1 0 68816 0 1 76573
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3208
timestamp 1649977179
transform 1 0 68816 0 1 75893
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3209
timestamp 1649977179
transform 1 0 68952 0 1 73173
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3210
timestamp 1649977179
transform 1 0 68952 0 1 75077
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3211
timestamp 1649977179
transform 1 0 76160 0 1 76573
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3212
timestamp 1649977179
transform 1 0 76160 0 1 75893
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3213
timestamp 1649977179
transform 1 0 68952 0 1 75213
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3214
timestamp 1649977179
transform 1 0 68952 0 1 77117
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3215
timestamp 1649977179
transform 1 0 73712 0 1 76573
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3216
timestamp 1649977179
transform 1 0 73712 0 1 75893
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3217
timestamp 1649977179
transform 1 0 75888 0 1 77117
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3218
timestamp 1649977179
transform 1 0 73576 0 1 77117
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3219
timestamp 1649977179
transform 1 0 70992 0 1 77117
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3220
timestamp 1649977179
transform 1 0 68544 0 1 77117
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3221
timestamp 1649977179
transform 1 0 71400 0 1 76573
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3222
timestamp 1649977179
transform 1 0 71400 0 1 75893
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3223
timestamp 1649977179
transform 1 0 71128 0 1 76573
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3224
timestamp 1649977179
transform 1 0 76432 0 1 73173
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3225
timestamp 1649977179
transform 1 0 76432 0 1 75077
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3226
timestamp 1649977179
transform 1 0 76432 0 1 75213
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3227
timestamp 1649977179
transform 1 0 76432 0 1 76981
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3228
timestamp 1649977179
transform 1 0 73984 0 1 73173
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3229
timestamp 1649977179
transform 1 0 73984 0 1 75077
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3230
timestamp 1649977179
transform 1 0 73848 0 1 75213
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3231
timestamp 1649977179
transform 1 0 73848 0 1 76981
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3232
timestamp 1649977179
transform 1 0 71400 0 1 73173
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3233
timestamp 1649977179
transform 1 0 71400 0 1 75077
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3234
timestamp 1649977179
transform 1 0 71264 0 1 75213
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3235
timestamp 1649977179
transform 1 0 71400 0 1 76981
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3236
timestamp 1649977179
transform 1 0 76160 0 1 82013
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3237
timestamp 1649977179
transform 1 0 76160 0 1 81469
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3238
timestamp 1649977179
transform 1 0 74392 0 1 82013
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3239
timestamp 1649977179
transform 1 0 74392 0 1 81469
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3240
timestamp 1649977179
transform 1 0 72624 0 1 82013
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3241
timestamp 1649977179
transform 1 0 72624 0 1 81469
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3242
timestamp 1649977179
transform 1 0 70856 0 1 82013
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3243
timestamp 1649977179
transform 1 0 70856 0 1 81469
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3244
timestamp 1649977179
transform 1 0 69224 0 1 82013
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3245
timestamp 1649977179
transform 1 0 69224 0 1 81469
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3246
timestamp 1649977179
transform 1 0 84456 0 1 82013
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3247
timestamp 1649977179
transform 1 0 84456 0 1 81469
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3248
timestamp 1649977179
transform 1 0 82688 0 1 82013
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3249
timestamp 1649977179
transform 1 0 82688 0 1 81469
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3250
timestamp 1649977179
transform 1 0 81328 0 1 82013
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3251
timestamp 1649977179
transform 1 0 81328 0 1 81469
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3252
timestamp 1649977179
transform 1 0 79424 0 1 82013
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3253
timestamp 1649977179
transform 1 0 77656 0 1 81469
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3254
timestamp 1649977179
transform 1 0 79424 0 1 81469
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3255
timestamp 1649977179
transform 1 0 77656 0 1 82013
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3256
timestamp 1649977179
transform 1 0 98600 0 1 76573
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3257
timestamp 1649977179
transform 1 0 101184 0 1 76573
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3258
timestamp 1649977179
transform 1 0 101184 0 1 75893
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3259
timestamp 1649977179
transform 1 0 96152 0 1 76573
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3260
timestamp 1649977179
transform 1 0 96152 0 1 75893
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3261
timestamp 1649977179
transform 1 0 98736 0 1 76573
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3262
timestamp 1649977179
transform 1 0 98736 0 1 75893
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3263
timestamp 1649977179
transform 1 0 101048 0 1 77117
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3264
timestamp 1649977179
transform 1 0 98464 0 1 77117
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3265
timestamp 1649977179
transform 1 0 96016 0 1 77117
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3266
timestamp 1649977179
transform 1 0 93840 0 1 76573
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3267
timestamp 1649977179
transform 1 0 93840 0 1 75893
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3268
timestamp 1649977179
transform 1 0 98600 0 1 75893
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3269
timestamp 1649977179
transform 1 0 101456 0 1 73173
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3270
timestamp 1649977179
transform 1 0 101456 0 1 75077
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3271
timestamp 1649977179
transform 1 0 101320 0 1 75213
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3272
timestamp 1649977179
transform 1 0 101320 0 1 76981
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3273
timestamp 1649977179
transform 1 0 98872 0 1 73173
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3274
timestamp 1649977179
transform 1 0 98872 0 1 75077
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3275
timestamp 1649977179
transform 1 0 98872 0 1 75213
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3276
timestamp 1649977179
transform 1 0 98872 0 1 76981
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3277
timestamp 1649977179
transform 1 0 96424 0 1 73173
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3278
timestamp 1649977179
transform 1 0 96424 0 1 75077
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3279
timestamp 1649977179
transform 1 0 96288 0 1 75213
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3280
timestamp 1649977179
transform 1 0 96288 0 1 76981
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3281
timestamp 1649977179
transform 1 0 93840 0 1 76981
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3282
timestamp 1649977179
transform 1 0 88808 0 1 76573
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3283
timestamp 1649977179
transform 1 0 88808 0 1 75893
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3284
timestamp 1649977179
transform 1 0 93568 0 1 75893
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3285
timestamp 1649977179
transform 1 0 93568 0 1 76573
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3286
timestamp 1649977179
transform 1 0 91392 0 1 76573
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3287
timestamp 1649977179
transform 1 0 91392 0 1 75893
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3288
timestamp 1649977179
transform 1 0 86360 0 1 76573
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3289
timestamp 1649977179
transform 1 0 86360 0 1 75893
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3290
timestamp 1649977179
transform 1 0 88536 0 1 76573
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3291
timestamp 1649977179
transform 1 0 93568 0 1 77117
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3292
timestamp 1649977179
transform 1 0 90984 0 1 77117
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3293
timestamp 1649977179
transform 1 0 88400 0 1 77117
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3294
timestamp 1649977179
transform 1 0 85952 0 1 77117
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3295
timestamp 1649977179
transform 1 0 93704 0 1 75213
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3296
timestamp 1649977179
transform 1 0 93704 0 1 75077
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3297
timestamp 1649977179
transform 1 0 93704 0 1 73173
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3298
timestamp 1649977179
transform 1 0 91392 0 1 73173
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3299
timestamp 1649977179
transform 1 0 91392 0 1 75077
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3300
timestamp 1649977179
transform 1 0 91256 0 1 75213
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3301
timestamp 1649977179
transform 1 0 91256 0 1 77117
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3302
timestamp 1649977179
transform 1 0 88944 0 1 73173
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3303
timestamp 1649977179
transform 1 0 88944 0 1 75077
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3304
timestamp 1649977179
transform 1 0 88944 0 1 75213
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3305
timestamp 1649977179
transform 1 0 88944 0 1 76981
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3306
timestamp 1649977179
transform 1 0 86496 0 1 73173
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3307
timestamp 1649977179
transform 1 0 86496 0 1 75077
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3308
timestamp 1649977179
transform 1 0 86224 0 1 75213
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3309
timestamp 1649977179
transform 1 0 86360 0 1 76981
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3310
timestamp 1649977179
transform 1 0 88536 0 1 75893
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3311
timestamp 1649977179
transform 1 0 92888 0 1 82013
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3312
timestamp 1649977179
transform 1 0 92888 0 1 81469
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3313
timestamp 1649977179
transform 1 0 91120 0 1 82013
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3314
timestamp 1649977179
transform 1 0 91120 0 1 81469
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3315
timestamp 1649977179
transform 1 0 89352 0 1 82013
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3316
timestamp 1649977179
transform 1 0 89352 0 1 81469
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3317
timestamp 1649977179
transform 1 0 87720 0 1 82013
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3318
timestamp 1649977179
transform 1 0 87720 0 1 81469
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3319
timestamp 1649977179
transform 1 0 86224 0 1 82013
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3320
timestamp 1649977179
transform 1 0 86224 0 1 81469
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3321
timestamp 1649977179
transform 1 0 94384 0 1 81469
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3322
timestamp 1649977179
transform 1 0 101320 0 1 82013
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3323
timestamp 1649977179
transform 1 0 101320 0 1 81469
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3324
timestamp 1649977179
transform 1 0 99688 0 1 82013
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3325
timestamp 1649977179
transform 1 0 99688 0 1 81469
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3326
timestamp 1649977179
transform 1 0 97920 0 1 82013
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3327
timestamp 1649977179
transform 1 0 97920 0 1 81469
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3328
timestamp 1649977179
transform 1 0 96288 0 1 82013
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3329
timestamp 1649977179
transform 1 0 96288 0 1 81469
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3330
timestamp 1649977179
transform 1 0 94384 0 1 82013
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3331
timestamp 1649977179
transform 1 0 135320 0 1 62429
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3332
timestamp 1649977179
transform 1 0 136000 0 1 64469
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3333
timestamp 1649977179
transform 1 0 133416 0 1 64197
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3334
timestamp 1649977179
transform 1 0 133144 0 1 67053
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3335
timestamp 1649977179
transform 1 0 132600 0 1 66917
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3336
timestamp 1649977179
transform 1 0 132600 0 1 64333
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3337
timestamp 1649977179
transform 1 0 135320 0 1 65829
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3338
timestamp 1649977179
transform 1 0 135320 0 1 64061
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3339
timestamp 1649977179
transform 1 0 122400 0 1 71405
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3340
timestamp 1649977179
transform 1 0 135320 0 1 70861
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3341
timestamp 1649977179
transform 1 0 133144 0 1 69773
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3342
timestamp 1649977179
transform 1 0 134776 0 1 70997
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3343
timestamp 1649977179
transform 1 0 134776 0 1 71269
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3344
timestamp 1649977179
transform 1 0 134776 0 1 69093
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3345
timestamp 1649977179
transform 1 0 134776 0 1 68549
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3346
timestamp 1649977179
transform 1 0 135320 0 1 69365
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3347
timestamp 1649977179
transform 1 0 134087 0 1 72293
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3348
timestamp 1649977179
transform 1 0 135320 0 1 72493
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3349
timestamp 1649977179
transform 1 0 135320 0 1 67597
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3350
timestamp 1649977179
transform 1 0 114376 0 1 65557
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3351
timestamp 1649977179
transform 1 0 114376 0 1 65965
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3352
timestamp 1649977179
transform 1 0 114376 0 1 65693
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3353
timestamp 1649977179
transform 1 0 115328 0 1 66101
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3354
timestamp 1649977179
transform 1 0 115328 0 1 66373
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3355
timestamp 1649977179
transform 1 0 115056 0 1 66101
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3356
timestamp 1649977179
transform 1 0 115056 0 1 66373
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3357
timestamp 1649977179
transform 1 0 115056 0 1 62565
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3358
timestamp 1649977179
transform 1 0 115056 0 1 62837
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3359
timestamp 1649977179
transform 1 0 115056 0 1 65149
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3360
timestamp 1649977179
transform 1 0 115056 0 1 64877
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3361
timestamp 1649977179
transform 1 0 115328 0 1 64061
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3362
timestamp 1649977179
transform 1 0 115328 0 1 64333
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3363
timestamp 1649977179
transform 1 0 114240 0 1 66101
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3364
timestamp 1649977179
transform 1 0 114240 0 1 66373
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3365
timestamp 1649977179
transform 1 0 115872 0 1 65285
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3366
timestamp 1649977179
transform 1 0 115872 0 1 65557
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3367
timestamp 1649977179
transform 1 0 114376 0 1 66781
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3368
timestamp 1649977179
transform 1 0 116008 0 1 67325
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3369
timestamp 1649977179
transform 1 0 114376 0 1 66509
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3370
timestamp 1649977179
transform 1 0 115600 0 1 66781
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3371
timestamp 1649977179
transform 1 0 115192 0 1 62429
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3372
timestamp 1649977179
transform 1 0 115600 0 1 66509
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3373
timestamp 1649977179
transform 1 0 116008 0 1 65693
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3374
timestamp 1649977179
transform 1 0 116008 0 1 65965
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3375
timestamp 1649977179
transform 1 0 116008 0 1 63789
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3376
timestamp 1649977179
transform 1 0 116008 0 1 64061
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3377
timestamp 1649977179
transform 1 0 115872 0 1 63653
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3378
timestamp 1649977179
transform 1 0 115872 0 1 63381
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3379
timestamp 1649977179
transform 1 0 116008 0 1 66101
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3380
timestamp 1649977179
transform 1 0 116008 0 1 66373
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3381
timestamp 1649977179
transform 1 0 115872 0 1 67189
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3382
timestamp 1649977179
transform 1 0 115872 0 1 66917
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3383
timestamp 1649977179
transform 1 0 115872 0 1 66509
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3384
timestamp 1649977179
transform 1 0 115872 0 1 66781
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3385
timestamp 1649977179
transform 1 0 116008 0 1 63245
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3386
timestamp 1649977179
transform 1 0 116008 0 1 62973
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3387
timestamp 1649977179
transform 1 0 115600 0 1 65693
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3388
timestamp 1649977179
transform 1 0 114240 0 1 64877
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3389
timestamp 1649977179
transform 1 0 114240 0 1 65149
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3390
timestamp 1649977179
transform 1 0 115872 0 1 62429
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3391
timestamp 1649977179
transform 1 0 115872 0 1 62837
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3392
timestamp 1649977179
transform 1 0 115872 0 1 62565
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3393
timestamp 1649977179
transform 1 0 114240 0 1 63245
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3394
timestamp 1649977179
transform 1 0 114240 0 1 62973
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3395
timestamp 1649977179
transform 1 0 115328 0 1 65285
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3396
timestamp 1649977179
transform 1 0 115328 0 1 65557
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3397
timestamp 1649977179
transform 1 0 114648 0 1 64469
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3398
timestamp 1649977179
transform 1 0 114648 0 1 64741
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3399
timestamp 1649977179
transform 1 0 114784 0 1 62429
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3400
timestamp 1649977179
transform 1 0 114648 0 1 62565
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3401
timestamp 1649977179
transform 1 0 114648 0 1 62837
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3402
timestamp 1649977179
transform 1 0 114240 0 1 62565
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3403
timestamp 1649977179
transform 1 0 114240 0 1 62837
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3404
timestamp 1649977179
transform 1 0 115600 0 1 65965
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3405
timestamp 1649977179
transform 1 0 115464 0 1 62837
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3406
timestamp 1649977179
transform 1 0 114784 0 1 62973
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3407
timestamp 1649977179
transform 1 0 114784 0 1 63245
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3408
timestamp 1649977179
transform 1 0 114376 0 1 62429
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3409
timestamp 1649977179
transform 1 0 115464 0 1 62565
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3410
timestamp 1649977179
transform 1 0 115464 0 1 65149
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3411
timestamp 1649977179
transform 1 0 115600 0 1 67325
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3412
timestamp 1649977179
transform 1 0 114648 0 1 65693
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3413
timestamp 1649977179
transform 1 0 114648 0 1 65965
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3414
timestamp 1649977179
transform 1 0 114784 0 1 66781
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3415
timestamp 1649977179
transform 1 0 114784 0 1 66509
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3416
timestamp 1649977179
transform 1 0 114648 0 1 66101
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3417
timestamp 1649977179
transform 1 0 114648 0 1 66373
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3418
timestamp 1649977179
transform 1 0 114648 0 1 64877
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3419
timestamp 1649977179
transform 1 0 114648 0 1 65149
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3420
timestamp 1649977179
transform 1 0 114648 0 1 65557
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3421
timestamp 1649977179
transform 1 0 114648 0 1 65285
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3422
timestamp 1649977179
transform 1 0 114648 0 1 66917
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3423
timestamp 1649977179
transform 1 0 114648 0 1 67189
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3424
timestamp 1649977179
transform 1 0 115192 0 1 65285
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3425
timestamp 1649977179
transform 1 0 115464 0 1 64877
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3426
timestamp 1649977179
transform 1 0 114376 0 1 64741
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3427
timestamp 1649977179
transform 1 0 114376 0 1 64469
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3428
timestamp 1649977179
transform 1 0 114376 0 1 67189
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3429
timestamp 1649977179
transform 1 0 114376 0 1 66917
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3430
timestamp 1649977179
transform 1 0 115464 0 1 63653
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3431
timestamp 1649977179
transform 1 0 115192 0 1 65557
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3432
timestamp 1649977179
transform 1 0 115464 0 1 63381
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3433
timestamp 1649977179
transform 1 0 114376 0 1 65285
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3434
timestamp 1649977179
transform 1 0 109344 0 1 67325
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3435
timestamp 1649977179
transform 1 0 109208 0 1 63925
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3436
timestamp 1649977179
transform 1 0 109208 0 1 63517
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3437
timestamp 1649977179
transform 1 0 109344 0 1 63789
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3438
timestamp 1649977179
transform 1 0 109344 0 1 63517
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3439
timestamp 1649977179
transform 1 0 109344 0 1 62565
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3440
timestamp 1649977179
transform 1 0 109480 0 1 63925
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3441
timestamp 1649977179
transform 1 0 109480 0 1 64197
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3442
timestamp 1649977179
transform 1 0 109480 0 1 67325
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3443
timestamp 1649977179
transform 1 0 109480 0 1 67053
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3444
timestamp 1649977179
transform 1 0 109344 0 1 64333
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3445
timestamp 1649977179
transform 1 0 109344 0 1 64741
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3446
timestamp 1649977179
transform 1 0 109480 0 1 67869
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3447
timestamp 1649977179
transform 1 0 109480 0 1 68141
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3448
timestamp 1649977179
transform 1 0 109616 0 1 70861
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3449
timestamp 1649977179
transform 1 0 106080 0 1 70997
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3450
timestamp 1649977179
transform 1 0 106080 0 1 71405
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3451
timestamp 1649977179
transform 1 0 110704 0 1 70589
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3452
timestamp 1649977179
transform 1 0 110704 0 1 70997
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3453
timestamp 1649977179
transform 1 0 108528 0 1 70997
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3454
timestamp 1649977179
transform 1 0 108528 0 1 71405
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3455
timestamp 1649977179
transform 1 0 104312 0 1 70997
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3456
timestamp 1649977179
transform 1 0 103632 0 1 71405
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3457
timestamp 1649977179
transform 1 0 107304 0 1 70997
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3458
timestamp 1649977179
transform 1 0 107304 0 1 71405
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3459
timestamp 1649977179
transform 1 0 105536 0 1 71405
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3460
timestamp 1649977179
transform 1 0 102408 0 1 70997
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3461
timestamp 1649977179
transform 1 0 103632 0 1 70997
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3462
timestamp 1649977179
transform 1 0 103088 0 1 71405
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3463
timestamp 1649977179
transform 1 0 105536 0 1 70997
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3464
timestamp 1649977179
transform 1 0 104856 0 1 70997
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3465
timestamp 1649977179
transform 1 0 104856 0 1 71405
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3466
timestamp 1649977179
transform 1 0 103088 0 1 70997
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3467
timestamp 1649977179
transform 1 0 102408 0 1 71405
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3468
timestamp 1649977179
transform 1 0 104312 0 1 71405
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3469
timestamp 1649977179
transform 1 0 109344 0 1 67733
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3470
timestamp 1649977179
transform 1 0 115328 0 1 69909
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3471
timestamp 1649977179
transform 1 0 115328 0 1 68277
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3472
timestamp 1649977179
transform 1 0 115328 0 1 68005
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3473
timestamp 1649977179
transform 1 0 115056 0 1 69501
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3474
timestamp 1649977179
transform 1 0 115056 0 1 69229
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3475
timestamp 1649977179
transform 1 0 116008 0 1 67597
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3476
timestamp 1649977179
transform 1 0 116008 0 1 68821
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3477
timestamp 1649977179
transform 1 0 116008 0 1 68549
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3478
timestamp 1649977179
transform 1 0 116008 0 1 69501
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3479
timestamp 1649977179
transform 1 0 116008 0 1 69229
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3480
timestamp 1649977179
transform 1 0 115192 0 1 69093
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3481
timestamp 1649977179
transform 1 0 115872 0 1 67733
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3482
timestamp 1649977179
transform 1 0 115872 0 1 68005
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3483
timestamp 1649977179
transform 1 0 115872 0 1 70045
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3484
timestamp 1649977179
transform 1 0 115192 0 1 68821
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3485
timestamp 1649977179
transform 1 0 114648 0 1 68685
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3486
timestamp 1649977179
transform 1 0 114648 0 1 68413
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3487
timestamp 1649977179
transform 1 0 114784 0 1 68821
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3488
timestamp 1649977179
transform 1 0 114784 0 1 69093
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3489
timestamp 1649977179
transform 1 0 114648 0 1 69909
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3490
timestamp 1649977179
transform 1 0 114648 0 1 69637
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3491
timestamp 1649977179
transform 1 0 114648 0 1 69229
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3492
timestamp 1649977179
transform 1 0 114648 0 1 69501
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3493
timestamp 1649977179
transform 1 0 114376 0 1 68413
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3494
timestamp 1649977179
transform 1 0 114376 0 1 68685
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3495
timestamp 1649977179
transform 1 0 114240 0 1 69501
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3496
timestamp 1649977179
transform 1 0 114240 0 1 69229
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3497
timestamp 1649977179
transform 1 0 114376 0 1 68821
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3498
timestamp 1649977179
transform 1 0 114376 0 1 69093
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3499
timestamp 1649977179
transform 1 0 114376 0 1 69637
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3500
timestamp 1649977179
transform 1 0 114376 0 1 69909
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3501
timestamp 1649977179
transform 1 0 115328 0 1 70589
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3502
timestamp 1649977179
transform 1 0 114240 0 1 70045
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3503
timestamp 1649977179
transform 1 0 114240 0 1 70453
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3504
timestamp 1649977179
transform 1 0 115600 0 1 67597
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3505
timestamp 1649977179
transform 1 0 115464 0 1 69909
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3506
timestamp 1649977179
transform 1 0 115464 0 1 69637
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3507
timestamp 1649977179
transform 1 0 115600 0 1 69501
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3508
timestamp 1649977179
transform 1 0 115600 0 1 69229
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3509
timestamp 1649977179
transform 1 0 115328 0 1 69637
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3510
timestamp 1649977179
transform 1 0 115872 0 1 72901
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3511
timestamp 1649977179
transform 1 0 115464 0 1 73037
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3512
timestamp 1649977179
transform 1 0 115464 0 1 75621
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3513
timestamp 1649977179
transform 1 0 115328 0 1 74397
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3514
timestamp 1649977179
transform 1 0 118048 0 1 77253
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3515
timestamp 1649977179
transform 1 0 116552 0 1 75893
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3516
timestamp 1649977179
transform 1 0 115328 0 1 77117
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3517
timestamp 1649977179
transform 1 0 115328 0 1 74261
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3518
timestamp 1649977179
transform 1 0 106352 0 1 76981
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3519
timestamp 1649977179
transform 1 0 103904 0 1 73173
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3520
timestamp 1649977179
transform 1 0 103904 0 1 75077
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3521
timestamp 1649977179
transform 1 0 103904 0 1 75213
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3522
timestamp 1649977179
transform 1 0 103904 0 1 77117
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3523
timestamp 1649977179
transform 1 0 106216 0 1 76573
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3524
timestamp 1649977179
transform 1 0 106216 0 1 75893
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3525
timestamp 1649977179
transform 1 0 106080 0 1 77117
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3526
timestamp 1649977179
transform 1 0 103768 0 1 76573
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3527
timestamp 1649977179
transform 1 0 103768 0 1 75893
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3528
timestamp 1649977179
transform 1 0 103360 0 1 77117
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3529
timestamp 1649977179
transform 1 0 109616 0 1 73037
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3530
timestamp 1649977179
transform 1 0 106352 0 1 73173
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3531
timestamp 1649977179
transform 1 0 106352 0 1 75077
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3532
timestamp 1649977179
transform 1 0 106352 0 1 75213
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3533
timestamp 1649977179
transform 1 0 109616 0 1 82013
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3534
timestamp 1649977179
transform 1 0 109616 0 1 81469
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3535
timestamp 1649977179
transform 1 0 107848 0 1 82013
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3536
timestamp 1649977179
transform 1 0 107848 0 1 81469
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3537
timestamp 1649977179
transform 1 0 106352 0 1 82013
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3538
timestamp 1649977179
transform 1 0 106352 0 1 81469
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3539
timestamp 1649977179
transform 1 0 104584 0 1 82013
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3540
timestamp 1649977179
transform 1 0 104584 0 1 81469
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3541
timestamp 1649977179
transform 1 0 102952 0 1 82013
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3542
timestamp 1649977179
transform 1 0 102952 0 1 81469
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3543
timestamp 1649977179
transform 1 0 118048 0 1 82693
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3544
timestamp 1649977179
transform 1 0 118048 0 1 80789
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3545
timestamp 1649977179
transform 1 0 117912 0 1 80653
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3546
timestamp 1649977179
transform 1 0 117912 0 1 78613
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3547
timestamp 1649977179
transform 1 0 116552 0 1 78477
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3548
timestamp 1649977179
transform 1 0 117912 0 1 82013
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3549
timestamp 1649977179
transform 1 0 117912 0 1 81469
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3550
timestamp 1649977179
transform 1 0 118184 0 1 79429
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3551
timestamp 1649977179
transform 1 0 118184 0 1 81333
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3552
timestamp 1649977179
transform 1 0 118048 0 1 79293
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3553
timestamp 1649977179
transform 1 0 116416 0 1 82013
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3554
timestamp 1649977179
transform 1 0 116416 0 1 81469
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3555
timestamp 1649977179
transform 1 0 114648 0 1 82013
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3556
timestamp 1649977179
transform 1 0 114648 0 1 81469
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3557
timestamp 1649977179
transform 1 0 112880 0 1 82013
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3558
timestamp 1649977179
transform 1 0 112880 0 1 81469
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3559
timestamp 1649977179
transform 1 0 111384 0 1 82013
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3560
timestamp 1649977179
transform 1 0 111384 0 1 81469
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3561
timestamp 1649977179
transform 1 0 118456 0 1 80245
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3562
timestamp 1649977179
transform 1 0 136000 0 1 72765
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3563
timestamp 1649977179
transform 1 0 135320 0 1 74125
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3564
timestamp 1649977179
transform 1 0 135320 0 1 77661
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3565
timestamp 1649977179
transform 1 0 135320 0 1 76029
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3566
timestamp 1649977179
transform 1 0 134776 0 1 77661
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3567
timestamp 1649977179
transform 1 0 122264 0 1 75621
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3568
timestamp 1649977179
transform 1 0 122400 0 1 76981
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3569
timestamp 1649977179
transform 1 0 122400 0 1 73989
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3570
timestamp 1649977179
transform 1 0 122400 0 1 76845
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3571
timestamp 1649977179
transform 1 0 122400 0 1 74261
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3572
timestamp 1649977179
transform 1 0 122264 0 1 75485
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3573
timestamp 1649977179
transform 1 0 122264 0 1 72765
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3574
timestamp 1649977179
transform 1 0 122400 0 1 79701
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3575
timestamp 1649977179
transform 1 0 122264 0 1 79837
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3576
timestamp 1649977179
transform 1 0 122264 0 1 80653
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3577
timestamp 1649977179
transform 1 0 126344 0 1 82013
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3578
timestamp 1649977179
transform 1 0 126344 0 1 81469
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3579
timestamp 1649977179
transform 1 0 124712 0 1 82013
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3580
timestamp 1649977179
transform 1 0 124712 0 1 81469
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3581
timestamp 1649977179
transform 1 0 123216 0 1 82013
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3582
timestamp 1649977179
transform 1 0 123216 0 1 81469
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3583
timestamp 1649977179
transform 1 0 122944 0 1 81333
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3584
timestamp 1649977179
transform 1 0 122944 0 1 78477
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3585
timestamp 1649977179
transform 1 0 122264 0 1 78341
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3586
timestamp 1649977179
transform 1 0 121448 0 1 82013
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3587
timestamp 1649977179
transform 1 0 121448 0 1 81469
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3588
timestamp 1649977179
transform 1 0 119544 0 1 82013
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3589
timestamp 1649977179
transform 1 0 119544 0 1 81469
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3590
timestamp 1649977179
transform 1 0 119680 0 1 80245
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3591
timestamp 1649977179
transform 1 0 136000 0 1 79837
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3592
timestamp 1649977179
transform 1 0 135320 0 1 79429
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3593
timestamp 1649977179
transform 1 0 134776 0 1 78341
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3594
timestamp 1649977179
transform 1 0 130832 0 1 79157
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3595
timestamp 1649977179
transform 1 0 131376 0 1 82013
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3596
timestamp 1649977179
transform 1 0 131376 0 1 81469
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3597
timestamp 1649977179
transform 1 0 129880 0 1 82013
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3598
timestamp 1649977179
transform 1 0 129880 0 1 81469
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3599
timestamp 1649977179
transform 1 0 128112 0 1 82013
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3600
timestamp 1649977179
transform 1 0 128112 0 1 81469
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3601
timestamp 1649977179
transform 1 0 135320 0 1 80925
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3602
timestamp 1649977179
transform 1 0 133144 0 1 82013
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3603
timestamp 1649977179
transform 1 0 133144 0 1 81469
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3604
timestamp 1649977179
transform 1 0 109344 0 1 62293
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3605
timestamp 1649977179
transform 1 0 115872 0 1 41621
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3606
timestamp 1649977179
transform 1 0 114784 0 1 41621
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3607
timestamp 1649977179
transform 1 0 22032 0 1 41621
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3608
timestamp 1649977179
transform 1 0 20808 0 1 41621
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3609
timestamp 1649977179
transform 1 0 115328 0 1 41621
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3610
timestamp 1649977179
transform 1 0 115192 0 1 41621
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3611
timestamp 1649977179
transform 1 0 114376 0 1 41621
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3612
timestamp 1649977179
transform 1 0 22440 0 1 41621
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3613
timestamp 1649977179
transform 1 0 21624 0 1 41621
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3614
timestamp 1649977179
transform 1 0 21216 0 1 41621
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3615
timestamp 1649977179
transform 1 0 68272 0 1 13061
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_38  sky130_sram_2kbyte_1rw1r_32x512_8_contact_38_0
timestamp 1649977179
transform 1 0 134776 0 1 1628
box 0 0 192 192
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_38  sky130_sram_2kbyte_1rw1r_32x512_8_contact_38_1
timestamp 1649977179
transform 1 0 1726 0 1 1628
box 0 0 192 192
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_38  sky130_sram_2kbyte_1rw1r_32x512_8_contact_38_2
timestamp 1649977179
transform 1 0 1726 0 1 81377
box 0 0 192 192
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_38  sky130_sram_2kbyte_1rw1r_32x512_8_contact_38_3
timestamp 1649977179
transform 1 0 134776 0 1 81377
box 0 0 192 192
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_39  sky130_sram_2kbyte_1rw1r_32x512_8_contact_39_0
timestamp 1649977179
transform 1 0 136000 0 1 413
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_39  sky130_sram_2kbyte_1rw1r_32x512_8_contact_39_1
timestamp 1649977179
transform 1 0 136272 0 1 413
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_39  sky130_sram_2kbyte_1rw1r_32x512_8_contact_39_2
timestamp 1649977179
transform 1 0 136136 0 1 549
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_39  sky130_sram_2kbyte_1rw1r_32x512_8_contact_39_3
timestamp 1649977179
transform 1 0 135592 0 1 1229
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_39  sky130_sram_2kbyte_1rw1r_32x512_8_contact_39_4
timestamp 1649977179
transform 1 0 135320 0 1 957
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_39  sky130_sram_2kbyte_1rw1r_32x512_8_contact_39_5
timestamp 1649977179
transform 1 0 135456 0 1 1229
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_39  sky130_sram_2kbyte_1rw1r_32x512_8_contact_39_6
timestamp 1649977179
transform 1 0 135592 0 1 1093
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_39  sky130_sram_2kbyte_1rw1r_32x512_8_contact_39_7
timestamp 1649977179
transform 1 0 135320 0 1 1229
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_39  sky130_sram_2kbyte_1rw1r_32x512_8_contact_39_8
timestamp 1649977179
transform 1 0 135456 0 1 957
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_39  sky130_sram_2kbyte_1rw1r_32x512_8_contact_39_9
timestamp 1649977179
transform 1 0 136272 0 1 277
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_39  sky130_sram_2kbyte_1rw1r_32x512_8_contact_39_10
timestamp 1649977179
transform 1 0 136000 0 1 277
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_39  sky130_sram_2kbyte_1rw1r_32x512_8_contact_39_11
timestamp 1649977179
transform 1 0 136272 0 1 549
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_39  sky130_sram_2kbyte_1rw1r_32x512_8_contact_39_12
timestamp 1649977179
transform 1 0 135456 0 1 1093
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_39  sky130_sram_2kbyte_1rw1r_32x512_8_contact_39_13
timestamp 1649977179
transform 1 0 136000 0 1 549
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_39  sky130_sram_2kbyte_1rw1r_32x512_8_contact_39_14
timestamp 1649977179
transform 1 0 135592 0 1 957
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_39  sky130_sram_2kbyte_1rw1r_32x512_8_contact_39_15
timestamp 1649977179
transform 1 0 135320 0 1 1093
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_39  sky130_sram_2kbyte_1rw1r_32x512_8_contact_39_16
timestamp 1649977179
transform 1 0 136136 0 1 277
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_39  sky130_sram_2kbyte_1rw1r_32x512_8_contact_39_17
timestamp 1649977179
transform 1 0 136136 0 1 413
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_39  sky130_sram_2kbyte_1rw1r_32x512_8_contact_39_18
timestamp 1649977179
transform 1 0 408 0 1 277
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_39  sky130_sram_2kbyte_1rw1r_32x512_8_contact_39_19
timestamp 1649977179
transform 1 0 544 0 1 277
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_39  sky130_sram_2kbyte_1rw1r_32x512_8_contact_39_20
timestamp 1649977179
transform 1 0 408 0 1 413
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_39  sky130_sram_2kbyte_1rw1r_32x512_8_contact_39_21
timestamp 1649977179
transform 1 0 544 0 1 549
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_39  sky130_sram_2kbyte_1rw1r_32x512_8_contact_39_22
timestamp 1649977179
transform 1 0 1224 0 1 1093
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_39  sky130_sram_2kbyte_1rw1r_32x512_8_contact_39_23
timestamp 1649977179
transform 1 0 952 0 1 1093
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_39  sky130_sram_2kbyte_1rw1r_32x512_8_contact_39_24
timestamp 1649977179
transform 1 0 952 0 1 1229
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_39  sky130_sram_2kbyte_1rw1r_32x512_8_contact_39_25
timestamp 1649977179
transform 1 0 1088 0 1 1229
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_39  sky130_sram_2kbyte_1rw1r_32x512_8_contact_39_26
timestamp 1649977179
transform 1 0 1088 0 1 1093
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_39  sky130_sram_2kbyte_1rw1r_32x512_8_contact_39_27
timestamp 1649977179
transform 1 0 408 0 1 549
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_39  sky130_sram_2kbyte_1rw1r_32x512_8_contact_39_28
timestamp 1649977179
transform 1 0 272 0 1 277
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_39  sky130_sram_2kbyte_1rw1r_32x512_8_contact_39_29
timestamp 1649977179
transform 1 0 1088 0 1 957
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_39  sky130_sram_2kbyte_1rw1r_32x512_8_contact_39_30
timestamp 1649977179
transform 1 0 1224 0 1 1229
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_39  sky130_sram_2kbyte_1rw1r_32x512_8_contact_39_31
timestamp 1649977179
transform 1 0 544 0 1 413
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_39  sky130_sram_2kbyte_1rw1r_32x512_8_contact_39_32
timestamp 1649977179
transform 1 0 1224 0 1 957
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_39  sky130_sram_2kbyte_1rw1r_32x512_8_contact_39_33
timestamp 1649977179
transform 1 0 952 0 1 957
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_39  sky130_sram_2kbyte_1rw1r_32x512_8_contact_39_34
timestamp 1649977179
transform 1 0 272 0 1 413
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_39  sky130_sram_2kbyte_1rw1r_32x512_8_contact_39_35
timestamp 1649977179
transform 1 0 272 0 1 549
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_39  sky130_sram_2kbyte_1rw1r_32x512_8_contact_39_36
timestamp 1649977179
transform 1 0 408 0 1 82829
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_39  sky130_sram_2kbyte_1rw1r_32x512_8_contact_39_37
timestamp 1649977179
transform 1 0 1224 0 1 82013
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_39  sky130_sram_2kbyte_1rw1r_32x512_8_contact_39_38
timestamp 1649977179
transform 1 0 272 0 1 82829
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_39  sky130_sram_2kbyte_1rw1r_32x512_8_contact_39_39
timestamp 1649977179
transform 1 0 544 0 1 82829
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_39  sky130_sram_2kbyte_1rw1r_32x512_8_contact_39_40
timestamp 1649977179
transform 1 0 1088 0 1 82285
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_39  sky130_sram_2kbyte_1rw1r_32x512_8_contact_39_41
timestamp 1649977179
transform 1 0 1224 0 1 82149
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_39  sky130_sram_2kbyte_1rw1r_32x512_8_contact_39_42
timestamp 1649977179
transform 1 0 952 0 1 82149
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_39  sky130_sram_2kbyte_1rw1r_32x512_8_contact_39_43
timestamp 1649977179
transform 1 0 952 0 1 82285
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_39  sky130_sram_2kbyte_1rw1r_32x512_8_contact_39_44
timestamp 1649977179
transform 1 0 272 0 1 82965
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_39  sky130_sram_2kbyte_1rw1r_32x512_8_contact_39_45
timestamp 1649977179
transform 1 0 544 0 1 82965
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_39  sky130_sram_2kbyte_1rw1r_32x512_8_contact_39_46
timestamp 1649977179
transform 1 0 1224 0 1 82285
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_39  sky130_sram_2kbyte_1rw1r_32x512_8_contact_39_47
timestamp 1649977179
transform 1 0 408 0 1 82693
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_39  sky130_sram_2kbyte_1rw1r_32x512_8_contact_39_48
timestamp 1649977179
transform 1 0 544 0 1 82693
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_39  sky130_sram_2kbyte_1rw1r_32x512_8_contact_39_49
timestamp 1649977179
transform 1 0 408 0 1 82965
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_39  sky130_sram_2kbyte_1rw1r_32x512_8_contact_39_50
timestamp 1649977179
transform 1 0 1088 0 1 82013
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_39  sky130_sram_2kbyte_1rw1r_32x512_8_contact_39_51
timestamp 1649977179
transform 1 0 952 0 1 82013
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_39  sky130_sram_2kbyte_1rw1r_32x512_8_contact_39_52
timestamp 1649977179
transform 1 0 272 0 1 82693
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_39  sky130_sram_2kbyte_1rw1r_32x512_8_contact_39_53
timestamp 1649977179
transform 1 0 1088 0 1 82149
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_39  sky130_sram_2kbyte_1rw1r_32x512_8_contact_39_54
timestamp 1649977179
transform 1 0 136000 0 1 82829
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_39  sky130_sram_2kbyte_1rw1r_32x512_8_contact_39_55
timestamp 1649977179
transform 1 0 136000 0 1 82693
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_39  sky130_sram_2kbyte_1rw1r_32x512_8_contact_39_56
timestamp 1649977179
transform 1 0 136272 0 1 82965
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_39  sky130_sram_2kbyte_1rw1r_32x512_8_contact_39_57
timestamp 1649977179
transform 1 0 136136 0 1 82829
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_39  sky130_sram_2kbyte_1rw1r_32x512_8_contact_39_58
timestamp 1649977179
transform 1 0 136000 0 1 82965
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_39  sky130_sram_2kbyte_1rw1r_32x512_8_contact_39_59
timestamp 1649977179
transform 1 0 136272 0 1 82693
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_39  sky130_sram_2kbyte_1rw1r_32x512_8_contact_39_60
timestamp 1649977179
transform 1 0 136272 0 1 82829
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_39  sky130_sram_2kbyte_1rw1r_32x512_8_contact_39_61
timestamp 1649977179
transform 1 0 136136 0 1 82965
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_39  sky130_sram_2kbyte_1rw1r_32x512_8_contact_39_62
timestamp 1649977179
transform 1 0 136136 0 1 82693
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_39  sky130_sram_2kbyte_1rw1r_32x512_8_contact_39_63
timestamp 1649977179
transform 1 0 135456 0 1 82285
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_39  sky130_sram_2kbyte_1rw1r_32x512_8_contact_39_64
timestamp 1649977179
transform 1 0 135592 0 1 82013
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_39  sky130_sram_2kbyte_1rw1r_32x512_8_contact_39_65
timestamp 1649977179
transform 1 0 135320 0 1 82149
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_39  sky130_sram_2kbyte_1rw1r_32x512_8_contact_39_66
timestamp 1649977179
transform 1 0 135456 0 1 82013
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_39  sky130_sram_2kbyte_1rw1r_32x512_8_contact_39_67
timestamp 1649977179
transform 1 0 135592 0 1 82285
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_39  sky130_sram_2kbyte_1rw1r_32x512_8_contact_39_68
timestamp 1649977179
transform 1 0 135320 0 1 82013
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_39  sky130_sram_2kbyte_1rw1r_32x512_8_contact_39_69
timestamp 1649977179
transform 1 0 135320 0 1 82285
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_39  sky130_sram_2kbyte_1rw1r_32x512_8_contact_39_70
timestamp 1649977179
transform 1 0 135456 0 1 82149
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_39  sky130_sram_2kbyte_1rw1r_32x512_8_contact_39_71
timestamp 1649977179
transform 1 0 135592 0 1 82149
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_control_logic_r  sky130_sram_2kbyte_1rw1r_32x512_8_control_logic_r_0
timestamp 1649977179
transform -1 0 134082 0 -1 79804
box -75 -49 11782 18431
use sky130_sram_2kbyte_1rw1r_32x512_8_control_logic_rw  sky130_sram_2kbyte_1rw1r_32x512_8_control_logic_rw_0
timestamp 1649977179
transform 1 0 2612 0 1 7620
box -75 -49 12082 18431
use sky130_sram_2kbyte_1rw1r_32x512_8_cr_3  sky130_sram_2kbyte_1rw1r_32x512_8_cr_3_0
timestamp 1649977179
transform 1 0 14862 0 1 9422
box 2083 -6379 5297 4372
use sky130_sram_2kbyte_1rw1r_32x512_8_cr_4  sky130_sram_2kbyte_1rw1r_32x512_8_cr_4_0
timestamp 1649977179
transform 1 0 14862 0 1 9422
box 4376 -6402 91393 1462
use sky130_sram_2kbyte_1rw1r_32x512_8_cr_5  sky130_sram_2kbyte_1rw1r_32x512_8_cr_5_0
timestamp 1649977179
transform 1 0 14862 0 1 9422
box 101765 67036 104019 70732
use sky130_sram_2kbyte_1rw1r_32x512_8_data_dff  sky130_sram_2kbyte_1rw1r_32x512_8_data_dff_0
timestamp 1649977179
transform 1 0 22870 0 1 2396
box -36 -49 37412 1467
use sky130_sram_2kbyte_1rw1r_32x512_8_row_addr_dff  sky130_sram_2kbyte_1rw1r_32x512_8_row_addr_dff_0
timestamp 1649977179
transform -1 0 123468 0 -1 19846
box -36 -49 1204 9951
use sky130_sram_2kbyte_1rw1r_32x512_8_row_addr_dff  sky130_sram_2kbyte_1rw1r_32x512_8_row_addr_dff_1
timestamp 1649977179
transform 1 0 13526 0 1 27746
box -36 -49 1204 9951
use sky130_sram_2kbyte_1rw1r_32x512_8_wmask_dff  sky130_sram_2kbyte_1rw1r_32x512_8_wmask_dff_0
timestamp 1649977179
transform 1 0 18198 0 1 2396
box -36 -49 4708 1467
<< labels >>
rlabel metal3 s 0 8024 212 8100 4 csb0
port 51 nsew default input
rlabel metal3 s 0 9928 212 10004 4 web0
port 53 nsew default input
rlabel metal3 s 0 8296 212 8372 4 clk0
port 54 nsew default input
rlabel metal3 s 0 28152 212 28228 4 addr0[2]
port 39 nsew default input
rlabel metal3 s 0 29920 212 29996 4 addr0[3]
port 38 nsew default input
rlabel metal3 s 0 31008 212 31084 4 addr0[4]
port 37 nsew default input
rlabel metal3 s 0 32776 212 32852 4 addr0[5]
port 36 nsew default input
rlabel metal3 s 0 33728 212 33804 4 addr0[6]
port 35 nsew default input
rlabel metal3 s 0 35904 212 35980 4 addr0[7]
port 34 nsew default input
rlabel metal3 s 0 36856 212 36932 4 addr0[8]
port 33 nsew default input
rlabel metal3 s 136408 79152 136620 79228 4 csb1
port 52 nsew default input
rlabel metal3 s 136408 19312 136620 19388 4 addr1[2]
port 48 nsew default input
rlabel metal3 s 136408 17680 136620 17756 4 addr1[3]
port 47 nsew default input
rlabel metal3 s 136408 16320 136620 16396 4 addr1[4]
port 46 nsew default input
rlabel metal3 s 136408 14824 136620 14900 4 addr1[5]
port 45 nsew default input
rlabel metal3 s 136408 13600 136620 13676 4 addr1[6]
port 44 nsew default input
rlabel metal3 s 952 82008 135668 82356 4 vccd1
port 124 nsew power bidirectional abutment
rlabel metal3 s 952 952 135668 1300 4 vccd1
port 124 nsew power bidirectional abutment
rlabel metal3 s 272 272 136348 620 4 vssd1
port 125 nsew ground bidirectional abutment
rlabel metal3 s 272 82688 136348 83036 4 vssd1
port 125 nsew ground bidirectional abutment
rlabel metal4 s 130832 83096 130908 83308 4 clk1
port 55 nsew default input
rlabel metal4 s 68544 83096 68620 83308 4 dout1[16]
port 107 nsew default output
rlabel metal4 s 70992 83096 71068 83308 4 dout1[17]
port 106 nsew default output
rlabel metal4 s 73576 83096 73652 83308 4 dout1[18]
port 105 nsew default output
rlabel metal4 s 75888 83096 75964 83308 4 dout1[19]
port 104 nsew default output
rlabel metal4 s 78608 83096 78684 83308 4 dout1[20]
port 103 nsew default output
rlabel metal4 s 81056 83096 81132 83308 4 dout1[21]
port 102 nsew default output
rlabel metal4 s 83504 83096 83580 83308 4 dout1[22]
port 101 nsew default output
rlabel metal4 s 85952 83096 86028 83308 4 dout1[23]
port 100 nsew default output
rlabel metal4 s 88400 83096 88476 83308 4 dout1[24]
port 99 nsew default output
rlabel metal4 s 90984 83096 91060 83308 4 dout1[25]
port 98 nsew default output
rlabel metal4 s 93568 83096 93644 83308 4 dout1[26]
port 97 nsew default output
rlabel metal4 s 96016 83096 96092 83308 4 dout1[27]
port 96 nsew default output
rlabel metal4 s 98464 83096 98540 83308 4 dout1[28]
port 95 nsew default output
rlabel metal4 s 101048 83096 101124 83308 4 dout1[29]
port 94 nsew default output
rlabel metal4 s 103360 83096 103436 83308 4 dout1[30]
port 93 nsew default output
rlabel metal4 s 106080 83096 106156 83308 4 dout1[31]
port 92 nsew default output
rlabel metal4 s 119680 83096 119756 83308 4 addr1[0]
port 50 nsew default input
rlabel metal4 s 118456 83096 118532 83308 4 addr1[1]
port 49 nsew default input
rlabel metal4 s 33456 83096 33532 83308 4 dout1[2]
port 121 nsew default output
rlabel metal4 s 36176 83096 36252 83308 4 dout1[3]
port 120 nsew default output
rlabel metal4 s 38488 83096 38564 83308 4 dout1[4]
port 119 nsew default output
rlabel metal4 s 41072 83096 41148 83308 4 dout1[5]
port 118 nsew default output
rlabel metal4 s 43520 83096 43596 83308 4 dout1[6]
port 117 nsew default output
rlabel metal4 s 46104 83096 46180 83308 4 dout1[7]
port 116 nsew default output
rlabel metal4 s 48552 83096 48628 83308 4 dout1[8]
port 115 nsew default output
rlabel metal4 s 51136 83096 51212 83308 4 dout1[9]
port 114 nsew default output
rlabel metal4 s 53584 83096 53660 83308 4 dout1[10]
port 113 nsew default output
rlabel metal4 s 56168 83096 56244 83308 4 dout1[11]
port 112 nsew default output
rlabel metal4 s 58480 83096 58556 83308 4 dout1[12]
port 111 nsew default output
rlabel metal4 s 60928 83096 61004 83308 4 dout1[13]
port 110 nsew default output
rlabel metal4 s 63648 83096 63724 83308 4 dout1[14]
port 109 nsew default output
rlabel metal4 s 66096 83096 66172 83308 4 dout1[15]
port 108 nsew default output
rlabel metal4 s 28696 83096 28772 83308 4 dout1[0]
port 123 nsew default output
rlabel metal4 s 31008 83096 31084 83308 4 dout1[1]
port 122 nsew default output
rlabel metal4 s 36040 0 36116 212 4 dout0[3]
port 88 nsew default output
rlabel metal4 s 38488 0 38564 212 4 dout0[4]
port 87 nsew default output
rlabel metal4 s 41072 0 41148 212 4 dout0[5]
port 86 nsew default output
rlabel metal4 s 43520 0 43596 212 4 dout0[6]
port 85 nsew default output
rlabel metal4 s 45968 0 46044 212 4 dout0[7]
port 84 nsew default output
rlabel metal4 s 48280 0 48356 212 4 dout0[8]
port 83 nsew default output
rlabel metal4 s 51000 0 51076 212 4 dout0[9]
port 82 nsew default output
rlabel metal4 s 53584 0 53660 212 4 dout0[10]
port 81 nsew default output
rlabel metal4 s 56032 0 56108 212 4 dout0[11]
port 80 nsew default output
rlabel metal4 s 58480 0 58556 212 4 dout0[12]
port 79 nsew default output
rlabel metal4 s 60928 0 61004 212 4 dout0[13]
port 78 nsew default output
rlabel metal4 s 63512 0 63588 212 4 dout0[14]
port 77 nsew default output
rlabel metal4 s 65960 0 66036 212 4 dout0[15]
port 76 nsew default output
rlabel metal4 s 68272 0 68348 212 4 dout0[16]
port 75 nsew default output
rlabel metal4 s 16048 0 16124 212 4 addr0[0]
port 41 nsew default input
rlabel metal4 s 17136 0 17212 212 4 addr0[1]
port 40 nsew default input
rlabel metal4 s 18224 0 18300 212 4 wmask0[0]
port 59 nsew default input
rlabel metal4 s 19584 0 19660 212 4 wmask0[1]
port 58 nsew default input
rlabel metal4 s 20536 0 20612 212 4 wmask0[2]
port 57 nsew default input
rlabel metal4 s 21760 0 21836 212 4 wmask0[3]
port 56 nsew default input
rlabel metal4 s 23120 0 23196 212 4 din0[0]
port 32 nsew default input
rlabel metal4 s 24208 0 24284 212 4 din0[1]
port 31 nsew default input
rlabel metal4 s 25432 0 25508 212 4 din0[2]
port 30 nsew default input
rlabel metal4 s 26520 0 26596 212 4 din0[3]
port 29 nsew default input
rlabel metal4 s 27608 0 27684 212 4 din0[4]
port 28 nsew default input
rlabel metal4 s 28696 0 28772 212 4 din0[5]
port 27 nsew default input
rlabel metal4 s 30056 0 30132 212 4 din0[6]
port 26 nsew default input
rlabel metal4 s 31280 0 31356 212 4 din0[7]
port 25 nsew default input
rlabel metal4 s 32368 0 32444 212 4 din0[8]
port 24 nsew default input
rlabel metal4 s 33456 0 33532 212 4 din0[9]
port 23 nsew default input
rlabel metal4 s 34544 0 34620 212 4 din0[10]
port 22 nsew default input
rlabel metal4 s 35904 0 35980 212 4 din0[11]
port 21 nsew default input
rlabel metal4 s 36992 0 37068 212 4 din0[12]
port 20 nsew default input
rlabel metal4 s 38080 0 38156 212 4 din0[13]
port 19 nsew default input
rlabel metal4 s 39440 0 39516 212 4 din0[14]
port 18 nsew default input
rlabel metal4 s 40664 0 40740 212 4 din0[15]
port 17 nsew default input
rlabel metal4 s 41752 0 41828 212 4 din0[16]
port 16 nsew default input
rlabel metal4 s 42840 0 42916 212 4 din0[17]
port 15 nsew default input
rlabel metal4 s 43928 0 44004 212 4 din0[18]
port 14 nsew default input
rlabel metal4 s 45288 0 45364 212 4 din0[19]
port 13 nsew default input
rlabel metal4 s 46376 0 46452 212 4 din0[20]
port 12 nsew default input
rlabel metal4 s 47600 0 47676 212 4 din0[21]
port 11 nsew default input
rlabel metal4 s 48688 0 48764 212 4 din0[22]
port 10 nsew default input
rlabel metal4 s 49776 0 49852 212 4 din0[23]
port 9 nsew default input
rlabel metal4 s 51136 0 51212 212 4 din0[24]
port 8 nsew default input
rlabel metal4 s 52224 0 52300 212 4 din0[25]
port 7 nsew default input
rlabel metal4 s 53312 0 53388 212 4 din0[26]
port 6 nsew default input
rlabel metal4 s 54400 0 54476 212 4 din0[27]
port 5 nsew default input
rlabel metal4 s 55760 0 55836 212 4 din0[28]
port 4 nsew default input
rlabel metal4 s 56984 0 57060 212 4 din0[29]
port 3 nsew default input
rlabel metal4 s 58072 0 58148 212 4 din0[30]
port 2 nsew default input
rlabel metal4 s 59160 0 59236 212 4 din0[31]
port 1 nsew default input
rlabel metal4 s 28288 0 28364 212 4 dout0[0]
port 91 nsew default output
rlabel metal4 s 30736 0 30812 212 4 dout0[1]
port 90 nsew default output
rlabel metal4 s 33592 0 33668 212 4 dout0[2]
port 89 nsew default output
rlabel metal4 s 952 952 1300 82356 4 vccd1
port 124 nsew power bidirectional abutment
rlabel metal4 s 272 272 620 83036 4 vssd1
port 125 nsew ground bidirectional abutment
rlabel metal4 s 103360 0 103436 212 4 dout0[30]
port 61 nsew default output
rlabel metal4 s 105944 0 106020 212 4 dout0[31]
port 60 nsew default output
rlabel metal4 s 70992 0 71068 212 4 dout0[17]
port 74 nsew default output
rlabel metal4 s 73440 0 73516 212 4 dout0[18]
port 73 nsew default output
rlabel metal4 s 75888 0 75964 212 4 dout0[19]
port 72 nsew default output
rlabel metal4 s 78472 0 78548 212 4 dout0[20]
port 71 nsew default output
rlabel metal4 s 80920 0 80996 212 4 dout0[21]
port 70 nsew default output
rlabel metal4 s 83504 0 83580 212 4 dout0[22]
port 69 nsew default output
rlabel metal4 s 85952 0 86028 212 4 dout0[23]
port 68 nsew default output
rlabel metal4 s 88536 0 88612 212 4 dout0[24]
port 67 nsew default output
rlabel metal4 s 90984 0 91060 212 4 dout0[25]
port 66 nsew default output
rlabel metal4 s 93432 0 93508 212 4 dout0[26]
port 65 nsew default output
rlabel metal4 s 95880 0 95956 212 4 dout0[27]
port 64 nsew default output
rlabel metal4 s 123216 0 123292 212 4 addr1[7]
port 43 nsew default input
rlabel metal4 s 123352 0 123428 212 4 addr1[8]
port 42 nsew default input
rlabel metal4 s 98464 0 98540 212 4 dout0[28]
port 63 nsew default output
rlabel metal4 s 135320 952 135668 82356 4 vccd1
port 124 nsew power bidirectional abutment
rlabel metal4 s 136000 272 136348 83036 4 vssd1
port 125 nsew ground bidirectional abutment
rlabel metal4 s 100912 0 100988 212 4 dout0[29]
port 62 nsew default output
<< properties >>
string FIXED_BBOX 0 0 136620 83308
string GDS_END 15213044
string GDS_FILE $PDKPATH/libs.ref/sky130_sram_macros/gds/sky130_sram_2kbyte_1rw1r_32x512_8.gds
string GDS_START 13196574
string LEFclass BLOCK
string LEFsymmetry X Y R90
<< end >>
